module basic_2500_25000_3000_5_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_2139,In_2478);
or U1 (N_1,In_329,In_1043);
xor U2 (N_2,In_1155,In_1976);
and U3 (N_3,In_1426,In_109);
nor U4 (N_4,In_1316,In_1248);
xnor U5 (N_5,In_2080,In_2346);
nor U6 (N_6,In_987,In_296);
nor U7 (N_7,In_2193,In_979);
nand U8 (N_8,In_390,In_357);
xnor U9 (N_9,In_980,In_1059);
nand U10 (N_10,In_153,In_1931);
or U11 (N_11,In_2076,In_2189);
nor U12 (N_12,In_2023,In_1821);
nor U13 (N_13,In_1932,In_1929);
or U14 (N_14,In_1991,In_1984);
nand U15 (N_15,In_1837,In_2200);
xor U16 (N_16,In_298,In_893);
xnor U17 (N_17,In_1681,In_2227);
or U18 (N_18,In_213,In_1975);
xnor U19 (N_19,In_185,In_2389);
and U20 (N_20,In_455,In_1690);
xor U21 (N_21,In_2220,In_1489);
and U22 (N_22,In_2349,In_2134);
nor U23 (N_23,In_1372,In_389);
and U24 (N_24,In_2020,In_2167);
and U25 (N_25,In_2415,In_2454);
nor U26 (N_26,In_741,In_70);
and U27 (N_27,In_281,In_355);
nor U28 (N_28,In_1635,In_302);
or U29 (N_29,In_328,In_396);
nor U30 (N_30,In_280,In_2051);
nand U31 (N_31,In_1729,In_1982);
and U32 (N_32,In_2041,In_1741);
or U33 (N_33,In_715,In_226);
and U34 (N_34,In_1742,In_1541);
or U35 (N_35,In_91,In_1539);
nor U36 (N_36,In_1421,In_1950);
xor U37 (N_37,In_1052,In_1567);
nand U38 (N_38,In_1503,In_2417);
or U39 (N_39,In_15,In_1359);
nor U40 (N_40,In_1985,In_1816);
nor U41 (N_41,In_1594,In_1619);
xnor U42 (N_42,In_1124,In_2018);
and U43 (N_43,In_1281,In_1679);
nand U44 (N_44,In_508,In_1517);
and U45 (N_45,In_1607,In_1666);
nor U46 (N_46,In_2197,In_519);
or U47 (N_47,In_1302,In_1630);
xnor U48 (N_48,In_850,In_2371);
nand U49 (N_49,In_598,In_362);
and U50 (N_50,In_1297,In_1417);
nor U51 (N_51,In_1076,In_2397);
xor U52 (N_52,In_76,In_452);
xnor U53 (N_53,In_2387,In_1069);
xor U54 (N_54,In_1363,In_2177);
or U55 (N_55,In_1809,In_648);
and U56 (N_56,In_545,In_251);
and U57 (N_57,In_1414,In_2121);
and U58 (N_58,In_2049,In_773);
or U59 (N_59,In_1538,In_1269);
nor U60 (N_60,In_748,In_1279);
nor U61 (N_61,In_29,In_1625);
nand U62 (N_62,In_1187,In_1340);
nor U63 (N_63,In_139,In_2317);
nand U64 (N_64,In_1788,In_166);
xor U65 (N_65,In_2108,In_1001);
nand U66 (N_66,In_607,In_1111);
xnor U67 (N_67,In_864,In_505);
or U68 (N_68,In_1531,In_44);
and U69 (N_69,In_899,In_399);
xor U70 (N_70,In_160,In_1331);
and U71 (N_71,In_54,In_616);
and U72 (N_72,In_2109,In_2077);
nor U73 (N_73,In_1728,In_241);
nand U74 (N_74,In_679,In_1794);
nand U75 (N_75,In_1475,In_2156);
xnor U76 (N_76,In_1587,In_564);
nor U77 (N_77,In_292,In_2323);
nand U78 (N_78,In_1257,In_1678);
xnor U79 (N_79,In_1899,In_591);
nand U80 (N_80,In_849,In_1156);
nor U81 (N_81,In_764,In_844);
xnor U82 (N_82,In_1448,In_1726);
nand U83 (N_83,In_1045,In_1926);
nand U84 (N_84,In_540,In_1874);
nand U85 (N_85,In_2033,In_2416);
and U86 (N_86,In_1940,In_2013);
or U87 (N_87,In_2101,In_1674);
nand U88 (N_88,In_1767,In_1467);
or U89 (N_89,In_1917,In_1776);
nand U90 (N_90,In_600,In_2017);
and U91 (N_91,In_919,In_413);
nor U92 (N_92,In_1849,In_1231);
or U93 (N_93,In_1171,In_141);
nor U94 (N_94,In_38,In_2026);
nor U95 (N_95,In_1575,In_82);
nor U96 (N_96,In_440,In_653);
nor U97 (N_97,In_22,In_1206);
and U98 (N_98,In_518,In_918);
nand U99 (N_99,In_2147,In_1751);
nand U100 (N_100,In_983,In_414);
or U101 (N_101,In_2246,In_1540);
and U102 (N_102,In_1096,In_633);
nand U103 (N_103,In_709,In_625);
and U104 (N_104,In_2363,In_96);
xor U105 (N_105,In_1165,In_1213);
and U106 (N_106,In_212,In_134);
or U107 (N_107,In_1964,In_632);
or U108 (N_108,In_1036,In_236);
or U109 (N_109,In_2123,In_841);
and U110 (N_110,In_894,In_1006);
nor U111 (N_111,In_1336,In_1164);
and U112 (N_112,In_194,In_1354);
nor U113 (N_113,In_675,In_1195);
nor U114 (N_114,In_579,In_187);
and U115 (N_115,In_1508,In_1110);
or U116 (N_116,In_766,In_1459);
xnor U117 (N_117,In_490,In_1157);
nand U118 (N_118,In_1119,In_668);
xnor U119 (N_119,In_780,In_2230);
or U120 (N_120,In_327,In_32);
xor U121 (N_121,In_813,In_1934);
xor U122 (N_122,In_2128,In_2178);
xor U123 (N_123,In_716,In_1677);
and U124 (N_124,In_963,In_925);
nand U125 (N_125,In_1659,In_808);
xnor U126 (N_126,In_201,In_1054);
nand U127 (N_127,In_1044,In_1038);
or U128 (N_128,In_1620,In_1115);
nor U129 (N_129,In_412,In_1709);
xor U130 (N_130,In_1974,In_199);
and U131 (N_131,In_9,In_101);
or U132 (N_132,In_288,In_1172);
or U133 (N_133,In_2199,In_311);
xor U134 (N_134,In_2437,In_868);
nand U135 (N_135,In_1662,In_278);
nor U136 (N_136,In_1647,In_496);
nand U137 (N_137,In_669,In_325);
and U138 (N_138,In_137,In_778);
nor U139 (N_139,In_1627,In_418);
xor U140 (N_140,In_1772,In_1324);
or U141 (N_141,In_2194,In_984);
and U142 (N_142,In_58,In_580);
or U143 (N_143,In_1078,In_1246);
nand U144 (N_144,In_1713,In_1745);
nand U145 (N_145,In_581,In_2324);
or U146 (N_146,In_1422,In_643);
nand U147 (N_147,In_996,In_2449);
or U148 (N_148,In_2262,In_936);
nor U149 (N_149,In_2340,In_811);
nor U150 (N_150,In_1273,In_95);
nand U151 (N_151,In_1787,In_1300);
nand U152 (N_152,In_334,In_2066);
xnor U153 (N_153,In_52,In_150);
or U154 (N_154,In_210,In_1261);
nand U155 (N_155,In_2241,In_1050);
nand U156 (N_156,In_1352,In_365);
nor U157 (N_157,In_363,In_1313);
or U158 (N_158,In_438,In_470);
xor U159 (N_159,In_1727,In_373);
or U160 (N_160,In_207,In_2245);
and U161 (N_161,In_2182,In_730);
or U162 (N_162,In_1074,In_1585);
xnor U163 (N_163,In_1186,In_842);
or U164 (N_164,In_477,In_1825);
nand U165 (N_165,In_2154,In_422);
or U166 (N_166,In_1371,In_970);
nand U167 (N_167,In_1838,In_164);
nand U168 (N_168,In_1801,In_295);
nand U169 (N_169,In_1218,In_1317);
and U170 (N_170,In_330,In_916);
or U171 (N_171,In_2451,In_2327);
or U172 (N_172,In_608,In_277);
xnor U173 (N_173,In_867,In_364);
and U174 (N_174,In_965,In_584);
nand U175 (N_175,In_2212,In_2420);
xor U176 (N_176,In_531,In_1335);
xnor U177 (N_177,In_2391,In_950);
nand U178 (N_178,In_624,In_1895);
nand U179 (N_179,In_548,In_907);
or U180 (N_180,In_1643,In_1373);
nor U181 (N_181,In_1958,In_1344);
nor U182 (N_182,In_2142,In_1210);
nand U183 (N_183,In_1428,In_1449);
nor U184 (N_184,In_416,In_588);
xor U185 (N_185,In_97,In_1460);
and U186 (N_186,In_771,In_1843);
and U187 (N_187,In_1031,In_1315);
nand U188 (N_188,In_1497,In_1131);
nand U189 (N_189,In_249,In_1379);
or U190 (N_190,In_886,In_1872);
nand U191 (N_191,In_276,In_2465);
or U192 (N_192,In_2224,In_1560);
nand U193 (N_193,In_806,In_1754);
or U194 (N_194,In_2221,In_2085);
xnor U195 (N_195,In_534,In_1628);
xnor U196 (N_196,In_1407,In_443);
and U197 (N_197,In_1536,In_989);
nand U198 (N_198,In_1008,In_1675);
nor U199 (N_199,In_246,In_1145);
nor U200 (N_200,In_180,In_721);
nor U201 (N_201,In_863,In_263);
xor U202 (N_202,In_1226,In_1040);
nand U203 (N_203,In_1477,In_673);
nor U204 (N_204,In_81,In_1798);
nand U205 (N_205,In_170,In_1887);
or U206 (N_206,In_130,In_1996);
or U207 (N_207,In_1660,In_1688);
or U208 (N_208,In_2072,In_1085);
and U209 (N_209,In_708,In_1683);
nor U210 (N_210,In_458,In_2052);
nand U211 (N_211,In_2028,In_410);
or U212 (N_212,In_374,In_1142);
nor U213 (N_213,In_2310,In_2119);
xor U214 (N_214,In_331,In_927);
and U215 (N_215,In_558,In_735);
nor U216 (N_216,In_234,In_66);
or U217 (N_217,In_1641,In_258);
nor U218 (N_218,In_2487,In_2097);
or U219 (N_219,In_734,In_2456);
nand U220 (N_220,In_2320,In_1533);
xnor U221 (N_221,In_94,In_441);
nand U222 (N_222,In_790,In_1135);
or U223 (N_223,In_1861,In_1309);
and U224 (N_224,In_428,In_2247);
nor U225 (N_225,In_2273,In_1463);
or U226 (N_226,In_1220,In_392);
xnor U227 (N_227,In_1377,In_468);
nand U228 (N_228,In_1270,In_369);
nand U229 (N_229,In_1446,In_400);
or U230 (N_230,In_1370,In_2486);
nand U231 (N_231,In_1584,In_2144);
nor U232 (N_232,In_1386,In_1480);
or U233 (N_233,In_1725,In_1501);
or U234 (N_234,In_1418,In_111);
xnor U235 (N_235,In_1733,In_831);
or U236 (N_236,In_1760,In_1307);
or U237 (N_237,In_1138,In_900);
nor U238 (N_238,In_812,In_2279);
nor U239 (N_239,In_656,In_905);
or U240 (N_240,In_2092,In_1884);
nor U241 (N_241,In_1048,In_1020);
nand U242 (N_242,In_2225,In_1438);
and U243 (N_243,In_1237,In_1254);
nand U244 (N_244,In_1440,In_2315);
or U245 (N_245,In_1267,In_1190);
or U246 (N_246,In_878,In_2057);
or U247 (N_247,In_1977,In_488);
nand U248 (N_248,In_1955,In_2396);
or U249 (N_249,In_1640,In_408);
or U250 (N_250,In_761,In_2412);
nor U251 (N_251,In_1437,In_404);
nand U252 (N_252,In_1482,In_1341);
nand U253 (N_253,In_717,In_421);
nor U254 (N_254,In_890,In_1384);
xnor U255 (N_255,In_682,In_1804);
nand U256 (N_256,In_239,In_1094);
nand U257 (N_257,In_1125,In_2024);
and U258 (N_258,In_1113,In_966);
xor U259 (N_259,In_2409,In_484);
nor U260 (N_260,In_274,In_286);
nor U261 (N_261,In_2118,In_1945);
or U262 (N_262,In_1841,In_462);
xor U263 (N_263,In_2325,In_1493);
or U264 (N_264,In_1399,In_2407);
nor U265 (N_265,In_1765,In_782);
nand U266 (N_266,In_1897,In_1972);
or U267 (N_267,In_924,In_1671);
and U268 (N_268,In_214,In_386);
xor U269 (N_269,In_1280,In_1935);
xor U270 (N_270,In_934,In_1944);
and U271 (N_271,In_2124,In_1579);
or U272 (N_272,In_1586,In_838);
xnor U273 (N_273,In_1290,In_7);
xnor U274 (N_274,In_1571,In_990);
nor U275 (N_275,In_1433,In_1104);
and U276 (N_276,In_2008,In_427);
or U277 (N_277,In_228,In_1060);
xnor U278 (N_278,In_1951,In_1966);
and U279 (N_279,In_1555,In_1092);
xnor U280 (N_280,In_1952,In_803);
and U281 (N_281,In_486,In_2330);
and U282 (N_282,In_2019,In_664);
nand U283 (N_283,In_1263,In_1021);
and U284 (N_284,In_937,In_2388);
and U285 (N_285,In_2381,In_2170);
nand U286 (N_286,In_1790,In_1087);
or U287 (N_287,In_2159,In_1238);
nor U288 (N_288,In_1349,In_393);
nor U289 (N_289,In_1920,In_127);
or U290 (N_290,In_1221,In_1327);
or U291 (N_291,In_74,In_1573);
nand U292 (N_292,In_459,In_999);
nand U293 (N_293,In_229,In_2140);
and U294 (N_294,In_662,In_2464);
nor U295 (N_295,In_1514,In_155);
xor U296 (N_296,In_426,In_480);
nor U297 (N_297,In_1667,In_420);
or U298 (N_298,In_2400,In_1707);
and U299 (N_299,In_1242,In_1163);
and U300 (N_300,In_1024,In_23);
and U301 (N_301,In_504,In_1922);
or U302 (N_302,In_401,In_405);
and U303 (N_303,In_382,In_2296);
xnor U304 (N_304,In_1906,In_2292);
xnor U305 (N_305,In_1046,In_1723);
xor U306 (N_306,In_435,In_2016);
nor U307 (N_307,In_2107,In_1326);
nor U308 (N_308,In_473,In_1771);
and U309 (N_309,In_498,In_941);
nand U310 (N_310,In_1240,In_2153);
and U311 (N_311,In_182,In_30);
nor U312 (N_312,In_884,In_1117);
xor U313 (N_313,In_169,In_825);
and U314 (N_314,In_1869,In_1432);
and U315 (N_315,In_2338,In_162);
and U316 (N_316,In_1227,In_342);
and U317 (N_317,In_1642,In_2260);
xnor U318 (N_318,In_1632,In_2459);
nor U319 (N_319,In_1605,In_1718);
and U320 (N_320,In_2267,In_2111);
nor U321 (N_321,In_751,In_528);
or U322 (N_322,In_354,In_492);
and U323 (N_323,In_259,In_1989);
nor U324 (N_324,In_1669,In_2091);
or U325 (N_325,In_1378,In_1484);
xor U326 (N_326,In_312,In_935);
nand U327 (N_327,In_1548,In_1894);
nor U328 (N_328,In_2335,In_221);
or U329 (N_329,In_931,In_644);
and U330 (N_330,In_2272,In_2084);
xor U331 (N_331,In_2264,In_1637);
or U332 (N_332,In_13,In_2138);
nand U333 (N_333,In_618,In_1805);
and U334 (N_334,In_196,In_407);
nor U335 (N_335,In_1737,In_2432);
or U336 (N_336,In_834,In_128);
nand U337 (N_337,In_1037,In_1470);
nor U338 (N_338,In_1409,In_163);
nand U339 (N_339,In_177,In_1782);
nand U340 (N_340,In_1530,In_2286);
nor U341 (N_341,In_2173,In_585);
nor U342 (N_342,In_2149,In_1488);
and U343 (N_343,In_674,In_240);
nor U344 (N_344,In_1562,In_513);
nor U345 (N_345,In_69,In_1106);
or U346 (N_346,In_1411,In_2314);
and U347 (N_347,In_2180,In_2425);
nand U348 (N_348,In_760,In_315);
or U349 (N_349,In_1056,In_1230);
nor U350 (N_350,In_2479,In_1457);
nor U351 (N_351,In_1916,In_772);
nor U352 (N_352,In_316,In_1763);
nand U353 (N_353,In_367,In_78);
nand U354 (N_354,In_2006,In_1905);
nor U355 (N_355,In_1262,In_1810);
xor U356 (N_356,In_2039,In_962);
xnor U357 (N_357,In_1986,In_2003);
or U358 (N_358,In_1464,In_807);
or U359 (N_359,In_2453,In_1755);
xor U360 (N_360,In_1051,In_879);
and U361 (N_361,In_2222,In_123);
nor U362 (N_362,In_2129,In_107);
nor U363 (N_363,In_1553,In_1880);
and U364 (N_364,In_1694,In_1631);
xor U365 (N_365,In_1817,In_339);
nand U366 (N_366,In_2448,In_1746);
xor U367 (N_367,In_2166,In_1717);
nor U368 (N_368,In_2086,In_1902);
or U369 (N_369,In_324,In_793);
nor U370 (N_370,In_467,In_1346);
and U371 (N_371,In_2214,In_1287);
xnor U372 (N_372,In_872,In_634);
and U373 (N_373,In_113,In_1770);
or U374 (N_374,In_1987,In_769);
nand U375 (N_375,In_1918,In_171);
xor U376 (N_376,In_1852,In_1615);
xnor U377 (N_377,In_220,In_1235);
and U378 (N_378,In_911,In_2047);
or U379 (N_379,In_809,In_2468);
or U380 (N_380,In_2263,In_1970);
or U381 (N_381,In_307,In_2036);
or U382 (N_382,In_657,In_725);
nor U383 (N_383,In_881,In_1842);
and U384 (N_384,In_1779,In_745);
xor U385 (N_385,In_507,In_297);
nor U386 (N_386,In_1042,In_739);
and U387 (N_387,In_1853,In_1193);
and U388 (N_388,In_695,In_1939);
nor U389 (N_389,In_969,In_713);
nand U390 (N_390,In_1919,In_85);
nor U391 (N_391,In_1668,In_1173);
xor U392 (N_392,In_1703,In_1212);
xnor U393 (N_393,In_1004,In_2361);
nand U394 (N_394,In_60,In_1786);
or U395 (N_395,In_1222,In_2205);
nand U396 (N_396,In_2010,In_1732);
or U397 (N_397,In_1828,In_757);
and U398 (N_398,In_1812,In_1967);
or U399 (N_399,In_1784,In_1785);
xor U400 (N_400,In_117,In_1522);
xor U401 (N_401,In_720,In_2476);
nor U402 (N_402,In_1581,In_6);
nand U403 (N_403,In_1547,In_2460);
nor U404 (N_404,In_124,In_1600);
nand U405 (N_405,In_703,In_2383);
nand U406 (N_406,In_1864,In_902);
nand U407 (N_407,In_112,In_854);
xor U408 (N_408,In_1780,In_1552);
and U409 (N_409,In_437,In_1469);
or U410 (N_410,In_291,In_1130);
and U411 (N_411,In_345,In_1695);
nand U412 (N_412,In_2424,In_2127);
nor U413 (N_413,In_2204,In_882);
nor U414 (N_414,In_711,In_906);
xor U415 (N_415,In_1799,In_2334);
nor U416 (N_416,In_843,In_230);
xnor U417 (N_417,In_1147,In_1323);
nand U418 (N_418,In_34,In_753);
and U419 (N_419,In_2283,In_1293);
and U420 (N_420,In_686,In_603);
or U421 (N_421,In_1266,In_651);
nand U422 (N_422,In_71,In_897);
xnor U423 (N_423,In_1258,In_756);
nand U424 (N_424,In_1132,In_2137);
nor U425 (N_425,In_1698,In_1198);
xor U426 (N_426,In_948,In_541);
nor U427 (N_427,In_179,In_572);
xor U428 (N_428,In_1978,In_895);
nand U429 (N_429,In_1330,In_216);
xor U430 (N_430,In_2494,In_671);
and U431 (N_431,In_2427,In_1445);
xnor U432 (N_432,In_2444,In_197);
nor U433 (N_433,In_789,In_2196);
and U434 (N_434,In_1829,In_2257);
or U435 (N_435,In_816,In_219);
and U436 (N_436,In_944,In_1364);
and U437 (N_437,In_235,In_57);
and U438 (N_438,In_566,In_1570);
or U439 (N_439,In_1822,In_2073);
xor U440 (N_440,In_660,In_1353);
nor U441 (N_441,In_544,In_1768);
nand U442 (N_442,In_105,In_2005);
xnor U443 (N_443,In_961,In_2302);
and U444 (N_444,In_784,In_231);
xnor U445 (N_445,In_289,In_442);
and U446 (N_446,In_1879,In_1007);
and U447 (N_447,In_306,In_173);
nand U448 (N_448,In_181,In_2288);
nor U449 (N_449,In_1891,In_300);
nor U450 (N_450,In_133,In_2443);
xnor U451 (N_451,In_2115,In_55);
nand U452 (N_452,In_1356,In_1516);
and U453 (N_453,In_1913,In_1844);
or U454 (N_454,In_1088,In_659);
nor U455 (N_455,In_1830,In_810);
and U456 (N_456,In_1093,In_515);
nor U457 (N_457,In_2089,In_1609);
and U458 (N_458,In_1528,In_99);
nor U459 (N_459,In_2390,In_1680);
nand U460 (N_460,In_209,In_1833);
nand U461 (N_461,In_1365,In_218);
xor U462 (N_462,In_1938,In_1590);
and U463 (N_463,In_143,In_158);
nand U464 (N_464,In_104,In_2278);
nor U465 (N_465,In_1299,In_463);
or U466 (N_466,In_1696,In_1691);
or U467 (N_467,In_140,In_1604);
nor U468 (N_468,In_2467,In_146);
nand U469 (N_469,In_1526,In_1022);
xor U470 (N_470,In_178,In_2291);
xnor U471 (N_471,In_1965,In_862);
and U472 (N_472,In_430,In_1710);
nand U473 (N_473,In_2295,In_747);
or U474 (N_474,In_2440,In_285);
nand U475 (N_475,In_1188,In_1520);
nor U476 (N_476,In_953,In_1818);
or U477 (N_477,In_244,In_1298);
or U478 (N_478,In_349,In_2305);
nand U479 (N_479,In_20,In_445);
nor U480 (N_480,In_2113,In_1606);
nor U481 (N_481,In_1578,In_2228);
nor U482 (N_482,In_304,In_2254);
xnor U483 (N_483,In_2452,In_204);
and U484 (N_484,In_1256,In_942);
nor U485 (N_485,In_1721,In_904);
or U486 (N_486,In_1439,In_2011);
and U487 (N_487,In_685,In_1140);
xnor U488 (N_488,In_1646,In_977);
or U489 (N_489,In_972,In_707);
xnor U490 (N_490,In_1182,In_471);
nor U491 (N_491,In_2054,In_1260);
and U492 (N_492,In_704,In_690);
nor U493 (N_493,In_2117,In_447);
or U494 (N_494,In_1223,In_1152);
nand U495 (N_495,In_631,In_1170);
xnor U496 (N_496,In_1629,In_1835);
or U497 (N_497,In_2174,In_1394);
nor U498 (N_498,In_1018,In_2007);
nand U499 (N_499,In_661,In_619);
xnor U500 (N_500,In_1761,In_1191);
and U501 (N_501,In_2438,In_947);
xor U502 (N_502,In_142,In_89);
and U503 (N_503,In_265,In_2014);
nand U504 (N_504,In_1211,In_652);
xor U505 (N_505,In_2164,In_2234);
or U506 (N_506,In_1101,In_2293);
and U507 (N_507,In_1375,In_946);
nor U508 (N_508,In_2053,In_1968);
nor U509 (N_509,In_824,In_1345);
nand U510 (N_510,In_1391,In_2242);
xnor U511 (N_511,In_2143,In_1143);
nor U512 (N_512,In_1648,In_2069);
nand U513 (N_513,In_1652,In_1988);
nand U514 (N_514,In_595,In_1062);
nand U515 (N_515,In_387,In_594);
xor U516 (N_516,In_2000,In_543);
and U517 (N_517,In_243,In_1963);
nor U518 (N_518,In_411,In_250);
and U519 (N_519,In_264,In_847);
nand U520 (N_520,In_2031,In_2360);
or U521 (N_521,In_1362,In_723);
nor U522 (N_522,In_2368,In_1228);
and U523 (N_523,In_1388,In_797);
nor U524 (N_524,In_2282,In_1347);
and U525 (N_525,In_1351,In_956);
or U526 (N_526,In_865,In_860);
nor U527 (N_527,In_320,In_1025);
nand U528 (N_528,In_955,In_1930);
and U529 (N_529,In_1750,In_2386);
nor U530 (N_530,In_176,In_2301);
or U531 (N_531,In_1283,In_1591);
or U532 (N_532,In_837,In_379);
xor U533 (N_533,In_2105,In_1275);
xnor U534 (N_534,In_424,In_875);
xor U535 (N_535,In_2233,In_976);
and U536 (N_536,In_1413,In_2074);
and U537 (N_537,In_1937,In_1824);
and U538 (N_538,In_1731,In_2252);
nand U539 (N_539,In_910,In_487);
and U540 (N_540,In_1355,In_303);
xnor U541 (N_541,In_2369,In_26);
nor U542 (N_542,In_1491,In_2044);
nand U543 (N_543,In_620,In_2078);
nand U544 (N_544,In_1102,In_1908);
xnor U545 (N_545,In_958,In_2378);
xor U546 (N_546,In_1781,In_2419);
or U547 (N_547,In_136,In_823);
nor U548 (N_548,In_2110,In_28);
nand U549 (N_549,In_1314,In_1715);
nor U550 (N_550,In_2308,In_2489);
xor U551 (N_551,In_586,In_260);
xnor U552 (N_552,In_982,In_1724);
xor U553 (N_553,In_1176,In_602);
xnor U554 (N_554,In_398,In_290);
or U555 (N_555,In_1689,In_1003);
and U556 (N_556,In_444,In_2068);
or U557 (N_557,In_475,In_1881);
or U558 (N_558,In_1487,In_859);
xnor U559 (N_559,In_1486,In_1942);
xor U560 (N_560,In_2075,In_1811);
and U561 (N_561,In_2155,In_189);
xnor U562 (N_562,In_2294,In_2152);
nand U563 (N_563,In_2484,In_2151);
nand U564 (N_564,In_1736,In_755);
or U565 (N_565,In_1960,In_2056);
xnor U566 (N_566,In_1588,In_195);
and U567 (N_567,In_2326,In_1333);
nor U568 (N_568,In_370,In_2219);
or U569 (N_569,In_1049,In_2211);
or U570 (N_570,In_1443,In_336);
nor U571 (N_571,In_1285,In_1095);
nand U572 (N_572,In_2087,In_397);
or U573 (N_573,In_2195,In_768);
nor U574 (N_574,In_2483,In_795);
or U575 (N_575,In_604,In_663);
and U576 (N_576,In_681,In_1622);
nor U577 (N_577,In_506,In_1306);
and U578 (N_578,In_434,In_192);
and U579 (N_579,In_350,In_1959);
or U580 (N_580,In_1507,In_1582);
and U581 (N_581,In_469,In_2354);
or U582 (N_582,In_521,In_2269);
or U583 (N_583,In_2112,In_1200);
or U584 (N_584,In_232,In_2165);
or U585 (N_585,In_729,In_2015);
or U586 (N_586,In_25,In_1803);
nand U587 (N_587,In_1807,In_1626);
xor U588 (N_588,In_2004,In_483);
xor U589 (N_589,In_871,In_777);
nor U590 (N_590,In_606,In_495);
nand U591 (N_591,In_317,In_2481);
nor U592 (N_592,In_2012,In_375);
nor U593 (N_593,In_1232,In_1867);
nand U594 (N_594,In_887,In_856);
nand U595 (N_595,In_658,In_630);
nor U596 (N_596,In_1969,In_1397);
or U597 (N_597,In_891,In_967);
or U598 (N_598,In_348,In_481);
nand U599 (N_599,In_568,In_1903);
xnor U600 (N_600,In_929,In_338);
xnor U601 (N_601,In_949,In_1483);
nor U602 (N_602,In_1856,In_131);
nor U603 (N_603,In_43,In_1057);
or U604 (N_604,In_640,In_1550);
and U605 (N_605,In_2090,In_1866);
nor U606 (N_606,In_1616,In_932);
or U607 (N_607,In_2318,In_322);
nand U608 (N_608,In_2380,In_2457);
nor U609 (N_609,In_2032,In_2116);
nor U610 (N_610,In_2331,In_2353);
nand U611 (N_611,In_489,In_1009);
or U612 (N_612,In_2098,In_590);
nand U613 (N_613,In_2034,In_72);
nand U614 (N_614,In_256,In_47);
xor U615 (N_615,In_1465,In_943);
nor U616 (N_616,In_2265,In_1367);
or U617 (N_617,In_913,In_1239);
or U618 (N_618,In_2046,In_1105);
and U619 (N_619,In_1682,In_1368);
nor U620 (N_620,In_565,In_273);
xnor U621 (N_621,In_570,In_356);
nor U622 (N_622,In_326,In_1328);
or U623 (N_623,In_378,In_1342);
or U624 (N_624,In_2307,In_524);
nand U625 (N_625,In_1686,In_2062);
and U626 (N_626,In_1740,In_2198);
nor U627 (N_627,In_262,In_2403);
or U628 (N_628,In_1308,In_1793);
nor U629 (N_629,In_994,In_2215);
xnor U630 (N_630,In_63,In_986);
nand U631 (N_631,In_641,In_1091);
nand U632 (N_632,In_1183,In_1034);
nand U633 (N_633,In_493,In_1137);
or U634 (N_634,In_945,In_1554);
xnor U635 (N_635,In_2497,In_346);
xnor U636 (N_636,In_1204,In_1035);
or U637 (N_637,In_959,In_2207);
nor U638 (N_638,In_1914,In_605);
and U639 (N_639,In_952,In_542);
xnor U640 (N_640,In_1845,In_2402);
and U641 (N_641,In_451,In_840);
xor U642 (N_642,In_978,In_2237);
and U643 (N_643,In_2306,In_1312);
and U644 (N_644,In_1318,In_2063);
or U645 (N_645,In_79,In_233);
xor U646 (N_646,In_1129,In_402);
and U647 (N_647,In_1196,In_100);
nor U648 (N_648,In_429,In_49);
nor U649 (N_649,In_649,In_1215);
nor U650 (N_650,In_688,In_1948);
nand U651 (N_651,In_1311,In_2045);
or U652 (N_652,In_926,In_2048);
nand U653 (N_653,In_914,In_1080);
xnor U654 (N_654,In_1542,In_559);
xor U655 (N_655,In_1524,In_2002);
or U656 (N_656,In_2188,In_861);
and U657 (N_657,In_1081,In_833);
nand U658 (N_658,In_1181,In_2406);
xor U659 (N_659,In_525,In_1099);
nor U660 (N_660,In_1334,In_538);
or U661 (N_661,In_1265,In_885);
xor U662 (N_662,In_2040,In_1995);
xnor U663 (N_663,In_1272,In_2);
nand U664 (N_664,In_815,In_1454);
nand U665 (N_665,In_676,In_750);
nand U666 (N_666,In_1700,In_787);
nand U667 (N_667,In_68,In_1225);
nand U668 (N_668,In_1769,In_549);
nor U669 (N_669,In_1893,In_805);
or U670 (N_670,In_762,In_746);
or U671 (N_671,In_737,In_988);
and U672 (N_672,In_973,In_1015);
or U673 (N_673,In_388,In_257);
and U674 (N_674,In_1079,In_67);
nand U675 (N_675,In_376,In_165);
or U676 (N_676,In_642,In_2037);
nor U677 (N_677,In_83,In_449);
nand U678 (N_678,In_0,In_1764);
and U679 (N_679,In_796,In_2300);
nand U680 (N_680,In_377,In_1158);
and U681 (N_681,In_2488,In_1067);
nand U682 (N_682,In_1634,In_2358);
or U683 (N_683,In_476,In_2431);
and U684 (N_684,In_1572,In_270);
nand U685 (N_685,In_1992,In_2093);
nand U686 (N_686,In_1244,In_1055);
nand U687 (N_687,In_2256,In_2103);
and U688 (N_688,In_271,In_964);
or U689 (N_689,In_655,In_1203);
or U690 (N_690,In_1858,In_2060);
xnor U691 (N_691,In_1650,In_61);
or U692 (N_692,In_722,In_1747);
xnor U693 (N_693,In_1883,In_995);
or U694 (N_694,In_2379,In_752);
nor U695 (N_695,In_1655,In_1241);
nand U696 (N_696,In_1017,In_147);
or U697 (N_697,In_215,In_1462);
and U698 (N_698,In_17,In_512);
and U699 (N_699,In_1556,In_2255);
nand U700 (N_700,In_612,In_1332);
xnor U701 (N_701,In_1148,In_188);
nand U702 (N_702,In_39,In_2482);
nand U703 (N_703,In_479,In_208);
or U704 (N_704,In_1954,In_2133);
xor U705 (N_705,In_678,In_557);
nand U706 (N_706,In_2364,In_1608);
and U707 (N_707,In_37,In_1656);
nor U708 (N_708,In_56,In_1633);
or U709 (N_709,In_2405,In_770);
nand U710 (N_710,In_759,In_1126);
nor U711 (N_711,In_2439,In_1150);
nand U712 (N_712,In_670,In_125);
nand U713 (N_713,In_1286,In_1180);
nand U714 (N_714,In_1875,In_2284);
and U715 (N_715,In_200,In_1603);
nor U716 (N_716,In_2359,In_1112);
nand U717 (N_717,In_1070,In_1673);
nor U718 (N_718,In_2146,In_692);
nand U719 (N_719,In_184,In_516);
and U720 (N_720,In_1670,In_997);
xor U721 (N_721,In_2226,In_203);
nor U722 (N_722,In_1398,In_1403);
or U723 (N_723,In_1502,In_2329);
nand U724 (N_724,In_1613,In_59);
nor U725 (N_725,In_1014,In_951);
nand U726 (N_726,In_1301,In_1128);
or U727 (N_727,In_1019,In_1453);
xor U728 (N_728,In_193,In_1521);
and U729 (N_729,In_2393,In_647);
or U730 (N_730,In_960,In_2352);
and U731 (N_731,In_2434,In_2462);
nand U732 (N_732,In_705,In_998);
and U733 (N_733,In_857,In_2009);
xnor U734 (N_734,In_940,In_792);
xnor U735 (N_735,In_774,In_1013);
and U736 (N_736,In_930,In_744);
or U737 (N_737,In_1162,In_877);
and U738 (N_738,In_2064,In_1481);
nand U739 (N_739,In_578,In_436);
xor U740 (N_740,In_546,In_2235);
nand U741 (N_741,In_2067,In_174);
or U742 (N_742,In_1946,In_1744);
xnor U743 (N_743,In_1645,In_1002);
and U744 (N_744,In_2304,In_2435);
and U745 (N_745,In_1161,In_503);
xnor U746 (N_746,In_992,In_1473);
nor U747 (N_747,In_217,In_1383);
nand U748 (N_748,In_1294,In_1990);
nor U749 (N_749,In_2471,In_3);
and U750 (N_750,In_1278,In_2100);
nor U751 (N_751,In_464,In_1205);
xor U752 (N_752,In_126,In_1855);
xor U753 (N_753,In_1510,In_1012);
or U754 (N_754,In_2176,In_2271);
nand U755 (N_755,In_380,In_132);
nor U756 (N_756,In_1458,In_2270);
or U757 (N_757,In_425,In_2382);
xor U758 (N_758,In_491,In_1596);
xnor U759 (N_759,In_801,In_2030);
and U760 (N_760,In_120,In_1292);
and U761 (N_761,In_1146,In_1123);
and U762 (N_762,In_2372,In_1826);
xor U763 (N_763,In_1819,In_332);
nand U764 (N_764,In_874,In_115);
nand U765 (N_765,In_573,In_2258);
nand U766 (N_766,In_1924,In_1395);
or U767 (N_767,In_1592,In_2160);
xor U768 (N_768,In_19,In_2042);
nor U769 (N_769,In_1429,In_1361);
xnor U770 (N_770,In_1083,In_1610);
and U771 (N_771,In_2442,In_2251);
or U772 (N_772,In_1077,In_1452);
nor U773 (N_773,In_2374,In_1863);
nor U774 (N_774,In_1425,In_2399);
nor U775 (N_775,In_623,In_2001);
and U776 (N_776,In_2367,In_383);
or U777 (N_777,In_21,In_1358);
nor U778 (N_778,In_1719,In_754);
nand U779 (N_779,In_636,In_1159);
nand U780 (N_780,In_1406,In_2277);
xnor U781 (N_781,In_45,In_321);
nor U782 (N_782,In_2059,In_245);
nor U783 (N_783,In_650,In_1597);
nor U784 (N_784,In_614,In_1276);
or U785 (N_785,In_791,In_2083);
and U786 (N_786,In_917,In_175);
or U787 (N_787,In_372,In_145);
or U788 (N_788,In_1400,In_149);
nor U789 (N_789,In_726,In_2395);
nor U790 (N_790,In_522,In_921);
or U791 (N_791,In_1589,In_876);
and U792 (N_792,In_223,In_2122);
or U793 (N_793,In_2385,In_1243);
xnor U794 (N_794,In_2275,In_563);
nor U795 (N_795,In_1624,In_991);
or U796 (N_796,In_2190,In_1498);
and U797 (N_797,In_1907,In_1513);
nor U798 (N_798,In_1569,In_119);
nand U799 (N_799,In_1350,In_2473);
nand U800 (N_800,In_560,In_283);
and U801 (N_801,In_2365,In_2218);
xor U802 (N_802,In_2357,In_1886);
nor U803 (N_803,In_702,In_108);
nor U804 (N_804,In_1033,In_2287);
nor U805 (N_805,In_1178,In_2096);
nand U806 (N_806,In_928,In_98);
xor U807 (N_807,In_1427,In_2299);
xor U808 (N_808,In_880,In_1901);
nand U809 (N_809,In_1133,In_2447);
nor U810 (N_810,In_1168,In_159);
or U811 (N_811,In_1757,In_198);
nand U812 (N_812,In_1039,In_1927);
and U813 (N_813,In_1325,In_1820);
nand U814 (N_814,In_2081,In_873);
nor U815 (N_815,In_1369,In_1665);
nand U816 (N_816,In_2421,In_2070);
xor U817 (N_817,In_714,In_2313);
nand U818 (N_818,In_2025,In_2203);
xor U819 (N_819,In_587,In_224);
nor U820 (N_820,In_1925,In_394);
nor U821 (N_821,In_1154,In_2297);
xnor U822 (N_822,In_2191,In_2311);
xnor U823 (N_823,In_775,In_1525);
nor U824 (N_824,In_1618,In_1971);
nor U825 (N_825,In_1752,In_2206);
or U826 (N_826,In_2470,In_2192);
or U827 (N_827,In_836,In_2210);
nand U828 (N_828,In_2351,In_706);
nand U829 (N_829,In_665,In_1028);
or U830 (N_830,In_822,In_1144);
nor U831 (N_831,In_361,In_2309);
and U832 (N_832,In_933,In_1865);
xnor U833 (N_833,In_1860,In_2082);
and U834 (N_834,In_1072,In_939);
nor U835 (N_835,In_482,In_275);
nand U836 (N_836,In_896,In_553);
nand U837 (N_837,In_1,In_1026);
or U838 (N_838,In_2341,In_46);
nand U839 (N_839,In_1456,In_892);
xnor U840 (N_840,In_2418,In_1499);
nand U841 (N_841,In_1684,In_1234);
and U842 (N_842,In_1169,In_1544);
and U843 (N_843,In_1549,In_2474);
nor U844 (N_844,In_333,In_1382);
or U845 (N_845,In_1716,In_501);
nand U846 (N_846,In_1068,In_1663);
or U847 (N_847,In_2375,In_1797);
nand U848 (N_848,In_853,In_2079);
and U849 (N_849,In_971,In_1202);
nor U850 (N_850,In_719,In_2333);
nand U851 (N_851,In_282,In_1871);
xor U852 (N_852,In_687,In_1509);
or U853 (N_853,In_1756,In_1360);
nor U854 (N_854,In_319,In_798);
xor U855 (N_855,In_1233,In_2135);
nand U856 (N_856,In_1563,In_1796);
nand U857 (N_857,In_1442,In_118);
nor U858 (N_858,In_1697,In_2239);
nand U859 (N_859,In_1831,In_2150);
and U860 (N_860,In_611,In_1167);
and U861 (N_861,In_156,In_2336);
nor U862 (N_862,In_1847,In_80);
and U863 (N_863,In_691,In_1743);
or U864 (N_864,In_415,In_1599);
nor U865 (N_865,In_786,In_2186);
and U866 (N_866,In_314,In_183);
or U867 (N_867,In_728,In_2414);
nand U868 (N_868,In_1441,In_536);
xnor U869 (N_869,In_1846,In_1711);
xor U870 (N_870,In_1357,In_2343);
nor U871 (N_871,In_733,In_2021);
or U872 (N_872,In_583,In_1274);
or U873 (N_873,In_1073,In_31);
xnor U874 (N_874,In_2071,In_1380);
nor U875 (N_875,In_2274,In_1904);
and U876 (N_876,In_2430,In_1532);
xor U877 (N_877,In_335,In_222);
or U878 (N_878,In_1778,In_294);
nor U879 (N_879,In_152,In_2332);
nand U880 (N_880,In_308,In_1506);
or U881 (N_881,In_1217,In_1374);
and U882 (N_882,In_654,In_1184);
nand U883 (N_883,In_2319,In_718);
nand U884 (N_884,In_385,In_151);
nand U885 (N_885,In_1827,In_12);
and U886 (N_886,In_1107,In_852);
and U887 (N_887,In_869,In_2495);
and U888 (N_888,In_2172,In_359);
or U889 (N_889,In_2130,In_1153);
nand U890 (N_890,In_1151,In_2285);
or U891 (N_891,In_106,In_1166);
nand U892 (N_892,In_116,In_1348);
nand U893 (N_893,In_571,In_2163);
or U894 (N_894,In_299,In_1199);
and U895 (N_895,In_2475,In_2342);
nand U896 (N_896,In_1461,In_1623);
xnor U897 (N_897,In_2038,In_547);
nand U898 (N_898,In_2175,In_954);
nand U899 (N_899,In_1577,In_1496);
or U900 (N_900,In_2493,In_1762);
nand U901 (N_901,In_2376,In_2229);
or U902 (N_902,In_2384,In_48);
and U903 (N_903,In_1999,In_968);
nand U904 (N_904,In_638,In_1702);
xor U905 (N_905,In_1450,In_1023);
nand U906 (N_906,In_1941,In_86);
nand U907 (N_907,In_510,In_1565);
and U908 (N_908,In_1505,In_261);
xor U909 (N_909,In_2355,In_1415);
nor U910 (N_910,In_2248,In_2347);
or U911 (N_911,In_617,In_1823);
xor U912 (N_912,In_1949,In_62);
nor U913 (N_913,In_597,In_736);
xor U914 (N_914,In_144,In_2428);
xnor U915 (N_915,In_526,In_353);
xnor U916 (N_916,In_779,In_1065);
or U917 (N_917,In_293,In_1114);
xor U918 (N_918,In_1714,In_2102);
xor U919 (N_919,In_938,In_2433);
nor U920 (N_920,In_238,In_698);
xnor U921 (N_921,In_35,In_1121);
and U922 (N_922,In_1758,In_2466);
xnor U923 (N_923,In_90,In_1583);
xnor U924 (N_924,In_697,In_1699);
or U925 (N_925,In_1047,In_1639);
nor U926 (N_926,In_1479,In_1504);
xor U927 (N_927,In_1259,In_1981);
nor U928 (N_928,In_237,In_689);
xnor U929 (N_929,In_1192,In_211);
or U930 (N_930,In_2125,In_2104);
xor U931 (N_931,In_626,In_2094);
and U932 (N_932,In_1515,In_1338);
and U933 (N_933,In_2120,In_2250);
nand U934 (N_934,In_432,In_1424);
and U935 (N_935,In_1685,In_1179);
and U936 (N_936,In_1649,In_1288);
and U937 (N_937,In_2145,In_511);
nor U938 (N_938,In_1561,In_1160);
nor U939 (N_939,In_1854,In_765);
xnor U940 (N_940,In_763,In_1512);
nand U941 (N_941,In_446,In_1947);
nand U942 (N_942,In_627,In_817);
and U943 (N_943,In_738,In_2148);
and U944 (N_944,In_1490,In_1434);
and U945 (N_945,In_1997,In_448);
nand U946 (N_946,In_1071,In_1289);
nor U947 (N_947,In_1430,In_2058);
nand U948 (N_948,In_1574,In_465);
or U949 (N_949,In_802,In_8);
nor U950 (N_950,In_539,In_2171);
and U951 (N_951,In_1658,In_776);
xor U952 (N_952,In_2131,In_1749);
or U953 (N_953,In_1953,In_1617);
xnor U954 (N_954,In_1687,In_310);
nor U955 (N_955,In_1936,In_253);
or U956 (N_956,In_2168,In_248);
and U957 (N_957,In_1268,In_993);
xor U958 (N_958,In_567,In_785);
nor U959 (N_959,In_1255,In_73);
or U960 (N_960,In_2446,In_1759);
or U961 (N_961,In_1896,In_1892);
xnor U962 (N_962,In_2463,In_2411);
and U963 (N_963,In_1264,In_1973);
xnor U964 (N_964,In_1519,In_1738);
nor U965 (N_965,In_1664,In_191);
or U966 (N_966,In_358,In_1010);
and U967 (N_967,In_788,In_922);
and U968 (N_968,In_1410,In_2298);
xor U969 (N_969,In_1814,In_268);
or U970 (N_970,In_1580,In_1075);
xor U971 (N_971,In_42,In_1385);
or U972 (N_972,In_269,In_533);
and U973 (N_973,In_1928,In_1730);
and U974 (N_974,In_637,In_1834);
xor U975 (N_975,In_114,In_2126);
and U976 (N_976,In_2348,In_724);
nand U977 (N_977,In_1122,In_2209);
or U978 (N_978,In_819,In_2472);
nand U979 (N_979,In_1109,In_381);
nand U980 (N_980,In_1053,In_301);
nor U981 (N_981,In_2217,In_1097);
xnor U982 (N_982,In_2027,In_157);
and U983 (N_983,In_323,In_360);
nand U984 (N_984,In_40,In_818);
and U985 (N_985,In_1636,In_2423);
nand U986 (N_986,In_1813,In_2088);
or U987 (N_987,In_2268,In_431);
nand U988 (N_988,In_2480,In_186);
xnor U989 (N_989,In_347,In_2339);
or U990 (N_990,In_1612,In_677);
or U991 (N_991,In_1802,In_1839);
nand U992 (N_992,In_2249,In_14);
and U993 (N_993,In_981,In_2398);
nand U994 (N_994,In_1923,In_1284);
or U995 (N_995,In_732,In_318);
and U996 (N_996,In_252,In_148);
and U997 (N_997,In_2029,In_1108);
nand U998 (N_998,In_1295,In_1189);
xnor U999 (N_999,In_11,In_1857);
nand U1000 (N_1000,In_1495,In_1621);
nor U1001 (N_1001,In_254,In_1310);
nor U1002 (N_1002,In_2259,In_1910);
xor U1003 (N_1003,In_1478,In_609);
nor U1004 (N_1004,In_1706,In_1993);
and U1005 (N_1005,In_2141,In_1319);
xnor U1006 (N_1006,In_1175,In_514);
xor U1007 (N_1007,In_103,In_1800);
or U1008 (N_1008,In_1576,In_693);
and U1009 (N_1009,In_577,In_1149);
xnor U1010 (N_1010,In_1773,In_523);
or U1011 (N_1011,In_1753,In_749);
and U1012 (N_1012,In_227,In_1090);
or U1013 (N_1013,In_161,In_1141);
or U1014 (N_1014,In_2232,In_1127);
nor U1015 (N_1015,In_1451,In_352);
nor U1016 (N_1016,In_1082,In_1708);
nand U1017 (N_1017,In_2394,In_371);
xnor U1018 (N_1018,In_135,In_2445);
nor U1019 (N_1019,In_1601,In_2161);
and U1020 (N_1020,In_1529,In_2208);
or U1021 (N_1021,In_450,In_1748);
nand U1022 (N_1022,In_574,In_93);
and U1023 (N_1023,In_1888,In_615);
nor U1024 (N_1024,In_2499,In_1651);
nor U1025 (N_1025,In_497,In_1543);
or U1026 (N_1026,In_1405,In_53);
xor U1027 (N_1027,In_2184,In_888);
nand U1028 (N_1028,In_1253,In_384);
or U1029 (N_1029,In_2169,In_731);
nand U1030 (N_1030,In_1247,In_821);
or U1031 (N_1031,In_1868,In_1389);
nand U1032 (N_1032,In_1654,In_92);
xor U1033 (N_1033,In_1224,In_2410);
or U1034 (N_1034,In_1089,In_1134);
or U1035 (N_1035,In_242,In_2490);
nand U1036 (N_1036,In_1568,In_2312);
and U1037 (N_1037,In_2213,In_1396);
and U1038 (N_1038,In_2187,In_2181);
nand U1039 (N_1039,In_1657,In_599);
nand U1040 (N_1040,In_460,In_1873);
nand U1041 (N_1041,In_77,In_202);
nand U1042 (N_1042,In_2132,In_832);
nand U1043 (N_1043,In_839,In_596);
nand U1044 (N_1044,In_206,In_439);
and U1045 (N_1045,In_255,In_457);
nand U1046 (N_1046,In_622,In_2345);
xor U1047 (N_1047,In_575,In_1197);
nor U1048 (N_1048,In_1420,In_1029);
nor U1049 (N_1049,In_1661,In_576);
xnor U1050 (N_1050,In_313,In_461);
nand U1051 (N_1051,In_1890,In_1271);
nor U1052 (N_1052,In_2289,In_1909);
nor U1053 (N_1053,In_1511,In_1956);
and U1054 (N_1054,In_474,In_667);
nand U1055 (N_1055,In_1174,In_2422);
nor U1056 (N_1056,In_2458,In_1774);
and U1057 (N_1057,In_423,In_24);
nor U1058 (N_1058,In_167,In_1392);
and U1059 (N_1059,In_1214,In_121);
nor U1060 (N_1060,In_672,In_102);
and U1061 (N_1061,In_1320,In_2095);
nand U1062 (N_1062,In_1889,In_499);
nor U1063 (N_1063,In_18,In_2106);
xnor U1064 (N_1064,In_2158,In_2231);
nand U1065 (N_1065,In_1840,In_1564);
nor U1066 (N_1066,In_1030,In_1870);
or U1067 (N_1067,In_41,In_829);
nor U1068 (N_1068,In_1139,In_64);
nand U1069 (N_1069,In_1208,In_2266);
or U1070 (N_1070,In_1712,In_889);
nor U1071 (N_1071,In_846,In_800);
nand U1072 (N_1072,In_1722,In_1957);
nand U1073 (N_1073,In_1321,In_2261);
xnor U1074 (N_1074,In_1832,In_138);
xor U1075 (N_1075,In_1466,In_2162);
or U1076 (N_1076,In_2392,In_247);
nor U1077 (N_1077,In_2350,In_110);
xor U1078 (N_1078,In_456,In_1943);
xor U1079 (N_1079,In_1474,In_1229);
xor U1080 (N_1080,In_908,In_2436);
and U1081 (N_1081,In_1701,In_1878);
or U1082 (N_1082,In_1704,In_975);
nand U1083 (N_1083,In_550,In_1494);
nor U1084 (N_1084,In_1252,In_517);
and U1085 (N_1085,In_1084,In_767);
and U1086 (N_1086,In_1322,In_2404);
nor U1087 (N_1087,In_340,In_835);
and U1088 (N_1088,In_696,In_845);
or U1089 (N_1089,In_1296,In_1016);
and U1090 (N_1090,In_1791,In_1766);
xnor U1091 (N_1091,In_903,In_1518);
and U1092 (N_1092,In_828,In_1401);
nand U1093 (N_1093,In_646,In_1245);
and U1094 (N_1094,In_1216,In_305);
nor U1095 (N_1095,In_1103,In_1476);
nand U1096 (N_1096,In_2179,In_1980);
nor U1097 (N_1097,In_1118,In_2322);
xor U1098 (N_1098,In_27,In_168);
or U1099 (N_1099,In_409,In_1795);
or U1100 (N_1100,In_1994,In_1404);
nand U1101 (N_1101,In_1559,In_84);
nand U1102 (N_1102,In_1933,In_1557);
xnor U1103 (N_1103,In_898,In_454);
xor U1104 (N_1104,In_1032,In_500);
nor U1105 (N_1105,In_2485,In_1381);
nor U1106 (N_1106,In_2202,In_1546);
nor U1107 (N_1107,In_2238,In_406);
or U1108 (N_1108,In_1376,In_2099);
nor U1109 (N_1109,In_2496,In_50);
xor U1110 (N_1110,In_1792,In_2280);
nand U1111 (N_1111,In_1282,In_1366);
nand U1112 (N_1112,In_225,In_1815);
nand U1113 (N_1113,In_1468,In_16);
xor U1114 (N_1114,In_1066,In_883);
xor U1115 (N_1115,In_2362,In_1593);
nand U1116 (N_1116,In_551,In_2240);
and U1117 (N_1117,In_2344,In_870);
and U1118 (N_1118,In_561,In_1595);
and U1119 (N_1119,In_701,In_915);
nor U1120 (N_1120,In_1915,In_1602);
nand U1121 (N_1121,In_1177,In_2183);
nor U1122 (N_1122,In_743,In_2216);
nand U1123 (N_1123,In_2461,In_368);
nor U1124 (N_1124,In_1250,In_266);
or U1125 (N_1125,In_2236,In_552);
and U1126 (N_1126,In_582,In_1412);
nor U1127 (N_1127,In_520,In_1061);
xnor U1128 (N_1128,In_830,In_1862);
nor U1129 (N_1129,In_1882,In_799);
and U1130 (N_1130,In_1291,In_556);
nor U1131 (N_1131,In_1249,In_1912);
xor U1132 (N_1132,In_2065,In_529);
nand U1133 (N_1133,In_1402,In_1911);
nand U1134 (N_1134,In_827,In_2243);
nand U1135 (N_1135,In_851,In_2316);
or U1136 (N_1136,In_1739,In_712);
or U1137 (N_1137,In_727,In_635);
nand U1138 (N_1138,In_1611,In_639);
nand U1139 (N_1139,In_190,In_2366);
and U1140 (N_1140,In_2201,In_629);
nand U1141 (N_1141,In_1735,In_1431);
or U1142 (N_1142,In_2303,In_742);
nand U1143 (N_1143,In_344,In_569);
nand U1144 (N_1144,In_494,In_88);
or U1145 (N_1145,In_645,In_2055);
nand U1146 (N_1146,In_1063,In_1116);
nor U1147 (N_1147,In_1447,In_172);
or U1148 (N_1148,In_2253,In_1207);
nand U1149 (N_1149,In_1435,In_2244);
xor U1150 (N_1150,In_87,In_453);
or U1151 (N_1151,In_272,In_2373);
or U1152 (N_1152,In_309,In_1219);
or U1153 (N_1153,In_343,In_610);
nor U1154 (N_1154,In_1236,In_820);
nand U1155 (N_1155,In_1100,In_2223);
or U1156 (N_1156,In_51,In_1551);
or U1157 (N_1157,In_1598,In_1343);
and U1158 (N_1158,In_527,In_1775);
and U1159 (N_1159,In_2491,In_1472);
nor U1160 (N_1160,In_36,In_2337);
nand U1161 (N_1161,In_555,In_781);
nand U1162 (N_1162,In_122,In_1638);
and U1163 (N_1163,In_804,In_1979);
nor U1164 (N_1164,In_284,In_1303);
and U1165 (N_1165,In_1339,In_2426);
nand U1166 (N_1166,In_2043,In_472);
xnor U1167 (N_1167,In_694,In_920);
and U1168 (N_1168,In_1492,In_593);
xor U1169 (N_1169,In_985,In_1777);
nand U1170 (N_1170,In_1848,In_2185);
nand U1171 (N_1171,In_1455,In_1921);
nor U1172 (N_1172,In_1734,In_509);
nand U1173 (N_1173,In_814,In_1720);
or U1174 (N_1174,In_909,In_1500);
or U1175 (N_1175,In_1789,In_419);
nor U1176 (N_1176,In_2114,In_1416);
and U1177 (N_1177,In_2290,In_1120);
and U1178 (N_1178,In_1672,In_783);
or U1179 (N_1179,In_351,In_1851);
nand U1180 (N_1180,In_601,In_403);
xor U1181 (N_1181,In_1387,In_974);
nor U1182 (N_1182,In_1653,In_2035);
xor U1183 (N_1183,In_740,In_1998);
xor U1184 (N_1184,In_2328,In_2492);
nor U1185 (N_1185,In_2050,In_758);
nand U1186 (N_1186,In_1329,In_2413);
and U1187 (N_1187,In_855,In_485);
and U1188 (N_1188,In_5,In_2441);
xor U1189 (N_1189,In_537,In_589);
xor U1190 (N_1190,In_433,In_1277);
xnor U1191 (N_1191,In_1423,In_65);
nor U1192 (N_1192,In_1537,In_10);
xnor U1193 (N_1193,In_337,In_1534);
or U1194 (N_1194,In_2450,In_1558);
nand U1195 (N_1195,In_2136,In_33);
nand U1196 (N_1196,In_1041,In_1644);
nand U1197 (N_1197,In_2061,In_1305);
xnor U1198 (N_1198,In_2370,In_267);
and U1199 (N_1199,In_466,In_1444);
and U1200 (N_1200,In_613,In_532);
and U1201 (N_1201,In_2429,In_1185);
nor U1202 (N_1202,In_1471,In_2498);
nand U1203 (N_1203,In_478,In_1876);
nand U1204 (N_1204,In_848,In_699);
nand U1205 (N_1205,In_1408,In_1885);
or U1206 (N_1206,In_923,In_1859);
xnor U1207 (N_1207,In_1251,In_1614);
or U1208 (N_1208,In_1393,In_279);
or U1209 (N_1209,In_957,In_562);
nor U1210 (N_1210,In_1304,In_1058);
nand U1211 (N_1211,In_341,In_1194);
and U1212 (N_1212,In_1676,In_1808);
nand U1213 (N_1213,In_683,In_554);
or U1214 (N_1214,In_2477,In_1485);
nor U1215 (N_1215,In_1064,In_1419);
and U1216 (N_1216,In_417,In_1877);
and U1217 (N_1217,In_1705,In_1011);
nor U1218 (N_1218,In_1961,In_1962);
or U1219 (N_1219,In_1983,In_395);
or U1220 (N_1220,In_1692,In_1027);
nor U1221 (N_1221,In_826,In_621);
and U1222 (N_1222,In_912,In_1806);
xor U1223 (N_1223,In_1136,In_530);
or U1224 (N_1224,In_1000,In_2321);
and U1225 (N_1225,In_700,In_628);
and U1226 (N_1226,In_1337,In_666);
nand U1227 (N_1227,In_1783,In_75);
or U1228 (N_1228,In_1566,In_1693);
or U1229 (N_1229,In_2469,In_2281);
nor U1230 (N_1230,In_901,In_2455);
nor U1231 (N_1231,In_1900,In_684);
and U1232 (N_1232,In_1436,In_535);
or U1233 (N_1233,In_1898,In_2401);
and U1234 (N_1234,In_858,In_680);
and U1235 (N_1235,In_1086,In_1005);
nand U1236 (N_1236,In_592,In_391);
xor U1237 (N_1237,In_502,In_866);
xnor U1238 (N_1238,In_129,In_1535);
xor U1239 (N_1239,In_710,In_1390);
nand U1240 (N_1240,In_1527,In_2022);
xnor U1241 (N_1241,In_205,In_1523);
nor U1242 (N_1242,In_1209,In_2157);
nor U1243 (N_1243,In_2408,In_1836);
and U1244 (N_1244,In_794,In_154);
or U1245 (N_1245,In_2377,In_287);
xor U1246 (N_1246,In_1201,In_1098);
xor U1247 (N_1247,In_1545,In_2276);
nand U1248 (N_1248,In_2356,In_4);
nand U1249 (N_1249,In_1850,In_366);
nand U1250 (N_1250,In_562,In_1733);
nor U1251 (N_1251,In_46,In_1837);
and U1252 (N_1252,In_1440,In_2136);
or U1253 (N_1253,In_13,In_253);
xor U1254 (N_1254,In_1853,In_2458);
xor U1255 (N_1255,In_113,In_841);
nand U1256 (N_1256,In_1994,In_918);
nor U1257 (N_1257,In_93,In_591);
nor U1258 (N_1258,In_1416,In_616);
or U1259 (N_1259,In_965,In_391);
nor U1260 (N_1260,In_1182,In_996);
xor U1261 (N_1261,In_1221,In_1020);
and U1262 (N_1262,In_1259,In_765);
nor U1263 (N_1263,In_763,In_799);
and U1264 (N_1264,In_936,In_737);
and U1265 (N_1265,In_357,In_2018);
and U1266 (N_1266,In_240,In_704);
and U1267 (N_1267,In_1557,In_2398);
nand U1268 (N_1268,In_1815,In_2238);
or U1269 (N_1269,In_1737,In_739);
nor U1270 (N_1270,In_94,In_2060);
and U1271 (N_1271,In_2207,In_22);
nor U1272 (N_1272,In_619,In_1892);
and U1273 (N_1273,In_2042,In_468);
or U1274 (N_1274,In_780,In_449);
xor U1275 (N_1275,In_2315,In_577);
xor U1276 (N_1276,In_2350,In_2285);
nor U1277 (N_1277,In_2228,In_21);
nand U1278 (N_1278,In_638,In_989);
nor U1279 (N_1279,In_567,In_1758);
nor U1280 (N_1280,In_1340,In_400);
nor U1281 (N_1281,In_771,In_2161);
xor U1282 (N_1282,In_2074,In_18);
or U1283 (N_1283,In_844,In_1769);
and U1284 (N_1284,In_2308,In_1589);
and U1285 (N_1285,In_1185,In_1927);
nor U1286 (N_1286,In_325,In_502);
xnor U1287 (N_1287,In_2113,In_857);
or U1288 (N_1288,In_1718,In_12);
or U1289 (N_1289,In_1743,In_1519);
and U1290 (N_1290,In_2350,In_1128);
nand U1291 (N_1291,In_2421,In_244);
or U1292 (N_1292,In_838,In_1974);
or U1293 (N_1293,In_1058,In_1660);
and U1294 (N_1294,In_2013,In_2057);
or U1295 (N_1295,In_1539,In_2319);
and U1296 (N_1296,In_1535,In_2289);
nor U1297 (N_1297,In_1096,In_2150);
nand U1298 (N_1298,In_354,In_999);
and U1299 (N_1299,In_1106,In_979);
nor U1300 (N_1300,In_264,In_2310);
nand U1301 (N_1301,In_1485,In_1578);
or U1302 (N_1302,In_1517,In_742);
nor U1303 (N_1303,In_1861,In_1282);
xor U1304 (N_1304,In_490,In_1413);
nand U1305 (N_1305,In_719,In_514);
and U1306 (N_1306,In_475,In_265);
xor U1307 (N_1307,In_1441,In_1408);
and U1308 (N_1308,In_174,In_2278);
or U1309 (N_1309,In_824,In_1583);
and U1310 (N_1310,In_1224,In_731);
and U1311 (N_1311,In_317,In_654);
nand U1312 (N_1312,In_1232,In_209);
xnor U1313 (N_1313,In_2159,In_1779);
or U1314 (N_1314,In_1946,In_1805);
and U1315 (N_1315,In_2396,In_981);
and U1316 (N_1316,In_1442,In_1846);
and U1317 (N_1317,In_2413,In_214);
nor U1318 (N_1318,In_486,In_1120);
nor U1319 (N_1319,In_255,In_1141);
or U1320 (N_1320,In_2178,In_1917);
or U1321 (N_1321,In_1139,In_956);
xor U1322 (N_1322,In_1202,In_560);
and U1323 (N_1323,In_1697,In_990);
nor U1324 (N_1324,In_1348,In_2385);
xnor U1325 (N_1325,In_1099,In_2335);
xnor U1326 (N_1326,In_679,In_681);
or U1327 (N_1327,In_318,In_1956);
and U1328 (N_1328,In_795,In_1286);
nor U1329 (N_1329,In_1518,In_471);
xnor U1330 (N_1330,In_16,In_755);
xnor U1331 (N_1331,In_2392,In_1840);
or U1332 (N_1332,In_2441,In_1506);
xnor U1333 (N_1333,In_768,In_24);
or U1334 (N_1334,In_1354,In_1355);
xnor U1335 (N_1335,In_2122,In_715);
nand U1336 (N_1336,In_526,In_493);
nor U1337 (N_1337,In_2381,In_2353);
xnor U1338 (N_1338,In_2022,In_181);
and U1339 (N_1339,In_2391,In_259);
xnor U1340 (N_1340,In_550,In_1061);
xnor U1341 (N_1341,In_32,In_2181);
nand U1342 (N_1342,In_541,In_2257);
nor U1343 (N_1343,In_971,In_183);
xor U1344 (N_1344,In_2450,In_197);
nor U1345 (N_1345,In_2213,In_262);
and U1346 (N_1346,In_1108,In_1801);
nor U1347 (N_1347,In_1280,In_2368);
or U1348 (N_1348,In_374,In_1189);
or U1349 (N_1349,In_784,In_658);
and U1350 (N_1350,In_1205,In_1138);
or U1351 (N_1351,In_21,In_2053);
or U1352 (N_1352,In_1927,In_2237);
and U1353 (N_1353,In_903,In_436);
or U1354 (N_1354,In_653,In_1826);
or U1355 (N_1355,In_243,In_1862);
nand U1356 (N_1356,In_1889,In_2328);
xor U1357 (N_1357,In_1632,In_1265);
nor U1358 (N_1358,In_2093,In_1722);
and U1359 (N_1359,In_1079,In_134);
and U1360 (N_1360,In_1316,In_1104);
or U1361 (N_1361,In_1690,In_2030);
nand U1362 (N_1362,In_1242,In_458);
nand U1363 (N_1363,In_1687,In_715);
or U1364 (N_1364,In_192,In_1288);
nand U1365 (N_1365,In_2268,In_557);
xnor U1366 (N_1366,In_422,In_2162);
nor U1367 (N_1367,In_1044,In_998);
nand U1368 (N_1368,In_2201,In_1514);
nand U1369 (N_1369,In_688,In_1909);
xnor U1370 (N_1370,In_536,In_361);
or U1371 (N_1371,In_1885,In_2220);
and U1372 (N_1372,In_1383,In_1819);
xor U1373 (N_1373,In_1883,In_1628);
nand U1374 (N_1374,In_793,In_1988);
and U1375 (N_1375,In_1621,In_1384);
nand U1376 (N_1376,In_565,In_358);
xnor U1377 (N_1377,In_789,In_1153);
nand U1378 (N_1378,In_1647,In_1662);
nand U1379 (N_1379,In_1725,In_1494);
and U1380 (N_1380,In_641,In_1748);
and U1381 (N_1381,In_959,In_1709);
nand U1382 (N_1382,In_2449,In_600);
and U1383 (N_1383,In_1758,In_1271);
nor U1384 (N_1384,In_1215,In_1184);
nand U1385 (N_1385,In_2381,In_2313);
or U1386 (N_1386,In_525,In_231);
and U1387 (N_1387,In_2446,In_1868);
nand U1388 (N_1388,In_1172,In_98);
nand U1389 (N_1389,In_2201,In_134);
or U1390 (N_1390,In_1529,In_76);
or U1391 (N_1391,In_660,In_31);
xor U1392 (N_1392,In_1432,In_389);
xnor U1393 (N_1393,In_928,In_370);
xor U1394 (N_1394,In_2115,In_1126);
nor U1395 (N_1395,In_1368,In_385);
or U1396 (N_1396,In_2347,In_1266);
and U1397 (N_1397,In_2291,In_142);
xor U1398 (N_1398,In_14,In_1781);
nand U1399 (N_1399,In_693,In_2096);
nand U1400 (N_1400,In_713,In_2093);
nand U1401 (N_1401,In_1261,In_1336);
xnor U1402 (N_1402,In_974,In_1052);
nor U1403 (N_1403,In_267,In_2409);
nand U1404 (N_1404,In_387,In_436);
nor U1405 (N_1405,In_1749,In_2133);
and U1406 (N_1406,In_731,In_2300);
and U1407 (N_1407,In_290,In_1729);
or U1408 (N_1408,In_1850,In_1924);
nor U1409 (N_1409,In_1831,In_671);
nor U1410 (N_1410,In_1007,In_1365);
nor U1411 (N_1411,In_1556,In_2208);
and U1412 (N_1412,In_1886,In_150);
and U1413 (N_1413,In_2199,In_1173);
xor U1414 (N_1414,In_2077,In_1779);
nor U1415 (N_1415,In_75,In_904);
and U1416 (N_1416,In_1942,In_370);
xnor U1417 (N_1417,In_1960,In_2461);
and U1418 (N_1418,In_1535,In_1588);
nand U1419 (N_1419,In_965,In_1768);
nor U1420 (N_1420,In_1523,In_298);
nor U1421 (N_1421,In_798,In_2189);
nand U1422 (N_1422,In_370,In_1204);
nand U1423 (N_1423,In_858,In_2224);
nor U1424 (N_1424,In_2446,In_846);
nor U1425 (N_1425,In_1283,In_458);
xor U1426 (N_1426,In_2189,In_583);
nor U1427 (N_1427,In_1745,In_1306);
nor U1428 (N_1428,In_2103,In_2398);
and U1429 (N_1429,In_787,In_1886);
and U1430 (N_1430,In_1866,In_1873);
and U1431 (N_1431,In_182,In_2237);
xor U1432 (N_1432,In_1275,In_991);
nand U1433 (N_1433,In_775,In_1200);
nand U1434 (N_1434,In_1477,In_289);
nand U1435 (N_1435,In_2044,In_1258);
nand U1436 (N_1436,In_2455,In_2471);
nor U1437 (N_1437,In_523,In_2284);
xor U1438 (N_1438,In_2145,In_1099);
or U1439 (N_1439,In_1195,In_184);
xnor U1440 (N_1440,In_1328,In_353);
nor U1441 (N_1441,In_2416,In_1701);
and U1442 (N_1442,In_1124,In_1663);
nor U1443 (N_1443,In_951,In_1808);
and U1444 (N_1444,In_1695,In_837);
and U1445 (N_1445,In_2413,In_1192);
nand U1446 (N_1446,In_1883,In_2491);
nand U1447 (N_1447,In_950,In_2065);
or U1448 (N_1448,In_1222,In_273);
and U1449 (N_1449,In_985,In_1926);
or U1450 (N_1450,In_2135,In_1146);
nor U1451 (N_1451,In_1275,In_1107);
or U1452 (N_1452,In_2150,In_1334);
and U1453 (N_1453,In_2075,In_959);
nor U1454 (N_1454,In_941,In_1905);
nand U1455 (N_1455,In_229,In_2258);
and U1456 (N_1456,In_97,In_692);
xnor U1457 (N_1457,In_952,In_1499);
and U1458 (N_1458,In_500,In_2282);
nor U1459 (N_1459,In_827,In_1671);
nand U1460 (N_1460,In_2211,In_572);
and U1461 (N_1461,In_460,In_877);
nor U1462 (N_1462,In_2358,In_2297);
xnor U1463 (N_1463,In_2259,In_249);
xnor U1464 (N_1464,In_26,In_336);
nor U1465 (N_1465,In_342,In_508);
nand U1466 (N_1466,In_1471,In_17);
xor U1467 (N_1467,In_237,In_959);
nand U1468 (N_1468,In_172,In_766);
and U1469 (N_1469,In_343,In_2203);
nand U1470 (N_1470,In_1986,In_1066);
nand U1471 (N_1471,In_347,In_3);
or U1472 (N_1472,In_1310,In_943);
and U1473 (N_1473,In_131,In_994);
and U1474 (N_1474,In_2303,In_734);
and U1475 (N_1475,In_2201,In_2439);
nor U1476 (N_1476,In_2488,In_409);
nor U1477 (N_1477,In_1265,In_2374);
nand U1478 (N_1478,In_1822,In_176);
nand U1479 (N_1479,In_1123,In_39);
or U1480 (N_1480,In_2014,In_487);
nand U1481 (N_1481,In_275,In_601);
nand U1482 (N_1482,In_2075,In_143);
xor U1483 (N_1483,In_2289,In_1848);
or U1484 (N_1484,In_766,In_1907);
nor U1485 (N_1485,In_1176,In_462);
nand U1486 (N_1486,In_924,In_1125);
xnor U1487 (N_1487,In_408,In_2003);
nand U1488 (N_1488,In_2026,In_981);
and U1489 (N_1489,In_129,In_349);
nand U1490 (N_1490,In_1222,In_672);
and U1491 (N_1491,In_295,In_432);
nor U1492 (N_1492,In_1881,In_1259);
nor U1493 (N_1493,In_1267,In_1737);
nand U1494 (N_1494,In_331,In_1779);
xor U1495 (N_1495,In_2023,In_478);
and U1496 (N_1496,In_1123,In_1790);
or U1497 (N_1497,In_2233,In_304);
and U1498 (N_1498,In_1787,In_263);
and U1499 (N_1499,In_768,In_1310);
nor U1500 (N_1500,In_1598,In_1211);
or U1501 (N_1501,In_889,In_1578);
nor U1502 (N_1502,In_81,In_2185);
xnor U1503 (N_1503,In_492,In_787);
nor U1504 (N_1504,In_2156,In_799);
or U1505 (N_1505,In_2052,In_254);
or U1506 (N_1506,In_217,In_1110);
and U1507 (N_1507,In_2029,In_1057);
nand U1508 (N_1508,In_221,In_2318);
nor U1509 (N_1509,In_469,In_885);
nand U1510 (N_1510,In_1290,In_976);
or U1511 (N_1511,In_2195,In_1291);
nand U1512 (N_1512,In_2070,In_1862);
xnor U1513 (N_1513,In_2209,In_1946);
xor U1514 (N_1514,In_2146,In_940);
or U1515 (N_1515,In_1500,In_2273);
or U1516 (N_1516,In_1840,In_552);
nor U1517 (N_1517,In_151,In_1703);
and U1518 (N_1518,In_378,In_2390);
nand U1519 (N_1519,In_1050,In_1230);
nor U1520 (N_1520,In_324,In_1516);
nand U1521 (N_1521,In_477,In_510);
xor U1522 (N_1522,In_2397,In_604);
nor U1523 (N_1523,In_2448,In_2104);
nand U1524 (N_1524,In_2226,In_1258);
and U1525 (N_1525,In_2465,In_898);
nand U1526 (N_1526,In_2390,In_1283);
xnor U1527 (N_1527,In_1438,In_519);
nor U1528 (N_1528,In_1557,In_1304);
nor U1529 (N_1529,In_1391,In_2333);
or U1530 (N_1530,In_1530,In_912);
nor U1531 (N_1531,In_720,In_2341);
nor U1532 (N_1532,In_2484,In_786);
nor U1533 (N_1533,In_916,In_2246);
or U1534 (N_1534,In_1412,In_432);
nor U1535 (N_1535,In_464,In_1686);
and U1536 (N_1536,In_2148,In_1527);
nand U1537 (N_1537,In_1953,In_2048);
nor U1538 (N_1538,In_2402,In_2038);
nor U1539 (N_1539,In_1898,In_2140);
nand U1540 (N_1540,In_1497,In_1725);
nor U1541 (N_1541,In_739,In_115);
or U1542 (N_1542,In_2009,In_1714);
xnor U1543 (N_1543,In_533,In_1506);
xnor U1544 (N_1544,In_678,In_723);
and U1545 (N_1545,In_1139,In_410);
xor U1546 (N_1546,In_2382,In_836);
xnor U1547 (N_1547,In_833,In_276);
nand U1548 (N_1548,In_1896,In_1040);
nor U1549 (N_1549,In_128,In_2185);
nand U1550 (N_1550,In_111,In_1526);
nor U1551 (N_1551,In_1223,In_2057);
or U1552 (N_1552,In_1745,In_2047);
or U1553 (N_1553,In_74,In_758);
xor U1554 (N_1554,In_1785,In_626);
and U1555 (N_1555,In_1781,In_210);
nor U1556 (N_1556,In_678,In_1025);
or U1557 (N_1557,In_1600,In_1395);
nor U1558 (N_1558,In_1451,In_1745);
xnor U1559 (N_1559,In_555,In_340);
nor U1560 (N_1560,In_742,In_1848);
nand U1561 (N_1561,In_274,In_109);
nor U1562 (N_1562,In_2329,In_119);
and U1563 (N_1563,In_1472,In_1116);
and U1564 (N_1564,In_2012,In_817);
or U1565 (N_1565,In_2497,In_2370);
nand U1566 (N_1566,In_1861,In_709);
xnor U1567 (N_1567,In_1309,In_2073);
nor U1568 (N_1568,In_1740,In_111);
nand U1569 (N_1569,In_1900,In_1570);
xnor U1570 (N_1570,In_2190,In_2224);
or U1571 (N_1571,In_522,In_19);
xnor U1572 (N_1572,In_303,In_1836);
nand U1573 (N_1573,In_1289,In_1762);
xnor U1574 (N_1574,In_2381,In_1310);
and U1575 (N_1575,In_586,In_2446);
nor U1576 (N_1576,In_2392,In_780);
nand U1577 (N_1577,In_2228,In_1472);
nor U1578 (N_1578,In_1664,In_754);
nor U1579 (N_1579,In_342,In_1110);
xnor U1580 (N_1580,In_755,In_1818);
nor U1581 (N_1581,In_5,In_1521);
nor U1582 (N_1582,In_958,In_389);
and U1583 (N_1583,In_1157,In_1801);
nand U1584 (N_1584,In_729,In_2023);
or U1585 (N_1585,In_1186,In_194);
and U1586 (N_1586,In_2242,In_2450);
nand U1587 (N_1587,In_1117,In_991);
and U1588 (N_1588,In_291,In_950);
and U1589 (N_1589,In_620,In_2322);
and U1590 (N_1590,In_2040,In_1745);
or U1591 (N_1591,In_2220,In_2165);
xnor U1592 (N_1592,In_779,In_1327);
or U1593 (N_1593,In_1731,In_1282);
and U1594 (N_1594,In_787,In_497);
xor U1595 (N_1595,In_746,In_2172);
and U1596 (N_1596,In_1715,In_2001);
nor U1597 (N_1597,In_716,In_1643);
nor U1598 (N_1598,In_1342,In_762);
nor U1599 (N_1599,In_2365,In_445);
nand U1600 (N_1600,In_1180,In_2116);
xnor U1601 (N_1601,In_1187,In_139);
and U1602 (N_1602,In_2355,In_969);
and U1603 (N_1603,In_1125,In_1273);
nor U1604 (N_1604,In_399,In_1961);
nor U1605 (N_1605,In_945,In_589);
nand U1606 (N_1606,In_2242,In_875);
and U1607 (N_1607,In_1569,In_2214);
nor U1608 (N_1608,In_1271,In_999);
xor U1609 (N_1609,In_1479,In_846);
or U1610 (N_1610,In_778,In_782);
nand U1611 (N_1611,In_918,In_848);
nand U1612 (N_1612,In_1284,In_1333);
or U1613 (N_1613,In_2112,In_1021);
nor U1614 (N_1614,In_1473,In_345);
nand U1615 (N_1615,In_1682,In_411);
nand U1616 (N_1616,In_1519,In_645);
or U1617 (N_1617,In_2222,In_494);
nor U1618 (N_1618,In_424,In_413);
and U1619 (N_1619,In_1306,In_313);
or U1620 (N_1620,In_2476,In_1616);
nor U1621 (N_1621,In_427,In_444);
xnor U1622 (N_1622,In_1008,In_1480);
nor U1623 (N_1623,In_395,In_2389);
and U1624 (N_1624,In_1131,In_244);
xor U1625 (N_1625,In_1388,In_947);
xor U1626 (N_1626,In_939,In_1430);
or U1627 (N_1627,In_1948,In_1731);
or U1628 (N_1628,In_80,In_2023);
or U1629 (N_1629,In_1064,In_2362);
and U1630 (N_1630,In_313,In_1271);
nand U1631 (N_1631,In_308,In_627);
nand U1632 (N_1632,In_2031,In_497);
nand U1633 (N_1633,In_2455,In_1550);
and U1634 (N_1634,In_1408,In_2049);
nor U1635 (N_1635,In_1983,In_2432);
nand U1636 (N_1636,In_666,In_631);
nand U1637 (N_1637,In_2128,In_2211);
nor U1638 (N_1638,In_379,In_522);
xnor U1639 (N_1639,In_825,In_321);
or U1640 (N_1640,In_1110,In_2111);
nand U1641 (N_1641,In_904,In_949);
and U1642 (N_1642,In_1872,In_1531);
or U1643 (N_1643,In_2130,In_12);
and U1644 (N_1644,In_2092,In_2282);
and U1645 (N_1645,In_55,In_2321);
nand U1646 (N_1646,In_569,In_862);
and U1647 (N_1647,In_1715,In_1246);
nand U1648 (N_1648,In_2160,In_1575);
nand U1649 (N_1649,In_303,In_1172);
nand U1650 (N_1650,In_1492,In_2461);
xnor U1651 (N_1651,In_2373,In_2212);
xnor U1652 (N_1652,In_1259,In_1651);
xnor U1653 (N_1653,In_843,In_2198);
nor U1654 (N_1654,In_1371,In_2484);
xnor U1655 (N_1655,In_1039,In_2460);
and U1656 (N_1656,In_986,In_1994);
xnor U1657 (N_1657,In_950,In_1013);
nor U1658 (N_1658,In_137,In_2309);
xor U1659 (N_1659,In_720,In_2142);
and U1660 (N_1660,In_179,In_1473);
xnor U1661 (N_1661,In_2157,In_1113);
nand U1662 (N_1662,In_810,In_1360);
nand U1663 (N_1663,In_1224,In_2033);
nor U1664 (N_1664,In_384,In_1331);
xor U1665 (N_1665,In_399,In_2297);
or U1666 (N_1666,In_1932,In_719);
nor U1667 (N_1667,In_2060,In_344);
or U1668 (N_1668,In_2276,In_858);
and U1669 (N_1669,In_226,In_2473);
or U1670 (N_1670,In_1863,In_237);
nor U1671 (N_1671,In_1344,In_78);
nor U1672 (N_1672,In_384,In_2324);
and U1673 (N_1673,In_834,In_1786);
xnor U1674 (N_1674,In_70,In_1827);
xor U1675 (N_1675,In_186,In_1730);
xnor U1676 (N_1676,In_681,In_1334);
nand U1677 (N_1677,In_1041,In_2329);
nor U1678 (N_1678,In_440,In_292);
and U1679 (N_1679,In_1166,In_657);
xnor U1680 (N_1680,In_2110,In_746);
or U1681 (N_1681,In_2477,In_814);
nand U1682 (N_1682,In_54,In_925);
or U1683 (N_1683,In_1910,In_1615);
nor U1684 (N_1684,In_580,In_560);
nor U1685 (N_1685,In_12,In_1994);
nor U1686 (N_1686,In_1545,In_1074);
xor U1687 (N_1687,In_243,In_461);
xor U1688 (N_1688,In_348,In_1648);
nand U1689 (N_1689,In_2132,In_227);
or U1690 (N_1690,In_90,In_1581);
nand U1691 (N_1691,In_1795,In_1928);
nand U1692 (N_1692,In_207,In_1122);
and U1693 (N_1693,In_126,In_1563);
xor U1694 (N_1694,In_1711,In_248);
xor U1695 (N_1695,In_852,In_1692);
and U1696 (N_1696,In_2378,In_1583);
xnor U1697 (N_1697,In_1170,In_1404);
and U1698 (N_1698,In_498,In_476);
and U1699 (N_1699,In_1335,In_2167);
or U1700 (N_1700,In_884,In_89);
nand U1701 (N_1701,In_1396,In_1670);
xor U1702 (N_1702,In_2402,In_1253);
nor U1703 (N_1703,In_922,In_1727);
xnor U1704 (N_1704,In_1567,In_1537);
nor U1705 (N_1705,In_302,In_474);
xnor U1706 (N_1706,In_1455,In_1959);
or U1707 (N_1707,In_2230,In_2411);
and U1708 (N_1708,In_1116,In_1497);
nor U1709 (N_1709,In_2091,In_1767);
or U1710 (N_1710,In_622,In_2141);
and U1711 (N_1711,In_859,In_1298);
or U1712 (N_1712,In_1212,In_2001);
nor U1713 (N_1713,In_1645,In_1935);
and U1714 (N_1714,In_627,In_1455);
or U1715 (N_1715,In_408,In_1256);
nand U1716 (N_1716,In_1494,In_1649);
and U1717 (N_1717,In_1283,In_330);
nor U1718 (N_1718,In_942,In_104);
nor U1719 (N_1719,In_284,In_832);
nand U1720 (N_1720,In_804,In_799);
xnor U1721 (N_1721,In_1657,In_2414);
and U1722 (N_1722,In_2068,In_2073);
nor U1723 (N_1723,In_1173,In_1729);
and U1724 (N_1724,In_1897,In_2118);
nand U1725 (N_1725,In_2376,In_1171);
nor U1726 (N_1726,In_1643,In_456);
and U1727 (N_1727,In_916,In_711);
nand U1728 (N_1728,In_2346,In_1205);
or U1729 (N_1729,In_1351,In_1658);
nand U1730 (N_1730,In_1211,In_1019);
or U1731 (N_1731,In_495,In_1239);
xnor U1732 (N_1732,In_672,In_711);
nor U1733 (N_1733,In_1153,In_2394);
or U1734 (N_1734,In_58,In_364);
nor U1735 (N_1735,In_1723,In_837);
and U1736 (N_1736,In_2305,In_2418);
nor U1737 (N_1737,In_2102,In_2378);
nor U1738 (N_1738,In_19,In_606);
xor U1739 (N_1739,In_1561,In_1689);
and U1740 (N_1740,In_1593,In_1994);
nand U1741 (N_1741,In_175,In_1973);
xnor U1742 (N_1742,In_1217,In_1387);
nor U1743 (N_1743,In_664,In_2003);
xor U1744 (N_1744,In_473,In_2428);
nand U1745 (N_1745,In_1389,In_1333);
and U1746 (N_1746,In_1573,In_1788);
or U1747 (N_1747,In_1842,In_1018);
and U1748 (N_1748,In_238,In_474);
nand U1749 (N_1749,In_548,In_639);
and U1750 (N_1750,In_1855,In_1919);
xor U1751 (N_1751,In_2463,In_1890);
nor U1752 (N_1752,In_562,In_1288);
xor U1753 (N_1753,In_176,In_219);
and U1754 (N_1754,In_1650,In_951);
nand U1755 (N_1755,In_1590,In_1674);
nor U1756 (N_1756,In_1383,In_2452);
or U1757 (N_1757,In_59,In_984);
and U1758 (N_1758,In_805,In_384);
or U1759 (N_1759,In_577,In_614);
nor U1760 (N_1760,In_1854,In_364);
or U1761 (N_1761,In_2249,In_665);
and U1762 (N_1762,In_1160,In_459);
or U1763 (N_1763,In_414,In_962);
or U1764 (N_1764,In_176,In_1304);
nand U1765 (N_1765,In_767,In_2011);
nand U1766 (N_1766,In_2073,In_2263);
and U1767 (N_1767,In_2113,In_1924);
or U1768 (N_1768,In_618,In_948);
xor U1769 (N_1769,In_2039,In_2295);
nand U1770 (N_1770,In_1207,In_408);
or U1771 (N_1771,In_231,In_1155);
nor U1772 (N_1772,In_47,In_2363);
nor U1773 (N_1773,In_480,In_868);
and U1774 (N_1774,In_2044,In_1899);
and U1775 (N_1775,In_1651,In_1147);
and U1776 (N_1776,In_1201,In_1890);
xnor U1777 (N_1777,In_129,In_1299);
xor U1778 (N_1778,In_1379,In_415);
nor U1779 (N_1779,In_2423,In_444);
nand U1780 (N_1780,In_1837,In_1346);
or U1781 (N_1781,In_1342,In_1425);
or U1782 (N_1782,In_2469,In_2498);
or U1783 (N_1783,In_2248,In_1194);
and U1784 (N_1784,In_1880,In_150);
nor U1785 (N_1785,In_1313,In_1017);
and U1786 (N_1786,In_172,In_877);
nor U1787 (N_1787,In_1159,In_1991);
or U1788 (N_1788,In_2178,In_560);
nor U1789 (N_1789,In_464,In_186);
or U1790 (N_1790,In_502,In_1250);
nor U1791 (N_1791,In_1439,In_2344);
nor U1792 (N_1792,In_151,In_860);
xor U1793 (N_1793,In_42,In_2334);
nand U1794 (N_1794,In_559,In_891);
and U1795 (N_1795,In_467,In_1052);
and U1796 (N_1796,In_63,In_994);
and U1797 (N_1797,In_941,In_1177);
xor U1798 (N_1798,In_2165,In_701);
or U1799 (N_1799,In_1800,In_10);
and U1800 (N_1800,In_889,In_1066);
xnor U1801 (N_1801,In_1319,In_1068);
and U1802 (N_1802,In_535,In_2200);
nor U1803 (N_1803,In_1382,In_1469);
nor U1804 (N_1804,In_395,In_703);
and U1805 (N_1805,In_1872,In_2414);
and U1806 (N_1806,In_646,In_95);
and U1807 (N_1807,In_344,In_52);
nor U1808 (N_1808,In_1516,In_1979);
nor U1809 (N_1809,In_304,In_663);
or U1810 (N_1810,In_618,In_805);
or U1811 (N_1811,In_334,In_1294);
nand U1812 (N_1812,In_1327,In_770);
nand U1813 (N_1813,In_968,In_1888);
xor U1814 (N_1814,In_2173,In_2012);
nand U1815 (N_1815,In_795,In_422);
nor U1816 (N_1816,In_1113,In_142);
and U1817 (N_1817,In_1154,In_2477);
xor U1818 (N_1818,In_1505,In_218);
xnor U1819 (N_1819,In_2263,In_601);
or U1820 (N_1820,In_366,In_1249);
or U1821 (N_1821,In_1285,In_986);
nand U1822 (N_1822,In_1857,In_2182);
xnor U1823 (N_1823,In_858,In_1659);
and U1824 (N_1824,In_1618,In_335);
and U1825 (N_1825,In_2157,In_1431);
or U1826 (N_1826,In_1965,In_2327);
and U1827 (N_1827,In_1820,In_900);
nand U1828 (N_1828,In_1155,In_1518);
nor U1829 (N_1829,In_396,In_1293);
or U1830 (N_1830,In_1491,In_426);
xor U1831 (N_1831,In_322,In_2107);
nand U1832 (N_1832,In_2479,In_1164);
and U1833 (N_1833,In_524,In_772);
xnor U1834 (N_1834,In_1108,In_944);
nand U1835 (N_1835,In_1428,In_507);
and U1836 (N_1836,In_560,In_1106);
xor U1837 (N_1837,In_43,In_897);
or U1838 (N_1838,In_1799,In_1778);
or U1839 (N_1839,In_1003,In_928);
or U1840 (N_1840,In_740,In_871);
or U1841 (N_1841,In_855,In_2356);
or U1842 (N_1842,In_729,In_2108);
and U1843 (N_1843,In_1100,In_630);
xor U1844 (N_1844,In_975,In_881);
xnor U1845 (N_1845,In_7,In_52);
xor U1846 (N_1846,In_2432,In_1306);
nor U1847 (N_1847,In_863,In_120);
and U1848 (N_1848,In_2496,In_204);
nor U1849 (N_1849,In_2212,In_429);
nor U1850 (N_1850,In_964,In_1444);
nand U1851 (N_1851,In_1829,In_548);
xor U1852 (N_1852,In_1667,In_1642);
xnor U1853 (N_1853,In_927,In_1867);
nor U1854 (N_1854,In_2395,In_2333);
nand U1855 (N_1855,In_1690,In_1767);
and U1856 (N_1856,In_1126,In_58);
xor U1857 (N_1857,In_1162,In_1144);
xor U1858 (N_1858,In_1362,In_1481);
xor U1859 (N_1859,In_1840,In_57);
nor U1860 (N_1860,In_1121,In_1470);
or U1861 (N_1861,In_2286,In_448);
nand U1862 (N_1862,In_507,In_2349);
or U1863 (N_1863,In_1126,In_931);
or U1864 (N_1864,In_2275,In_2359);
nand U1865 (N_1865,In_1298,In_39);
nand U1866 (N_1866,In_461,In_385);
or U1867 (N_1867,In_1230,In_959);
nand U1868 (N_1868,In_2409,In_1674);
or U1869 (N_1869,In_2396,In_2432);
or U1870 (N_1870,In_412,In_1276);
xor U1871 (N_1871,In_2062,In_165);
xnor U1872 (N_1872,In_1356,In_589);
and U1873 (N_1873,In_163,In_1671);
nand U1874 (N_1874,In_579,In_756);
or U1875 (N_1875,In_409,In_412);
xnor U1876 (N_1876,In_258,In_43);
or U1877 (N_1877,In_1673,In_1944);
nand U1878 (N_1878,In_2393,In_1206);
nor U1879 (N_1879,In_2083,In_1702);
nor U1880 (N_1880,In_345,In_984);
or U1881 (N_1881,In_32,In_480);
xnor U1882 (N_1882,In_2063,In_376);
nor U1883 (N_1883,In_2132,In_985);
nor U1884 (N_1884,In_1817,In_1399);
nor U1885 (N_1885,In_1453,In_1201);
or U1886 (N_1886,In_222,In_321);
and U1887 (N_1887,In_2213,In_2350);
and U1888 (N_1888,In_2149,In_2195);
and U1889 (N_1889,In_478,In_2092);
and U1890 (N_1890,In_180,In_218);
xor U1891 (N_1891,In_1020,In_2192);
nand U1892 (N_1892,In_1326,In_2258);
and U1893 (N_1893,In_499,In_1841);
nand U1894 (N_1894,In_2150,In_2405);
or U1895 (N_1895,In_503,In_2295);
and U1896 (N_1896,In_1806,In_1236);
nor U1897 (N_1897,In_28,In_1151);
and U1898 (N_1898,In_1388,In_529);
xor U1899 (N_1899,In_2115,In_2106);
nor U1900 (N_1900,In_1672,In_199);
or U1901 (N_1901,In_1854,In_2125);
xor U1902 (N_1902,In_785,In_834);
xor U1903 (N_1903,In_1909,In_1838);
nand U1904 (N_1904,In_2404,In_1192);
nand U1905 (N_1905,In_2265,In_2137);
xor U1906 (N_1906,In_392,In_1157);
nand U1907 (N_1907,In_35,In_885);
nor U1908 (N_1908,In_2219,In_1906);
nor U1909 (N_1909,In_1839,In_1936);
xnor U1910 (N_1910,In_557,In_1988);
nor U1911 (N_1911,In_1284,In_2280);
nor U1912 (N_1912,In_1684,In_2381);
xor U1913 (N_1913,In_1884,In_17);
nor U1914 (N_1914,In_1590,In_1316);
nor U1915 (N_1915,In_437,In_1012);
nand U1916 (N_1916,In_245,In_501);
xnor U1917 (N_1917,In_1261,In_1601);
xor U1918 (N_1918,In_614,In_1395);
xor U1919 (N_1919,In_413,In_22);
nor U1920 (N_1920,In_1941,In_813);
xor U1921 (N_1921,In_2276,In_629);
xor U1922 (N_1922,In_2033,In_121);
xor U1923 (N_1923,In_132,In_2008);
nand U1924 (N_1924,In_1663,In_2343);
and U1925 (N_1925,In_978,In_566);
or U1926 (N_1926,In_766,In_893);
nor U1927 (N_1927,In_820,In_1897);
or U1928 (N_1928,In_605,In_2214);
or U1929 (N_1929,In_674,In_2304);
xnor U1930 (N_1930,In_775,In_465);
nor U1931 (N_1931,In_19,In_547);
and U1932 (N_1932,In_2079,In_110);
and U1933 (N_1933,In_2304,In_195);
nor U1934 (N_1934,In_1643,In_1438);
xnor U1935 (N_1935,In_575,In_1650);
nand U1936 (N_1936,In_2190,In_627);
or U1937 (N_1937,In_773,In_1061);
or U1938 (N_1938,In_1394,In_1940);
nor U1939 (N_1939,In_544,In_2115);
or U1940 (N_1940,In_1227,In_2215);
nand U1941 (N_1941,In_1496,In_343);
xnor U1942 (N_1942,In_1669,In_335);
nor U1943 (N_1943,In_78,In_2262);
and U1944 (N_1944,In_2107,In_1440);
nor U1945 (N_1945,In_343,In_1321);
and U1946 (N_1946,In_1913,In_1019);
xor U1947 (N_1947,In_1856,In_1802);
xnor U1948 (N_1948,In_1742,In_473);
nor U1949 (N_1949,In_1254,In_1547);
and U1950 (N_1950,In_595,In_1056);
xor U1951 (N_1951,In_1627,In_1928);
nand U1952 (N_1952,In_1627,In_1105);
nand U1953 (N_1953,In_2335,In_747);
and U1954 (N_1954,In_2040,In_205);
and U1955 (N_1955,In_2311,In_536);
xnor U1956 (N_1956,In_1298,In_2470);
or U1957 (N_1957,In_1877,In_1738);
xnor U1958 (N_1958,In_2284,In_2319);
or U1959 (N_1959,In_2168,In_729);
nand U1960 (N_1960,In_1984,In_940);
xnor U1961 (N_1961,In_1905,In_1944);
or U1962 (N_1962,In_2317,In_206);
xor U1963 (N_1963,In_769,In_2130);
nand U1964 (N_1964,In_704,In_1606);
and U1965 (N_1965,In_1194,In_424);
nor U1966 (N_1966,In_2214,In_910);
nand U1967 (N_1967,In_1332,In_2143);
nand U1968 (N_1968,In_289,In_2126);
and U1969 (N_1969,In_573,In_503);
nand U1970 (N_1970,In_1901,In_628);
nand U1971 (N_1971,In_1063,In_2458);
nor U1972 (N_1972,In_176,In_82);
nand U1973 (N_1973,In_1629,In_694);
nand U1974 (N_1974,In_1935,In_91);
nor U1975 (N_1975,In_387,In_344);
nand U1976 (N_1976,In_1003,In_143);
xnor U1977 (N_1977,In_1370,In_1998);
and U1978 (N_1978,In_1379,In_2355);
nand U1979 (N_1979,In_1862,In_1379);
and U1980 (N_1980,In_1329,In_580);
xor U1981 (N_1981,In_1637,In_1071);
nand U1982 (N_1982,In_382,In_22);
xnor U1983 (N_1983,In_1192,In_820);
and U1984 (N_1984,In_601,In_2388);
and U1985 (N_1985,In_2449,In_2355);
and U1986 (N_1986,In_2458,In_1235);
nand U1987 (N_1987,In_1869,In_1428);
or U1988 (N_1988,In_2248,In_1114);
and U1989 (N_1989,In_511,In_1486);
xnor U1990 (N_1990,In_1087,In_628);
nand U1991 (N_1991,In_2291,In_2227);
xor U1992 (N_1992,In_1285,In_377);
and U1993 (N_1993,In_683,In_1072);
or U1994 (N_1994,In_2130,In_1985);
nor U1995 (N_1995,In_2290,In_2195);
or U1996 (N_1996,In_558,In_2055);
nor U1997 (N_1997,In_794,In_789);
nand U1998 (N_1998,In_1770,In_1711);
nand U1999 (N_1999,In_1327,In_1576);
xor U2000 (N_2000,In_891,In_1703);
nor U2001 (N_2001,In_580,In_1298);
nor U2002 (N_2002,In_450,In_1909);
or U2003 (N_2003,In_677,In_1672);
xnor U2004 (N_2004,In_18,In_33);
nor U2005 (N_2005,In_826,In_1025);
and U2006 (N_2006,In_1336,In_1176);
xor U2007 (N_2007,In_319,In_671);
and U2008 (N_2008,In_172,In_116);
nor U2009 (N_2009,In_1222,In_329);
nand U2010 (N_2010,In_522,In_1971);
and U2011 (N_2011,In_2234,In_531);
nand U2012 (N_2012,In_393,In_1648);
and U2013 (N_2013,In_1977,In_2105);
nor U2014 (N_2014,In_1059,In_294);
nand U2015 (N_2015,In_1823,In_336);
nand U2016 (N_2016,In_940,In_934);
nor U2017 (N_2017,In_744,In_1417);
or U2018 (N_2018,In_488,In_1499);
or U2019 (N_2019,In_1357,In_1381);
nand U2020 (N_2020,In_431,In_17);
or U2021 (N_2021,In_2302,In_1410);
and U2022 (N_2022,In_1468,In_737);
nor U2023 (N_2023,In_2470,In_550);
xor U2024 (N_2024,In_1426,In_2020);
xor U2025 (N_2025,In_1676,In_412);
nor U2026 (N_2026,In_972,In_1041);
nor U2027 (N_2027,In_1206,In_2262);
and U2028 (N_2028,In_605,In_1053);
xor U2029 (N_2029,In_1229,In_2142);
nand U2030 (N_2030,In_1826,In_2419);
or U2031 (N_2031,In_1724,In_12);
xor U2032 (N_2032,In_1576,In_2258);
nand U2033 (N_2033,In_1841,In_267);
or U2034 (N_2034,In_1059,In_1244);
or U2035 (N_2035,In_2053,In_1798);
nand U2036 (N_2036,In_1211,In_1086);
and U2037 (N_2037,In_1673,In_2490);
xor U2038 (N_2038,In_2089,In_1083);
and U2039 (N_2039,In_1898,In_800);
xnor U2040 (N_2040,In_128,In_2462);
or U2041 (N_2041,In_1356,In_55);
xnor U2042 (N_2042,In_254,In_687);
or U2043 (N_2043,In_992,In_1214);
and U2044 (N_2044,In_508,In_1431);
nor U2045 (N_2045,In_1273,In_722);
nor U2046 (N_2046,In_280,In_2183);
or U2047 (N_2047,In_2456,In_507);
nor U2048 (N_2048,In_181,In_243);
and U2049 (N_2049,In_1012,In_857);
nor U2050 (N_2050,In_1889,In_2202);
or U2051 (N_2051,In_310,In_1719);
nor U2052 (N_2052,In_994,In_638);
and U2053 (N_2053,In_1032,In_535);
or U2054 (N_2054,In_29,In_2417);
or U2055 (N_2055,In_871,In_2213);
or U2056 (N_2056,In_69,In_371);
nand U2057 (N_2057,In_1146,In_2161);
or U2058 (N_2058,In_82,In_1787);
or U2059 (N_2059,In_1249,In_170);
nand U2060 (N_2060,In_210,In_1371);
xor U2061 (N_2061,In_793,In_1604);
nand U2062 (N_2062,In_1065,In_1028);
xor U2063 (N_2063,In_2474,In_2196);
nand U2064 (N_2064,In_204,In_1134);
xnor U2065 (N_2065,In_917,In_1265);
xor U2066 (N_2066,In_607,In_2018);
nand U2067 (N_2067,In_1812,In_1323);
xor U2068 (N_2068,In_1789,In_567);
or U2069 (N_2069,In_2375,In_67);
nor U2070 (N_2070,In_1738,In_1813);
xnor U2071 (N_2071,In_326,In_1732);
xor U2072 (N_2072,In_441,In_2088);
xor U2073 (N_2073,In_86,In_1706);
nand U2074 (N_2074,In_2252,In_1056);
nand U2075 (N_2075,In_2097,In_1961);
and U2076 (N_2076,In_1903,In_132);
nand U2077 (N_2077,In_1596,In_1853);
and U2078 (N_2078,In_1354,In_423);
and U2079 (N_2079,In_401,In_750);
and U2080 (N_2080,In_2113,In_2167);
nand U2081 (N_2081,In_1418,In_2141);
and U2082 (N_2082,In_2466,In_294);
or U2083 (N_2083,In_59,In_655);
and U2084 (N_2084,In_1863,In_933);
or U2085 (N_2085,In_1058,In_624);
nor U2086 (N_2086,In_1908,In_103);
nor U2087 (N_2087,In_821,In_604);
or U2088 (N_2088,In_2089,In_1569);
and U2089 (N_2089,In_739,In_957);
and U2090 (N_2090,In_2316,In_670);
or U2091 (N_2091,In_1643,In_714);
or U2092 (N_2092,In_2352,In_34);
xnor U2093 (N_2093,In_1421,In_1269);
nand U2094 (N_2094,In_1069,In_984);
nor U2095 (N_2095,In_1843,In_329);
and U2096 (N_2096,In_2488,In_2451);
nor U2097 (N_2097,In_398,In_1701);
or U2098 (N_2098,In_2157,In_1111);
and U2099 (N_2099,In_1230,In_1139);
nor U2100 (N_2100,In_925,In_209);
and U2101 (N_2101,In_2046,In_2181);
nand U2102 (N_2102,In_1344,In_536);
nand U2103 (N_2103,In_225,In_1023);
nor U2104 (N_2104,In_495,In_67);
nand U2105 (N_2105,In_1468,In_1385);
and U2106 (N_2106,In_1338,In_137);
nand U2107 (N_2107,In_2329,In_669);
and U2108 (N_2108,In_1243,In_2335);
and U2109 (N_2109,In_618,In_1536);
nand U2110 (N_2110,In_1499,In_1326);
or U2111 (N_2111,In_1331,In_1413);
nor U2112 (N_2112,In_341,In_2427);
nor U2113 (N_2113,In_1609,In_1050);
or U2114 (N_2114,In_819,In_2344);
and U2115 (N_2115,In_371,In_1153);
and U2116 (N_2116,In_1416,In_2224);
nor U2117 (N_2117,In_2275,In_2379);
nand U2118 (N_2118,In_866,In_1063);
nand U2119 (N_2119,In_2247,In_1768);
xnor U2120 (N_2120,In_765,In_199);
xor U2121 (N_2121,In_1178,In_1922);
nand U2122 (N_2122,In_866,In_865);
nand U2123 (N_2123,In_1033,In_1540);
xor U2124 (N_2124,In_1088,In_1622);
xnor U2125 (N_2125,In_857,In_1375);
nor U2126 (N_2126,In_2109,In_1130);
xor U2127 (N_2127,In_1449,In_1941);
nand U2128 (N_2128,In_102,In_196);
nor U2129 (N_2129,In_1931,In_1204);
and U2130 (N_2130,In_1424,In_2042);
nand U2131 (N_2131,In_2435,In_1440);
xnor U2132 (N_2132,In_1551,In_2233);
or U2133 (N_2133,In_887,In_523);
and U2134 (N_2134,In_299,In_1423);
xor U2135 (N_2135,In_1443,In_1339);
nand U2136 (N_2136,In_1619,In_237);
nand U2137 (N_2137,In_8,In_23);
xnor U2138 (N_2138,In_1991,In_2053);
nor U2139 (N_2139,In_1502,In_2413);
xor U2140 (N_2140,In_159,In_241);
nand U2141 (N_2141,In_384,In_1920);
or U2142 (N_2142,In_1059,In_1058);
nand U2143 (N_2143,In_1787,In_446);
nor U2144 (N_2144,In_202,In_2356);
or U2145 (N_2145,In_166,In_2117);
or U2146 (N_2146,In_89,In_886);
and U2147 (N_2147,In_2157,In_434);
nor U2148 (N_2148,In_2041,In_2451);
nand U2149 (N_2149,In_1223,In_1702);
nor U2150 (N_2150,In_1453,In_1116);
xnor U2151 (N_2151,In_1407,In_1801);
or U2152 (N_2152,In_143,In_1369);
nand U2153 (N_2153,In_940,In_1681);
or U2154 (N_2154,In_1927,In_2436);
nand U2155 (N_2155,In_1922,In_1073);
xor U2156 (N_2156,In_657,In_1246);
or U2157 (N_2157,In_1658,In_838);
or U2158 (N_2158,In_2428,In_1123);
and U2159 (N_2159,In_1679,In_2109);
or U2160 (N_2160,In_1914,In_296);
nor U2161 (N_2161,In_2114,In_1500);
and U2162 (N_2162,In_2429,In_504);
nor U2163 (N_2163,In_1681,In_580);
nor U2164 (N_2164,In_1367,In_23);
xnor U2165 (N_2165,In_1244,In_2273);
and U2166 (N_2166,In_2373,In_78);
nor U2167 (N_2167,In_495,In_620);
or U2168 (N_2168,In_2137,In_94);
nor U2169 (N_2169,In_2304,In_1379);
nand U2170 (N_2170,In_2436,In_2093);
and U2171 (N_2171,In_1417,In_2225);
and U2172 (N_2172,In_85,In_767);
xnor U2173 (N_2173,In_2155,In_1408);
nor U2174 (N_2174,In_938,In_1391);
nand U2175 (N_2175,In_2474,In_2105);
or U2176 (N_2176,In_1061,In_1648);
and U2177 (N_2177,In_1317,In_218);
nand U2178 (N_2178,In_1397,In_1263);
xor U2179 (N_2179,In_1659,In_1656);
nor U2180 (N_2180,In_2262,In_1903);
and U2181 (N_2181,In_1129,In_673);
xor U2182 (N_2182,In_1292,In_1030);
and U2183 (N_2183,In_789,In_718);
nor U2184 (N_2184,In_313,In_1182);
xor U2185 (N_2185,In_417,In_1653);
nor U2186 (N_2186,In_145,In_397);
and U2187 (N_2187,In_2446,In_2346);
or U2188 (N_2188,In_578,In_2397);
xnor U2189 (N_2189,In_557,In_1351);
or U2190 (N_2190,In_74,In_1793);
or U2191 (N_2191,In_1216,In_2195);
and U2192 (N_2192,In_1868,In_1233);
or U2193 (N_2193,In_750,In_47);
xnor U2194 (N_2194,In_855,In_596);
nor U2195 (N_2195,In_1691,In_2094);
or U2196 (N_2196,In_1182,In_385);
and U2197 (N_2197,In_252,In_980);
or U2198 (N_2198,In_910,In_997);
and U2199 (N_2199,In_1039,In_100);
nor U2200 (N_2200,In_1437,In_1636);
or U2201 (N_2201,In_1109,In_583);
xor U2202 (N_2202,In_2281,In_1897);
xnor U2203 (N_2203,In_1490,In_991);
nand U2204 (N_2204,In_865,In_1659);
nand U2205 (N_2205,In_2163,In_35);
xor U2206 (N_2206,In_1440,In_1978);
xnor U2207 (N_2207,In_2032,In_1741);
nand U2208 (N_2208,In_1359,In_1946);
or U2209 (N_2209,In_2035,In_1722);
xor U2210 (N_2210,In_906,In_614);
and U2211 (N_2211,In_2039,In_1203);
nor U2212 (N_2212,In_532,In_761);
xor U2213 (N_2213,In_400,In_2167);
xor U2214 (N_2214,In_1282,In_1736);
nand U2215 (N_2215,In_2402,In_142);
xnor U2216 (N_2216,In_59,In_970);
nand U2217 (N_2217,In_480,In_126);
nand U2218 (N_2218,In_1578,In_1777);
xnor U2219 (N_2219,In_404,In_160);
nand U2220 (N_2220,In_1590,In_1266);
nor U2221 (N_2221,In_2476,In_1207);
and U2222 (N_2222,In_1534,In_2067);
xnor U2223 (N_2223,In_1138,In_1570);
or U2224 (N_2224,In_2230,In_526);
or U2225 (N_2225,In_1782,In_1980);
or U2226 (N_2226,In_645,In_2277);
nor U2227 (N_2227,In_1905,In_2102);
nor U2228 (N_2228,In_189,In_1165);
nand U2229 (N_2229,In_692,In_1303);
and U2230 (N_2230,In_1510,In_2275);
nand U2231 (N_2231,In_1228,In_939);
or U2232 (N_2232,In_1413,In_2152);
and U2233 (N_2233,In_1639,In_435);
or U2234 (N_2234,In_2088,In_1347);
xnor U2235 (N_2235,In_1662,In_970);
or U2236 (N_2236,In_1725,In_720);
and U2237 (N_2237,In_551,In_1006);
nor U2238 (N_2238,In_2475,In_886);
and U2239 (N_2239,In_1115,In_287);
xor U2240 (N_2240,In_724,In_1896);
xor U2241 (N_2241,In_543,In_212);
xor U2242 (N_2242,In_495,In_273);
or U2243 (N_2243,In_1538,In_2326);
or U2244 (N_2244,In_966,In_2112);
xor U2245 (N_2245,In_357,In_155);
nor U2246 (N_2246,In_1977,In_1127);
or U2247 (N_2247,In_1360,In_1585);
nor U2248 (N_2248,In_1550,In_705);
xor U2249 (N_2249,In_1472,In_6);
nor U2250 (N_2250,In_98,In_1545);
or U2251 (N_2251,In_5,In_2159);
and U2252 (N_2252,In_856,In_1476);
nand U2253 (N_2253,In_329,In_913);
nand U2254 (N_2254,In_2345,In_1366);
and U2255 (N_2255,In_530,In_2322);
and U2256 (N_2256,In_342,In_1240);
xnor U2257 (N_2257,In_609,In_2053);
xnor U2258 (N_2258,In_2119,In_67);
xor U2259 (N_2259,In_843,In_1442);
and U2260 (N_2260,In_207,In_1070);
and U2261 (N_2261,In_1123,In_2037);
and U2262 (N_2262,In_1963,In_854);
xor U2263 (N_2263,In_684,In_1249);
and U2264 (N_2264,In_2209,In_290);
nor U2265 (N_2265,In_1518,In_2222);
xor U2266 (N_2266,In_1508,In_2426);
or U2267 (N_2267,In_1090,In_1591);
or U2268 (N_2268,In_1718,In_2303);
and U2269 (N_2269,In_2126,In_406);
nand U2270 (N_2270,In_1025,In_1755);
and U2271 (N_2271,In_114,In_1672);
nor U2272 (N_2272,In_679,In_2185);
and U2273 (N_2273,In_327,In_1615);
xor U2274 (N_2274,In_577,In_495);
and U2275 (N_2275,In_819,In_1251);
nand U2276 (N_2276,In_679,In_856);
or U2277 (N_2277,In_1775,In_2451);
nor U2278 (N_2278,In_707,In_1831);
and U2279 (N_2279,In_167,In_2368);
nand U2280 (N_2280,In_1009,In_685);
and U2281 (N_2281,In_915,In_604);
nand U2282 (N_2282,In_2181,In_125);
xnor U2283 (N_2283,In_1471,In_1947);
and U2284 (N_2284,In_74,In_1387);
or U2285 (N_2285,In_397,In_1851);
xor U2286 (N_2286,In_738,In_2037);
xnor U2287 (N_2287,In_1750,In_912);
or U2288 (N_2288,In_1143,In_1246);
and U2289 (N_2289,In_357,In_1171);
nand U2290 (N_2290,In_2191,In_819);
nor U2291 (N_2291,In_264,In_1418);
xnor U2292 (N_2292,In_1380,In_996);
nand U2293 (N_2293,In_1020,In_1864);
and U2294 (N_2294,In_86,In_2085);
xor U2295 (N_2295,In_440,In_1623);
or U2296 (N_2296,In_2397,In_1553);
and U2297 (N_2297,In_1345,In_2117);
nor U2298 (N_2298,In_280,In_1305);
nor U2299 (N_2299,In_1357,In_1694);
or U2300 (N_2300,In_398,In_2477);
and U2301 (N_2301,In_1262,In_1409);
or U2302 (N_2302,In_1063,In_850);
or U2303 (N_2303,In_1256,In_1248);
or U2304 (N_2304,In_778,In_1502);
xor U2305 (N_2305,In_1570,In_1203);
and U2306 (N_2306,In_1851,In_156);
or U2307 (N_2307,In_353,In_1099);
xor U2308 (N_2308,In_421,In_1812);
or U2309 (N_2309,In_570,In_715);
or U2310 (N_2310,In_2146,In_919);
xor U2311 (N_2311,In_2368,In_856);
xnor U2312 (N_2312,In_1471,In_621);
nor U2313 (N_2313,In_2285,In_323);
and U2314 (N_2314,In_1265,In_1428);
or U2315 (N_2315,In_472,In_2450);
xnor U2316 (N_2316,In_1600,In_1163);
nand U2317 (N_2317,In_422,In_1383);
nor U2318 (N_2318,In_1274,In_528);
nor U2319 (N_2319,In_365,In_2031);
or U2320 (N_2320,In_974,In_1144);
or U2321 (N_2321,In_983,In_579);
xnor U2322 (N_2322,In_2296,In_77);
nor U2323 (N_2323,In_2029,In_516);
xor U2324 (N_2324,In_660,In_271);
and U2325 (N_2325,In_412,In_1044);
and U2326 (N_2326,In_1550,In_1139);
xor U2327 (N_2327,In_863,In_218);
nand U2328 (N_2328,In_743,In_1495);
or U2329 (N_2329,In_854,In_966);
nand U2330 (N_2330,In_618,In_576);
and U2331 (N_2331,In_483,In_1592);
xnor U2332 (N_2332,In_88,In_203);
and U2333 (N_2333,In_2283,In_165);
nand U2334 (N_2334,In_149,In_1399);
and U2335 (N_2335,In_1304,In_1141);
xnor U2336 (N_2336,In_2023,In_1526);
nand U2337 (N_2337,In_205,In_1552);
and U2338 (N_2338,In_939,In_879);
or U2339 (N_2339,In_1892,In_2491);
nand U2340 (N_2340,In_494,In_981);
or U2341 (N_2341,In_131,In_947);
nand U2342 (N_2342,In_2374,In_1651);
or U2343 (N_2343,In_212,In_940);
nand U2344 (N_2344,In_1496,In_1184);
xor U2345 (N_2345,In_1647,In_1523);
or U2346 (N_2346,In_2103,In_100);
and U2347 (N_2347,In_944,In_89);
nor U2348 (N_2348,In_997,In_1906);
xnor U2349 (N_2349,In_600,In_106);
nand U2350 (N_2350,In_325,In_1862);
nor U2351 (N_2351,In_970,In_68);
and U2352 (N_2352,In_1605,In_1590);
and U2353 (N_2353,In_8,In_1697);
and U2354 (N_2354,In_1594,In_1436);
nor U2355 (N_2355,In_738,In_1649);
nor U2356 (N_2356,In_1624,In_16);
or U2357 (N_2357,In_1864,In_1276);
nor U2358 (N_2358,In_1073,In_992);
and U2359 (N_2359,In_2403,In_566);
nand U2360 (N_2360,In_377,In_455);
nor U2361 (N_2361,In_918,In_297);
or U2362 (N_2362,In_2011,In_2068);
nor U2363 (N_2363,In_1107,In_1622);
nand U2364 (N_2364,In_1642,In_2475);
nor U2365 (N_2365,In_2271,In_1742);
or U2366 (N_2366,In_1462,In_88);
xnor U2367 (N_2367,In_1046,In_1820);
nand U2368 (N_2368,In_1941,In_1729);
or U2369 (N_2369,In_199,In_396);
and U2370 (N_2370,In_152,In_1329);
or U2371 (N_2371,In_2130,In_847);
xor U2372 (N_2372,In_749,In_2218);
nor U2373 (N_2373,In_1114,In_334);
xor U2374 (N_2374,In_94,In_1584);
xnor U2375 (N_2375,In_168,In_2061);
nand U2376 (N_2376,In_1533,In_1584);
or U2377 (N_2377,In_978,In_230);
or U2378 (N_2378,In_941,In_1790);
nor U2379 (N_2379,In_145,In_1006);
xor U2380 (N_2380,In_550,In_883);
nor U2381 (N_2381,In_1121,In_12);
xor U2382 (N_2382,In_1312,In_2041);
or U2383 (N_2383,In_1072,In_1027);
nor U2384 (N_2384,In_647,In_512);
and U2385 (N_2385,In_32,In_395);
xnor U2386 (N_2386,In_303,In_1103);
and U2387 (N_2387,In_1963,In_2317);
xor U2388 (N_2388,In_689,In_1);
nor U2389 (N_2389,In_91,In_1845);
xor U2390 (N_2390,In_804,In_2157);
and U2391 (N_2391,In_248,In_2186);
and U2392 (N_2392,In_240,In_1587);
nor U2393 (N_2393,In_1013,In_266);
xor U2394 (N_2394,In_1010,In_1954);
nor U2395 (N_2395,In_1309,In_1698);
nor U2396 (N_2396,In_1667,In_229);
nor U2397 (N_2397,In_1636,In_1047);
nand U2398 (N_2398,In_1805,In_1153);
nor U2399 (N_2399,In_1155,In_1355);
or U2400 (N_2400,In_1233,In_490);
xnor U2401 (N_2401,In_102,In_963);
nor U2402 (N_2402,In_994,In_1732);
nor U2403 (N_2403,In_583,In_2365);
or U2404 (N_2404,In_361,In_1589);
nor U2405 (N_2405,In_506,In_1728);
nor U2406 (N_2406,In_1101,In_2454);
nor U2407 (N_2407,In_1249,In_1965);
or U2408 (N_2408,In_2063,In_149);
and U2409 (N_2409,In_2205,In_882);
xnor U2410 (N_2410,In_246,In_1746);
nor U2411 (N_2411,In_981,In_2084);
or U2412 (N_2412,In_126,In_555);
or U2413 (N_2413,In_259,In_80);
or U2414 (N_2414,In_261,In_836);
and U2415 (N_2415,In_115,In_2498);
xnor U2416 (N_2416,In_879,In_520);
nand U2417 (N_2417,In_1061,In_102);
and U2418 (N_2418,In_825,In_163);
or U2419 (N_2419,In_2444,In_612);
xnor U2420 (N_2420,In_391,In_1636);
or U2421 (N_2421,In_437,In_2053);
nand U2422 (N_2422,In_1855,In_1472);
nor U2423 (N_2423,In_148,In_2478);
nand U2424 (N_2424,In_2346,In_1190);
or U2425 (N_2425,In_138,In_1933);
nand U2426 (N_2426,In_1727,In_1386);
nor U2427 (N_2427,In_2070,In_27);
xnor U2428 (N_2428,In_1236,In_1519);
xnor U2429 (N_2429,In_68,In_1985);
nand U2430 (N_2430,In_1032,In_2232);
xnor U2431 (N_2431,In_2414,In_406);
or U2432 (N_2432,In_1037,In_645);
or U2433 (N_2433,In_2127,In_1194);
nand U2434 (N_2434,In_1913,In_2042);
or U2435 (N_2435,In_1198,In_697);
and U2436 (N_2436,In_2073,In_1438);
and U2437 (N_2437,In_398,In_585);
xor U2438 (N_2438,In_72,In_899);
nor U2439 (N_2439,In_2002,In_1748);
or U2440 (N_2440,In_873,In_2189);
and U2441 (N_2441,In_2069,In_1666);
and U2442 (N_2442,In_2460,In_231);
and U2443 (N_2443,In_1540,In_136);
nor U2444 (N_2444,In_607,In_2026);
or U2445 (N_2445,In_1098,In_36);
nand U2446 (N_2446,In_1169,In_1220);
xor U2447 (N_2447,In_369,In_803);
nor U2448 (N_2448,In_2048,In_579);
and U2449 (N_2449,In_2165,In_1608);
xor U2450 (N_2450,In_774,In_1867);
and U2451 (N_2451,In_898,In_2326);
nand U2452 (N_2452,In_787,In_476);
or U2453 (N_2453,In_1883,In_2019);
and U2454 (N_2454,In_1252,In_437);
or U2455 (N_2455,In_360,In_2042);
nand U2456 (N_2456,In_819,In_1241);
xnor U2457 (N_2457,In_1259,In_2361);
xnor U2458 (N_2458,In_1847,In_58);
and U2459 (N_2459,In_1155,In_31);
or U2460 (N_2460,In_1025,In_1237);
nor U2461 (N_2461,In_1281,In_134);
and U2462 (N_2462,In_1210,In_252);
nor U2463 (N_2463,In_542,In_1102);
nand U2464 (N_2464,In_659,In_1546);
nand U2465 (N_2465,In_416,In_188);
nand U2466 (N_2466,In_482,In_1840);
xnor U2467 (N_2467,In_1552,In_716);
xor U2468 (N_2468,In_1601,In_1975);
nand U2469 (N_2469,In_1271,In_380);
nand U2470 (N_2470,In_2422,In_2306);
nor U2471 (N_2471,In_2368,In_1428);
or U2472 (N_2472,In_1718,In_987);
xor U2473 (N_2473,In_2150,In_339);
or U2474 (N_2474,In_1244,In_877);
and U2475 (N_2475,In_1190,In_1535);
xnor U2476 (N_2476,In_2000,In_347);
nand U2477 (N_2477,In_1441,In_995);
and U2478 (N_2478,In_240,In_47);
or U2479 (N_2479,In_1395,In_942);
xor U2480 (N_2480,In_377,In_540);
nand U2481 (N_2481,In_375,In_715);
nand U2482 (N_2482,In_1702,In_1622);
nand U2483 (N_2483,In_357,In_161);
nor U2484 (N_2484,In_39,In_510);
and U2485 (N_2485,In_977,In_2447);
xnor U2486 (N_2486,In_2101,In_428);
nor U2487 (N_2487,In_267,In_444);
xnor U2488 (N_2488,In_160,In_1000);
xor U2489 (N_2489,In_472,In_676);
or U2490 (N_2490,In_1360,In_1754);
or U2491 (N_2491,In_400,In_2154);
xnor U2492 (N_2492,In_2244,In_1063);
xnor U2493 (N_2493,In_199,In_2300);
nand U2494 (N_2494,In_241,In_1454);
nor U2495 (N_2495,In_2078,In_1909);
and U2496 (N_2496,In_1135,In_2355);
or U2497 (N_2497,In_1637,In_1843);
or U2498 (N_2498,In_2324,In_1846);
xnor U2499 (N_2499,In_1455,In_746);
nor U2500 (N_2500,In_1008,In_1927);
nand U2501 (N_2501,In_2395,In_1159);
and U2502 (N_2502,In_524,In_1008);
nor U2503 (N_2503,In_147,In_1332);
nand U2504 (N_2504,In_1278,In_1733);
nand U2505 (N_2505,In_817,In_638);
nor U2506 (N_2506,In_2492,In_2006);
xnor U2507 (N_2507,In_2380,In_1702);
or U2508 (N_2508,In_865,In_2499);
nand U2509 (N_2509,In_252,In_215);
xor U2510 (N_2510,In_1625,In_998);
nand U2511 (N_2511,In_1819,In_2055);
nor U2512 (N_2512,In_627,In_2302);
nor U2513 (N_2513,In_1402,In_2358);
nor U2514 (N_2514,In_1432,In_1294);
nor U2515 (N_2515,In_238,In_2165);
or U2516 (N_2516,In_1896,In_2136);
or U2517 (N_2517,In_689,In_1504);
xor U2518 (N_2518,In_1210,In_2167);
or U2519 (N_2519,In_674,In_1124);
or U2520 (N_2520,In_396,In_1186);
or U2521 (N_2521,In_295,In_979);
or U2522 (N_2522,In_1894,In_974);
and U2523 (N_2523,In_2128,In_1337);
xor U2524 (N_2524,In_2118,In_2396);
xnor U2525 (N_2525,In_199,In_388);
nor U2526 (N_2526,In_2389,In_1759);
or U2527 (N_2527,In_508,In_1029);
nor U2528 (N_2528,In_914,In_583);
and U2529 (N_2529,In_591,In_163);
nand U2530 (N_2530,In_200,In_1099);
and U2531 (N_2531,In_1210,In_1402);
or U2532 (N_2532,In_2019,In_2486);
xnor U2533 (N_2533,In_1449,In_1347);
nor U2534 (N_2534,In_932,In_665);
or U2535 (N_2535,In_1897,In_425);
and U2536 (N_2536,In_139,In_961);
nor U2537 (N_2537,In_181,In_1060);
nor U2538 (N_2538,In_1071,In_373);
xnor U2539 (N_2539,In_1710,In_1104);
or U2540 (N_2540,In_2302,In_2409);
xnor U2541 (N_2541,In_286,In_344);
nor U2542 (N_2542,In_2329,In_165);
nand U2543 (N_2543,In_529,In_649);
or U2544 (N_2544,In_1215,In_1634);
or U2545 (N_2545,In_2492,In_618);
and U2546 (N_2546,In_806,In_602);
or U2547 (N_2547,In_2090,In_1915);
or U2548 (N_2548,In_2393,In_80);
xor U2549 (N_2549,In_445,In_1791);
nor U2550 (N_2550,In_1110,In_1784);
or U2551 (N_2551,In_299,In_1394);
nand U2552 (N_2552,In_162,In_911);
or U2553 (N_2553,In_1391,In_1979);
or U2554 (N_2554,In_201,In_1279);
and U2555 (N_2555,In_1084,In_1771);
xnor U2556 (N_2556,In_1875,In_1565);
nand U2557 (N_2557,In_484,In_1260);
xnor U2558 (N_2558,In_2023,In_1084);
or U2559 (N_2559,In_2408,In_1043);
xnor U2560 (N_2560,In_1287,In_1125);
and U2561 (N_2561,In_434,In_2194);
or U2562 (N_2562,In_1564,In_2401);
xor U2563 (N_2563,In_397,In_1251);
xnor U2564 (N_2564,In_1848,In_200);
nor U2565 (N_2565,In_2256,In_1747);
and U2566 (N_2566,In_1070,In_72);
or U2567 (N_2567,In_269,In_1219);
and U2568 (N_2568,In_1981,In_1588);
and U2569 (N_2569,In_2277,In_94);
nor U2570 (N_2570,In_499,In_158);
or U2571 (N_2571,In_1785,In_1520);
and U2572 (N_2572,In_2204,In_1842);
or U2573 (N_2573,In_612,In_564);
or U2574 (N_2574,In_2420,In_1084);
nor U2575 (N_2575,In_2065,In_394);
xor U2576 (N_2576,In_1267,In_118);
or U2577 (N_2577,In_1245,In_1418);
nand U2578 (N_2578,In_569,In_1125);
or U2579 (N_2579,In_2318,In_252);
nor U2580 (N_2580,In_1736,In_2041);
nor U2581 (N_2581,In_2479,In_853);
nand U2582 (N_2582,In_2474,In_534);
xor U2583 (N_2583,In_2319,In_743);
xor U2584 (N_2584,In_1114,In_1243);
xor U2585 (N_2585,In_1289,In_993);
or U2586 (N_2586,In_1085,In_711);
nor U2587 (N_2587,In_678,In_602);
xnor U2588 (N_2588,In_1275,In_1686);
xnor U2589 (N_2589,In_911,In_551);
or U2590 (N_2590,In_435,In_2324);
nor U2591 (N_2591,In_824,In_1674);
nor U2592 (N_2592,In_677,In_2380);
nand U2593 (N_2593,In_220,In_689);
xnor U2594 (N_2594,In_2201,In_513);
nand U2595 (N_2595,In_2100,In_2498);
xnor U2596 (N_2596,In_386,In_587);
and U2597 (N_2597,In_1827,In_986);
nor U2598 (N_2598,In_2258,In_2426);
nor U2599 (N_2599,In_227,In_1215);
nand U2600 (N_2600,In_594,In_2398);
or U2601 (N_2601,In_224,In_1536);
xnor U2602 (N_2602,In_1993,In_1711);
or U2603 (N_2603,In_1604,In_2467);
or U2604 (N_2604,In_259,In_371);
or U2605 (N_2605,In_286,In_560);
nand U2606 (N_2606,In_1301,In_2275);
and U2607 (N_2607,In_2117,In_126);
or U2608 (N_2608,In_1837,In_1519);
or U2609 (N_2609,In_888,In_1477);
nand U2610 (N_2610,In_2164,In_2131);
or U2611 (N_2611,In_1104,In_2195);
and U2612 (N_2612,In_656,In_1863);
or U2613 (N_2613,In_1069,In_846);
or U2614 (N_2614,In_1333,In_34);
nand U2615 (N_2615,In_1737,In_727);
nor U2616 (N_2616,In_313,In_627);
nand U2617 (N_2617,In_21,In_1337);
nand U2618 (N_2618,In_1535,In_398);
nand U2619 (N_2619,In_617,In_2177);
and U2620 (N_2620,In_1939,In_798);
and U2621 (N_2621,In_893,In_915);
nor U2622 (N_2622,In_5,In_1744);
and U2623 (N_2623,In_2339,In_1047);
nor U2624 (N_2624,In_2243,In_2458);
xor U2625 (N_2625,In_1231,In_2274);
and U2626 (N_2626,In_712,In_193);
or U2627 (N_2627,In_2498,In_1307);
or U2628 (N_2628,In_366,In_161);
nand U2629 (N_2629,In_889,In_2137);
xor U2630 (N_2630,In_408,In_1641);
nor U2631 (N_2631,In_1622,In_190);
nor U2632 (N_2632,In_2328,In_2288);
nor U2633 (N_2633,In_1009,In_992);
nand U2634 (N_2634,In_2444,In_572);
and U2635 (N_2635,In_1394,In_1778);
nor U2636 (N_2636,In_1703,In_0);
and U2637 (N_2637,In_477,In_1885);
nand U2638 (N_2638,In_1548,In_2099);
or U2639 (N_2639,In_310,In_104);
or U2640 (N_2640,In_576,In_768);
xnor U2641 (N_2641,In_1027,In_1679);
or U2642 (N_2642,In_1065,In_1528);
xor U2643 (N_2643,In_182,In_1055);
xnor U2644 (N_2644,In_926,In_438);
xor U2645 (N_2645,In_2315,In_641);
nand U2646 (N_2646,In_2489,In_2248);
and U2647 (N_2647,In_476,In_1889);
and U2648 (N_2648,In_1867,In_894);
or U2649 (N_2649,In_2205,In_150);
xnor U2650 (N_2650,In_1215,In_1218);
or U2651 (N_2651,In_1085,In_687);
nand U2652 (N_2652,In_1120,In_936);
nor U2653 (N_2653,In_1733,In_1588);
and U2654 (N_2654,In_1381,In_2473);
nand U2655 (N_2655,In_1561,In_1913);
and U2656 (N_2656,In_456,In_1398);
nor U2657 (N_2657,In_1284,In_608);
nand U2658 (N_2658,In_2244,In_110);
and U2659 (N_2659,In_777,In_303);
nor U2660 (N_2660,In_1497,In_659);
nand U2661 (N_2661,In_642,In_1979);
xor U2662 (N_2662,In_1984,In_1694);
or U2663 (N_2663,In_1383,In_2109);
nand U2664 (N_2664,In_691,In_775);
nand U2665 (N_2665,In_2159,In_1509);
and U2666 (N_2666,In_634,In_533);
nor U2667 (N_2667,In_2056,In_833);
or U2668 (N_2668,In_1584,In_1278);
xor U2669 (N_2669,In_1726,In_1896);
nand U2670 (N_2670,In_1150,In_394);
or U2671 (N_2671,In_2151,In_2087);
nand U2672 (N_2672,In_2133,In_631);
nand U2673 (N_2673,In_431,In_1855);
xor U2674 (N_2674,In_2011,In_463);
xnor U2675 (N_2675,In_481,In_1708);
and U2676 (N_2676,In_1858,In_549);
nand U2677 (N_2677,In_1335,In_666);
nand U2678 (N_2678,In_1249,In_2425);
nand U2679 (N_2679,In_1401,In_1867);
or U2680 (N_2680,In_2120,In_759);
and U2681 (N_2681,In_138,In_2472);
and U2682 (N_2682,In_1828,In_1057);
nand U2683 (N_2683,In_1734,In_1329);
or U2684 (N_2684,In_815,In_1578);
xor U2685 (N_2685,In_1599,In_1523);
xnor U2686 (N_2686,In_451,In_332);
and U2687 (N_2687,In_1356,In_2192);
xor U2688 (N_2688,In_1904,In_250);
or U2689 (N_2689,In_2082,In_1553);
and U2690 (N_2690,In_2431,In_436);
and U2691 (N_2691,In_2462,In_18);
or U2692 (N_2692,In_2084,In_163);
xnor U2693 (N_2693,In_1197,In_1140);
nand U2694 (N_2694,In_108,In_2036);
nand U2695 (N_2695,In_10,In_1334);
nand U2696 (N_2696,In_1028,In_2056);
or U2697 (N_2697,In_961,In_2313);
or U2698 (N_2698,In_642,In_566);
and U2699 (N_2699,In_241,In_927);
and U2700 (N_2700,In_1879,In_820);
nor U2701 (N_2701,In_198,In_17);
or U2702 (N_2702,In_84,In_967);
and U2703 (N_2703,In_1744,In_1549);
or U2704 (N_2704,In_2248,In_964);
xnor U2705 (N_2705,In_1678,In_1948);
and U2706 (N_2706,In_309,In_1988);
nor U2707 (N_2707,In_672,In_100);
and U2708 (N_2708,In_1709,In_2005);
and U2709 (N_2709,In_328,In_1616);
xor U2710 (N_2710,In_1578,In_2396);
and U2711 (N_2711,In_11,In_454);
xor U2712 (N_2712,In_121,In_1373);
nand U2713 (N_2713,In_1188,In_2388);
xnor U2714 (N_2714,In_2284,In_236);
or U2715 (N_2715,In_1348,In_1684);
and U2716 (N_2716,In_2234,In_1135);
xor U2717 (N_2717,In_1628,In_2158);
and U2718 (N_2718,In_116,In_2272);
nor U2719 (N_2719,In_1818,In_1898);
nand U2720 (N_2720,In_2077,In_76);
nand U2721 (N_2721,In_1437,In_848);
nor U2722 (N_2722,In_2210,In_189);
nor U2723 (N_2723,In_1967,In_2261);
and U2724 (N_2724,In_1670,In_2417);
xor U2725 (N_2725,In_2424,In_635);
nand U2726 (N_2726,In_2417,In_2197);
nor U2727 (N_2727,In_104,In_398);
xor U2728 (N_2728,In_1034,In_1236);
xor U2729 (N_2729,In_483,In_1677);
and U2730 (N_2730,In_1911,In_52);
or U2731 (N_2731,In_1195,In_1666);
xnor U2732 (N_2732,In_1387,In_2427);
and U2733 (N_2733,In_1060,In_874);
nand U2734 (N_2734,In_1662,In_965);
nor U2735 (N_2735,In_38,In_1563);
nor U2736 (N_2736,In_2044,In_310);
nand U2737 (N_2737,In_96,In_1651);
and U2738 (N_2738,In_846,In_673);
and U2739 (N_2739,In_1211,In_2335);
or U2740 (N_2740,In_281,In_595);
or U2741 (N_2741,In_291,In_417);
or U2742 (N_2742,In_2397,In_1033);
xor U2743 (N_2743,In_1782,In_335);
and U2744 (N_2744,In_2110,In_1252);
nor U2745 (N_2745,In_662,In_2145);
nand U2746 (N_2746,In_2368,In_292);
and U2747 (N_2747,In_1256,In_2464);
nand U2748 (N_2748,In_1135,In_342);
or U2749 (N_2749,In_1707,In_2171);
or U2750 (N_2750,In_992,In_501);
or U2751 (N_2751,In_267,In_639);
or U2752 (N_2752,In_454,In_1071);
or U2753 (N_2753,In_256,In_1026);
nor U2754 (N_2754,In_1637,In_1157);
and U2755 (N_2755,In_1485,In_1988);
and U2756 (N_2756,In_2282,In_113);
xnor U2757 (N_2757,In_2210,In_37);
or U2758 (N_2758,In_156,In_1118);
nor U2759 (N_2759,In_2093,In_377);
xnor U2760 (N_2760,In_2416,In_477);
nand U2761 (N_2761,In_667,In_1998);
xnor U2762 (N_2762,In_168,In_1180);
nand U2763 (N_2763,In_1080,In_2391);
xor U2764 (N_2764,In_355,In_900);
xor U2765 (N_2765,In_1555,In_2168);
and U2766 (N_2766,In_1192,In_968);
xnor U2767 (N_2767,In_843,In_380);
and U2768 (N_2768,In_2260,In_1912);
or U2769 (N_2769,In_1874,In_967);
or U2770 (N_2770,In_1306,In_556);
and U2771 (N_2771,In_1934,In_2300);
and U2772 (N_2772,In_1274,In_1646);
nand U2773 (N_2773,In_2457,In_454);
nor U2774 (N_2774,In_664,In_487);
or U2775 (N_2775,In_2003,In_1255);
and U2776 (N_2776,In_1904,In_1069);
and U2777 (N_2777,In_901,In_1269);
nor U2778 (N_2778,In_2246,In_2139);
xor U2779 (N_2779,In_356,In_2455);
and U2780 (N_2780,In_809,In_1778);
xnor U2781 (N_2781,In_169,In_1793);
xnor U2782 (N_2782,In_2098,In_1640);
xnor U2783 (N_2783,In_2421,In_1973);
nor U2784 (N_2784,In_2273,In_1711);
and U2785 (N_2785,In_1946,In_768);
or U2786 (N_2786,In_503,In_627);
or U2787 (N_2787,In_1565,In_2472);
nor U2788 (N_2788,In_2214,In_1580);
nor U2789 (N_2789,In_432,In_90);
xor U2790 (N_2790,In_2033,In_1109);
or U2791 (N_2791,In_2291,In_2013);
or U2792 (N_2792,In_800,In_2490);
or U2793 (N_2793,In_207,In_319);
or U2794 (N_2794,In_2338,In_277);
or U2795 (N_2795,In_13,In_1166);
or U2796 (N_2796,In_2333,In_1308);
nand U2797 (N_2797,In_952,In_2000);
xor U2798 (N_2798,In_1403,In_2287);
nand U2799 (N_2799,In_505,In_110);
xnor U2800 (N_2800,In_1364,In_320);
and U2801 (N_2801,In_1258,In_1689);
xor U2802 (N_2802,In_74,In_631);
nand U2803 (N_2803,In_428,In_133);
nand U2804 (N_2804,In_970,In_399);
and U2805 (N_2805,In_2436,In_1902);
xnor U2806 (N_2806,In_543,In_1440);
xor U2807 (N_2807,In_2442,In_1089);
and U2808 (N_2808,In_2067,In_420);
nor U2809 (N_2809,In_498,In_1657);
and U2810 (N_2810,In_1641,In_728);
xnor U2811 (N_2811,In_1803,In_2263);
xnor U2812 (N_2812,In_1877,In_1629);
xor U2813 (N_2813,In_962,In_1850);
nor U2814 (N_2814,In_2381,In_1276);
or U2815 (N_2815,In_1889,In_1864);
and U2816 (N_2816,In_2352,In_1718);
or U2817 (N_2817,In_977,In_888);
and U2818 (N_2818,In_1251,In_793);
xor U2819 (N_2819,In_784,In_1445);
xnor U2820 (N_2820,In_2052,In_601);
nor U2821 (N_2821,In_773,In_1539);
nand U2822 (N_2822,In_770,In_2367);
nand U2823 (N_2823,In_1506,In_1155);
xnor U2824 (N_2824,In_392,In_2372);
nor U2825 (N_2825,In_554,In_2160);
nor U2826 (N_2826,In_1106,In_2115);
nor U2827 (N_2827,In_1510,In_941);
nor U2828 (N_2828,In_29,In_1651);
nor U2829 (N_2829,In_2179,In_246);
xnor U2830 (N_2830,In_467,In_232);
or U2831 (N_2831,In_2004,In_1592);
nand U2832 (N_2832,In_1716,In_66);
or U2833 (N_2833,In_350,In_1468);
xor U2834 (N_2834,In_1403,In_1013);
xnor U2835 (N_2835,In_285,In_82);
or U2836 (N_2836,In_1018,In_1874);
nor U2837 (N_2837,In_1783,In_556);
nor U2838 (N_2838,In_1369,In_590);
nor U2839 (N_2839,In_1154,In_1720);
and U2840 (N_2840,In_896,In_10);
nand U2841 (N_2841,In_1514,In_1101);
nand U2842 (N_2842,In_1966,In_2349);
nor U2843 (N_2843,In_200,In_497);
nand U2844 (N_2844,In_1336,In_1348);
nand U2845 (N_2845,In_1525,In_1816);
nor U2846 (N_2846,In_364,In_111);
nand U2847 (N_2847,In_20,In_813);
and U2848 (N_2848,In_149,In_9);
and U2849 (N_2849,In_784,In_596);
and U2850 (N_2850,In_301,In_21);
nor U2851 (N_2851,In_2386,In_1588);
xnor U2852 (N_2852,In_1021,In_546);
or U2853 (N_2853,In_899,In_1595);
nand U2854 (N_2854,In_2173,In_1271);
and U2855 (N_2855,In_2464,In_756);
or U2856 (N_2856,In_899,In_1926);
xor U2857 (N_2857,In_1037,In_382);
or U2858 (N_2858,In_995,In_938);
and U2859 (N_2859,In_1500,In_1350);
xor U2860 (N_2860,In_2134,In_2449);
and U2861 (N_2861,In_64,In_390);
nor U2862 (N_2862,In_492,In_2257);
nand U2863 (N_2863,In_2077,In_407);
nand U2864 (N_2864,In_1275,In_328);
nand U2865 (N_2865,In_2204,In_2375);
or U2866 (N_2866,In_166,In_2079);
xnor U2867 (N_2867,In_837,In_1827);
or U2868 (N_2868,In_1254,In_1597);
xor U2869 (N_2869,In_2005,In_1295);
and U2870 (N_2870,In_1483,In_1135);
nand U2871 (N_2871,In_361,In_847);
xnor U2872 (N_2872,In_1042,In_418);
xnor U2873 (N_2873,In_2027,In_1535);
nand U2874 (N_2874,In_2067,In_1898);
and U2875 (N_2875,In_1602,In_1978);
nand U2876 (N_2876,In_1450,In_1147);
nand U2877 (N_2877,In_298,In_2419);
nand U2878 (N_2878,In_961,In_1017);
or U2879 (N_2879,In_2457,In_107);
nand U2880 (N_2880,In_1710,In_1001);
and U2881 (N_2881,In_570,In_1105);
nor U2882 (N_2882,In_73,In_511);
or U2883 (N_2883,In_1057,In_1022);
and U2884 (N_2884,In_2367,In_37);
nor U2885 (N_2885,In_1876,In_1049);
and U2886 (N_2886,In_53,In_1094);
and U2887 (N_2887,In_312,In_1522);
nand U2888 (N_2888,In_885,In_800);
nand U2889 (N_2889,In_338,In_1618);
nor U2890 (N_2890,In_241,In_1509);
nand U2891 (N_2891,In_2274,In_1842);
nand U2892 (N_2892,In_554,In_1515);
nor U2893 (N_2893,In_78,In_1794);
and U2894 (N_2894,In_486,In_579);
nor U2895 (N_2895,In_1647,In_1218);
nor U2896 (N_2896,In_1880,In_1541);
or U2897 (N_2897,In_869,In_1151);
or U2898 (N_2898,In_247,In_1135);
nand U2899 (N_2899,In_577,In_1867);
or U2900 (N_2900,In_1173,In_189);
xnor U2901 (N_2901,In_99,In_1248);
nand U2902 (N_2902,In_1858,In_1396);
nand U2903 (N_2903,In_2127,In_860);
xor U2904 (N_2904,In_1580,In_2162);
and U2905 (N_2905,In_104,In_2099);
and U2906 (N_2906,In_510,In_1499);
and U2907 (N_2907,In_814,In_1349);
or U2908 (N_2908,In_1384,In_236);
xor U2909 (N_2909,In_544,In_2392);
and U2910 (N_2910,In_1553,In_18);
nand U2911 (N_2911,In_1785,In_1010);
or U2912 (N_2912,In_420,In_1826);
nand U2913 (N_2913,In_395,In_642);
and U2914 (N_2914,In_582,In_576);
nor U2915 (N_2915,In_1431,In_1661);
nand U2916 (N_2916,In_2327,In_259);
nor U2917 (N_2917,In_579,In_2162);
or U2918 (N_2918,In_1975,In_1159);
and U2919 (N_2919,In_2250,In_1058);
and U2920 (N_2920,In_531,In_2197);
nor U2921 (N_2921,In_492,In_311);
xor U2922 (N_2922,In_2456,In_337);
xor U2923 (N_2923,In_358,In_1979);
nor U2924 (N_2924,In_408,In_2442);
and U2925 (N_2925,In_349,In_1541);
and U2926 (N_2926,In_361,In_1969);
xor U2927 (N_2927,In_441,In_724);
nand U2928 (N_2928,In_1564,In_2354);
and U2929 (N_2929,In_1136,In_1119);
or U2930 (N_2930,In_2044,In_1675);
and U2931 (N_2931,In_1979,In_1005);
and U2932 (N_2932,In_2361,In_275);
nand U2933 (N_2933,In_433,In_2442);
or U2934 (N_2934,In_2418,In_461);
nand U2935 (N_2935,In_1167,In_1726);
nor U2936 (N_2936,In_1335,In_104);
xor U2937 (N_2937,In_293,In_1862);
nand U2938 (N_2938,In_2407,In_2071);
nor U2939 (N_2939,In_2429,In_97);
or U2940 (N_2940,In_1189,In_1779);
nor U2941 (N_2941,In_370,In_1377);
xnor U2942 (N_2942,In_2438,In_631);
xor U2943 (N_2943,In_1467,In_964);
and U2944 (N_2944,In_48,In_1508);
and U2945 (N_2945,In_181,In_1165);
and U2946 (N_2946,In_868,In_2015);
xnor U2947 (N_2947,In_925,In_231);
or U2948 (N_2948,In_2276,In_1381);
and U2949 (N_2949,In_541,In_1831);
nor U2950 (N_2950,In_2123,In_289);
nand U2951 (N_2951,In_1087,In_438);
and U2952 (N_2952,In_1409,In_1065);
xor U2953 (N_2953,In_935,In_864);
nand U2954 (N_2954,In_895,In_716);
nor U2955 (N_2955,In_1637,In_1260);
or U2956 (N_2956,In_1506,In_77);
nand U2957 (N_2957,In_1751,In_1446);
nor U2958 (N_2958,In_605,In_1558);
or U2959 (N_2959,In_989,In_1783);
and U2960 (N_2960,In_2064,In_184);
and U2961 (N_2961,In_44,In_1032);
nand U2962 (N_2962,In_1904,In_50);
and U2963 (N_2963,In_642,In_498);
and U2964 (N_2964,In_615,In_666);
xor U2965 (N_2965,In_1395,In_195);
or U2966 (N_2966,In_815,In_2151);
or U2967 (N_2967,In_1569,In_2286);
nand U2968 (N_2968,In_386,In_968);
or U2969 (N_2969,In_525,In_2286);
nor U2970 (N_2970,In_1233,In_215);
nor U2971 (N_2971,In_2203,In_1769);
nand U2972 (N_2972,In_2067,In_572);
and U2973 (N_2973,In_399,In_1828);
xnor U2974 (N_2974,In_2439,In_291);
xor U2975 (N_2975,In_1091,In_2426);
and U2976 (N_2976,In_2212,In_408);
xor U2977 (N_2977,In_1605,In_376);
and U2978 (N_2978,In_1672,In_303);
nor U2979 (N_2979,In_1691,In_1129);
or U2980 (N_2980,In_30,In_1228);
xnor U2981 (N_2981,In_2419,In_1995);
and U2982 (N_2982,In_2052,In_2034);
xnor U2983 (N_2983,In_448,In_1529);
or U2984 (N_2984,In_634,In_1463);
nor U2985 (N_2985,In_830,In_1209);
xor U2986 (N_2986,In_2466,In_1634);
or U2987 (N_2987,In_275,In_1804);
or U2988 (N_2988,In_2455,In_1513);
and U2989 (N_2989,In_974,In_305);
xnor U2990 (N_2990,In_1235,In_2238);
and U2991 (N_2991,In_283,In_11);
xnor U2992 (N_2992,In_1805,In_328);
nor U2993 (N_2993,In_2093,In_1314);
and U2994 (N_2994,In_2076,In_1444);
xor U2995 (N_2995,In_1191,In_194);
or U2996 (N_2996,In_2191,In_169);
xnor U2997 (N_2997,In_1845,In_1503);
nand U2998 (N_2998,In_1277,In_2007);
nor U2999 (N_2999,In_1691,In_50);
and U3000 (N_3000,In_1744,In_1713);
nand U3001 (N_3001,In_1110,In_768);
nand U3002 (N_3002,In_757,In_481);
nor U3003 (N_3003,In_2420,In_1125);
nor U3004 (N_3004,In_476,In_900);
xnor U3005 (N_3005,In_2108,In_543);
or U3006 (N_3006,In_653,In_2225);
and U3007 (N_3007,In_2175,In_1185);
nand U3008 (N_3008,In_93,In_359);
and U3009 (N_3009,In_1633,In_1359);
or U3010 (N_3010,In_1134,In_2460);
xor U3011 (N_3011,In_577,In_571);
nor U3012 (N_3012,In_94,In_277);
and U3013 (N_3013,In_483,In_1186);
or U3014 (N_3014,In_1134,In_1137);
xor U3015 (N_3015,In_549,In_547);
and U3016 (N_3016,In_2056,In_1985);
xnor U3017 (N_3017,In_1964,In_2130);
or U3018 (N_3018,In_65,In_2252);
nand U3019 (N_3019,In_613,In_680);
nand U3020 (N_3020,In_1201,In_273);
or U3021 (N_3021,In_2379,In_727);
and U3022 (N_3022,In_1082,In_1830);
nand U3023 (N_3023,In_1313,In_1585);
nor U3024 (N_3024,In_2487,In_1971);
or U3025 (N_3025,In_2384,In_748);
xnor U3026 (N_3026,In_1368,In_797);
and U3027 (N_3027,In_1164,In_1964);
nor U3028 (N_3028,In_906,In_856);
or U3029 (N_3029,In_1829,In_169);
xor U3030 (N_3030,In_2137,In_1561);
or U3031 (N_3031,In_427,In_1061);
and U3032 (N_3032,In_208,In_2220);
xnor U3033 (N_3033,In_1953,In_1995);
nor U3034 (N_3034,In_1193,In_2039);
and U3035 (N_3035,In_2192,In_1541);
or U3036 (N_3036,In_104,In_2415);
or U3037 (N_3037,In_640,In_1336);
or U3038 (N_3038,In_2439,In_771);
xnor U3039 (N_3039,In_1081,In_1920);
xor U3040 (N_3040,In_545,In_1574);
nor U3041 (N_3041,In_497,In_1924);
nor U3042 (N_3042,In_2483,In_1605);
or U3043 (N_3043,In_1782,In_1064);
nand U3044 (N_3044,In_949,In_2297);
xor U3045 (N_3045,In_867,In_1831);
nand U3046 (N_3046,In_1060,In_2291);
or U3047 (N_3047,In_2354,In_2047);
nor U3048 (N_3048,In_1374,In_924);
nand U3049 (N_3049,In_398,In_1125);
nor U3050 (N_3050,In_336,In_2259);
nor U3051 (N_3051,In_212,In_379);
nor U3052 (N_3052,In_493,In_1810);
xnor U3053 (N_3053,In_806,In_981);
or U3054 (N_3054,In_1376,In_958);
or U3055 (N_3055,In_1092,In_1987);
nor U3056 (N_3056,In_1139,In_1123);
or U3057 (N_3057,In_2275,In_1640);
nor U3058 (N_3058,In_1076,In_2227);
nor U3059 (N_3059,In_1506,In_2119);
nand U3060 (N_3060,In_1243,In_796);
xor U3061 (N_3061,In_2174,In_678);
nor U3062 (N_3062,In_238,In_1084);
and U3063 (N_3063,In_909,In_2228);
or U3064 (N_3064,In_2169,In_1171);
xor U3065 (N_3065,In_597,In_107);
and U3066 (N_3066,In_475,In_1584);
nor U3067 (N_3067,In_791,In_2250);
and U3068 (N_3068,In_708,In_1856);
nor U3069 (N_3069,In_514,In_285);
nor U3070 (N_3070,In_209,In_941);
or U3071 (N_3071,In_1879,In_792);
xnor U3072 (N_3072,In_131,In_1119);
nand U3073 (N_3073,In_2266,In_1413);
nor U3074 (N_3074,In_740,In_211);
or U3075 (N_3075,In_1994,In_1235);
nand U3076 (N_3076,In_56,In_1263);
nor U3077 (N_3077,In_1222,In_2120);
nor U3078 (N_3078,In_971,In_2069);
or U3079 (N_3079,In_588,In_1348);
nand U3080 (N_3080,In_24,In_164);
nor U3081 (N_3081,In_1583,In_2030);
or U3082 (N_3082,In_195,In_1109);
and U3083 (N_3083,In_941,In_1842);
nor U3084 (N_3084,In_1287,In_566);
nor U3085 (N_3085,In_303,In_1950);
or U3086 (N_3086,In_128,In_1328);
nor U3087 (N_3087,In_681,In_438);
xor U3088 (N_3088,In_348,In_2051);
nand U3089 (N_3089,In_426,In_1283);
and U3090 (N_3090,In_2415,In_2168);
nand U3091 (N_3091,In_965,In_1788);
or U3092 (N_3092,In_1706,In_1936);
nor U3093 (N_3093,In_1985,In_1825);
and U3094 (N_3094,In_950,In_1918);
xor U3095 (N_3095,In_1805,In_1601);
or U3096 (N_3096,In_867,In_127);
nor U3097 (N_3097,In_1776,In_870);
xor U3098 (N_3098,In_898,In_1086);
nor U3099 (N_3099,In_2164,In_1389);
nand U3100 (N_3100,In_157,In_1881);
nand U3101 (N_3101,In_441,In_11);
or U3102 (N_3102,In_2437,In_562);
nand U3103 (N_3103,In_1297,In_1507);
nor U3104 (N_3104,In_1257,In_2177);
nand U3105 (N_3105,In_1067,In_575);
or U3106 (N_3106,In_287,In_205);
nor U3107 (N_3107,In_521,In_540);
xor U3108 (N_3108,In_2452,In_1574);
nor U3109 (N_3109,In_1761,In_437);
or U3110 (N_3110,In_2142,In_2066);
nor U3111 (N_3111,In_1562,In_2303);
nor U3112 (N_3112,In_768,In_289);
and U3113 (N_3113,In_27,In_842);
or U3114 (N_3114,In_1122,In_1378);
nand U3115 (N_3115,In_2118,In_2084);
xnor U3116 (N_3116,In_1064,In_1474);
or U3117 (N_3117,In_2390,In_1857);
and U3118 (N_3118,In_2203,In_1466);
nand U3119 (N_3119,In_871,In_2151);
nand U3120 (N_3120,In_1083,In_229);
nand U3121 (N_3121,In_2065,In_1510);
nand U3122 (N_3122,In_1796,In_1277);
nor U3123 (N_3123,In_908,In_423);
and U3124 (N_3124,In_384,In_1263);
and U3125 (N_3125,In_1535,In_2249);
nand U3126 (N_3126,In_202,In_717);
nor U3127 (N_3127,In_2096,In_729);
nand U3128 (N_3128,In_1550,In_1049);
and U3129 (N_3129,In_2314,In_898);
nand U3130 (N_3130,In_1807,In_1729);
nand U3131 (N_3131,In_425,In_2184);
nor U3132 (N_3132,In_13,In_1342);
nand U3133 (N_3133,In_1467,In_639);
or U3134 (N_3134,In_1483,In_193);
nor U3135 (N_3135,In_1439,In_1468);
or U3136 (N_3136,In_1239,In_1139);
nor U3137 (N_3137,In_402,In_1635);
nor U3138 (N_3138,In_1668,In_850);
nand U3139 (N_3139,In_2150,In_2216);
and U3140 (N_3140,In_1685,In_2191);
or U3141 (N_3141,In_475,In_239);
and U3142 (N_3142,In_1978,In_94);
or U3143 (N_3143,In_1511,In_2496);
and U3144 (N_3144,In_1205,In_2236);
or U3145 (N_3145,In_135,In_266);
or U3146 (N_3146,In_1799,In_1554);
nor U3147 (N_3147,In_1321,In_1124);
nor U3148 (N_3148,In_2495,In_1798);
nand U3149 (N_3149,In_2476,In_1880);
and U3150 (N_3150,In_765,In_1110);
nand U3151 (N_3151,In_384,In_956);
nand U3152 (N_3152,In_1141,In_1603);
nand U3153 (N_3153,In_1577,In_1329);
or U3154 (N_3154,In_595,In_1937);
nor U3155 (N_3155,In_1815,In_731);
and U3156 (N_3156,In_114,In_490);
nand U3157 (N_3157,In_517,In_2346);
nor U3158 (N_3158,In_1724,In_780);
xor U3159 (N_3159,In_938,In_2274);
or U3160 (N_3160,In_345,In_277);
xor U3161 (N_3161,In_784,In_1280);
nand U3162 (N_3162,In_1663,In_1016);
xnor U3163 (N_3163,In_2111,In_2339);
nor U3164 (N_3164,In_202,In_1795);
and U3165 (N_3165,In_1847,In_1914);
xnor U3166 (N_3166,In_1979,In_1661);
and U3167 (N_3167,In_1535,In_2329);
or U3168 (N_3168,In_790,In_1535);
or U3169 (N_3169,In_680,In_2097);
nand U3170 (N_3170,In_1145,In_323);
nand U3171 (N_3171,In_1424,In_1675);
and U3172 (N_3172,In_2019,In_2237);
and U3173 (N_3173,In_10,In_912);
or U3174 (N_3174,In_1915,In_1150);
nor U3175 (N_3175,In_323,In_262);
xor U3176 (N_3176,In_1220,In_1628);
xnor U3177 (N_3177,In_905,In_1394);
nor U3178 (N_3178,In_67,In_1232);
nand U3179 (N_3179,In_2000,In_1408);
nand U3180 (N_3180,In_2316,In_337);
and U3181 (N_3181,In_2253,In_1286);
and U3182 (N_3182,In_1129,In_1912);
nand U3183 (N_3183,In_1213,In_56);
nor U3184 (N_3184,In_2288,In_2255);
nor U3185 (N_3185,In_1012,In_1967);
or U3186 (N_3186,In_1771,In_1211);
nor U3187 (N_3187,In_1577,In_1364);
xnor U3188 (N_3188,In_308,In_331);
nand U3189 (N_3189,In_2418,In_340);
and U3190 (N_3190,In_1253,In_2281);
nand U3191 (N_3191,In_2063,In_1760);
and U3192 (N_3192,In_1505,In_532);
xor U3193 (N_3193,In_1819,In_1004);
nand U3194 (N_3194,In_1538,In_1499);
xnor U3195 (N_3195,In_2456,In_1744);
or U3196 (N_3196,In_926,In_1311);
nor U3197 (N_3197,In_1247,In_812);
nand U3198 (N_3198,In_543,In_91);
nor U3199 (N_3199,In_416,In_1697);
nand U3200 (N_3200,In_741,In_2050);
xor U3201 (N_3201,In_1744,In_2343);
and U3202 (N_3202,In_39,In_844);
or U3203 (N_3203,In_1145,In_1888);
nor U3204 (N_3204,In_884,In_810);
xnor U3205 (N_3205,In_1630,In_2301);
nand U3206 (N_3206,In_1591,In_1);
or U3207 (N_3207,In_709,In_1495);
and U3208 (N_3208,In_1747,In_431);
nor U3209 (N_3209,In_1059,In_357);
or U3210 (N_3210,In_1782,In_1593);
nor U3211 (N_3211,In_1540,In_1972);
xnor U3212 (N_3212,In_504,In_1981);
nor U3213 (N_3213,In_2333,In_675);
xor U3214 (N_3214,In_1996,In_2151);
nand U3215 (N_3215,In_1067,In_1557);
and U3216 (N_3216,In_34,In_19);
or U3217 (N_3217,In_64,In_2336);
and U3218 (N_3218,In_129,In_2294);
nor U3219 (N_3219,In_522,In_1386);
nor U3220 (N_3220,In_1590,In_472);
nand U3221 (N_3221,In_1028,In_1006);
and U3222 (N_3222,In_181,In_665);
and U3223 (N_3223,In_470,In_274);
nor U3224 (N_3224,In_2276,In_508);
and U3225 (N_3225,In_223,In_881);
nand U3226 (N_3226,In_619,In_1117);
and U3227 (N_3227,In_1977,In_489);
nor U3228 (N_3228,In_884,In_2284);
and U3229 (N_3229,In_2103,In_977);
xnor U3230 (N_3230,In_2478,In_644);
nor U3231 (N_3231,In_1618,In_89);
and U3232 (N_3232,In_55,In_373);
or U3233 (N_3233,In_2039,In_727);
and U3234 (N_3234,In_634,In_317);
nor U3235 (N_3235,In_2255,In_1414);
or U3236 (N_3236,In_1748,In_1824);
nand U3237 (N_3237,In_1844,In_1537);
and U3238 (N_3238,In_82,In_2430);
and U3239 (N_3239,In_2108,In_1039);
or U3240 (N_3240,In_1832,In_1801);
xnor U3241 (N_3241,In_1552,In_785);
nand U3242 (N_3242,In_1796,In_1318);
nor U3243 (N_3243,In_2179,In_2355);
nor U3244 (N_3244,In_2472,In_1501);
nand U3245 (N_3245,In_1581,In_2182);
nand U3246 (N_3246,In_395,In_1952);
and U3247 (N_3247,In_56,In_1901);
xnor U3248 (N_3248,In_2237,In_931);
xor U3249 (N_3249,In_803,In_1293);
nand U3250 (N_3250,In_2400,In_1617);
or U3251 (N_3251,In_1290,In_1553);
xnor U3252 (N_3252,In_2368,In_42);
and U3253 (N_3253,In_541,In_1886);
nand U3254 (N_3254,In_1066,In_1656);
nor U3255 (N_3255,In_13,In_1439);
nor U3256 (N_3256,In_425,In_933);
nor U3257 (N_3257,In_347,In_427);
xor U3258 (N_3258,In_1128,In_758);
nor U3259 (N_3259,In_1908,In_1544);
xor U3260 (N_3260,In_2395,In_1717);
nor U3261 (N_3261,In_1083,In_877);
and U3262 (N_3262,In_2419,In_947);
xor U3263 (N_3263,In_1730,In_136);
nor U3264 (N_3264,In_153,In_165);
nand U3265 (N_3265,In_936,In_452);
and U3266 (N_3266,In_153,In_1173);
nand U3267 (N_3267,In_932,In_1048);
or U3268 (N_3268,In_1896,In_1575);
and U3269 (N_3269,In_667,In_431);
or U3270 (N_3270,In_2175,In_2278);
or U3271 (N_3271,In_211,In_4);
and U3272 (N_3272,In_865,In_690);
or U3273 (N_3273,In_586,In_894);
and U3274 (N_3274,In_1257,In_920);
nand U3275 (N_3275,In_2111,In_2081);
and U3276 (N_3276,In_2114,In_156);
nor U3277 (N_3277,In_1162,In_2088);
xor U3278 (N_3278,In_2078,In_947);
or U3279 (N_3279,In_1765,In_724);
xnor U3280 (N_3280,In_941,In_435);
xor U3281 (N_3281,In_1636,In_2379);
nor U3282 (N_3282,In_1657,In_999);
or U3283 (N_3283,In_1601,In_1447);
xor U3284 (N_3284,In_928,In_2000);
nor U3285 (N_3285,In_1086,In_1996);
nand U3286 (N_3286,In_2162,In_2328);
xor U3287 (N_3287,In_921,In_1356);
nand U3288 (N_3288,In_320,In_1731);
or U3289 (N_3289,In_2087,In_2170);
and U3290 (N_3290,In_383,In_973);
nand U3291 (N_3291,In_2494,In_91);
nor U3292 (N_3292,In_560,In_1376);
and U3293 (N_3293,In_1133,In_842);
xor U3294 (N_3294,In_113,In_703);
nor U3295 (N_3295,In_347,In_429);
nand U3296 (N_3296,In_1396,In_2473);
and U3297 (N_3297,In_2311,In_1973);
or U3298 (N_3298,In_595,In_459);
nand U3299 (N_3299,In_342,In_2195);
xnor U3300 (N_3300,In_129,In_2327);
nand U3301 (N_3301,In_2025,In_690);
nand U3302 (N_3302,In_901,In_137);
nand U3303 (N_3303,In_2035,In_1701);
xor U3304 (N_3304,In_657,In_41);
nand U3305 (N_3305,In_1819,In_217);
xor U3306 (N_3306,In_2363,In_118);
xor U3307 (N_3307,In_1456,In_1363);
xnor U3308 (N_3308,In_2143,In_2401);
and U3309 (N_3309,In_1238,In_648);
and U3310 (N_3310,In_527,In_2332);
and U3311 (N_3311,In_634,In_1156);
nor U3312 (N_3312,In_940,In_682);
or U3313 (N_3313,In_1632,In_2277);
xnor U3314 (N_3314,In_1233,In_1580);
nand U3315 (N_3315,In_2288,In_1659);
nand U3316 (N_3316,In_1302,In_2172);
nor U3317 (N_3317,In_844,In_2260);
and U3318 (N_3318,In_2119,In_1754);
xnor U3319 (N_3319,In_772,In_405);
or U3320 (N_3320,In_868,In_548);
nand U3321 (N_3321,In_290,In_1102);
and U3322 (N_3322,In_673,In_162);
nor U3323 (N_3323,In_541,In_1724);
or U3324 (N_3324,In_1338,In_2134);
nand U3325 (N_3325,In_2183,In_2158);
xor U3326 (N_3326,In_629,In_2200);
or U3327 (N_3327,In_1657,In_2254);
xor U3328 (N_3328,In_990,In_1876);
xor U3329 (N_3329,In_198,In_1407);
and U3330 (N_3330,In_764,In_1691);
or U3331 (N_3331,In_1136,In_831);
or U3332 (N_3332,In_1000,In_565);
xnor U3333 (N_3333,In_1261,In_477);
or U3334 (N_3334,In_1425,In_1958);
and U3335 (N_3335,In_1066,In_689);
nand U3336 (N_3336,In_172,In_2096);
nor U3337 (N_3337,In_607,In_2477);
nand U3338 (N_3338,In_870,In_664);
or U3339 (N_3339,In_1134,In_1130);
and U3340 (N_3340,In_1169,In_2027);
and U3341 (N_3341,In_2170,In_657);
and U3342 (N_3342,In_146,In_1766);
and U3343 (N_3343,In_1247,In_440);
xor U3344 (N_3344,In_962,In_9);
and U3345 (N_3345,In_1541,In_321);
xor U3346 (N_3346,In_985,In_2313);
nand U3347 (N_3347,In_1473,In_335);
nor U3348 (N_3348,In_1425,In_471);
and U3349 (N_3349,In_1337,In_255);
nor U3350 (N_3350,In_1663,In_741);
and U3351 (N_3351,In_688,In_2072);
nor U3352 (N_3352,In_524,In_881);
xor U3353 (N_3353,In_907,In_1007);
nor U3354 (N_3354,In_1814,In_1989);
and U3355 (N_3355,In_1345,In_2150);
xnor U3356 (N_3356,In_1947,In_1560);
or U3357 (N_3357,In_1388,In_3);
and U3358 (N_3358,In_468,In_2234);
nand U3359 (N_3359,In_2024,In_1381);
xor U3360 (N_3360,In_1882,In_517);
nand U3361 (N_3361,In_2370,In_1188);
nand U3362 (N_3362,In_1005,In_1228);
and U3363 (N_3363,In_1328,In_2270);
xnor U3364 (N_3364,In_1078,In_1582);
and U3365 (N_3365,In_257,In_1001);
or U3366 (N_3366,In_1770,In_707);
xnor U3367 (N_3367,In_1328,In_1310);
xor U3368 (N_3368,In_1732,In_148);
or U3369 (N_3369,In_2041,In_2096);
xnor U3370 (N_3370,In_2286,In_1913);
nor U3371 (N_3371,In_1440,In_36);
xnor U3372 (N_3372,In_1166,In_993);
and U3373 (N_3373,In_17,In_1754);
and U3374 (N_3374,In_1486,In_1751);
and U3375 (N_3375,In_1527,In_1242);
nor U3376 (N_3376,In_407,In_348);
nand U3377 (N_3377,In_1006,In_588);
nor U3378 (N_3378,In_180,In_2304);
xor U3379 (N_3379,In_44,In_1354);
and U3380 (N_3380,In_633,In_1528);
nand U3381 (N_3381,In_2065,In_1794);
and U3382 (N_3382,In_1479,In_1949);
nand U3383 (N_3383,In_2362,In_1148);
nand U3384 (N_3384,In_683,In_2408);
xnor U3385 (N_3385,In_702,In_159);
nor U3386 (N_3386,In_2066,In_724);
or U3387 (N_3387,In_1026,In_1666);
nand U3388 (N_3388,In_1846,In_1065);
xor U3389 (N_3389,In_81,In_733);
and U3390 (N_3390,In_864,In_1345);
or U3391 (N_3391,In_167,In_1405);
xor U3392 (N_3392,In_2191,In_2182);
nand U3393 (N_3393,In_844,In_1629);
xnor U3394 (N_3394,In_404,In_2357);
nand U3395 (N_3395,In_1125,In_2257);
nor U3396 (N_3396,In_293,In_590);
xor U3397 (N_3397,In_330,In_1958);
and U3398 (N_3398,In_1060,In_1569);
xnor U3399 (N_3399,In_2122,In_1196);
and U3400 (N_3400,In_993,In_1214);
or U3401 (N_3401,In_142,In_853);
xnor U3402 (N_3402,In_2367,In_877);
and U3403 (N_3403,In_89,In_154);
nand U3404 (N_3404,In_2341,In_357);
nor U3405 (N_3405,In_210,In_463);
nand U3406 (N_3406,In_923,In_1502);
nand U3407 (N_3407,In_122,In_548);
nand U3408 (N_3408,In_2098,In_837);
nand U3409 (N_3409,In_41,In_1017);
xnor U3410 (N_3410,In_1291,In_1836);
nor U3411 (N_3411,In_230,In_1214);
xor U3412 (N_3412,In_1970,In_1339);
nand U3413 (N_3413,In_468,In_611);
or U3414 (N_3414,In_420,In_1716);
or U3415 (N_3415,In_306,In_1904);
nand U3416 (N_3416,In_248,In_938);
nand U3417 (N_3417,In_1047,In_1976);
or U3418 (N_3418,In_2044,In_2405);
xor U3419 (N_3419,In_279,In_959);
xnor U3420 (N_3420,In_674,In_1370);
and U3421 (N_3421,In_162,In_172);
nor U3422 (N_3422,In_35,In_767);
xor U3423 (N_3423,In_2117,In_868);
and U3424 (N_3424,In_1883,In_2451);
nor U3425 (N_3425,In_1399,In_991);
or U3426 (N_3426,In_1895,In_2463);
or U3427 (N_3427,In_2337,In_184);
and U3428 (N_3428,In_1977,In_2021);
nand U3429 (N_3429,In_2282,In_2405);
xor U3430 (N_3430,In_286,In_2012);
nor U3431 (N_3431,In_1889,In_1078);
and U3432 (N_3432,In_1807,In_2485);
and U3433 (N_3433,In_1416,In_1015);
xnor U3434 (N_3434,In_1200,In_2123);
and U3435 (N_3435,In_24,In_1400);
nand U3436 (N_3436,In_186,In_1985);
xor U3437 (N_3437,In_17,In_1917);
xnor U3438 (N_3438,In_308,In_65);
xnor U3439 (N_3439,In_188,In_614);
xor U3440 (N_3440,In_2285,In_1357);
or U3441 (N_3441,In_937,In_1893);
nand U3442 (N_3442,In_160,In_1008);
or U3443 (N_3443,In_1547,In_2364);
and U3444 (N_3444,In_967,In_685);
nor U3445 (N_3445,In_217,In_1941);
nor U3446 (N_3446,In_952,In_1640);
nand U3447 (N_3447,In_778,In_1257);
nand U3448 (N_3448,In_1184,In_2269);
xor U3449 (N_3449,In_1456,In_2069);
or U3450 (N_3450,In_2095,In_440);
nor U3451 (N_3451,In_247,In_1131);
nand U3452 (N_3452,In_2059,In_132);
or U3453 (N_3453,In_1503,In_1405);
and U3454 (N_3454,In_1145,In_1011);
xnor U3455 (N_3455,In_250,In_284);
nand U3456 (N_3456,In_2018,In_61);
nor U3457 (N_3457,In_2255,In_2039);
nor U3458 (N_3458,In_1236,In_2470);
nor U3459 (N_3459,In_1529,In_1797);
nand U3460 (N_3460,In_1985,In_1324);
nor U3461 (N_3461,In_2072,In_1855);
nand U3462 (N_3462,In_2130,In_688);
nor U3463 (N_3463,In_1519,In_1916);
or U3464 (N_3464,In_323,In_48);
xor U3465 (N_3465,In_492,In_507);
xnor U3466 (N_3466,In_289,In_2385);
nor U3467 (N_3467,In_397,In_1579);
xor U3468 (N_3468,In_293,In_752);
or U3469 (N_3469,In_1842,In_2283);
and U3470 (N_3470,In_1352,In_2349);
and U3471 (N_3471,In_713,In_387);
nand U3472 (N_3472,In_437,In_1856);
nand U3473 (N_3473,In_744,In_1895);
xnor U3474 (N_3474,In_332,In_1694);
xor U3475 (N_3475,In_576,In_2442);
or U3476 (N_3476,In_397,In_608);
nand U3477 (N_3477,In_2249,In_798);
nand U3478 (N_3478,In_107,In_666);
nand U3479 (N_3479,In_824,In_2061);
nand U3480 (N_3480,In_1849,In_2357);
nor U3481 (N_3481,In_2306,In_2486);
xnor U3482 (N_3482,In_156,In_2425);
nor U3483 (N_3483,In_10,In_252);
and U3484 (N_3484,In_389,In_561);
nand U3485 (N_3485,In_931,In_1296);
xnor U3486 (N_3486,In_12,In_1195);
or U3487 (N_3487,In_5,In_116);
and U3488 (N_3488,In_448,In_908);
and U3489 (N_3489,In_2129,In_1949);
or U3490 (N_3490,In_1872,In_1343);
nor U3491 (N_3491,In_606,In_555);
nor U3492 (N_3492,In_462,In_1672);
or U3493 (N_3493,In_1845,In_2010);
xor U3494 (N_3494,In_1385,In_2094);
nand U3495 (N_3495,In_1652,In_1231);
nand U3496 (N_3496,In_564,In_1042);
nand U3497 (N_3497,In_957,In_2167);
and U3498 (N_3498,In_380,In_1595);
nand U3499 (N_3499,In_951,In_1089);
nor U3500 (N_3500,In_133,In_2437);
xor U3501 (N_3501,In_337,In_2413);
nor U3502 (N_3502,In_808,In_56);
xnor U3503 (N_3503,In_1130,In_164);
and U3504 (N_3504,In_968,In_2257);
and U3505 (N_3505,In_325,In_1794);
and U3506 (N_3506,In_1416,In_867);
or U3507 (N_3507,In_1085,In_239);
and U3508 (N_3508,In_630,In_484);
or U3509 (N_3509,In_164,In_487);
nand U3510 (N_3510,In_1968,In_1954);
nand U3511 (N_3511,In_2184,In_83);
or U3512 (N_3512,In_66,In_1823);
nand U3513 (N_3513,In_1760,In_280);
and U3514 (N_3514,In_719,In_1465);
or U3515 (N_3515,In_1832,In_1078);
nand U3516 (N_3516,In_1844,In_2332);
nand U3517 (N_3517,In_788,In_1178);
and U3518 (N_3518,In_644,In_1324);
xor U3519 (N_3519,In_1004,In_1632);
and U3520 (N_3520,In_1168,In_2086);
and U3521 (N_3521,In_2078,In_861);
nor U3522 (N_3522,In_554,In_409);
or U3523 (N_3523,In_468,In_1670);
xnor U3524 (N_3524,In_2347,In_2062);
xnor U3525 (N_3525,In_1609,In_162);
nand U3526 (N_3526,In_2241,In_1275);
xnor U3527 (N_3527,In_1694,In_537);
and U3528 (N_3528,In_1897,In_2035);
and U3529 (N_3529,In_2052,In_1884);
nor U3530 (N_3530,In_1674,In_1302);
xnor U3531 (N_3531,In_2424,In_792);
and U3532 (N_3532,In_1383,In_414);
xnor U3533 (N_3533,In_2387,In_1366);
or U3534 (N_3534,In_1178,In_706);
xnor U3535 (N_3535,In_617,In_2294);
nand U3536 (N_3536,In_2033,In_2223);
xor U3537 (N_3537,In_1159,In_334);
nand U3538 (N_3538,In_804,In_1997);
nor U3539 (N_3539,In_1005,In_1100);
nor U3540 (N_3540,In_215,In_2286);
xnor U3541 (N_3541,In_151,In_2153);
and U3542 (N_3542,In_358,In_1566);
nand U3543 (N_3543,In_1076,In_1275);
and U3544 (N_3544,In_1974,In_1988);
xnor U3545 (N_3545,In_2401,In_589);
nor U3546 (N_3546,In_1771,In_1226);
nor U3547 (N_3547,In_2311,In_586);
or U3548 (N_3548,In_807,In_1339);
and U3549 (N_3549,In_1427,In_1120);
and U3550 (N_3550,In_782,In_991);
nand U3551 (N_3551,In_1076,In_1747);
or U3552 (N_3552,In_1488,In_2188);
and U3553 (N_3553,In_1788,In_1229);
or U3554 (N_3554,In_1302,In_2198);
nor U3555 (N_3555,In_2349,In_2347);
nand U3556 (N_3556,In_561,In_2316);
and U3557 (N_3557,In_1327,In_2308);
and U3558 (N_3558,In_772,In_1049);
xor U3559 (N_3559,In_6,In_1048);
xnor U3560 (N_3560,In_1617,In_2468);
nand U3561 (N_3561,In_403,In_2443);
xnor U3562 (N_3562,In_1039,In_2232);
nand U3563 (N_3563,In_2417,In_2385);
nor U3564 (N_3564,In_1612,In_1513);
nand U3565 (N_3565,In_1021,In_961);
xor U3566 (N_3566,In_1722,In_1719);
nand U3567 (N_3567,In_1578,In_2124);
nor U3568 (N_3568,In_1264,In_1220);
nor U3569 (N_3569,In_986,In_1244);
nor U3570 (N_3570,In_1316,In_1603);
or U3571 (N_3571,In_1392,In_1892);
nor U3572 (N_3572,In_1032,In_2042);
nor U3573 (N_3573,In_1885,In_2360);
or U3574 (N_3574,In_599,In_2134);
or U3575 (N_3575,In_1437,In_1514);
nand U3576 (N_3576,In_1566,In_1174);
or U3577 (N_3577,In_1380,In_1341);
and U3578 (N_3578,In_1083,In_560);
or U3579 (N_3579,In_502,In_1226);
nand U3580 (N_3580,In_431,In_1587);
and U3581 (N_3581,In_894,In_2019);
nor U3582 (N_3582,In_241,In_307);
nor U3583 (N_3583,In_569,In_1028);
or U3584 (N_3584,In_2289,In_494);
nand U3585 (N_3585,In_668,In_1505);
nand U3586 (N_3586,In_252,In_511);
and U3587 (N_3587,In_672,In_1946);
or U3588 (N_3588,In_2359,In_539);
xor U3589 (N_3589,In_1443,In_1024);
nor U3590 (N_3590,In_430,In_2203);
xnor U3591 (N_3591,In_2062,In_1168);
nor U3592 (N_3592,In_1308,In_1167);
or U3593 (N_3593,In_1860,In_657);
or U3594 (N_3594,In_382,In_1995);
nor U3595 (N_3595,In_2465,In_1778);
nor U3596 (N_3596,In_404,In_2490);
nand U3597 (N_3597,In_2108,In_1076);
and U3598 (N_3598,In_382,In_1928);
and U3599 (N_3599,In_939,In_1203);
and U3600 (N_3600,In_518,In_1461);
and U3601 (N_3601,In_2250,In_2101);
nor U3602 (N_3602,In_1995,In_249);
and U3603 (N_3603,In_347,In_290);
nand U3604 (N_3604,In_733,In_1651);
nor U3605 (N_3605,In_2278,In_473);
or U3606 (N_3606,In_1314,In_1140);
or U3607 (N_3607,In_1831,In_65);
xor U3608 (N_3608,In_843,In_2496);
and U3609 (N_3609,In_2257,In_1028);
xnor U3610 (N_3610,In_1282,In_2282);
xor U3611 (N_3611,In_2368,In_2447);
xnor U3612 (N_3612,In_1242,In_1227);
and U3613 (N_3613,In_669,In_448);
nand U3614 (N_3614,In_257,In_2466);
or U3615 (N_3615,In_2470,In_44);
nand U3616 (N_3616,In_448,In_821);
or U3617 (N_3617,In_2497,In_1824);
xor U3618 (N_3618,In_72,In_832);
xor U3619 (N_3619,In_231,In_1444);
xnor U3620 (N_3620,In_1084,In_1678);
and U3621 (N_3621,In_1849,In_27);
nand U3622 (N_3622,In_177,In_1991);
and U3623 (N_3623,In_50,In_2322);
or U3624 (N_3624,In_1796,In_1415);
and U3625 (N_3625,In_1936,In_385);
xnor U3626 (N_3626,In_226,In_2124);
or U3627 (N_3627,In_463,In_135);
xnor U3628 (N_3628,In_919,In_2210);
and U3629 (N_3629,In_1107,In_218);
xor U3630 (N_3630,In_1791,In_2111);
and U3631 (N_3631,In_1584,In_124);
or U3632 (N_3632,In_2249,In_416);
nor U3633 (N_3633,In_935,In_686);
xnor U3634 (N_3634,In_79,In_243);
or U3635 (N_3635,In_1456,In_1923);
and U3636 (N_3636,In_2346,In_1637);
nor U3637 (N_3637,In_1264,In_1875);
nand U3638 (N_3638,In_725,In_1868);
or U3639 (N_3639,In_1448,In_2146);
nor U3640 (N_3640,In_138,In_53);
and U3641 (N_3641,In_1254,In_331);
or U3642 (N_3642,In_81,In_2172);
xor U3643 (N_3643,In_733,In_930);
xnor U3644 (N_3644,In_1648,In_1790);
and U3645 (N_3645,In_1837,In_1427);
nand U3646 (N_3646,In_627,In_1177);
and U3647 (N_3647,In_478,In_1212);
xor U3648 (N_3648,In_1183,In_568);
and U3649 (N_3649,In_1563,In_1591);
xnor U3650 (N_3650,In_187,In_1324);
nand U3651 (N_3651,In_535,In_1320);
nand U3652 (N_3652,In_1113,In_2221);
xor U3653 (N_3653,In_1671,In_2126);
and U3654 (N_3654,In_2133,In_541);
nor U3655 (N_3655,In_784,In_2356);
nand U3656 (N_3656,In_1740,In_1376);
or U3657 (N_3657,In_1761,In_1795);
nand U3658 (N_3658,In_1042,In_1177);
and U3659 (N_3659,In_454,In_397);
nand U3660 (N_3660,In_1422,In_349);
nor U3661 (N_3661,In_1738,In_2239);
xor U3662 (N_3662,In_787,In_2338);
xnor U3663 (N_3663,In_1504,In_1697);
or U3664 (N_3664,In_2119,In_1965);
or U3665 (N_3665,In_2103,In_590);
and U3666 (N_3666,In_1225,In_1118);
and U3667 (N_3667,In_521,In_79);
or U3668 (N_3668,In_799,In_1876);
and U3669 (N_3669,In_257,In_1804);
or U3670 (N_3670,In_1053,In_1199);
or U3671 (N_3671,In_2348,In_2417);
nand U3672 (N_3672,In_650,In_1784);
and U3673 (N_3673,In_864,In_916);
or U3674 (N_3674,In_556,In_1446);
nand U3675 (N_3675,In_2121,In_199);
and U3676 (N_3676,In_275,In_98);
xnor U3677 (N_3677,In_1976,In_54);
or U3678 (N_3678,In_156,In_103);
and U3679 (N_3679,In_2137,In_741);
xor U3680 (N_3680,In_472,In_1372);
xor U3681 (N_3681,In_1527,In_555);
or U3682 (N_3682,In_1645,In_2456);
nor U3683 (N_3683,In_298,In_617);
or U3684 (N_3684,In_2310,In_341);
and U3685 (N_3685,In_1504,In_255);
nand U3686 (N_3686,In_550,In_1328);
xor U3687 (N_3687,In_1188,In_1675);
nor U3688 (N_3688,In_983,In_655);
and U3689 (N_3689,In_1906,In_342);
nor U3690 (N_3690,In_1009,In_1750);
and U3691 (N_3691,In_960,In_2390);
nor U3692 (N_3692,In_535,In_2477);
xor U3693 (N_3693,In_117,In_2127);
nand U3694 (N_3694,In_2371,In_1101);
nand U3695 (N_3695,In_1986,In_2048);
and U3696 (N_3696,In_1089,In_656);
nand U3697 (N_3697,In_32,In_550);
or U3698 (N_3698,In_32,In_956);
or U3699 (N_3699,In_360,In_1792);
xor U3700 (N_3700,In_1411,In_1883);
nand U3701 (N_3701,In_869,In_2118);
xnor U3702 (N_3702,In_930,In_889);
nand U3703 (N_3703,In_19,In_1808);
xor U3704 (N_3704,In_1834,In_2321);
or U3705 (N_3705,In_2050,In_1657);
and U3706 (N_3706,In_1641,In_843);
xor U3707 (N_3707,In_1950,In_1457);
and U3708 (N_3708,In_118,In_760);
nand U3709 (N_3709,In_28,In_2158);
nand U3710 (N_3710,In_1099,In_1538);
or U3711 (N_3711,In_1989,In_2455);
and U3712 (N_3712,In_1175,In_1312);
and U3713 (N_3713,In_126,In_1208);
and U3714 (N_3714,In_1341,In_1176);
and U3715 (N_3715,In_2491,In_1347);
xor U3716 (N_3716,In_1463,In_2083);
and U3717 (N_3717,In_578,In_2289);
nor U3718 (N_3718,In_723,In_1872);
or U3719 (N_3719,In_925,In_690);
nor U3720 (N_3720,In_2078,In_430);
nor U3721 (N_3721,In_686,In_2291);
and U3722 (N_3722,In_1470,In_1449);
nor U3723 (N_3723,In_1110,In_1425);
and U3724 (N_3724,In_1533,In_254);
or U3725 (N_3725,In_2481,In_2358);
and U3726 (N_3726,In_632,In_68);
nand U3727 (N_3727,In_1072,In_438);
nor U3728 (N_3728,In_192,In_155);
nand U3729 (N_3729,In_66,In_837);
nor U3730 (N_3730,In_449,In_368);
nand U3731 (N_3731,In_2147,In_2327);
and U3732 (N_3732,In_1052,In_2084);
xnor U3733 (N_3733,In_933,In_404);
and U3734 (N_3734,In_1831,In_1361);
xnor U3735 (N_3735,In_2307,In_170);
and U3736 (N_3736,In_1235,In_2069);
xnor U3737 (N_3737,In_1018,In_1361);
and U3738 (N_3738,In_1838,In_1198);
xor U3739 (N_3739,In_2435,In_208);
xor U3740 (N_3740,In_1466,In_398);
or U3741 (N_3741,In_439,In_1877);
or U3742 (N_3742,In_394,In_860);
xor U3743 (N_3743,In_1484,In_2147);
nand U3744 (N_3744,In_484,In_525);
and U3745 (N_3745,In_1566,In_946);
nor U3746 (N_3746,In_94,In_1059);
and U3747 (N_3747,In_1955,In_934);
nor U3748 (N_3748,In_1655,In_1446);
and U3749 (N_3749,In_1131,In_178);
or U3750 (N_3750,In_621,In_1844);
nor U3751 (N_3751,In_596,In_2481);
or U3752 (N_3752,In_1406,In_1652);
or U3753 (N_3753,In_1946,In_884);
nand U3754 (N_3754,In_229,In_280);
or U3755 (N_3755,In_512,In_1232);
nand U3756 (N_3756,In_1877,In_875);
and U3757 (N_3757,In_2193,In_1263);
and U3758 (N_3758,In_2201,In_758);
or U3759 (N_3759,In_2323,In_2247);
xor U3760 (N_3760,In_772,In_1279);
nand U3761 (N_3761,In_2018,In_511);
or U3762 (N_3762,In_1176,In_1161);
and U3763 (N_3763,In_1648,In_71);
and U3764 (N_3764,In_1513,In_1962);
nor U3765 (N_3765,In_2285,In_31);
xnor U3766 (N_3766,In_129,In_277);
or U3767 (N_3767,In_428,In_102);
nand U3768 (N_3768,In_903,In_949);
and U3769 (N_3769,In_1584,In_1714);
or U3770 (N_3770,In_781,In_1556);
and U3771 (N_3771,In_1876,In_1448);
xor U3772 (N_3772,In_279,In_1465);
xor U3773 (N_3773,In_886,In_2092);
nor U3774 (N_3774,In_1007,In_1164);
xor U3775 (N_3775,In_1564,In_1773);
nor U3776 (N_3776,In_1376,In_1605);
or U3777 (N_3777,In_1443,In_1565);
or U3778 (N_3778,In_1689,In_2047);
and U3779 (N_3779,In_1072,In_2482);
xnor U3780 (N_3780,In_1331,In_441);
or U3781 (N_3781,In_935,In_1036);
or U3782 (N_3782,In_133,In_1280);
or U3783 (N_3783,In_2425,In_1942);
xnor U3784 (N_3784,In_1090,In_2217);
nand U3785 (N_3785,In_2461,In_2137);
or U3786 (N_3786,In_1064,In_668);
or U3787 (N_3787,In_1687,In_270);
and U3788 (N_3788,In_106,In_1227);
nor U3789 (N_3789,In_223,In_2437);
nand U3790 (N_3790,In_2449,In_2427);
or U3791 (N_3791,In_1254,In_1751);
nand U3792 (N_3792,In_1714,In_1164);
xnor U3793 (N_3793,In_782,In_566);
or U3794 (N_3794,In_1146,In_1800);
nand U3795 (N_3795,In_1192,In_1719);
nor U3796 (N_3796,In_1485,In_1493);
nand U3797 (N_3797,In_1474,In_910);
xnor U3798 (N_3798,In_627,In_1496);
nor U3799 (N_3799,In_1713,In_2411);
nor U3800 (N_3800,In_2006,In_2336);
and U3801 (N_3801,In_887,In_1292);
or U3802 (N_3802,In_674,In_407);
and U3803 (N_3803,In_646,In_1579);
xor U3804 (N_3804,In_727,In_1327);
nor U3805 (N_3805,In_2418,In_1477);
nor U3806 (N_3806,In_1860,In_688);
or U3807 (N_3807,In_2405,In_1549);
nor U3808 (N_3808,In_2139,In_650);
nor U3809 (N_3809,In_2163,In_586);
xnor U3810 (N_3810,In_1875,In_2326);
nor U3811 (N_3811,In_1440,In_589);
or U3812 (N_3812,In_413,In_1002);
xnor U3813 (N_3813,In_2021,In_1754);
and U3814 (N_3814,In_1655,In_26);
xnor U3815 (N_3815,In_533,In_424);
nor U3816 (N_3816,In_492,In_2469);
xnor U3817 (N_3817,In_337,In_1792);
xor U3818 (N_3818,In_611,In_1022);
nor U3819 (N_3819,In_2240,In_1735);
nand U3820 (N_3820,In_1905,In_1398);
and U3821 (N_3821,In_2184,In_596);
and U3822 (N_3822,In_78,In_364);
and U3823 (N_3823,In_2453,In_2182);
nor U3824 (N_3824,In_50,In_252);
nand U3825 (N_3825,In_1014,In_688);
xor U3826 (N_3826,In_2447,In_462);
and U3827 (N_3827,In_1440,In_1378);
xor U3828 (N_3828,In_879,In_1149);
nor U3829 (N_3829,In_152,In_1982);
nand U3830 (N_3830,In_1736,In_2325);
xor U3831 (N_3831,In_1780,In_2495);
nor U3832 (N_3832,In_2131,In_1006);
nor U3833 (N_3833,In_186,In_756);
or U3834 (N_3834,In_798,In_1842);
nand U3835 (N_3835,In_1913,In_2230);
nand U3836 (N_3836,In_518,In_579);
xor U3837 (N_3837,In_2036,In_1523);
xor U3838 (N_3838,In_2436,In_1625);
nor U3839 (N_3839,In_721,In_600);
nand U3840 (N_3840,In_335,In_624);
xnor U3841 (N_3841,In_65,In_172);
xor U3842 (N_3842,In_836,In_1225);
or U3843 (N_3843,In_1522,In_1855);
or U3844 (N_3844,In_1584,In_1683);
nor U3845 (N_3845,In_670,In_1509);
xnor U3846 (N_3846,In_117,In_1396);
xnor U3847 (N_3847,In_1219,In_1032);
and U3848 (N_3848,In_1831,In_1697);
and U3849 (N_3849,In_318,In_98);
nor U3850 (N_3850,In_1587,In_1542);
and U3851 (N_3851,In_916,In_1477);
nand U3852 (N_3852,In_118,In_309);
nand U3853 (N_3853,In_2354,In_1948);
and U3854 (N_3854,In_1386,In_1608);
nor U3855 (N_3855,In_1784,In_1767);
or U3856 (N_3856,In_2026,In_198);
xnor U3857 (N_3857,In_2174,In_0);
or U3858 (N_3858,In_2166,In_167);
and U3859 (N_3859,In_2306,In_2475);
nor U3860 (N_3860,In_2114,In_1836);
nor U3861 (N_3861,In_1654,In_1354);
xor U3862 (N_3862,In_1507,In_1479);
or U3863 (N_3863,In_2364,In_2144);
xor U3864 (N_3864,In_1842,In_2355);
nand U3865 (N_3865,In_1184,In_876);
and U3866 (N_3866,In_626,In_342);
or U3867 (N_3867,In_245,In_37);
xor U3868 (N_3868,In_726,In_1219);
and U3869 (N_3869,In_2043,In_2150);
or U3870 (N_3870,In_2071,In_2228);
nor U3871 (N_3871,In_75,In_2122);
or U3872 (N_3872,In_1317,In_74);
nand U3873 (N_3873,In_2330,In_755);
and U3874 (N_3874,In_2375,In_1506);
and U3875 (N_3875,In_35,In_950);
xor U3876 (N_3876,In_1533,In_712);
or U3877 (N_3877,In_2268,In_281);
nand U3878 (N_3878,In_1427,In_676);
xnor U3879 (N_3879,In_2231,In_1323);
nand U3880 (N_3880,In_2284,In_482);
and U3881 (N_3881,In_393,In_244);
and U3882 (N_3882,In_1261,In_237);
or U3883 (N_3883,In_2195,In_589);
nor U3884 (N_3884,In_2430,In_312);
or U3885 (N_3885,In_979,In_1670);
nand U3886 (N_3886,In_339,In_1556);
xor U3887 (N_3887,In_2250,In_74);
nor U3888 (N_3888,In_2358,In_2082);
and U3889 (N_3889,In_1590,In_83);
xnor U3890 (N_3890,In_1508,In_1635);
and U3891 (N_3891,In_1577,In_576);
nor U3892 (N_3892,In_1880,In_1704);
nand U3893 (N_3893,In_1249,In_2133);
nand U3894 (N_3894,In_1288,In_1645);
nand U3895 (N_3895,In_659,In_77);
and U3896 (N_3896,In_993,In_2184);
xor U3897 (N_3897,In_819,In_944);
xor U3898 (N_3898,In_438,In_1512);
xnor U3899 (N_3899,In_1699,In_2320);
and U3900 (N_3900,In_1502,In_1743);
nand U3901 (N_3901,In_526,In_964);
nand U3902 (N_3902,In_866,In_2396);
nor U3903 (N_3903,In_2372,In_559);
xor U3904 (N_3904,In_449,In_851);
nand U3905 (N_3905,In_1861,In_1084);
nor U3906 (N_3906,In_409,In_1342);
nor U3907 (N_3907,In_2401,In_446);
xor U3908 (N_3908,In_343,In_607);
and U3909 (N_3909,In_1389,In_725);
nor U3910 (N_3910,In_453,In_1680);
nand U3911 (N_3911,In_991,In_1159);
nor U3912 (N_3912,In_1084,In_2076);
and U3913 (N_3913,In_1539,In_432);
nor U3914 (N_3914,In_2158,In_1605);
xor U3915 (N_3915,In_503,In_500);
nor U3916 (N_3916,In_720,In_869);
nor U3917 (N_3917,In_1301,In_1932);
xnor U3918 (N_3918,In_1911,In_2474);
nand U3919 (N_3919,In_571,In_2398);
nand U3920 (N_3920,In_100,In_1020);
and U3921 (N_3921,In_762,In_1734);
and U3922 (N_3922,In_715,In_1244);
nand U3923 (N_3923,In_2066,In_1488);
nor U3924 (N_3924,In_1147,In_1986);
and U3925 (N_3925,In_1887,In_1064);
and U3926 (N_3926,In_1837,In_542);
nor U3927 (N_3927,In_1882,In_1841);
xnor U3928 (N_3928,In_853,In_2016);
and U3929 (N_3929,In_1751,In_1946);
or U3930 (N_3930,In_837,In_2276);
nand U3931 (N_3931,In_965,In_1540);
nand U3932 (N_3932,In_413,In_422);
and U3933 (N_3933,In_2032,In_782);
xor U3934 (N_3934,In_1862,In_510);
nor U3935 (N_3935,In_1165,In_250);
nand U3936 (N_3936,In_2240,In_43);
nand U3937 (N_3937,In_1501,In_2209);
or U3938 (N_3938,In_1566,In_0);
nand U3939 (N_3939,In_1762,In_1931);
nand U3940 (N_3940,In_1413,In_779);
nand U3941 (N_3941,In_2245,In_942);
and U3942 (N_3942,In_1468,In_901);
nand U3943 (N_3943,In_2195,In_683);
xor U3944 (N_3944,In_516,In_1407);
and U3945 (N_3945,In_109,In_1550);
or U3946 (N_3946,In_1944,In_854);
and U3947 (N_3947,In_1257,In_424);
and U3948 (N_3948,In_2019,In_1315);
nor U3949 (N_3949,In_984,In_1176);
and U3950 (N_3950,In_938,In_108);
nor U3951 (N_3951,In_752,In_169);
or U3952 (N_3952,In_1462,In_755);
and U3953 (N_3953,In_2343,In_12);
or U3954 (N_3954,In_1465,In_1396);
and U3955 (N_3955,In_1368,In_664);
xor U3956 (N_3956,In_1457,In_892);
nand U3957 (N_3957,In_1854,In_2260);
xnor U3958 (N_3958,In_1323,In_1517);
nor U3959 (N_3959,In_1936,In_1374);
nand U3960 (N_3960,In_1090,In_1566);
xor U3961 (N_3961,In_1002,In_253);
xnor U3962 (N_3962,In_2327,In_268);
nand U3963 (N_3963,In_1950,In_1113);
nor U3964 (N_3964,In_502,In_93);
nor U3965 (N_3965,In_2308,In_2);
xnor U3966 (N_3966,In_486,In_444);
nand U3967 (N_3967,In_712,In_1733);
xnor U3968 (N_3968,In_176,In_425);
nand U3969 (N_3969,In_2113,In_1078);
nor U3970 (N_3970,In_434,In_521);
nand U3971 (N_3971,In_614,In_369);
and U3972 (N_3972,In_685,In_2190);
nor U3973 (N_3973,In_738,In_743);
nand U3974 (N_3974,In_605,In_846);
and U3975 (N_3975,In_394,In_4);
or U3976 (N_3976,In_140,In_101);
nor U3977 (N_3977,In_476,In_622);
nor U3978 (N_3978,In_2068,In_1074);
and U3979 (N_3979,In_1013,In_387);
xnor U3980 (N_3980,In_885,In_2412);
nand U3981 (N_3981,In_314,In_820);
xnor U3982 (N_3982,In_2065,In_1565);
nand U3983 (N_3983,In_1746,In_770);
xnor U3984 (N_3984,In_2052,In_158);
nand U3985 (N_3985,In_741,In_244);
nand U3986 (N_3986,In_1834,In_875);
and U3987 (N_3987,In_1953,In_1623);
nand U3988 (N_3988,In_36,In_1676);
and U3989 (N_3989,In_1862,In_1460);
or U3990 (N_3990,In_2441,In_12);
and U3991 (N_3991,In_82,In_643);
nor U3992 (N_3992,In_1579,In_1530);
or U3993 (N_3993,In_762,In_1398);
or U3994 (N_3994,In_1997,In_1424);
nand U3995 (N_3995,In_1551,In_790);
and U3996 (N_3996,In_1859,In_2248);
or U3997 (N_3997,In_1440,In_1591);
xor U3998 (N_3998,In_85,In_1681);
or U3999 (N_3999,In_600,In_785);
and U4000 (N_4000,In_1817,In_848);
nor U4001 (N_4001,In_1296,In_769);
nor U4002 (N_4002,In_1776,In_2473);
nor U4003 (N_4003,In_547,In_1982);
nand U4004 (N_4004,In_112,In_2121);
nor U4005 (N_4005,In_2111,In_248);
and U4006 (N_4006,In_618,In_2420);
and U4007 (N_4007,In_396,In_2108);
xnor U4008 (N_4008,In_224,In_487);
xnor U4009 (N_4009,In_678,In_2075);
nor U4010 (N_4010,In_133,In_2153);
and U4011 (N_4011,In_1925,In_2047);
or U4012 (N_4012,In_2463,In_921);
nor U4013 (N_4013,In_407,In_2278);
nor U4014 (N_4014,In_2141,In_2304);
nor U4015 (N_4015,In_1164,In_991);
nor U4016 (N_4016,In_193,In_2184);
and U4017 (N_4017,In_2301,In_2264);
or U4018 (N_4018,In_867,In_1953);
nand U4019 (N_4019,In_628,In_66);
and U4020 (N_4020,In_2084,In_661);
nor U4021 (N_4021,In_2021,In_2300);
and U4022 (N_4022,In_2155,In_1359);
xor U4023 (N_4023,In_863,In_1943);
xor U4024 (N_4024,In_731,In_898);
xnor U4025 (N_4025,In_2139,In_2332);
xnor U4026 (N_4026,In_2372,In_737);
nand U4027 (N_4027,In_2184,In_2044);
nor U4028 (N_4028,In_2360,In_1898);
nor U4029 (N_4029,In_1395,In_215);
nor U4030 (N_4030,In_1695,In_2465);
xor U4031 (N_4031,In_331,In_49);
nand U4032 (N_4032,In_1453,In_706);
or U4033 (N_4033,In_1571,In_1849);
and U4034 (N_4034,In_1747,In_2443);
xnor U4035 (N_4035,In_186,In_1205);
xor U4036 (N_4036,In_2464,In_295);
and U4037 (N_4037,In_1914,In_346);
xor U4038 (N_4038,In_1563,In_677);
nor U4039 (N_4039,In_2,In_963);
nand U4040 (N_4040,In_1762,In_1151);
or U4041 (N_4041,In_588,In_2314);
or U4042 (N_4042,In_1506,In_556);
nand U4043 (N_4043,In_427,In_157);
xnor U4044 (N_4044,In_1590,In_2077);
and U4045 (N_4045,In_70,In_2022);
xnor U4046 (N_4046,In_725,In_1607);
or U4047 (N_4047,In_2326,In_2084);
xnor U4048 (N_4048,In_13,In_2488);
xnor U4049 (N_4049,In_1924,In_1411);
or U4050 (N_4050,In_571,In_217);
or U4051 (N_4051,In_678,In_1484);
nand U4052 (N_4052,In_1517,In_721);
nand U4053 (N_4053,In_1349,In_28);
nor U4054 (N_4054,In_1762,In_783);
or U4055 (N_4055,In_2212,In_238);
nand U4056 (N_4056,In_113,In_2299);
nor U4057 (N_4057,In_1309,In_1074);
nor U4058 (N_4058,In_2326,In_2394);
xnor U4059 (N_4059,In_1402,In_1269);
nor U4060 (N_4060,In_2331,In_1444);
nand U4061 (N_4061,In_2467,In_2497);
nor U4062 (N_4062,In_717,In_2346);
nor U4063 (N_4063,In_1546,In_189);
nor U4064 (N_4064,In_212,In_1289);
xnor U4065 (N_4065,In_1522,In_1728);
xor U4066 (N_4066,In_640,In_2133);
xnor U4067 (N_4067,In_237,In_804);
or U4068 (N_4068,In_607,In_888);
or U4069 (N_4069,In_196,In_1835);
and U4070 (N_4070,In_1821,In_453);
xor U4071 (N_4071,In_421,In_2225);
nand U4072 (N_4072,In_2321,In_805);
xor U4073 (N_4073,In_1754,In_1826);
xor U4074 (N_4074,In_1391,In_482);
or U4075 (N_4075,In_460,In_231);
nand U4076 (N_4076,In_1473,In_1074);
xnor U4077 (N_4077,In_1918,In_812);
nand U4078 (N_4078,In_37,In_1718);
nand U4079 (N_4079,In_40,In_1897);
nand U4080 (N_4080,In_154,In_946);
nor U4081 (N_4081,In_2420,In_1224);
or U4082 (N_4082,In_2154,In_387);
xnor U4083 (N_4083,In_1028,In_1617);
nand U4084 (N_4084,In_1597,In_1213);
or U4085 (N_4085,In_777,In_1281);
xnor U4086 (N_4086,In_621,In_172);
and U4087 (N_4087,In_712,In_1398);
nand U4088 (N_4088,In_1480,In_1625);
nand U4089 (N_4089,In_1413,In_418);
xor U4090 (N_4090,In_1248,In_1906);
and U4091 (N_4091,In_1373,In_488);
nand U4092 (N_4092,In_1156,In_303);
xor U4093 (N_4093,In_2005,In_2403);
nor U4094 (N_4094,In_1085,In_1794);
or U4095 (N_4095,In_47,In_216);
nor U4096 (N_4096,In_954,In_1343);
and U4097 (N_4097,In_100,In_893);
nor U4098 (N_4098,In_1277,In_1290);
or U4099 (N_4099,In_2473,In_194);
and U4100 (N_4100,In_817,In_53);
and U4101 (N_4101,In_2212,In_1827);
or U4102 (N_4102,In_428,In_419);
or U4103 (N_4103,In_300,In_577);
and U4104 (N_4104,In_2216,In_214);
xnor U4105 (N_4105,In_556,In_612);
nor U4106 (N_4106,In_1080,In_2265);
and U4107 (N_4107,In_528,In_2040);
nand U4108 (N_4108,In_926,In_2234);
or U4109 (N_4109,In_2355,In_733);
and U4110 (N_4110,In_245,In_2399);
or U4111 (N_4111,In_1265,In_954);
or U4112 (N_4112,In_45,In_2269);
or U4113 (N_4113,In_1999,In_772);
nand U4114 (N_4114,In_1896,In_755);
and U4115 (N_4115,In_2113,In_1822);
nand U4116 (N_4116,In_2075,In_531);
or U4117 (N_4117,In_2167,In_760);
or U4118 (N_4118,In_2033,In_1051);
or U4119 (N_4119,In_251,In_699);
or U4120 (N_4120,In_1080,In_1525);
and U4121 (N_4121,In_2443,In_848);
xnor U4122 (N_4122,In_106,In_462);
and U4123 (N_4123,In_2161,In_1870);
xnor U4124 (N_4124,In_392,In_1606);
and U4125 (N_4125,In_1159,In_148);
and U4126 (N_4126,In_2247,In_2063);
nand U4127 (N_4127,In_1741,In_576);
nand U4128 (N_4128,In_1716,In_1088);
nand U4129 (N_4129,In_529,In_2187);
nor U4130 (N_4130,In_2451,In_1822);
nand U4131 (N_4131,In_1338,In_166);
nor U4132 (N_4132,In_217,In_331);
xor U4133 (N_4133,In_1809,In_1620);
nand U4134 (N_4134,In_1921,In_1251);
nand U4135 (N_4135,In_1257,In_121);
and U4136 (N_4136,In_667,In_2382);
nor U4137 (N_4137,In_1337,In_886);
and U4138 (N_4138,In_1613,In_1293);
nand U4139 (N_4139,In_1306,In_113);
and U4140 (N_4140,In_1552,In_1881);
and U4141 (N_4141,In_2319,In_1434);
nor U4142 (N_4142,In_216,In_1290);
and U4143 (N_4143,In_1710,In_1942);
or U4144 (N_4144,In_1491,In_2169);
xnor U4145 (N_4145,In_595,In_1392);
and U4146 (N_4146,In_1424,In_1127);
or U4147 (N_4147,In_1863,In_1465);
or U4148 (N_4148,In_1337,In_662);
nand U4149 (N_4149,In_406,In_2287);
and U4150 (N_4150,In_973,In_482);
and U4151 (N_4151,In_676,In_1886);
or U4152 (N_4152,In_1799,In_1890);
or U4153 (N_4153,In_755,In_871);
nor U4154 (N_4154,In_239,In_2223);
nor U4155 (N_4155,In_1962,In_2234);
and U4156 (N_4156,In_1115,In_774);
xor U4157 (N_4157,In_591,In_290);
xnor U4158 (N_4158,In_1765,In_424);
and U4159 (N_4159,In_2351,In_2412);
and U4160 (N_4160,In_619,In_231);
or U4161 (N_4161,In_337,In_1912);
nor U4162 (N_4162,In_57,In_1715);
nand U4163 (N_4163,In_560,In_47);
and U4164 (N_4164,In_167,In_2192);
xor U4165 (N_4165,In_1848,In_120);
and U4166 (N_4166,In_541,In_1026);
or U4167 (N_4167,In_2358,In_541);
nor U4168 (N_4168,In_56,In_1373);
and U4169 (N_4169,In_659,In_1483);
or U4170 (N_4170,In_237,In_977);
xor U4171 (N_4171,In_125,In_1096);
and U4172 (N_4172,In_184,In_1078);
xnor U4173 (N_4173,In_2169,In_2406);
and U4174 (N_4174,In_907,In_1673);
nand U4175 (N_4175,In_959,In_2287);
nand U4176 (N_4176,In_926,In_345);
xor U4177 (N_4177,In_454,In_2123);
xnor U4178 (N_4178,In_1874,In_2176);
and U4179 (N_4179,In_1753,In_2223);
nor U4180 (N_4180,In_1234,In_263);
nand U4181 (N_4181,In_2488,In_2188);
and U4182 (N_4182,In_1922,In_146);
nand U4183 (N_4183,In_1379,In_1628);
nand U4184 (N_4184,In_2278,In_2101);
nor U4185 (N_4185,In_169,In_297);
xnor U4186 (N_4186,In_1268,In_997);
nand U4187 (N_4187,In_2300,In_1244);
xnor U4188 (N_4188,In_50,In_2140);
nand U4189 (N_4189,In_1995,In_2312);
or U4190 (N_4190,In_432,In_1572);
xor U4191 (N_4191,In_1345,In_874);
and U4192 (N_4192,In_1712,In_2239);
and U4193 (N_4193,In_2048,In_1510);
nand U4194 (N_4194,In_564,In_1955);
nand U4195 (N_4195,In_276,In_66);
nor U4196 (N_4196,In_2384,In_405);
xnor U4197 (N_4197,In_2212,In_343);
nor U4198 (N_4198,In_1735,In_479);
xor U4199 (N_4199,In_2352,In_243);
nor U4200 (N_4200,In_1654,In_263);
nor U4201 (N_4201,In_2005,In_1104);
nand U4202 (N_4202,In_1538,In_1747);
xor U4203 (N_4203,In_2317,In_886);
nor U4204 (N_4204,In_1857,In_1792);
and U4205 (N_4205,In_2257,In_2278);
and U4206 (N_4206,In_951,In_1710);
nand U4207 (N_4207,In_2110,In_993);
nand U4208 (N_4208,In_2363,In_1790);
or U4209 (N_4209,In_1415,In_2006);
and U4210 (N_4210,In_271,In_1274);
or U4211 (N_4211,In_1055,In_2125);
and U4212 (N_4212,In_210,In_2498);
and U4213 (N_4213,In_1194,In_1568);
and U4214 (N_4214,In_447,In_1697);
xnor U4215 (N_4215,In_2422,In_1188);
nand U4216 (N_4216,In_2470,In_1994);
nand U4217 (N_4217,In_759,In_1641);
nand U4218 (N_4218,In_2459,In_1697);
xor U4219 (N_4219,In_1648,In_2049);
xor U4220 (N_4220,In_2168,In_134);
xor U4221 (N_4221,In_897,In_163);
nand U4222 (N_4222,In_173,In_1163);
or U4223 (N_4223,In_1914,In_262);
and U4224 (N_4224,In_220,In_233);
nand U4225 (N_4225,In_184,In_1574);
nand U4226 (N_4226,In_1884,In_2279);
xor U4227 (N_4227,In_913,In_2316);
and U4228 (N_4228,In_391,In_1545);
or U4229 (N_4229,In_1067,In_337);
nand U4230 (N_4230,In_2474,In_1920);
or U4231 (N_4231,In_758,In_1063);
or U4232 (N_4232,In_2173,In_1982);
and U4233 (N_4233,In_594,In_221);
nand U4234 (N_4234,In_1420,In_1470);
xor U4235 (N_4235,In_1119,In_2292);
nand U4236 (N_4236,In_534,In_861);
or U4237 (N_4237,In_1544,In_899);
xor U4238 (N_4238,In_2128,In_330);
and U4239 (N_4239,In_475,In_1337);
and U4240 (N_4240,In_995,In_699);
nor U4241 (N_4241,In_1452,In_1109);
or U4242 (N_4242,In_721,In_1463);
nand U4243 (N_4243,In_1846,In_1590);
or U4244 (N_4244,In_917,In_2066);
or U4245 (N_4245,In_2208,In_1440);
xnor U4246 (N_4246,In_1525,In_1025);
nand U4247 (N_4247,In_1995,In_192);
and U4248 (N_4248,In_2474,In_452);
xnor U4249 (N_4249,In_2159,In_1849);
or U4250 (N_4250,In_1441,In_1727);
nor U4251 (N_4251,In_1513,In_2033);
nor U4252 (N_4252,In_538,In_1417);
nor U4253 (N_4253,In_1388,In_789);
and U4254 (N_4254,In_316,In_1840);
or U4255 (N_4255,In_2403,In_968);
and U4256 (N_4256,In_654,In_1149);
and U4257 (N_4257,In_1273,In_1280);
xnor U4258 (N_4258,In_711,In_1300);
xor U4259 (N_4259,In_2198,In_1129);
nand U4260 (N_4260,In_2127,In_68);
xnor U4261 (N_4261,In_90,In_2298);
nor U4262 (N_4262,In_849,In_2046);
and U4263 (N_4263,In_2474,In_623);
nand U4264 (N_4264,In_813,In_597);
nand U4265 (N_4265,In_1068,In_2396);
xnor U4266 (N_4266,In_1042,In_11);
and U4267 (N_4267,In_746,In_2385);
and U4268 (N_4268,In_2336,In_2009);
and U4269 (N_4269,In_1468,In_2039);
nor U4270 (N_4270,In_2182,In_12);
xnor U4271 (N_4271,In_347,In_2472);
xnor U4272 (N_4272,In_2184,In_344);
nor U4273 (N_4273,In_2480,In_2303);
xor U4274 (N_4274,In_313,In_1939);
and U4275 (N_4275,In_2145,In_1661);
nand U4276 (N_4276,In_596,In_232);
or U4277 (N_4277,In_690,In_428);
nor U4278 (N_4278,In_2063,In_37);
and U4279 (N_4279,In_2023,In_684);
xor U4280 (N_4280,In_2128,In_1750);
xnor U4281 (N_4281,In_1728,In_602);
xor U4282 (N_4282,In_1790,In_399);
nor U4283 (N_4283,In_415,In_1159);
nor U4284 (N_4284,In_1786,In_1699);
or U4285 (N_4285,In_1294,In_2288);
and U4286 (N_4286,In_1093,In_116);
nand U4287 (N_4287,In_263,In_1317);
nor U4288 (N_4288,In_850,In_2069);
xor U4289 (N_4289,In_1952,In_891);
nand U4290 (N_4290,In_1315,In_2190);
or U4291 (N_4291,In_1606,In_1004);
nand U4292 (N_4292,In_2288,In_255);
or U4293 (N_4293,In_195,In_764);
or U4294 (N_4294,In_2371,In_573);
nand U4295 (N_4295,In_423,In_1646);
nor U4296 (N_4296,In_1250,In_683);
and U4297 (N_4297,In_429,In_1101);
or U4298 (N_4298,In_176,In_0);
and U4299 (N_4299,In_798,In_1184);
or U4300 (N_4300,In_759,In_940);
or U4301 (N_4301,In_172,In_376);
and U4302 (N_4302,In_833,In_2182);
or U4303 (N_4303,In_2386,In_1374);
nand U4304 (N_4304,In_999,In_32);
nor U4305 (N_4305,In_1578,In_1125);
nand U4306 (N_4306,In_2438,In_538);
and U4307 (N_4307,In_535,In_1660);
nor U4308 (N_4308,In_2082,In_680);
nand U4309 (N_4309,In_875,In_2264);
nand U4310 (N_4310,In_1543,In_479);
xor U4311 (N_4311,In_2322,In_645);
xnor U4312 (N_4312,In_2070,In_40);
and U4313 (N_4313,In_1267,In_2192);
xor U4314 (N_4314,In_656,In_171);
xor U4315 (N_4315,In_1982,In_909);
or U4316 (N_4316,In_620,In_1467);
nand U4317 (N_4317,In_2431,In_2055);
nor U4318 (N_4318,In_1166,In_2490);
or U4319 (N_4319,In_2061,In_2024);
xor U4320 (N_4320,In_1453,In_1130);
or U4321 (N_4321,In_1416,In_11);
nor U4322 (N_4322,In_2203,In_2143);
or U4323 (N_4323,In_305,In_408);
xnor U4324 (N_4324,In_1872,In_989);
nor U4325 (N_4325,In_1397,In_1048);
or U4326 (N_4326,In_24,In_989);
and U4327 (N_4327,In_2423,In_2118);
nor U4328 (N_4328,In_999,In_1778);
or U4329 (N_4329,In_122,In_2300);
xor U4330 (N_4330,In_1260,In_401);
nand U4331 (N_4331,In_1281,In_1424);
xnor U4332 (N_4332,In_2312,In_1291);
nand U4333 (N_4333,In_600,In_1153);
xor U4334 (N_4334,In_325,In_781);
nand U4335 (N_4335,In_891,In_265);
xor U4336 (N_4336,In_276,In_1284);
nor U4337 (N_4337,In_1535,In_1063);
nand U4338 (N_4338,In_1718,In_491);
and U4339 (N_4339,In_2429,In_1496);
nor U4340 (N_4340,In_1113,In_2068);
or U4341 (N_4341,In_209,In_798);
xnor U4342 (N_4342,In_1249,In_710);
nor U4343 (N_4343,In_182,In_1038);
and U4344 (N_4344,In_822,In_671);
and U4345 (N_4345,In_1231,In_1882);
nand U4346 (N_4346,In_2160,In_1234);
and U4347 (N_4347,In_1755,In_1842);
nor U4348 (N_4348,In_1749,In_2221);
and U4349 (N_4349,In_2466,In_2207);
nand U4350 (N_4350,In_1901,In_298);
nor U4351 (N_4351,In_889,In_1881);
and U4352 (N_4352,In_138,In_2371);
or U4353 (N_4353,In_1328,In_1317);
and U4354 (N_4354,In_1584,In_568);
xor U4355 (N_4355,In_1556,In_1101);
and U4356 (N_4356,In_724,In_2087);
xnor U4357 (N_4357,In_1807,In_1140);
xor U4358 (N_4358,In_2134,In_111);
xnor U4359 (N_4359,In_1281,In_156);
or U4360 (N_4360,In_811,In_779);
nand U4361 (N_4361,In_1445,In_1884);
or U4362 (N_4362,In_2315,In_2258);
or U4363 (N_4363,In_2150,In_1444);
or U4364 (N_4364,In_1075,In_1700);
or U4365 (N_4365,In_2115,In_2234);
nand U4366 (N_4366,In_543,In_71);
and U4367 (N_4367,In_777,In_218);
nor U4368 (N_4368,In_1129,In_1032);
and U4369 (N_4369,In_2251,In_198);
and U4370 (N_4370,In_691,In_1095);
xnor U4371 (N_4371,In_217,In_2425);
or U4372 (N_4372,In_2378,In_1001);
and U4373 (N_4373,In_592,In_1722);
and U4374 (N_4374,In_1251,In_674);
or U4375 (N_4375,In_522,In_1805);
or U4376 (N_4376,In_1347,In_2052);
nand U4377 (N_4377,In_410,In_44);
nand U4378 (N_4378,In_2281,In_1945);
xnor U4379 (N_4379,In_1220,In_1350);
nand U4380 (N_4380,In_765,In_1646);
xor U4381 (N_4381,In_98,In_1818);
nor U4382 (N_4382,In_2260,In_751);
nand U4383 (N_4383,In_1228,In_440);
or U4384 (N_4384,In_584,In_1546);
or U4385 (N_4385,In_2107,In_1206);
and U4386 (N_4386,In_2399,In_593);
nand U4387 (N_4387,In_1912,In_2086);
or U4388 (N_4388,In_604,In_302);
nor U4389 (N_4389,In_830,In_2229);
and U4390 (N_4390,In_1825,In_2298);
nor U4391 (N_4391,In_431,In_2025);
nand U4392 (N_4392,In_1861,In_128);
nand U4393 (N_4393,In_2077,In_98);
xnor U4394 (N_4394,In_2082,In_1642);
nand U4395 (N_4395,In_1769,In_814);
nor U4396 (N_4396,In_897,In_1277);
xnor U4397 (N_4397,In_516,In_146);
and U4398 (N_4398,In_613,In_2234);
nor U4399 (N_4399,In_619,In_1229);
nor U4400 (N_4400,In_1942,In_1332);
or U4401 (N_4401,In_1896,In_1374);
xor U4402 (N_4402,In_447,In_908);
xor U4403 (N_4403,In_193,In_871);
xor U4404 (N_4404,In_1888,In_323);
nor U4405 (N_4405,In_990,In_1505);
xnor U4406 (N_4406,In_2427,In_573);
xor U4407 (N_4407,In_899,In_258);
or U4408 (N_4408,In_1561,In_1246);
nand U4409 (N_4409,In_1581,In_52);
or U4410 (N_4410,In_1682,In_1356);
or U4411 (N_4411,In_1596,In_716);
nor U4412 (N_4412,In_1818,In_2370);
nor U4413 (N_4413,In_79,In_1952);
xor U4414 (N_4414,In_1627,In_1562);
nor U4415 (N_4415,In_889,In_383);
and U4416 (N_4416,In_2294,In_1192);
or U4417 (N_4417,In_2099,In_1420);
nor U4418 (N_4418,In_692,In_1035);
or U4419 (N_4419,In_2222,In_1373);
and U4420 (N_4420,In_1234,In_782);
and U4421 (N_4421,In_1117,In_1003);
and U4422 (N_4422,In_1536,In_1614);
and U4423 (N_4423,In_2418,In_970);
nand U4424 (N_4424,In_329,In_325);
xor U4425 (N_4425,In_1242,In_2004);
or U4426 (N_4426,In_1725,In_1861);
nand U4427 (N_4427,In_200,In_1310);
and U4428 (N_4428,In_280,In_2431);
nand U4429 (N_4429,In_1771,In_367);
nor U4430 (N_4430,In_1280,In_1871);
xor U4431 (N_4431,In_1266,In_406);
and U4432 (N_4432,In_1184,In_491);
nor U4433 (N_4433,In_879,In_318);
xor U4434 (N_4434,In_1617,In_1815);
or U4435 (N_4435,In_712,In_0);
nand U4436 (N_4436,In_1141,In_1757);
nand U4437 (N_4437,In_253,In_1187);
nand U4438 (N_4438,In_1382,In_551);
nand U4439 (N_4439,In_2202,In_766);
or U4440 (N_4440,In_1352,In_2282);
xnor U4441 (N_4441,In_396,In_1393);
and U4442 (N_4442,In_1729,In_125);
or U4443 (N_4443,In_589,In_2249);
or U4444 (N_4444,In_2385,In_1167);
or U4445 (N_4445,In_571,In_1324);
and U4446 (N_4446,In_1505,In_529);
nand U4447 (N_4447,In_1040,In_129);
nand U4448 (N_4448,In_1803,In_558);
nand U4449 (N_4449,In_1707,In_1572);
nand U4450 (N_4450,In_1090,In_2049);
and U4451 (N_4451,In_569,In_803);
nor U4452 (N_4452,In_2052,In_275);
nor U4453 (N_4453,In_677,In_848);
nand U4454 (N_4454,In_1697,In_293);
nor U4455 (N_4455,In_2383,In_1222);
xnor U4456 (N_4456,In_792,In_1489);
nor U4457 (N_4457,In_1646,In_267);
nand U4458 (N_4458,In_1750,In_2161);
nand U4459 (N_4459,In_845,In_497);
xor U4460 (N_4460,In_1367,In_693);
nand U4461 (N_4461,In_152,In_1134);
and U4462 (N_4462,In_1549,In_1103);
and U4463 (N_4463,In_1125,In_829);
xnor U4464 (N_4464,In_1127,In_1183);
and U4465 (N_4465,In_1066,In_505);
xnor U4466 (N_4466,In_784,In_1539);
and U4467 (N_4467,In_707,In_2317);
or U4468 (N_4468,In_434,In_1254);
or U4469 (N_4469,In_331,In_1231);
or U4470 (N_4470,In_1260,In_473);
and U4471 (N_4471,In_241,In_261);
and U4472 (N_4472,In_1173,In_1342);
xnor U4473 (N_4473,In_1404,In_1420);
and U4474 (N_4474,In_594,In_833);
or U4475 (N_4475,In_1864,In_2163);
nor U4476 (N_4476,In_366,In_1072);
and U4477 (N_4477,In_76,In_1175);
xor U4478 (N_4478,In_342,In_844);
and U4479 (N_4479,In_282,In_1425);
and U4480 (N_4480,In_1757,In_1214);
and U4481 (N_4481,In_216,In_1827);
or U4482 (N_4482,In_465,In_1312);
and U4483 (N_4483,In_97,In_535);
nor U4484 (N_4484,In_603,In_2143);
xor U4485 (N_4485,In_1334,In_1471);
nand U4486 (N_4486,In_1013,In_395);
nand U4487 (N_4487,In_1826,In_146);
nor U4488 (N_4488,In_315,In_2177);
and U4489 (N_4489,In_1413,In_156);
nor U4490 (N_4490,In_344,In_2051);
nor U4491 (N_4491,In_2445,In_1359);
and U4492 (N_4492,In_201,In_814);
nand U4493 (N_4493,In_1495,In_2203);
and U4494 (N_4494,In_873,In_616);
nand U4495 (N_4495,In_1305,In_399);
or U4496 (N_4496,In_2117,In_2059);
nand U4497 (N_4497,In_2379,In_593);
or U4498 (N_4498,In_2489,In_2165);
or U4499 (N_4499,In_48,In_1092);
xnor U4500 (N_4500,In_741,In_638);
or U4501 (N_4501,In_1238,In_1743);
or U4502 (N_4502,In_1101,In_1285);
or U4503 (N_4503,In_102,In_1476);
nor U4504 (N_4504,In_1930,In_743);
nand U4505 (N_4505,In_523,In_1071);
nand U4506 (N_4506,In_747,In_1631);
and U4507 (N_4507,In_654,In_453);
nand U4508 (N_4508,In_1783,In_1377);
xor U4509 (N_4509,In_2363,In_301);
nand U4510 (N_4510,In_1048,In_2108);
and U4511 (N_4511,In_133,In_1529);
nor U4512 (N_4512,In_1120,In_92);
nor U4513 (N_4513,In_1147,In_307);
nor U4514 (N_4514,In_1823,In_2180);
or U4515 (N_4515,In_203,In_2142);
xor U4516 (N_4516,In_193,In_1757);
or U4517 (N_4517,In_2110,In_2417);
and U4518 (N_4518,In_2456,In_358);
and U4519 (N_4519,In_2139,In_2102);
xor U4520 (N_4520,In_258,In_767);
or U4521 (N_4521,In_1995,In_818);
or U4522 (N_4522,In_1977,In_961);
and U4523 (N_4523,In_1409,In_1906);
nor U4524 (N_4524,In_585,In_470);
and U4525 (N_4525,In_1334,In_660);
or U4526 (N_4526,In_968,In_1728);
or U4527 (N_4527,In_2420,In_1601);
and U4528 (N_4528,In_643,In_827);
or U4529 (N_4529,In_725,In_386);
or U4530 (N_4530,In_1226,In_1429);
or U4531 (N_4531,In_1581,In_425);
or U4532 (N_4532,In_319,In_304);
or U4533 (N_4533,In_100,In_2011);
nor U4534 (N_4534,In_2307,In_707);
nor U4535 (N_4535,In_2033,In_1448);
xnor U4536 (N_4536,In_1864,In_2406);
and U4537 (N_4537,In_1328,In_2348);
nor U4538 (N_4538,In_1736,In_1450);
nor U4539 (N_4539,In_2479,In_334);
nor U4540 (N_4540,In_200,In_2258);
nor U4541 (N_4541,In_406,In_669);
or U4542 (N_4542,In_1078,In_2244);
nor U4543 (N_4543,In_1086,In_913);
or U4544 (N_4544,In_1798,In_928);
nand U4545 (N_4545,In_674,In_1848);
nor U4546 (N_4546,In_1440,In_843);
or U4547 (N_4547,In_1614,In_2000);
nor U4548 (N_4548,In_1058,In_2106);
nand U4549 (N_4549,In_2156,In_305);
nand U4550 (N_4550,In_2442,In_2026);
nor U4551 (N_4551,In_2439,In_1090);
or U4552 (N_4552,In_1792,In_7);
and U4553 (N_4553,In_1449,In_197);
nor U4554 (N_4554,In_1707,In_2227);
or U4555 (N_4555,In_1595,In_2163);
nor U4556 (N_4556,In_2040,In_65);
nor U4557 (N_4557,In_1751,In_2041);
or U4558 (N_4558,In_449,In_271);
and U4559 (N_4559,In_1377,In_91);
or U4560 (N_4560,In_1393,In_795);
or U4561 (N_4561,In_526,In_643);
nand U4562 (N_4562,In_1221,In_1585);
or U4563 (N_4563,In_2143,In_1057);
and U4564 (N_4564,In_1426,In_2295);
or U4565 (N_4565,In_1794,In_1419);
nand U4566 (N_4566,In_1371,In_2060);
or U4567 (N_4567,In_1739,In_84);
and U4568 (N_4568,In_442,In_1164);
or U4569 (N_4569,In_717,In_952);
or U4570 (N_4570,In_287,In_1907);
nor U4571 (N_4571,In_2087,In_1995);
and U4572 (N_4572,In_457,In_1676);
and U4573 (N_4573,In_300,In_831);
nor U4574 (N_4574,In_159,In_608);
xnor U4575 (N_4575,In_96,In_587);
nor U4576 (N_4576,In_1110,In_791);
or U4577 (N_4577,In_2303,In_1546);
nand U4578 (N_4578,In_847,In_1075);
nand U4579 (N_4579,In_2078,In_872);
nand U4580 (N_4580,In_1802,In_2039);
or U4581 (N_4581,In_2290,In_780);
or U4582 (N_4582,In_2246,In_2146);
xnor U4583 (N_4583,In_1698,In_342);
nor U4584 (N_4584,In_1850,In_1465);
nor U4585 (N_4585,In_2075,In_348);
and U4586 (N_4586,In_30,In_177);
nor U4587 (N_4587,In_436,In_497);
or U4588 (N_4588,In_2173,In_783);
xnor U4589 (N_4589,In_1045,In_789);
and U4590 (N_4590,In_142,In_1610);
nand U4591 (N_4591,In_2166,In_178);
nor U4592 (N_4592,In_891,In_1146);
xnor U4593 (N_4593,In_333,In_1794);
nor U4594 (N_4594,In_2098,In_1759);
xnor U4595 (N_4595,In_1855,In_1120);
xor U4596 (N_4596,In_1086,In_84);
or U4597 (N_4597,In_1533,In_685);
nor U4598 (N_4598,In_1983,In_229);
nand U4599 (N_4599,In_1012,In_656);
xor U4600 (N_4600,In_1644,In_615);
and U4601 (N_4601,In_770,In_1750);
nand U4602 (N_4602,In_2051,In_477);
nor U4603 (N_4603,In_1447,In_1115);
nor U4604 (N_4604,In_2473,In_1694);
or U4605 (N_4605,In_1867,In_1828);
nor U4606 (N_4606,In_2283,In_1838);
xor U4607 (N_4607,In_1595,In_1055);
xor U4608 (N_4608,In_870,In_365);
and U4609 (N_4609,In_1144,In_820);
or U4610 (N_4610,In_616,In_2262);
xor U4611 (N_4611,In_505,In_885);
xnor U4612 (N_4612,In_772,In_1045);
nor U4613 (N_4613,In_1836,In_2400);
or U4614 (N_4614,In_1434,In_754);
and U4615 (N_4615,In_1295,In_1468);
nand U4616 (N_4616,In_234,In_1862);
or U4617 (N_4617,In_678,In_1699);
nor U4618 (N_4618,In_2192,In_200);
nor U4619 (N_4619,In_1402,In_2067);
nand U4620 (N_4620,In_2281,In_210);
nor U4621 (N_4621,In_60,In_966);
or U4622 (N_4622,In_1023,In_1650);
and U4623 (N_4623,In_1625,In_171);
nor U4624 (N_4624,In_1925,In_14);
and U4625 (N_4625,In_1280,In_1197);
and U4626 (N_4626,In_1342,In_336);
and U4627 (N_4627,In_2182,In_1085);
nor U4628 (N_4628,In_2035,In_1420);
nand U4629 (N_4629,In_264,In_2057);
nor U4630 (N_4630,In_1573,In_385);
nand U4631 (N_4631,In_309,In_2368);
and U4632 (N_4632,In_1387,In_2471);
nand U4633 (N_4633,In_2357,In_2354);
xor U4634 (N_4634,In_1521,In_390);
and U4635 (N_4635,In_284,In_1047);
xor U4636 (N_4636,In_491,In_1049);
nor U4637 (N_4637,In_1983,In_827);
nand U4638 (N_4638,In_2498,In_1554);
or U4639 (N_4639,In_1365,In_1373);
nand U4640 (N_4640,In_1113,In_1013);
or U4641 (N_4641,In_463,In_2449);
or U4642 (N_4642,In_1119,In_10);
nand U4643 (N_4643,In_2217,In_67);
or U4644 (N_4644,In_966,In_242);
or U4645 (N_4645,In_842,In_1436);
nor U4646 (N_4646,In_1264,In_1490);
nor U4647 (N_4647,In_525,In_1929);
or U4648 (N_4648,In_195,In_1120);
nor U4649 (N_4649,In_1630,In_2143);
nor U4650 (N_4650,In_1202,In_837);
nor U4651 (N_4651,In_779,In_1718);
and U4652 (N_4652,In_1969,In_1044);
and U4653 (N_4653,In_1733,In_1209);
or U4654 (N_4654,In_2092,In_318);
and U4655 (N_4655,In_889,In_76);
nor U4656 (N_4656,In_468,In_903);
and U4657 (N_4657,In_194,In_617);
or U4658 (N_4658,In_1145,In_2417);
or U4659 (N_4659,In_2228,In_997);
and U4660 (N_4660,In_1982,In_633);
xnor U4661 (N_4661,In_165,In_2145);
and U4662 (N_4662,In_1217,In_88);
nand U4663 (N_4663,In_2231,In_1539);
or U4664 (N_4664,In_772,In_1443);
or U4665 (N_4665,In_297,In_2092);
or U4666 (N_4666,In_266,In_1703);
nand U4667 (N_4667,In_1133,In_2351);
and U4668 (N_4668,In_4,In_835);
nor U4669 (N_4669,In_1779,In_790);
and U4670 (N_4670,In_785,In_118);
nor U4671 (N_4671,In_307,In_1792);
xor U4672 (N_4672,In_202,In_2042);
and U4673 (N_4673,In_1358,In_2266);
xnor U4674 (N_4674,In_838,In_1575);
xnor U4675 (N_4675,In_1678,In_556);
and U4676 (N_4676,In_1423,In_2212);
xnor U4677 (N_4677,In_1284,In_1494);
and U4678 (N_4678,In_2172,In_2101);
or U4679 (N_4679,In_272,In_1168);
nor U4680 (N_4680,In_1372,In_856);
xnor U4681 (N_4681,In_1303,In_1533);
nand U4682 (N_4682,In_624,In_1926);
or U4683 (N_4683,In_1865,In_2409);
nor U4684 (N_4684,In_68,In_1888);
xnor U4685 (N_4685,In_1389,In_1560);
nand U4686 (N_4686,In_938,In_554);
or U4687 (N_4687,In_2138,In_1869);
and U4688 (N_4688,In_2483,In_1422);
nand U4689 (N_4689,In_2267,In_1162);
nor U4690 (N_4690,In_2457,In_344);
or U4691 (N_4691,In_946,In_1877);
nor U4692 (N_4692,In_745,In_2433);
nor U4693 (N_4693,In_2170,In_587);
and U4694 (N_4694,In_1179,In_1511);
or U4695 (N_4695,In_49,In_161);
nand U4696 (N_4696,In_2392,In_1773);
xor U4697 (N_4697,In_567,In_143);
xnor U4698 (N_4698,In_1285,In_419);
nor U4699 (N_4699,In_430,In_2137);
nand U4700 (N_4700,In_1636,In_279);
xnor U4701 (N_4701,In_658,In_627);
and U4702 (N_4702,In_464,In_57);
nor U4703 (N_4703,In_2382,In_1700);
xor U4704 (N_4704,In_846,In_910);
and U4705 (N_4705,In_2196,In_259);
xnor U4706 (N_4706,In_1582,In_1822);
nand U4707 (N_4707,In_2173,In_1289);
nor U4708 (N_4708,In_1581,In_2058);
nand U4709 (N_4709,In_303,In_1581);
or U4710 (N_4710,In_1264,In_382);
or U4711 (N_4711,In_101,In_1208);
or U4712 (N_4712,In_2092,In_2120);
nand U4713 (N_4713,In_1409,In_2486);
nor U4714 (N_4714,In_1393,In_2137);
or U4715 (N_4715,In_2318,In_1605);
and U4716 (N_4716,In_1436,In_556);
nand U4717 (N_4717,In_213,In_2006);
xnor U4718 (N_4718,In_1857,In_321);
and U4719 (N_4719,In_1218,In_1751);
nand U4720 (N_4720,In_2307,In_795);
or U4721 (N_4721,In_1961,In_729);
and U4722 (N_4722,In_1122,In_682);
or U4723 (N_4723,In_1966,In_2336);
or U4724 (N_4724,In_469,In_948);
or U4725 (N_4725,In_1694,In_2135);
xor U4726 (N_4726,In_1378,In_1408);
nand U4727 (N_4727,In_1208,In_1044);
nand U4728 (N_4728,In_1248,In_359);
nor U4729 (N_4729,In_1897,In_2172);
nor U4730 (N_4730,In_712,In_2189);
nand U4731 (N_4731,In_1157,In_341);
xor U4732 (N_4732,In_1553,In_1308);
or U4733 (N_4733,In_2358,In_318);
nand U4734 (N_4734,In_1777,In_689);
and U4735 (N_4735,In_2464,In_1613);
nand U4736 (N_4736,In_633,In_360);
or U4737 (N_4737,In_1256,In_322);
or U4738 (N_4738,In_1954,In_1030);
xnor U4739 (N_4739,In_603,In_620);
xor U4740 (N_4740,In_470,In_405);
or U4741 (N_4741,In_858,In_2482);
or U4742 (N_4742,In_2344,In_684);
and U4743 (N_4743,In_1667,In_1834);
or U4744 (N_4744,In_1429,In_1283);
xnor U4745 (N_4745,In_29,In_1815);
xnor U4746 (N_4746,In_1200,In_154);
nand U4747 (N_4747,In_72,In_1836);
xnor U4748 (N_4748,In_253,In_1314);
nor U4749 (N_4749,In_45,In_2383);
and U4750 (N_4750,In_1277,In_678);
nand U4751 (N_4751,In_962,In_266);
nor U4752 (N_4752,In_2399,In_350);
or U4753 (N_4753,In_1155,In_2244);
or U4754 (N_4754,In_2078,In_2025);
nand U4755 (N_4755,In_2013,In_502);
nor U4756 (N_4756,In_1645,In_1989);
nor U4757 (N_4757,In_2037,In_2294);
nor U4758 (N_4758,In_1643,In_47);
and U4759 (N_4759,In_1298,In_1862);
xnor U4760 (N_4760,In_947,In_470);
nor U4761 (N_4761,In_2270,In_628);
nand U4762 (N_4762,In_714,In_1880);
and U4763 (N_4763,In_1034,In_1688);
nor U4764 (N_4764,In_2279,In_1838);
xnor U4765 (N_4765,In_623,In_332);
and U4766 (N_4766,In_445,In_1977);
xor U4767 (N_4767,In_2386,In_2057);
nand U4768 (N_4768,In_2130,In_2156);
xnor U4769 (N_4769,In_159,In_1114);
and U4770 (N_4770,In_289,In_1925);
xor U4771 (N_4771,In_1114,In_2281);
nand U4772 (N_4772,In_1894,In_1233);
xor U4773 (N_4773,In_658,In_1030);
and U4774 (N_4774,In_694,In_635);
xnor U4775 (N_4775,In_1289,In_2144);
nand U4776 (N_4776,In_1457,In_2287);
nor U4777 (N_4777,In_66,In_612);
or U4778 (N_4778,In_1944,In_1224);
nor U4779 (N_4779,In_2484,In_1557);
and U4780 (N_4780,In_658,In_1741);
and U4781 (N_4781,In_1271,In_1775);
nor U4782 (N_4782,In_1442,In_373);
nand U4783 (N_4783,In_2468,In_195);
nor U4784 (N_4784,In_260,In_920);
xnor U4785 (N_4785,In_183,In_2056);
nand U4786 (N_4786,In_1806,In_980);
nand U4787 (N_4787,In_1331,In_1844);
nor U4788 (N_4788,In_642,In_112);
nand U4789 (N_4789,In_2166,In_656);
nor U4790 (N_4790,In_760,In_1803);
nor U4791 (N_4791,In_1881,In_1673);
and U4792 (N_4792,In_1843,In_108);
xor U4793 (N_4793,In_1232,In_1417);
or U4794 (N_4794,In_1616,In_557);
nand U4795 (N_4795,In_929,In_2314);
and U4796 (N_4796,In_2381,In_1482);
xnor U4797 (N_4797,In_1429,In_905);
and U4798 (N_4798,In_1480,In_662);
and U4799 (N_4799,In_2484,In_120);
nand U4800 (N_4800,In_109,In_914);
nand U4801 (N_4801,In_59,In_830);
nand U4802 (N_4802,In_2432,In_1209);
or U4803 (N_4803,In_2420,In_1986);
xor U4804 (N_4804,In_2296,In_354);
or U4805 (N_4805,In_1248,In_457);
xor U4806 (N_4806,In_1138,In_1310);
and U4807 (N_4807,In_1186,In_788);
nor U4808 (N_4808,In_457,In_895);
xnor U4809 (N_4809,In_1192,In_544);
or U4810 (N_4810,In_1038,In_1530);
nor U4811 (N_4811,In_1912,In_1609);
or U4812 (N_4812,In_648,In_1351);
and U4813 (N_4813,In_63,In_1953);
xor U4814 (N_4814,In_463,In_1786);
nor U4815 (N_4815,In_618,In_1512);
or U4816 (N_4816,In_444,In_1843);
xor U4817 (N_4817,In_2422,In_2378);
nor U4818 (N_4818,In_2221,In_1213);
nand U4819 (N_4819,In_1116,In_914);
nand U4820 (N_4820,In_1350,In_280);
nor U4821 (N_4821,In_1379,In_795);
xnor U4822 (N_4822,In_1114,In_1218);
and U4823 (N_4823,In_958,In_1423);
nor U4824 (N_4824,In_1331,In_317);
xnor U4825 (N_4825,In_765,In_606);
nand U4826 (N_4826,In_2189,In_525);
xnor U4827 (N_4827,In_619,In_463);
or U4828 (N_4828,In_1817,In_658);
xor U4829 (N_4829,In_225,In_2285);
and U4830 (N_4830,In_1899,In_1853);
nand U4831 (N_4831,In_2213,In_1632);
xnor U4832 (N_4832,In_1039,In_1815);
or U4833 (N_4833,In_1512,In_1753);
nand U4834 (N_4834,In_1791,In_1160);
nor U4835 (N_4835,In_305,In_1716);
and U4836 (N_4836,In_458,In_386);
nor U4837 (N_4837,In_2099,In_772);
and U4838 (N_4838,In_178,In_1663);
xor U4839 (N_4839,In_810,In_422);
or U4840 (N_4840,In_432,In_472);
or U4841 (N_4841,In_531,In_1035);
nand U4842 (N_4842,In_32,In_47);
or U4843 (N_4843,In_169,In_2484);
xnor U4844 (N_4844,In_1935,In_874);
nand U4845 (N_4845,In_1941,In_1505);
and U4846 (N_4846,In_2299,In_1755);
nor U4847 (N_4847,In_1197,In_906);
nor U4848 (N_4848,In_1144,In_1046);
nand U4849 (N_4849,In_786,In_1223);
and U4850 (N_4850,In_1008,In_482);
nand U4851 (N_4851,In_2128,In_2160);
or U4852 (N_4852,In_274,In_956);
xnor U4853 (N_4853,In_1599,In_1013);
nand U4854 (N_4854,In_537,In_1460);
nor U4855 (N_4855,In_1540,In_62);
nand U4856 (N_4856,In_1508,In_196);
xor U4857 (N_4857,In_2174,In_2357);
nor U4858 (N_4858,In_2258,In_342);
or U4859 (N_4859,In_2198,In_1813);
and U4860 (N_4860,In_169,In_423);
nand U4861 (N_4861,In_950,In_1023);
or U4862 (N_4862,In_386,In_2301);
nand U4863 (N_4863,In_391,In_2169);
xor U4864 (N_4864,In_1438,In_2115);
and U4865 (N_4865,In_1569,In_296);
xor U4866 (N_4866,In_2086,In_202);
or U4867 (N_4867,In_1137,In_776);
and U4868 (N_4868,In_844,In_584);
and U4869 (N_4869,In_28,In_840);
xor U4870 (N_4870,In_818,In_729);
or U4871 (N_4871,In_1155,In_1147);
xnor U4872 (N_4872,In_2415,In_923);
xor U4873 (N_4873,In_326,In_1424);
xor U4874 (N_4874,In_760,In_899);
nor U4875 (N_4875,In_2132,In_1200);
or U4876 (N_4876,In_1087,In_444);
nand U4877 (N_4877,In_1603,In_154);
and U4878 (N_4878,In_918,In_1764);
nor U4879 (N_4879,In_1706,In_278);
or U4880 (N_4880,In_1165,In_1335);
or U4881 (N_4881,In_864,In_1228);
or U4882 (N_4882,In_1498,In_541);
nor U4883 (N_4883,In_608,In_1794);
nand U4884 (N_4884,In_242,In_572);
or U4885 (N_4885,In_2444,In_2474);
and U4886 (N_4886,In_732,In_909);
xor U4887 (N_4887,In_1341,In_807);
and U4888 (N_4888,In_2399,In_1736);
nand U4889 (N_4889,In_1558,In_351);
nand U4890 (N_4890,In_1884,In_2228);
or U4891 (N_4891,In_1779,In_394);
or U4892 (N_4892,In_1030,In_298);
and U4893 (N_4893,In_1979,In_239);
or U4894 (N_4894,In_1101,In_2186);
or U4895 (N_4895,In_2034,In_2271);
and U4896 (N_4896,In_1402,In_516);
and U4897 (N_4897,In_1192,In_1849);
nand U4898 (N_4898,In_605,In_85);
nand U4899 (N_4899,In_2463,In_1602);
xnor U4900 (N_4900,In_1103,In_1544);
xor U4901 (N_4901,In_2443,In_459);
nor U4902 (N_4902,In_1895,In_58);
or U4903 (N_4903,In_1059,In_524);
and U4904 (N_4904,In_1117,In_915);
or U4905 (N_4905,In_1892,In_605);
or U4906 (N_4906,In_2319,In_1791);
or U4907 (N_4907,In_2064,In_674);
xor U4908 (N_4908,In_2268,In_1613);
nor U4909 (N_4909,In_2487,In_1657);
nor U4910 (N_4910,In_1198,In_1733);
and U4911 (N_4911,In_696,In_1313);
and U4912 (N_4912,In_2296,In_2069);
xor U4913 (N_4913,In_370,In_2459);
nor U4914 (N_4914,In_1495,In_2284);
xor U4915 (N_4915,In_1393,In_1165);
xor U4916 (N_4916,In_2306,In_1918);
nor U4917 (N_4917,In_49,In_1207);
and U4918 (N_4918,In_810,In_218);
nand U4919 (N_4919,In_2387,In_1508);
nand U4920 (N_4920,In_2245,In_1573);
or U4921 (N_4921,In_1144,In_1208);
nor U4922 (N_4922,In_1334,In_43);
or U4923 (N_4923,In_1350,In_2044);
nor U4924 (N_4924,In_2122,In_1931);
xnor U4925 (N_4925,In_973,In_1327);
and U4926 (N_4926,In_1664,In_2159);
nor U4927 (N_4927,In_1973,In_1493);
or U4928 (N_4928,In_202,In_56);
xnor U4929 (N_4929,In_2094,In_752);
xnor U4930 (N_4930,In_676,In_1861);
and U4931 (N_4931,In_13,In_838);
and U4932 (N_4932,In_1542,In_1701);
and U4933 (N_4933,In_1788,In_2370);
or U4934 (N_4934,In_2230,In_249);
xnor U4935 (N_4935,In_469,In_390);
and U4936 (N_4936,In_953,In_285);
or U4937 (N_4937,In_1932,In_108);
xor U4938 (N_4938,In_699,In_471);
nand U4939 (N_4939,In_890,In_1264);
nor U4940 (N_4940,In_1505,In_1154);
or U4941 (N_4941,In_13,In_971);
and U4942 (N_4942,In_2058,In_930);
nor U4943 (N_4943,In_2087,In_1625);
nand U4944 (N_4944,In_1135,In_94);
xnor U4945 (N_4945,In_1328,In_1774);
or U4946 (N_4946,In_874,In_785);
xnor U4947 (N_4947,In_2288,In_929);
or U4948 (N_4948,In_270,In_1592);
xnor U4949 (N_4949,In_654,In_1345);
or U4950 (N_4950,In_94,In_2057);
and U4951 (N_4951,In_2255,In_908);
and U4952 (N_4952,In_2005,In_2157);
or U4953 (N_4953,In_1811,In_816);
and U4954 (N_4954,In_2343,In_612);
xnor U4955 (N_4955,In_1694,In_947);
and U4956 (N_4956,In_25,In_1513);
nor U4957 (N_4957,In_1307,In_1582);
xnor U4958 (N_4958,In_480,In_471);
or U4959 (N_4959,In_1937,In_1587);
nor U4960 (N_4960,In_575,In_2135);
or U4961 (N_4961,In_1810,In_1108);
or U4962 (N_4962,In_788,In_1832);
nand U4963 (N_4963,In_1196,In_339);
xor U4964 (N_4964,In_1717,In_413);
nor U4965 (N_4965,In_1303,In_1501);
or U4966 (N_4966,In_1083,In_2192);
xor U4967 (N_4967,In_834,In_2255);
xor U4968 (N_4968,In_2428,In_199);
xnor U4969 (N_4969,In_404,In_2295);
and U4970 (N_4970,In_1574,In_791);
nand U4971 (N_4971,In_1554,In_888);
nand U4972 (N_4972,In_259,In_1639);
and U4973 (N_4973,In_329,In_1975);
or U4974 (N_4974,In_491,In_2480);
nor U4975 (N_4975,In_761,In_1471);
nand U4976 (N_4976,In_1768,In_641);
nor U4977 (N_4977,In_1184,In_587);
nand U4978 (N_4978,In_1129,In_396);
or U4979 (N_4979,In_729,In_728);
nand U4980 (N_4980,In_360,In_703);
or U4981 (N_4981,In_1094,In_2340);
and U4982 (N_4982,In_2143,In_423);
or U4983 (N_4983,In_2457,In_1768);
or U4984 (N_4984,In_1606,In_2052);
or U4985 (N_4985,In_653,In_1066);
or U4986 (N_4986,In_33,In_743);
and U4987 (N_4987,In_274,In_951);
nor U4988 (N_4988,In_810,In_1091);
nand U4989 (N_4989,In_1762,In_2152);
nand U4990 (N_4990,In_2101,In_368);
or U4991 (N_4991,In_1879,In_1121);
xnor U4992 (N_4992,In_90,In_1317);
nor U4993 (N_4993,In_1455,In_2380);
xnor U4994 (N_4994,In_2484,In_1060);
and U4995 (N_4995,In_2211,In_1655);
and U4996 (N_4996,In_1328,In_1745);
nand U4997 (N_4997,In_42,In_12);
nor U4998 (N_4998,In_710,In_1804);
xnor U4999 (N_4999,In_645,In_1915);
nor U5000 (N_5000,N_1193,N_1332);
xnor U5001 (N_5001,N_497,N_297);
nand U5002 (N_5002,N_4808,N_2507);
nor U5003 (N_5003,N_1753,N_1173);
and U5004 (N_5004,N_4497,N_663);
xor U5005 (N_5005,N_1300,N_2910);
xnor U5006 (N_5006,N_3019,N_2562);
or U5007 (N_5007,N_2086,N_1172);
nand U5008 (N_5008,N_706,N_1983);
nand U5009 (N_5009,N_2206,N_2463);
and U5010 (N_5010,N_1096,N_4614);
xnor U5011 (N_5011,N_1415,N_4721);
nand U5012 (N_5012,N_2754,N_2572);
nand U5013 (N_5013,N_3915,N_4225);
nor U5014 (N_5014,N_3588,N_4233);
and U5015 (N_5015,N_2947,N_664);
nand U5016 (N_5016,N_4561,N_2822);
nor U5017 (N_5017,N_2743,N_236);
and U5018 (N_5018,N_2324,N_4547);
xor U5019 (N_5019,N_3168,N_3766);
nand U5020 (N_5020,N_4610,N_371);
xor U5021 (N_5021,N_1842,N_98);
nand U5022 (N_5022,N_1976,N_2759);
or U5023 (N_5023,N_112,N_3305);
and U5024 (N_5024,N_1135,N_3602);
nor U5025 (N_5025,N_3357,N_2081);
or U5026 (N_5026,N_567,N_3180);
nand U5027 (N_5027,N_528,N_3798);
or U5028 (N_5028,N_515,N_2912);
xnor U5029 (N_5029,N_3010,N_2604);
nand U5030 (N_5030,N_4831,N_3757);
nor U5031 (N_5031,N_4968,N_1065);
or U5032 (N_5032,N_3770,N_1245);
or U5033 (N_5033,N_44,N_4403);
or U5034 (N_5034,N_2127,N_2727);
nand U5035 (N_5035,N_352,N_4441);
or U5036 (N_5036,N_819,N_3254);
nor U5037 (N_5037,N_388,N_2358);
or U5038 (N_5038,N_4907,N_2907);
or U5039 (N_5039,N_3186,N_517);
xnor U5040 (N_5040,N_601,N_1435);
nor U5041 (N_5041,N_2030,N_1267);
nand U5042 (N_5042,N_1940,N_1461);
and U5043 (N_5043,N_662,N_4582);
and U5044 (N_5044,N_3153,N_1880);
and U5045 (N_5045,N_918,N_4733);
nor U5046 (N_5046,N_3948,N_3999);
nand U5047 (N_5047,N_1911,N_4558);
nor U5048 (N_5048,N_4608,N_2034);
nor U5049 (N_5049,N_3835,N_4754);
and U5050 (N_5050,N_2270,N_2342);
or U5051 (N_5051,N_877,N_4103);
xnor U5052 (N_5052,N_3709,N_250);
nor U5053 (N_5053,N_999,N_892);
nand U5054 (N_5054,N_3860,N_2302);
or U5055 (N_5055,N_1817,N_1353);
nand U5056 (N_5056,N_2273,N_874);
xor U5057 (N_5057,N_4868,N_990);
xnor U5058 (N_5058,N_4650,N_3544);
or U5059 (N_5059,N_4259,N_4163);
or U5060 (N_5060,N_4605,N_1177);
nor U5061 (N_5061,N_271,N_657);
nand U5062 (N_5062,N_2343,N_3490);
and U5063 (N_5063,N_0,N_2462);
nand U5064 (N_5064,N_249,N_2811);
nor U5065 (N_5065,N_2998,N_3997);
nor U5066 (N_5066,N_3464,N_153);
xor U5067 (N_5067,N_4056,N_1071);
xnor U5068 (N_5068,N_3515,N_1971);
nor U5069 (N_5069,N_2381,N_4176);
xor U5070 (N_5070,N_2646,N_4729);
or U5071 (N_5071,N_4366,N_1199);
nor U5072 (N_5072,N_1164,N_3146);
and U5073 (N_5073,N_3197,N_3669);
xnor U5074 (N_5074,N_356,N_2055);
nor U5075 (N_5075,N_1969,N_2064);
xor U5076 (N_5076,N_597,N_4293);
nand U5077 (N_5077,N_474,N_2684);
nor U5078 (N_5078,N_2746,N_855);
nor U5079 (N_5079,N_4381,N_4736);
xnor U5080 (N_5080,N_45,N_1308);
xnor U5081 (N_5081,N_4095,N_1997);
xnor U5082 (N_5082,N_3039,N_2103);
and U5083 (N_5083,N_703,N_2515);
xnor U5084 (N_5084,N_4182,N_4632);
xor U5085 (N_5085,N_2609,N_4607);
or U5086 (N_5086,N_4150,N_3514);
and U5087 (N_5087,N_133,N_978);
or U5088 (N_5088,N_274,N_4580);
xnor U5089 (N_5089,N_1121,N_4322);
nor U5090 (N_5090,N_1742,N_4341);
nand U5091 (N_5091,N_50,N_3119);
and U5092 (N_5092,N_4778,N_3346);
or U5093 (N_5093,N_3638,N_3616);
nand U5094 (N_5094,N_408,N_750);
or U5095 (N_5095,N_2553,N_132);
xor U5096 (N_5096,N_1212,N_862);
and U5097 (N_5097,N_3995,N_4804);
xnor U5098 (N_5098,N_4200,N_3540);
and U5099 (N_5099,N_839,N_1347);
or U5100 (N_5100,N_796,N_1662);
nand U5101 (N_5101,N_4207,N_749);
nand U5102 (N_5102,N_4934,N_4890);
or U5103 (N_5103,N_4058,N_4642);
xnor U5104 (N_5104,N_1740,N_1496);
nand U5105 (N_5105,N_3430,N_4395);
and U5106 (N_5106,N_287,N_1034);
nand U5107 (N_5107,N_852,N_3134);
and U5108 (N_5108,N_3319,N_2292);
xnor U5109 (N_5109,N_4107,N_4476);
nor U5110 (N_5110,N_4284,N_1312);
nor U5111 (N_5111,N_1592,N_1925);
or U5112 (N_5112,N_1487,N_2079);
or U5113 (N_5113,N_1543,N_4555);
nor U5114 (N_5114,N_396,N_2364);
nand U5115 (N_5115,N_3905,N_123);
and U5116 (N_5116,N_4835,N_1708);
and U5117 (N_5117,N_970,N_3608);
and U5118 (N_5118,N_816,N_806);
nand U5119 (N_5119,N_2368,N_155);
xor U5120 (N_5120,N_3362,N_2038);
xor U5121 (N_5121,N_679,N_4922);
or U5122 (N_5122,N_3879,N_4459);
nand U5123 (N_5123,N_4693,N_1362);
nor U5124 (N_5124,N_2047,N_3828);
nor U5125 (N_5125,N_4826,N_4675);
xor U5126 (N_5126,N_2724,N_110);
nor U5127 (N_5127,N_3469,N_307);
nand U5128 (N_5128,N_223,N_508);
nand U5129 (N_5129,N_4572,N_2330);
and U5130 (N_5130,N_2471,N_797);
xor U5131 (N_5131,N_1499,N_3106);
or U5132 (N_5132,N_3491,N_351);
nor U5133 (N_5133,N_1946,N_1115);
and U5134 (N_5134,N_4914,N_4856);
nor U5135 (N_5135,N_4997,N_3715);
xnor U5136 (N_5136,N_4251,N_1625);
or U5137 (N_5137,N_606,N_808);
nand U5138 (N_5138,N_4453,N_2749);
or U5139 (N_5139,N_3800,N_1399);
nand U5140 (N_5140,N_4878,N_1994);
and U5141 (N_5141,N_678,N_3893);
nor U5142 (N_5142,N_4113,N_1766);
and U5143 (N_5143,N_926,N_1989);
xor U5144 (N_5144,N_947,N_4475);
and U5145 (N_5145,N_730,N_4981);
xnor U5146 (N_5146,N_2989,N_1931);
and U5147 (N_5147,N_1757,N_3269);
nor U5148 (N_5148,N_3143,N_3156);
or U5149 (N_5149,N_3232,N_1980);
xor U5150 (N_5150,N_290,N_2802);
nor U5151 (N_5151,N_192,N_804);
nand U5152 (N_5152,N_183,N_2964);
xor U5153 (N_5153,N_2588,N_2888);
xnor U5154 (N_5154,N_1908,N_2493);
xnor U5155 (N_5155,N_1301,N_1630);
xor U5156 (N_5156,N_910,N_1844);
nand U5157 (N_5157,N_1862,N_2542);
nor U5158 (N_5158,N_2044,N_1137);
nand U5159 (N_5159,N_1049,N_3850);
and U5160 (N_5160,N_848,N_716);
xnor U5161 (N_5161,N_4101,N_1785);
or U5162 (N_5162,N_1494,N_4351);
xnor U5163 (N_5163,N_4513,N_361);
and U5164 (N_5164,N_1101,N_3301);
nand U5165 (N_5165,N_2495,N_4481);
nor U5166 (N_5166,N_1829,N_4278);
nor U5167 (N_5167,N_4415,N_437);
and U5168 (N_5168,N_824,N_4119);
nand U5169 (N_5169,N_2382,N_770);
nand U5170 (N_5170,N_3685,N_2611);
or U5171 (N_5171,N_3023,N_1944);
and U5172 (N_5172,N_4483,N_232);
xnor U5173 (N_5173,N_717,N_4390);
nor U5174 (N_5174,N_1040,N_1967);
or U5175 (N_5175,N_2862,N_1283);
or U5176 (N_5176,N_4719,N_196);
nor U5177 (N_5177,N_1070,N_1392);
nor U5178 (N_5178,N_1787,N_1006);
nor U5179 (N_5179,N_4815,N_2234);
nor U5180 (N_5180,N_36,N_91);
nor U5181 (N_5181,N_2657,N_2698);
nand U5182 (N_5182,N_4268,N_3922);
or U5183 (N_5183,N_4557,N_1727);
xor U5184 (N_5184,N_540,N_4140);
nand U5185 (N_5185,N_4895,N_3107);
and U5186 (N_5186,N_3159,N_4179);
nor U5187 (N_5187,N_4175,N_1521);
xnor U5188 (N_5188,N_2735,N_1603);
nor U5189 (N_5189,N_1018,N_4180);
or U5190 (N_5190,N_379,N_284);
nand U5191 (N_5191,N_3916,N_3487);
nor U5192 (N_5192,N_3006,N_3007);
xor U5193 (N_5193,N_680,N_1161);
nand U5194 (N_5194,N_2530,N_1036);
and U5195 (N_5195,N_511,N_1390);
nor U5196 (N_5196,N_1002,N_4944);
xnor U5197 (N_5197,N_1935,N_1743);
and U5198 (N_5198,N_2610,N_1099);
or U5199 (N_5199,N_519,N_4703);
or U5200 (N_5200,N_4374,N_4325);
and U5201 (N_5201,N_4688,N_60);
or U5202 (N_5202,N_1821,N_1500);
xor U5203 (N_5203,N_4857,N_2316);
xor U5204 (N_5204,N_2080,N_1294);
or U5205 (N_5205,N_2601,N_3118);
xor U5206 (N_5206,N_3804,N_3943);
nor U5207 (N_5207,N_2276,N_4346);
and U5208 (N_5208,N_46,N_4683);
nand U5209 (N_5209,N_2459,N_1641);
xnor U5210 (N_5210,N_2250,N_3355);
nand U5211 (N_5211,N_1827,N_3574);
xnor U5212 (N_5212,N_4108,N_4472);
or U5213 (N_5213,N_4774,N_2804);
nor U5214 (N_5214,N_1030,N_2776);
nand U5215 (N_5215,N_1277,N_482);
xnor U5216 (N_5216,N_3296,N_1819);
nor U5217 (N_5217,N_368,N_4256);
nand U5218 (N_5218,N_269,N_1850);
or U5219 (N_5219,N_4811,N_1326);
and U5220 (N_5220,N_230,N_2446);
nor U5221 (N_5221,N_2496,N_4963);
xnor U5222 (N_5222,N_4442,N_4541);
nand U5223 (N_5223,N_4131,N_3421);
nor U5224 (N_5224,N_201,N_3891);
nor U5225 (N_5225,N_3960,N_3216);
or U5226 (N_5226,N_3837,N_4885);
nand U5227 (N_5227,N_849,N_2997);
nor U5228 (N_5228,N_383,N_2608);
nor U5229 (N_5229,N_596,N_3295);
or U5230 (N_5230,N_3895,N_988);
and U5231 (N_5231,N_996,N_1810);
and U5232 (N_5232,N_1473,N_602);
xnor U5233 (N_5233,N_2213,N_3687);
or U5234 (N_5234,N_4559,N_2356);
nor U5235 (N_5235,N_835,N_4470);
xor U5236 (N_5236,N_1108,N_1576);
or U5237 (N_5237,N_2453,N_260);
nand U5238 (N_5238,N_4518,N_579);
xor U5239 (N_5239,N_4957,N_3692);
and U5240 (N_5240,N_1462,N_2875);
xnor U5241 (N_5241,N_1750,N_3397);
or U5242 (N_5242,N_3841,N_3273);
and U5243 (N_5243,N_1234,N_4405);
nand U5244 (N_5244,N_1680,N_4170);
and U5245 (N_5245,N_2879,N_2991);
or U5246 (N_5246,N_4964,N_1544);
xor U5247 (N_5247,N_1755,N_1875);
or U5248 (N_5248,N_479,N_413);
or U5249 (N_5249,N_2861,N_4508);
or U5250 (N_5250,N_3055,N_2181);
xor U5251 (N_5251,N_3166,N_2265);
or U5252 (N_5252,N_2001,N_3827);
and U5253 (N_5253,N_1444,N_1736);
or U5254 (N_5254,N_2674,N_1688);
and U5255 (N_5255,N_1586,N_2826);
or U5256 (N_5256,N_3548,N_4905);
nor U5257 (N_5257,N_4660,N_647);
nor U5258 (N_5258,N_247,N_3356);
xnor U5259 (N_5259,N_4297,N_377);
xnor U5260 (N_5260,N_401,N_3767);
or U5261 (N_5261,N_1182,N_2742);
nand U5262 (N_5262,N_3476,N_3780);
nand U5263 (N_5263,N_3625,N_2501);
or U5264 (N_5264,N_3512,N_1606);
or U5265 (N_5265,N_1329,N_292);
or U5266 (N_5266,N_3302,N_4375);
or U5267 (N_5267,N_720,N_2550);
xor U5268 (N_5268,N_4564,N_1163);
or U5269 (N_5269,N_3676,N_2426);
xor U5270 (N_5270,N_3130,N_3103);
nor U5271 (N_5271,N_4621,N_2868);
nor U5272 (N_5272,N_4234,N_4389);
nand U5273 (N_5273,N_2685,N_2993);
and U5274 (N_5274,N_2143,N_3444);
nand U5275 (N_5275,N_2720,N_618);
xnor U5276 (N_5276,N_3405,N_4);
nor U5277 (N_5277,N_886,N_1056);
xor U5278 (N_5278,N_4120,N_2218);
nor U5279 (N_5279,N_2896,N_3152);
xnor U5280 (N_5280,N_293,N_2622);
nor U5281 (N_5281,N_3101,N_2521);
nand U5282 (N_5282,N_870,N_860);
nand U5283 (N_5283,N_3223,N_4695);
and U5284 (N_5284,N_4926,N_3597);
nor U5285 (N_5285,N_4345,N_635);
nor U5286 (N_5286,N_424,N_3084);
nand U5287 (N_5287,N_2014,N_1644);
nand U5288 (N_5288,N_2546,N_4362);
xor U5289 (N_5289,N_2642,N_2526);
xor U5290 (N_5290,N_4332,N_4622);
or U5291 (N_5291,N_4039,N_1781);
xor U5292 (N_5292,N_2536,N_3598);
nor U5293 (N_5293,N_4370,N_4435);
nand U5294 (N_5294,N_4872,N_1721);
xnor U5295 (N_5295,N_4024,N_4059);
and U5296 (N_5296,N_2589,N_4333);
nand U5297 (N_5297,N_2728,N_908);
and U5298 (N_5298,N_2543,N_4277);
and U5299 (N_5299,N_4275,N_551);
xnor U5300 (N_5300,N_2154,N_215);
xnor U5301 (N_5301,N_117,N_3198);
xnor U5302 (N_5302,N_1713,N_1367);
and U5303 (N_5303,N_4003,N_3163);
xnor U5304 (N_5304,N_1229,N_3516);
nor U5305 (N_5305,N_3316,N_2114);
and U5306 (N_5306,N_4576,N_100);
nor U5307 (N_5307,N_4080,N_4388);
nand U5308 (N_5308,N_1015,N_699);
xor U5309 (N_5309,N_1147,N_2920);
xnor U5310 (N_5310,N_4735,N_1620);
xor U5311 (N_5311,N_1134,N_1937);
and U5312 (N_5312,N_2965,N_4502);
and U5313 (N_5313,N_3085,N_2577);
or U5314 (N_5314,N_503,N_188);
nor U5315 (N_5315,N_4889,N_654);
nor U5316 (N_5316,N_2475,N_4156);
and U5317 (N_5317,N_739,N_3169);
nor U5318 (N_5318,N_2448,N_3799);
or U5319 (N_5319,N_2950,N_574);
or U5320 (N_5320,N_1657,N_820);
xor U5321 (N_5321,N_1816,N_4193);
xor U5322 (N_5322,N_3953,N_3199);
and U5323 (N_5323,N_2350,N_409);
nand U5324 (N_5324,N_4891,N_769);
or U5325 (N_5325,N_4698,N_2231);
or U5326 (N_5326,N_2522,N_2829);
nand U5327 (N_5327,N_3195,N_1441);
and U5328 (N_5328,N_2474,N_2789);
or U5329 (N_5329,N_1954,N_1923);
nand U5330 (N_5330,N_861,N_294);
and U5331 (N_5331,N_4218,N_1695);
and U5332 (N_5332,N_4537,N_4169);
or U5333 (N_5333,N_4069,N_2666);
and U5334 (N_5334,N_1434,N_334);
nand U5335 (N_5335,N_812,N_52);
nor U5336 (N_5336,N_1324,N_3314);
nand U5337 (N_5337,N_283,N_1658);
and U5338 (N_5338,N_2219,N_4480);
and U5339 (N_5339,N_887,N_1951);
or U5340 (N_5340,N_2513,N_3745);
xor U5341 (N_5341,N_4443,N_495);
or U5342 (N_5342,N_3695,N_2373);
nor U5343 (N_5343,N_3786,N_533);
xnor U5344 (N_5344,N_3499,N_3610);
xnor U5345 (N_5345,N_1457,N_2053);
nor U5346 (N_5346,N_4604,N_4625);
and U5347 (N_5347,N_1014,N_3329);
nand U5348 (N_5348,N_2878,N_732);
xnor U5349 (N_5349,N_811,N_1280);
nand U5350 (N_5350,N_1282,N_914);
xnor U5351 (N_5351,N_2605,N_1366);
and U5352 (N_5352,N_3782,N_130);
nor U5353 (N_5353,N_1260,N_1802);
or U5354 (N_5354,N_411,N_4496);
xor U5355 (N_5355,N_2959,N_4684);
xor U5356 (N_5356,N_165,N_3322);
or U5357 (N_5357,N_414,N_360);
nor U5358 (N_5358,N_2036,N_254);
or U5359 (N_5359,N_2396,N_4252);
nand U5360 (N_5360,N_2800,N_4751);
xor U5361 (N_5361,N_2421,N_4993);
or U5362 (N_5362,N_4711,N_2004);
or U5363 (N_5363,N_1681,N_3582);
and U5364 (N_5364,N_4772,N_3251);
xnor U5365 (N_5365,N_4230,N_1542);
nor U5366 (N_5366,N_4227,N_4368);
nand U5367 (N_5367,N_3126,N_4187);
nor U5368 (N_5368,N_4847,N_2435);
nand U5369 (N_5369,N_3214,N_1965);
nor U5370 (N_5370,N_932,N_1472);
xor U5371 (N_5371,N_4318,N_1811);
or U5372 (N_5372,N_1384,N_4875);
or U5373 (N_5373,N_3545,N_628);
nor U5374 (N_5374,N_1189,N_2297);
nand U5375 (N_5375,N_2656,N_394);
or U5376 (N_5376,N_1518,N_2897);
xnor U5377 (N_5377,N_974,N_3537);
nor U5378 (N_5378,N_3215,N_4616);
nor U5379 (N_5379,N_3517,N_4001);
nor U5380 (N_5380,N_3492,N_373);
and U5381 (N_5381,N_1535,N_453);
nand U5382 (N_5382,N_1635,N_4672);
nor U5383 (N_5383,N_3580,N_2602);
nand U5384 (N_5384,N_997,N_1433);
and U5385 (N_5385,N_1171,N_4881);
xnor U5386 (N_5386,N_3595,N_3586);
xor U5387 (N_5387,N_937,N_1223);
nor U5388 (N_5388,N_3263,N_4064);
nand U5389 (N_5389,N_3628,N_126);
and U5390 (N_5390,N_2042,N_2241);
xnor U5391 (N_5391,N_4601,N_1388);
nand U5392 (N_5392,N_466,N_4617);
nor U5393 (N_5393,N_2107,N_821);
xor U5394 (N_5394,N_3775,N_1920);
and U5395 (N_5395,N_4093,N_1477);
and U5396 (N_5396,N_1091,N_4042);
and U5397 (N_5397,N_4488,N_2909);
nor U5398 (N_5398,N_4904,N_2621);
nor U5399 (N_5399,N_948,N_1834);
xor U5400 (N_5400,N_2980,N_3201);
and U5401 (N_5401,N_2180,N_275);
xor U5402 (N_5402,N_4264,N_3090);
nor U5403 (N_5403,N_1889,N_3935);
and U5404 (N_5404,N_566,N_4279);
and U5405 (N_5405,N_1109,N_3032);
nand U5406 (N_5406,N_3002,N_4897);
xnor U5407 (N_5407,N_3477,N_2843);
or U5408 (N_5408,N_2708,N_242);
nand U5409 (N_5409,N_4896,N_1587);
nor U5410 (N_5410,N_2258,N_2625);
nand U5411 (N_5411,N_2520,N_4829);
and U5412 (N_5412,N_3121,N_4399);
nand U5413 (N_5413,N_4830,N_4006);
xnor U5414 (N_5414,N_2845,N_4340);
or U5415 (N_5415,N_728,N_878);
nand U5416 (N_5416,N_3479,N_2628);
xnor U5417 (N_5417,N_70,N_3063);
nand U5418 (N_5418,N_3035,N_291);
or U5419 (N_5419,N_1386,N_2403);
nor U5420 (N_5420,N_3435,N_4552);
and U5421 (N_5421,N_3964,N_3171);
and U5422 (N_5422,N_428,N_1626);
and U5423 (N_5423,N_96,N_3542);
nand U5424 (N_5424,N_238,N_4285);
xor U5425 (N_5425,N_653,N_1675);
or U5426 (N_5426,N_4612,N_3061);
nand U5427 (N_5427,N_4681,N_1395);
nor U5428 (N_5428,N_2516,N_2860);
nand U5429 (N_5429,N_3287,N_898);
and U5430 (N_5430,N_1770,N_696);
and U5431 (N_5431,N_941,N_4429);
and U5432 (N_5432,N_1170,N_4969);
nand U5433 (N_5433,N_311,N_1640);
nand U5434 (N_5434,N_2949,N_4495);
xor U5435 (N_5435,N_3406,N_1155);
nand U5436 (N_5436,N_2925,N_4456);
nand U5437 (N_5437,N_4018,N_4977);
xor U5438 (N_5438,N_3965,N_4474);
nand U5439 (N_5439,N_3870,N_3177);
nor U5440 (N_5440,N_4664,N_319);
xor U5441 (N_5441,N_57,N_4742);
or U5442 (N_5442,N_2346,N_829);
and U5443 (N_5443,N_2506,N_975);
nor U5444 (N_5444,N_3728,N_1579);
nand U5445 (N_5445,N_3690,N_4532);
and U5446 (N_5446,N_787,N_2633);
xor U5447 (N_5447,N_768,N_3579);
or U5448 (N_5448,N_4391,N_4756);
nand U5449 (N_5449,N_2834,N_659);
and U5450 (N_5450,N_4009,N_4945);
or U5451 (N_5451,N_921,N_1162);
nor U5452 (N_5452,N_3466,N_2869);
xor U5453 (N_5453,N_665,N_3937);
and U5454 (N_5454,N_4026,N_30);
or U5455 (N_5455,N_2018,N_489);
nor U5456 (N_5456,N_2420,N_1719);
or U5457 (N_5457,N_1097,N_3184);
and U5458 (N_5458,N_2831,N_4079);
or U5459 (N_5459,N_3137,N_506);
nor U5460 (N_5460,N_1144,N_4249);
and U5461 (N_5461,N_2818,N_4398);
nand U5462 (N_5462,N_4186,N_444);
nand U5463 (N_5463,N_4543,N_697);
nor U5464 (N_5464,N_854,N_2113);
and U5465 (N_5465,N_4289,N_2808);
xor U5466 (N_5466,N_2284,N_4837);
and U5467 (N_5467,N_4995,N_2527);
nor U5468 (N_5468,N_3732,N_669);
and U5469 (N_5469,N_4750,N_4935);
and U5470 (N_5470,N_2574,N_1682);
nand U5471 (N_5471,N_4846,N_507);
or U5472 (N_5472,N_1341,N_3459);
nand U5473 (N_5473,N_4933,N_742);
and U5474 (N_5474,N_4797,N_4425);
nor U5475 (N_5475,N_564,N_2287);
and U5476 (N_5476,N_4724,N_2007);
nand U5477 (N_5477,N_3705,N_3067);
nand U5478 (N_5478,N_2214,N_299);
xor U5479 (N_5479,N_29,N_512);
and U5480 (N_5480,N_3557,N_2926);
nor U5481 (N_5481,N_2406,N_2409);
and U5482 (N_5482,N_1001,N_4372);
and U5483 (N_5483,N_4396,N_2732);
nand U5484 (N_5484,N_3125,N_3613);
or U5485 (N_5485,N_3122,N_4028);
and U5486 (N_5486,N_370,N_3707);
nand U5487 (N_5487,N_4825,N_3139);
nand U5488 (N_5488,N_800,N_3497);
xor U5489 (N_5489,N_3666,N_3266);
xor U5490 (N_5490,N_4581,N_2511);
nor U5491 (N_5491,N_4955,N_3878);
and U5492 (N_5492,N_3919,N_960);
nand U5493 (N_5493,N_2846,N_1263);
nand U5494 (N_5494,N_585,N_330);
and U5495 (N_5495,N_3294,N_2224);
nand U5496 (N_5496,N_3529,N_4084);
nor U5497 (N_5497,N_1039,N_88);
xnor U5498 (N_5498,N_1082,N_2207);
nand U5499 (N_5499,N_828,N_1219);
or U5500 (N_5500,N_4114,N_2627);
xor U5501 (N_5501,N_1236,N_3655);
or U5502 (N_5502,N_2539,N_2745);
and U5503 (N_5503,N_704,N_3437);
xor U5504 (N_5504,N_118,N_4584);
nor U5505 (N_5505,N_879,N_2354);
nand U5506 (N_5506,N_756,N_648);
nor U5507 (N_5507,N_3932,N_461);
nor U5508 (N_5508,N_936,N_858);
nor U5509 (N_5509,N_3076,N_876);
or U5510 (N_5510,N_2575,N_2271);
nand U5511 (N_5511,N_3942,N_3069);
or U5512 (N_5512,N_607,N_3270);
nor U5513 (N_5513,N_2132,N_20);
and U5514 (N_5514,N_255,N_1309);
nor U5515 (N_5515,N_4164,N_1737);
nor U5516 (N_5516,N_2630,N_2478);
or U5517 (N_5517,N_472,N_1936);
xnor U5518 (N_5518,N_4801,N_4671);
and U5519 (N_5519,N_1207,N_1958);
or U5520 (N_5520,N_1432,N_1202);
and U5521 (N_5521,N_3996,N_2801);
or U5522 (N_5522,N_1933,N_3576);
or U5523 (N_5523,N_2596,N_4373);
and U5524 (N_5524,N_3867,N_4401);
nor U5525 (N_5525,N_2904,N_3864);
nor U5526 (N_5526,N_4707,N_2927);
xnor U5527 (N_5527,N_3846,N_1809);
or U5528 (N_5528,N_1796,N_1602);
xor U5529 (N_5529,N_3806,N_3658);
nor U5530 (N_5530,N_3872,N_4212);
and U5531 (N_5531,N_32,N_2104);
or U5532 (N_5532,N_939,N_2710);
or U5533 (N_5533,N_617,N_3325);
nor U5534 (N_5534,N_4646,N_2844);
nand U5535 (N_5535,N_4002,N_3472);
or U5536 (N_5536,N_2617,N_522);
or U5537 (N_5537,N_2072,N_1637);
nand U5538 (N_5538,N_4298,N_1720);
nand U5539 (N_5539,N_2118,N_1328);
or U5540 (N_5540,N_1124,N_3131);
and U5541 (N_5541,N_3368,N_3618);
and U5542 (N_5542,N_1381,N_1927);
and U5543 (N_5543,N_4795,N_2531);
xnor U5544 (N_5544,N_2122,N_526);
nor U5545 (N_5545,N_344,N_989);
nor U5546 (N_5546,N_3013,N_872);
and U5547 (N_5547,N_2901,N_616);
nor U5548 (N_5548,N_3857,N_4177);
or U5549 (N_5549,N_3181,N_2447);
and U5550 (N_5550,N_1669,N_1100);
xnor U5551 (N_5551,N_2172,N_2415);
or U5552 (N_5552,N_120,N_3809);
nor U5553 (N_5553,N_1303,N_1254);
nor U5554 (N_5554,N_1043,N_4549);
xor U5555 (N_5555,N_263,N_4085);
or U5556 (N_5556,N_1511,N_107);
or U5557 (N_5557,N_4255,N_2886);
nand U5558 (N_5558,N_2972,N_2786);
or U5559 (N_5559,N_4406,N_1596);
nand U5560 (N_5560,N_4832,N_280);
nand U5561 (N_5561,N_3550,N_2394);
nor U5562 (N_5562,N_1532,N_2145);
and U5563 (N_5563,N_563,N_3249);
nor U5564 (N_5564,N_3716,N_3981);
nand U5565 (N_5565,N_2955,N_3604);
nor U5566 (N_5566,N_3673,N_2963);
xnor U5567 (N_5567,N_4173,N_916);
or U5568 (N_5568,N_220,N_1313);
or U5569 (N_5569,N_3231,N_4840);
nand U5570 (N_5570,N_2318,N_1387);
or U5571 (N_5571,N_4434,N_4263);
nand U5572 (N_5572,N_943,N_2467);
and U5573 (N_5573,N_2248,N_205);
nand U5574 (N_5574,N_2940,N_3918);
xnor U5575 (N_5575,N_4515,N_171);
or U5576 (N_5576,N_4148,N_2876);
and U5577 (N_5577,N_4426,N_3114);
nand U5578 (N_5578,N_4126,N_1031);
nor U5579 (N_5579,N_3742,N_4539);
nand U5580 (N_5580,N_4863,N_405);
or U5581 (N_5581,N_2524,N_4652);
nand U5582 (N_5582,N_3717,N_3719);
nand U5583 (N_5583,N_3417,N_4892);
xor U5584 (N_5584,N_2649,N_3611);
xnor U5585 (N_5585,N_4134,N_1611);
and U5586 (N_5586,N_4634,N_1698);
nand U5587 (N_5587,N_2594,N_4228);
nor U5588 (N_5588,N_1815,N_4143);
xnor U5589 (N_5589,N_2005,N_976);
or U5590 (N_5590,N_257,N_1201);
nor U5591 (N_5591,N_2523,N_502);
or U5592 (N_5592,N_406,N_3042);
and U5593 (N_5593,N_3053,N_4096);
and U5594 (N_5594,N_3764,N_2158);
and U5595 (N_5595,N_2854,N_1333);
and U5596 (N_5596,N_2099,N_1685);
nor U5597 (N_5597,N_3513,N_315);
xor U5598 (N_5598,N_4136,N_4133);
xor U5599 (N_5599,N_3015,N_2059);
or U5600 (N_5600,N_2279,N_4708);
nor U5601 (N_5601,N_2995,N_3718);
and U5602 (N_5602,N_3004,N_4974);
nor U5603 (N_5603,N_3978,N_2212);
and U5604 (N_5604,N_4999,N_4137);
and U5605 (N_5605,N_1619,N_4432);
or U5606 (N_5606,N_2499,N_3522);
nor U5607 (N_5607,N_480,N_4141);
xor U5608 (N_5608,N_3113,N_3889);
and U5609 (N_5609,N_1420,N_928);
nor U5610 (N_5610,N_4507,N_1756);
or U5611 (N_5611,N_3262,N_1464);
and U5612 (N_5612,N_1168,N_4741);
and U5613 (N_5613,N_3921,N_457);
and U5614 (N_5614,N_2117,N_4211);
nor U5615 (N_5615,N_267,N_452);
and U5616 (N_5616,N_4519,N_709);
and U5617 (N_5617,N_3982,N_4512);
and U5618 (N_5618,N_2559,N_1707);
nor U5619 (N_5619,N_3614,N_1588);
nand U5620 (N_5620,N_4917,N_2957);
and U5621 (N_5621,N_4030,N_1174);
xnor U5622 (N_5622,N_3074,N_4221);
xnor U5623 (N_5623,N_2123,N_3558);
xnor U5624 (N_5624,N_1293,N_2755);
or U5625 (N_5625,N_3571,N_2919);
and U5626 (N_5626,N_4242,N_1232);
nand U5627 (N_5627,N_923,N_2662);
or U5628 (N_5628,N_2882,N_1972);
nor U5629 (N_5629,N_4870,N_4589);
or U5630 (N_5630,N_3698,N_1835);
or U5631 (N_5631,N_3855,N_3939);
xnor U5632 (N_5632,N_927,N_3772);
nor U5633 (N_5633,N_22,N_1479);
nor U5634 (N_5634,N_2344,N_2733);
nand U5635 (N_5635,N_2937,N_4692);
and U5636 (N_5636,N_856,N_1154);
or U5637 (N_5637,N_2407,N_3738);
xnor U5638 (N_5638,N_837,N_3994);
xnor U5639 (N_5639,N_3931,N_4544);
nand U5640 (N_5640,N_4588,N_1148);
or U5641 (N_5641,N_4998,N_2242);
nor U5642 (N_5642,N_2544,N_1383);
and U5643 (N_5643,N_1649,N_3756);
xor U5644 (N_5644,N_2564,N_4670);
or U5645 (N_5645,N_3257,N_1139);
and U5646 (N_5646,N_4822,N_1012);
nor U5647 (N_5647,N_2765,N_3009);
nand U5648 (N_5648,N_1565,N_3744);
xnor U5649 (N_5649,N_900,N_2183);
nor U5650 (N_5650,N_1463,N_3880);
or U5651 (N_5651,N_1772,N_646);
nor U5652 (N_5652,N_4697,N_3358);
or U5653 (N_5653,N_1798,N_1491);
xnor U5654 (N_5654,N_2996,N_3438);
xor U5655 (N_5655,N_4044,N_3432);
or U5656 (N_5656,N_3674,N_4115);
or U5657 (N_5657,N_934,N_2092);
xor U5658 (N_5658,N_4288,N_3383);
nor U5659 (N_5659,N_4445,N_4685);
and U5660 (N_5660,N_813,N_363);
nand U5661 (N_5661,N_1348,N_783);
nand U5662 (N_5662,N_4147,N_2640);
and U5663 (N_5663,N_2748,N_818);
xor U5664 (N_5664,N_2715,N_102);
and U5665 (N_5665,N_3549,N_3887);
nor U5666 (N_5666,N_3157,N_4359);
and U5667 (N_5667,N_2794,N_384);
nand U5668 (N_5668,N_3958,N_4492);
and U5669 (N_5669,N_4571,N_4594);
xnor U5670 (N_5670,N_4419,N_1128);
or U5671 (N_5671,N_359,N_4236);
xnor U5672 (N_5672,N_598,N_4408);
nor U5673 (N_5673,N_2352,N_2855);
nand U5674 (N_5674,N_3408,N_1355);
nand U5675 (N_5675,N_81,N_2714);
nor U5676 (N_5676,N_4290,N_2606);
nor U5677 (N_5677,N_1624,N_1514);
xnor U5678 (N_5678,N_3108,N_1374);
or U5679 (N_5679,N_3178,N_1830);
nor U5680 (N_5680,N_2857,N_4879);
nand U5681 (N_5681,N_1138,N_4834);
nand U5682 (N_5682,N_1647,N_1502);
and U5683 (N_5683,N_1975,N_1702);
xnor U5684 (N_5684,N_403,N_4587);
or U5685 (N_5685,N_1704,N_4162);
nand U5686 (N_5686,N_4653,N_3486);
nor U5687 (N_5687,N_3840,N_501);
and U5688 (N_5688,N_755,N_521);
or U5689 (N_5689,N_1831,N_3309);
nor U5690 (N_5690,N_2223,N_3765);
nor U5691 (N_5691,N_520,N_840);
nand U5692 (N_5692,N_1510,N_2824);
and U5693 (N_5693,N_2147,N_1020);
or U5694 (N_5694,N_3268,N_2339);
nand U5695 (N_5695,N_3633,N_4145);
nor U5696 (N_5696,N_2402,N_621);
nor U5697 (N_5697,N_1690,N_671);
and U5698 (N_5698,N_1307,N_3436);
nor U5699 (N_5699,N_2781,N_2061);
xnor U5700 (N_5700,N_683,N_4273);
xnor U5701 (N_5701,N_2970,N_2027);
or U5702 (N_5702,N_4991,N_14);
or U5703 (N_5703,N_447,N_3278);
and U5704 (N_5704,N_1665,N_312);
xnor U5705 (N_5705,N_3474,N_1964);
or U5706 (N_5706,N_765,N_178);
nor U5707 (N_5707,N_1941,N_3621);
xor U5708 (N_5708,N_2740,N_2973);
xor U5709 (N_5709,N_1022,N_3338);
nor U5710 (N_5710,N_2851,N_1237);
nor U5711 (N_5711,N_5,N_4932);
and U5712 (N_5712,N_3810,N_3834);
xor U5713 (N_5713,N_2968,N_1549);
nand U5714 (N_5714,N_3145,N_1848);
nand U5715 (N_5715,N_1000,N_3814);
or U5716 (N_5716,N_3029,N_2362);
and U5717 (N_5717,N_543,N_2020);
and U5718 (N_5718,N_4709,N_4908);
nor U5719 (N_5719,N_13,N_4302);
and U5720 (N_5720,N_2136,N_3483);
or U5721 (N_5721,N_4768,N_3078);
nor U5722 (N_5722,N_634,N_4206);
or U5723 (N_5723,N_736,N_2651);
or U5724 (N_5724,N_2895,N_3244);
nor U5725 (N_5725,N_4844,N_2000);
nand U5726 (N_5726,N_3261,N_7);
xor U5727 (N_5727,N_4560,N_3976);
and U5728 (N_5728,N_3112,N_1349);
xnor U5729 (N_5729,N_4104,N_1849);
xor U5730 (N_5730,N_2049,N_3975);
nor U5731 (N_5731,N_2274,N_4016);
or U5732 (N_5732,N_1452,N_2525);
nand U5733 (N_5733,N_3636,N_4850);
xnor U5734 (N_5734,N_1215,N_883);
and U5735 (N_5735,N_4240,N_2465);
and U5736 (N_5736,N_4824,N_1026);
nand U5737 (N_5737,N_3670,N_1278);
nand U5738 (N_5738,N_4110,N_3304);
xnor U5739 (N_5739,N_4219,N_2547);
and U5740 (N_5740,N_1893,N_1498);
and U5741 (N_5741,N_4954,N_4710);
or U5742 (N_5742,N_2812,N_2615);
xnor U5743 (N_5743,N_1912,N_1621);
or U5744 (N_5744,N_2758,N_3335);
or U5745 (N_5745,N_1013,N_2039);
nor U5746 (N_5746,N_4317,N_2678);
or U5747 (N_5747,N_4836,N_933);
nand U5748 (N_5748,N_1112,N_4925);
and U5749 (N_5749,N_3008,N_3056);
xnor U5750 (N_5750,N_1536,N_4354);
nor U5751 (N_5751,N_953,N_3647);
nor U5752 (N_5752,N_4758,N_1528);
nand U5753 (N_5753,N_1723,N_4668);
xor U5754 (N_5754,N_440,N_1468);
nor U5755 (N_5755,N_2303,N_781);
and U5756 (N_5756,N_2466,N_2905);
nor U5757 (N_5757,N_84,N_3445);
and U5758 (N_5758,N_4522,N_802);
nand U5759 (N_5759,N_2095,N_2683);
or U5760 (N_5760,N_4624,N_4620);
xor U5761 (N_5761,N_2268,N_2111);
nor U5762 (N_5762,N_631,N_364);
nand U5763 (N_5763,N_3531,N_4739);
nand U5764 (N_5764,N_4953,N_67);
and U5765 (N_5765,N_4000,N_2747);
nand U5766 (N_5766,N_4204,N_1242);
or U5767 (N_5767,N_3569,N_3470);
nor U5768 (N_5768,N_4586,N_381);
and U5769 (N_5769,N_1870,N_1639);
and U5770 (N_5770,N_2723,N_737);
xnor U5771 (N_5771,N_2647,N_1864);
and U5772 (N_5772,N_2253,N_4184);
and U5773 (N_5773,N_1141,N_39);
nand U5774 (N_5774,N_1460,N_427);
xnor U5775 (N_5775,N_3720,N_1915);
and U5776 (N_5776,N_1728,N_4365);
and U5777 (N_5777,N_4902,N_1668);
xor U5778 (N_5778,N_3333,N_185);
nand U5779 (N_5779,N_3797,N_2704);
nand U5780 (N_5780,N_3565,N_303);
or U5781 (N_5781,N_4449,N_1607);
or U5782 (N_5782,N_1480,N_92);
or U5783 (N_5783,N_2335,N_3339);
nor U5784 (N_5784,N_793,N_3381);
nor U5785 (N_5785,N_3372,N_727);
or U5786 (N_5786,N_4551,N_3073);
or U5787 (N_5787,N_3149,N_1266);
or U5788 (N_5788,N_2533,N_2164);
and U5789 (N_5789,N_2228,N_4816);
nand U5790 (N_5790,N_2832,N_3632);
nand U5791 (N_5791,N_2267,N_1745);
nor U5792 (N_5792,N_10,N_949);
nor U5793 (N_5793,N_2294,N_3938);
nand U5794 (N_5794,N_3763,N_4570);
nor U5795 (N_5795,N_1652,N_2306);
or U5796 (N_5796,N_3027,N_4216);
or U5797 (N_5797,N_3203,N_2311);
xnor U5798 (N_5798,N_207,N_2703);
nor U5799 (N_5799,N_3693,N_1765);
nor U5800 (N_5800,N_2839,N_2696);
or U5801 (N_5801,N_3784,N_4796);
nand U5802 (N_5802,N_241,N_1042);
xnor U5803 (N_5803,N_1513,N_1418);
or U5804 (N_5804,N_4686,N_547);
or U5805 (N_5805,N_3955,N_4311);
and U5806 (N_5806,N_4538,N_4066);
and U5807 (N_5807,N_700,N_4383);
xnor U5808 (N_5808,N_2767,N_4004);
or U5809 (N_5809,N_456,N_645);
or U5810 (N_5810,N_4461,N_2450);
xor U5811 (N_5811,N_4217,N_2216);
nand U5812 (N_5812,N_2184,N_4316);
and U5813 (N_5813,N_3777,N_3402);
and U5814 (N_5814,N_328,N_3482);
and U5815 (N_5815,N_1051,N_122);
and U5816 (N_5816,N_694,N_3503);
and U5817 (N_5817,N_1557,N_467);
xnor U5818 (N_5818,N_154,N_524);
and U5819 (N_5819,N_3105,N_1192);
and U5820 (N_5820,N_1361,N_4949);
xnor U5821 (N_5821,N_3552,N_917);
or U5822 (N_5822,N_94,N_1982);
and U5823 (N_5823,N_3635,N_4334);
or U5824 (N_5824,N_2936,N_2653);
nand U5825 (N_5825,N_4673,N_3680);
xnor U5826 (N_5826,N_3733,N_89);
nor U5827 (N_5827,N_1823,N_1820);
xor U5828 (N_5828,N_4894,N_4460);
nor U5829 (N_5829,N_1029,N_912);
xor U5830 (N_5830,N_780,N_2193);
and U5831 (N_5831,N_3825,N_498);
and U5832 (N_5832,N_1443,N_3699);
and U5833 (N_5833,N_308,N_791);
or U5834 (N_5834,N_2296,N_2623);
and U5835 (N_5835,N_3801,N_1107);
nand U5836 (N_5836,N_4308,N_560);
nor U5837 (N_5837,N_3299,N_42);
nor U5838 (N_5838,N_2322,N_4257);
or U5839 (N_5839,N_2130,N_4800);
and U5840 (N_5840,N_4845,N_4674);
and U5841 (N_5841,N_4404,N_3852);
xor U5842 (N_5842,N_761,N_2810);
or U5843 (N_5843,N_1322,N_4909);
nand U5844 (N_5844,N_4139,N_2585);
and U5845 (N_5845,N_906,N_3607);
xnor U5846 (N_5846,N_1130,N_3907);
and U5847 (N_5847,N_2680,N_4247);
and U5848 (N_5848,N_4701,N_58);
and U5849 (N_5849,N_1732,N_3123);
xor U5850 (N_5850,N_4335,N_4960);
and U5851 (N_5851,N_4410,N_2454);
nand U5852 (N_5852,N_1072,N_925);
xor U5853 (N_5853,N_2378,N_259);
or U5854 (N_5854,N_2751,N_3533);
nor U5855 (N_5855,N_1190,N_1019);
nand U5856 (N_5856,N_1221,N_3327);
xor U5857 (N_5857,N_2676,N_268);
nor U5858 (N_5858,N_1288,N_4438);
or U5859 (N_5859,N_3617,N_262);
nor U5860 (N_5860,N_2260,N_4327);
xor U5861 (N_5861,N_108,N_1380);
nor U5862 (N_5862,N_3148,N_3285);
xor U5863 (N_5863,N_1773,N_347);
xor U5864 (N_5864,N_4579,N_54);
or U5865 (N_5865,N_305,N_324);
or U5866 (N_5866,N_4132,N_1119);
xnor U5867 (N_5867,N_1486,N_3310);
nor U5868 (N_5868,N_1774,N_2958);
or U5869 (N_5869,N_956,N_1726);
or U5870 (N_5870,N_2264,N_2866);
nor U5871 (N_5871,N_2534,N_3581);
or U5872 (N_5872,N_73,N_1391);
and U5873 (N_5873,N_2570,N_4057);
nand U5874 (N_5874,N_2718,N_4301);
or U5875 (N_5875,N_2110,N_4248);
xnor U5876 (N_5876,N_4241,N_2932);
and U5877 (N_5877,N_2616,N_4303);
nor U5878 (N_5878,N_4883,N_3897);
nor U5879 (N_5879,N_772,N_3208);
nor U5880 (N_5880,N_233,N_4803);
or U5881 (N_5881,N_2011,N_2280);
nor U5882 (N_5882,N_2752,N_4339);
xor U5883 (N_5883,N_2569,N_4659);
xor U5884 (N_5884,N_2051,N_2582);
nand U5885 (N_5885,N_189,N_1791);
nor U5886 (N_5886,N_3813,N_3080);
xnor U5887 (N_5887,N_4367,N_3132);
nand U5888 (N_5888,N_966,N_2169);
nor U5889 (N_5889,N_3211,N_4213);
or U5890 (N_5890,N_3065,N_4725);
nor U5891 (N_5891,N_4469,N_3187);
or U5892 (N_5892,N_1466,N_1084);
nand U5893 (N_5893,N_1959,N_2455);
nand U5894 (N_5894,N_3822,N_1241);
or U5895 (N_5895,N_3908,N_1195);
xnor U5896 (N_5896,N_2395,N_1449);
nand U5897 (N_5897,N_4479,N_823);
xnor U5898 (N_5898,N_1605,N_3191);
or U5899 (N_5899,N_632,N_4347);
or U5900 (N_5900,N_582,N_2383);
nand U5901 (N_5901,N_676,N_2655);
and U5902 (N_5902,N_174,N_2650);
and U5903 (N_5903,N_1999,N_3749);
xnor U5904 (N_5904,N_2298,N_3311);
and U5905 (N_5905,N_588,N_2637);
nand U5906 (N_5906,N_1546,N_2048);
xor U5907 (N_5907,N_4157,N_3861);
xnor U5908 (N_5908,N_3183,N_1411);
nand U5909 (N_5909,N_1185,N_286);
nand U5910 (N_5910,N_1856,N_3081);
xnor U5911 (N_5911,N_4516,N_4814);
nor U5912 (N_5912,N_2485,N_2847);
or U5913 (N_5913,N_4074,N_3596);
or U5914 (N_5914,N_4988,N_3672);
or U5915 (N_5915,N_2060,N_4489);
xnor U5916 (N_5916,N_771,N_3237);
xor U5917 (N_5917,N_1493,N_1751);
or U5918 (N_5918,N_4411,N_3127);
xor U5919 (N_5919,N_4214,N_2734);
or U5920 (N_5920,N_1524,N_3600);
and U5921 (N_5921,N_1132,N_2046);
or U5922 (N_5922,N_987,N_4326);
and U5923 (N_5923,N_4700,N_3259);
nand U5924 (N_5924,N_4270,N_206);
and U5925 (N_5925,N_3315,N_3274);
nand U5926 (N_5926,N_3275,N_1009);
nor U5927 (N_5927,N_1679,N_3233);
or U5928 (N_5928,N_4818,N_1929);
and U5929 (N_5929,N_33,N_3691);
and U5930 (N_5930,N_4849,N_4220);
or U5931 (N_5931,N_4535,N_2902);
nand U5932 (N_5932,N_4567,N_1344);
nand U5933 (N_5933,N_3467,N_782);
xor U5934 (N_5934,N_1220,N_4971);
nor U5935 (N_5935,N_3429,N_4992);
and U5936 (N_5936,N_2244,N_1310);
or U5937 (N_5937,N_3225,N_1793);
nor U5938 (N_5938,N_3446,N_603);
nand U5939 (N_5939,N_4014,N_3998);
nor U5940 (N_5940,N_3662,N_3129);
nand U5941 (N_5941,N_1209,N_3473);
nor U5942 (N_5942,N_3265,N_3284);
nand U5943 (N_5943,N_3794,N_2816);
or U5944 (N_5944,N_354,N_4526);
or U5945 (N_5945,N_2178,N_2075);
nand U5946 (N_5946,N_3683,N_611);
or U5947 (N_5947,N_1382,N_4611);
xnor U5948 (N_5948,N_4819,N_2660);
or U5949 (N_5949,N_470,N_981);
nand U5950 (N_5950,N_1272,N_4591);
nand U5951 (N_5951,N_3453,N_4871);
or U5952 (N_5952,N_4728,N_3750);
and U5953 (N_5953,N_4047,N_1861);
or U5954 (N_5954,N_1450,N_2593);
xor U5955 (N_5955,N_2144,N_1077);
nand U5956 (N_5956,N_4201,N_3612);
and U5957 (N_5957,N_904,N_891);
and U5958 (N_5958,N_2230,N_3228);
or U5959 (N_5959,N_3109,N_1083);
or U5960 (N_5960,N_1504,N_1123);
and U5961 (N_5961,N_3817,N_204);
nor U5962 (N_5962,N_1055,N_3342);
nor U5963 (N_5963,N_4258,N_626);
nand U5964 (N_5964,N_4130,N_4996);
nand U5965 (N_5965,N_4433,N_972);
or U5966 (N_5966,N_1459,N_2309);
nand U5967 (N_5967,N_951,N_4790);
xnor U5968 (N_5968,N_463,N_1539);
nor U5969 (N_5969,N_1389,N_69);
xor U5970 (N_5970,N_1922,N_4786);
and U5971 (N_5971,N_3360,N_1085);
nand U5972 (N_5972,N_2040,N_2541);
nand U5973 (N_5973,N_1412,N_745);
nand U5974 (N_5974,N_2540,N_857);
xnor U5975 (N_5975,N_2554,N_4199);
or U5976 (N_5976,N_4680,N_157);
and U5977 (N_5977,N_2567,N_2401);
xor U5978 (N_5978,N_4713,N_1230);
and U5979 (N_5979,N_4876,N_4730);
xnor U5980 (N_5980,N_2150,N_306);
xnor U5981 (N_5981,N_4636,N_4658);
and U5982 (N_5982,N_1393,N_59);
nand U5983 (N_5983,N_1733,N_2128);
or U5984 (N_5984,N_3877,N_2624);
or U5985 (N_5985,N_846,N_2681);
or U5986 (N_5986,N_2483,N_418);
xor U5987 (N_5987,N_2037,N_1191);
nand U5988 (N_5988,N_1661,N_902);
or U5989 (N_5989,N_1304,N_2129);
nor U5990 (N_5990,N_3648,N_404);
or U5991 (N_5991,N_1655,N_3627);
xor U5992 (N_5992,N_2983,N_2503);
nor U5993 (N_5993,N_1832,N_3252);
xor U5994 (N_5994,N_1771,N_833);
or U5995 (N_5995,N_1899,N_2473);
or U5996 (N_5996,N_1305,N_150);
or U5997 (N_5997,N_97,N_3973);
xor U5998 (N_5998,N_2225,N_2168);
nor U5999 (N_5999,N_565,N_516);
nand U6000 (N_6000,N_3449,N_2305);
xor U6001 (N_6001,N_3377,N_3373);
xnor U6002 (N_6002,N_4422,N_983);
xor U6003 (N_6003,N_3901,N_1520);
nand U6004 (N_6004,N_3343,N_2792);
nand U6005 (N_6005,N_3760,N_4603);
nor U6006 (N_6006,N_1523,N_1239);
or U6007 (N_6007,N_1739,N_4643);
nor U6008 (N_6008,N_1198,N_1136);
xor U6009 (N_6009,N_571,N_4155);
or U6010 (N_6010,N_244,N_4352);
and U6011 (N_6011,N_729,N_3419);
nand U6012 (N_6012,N_3095,N_197);
or U6013 (N_6013,N_3723,N_2620);
nand U6014 (N_6014,N_2433,N_1526);
or U6015 (N_6015,N_2156,N_385);
or U6016 (N_6016,N_4888,N_3591);
and U6017 (N_6017,N_4970,N_3051);
xor U6018 (N_6018,N_4117,N_3267);
and U6019 (N_6019,N_2667,N_1799);
or U6020 (N_6020,N_2756,N_532);
and U6021 (N_6021,N_1376,N_3321);
or U6022 (N_6022,N_4906,N_2966);
or U6023 (N_6023,N_2780,N_2835);
nor U6024 (N_6024,N_909,N_1093);
nor U6025 (N_6025,N_445,N_3677);
nand U6026 (N_6026,N_1447,N_4752);
nand U6027 (N_6027,N_2282,N_4129);
nor U6028 (N_6028,N_586,N_1746);
or U6029 (N_6029,N_1364,N_3594);
or U6030 (N_6030,N_1054,N_2052);
nor U6031 (N_6031,N_3033,N_3977);
xnor U6032 (N_6032,N_2914,N_627);
nand U6033 (N_6033,N_3896,N_4644);
or U6034 (N_6034,N_4984,N_3783);
and U6035 (N_6035,N_2389,N_1717);
or U6036 (N_6036,N_2887,N_3091);
nor U6037 (N_6037,N_1268,N_589);
and U6038 (N_6038,N_4344,N_4161);
nor U6039 (N_6039,N_529,N_2636);
nor U6040 (N_6040,N_2934,N_1371);
xnor U6041 (N_6041,N_775,N_637);
xnor U6042 (N_6042,N_4491,N_3224);
or U6043 (N_6043,N_2009,N_1867);
or U6044 (N_6044,N_944,N_3158);
or U6045 (N_6045,N_957,N_2423);
nor U6046 (N_6046,N_3099,N_3434);
or U6047 (N_6047,N_3902,N_2986);
nand U6048 (N_6048,N_538,N_3967);
and U6049 (N_6049,N_3172,N_4976);
or U6050 (N_6050,N_1475,N_111);
nand U6051 (N_6051,N_4231,N_2291);
xor U6052 (N_6052,N_4929,N_2494);
nor U6053 (N_6053,N_3374,N_4223);
or U6054 (N_6054,N_1869,N_735);
nand U6055 (N_6055,N_4921,N_1408);
and U6056 (N_6056,N_228,N_1627);
nor U6057 (N_6057,N_3630,N_986);
or U6058 (N_6058,N_4802,N_1439);
xnor U6059 (N_6059,N_1916,N_548);
nor U6060 (N_6060,N_971,N_1609);
or U6061 (N_6061,N_3072,N_2641);
and U6062 (N_6062,N_656,N_4542);
nand U6063 (N_6063,N_2238,N_179);
nor U6064 (N_6064,N_622,N_1977);
nor U6065 (N_6065,N_1990,N_261);
nand U6066 (N_6066,N_553,N_3226);
or U6067 (N_6067,N_4077,N_2247);
xnor U6068 (N_6068,N_3681,N_2917);
nand U6069 (N_6069,N_3307,N_4556);
xnor U6070 (N_6070,N_309,N_903);
nor U6071 (N_6071,N_31,N_4931);
xnor U6072 (N_6072,N_1897,N_2951);
nand U6073 (N_6073,N_4309,N_1111);
xor U6074 (N_6074,N_2239,N_1421);
xor U6075 (N_6075,N_3572,N_578);
nand U6076 (N_6076,N_2870,N_442);
nand U6077 (N_6077,N_1818,N_1503);
and U6078 (N_6078,N_2579,N_1653);
and U6079 (N_6079,N_3601,N_1845);
nor U6080 (N_6080,N_1501,N_2016);
nor U6081 (N_6081,N_2019,N_1594);
nand U6082 (N_6082,N_2235,N_1904);
nand U6083 (N_6083,N_3375,N_4324);
or U6084 (N_6084,N_3629,N_4031);
nor U6085 (N_6085,N_1678,N_4565);
xor U6086 (N_6086,N_3330,N_4142);
xnor U6087 (N_6087,N_4286,N_2899);
xor U6088 (N_6088,N_3924,N_1932);
or U6089 (N_6089,N_301,N_4261);
xnor U6090 (N_6090,N_4727,N_1249);
xnor U6091 (N_6091,N_705,N_3858);
and U6092 (N_6092,N_76,N_4052);
xnor U6093 (N_6093,N_3646,N_3506);
nand U6094 (N_6094,N_2510,N_4901);
and U6095 (N_6095,N_2969,N_3240);
xor U6096 (N_6096,N_2889,N_1325);
nor U6097 (N_6097,N_2054,N_74);
nand U6098 (N_6098,N_1711,N_376);
nor U6099 (N_6099,N_1987,N_1676);
nand U6100 (N_6100,N_1338,N_1010);
or U6101 (N_6101,N_4689,N_3578);
or U6102 (N_6102,N_744,N_3993);
or U6103 (N_6103,N_3207,N_1409);
nand U6104 (N_6104,N_3463,N_2090);
xnor U6105 (N_6105,N_106,N_1876);
nand U6106 (N_6106,N_4506,N_2739);
nand U6107 (N_6107,N_1197,N_71);
nand U6108 (N_6108,N_2325,N_1558);
xor U6109 (N_6109,N_3401,N_2003);
xor U6110 (N_6110,N_194,N_3276);
nor U6111 (N_6111,N_1571,N_955);
nand U6112 (N_6112,N_1956,N_2690);
nand U6113 (N_6113,N_4886,N_2300);
nor U6114 (N_6114,N_24,N_3890);
or U6115 (N_6115,N_2974,N_4738);
xnor U6116 (N_6116,N_1027,N_4596);
nor U6117 (N_6117,N_867,N_2551);
xnor U6118 (N_6118,N_3416,N_214);
nand U6119 (N_6119,N_773,N_4116);
and U6120 (N_6120,N_1613,N_1142);
nand U6121 (N_6121,N_68,N_2412);
nand U6122 (N_6122,N_2631,N_465);
or U6123 (N_6123,N_4677,N_4500);
xnor U6124 (N_6124,N_1429,N_2773);
and U6125 (N_6125,N_753,N_4061);
xor U6126 (N_6126,N_901,N_186);
nand U6127 (N_6127,N_3366,N_26);
nor U6128 (N_6128,N_367,N_4283);
and U6129 (N_6129,N_1080,N_1454);
xnor U6130 (N_6130,N_1281,N_2788);
nor U6131 (N_6131,N_4699,N_3098);
or U6132 (N_6132,N_1616,N_2151);
nand U6133 (N_6133,N_661,N_4321);
and U6134 (N_6134,N_227,N_3962);
nor U6135 (N_6135,N_2480,N_600);
nor U6136 (N_6136,N_4073,N_4458);
nor U6137 (N_6137,N_1953,N_3710);
nand U6138 (N_6138,N_85,N_1078);
or U6139 (N_6139,N_1730,N_4600);
nor U6140 (N_6140,N_2252,N_629);
xor U6141 (N_6141,N_2174,N_3553);
xor U6142 (N_6142,N_544,N_866);
nor U6143 (N_6143,N_4755,N_2203);
nand U6144 (N_6144,N_3671,N_4451);
xnor U6145 (N_6145,N_911,N_127);
or U6146 (N_6146,N_2805,N_433);
or U6147 (N_6147,N_4168,N_865);
and U6148 (N_6148,N_2929,N_1788);
nor U6149 (N_6149,N_4146,N_375);
xnor U6150 (N_6150,N_3771,N_4990);
nand U6151 (N_6151,N_1551,N_3868);
nor U6152 (N_6152,N_3212,N_4012);
and U6153 (N_6153,N_1419,N_1574);
or U6154 (N_6154,N_3668,N_722);
nand U6155 (N_6155,N_1891,N_1659);
nand U6156 (N_6156,N_3026,N_355);
or U6157 (N_6157,N_505,N_4208);
xnor U6158 (N_6158,N_644,N_2100);
xor U6159 (N_6159,N_3344,N_3970);
nor U6160 (N_6160,N_4128,N_959);
or U6161 (N_6161,N_4764,N_682);
or U6162 (N_6162,N_4784,N_4154);
nor U6163 (N_6163,N_3471,N_2024);
nand U6164 (N_6164,N_1759,N_569);
nand U6165 (N_6165,N_3521,N_4841);
nand U6166 (N_6166,N_1385,N_2836);
nor U6167 (N_6167,N_3317,N_1317);
and U6168 (N_6168,N_4504,N_1474);
and U6169 (N_6169,N_1400,N_101);
xor U6170 (N_6170,N_859,N_4782);
nand U6171 (N_6171,N_1979,N_87);
nor U6172 (N_6172,N_417,N_146);
or U6173 (N_6173,N_2259,N_3481);
or U6174 (N_6174,N_4903,N_2177);
or U6175 (N_6175,N_421,N_2548);
nor U6176 (N_6176,N_4762,N_1554);
and U6177 (N_6177,N_1919,N_216);
and U6178 (N_6178,N_4936,N_162);
nor U6179 (N_6179,N_1095,N_3071);
and U6180 (N_6180,N_121,N_555);
and U6181 (N_6181,N_2334,N_415);
nand U6182 (N_6182,N_3527,N_1228);
or U6183 (N_6183,N_2853,N_945);
and U6184 (N_6184,N_4209,N_2908);
nor U6185 (N_6185,N_1045,N_273);
nand U6186 (N_6186,N_1323,N_3336);
and U6187 (N_6187,N_1032,N_18);
nand U6188 (N_6188,N_3979,N_2990);
nand U6189 (N_6189,N_4972,N_2093);
nand U6190 (N_6190,N_2591,N_4127);
xor U6191 (N_6191,N_2827,N_2782);
xor U6192 (N_6192,N_2944,N_1632);
xor U6193 (N_6193,N_4939,N_4527);
xor U6194 (N_6194,N_652,N_3679);
nor U6195 (N_6195,N_2504,N_4281);
nor U6196 (N_6196,N_3535,N_139);
or U6197 (N_6197,N_3264,N_3985);
nor U6198 (N_6198,N_3762,N_1073);
or U6199 (N_6199,N_1297,N_3585);
xnor U6200 (N_6200,N_1453,N_3928);
xnor U6201 (N_6201,N_1775,N_219);
nor U6202 (N_6202,N_1852,N_3227);
and U6203 (N_6203,N_3866,N_2783);
and U6204 (N_6204,N_4827,N_613);
nand U6205 (N_6205,N_1321,N_64);
or U6206 (N_6206,N_2376,N_3869);
or U6207 (N_6207,N_2405,N_3196);
nor U6208 (N_6208,N_3185,N_3643);
nor U6209 (N_6209,N_4416,N_4029);
xnor U6210 (N_6210,N_605,N_3768);
or U6211 (N_6211,N_1069,N_4867);
xnor U6212 (N_6212,N_3875,N_4384);
nor U6213 (N_6213,N_2091,N_3844);
nor U6214 (N_6214,N_3220,N_4430);
nor U6215 (N_6215,N_3945,N_4159);
xor U6216 (N_6216,N_252,N_3018);
nor U6217 (N_6217,N_2675,N_2833);
nand U6218 (N_6218,N_4106,N_3403);
nand U6219 (N_6219,N_2488,N_4098);
or U6220 (N_6220,N_4356,N_2717);
and U6221 (N_6221,N_504,N_4158);
or U6222 (N_6222,N_4412,N_491);
nor U6223 (N_6223,N_339,N_4779);
or U6224 (N_6224,N_594,N_4864);
xor U6225 (N_6225,N_4205,N_763);
nor U6226 (N_6226,N_1909,N_1345);
or U6227 (N_6227,N_2418,N_4312);
nand U6228 (N_6228,N_436,N_731);
and U6229 (N_6229,N_1938,N_3411);
or U6230 (N_6230,N_1928,N_235);
or U6231 (N_6231,N_1888,N_2819);
or U6232 (N_6232,N_743,N_3863);
and U6233 (N_6233,N_2286,N_776);
and U6234 (N_6234,N_4962,N_4690);
nor U6235 (N_6235,N_3736,N_1986);
or U6236 (N_6236,N_1988,N_3847);
nor U6237 (N_6237,N_3812,N_1628);
or U6238 (N_6238,N_684,N_3282);
nor U6239 (N_6239,N_3909,N_922);
and U6240 (N_6240,N_2353,N_4041);
nand U6241 (N_6241,N_4869,N_2067);
xor U6242 (N_6242,N_2070,N_3115);
or U6243 (N_6243,N_1577,N_1334);
xor U6244 (N_6244,N_2671,N_1656);
nor U6245 (N_6245,N_2348,N_1714);
nor U6246 (N_6246,N_2404,N_4791);
xor U6247 (N_6247,N_1037,N_2669);
or U6248 (N_6248,N_4319,N_63);
nor U6249 (N_6249,N_1677,N_1224);
nor U6250 (N_6250,N_459,N_1786);
nand U6251 (N_6251,N_3972,N_3761);
xnor U6252 (N_6252,N_4135,N_4956);
nor U6253 (N_6253,N_3819,N_2417);
and U6254 (N_6254,N_12,N_2195);
and U6255 (N_6255,N_4021,N_160);
nand U6256 (N_6256,N_4342,N_4812);
nand U6257 (N_6257,N_2326,N_3291);
nor U6258 (N_6258,N_3807,N_3391);
or U6259 (N_6259,N_2580,N_72);
nor U6260 (N_6260,N_158,N_880);
nor U6261 (N_6261,N_2699,N_2377);
or U6262 (N_6262,N_2705,N_3234);
nand U6263 (N_6263,N_2730,N_4942);
or U6264 (N_6264,N_3306,N_2928);
and U6265 (N_6265,N_3104,N_4789);
or U6266 (N_6266,N_4245,N_2863);
nor U6267 (N_6267,N_310,N_460);
nand U6268 (N_6268,N_4994,N_3202);
xor U6269 (N_6269,N_198,N_2266);
xnor U6270 (N_6270,N_2153,N_4269);
and U6271 (N_6271,N_3052,N_15);
nor U6272 (N_6272,N_1805,N_556);
or U6273 (N_6273,N_2790,N_1327);
xor U6274 (N_6274,N_3349,N_1129);
nand U6275 (N_6275,N_1840,N_688);
nand U6276 (N_6276,N_2512,N_1140);
nand U6277 (N_6277,N_3087,N_4748);
or U6278 (N_6278,N_1512,N_2476);
nand U6279 (N_6279,N_321,N_4530);
xor U6280 (N_6280,N_2892,N_2025);
nand U6281 (N_6281,N_608,N_1186);
nor U6282 (N_6282,N_1290,N_3120);
nor U6283 (N_6283,N_1117,N_134);
nor U6284 (N_6284,N_4627,N_2439);
or U6285 (N_6285,N_3047,N_3364);
and U6286 (N_6286,N_3176,N_1044);
nor U6287 (N_6287,N_1257,N_3337);
or U6288 (N_6288,N_318,N_4694);
and U6289 (N_6289,N_93,N_3400);
or U6290 (N_6290,N_43,N_4274);
nand U6291 (N_6291,N_468,N_2452);
and U6292 (N_6292,N_3980,N_977);
nor U6293 (N_6293,N_4833,N_1942);
nor U6294 (N_6294,N_4726,N_1431);
or U6295 (N_6295,N_1779,N_1352);
xor U6296 (N_6296,N_1752,N_1058);
nand U6297 (N_6297,N_1279,N_1360);
nand U6298 (N_6298,N_1921,N_3845);
and U6299 (N_6299,N_451,N_147);
or U6300 (N_6300,N_4191,N_3458);
nor U6301 (N_6301,N_899,N_2500);
and U6302 (N_6302,N_1761,N_672);
nand U6303 (N_6303,N_2464,N_995);
and U6304 (N_6304,N_1021,N_2549);
xnor U6305 (N_6305,N_4637,N_2056);
or U6306 (N_6306,N_4421,N_1562);
or U6307 (N_6307,N_170,N_3041);
and U6308 (N_6308,N_3963,N_4005);
nor U6309 (N_6309,N_4884,N_342);
nor U6310 (N_6310,N_1806,N_3675);
and U6311 (N_6311,N_952,N_929);
nor U6312 (N_6312,N_1410,N_2576);
nand U6313 (N_6313,N_399,N_1024);
nand U6314 (N_6314,N_1825,N_3833);
xnor U6315 (N_6315,N_1981,N_3218);
or U6316 (N_6316,N_4371,N_3092);
nand U6317 (N_6317,N_2992,N_2885);
nor U6318 (N_6318,N_4413,N_1615);
nor U6319 (N_6319,N_873,N_2560);
or U6320 (N_6320,N_314,N_4798);
or U6321 (N_6321,N_2190,N_1973);
and U6322 (N_6322,N_4880,N_1913);
xnor U6323 (N_6323,N_1150,N_4271);
and U6324 (N_6324,N_2436,N_1691);
or U6325 (N_6325,N_760,N_3987);
nand U6326 (N_6326,N_2726,N_642);
nand U6327 (N_6327,N_4171,N_1451);
and U6328 (N_6328,N_3774,N_4546);
or U6329 (N_6329,N_557,N_3722);
or U6330 (N_6330,N_537,N_1716);
nor U6331 (N_6331,N_1243,N_2509);
or U6332 (N_6332,N_4536,N_2791);
or U6333 (N_6333,N_1053,N_2026);
nand U6334 (N_6334,N_1905,N_320);
nor U6335 (N_6335,N_3034,N_1784);
xor U6336 (N_6336,N_1120,N_3250);
and U6337 (N_6337,N_3000,N_3455);
and U6338 (N_6338,N_1930,N_1187);
and U6339 (N_6339,N_4740,N_313);
or U6340 (N_6340,N_1436,N_3388);
or U6341 (N_6341,N_884,N_871);
xor U6342 (N_6342,N_288,N_103);
or U6343 (N_6343,N_1924,N_2385);
xnor U6344 (N_6344,N_655,N_3966);
and U6345 (N_6345,N_2918,N_105);
or U6346 (N_6346,N_3620,N_2050);
or U6347 (N_6347,N_3100,N_4520);
and U6348 (N_6348,N_4706,N_2240);
xnor U6349 (N_6349,N_591,N_2999);
nand U6350 (N_6350,N_686,N_3348);
nand U6351 (N_6351,N_4355,N_850);
nand U6352 (N_6352,N_752,N_2188);
nand U6353 (N_6353,N_2859,N_2597);
nand U6354 (N_6354,N_4769,N_1517);
nor U6355 (N_6355,N_4577,N_3645);
xnor U6356 (N_6356,N_2327,N_1871);
xor U6357 (N_6357,N_967,N_3209);
xnor U6358 (N_6358,N_795,N_2795);
xor U6359 (N_6359,N_822,N_1465);
nand U6360 (N_6360,N_3420,N_234);
nand U6361 (N_6361,N_1401,N_1505);
xnor U6362 (N_6362,N_3238,N_805);
or U6363 (N_6363,N_3312,N_3017);
and U6364 (N_6364,N_2249,N_135);
or U6365 (N_6365,N_1169,N_3161);
xor U6366 (N_6366,N_4799,N_2694);
xnor U6367 (N_6367,N_1598,N_723);
or U6368 (N_6368,N_2890,N_758);
and U6369 (N_6369,N_930,N_3200);
and U6370 (N_6370,N_2449,N_1456);
nand U6371 (N_6371,N_3457,N_3874);
xnor U6372 (N_6372,N_2880,N_3986);
xor U6373 (N_6373,N_2852,N_4592);
nand U6374 (N_6374,N_253,N_2517);
and U6375 (N_6375,N_95,N_2738);
xor U6376 (N_6376,N_3714,N_3448);
and U6377 (N_6377,N_1687,N_1424);
and U6378 (N_6378,N_4639,N_4961);
or U6379 (N_6379,N_4641,N_979);
nand U6380 (N_6380,N_3708,N_4463);
xnor U6381 (N_6381,N_1590,N_1226);
nand U6382 (N_6382,N_1854,N_438);
nor U6383 (N_6383,N_1175,N_410);
xor U6384 (N_6384,N_2716,N_1828);
xor U6385 (N_6385,N_1575,N_2232);
or U6386 (N_6386,N_2985,N_2673);
xnor U6387 (N_6387,N_3561,N_1879);
and U6388 (N_6388,N_4377,N_1722);
nand U6389 (N_6389,N_374,N_2440);
nand U6390 (N_6390,N_4763,N_2884);
and U6391 (N_6391,N_2468,N_2002);
or U6392 (N_6392,N_2163,N_4805);
nor U6393 (N_6393,N_323,N_2359);
xor U6394 (N_6394,N_2491,N_2772);
nor U6395 (N_6395,N_1350,N_1233);
nand U6396 (N_6396,N_4197,N_3011);
nor U6397 (N_6397,N_4887,N_4452);
nor U6398 (N_6398,N_1068,N_3059);
or U6399 (N_6399,N_552,N_3485);
nand U6400 (N_6400,N_500,N_2923);
or U6401 (N_6401,N_1025,N_4239);
or U6402 (N_6402,N_834,N_166);
nor U6403 (N_6403,N_4919,N_2010);
or U6404 (N_6404,N_4265,N_1059);
nand U6405 (N_6405,N_2097,N_931);
nor U6406 (N_6406,N_484,N_3917);
nor U6407 (N_6407,N_509,N_1028);
xor U6408 (N_6408,N_3853,N_258);
xnor U6409 (N_6409,N_2924,N_1011);
or U6410 (N_6410,N_4386,N_4294);
nor U6411 (N_6411,N_4394,N_1214);
nand U6412 (N_6412,N_604,N_842);
nand U6413 (N_6413,N_3380,N_573);
and U6414 (N_6414,N_2071,N_3568);
nand U6415 (N_6415,N_2199,N_1693);
or U6416 (N_6416,N_3014,N_2978);
xor U6417 (N_6417,N_2961,N_1204);
xor U6418 (N_6418,N_810,N_1902);
xor U6419 (N_6419,N_3068,N_21);
nor U6420 (N_6420,N_1978,N_2583);
or U6421 (N_6421,N_3605,N_982);
and U6422 (N_6422,N_2209,N_1782);
and U6423 (N_6423,N_212,N_163);
nand U6424 (N_6424,N_895,N_3832);
nor U6425 (N_6425,N_2331,N_2068);
and U6426 (N_6426,N_2251,N_1240);
and U6427 (N_6427,N_1758,N_3089);
nor U6428 (N_6428,N_2290,N_2614);
and U6429 (N_6429,N_2384,N_2638);
xor U6430 (N_6430,N_2558,N_2941);
nor U6431 (N_6431,N_2288,N_2769);
nor U6432 (N_6432,N_3393,N_4575);
or U6433 (N_6433,N_4323,N_2807);
xnor U6434 (N_6434,N_630,N_919);
nand U6435 (N_6435,N_4086,N_3530);
and U6436 (N_6436,N_3150,N_2842);
and U6437 (N_6437,N_633,N_1595);
xor U6438 (N_6438,N_1105,N_3352);
or U6439 (N_6439,N_4574,N_4457);
nand U6440 (N_6440,N_322,N_2443);
and U6441 (N_6441,N_830,N_2197);
nand U6442 (N_6442,N_2215,N_2285);
nand U6443 (N_6443,N_4081,N_369);
and U6444 (N_6444,N_4315,N_3554);
xor U6445 (N_6445,N_1778,N_1747);
or U6446 (N_6446,N_1895,N_49);
or U6447 (N_6447,N_2981,N_2392);
xor U6448 (N_6448,N_2634,N_4524);
nor U6449 (N_6449,N_3746,N_3747);
and U6450 (N_6450,N_300,N_3689);
nor U6451 (N_6451,N_4387,N_2573);
and U6452 (N_6452,N_1076,N_4296);
and U6453 (N_6453,N_2115,N_3409);
xor U6454 (N_6454,N_239,N_246);
nor U6455 (N_6455,N_51,N_2545);
and U6456 (N_6456,N_767,N_3703);
and U6457 (N_6457,N_2332,N_1963);
nand U6458 (N_6458,N_477,N_2283);
or U6459 (N_6459,N_4035,N_4439);
nor U6460 (N_6460,N_4787,N_1004);
nor U6461 (N_6461,N_1645,N_4985);
nor U6462 (N_6462,N_2349,N_2233);
nand U6463 (N_6463,N_2008,N_3946);
nand U6464 (N_6464,N_1812,N_1507);
and U6465 (N_6465,N_1508,N_809);
xnor U6466 (N_6466,N_2603,N_2293);
or U6467 (N_6467,N_3354,N_2210);
nand U6468 (N_6468,N_1749,N_337);
nand U6469 (N_6469,N_3524,N_2196);
and U6470 (N_6470,N_1351,N_4015);
nand U6471 (N_6471,N_8,N_2170);
nor U6472 (N_6472,N_2598,N_4194);
nand U6473 (N_6473,N_4663,N_3721);
and U6474 (N_6474,N_3162,N_1926);
xnor U6475 (N_6475,N_4153,N_1337);
and U6476 (N_6476,N_2481,N_3816);
nor U6477 (N_6477,N_587,N_2775);
nand U6478 (N_6478,N_2537,N_1567);
nor U6479 (N_6479,N_1530,N_3116);
xor U6480 (N_6480,N_881,N_4331);
nor U6481 (N_6481,N_1225,N_3423);
or U6482 (N_6482,N_868,N_1088);
xnor U6483 (N_6483,N_4950,N_218);
or U6484 (N_6484,N_2269,N_2713);
nand U6485 (N_6485,N_1664,N_184);
nand U6486 (N_6486,N_2141,N_3077);
nor U6487 (N_6487,N_2881,N_1342);
or U6488 (N_6488,N_28,N_4238);
and U6489 (N_6489,N_1966,N_3667);
xor U6490 (N_6490,N_2155,N_3379);
xor U6491 (N_6491,N_1608,N_2946);
or U6492 (N_6492,N_3155,N_1261);
or U6493 (N_6493,N_1357,N_329);
xor U6494 (N_6494,N_3639,N_954);
or U6495 (N_6495,N_3686,N_3778);
or U6496 (N_6496,N_844,N_3142);
nand U6497 (N_6497,N_4669,N_992);
and U6498 (N_6498,N_1416,N_3384);
xor U6499 (N_6499,N_1968,N_104);
and U6500 (N_6500,N_3951,N_3983);
nor U6501 (N_6501,N_435,N_3426);
nand U6502 (N_6502,N_4464,N_2768);
and U6503 (N_6503,N_2189,N_4111);
or U6504 (N_6504,N_4657,N_785);
and U6505 (N_6505,N_3929,N_4852);
xor U6506 (N_6506,N_3245,N_3219);
xnor U6507 (N_6507,N_1686,N_1118);
nor U6508 (N_6508,N_4266,N_527);
nor U6509 (N_6509,N_3392,N_2581);
or U6510 (N_6510,N_4533,N_1314);
nand U6511 (N_6511,N_4731,N_609);
nand U6512 (N_6512,N_4037,N_226);
and U6513 (N_6513,N_1425,N_164);
and U6514 (N_6514,N_4973,N_3093);
or U6515 (N_6515,N_1570,N_3884);
nor U6516 (N_6516,N_701,N_2159);
or U6517 (N_6517,N_2393,N_3399);
nor U6518 (N_6518,N_496,N_3303);
xor U6519 (N_6519,N_1482,N_4851);
and U6520 (N_6520,N_3936,N_3735);
and U6521 (N_6521,N_942,N_1478);
nor U6522 (N_6522,N_2777,N_3428);
xnor U6523 (N_6523,N_1541,N_1110);
nor U6524 (N_6524,N_1629,N_4776);
xor U6525 (N_6525,N_3318,N_4330);
or U6526 (N_6526,N_1180,N_4112);
or U6527 (N_6527,N_3450,N_1800);
and U6528 (N_6528,N_1881,N_4486);
and U6529 (N_6529,N_1057,N_1943);
and U6530 (N_6530,N_331,N_847);
xor U6531 (N_6531,N_590,N_3706);
or U6532 (N_6532,N_3930,N_3650);
nand U6533 (N_6533,N_817,N_4854);
xor U6534 (N_6534,N_2157,N_4583);
and U6535 (N_6535,N_2281,N_4022);
nand U6536 (N_6536,N_1417,N_1316);
xor U6537 (N_6537,N_2333,N_3326);
and U6538 (N_6538,N_4065,N_4986);
or U6539 (N_6539,N_4068,N_1519);
and U6540 (N_6540,N_1715,N_1336);
or U6541 (N_6541,N_2556,N_4510);
xor U6542 (N_6542,N_2687,N_2813);
xnor U6543 (N_6543,N_3914,N_584);
nand U6544 (N_6544,N_4691,N_4099);
and U6545 (N_6545,N_4272,N_237);
and U6546 (N_6546,N_4665,N_4053);
nand U6547 (N_6547,N_1060,N_4745);
and U6548 (N_6548,N_1222,N_4514);
nand U6549 (N_6549,N_897,N_539);
xor U6550 (N_6550,N_2930,N_485);
nand U6551 (N_6551,N_4392,N_3359);
or U6552 (N_6552,N_4793,N_546);
nand U6553 (N_6553,N_1273,N_1256);
nor U6554 (N_6554,N_289,N_3230);
xor U6555 (N_6555,N_3345,N_882);
nor U6556 (N_6556,N_1760,N_4595);
xnor U6557 (N_6557,N_3567,N_1744);
or U6558 (N_6558,N_3021,N_3454);
nor U6559 (N_6559,N_395,N_416);
or U6560 (N_6560,N_182,N_3117);
xor U6561 (N_6561,N_869,N_387);
or U6562 (N_6562,N_2737,N_3821);
nand U6563 (N_6563,N_4165,N_757);
and U6564 (N_6564,N_426,N_4254);
and U6565 (N_6565,N_4773,N_3758);
and U6566 (N_6566,N_1151,N_3701);
nand U6567 (N_6567,N_4714,N_4975);
nand U6568 (N_6568,N_3431,N_4747);
and U6569 (N_6569,N_2301,N_224);
or U6570 (N_6570,N_3044,N_4615);
nand U6571 (N_6571,N_200,N_4402);
xnor U6572 (N_6572,N_1497,N_4287);
nor U6573 (N_6573,N_774,N_674);
xor U6574 (N_6574,N_2568,N_3412);
nand U6575 (N_6575,N_4705,N_3193);
or U6576 (N_6576,N_27,N_2741);
nor U6577 (N_6577,N_2126,N_2);
xnor U6578 (N_6578,N_1841,N_3083);
nor U6579 (N_6579,N_55,N_4813);
xnor U6580 (N_6580,N_3615,N_4649);
xnor U6581 (N_6581,N_3899,N_1623);
or U6582 (N_6582,N_1271,N_708);
and U6583 (N_6583,N_1568,N_2900);
or U6584 (N_6584,N_3626,N_754);
nand U6585 (N_6585,N_2328,N_2913);
nor U6586 (N_6586,N_559,N_2138);
xor U6587 (N_6587,N_1372,N_2729);
and U6588 (N_6588,N_2587,N_211);
nand U6589 (N_6589,N_4124,N_3020);
nor U6590 (N_6590,N_4828,N_1948);
and U6591 (N_6591,N_4638,N_2979);
and U6592 (N_6592,N_4027,N_973);
nand U6593 (N_6593,N_2938,N_3659);
or U6594 (N_6594,N_2988,N_4562);
xor U6595 (N_6595,N_2677,N_2849);
or U6596 (N_6596,N_1365,N_1538);
xor U6597 (N_6597,N_3164,N_4785);
nor U6598 (N_6598,N_2815,N_3536);
xnor U6599 (N_6599,N_2770,N_4414);
xor U6600 (N_6600,N_2208,N_3811);
xor U6601 (N_6601,N_2222,N_3792);
or U6602 (N_6602,N_1995,N_1331);
xnor U6603 (N_6603,N_1269,N_203);
nand U6604 (N_6604,N_3057,N_397);
xor U6605 (N_6605,N_1094,N_2692);
nand U6606 (N_6606,N_1803,N_2490);
or U6607 (N_6607,N_825,N_4226);
nand U6608 (N_6608,N_4941,N_690);
and U6609 (N_6609,N_1181,N_2679);
xor U6610 (N_6610,N_2508,N_3096);
and U6611 (N_6611,N_549,N_19);
or U6612 (N_6612,N_1063,N_2809);
nand U6613 (N_6613,N_3952,N_1048);
xnor U6614 (N_6614,N_963,N_3447);
nor U6615 (N_6615,N_3739,N_4190);
xnor U6616 (N_6616,N_1706,N_2766);
or U6617 (N_6617,N_4036,N_1087);
nand U6618 (N_6618,N_3182,N_3367);
and U6619 (N_6619,N_1878,N_1814);
and U6620 (N_6620,N_1582,N_3206);
and U6621 (N_6621,N_455,N_2202);
nor U6622 (N_6622,N_4224,N_316);
and U6623 (N_6623,N_2850,N_1684);
xor U6624 (N_6624,N_2652,N_1857);
nor U6625 (N_6625,N_4860,N_2502);
xnor U6626 (N_6626,N_35,N_4125);
and U6627 (N_6627,N_2094,N_2012);
xnor U6628 (N_6628,N_1437,N_3843);
nor U6629 (N_6629,N_2688,N_4307);
nand U6630 (N_6630,N_2386,N_488);
xor U6631 (N_6631,N_2945,N_3892);
xor U6632 (N_6632,N_3133,N_199);
nand U6633 (N_6633,N_2031,N_432);
or U6634 (N_6634,N_3603,N_3281);
or U6635 (N_6635,N_3313,N_2736);
nor U6636 (N_6636,N_4777,N_3913);
or U6637 (N_6637,N_1584,N_4102);
nand U6638 (N_6638,N_1455,N_3661);
and U6639 (N_6639,N_1643,N_2229);
and U6640 (N_6640,N_695,N_25);
nand U6641 (N_6641,N_1089,N_3300);
or U6642 (N_6642,N_3297,N_864);
xnor U6643 (N_6643,N_1404,N_4898);
or U6644 (N_6644,N_2613,N_3634);
xor U6645 (N_6645,N_431,N_4477);
xnor U6646 (N_6646,N_4083,N_1578);
or U6647 (N_6647,N_920,N_3592);
nand U6648 (N_6648,N_1127,N_3631);
and U6649 (N_6649,N_1133,N_4820);
nand U6650 (N_6650,N_3949,N_3427);
nor U6651 (N_6651,N_1292,N_1285);
and U6652 (N_6652,N_513,N_2360);
xor U6653 (N_6653,N_2035,N_1038);
nand U6654 (N_6654,N_1438,N_3583);
nor U6655 (N_6655,N_4019,N_3347);
nand U6656 (N_6656,N_3442,N_2256);
and U6657 (N_6657,N_4900,N_2915);
xor U6658 (N_6658,N_1394,N_1547);
nor U6659 (N_6659,N_4314,N_4075);
xor U6660 (N_6660,N_838,N_4493);
and U6661 (N_6661,N_3904,N_4350);
nand U6662 (N_6662,N_1116,N_3495);
and U6663 (N_6663,N_4436,N_3954);
nor U6664 (N_6664,N_1396,N_3785);
xor U6665 (N_6665,N_4121,N_3288);
and U6666 (N_6666,N_2486,N_1866);
nor U6667 (N_6667,N_4337,N_1253);
and U6668 (N_6668,N_2971,N_1741);
nand U6669 (N_6669,N_4656,N_4761);
nand U6670 (N_6670,N_4450,N_4678);
nor U6671 (N_6671,N_2133,N_541);
xor U6672 (N_6672,N_4633,N_4913);
or U6673 (N_6673,N_4379,N_2257);
nor U6674 (N_6674,N_3941,N_2916);
or U6675 (N_6675,N_4338,N_3818);
nor U6676 (N_6676,N_4930,N_336);
xnor U6677 (N_6677,N_2304,N_3043);
xor U6678 (N_6678,N_2519,N_3665);
and U6679 (N_6679,N_2379,N_4440);
and U6680 (N_6680,N_1873,N_131);
nand U6681 (N_6681,N_890,N_1984);
nand U6682 (N_6682,N_4794,N_620);
nand U6683 (N_6683,N_1330,N_4087);
nand U6684 (N_6684,N_1764,N_1839);
nor U6685 (N_6685,N_302,N_4965);
or U6686 (N_6686,N_446,N_3271);
nand U6687 (N_6687,N_3046,N_83);
or U6688 (N_6688,N_2112,N_2864);
or U6689 (N_6689,N_2538,N_3353);
and U6690 (N_6690,N_2906,N_980);
or U6691 (N_6691,N_1251,N_3751);
or U6692 (N_6692,N_1667,N_1768);
and U6693 (N_6693,N_4529,N_1146);
nand U6694 (N_6694,N_4979,N_1430);
or U6695 (N_6695,N_1522,N_2341);
xnor U6696 (N_6696,N_4152,N_2709);
xnor U6697 (N_6697,N_4048,N_1794);
and U6698 (N_6698,N_137,N_536);
nor U6699 (N_6699,N_1540,N_4554);
and U6700 (N_6700,N_2952,N_1614);
nor U6701 (N_6701,N_4548,N_1183);
and U6702 (N_6702,N_279,N_4912);
and U6703 (N_6703,N_362,N_814);
xnor U6704 (N_6704,N_4250,N_2045);
xnor U6705 (N_6705,N_2779,N_1961);
nor U6706 (N_6706,N_4378,N_3221);
xnor U6707 (N_6707,N_2125,N_2096);
xor U6708 (N_6708,N_2498,N_1622);
and U6709 (N_6709,N_1955,N_4088);
xor U6710 (N_6710,N_3376,N_3461);
nor U6711 (N_6711,N_1167,N_4720);
nand U6712 (N_6712,N_1286,N_689);
xor U6713 (N_6713,N_1654,N_3911);
and U6714 (N_6714,N_1555,N_119);
nand U6715 (N_6715,N_3856,N_1858);
nand U6716 (N_6716,N_3277,N_3058);
nand U6717 (N_6717,N_3990,N_4092);
or U6718 (N_6718,N_1877,N_4363);
or U6719 (N_6719,N_251,N_2013);
xor U6720 (N_6720,N_3791,N_3189);
and U6721 (N_6721,N_2387,N_1892);
nor U6722 (N_6722,N_3753,N_3563);
nand U6723 (N_6723,N_2618,N_4568);
nor U6724 (N_6724,N_4202,N_1262);
nor U6725 (N_6725,N_3838,N_4427);
and U6726 (N_6726,N_946,N_4262);
or U6727 (N_6727,N_4952,N_1252);
and U6728 (N_6728,N_4185,N_3920);
or U6729 (N_6729,N_4911,N_1692);
nor U6730 (N_6730,N_140,N_1591);
and U6731 (N_6731,N_402,N_3003);
or U6732 (N_6732,N_4809,N_16);
xnor U6733 (N_6733,N_1428,N_1373);
and U6734 (N_6734,N_2865,N_2994);
nand U6735 (N_6735,N_915,N_3926);
or U6736 (N_6736,N_2607,N_180);
or U6737 (N_6737,N_222,N_1407);
nand U6738 (N_6738,N_1413,N_3110);
nor U6739 (N_6739,N_2838,N_1244);
or U6740 (N_6740,N_1426,N_1363);
xor U6741 (N_6741,N_3664,N_2982);
or U6742 (N_6742,N_3028,N_161);
and U6743 (N_6743,N_968,N_1370);
nand U6744 (N_6744,N_4011,N_2877);
nor U6745 (N_6745,N_649,N_3609);
xnor U6746 (N_6746,N_2063,N_4328);
or U6747 (N_6747,N_3341,N_1673);
xor U6748 (N_6748,N_3280,N_3593);
nor U6749 (N_6749,N_1859,N_2948);
nand U6750 (N_6750,N_4718,N_4423);
xnor U6751 (N_6751,N_1957,N_961);
and U6752 (N_6752,N_4661,N_3560);
xnor U6753 (N_6753,N_365,N_2205);
xnor U6754 (N_6754,N_4183,N_229);
nand U6755 (N_6755,N_3787,N_1824);
xnor U6756 (N_6756,N_3830,N_1672);
or U6757 (N_6757,N_4215,N_3759);
nand U6758 (N_6758,N_3862,N_4465);
or U6759 (N_6759,N_2987,N_2255);
xor U6760 (N_6760,N_3246,N_434);
nor U6761 (N_6761,N_1276,N_4877);
nand U6762 (N_6762,N_826,N_3551);
nor U6763 (N_6763,N_124,N_3888);
or U6764 (N_6764,N_3793,N_80);
xor U6765 (N_6765,N_3547,N_3170);
nor U6766 (N_6766,N_4045,N_3575);
or U6767 (N_6767,N_38,N_1270);
nand U6768 (N_6768,N_2032,N_3642);
nor U6769 (N_6769,N_2187,N_3060);
or U6770 (N_6770,N_2771,N_4966);
nor U6771 (N_6771,N_2442,N_109);
and U6772 (N_6772,N_443,N_3624);
nor U6773 (N_6773,N_1729,N_4550);
nor U6774 (N_6774,N_3468,N_2434);
xor U6775 (N_6775,N_738,N_3957);
or U6776 (N_6776,N_2098,N_4505);
nor U6777 (N_6777,N_1670,N_2142);
and U6778 (N_6778,N_3871,N_668);
xor U6779 (N_6779,N_48,N_3971);
or U6780 (N_6780,N_1156,N_2487);
xnor U6781 (N_6781,N_3906,N_2374);
nor U6782 (N_6782,N_2365,N_4360);
xnor U6783 (N_6783,N_53,N_3823);
nand U6784 (N_6784,N_4049,N_1339);
and U6785 (N_6785,N_471,N_1079);
xor U6786 (N_6786,N_4702,N_2528);
nand U6787 (N_6787,N_2872,N_2073);
xor U6788 (N_6788,N_3526,N_3654);
nor U6789 (N_6789,N_3260,N_3365);
nor U6790 (N_6790,N_784,N_514);
and U6791 (N_6791,N_2665,N_1104);
or U6792 (N_6792,N_3727,N_658);
nor U6793 (N_6793,N_4023,N_3730);
nand U6794 (N_6794,N_4385,N_1699);
nor U6795 (N_6795,N_583,N_4007);
nor U6796 (N_6796,N_4313,N_1440);
or U6797 (N_6797,N_4679,N_296);
or U6798 (N_6798,N_2077,N_1573);
nor U6799 (N_6799,N_1837,N_3851);
nor U6800 (N_6800,N_2312,N_4810);
nand U6801 (N_6801,N_1566,N_4244);
nand U6802 (N_6802,N_3272,N_2661);
and U6803 (N_6803,N_4743,N_4446);
and U6804 (N_6804,N_2121,N_2645);
nor U6805 (N_6805,N_801,N_3519);
and U6806 (N_6806,N_1618,N_493);
or U6807 (N_6807,N_47,N_4300);
or U6808 (N_6808,N_4336,N_4499);
and U6809 (N_6809,N_3079,N_1481);
nor U6810 (N_6810,N_2898,N_2821);
xor U6811 (N_6811,N_715,N_3590);
and U6812 (N_6812,N_2663,N_530);
and U6813 (N_6813,N_639,N_1358);
or U6814 (N_6814,N_2954,N_4051);
and U6815 (N_6815,N_4817,N_3989);
xnor U6816 (N_6816,N_3900,N_338);
or U6817 (N_6817,N_3974,N_1865);
or U6818 (N_6818,N_2370,N_1122);
xnor U6819 (N_6819,N_187,N_1050);
nor U6820 (N_6820,N_2338,N_1178);
nand U6821 (N_6821,N_1061,N_3984);
or U6822 (N_6822,N_2428,N_687);
xnor U6823 (N_6823,N_3075,N_2518);
nand U6824 (N_6824,N_4517,N_1299);
and U6825 (N_6825,N_3910,N_3940);
and U6826 (N_6826,N_357,N_4400);
or U6827 (N_6827,N_1103,N_2721);
nor U6828 (N_6828,N_3135,N_4578);
nor U6829 (N_6829,N_3694,N_4060);
or U6830 (N_6830,N_1210,N_2315);
nand U6831 (N_6831,N_1795,N_2659);
nor U6832 (N_6832,N_4082,N_851);
and U6833 (N_6833,N_1712,N_2345);
nor U6834 (N_6834,N_3713,N_3505);
xnor U6835 (N_6835,N_1484,N_2106);
xor U6836 (N_6836,N_2670,N_3923);
nand U6837 (N_6837,N_2245,N_40);
and U6838 (N_6838,N_4397,N_4418);
or U6839 (N_6839,N_762,N_888);
nor U6840 (N_6840,N_1599,N_2760);
and U6841 (N_6841,N_332,N_1906);
or U6842 (N_6842,N_3144,N_2124);
nor U6843 (N_6843,N_2682,N_1769);
or U6844 (N_6844,N_4144,N_3682);
or U6845 (N_6845,N_3653,N_2793);
and U6846 (N_6846,N_3729,N_4749);
nor U6847 (N_6847,N_4916,N_670);
and U6848 (N_6848,N_4447,N_1569);
xnor U6849 (N_6849,N_673,N_1683);
and U6850 (N_6850,N_542,N_1340);
nand U6851 (N_6851,N_3217,N_1302);
and U6852 (N_6852,N_1035,N_2612);
xnor U6853 (N_6853,N_3370,N_3236);
and U6854 (N_6854,N_964,N_3849);
nand U6855 (N_6855,N_1646,N_3243);
and U6856 (N_6856,N_2236,N_2858);
nor U6857 (N_6857,N_1047,N_1970);
nand U6858 (N_6858,N_3781,N_56);
or U6859 (N_6859,N_62,N_3881);
and U6860 (N_6860,N_173,N_4280);
or U6861 (N_6861,N_3443,N_2707);
or U6862 (N_6862,N_1531,N_1872);
xnor U6863 (N_6863,N_2472,N_1378);
nand U6864 (N_6864,N_1777,N_2697);
nand U6865 (N_6865,N_2437,N_4070);
and U6866 (N_6866,N_2477,N_141);
nand U6867 (N_6867,N_4781,N_389);
or U6868 (N_6868,N_3290,N_129);
nor U6869 (N_6869,N_778,N_1489);
and U6870 (N_6870,N_1561,N_3025);
nand U6871 (N_6871,N_2041,N_2400);
or U6872 (N_6872,N_4409,N_3700);
and U6873 (N_6873,N_4918,N_4806);
xnor U6874 (N_6874,N_1610,N_2693);
or U6875 (N_6875,N_1356,N_2691);
or U6876 (N_6876,N_1081,N_4865);
and U6877 (N_6877,N_3925,N_3398);
or U6878 (N_6878,N_2320,N_3555);
nand U6879 (N_6879,N_792,N_4618);
nand U6880 (N_6880,N_3094,N_3256);
and U6881 (N_6881,N_993,N_1062);
nor U6882 (N_6882,N_423,N_3769);
xor U6883 (N_6883,N_3147,N_1674);
or U6884 (N_6884,N_327,N_4525);
nand U6885 (N_6885,N_2391,N_3279);
and U6886 (N_6886,N_2820,N_3566);
nand U6887 (N_6887,N_1284,N_2221);
and U6888 (N_6888,N_3961,N_4978);
or U6889 (N_6889,N_3711,N_2700);
and U6890 (N_6890,N_3697,N_2329);
or U6891 (N_6891,N_1149,N_4455);
xnor U6892 (N_6892,N_4349,N_2246);
or U6893 (N_6893,N_3508,N_2763);
xor U6894 (N_6894,N_3501,N_4188);
nor U6895 (N_6895,N_2408,N_2105);
or U6896 (N_6896,N_1767,N_1792);
xor U6897 (N_6897,N_326,N_2432);
xnor U6898 (N_6898,N_2672,N_619);
xor U6899 (N_6899,N_4937,N_3539);
nand U6900 (N_6900,N_3789,N_2565);
nor U6901 (N_6901,N_3743,N_3030);
xor U6902 (N_6902,N_2321,N_1612);
and U6903 (N_6903,N_2399,N_473);
and U6904 (N_6904,N_34,N_3912);
and U6905 (N_6905,N_1106,N_3229);
and U6906 (N_6906,N_392,N_1516);
and U6907 (N_6907,N_4569,N_4369);
and U6908 (N_6908,N_1354,N_1448);
xnor U6909 (N_6909,N_3088,N_4767);
nand U6910 (N_6910,N_1763,N_1838);
and U6911 (N_6911,N_3988,N_4734);
xor U6912 (N_6912,N_4482,N_568);
nor U6913 (N_6913,N_2514,N_2380);
or U6914 (N_6914,N_430,N_272);
nor U6915 (N_6915,N_4983,N_2960);
and U6916 (N_6916,N_2976,N_638);
nand U6917 (N_6917,N_3754,N_2785);
and U6918 (N_6918,N_3829,N_3969);
nand U6919 (N_6919,N_4417,N_4843);
nand U6920 (N_6920,N_2984,N_3622);
and U6921 (N_6921,N_4020,N_1804);
nor U6922 (N_6922,N_475,N_2429);
xnor U6923 (N_6923,N_1379,N_3657);
xnor U6924 (N_6924,N_2084,N_3992);
xnor U6925 (N_6925,N_3831,N_2369);
nor U6926 (N_6926,N_807,N_4899);
nor U6927 (N_6927,N_2445,N_4310);
xnor U6928 (N_6928,N_2372,N_2131);
xor U6929 (N_6929,N_210,N_4722);
xnor U6930 (N_6930,N_464,N_2451);
or U6931 (N_6931,N_116,N_2823);
nand U6932 (N_6932,N_265,N_142);
xor U6933 (N_6933,N_1208,N_1991);
and U6934 (N_6934,N_3361,N_1160);
nand U6935 (N_6935,N_599,N_4943);
nand U6936 (N_6936,N_3175,N_562);
xnor U6937 (N_6937,N_4553,N_4967);
or U6938 (N_6938,N_1952,N_4050);
nor U6939 (N_6939,N_2160,N_2323);
or U6940 (N_6940,N_1064,N_425);
xnor U6941 (N_6941,N_3040,N_4783);
nand U6942 (N_6942,N_3070,N_407);
nor U6943 (N_6943,N_4842,N_1005);
and U6944 (N_6944,N_3702,N_343);
nor U6945 (N_6945,N_2438,N_4210);
or U6946 (N_6946,N_11,N_3678);
nor U6947 (N_6947,N_3644,N_1335);
nand U6948 (N_6948,N_2220,N_798);
nand U6949 (N_6949,N_788,N_3167);
or U6950 (N_6950,N_1176,N_1492);
nand U6951 (N_6951,N_510,N_1016);
nor U6952 (N_6952,N_6,N_2137);
or U6953 (N_6953,N_2278,N_1188);
xnor U6954 (N_6954,N_1377,N_231);
xnor U6955 (N_6955,N_913,N_4540);
nand U6956 (N_6956,N_3520,N_3410);
xnor U6957 (N_6957,N_3502,N_159);
or U6958 (N_6958,N_1359,N_3086);
nor U6959 (N_6959,N_2555,N_1631);
or U6960 (N_6960,N_2078,N_3820);
and U6961 (N_6961,N_4473,N_240);
nor U6962 (N_6962,N_2873,N_2722);
and U6963 (N_6963,N_393,N_2744);
nand U6964 (N_6964,N_217,N_1476);
or U6965 (N_6965,N_2689,N_469);
xnor U6966 (N_6966,N_3589,N_734);
nand U6967 (N_6967,N_4915,N_350);
and U6968 (N_6968,N_4038,N_3959);
nor U6969 (N_6969,N_2828,N_3651);
or U6970 (N_6970,N_2590,N_346);
or U6971 (N_6971,N_3194,N_643);
and U6972 (N_6972,N_1041,N_1427);
nor U6973 (N_6973,N_1527,N_747);
nor U6974 (N_6974,N_3241,N_681);
xnor U6975 (N_6975,N_2397,N_1405);
xor U6976 (N_6976,N_4364,N_23);
or U6977 (N_6977,N_1052,N_1604);
nor U6978 (N_6978,N_2295,N_77);
and U6979 (N_6979,N_3947,N_4094);
or U6980 (N_6980,N_4253,N_499);
nor U6981 (N_6981,N_1552,N_3956);
nand U6982 (N_6982,N_3564,N_281);
nand U6983 (N_6983,N_4420,N_2062);
and U6984 (N_6984,N_2595,N_3991);
nor U6985 (N_6985,N_1884,N_143);
xor U6986 (N_6986,N_3525,N_4640);
and U6987 (N_6987,N_2109,N_4299);
or U6988 (N_6988,N_151,N_3066);
and U6989 (N_6989,N_4528,N_65);
nor U6990 (N_6990,N_845,N_2648);
and U6991 (N_6991,N_4667,N_4071);
xnor U6992 (N_6992,N_2082,N_1529);
or U6993 (N_6993,N_78,N_2497);
or U6994 (N_6994,N_3,N_4861);
or U6995 (N_6995,N_348,N_2102);
nand U6996 (N_6996,N_1874,N_4946);
and U6997 (N_6997,N_3532,N_3049);
and U6998 (N_6998,N_1836,N_1671);
nor U6999 (N_6999,N_4189,N_4243);
xnor U7000 (N_7000,N_2173,N_1289);
xor U7001 (N_7001,N_4358,N_2796);
nor U7002 (N_7002,N_577,N_1950);
and U7003 (N_7003,N_3836,N_3111);
xor U7004 (N_7004,N_2366,N_177);
xor U7005 (N_7005,N_3696,N_1258);
nor U7006 (N_7006,N_208,N_1705);
xnor U7007 (N_7007,N_2658,N_1247);
or U7008 (N_7008,N_4235,N_1406);
nand U7009 (N_7009,N_3452,N_4509);
or U7010 (N_7010,N_4623,N_4599);
nand U7011 (N_7011,N_3174,N_114);
nor U7012 (N_7012,N_86,N_1179);
and U7013 (N_7013,N_2441,N_965);
or U7014 (N_7014,N_764,N_1008);
nand U7015 (N_7015,N_2894,N_2416);
nor U7016 (N_7016,N_2922,N_2375);
xor U7017 (N_7017,N_2277,N_3927);
nor U7018 (N_7018,N_4237,N_2711);
nor U7019 (N_7019,N_2814,N_4606);
and U7020 (N_7020,N_2390,N_1807);
and U7021 (N_7021,N_3538,N_448);
xnor U7022 (N_7022,N_893,N_863);
nand U7023 (N_7023,N_1860,N_4882);
nor U7024 (N_7024,N_4521,N_1194);
xnor U7025 (N_7025,N_476,N_4267);
or U7026 (N_7026,N_1843,N_4628);
xor U7027 (N_7027,N_1485,N_3950);
xor U7028 (N_7028,N_4948,N_1589);
nor U7029 (N_7029,N_2171,N_1368);
and U7030 (N_7030,N_138,N_4468);
nor U7031 (N_7031,N_1217,N_790);
nand U7032 (N_7032,N_4766,N_4462);
xnor U7033 (N_7033,N_3933,N_1506);
or U7034 (N_7034,N_3528,N_2461);
or U7035 (N_7035,N_1098,N_4563);
nand U7036 (N_7036,N_2706,N_61);
or U7037 (N_7037,N_3803,N_1724);
and U7038 (N_7038,N_2505,N_1414);
and U7039 (N_7039,N_3790,N_2028);
nand U7040 (N_7040,N_2116,N_3475);
or U7041 (N_7041,N_256,N_2935);
or U7042 (N_7042,N_1851,N_3190);
xnor U7043 (N_7043,N_3038,N_4920);
nand U7044 (N_7044,N_270,N_1633);
nand U7045 (N_7045,N_1445,N_372);
nand U7046 (N_7046,N_4222,N_550);
xor U7047 (N_7047,N_4987,N_2798);
or U7048 (N_7048,N_1250,N_4393);
nand U7049 (N_7049,N_2076,N_938);
and U7050 (N_7050,N_2639,N_3641);
nor U7051 (N_7051,N_1287,N_1648);
or U7052 (N_7052,N_4687,N_2101);
nor U7053 (N_7053,N_721,N_3883);
or U7054 (N_7054,N_3511,N_4348);
or U7055 (N_7055,N_3192,N_1808);
nand U7056 (N_7056,N_1939,N_2764);
or U7057 (N_7057,N_1143,N_3102);
or U7058 (N_7058,N_2186,N_152);
nor U7059 (N_7059,N_4054,N_3064);
nand U7060 (N_7060,N_2931,N_2750);
xor U7061 (N_7061,N_3752,N_2817);
nand U7062 (N_7062,N_815,N_225);
xnor U7063 (N_7063,N_4712,N_2194);
or U7064 (N_7064,N_148,N_1483);
or U7065 (N_7065,N_4196,N_3124);
xor U7066 (N_7066,N_3289,N_751);
xnor U7067 (N_7067,N_2065,N_2489);
xor U7068 (N_7068,N_2139,N_4655);
and U7069 (N_7069,N_2778,N_282);
xnor U7070 (N_7070,N_1515,N_382);
nand U7071 (N_7071,N_4192,N_1666);
nor U7072 (N_7072,N_4732,N_3328);
xor U7073 (N_7073,N_3934,N_2695);
or U7074 (N_7074,N_2015,N_2644);
or U7075 (N_7075,N_2942,N_2182);
or U7076 (N_7076,N_1553,N_4585);
nand U7077 (N_7077,N_4855,N_853);
or U7078 (N_7078,N_593,N_3873);
or U7079 (N_7079,N_1152,N_2492);
nor U7080 (N_7080,N_3824,N_1993);
and U7081 (N_7081,N_128,N_1227);
nor U7082 (N_7082,N_2367,N_1033);
or U7083 (N_7083,N_1216,N_3424);
xor U7084 (N_7084,N_4329,N_4923);
xor U7085 (N_7085,N_624,N_1738);
nor U7086 (N_7086,N_4484,N_3510);
nor U7087 (N_7087,N_3898,N_1102);
xnor U7088 (N_7088,N_3584,N_3795);
nor U7089 (N_7089,N_478,N_1709);
nand U7090 (N_7090,N_398,N_614);
or U7091 (N_7091,N_1642,N_3390);
or U7092 (N_7092,N_4487,N_4757);
nor U7093 (N_7093,N_4380,N_2668);
nor U7094 (N_7094,N_4431,N_595);
nor U7095 (N_7095,N_1203,N_1780);
or U7096 (N_7096,N_4989,N_2841);
and U7097 (N_7097,N_1534,N_264);
xnor U7098 (N_7098,N_1689,N_1066);
and U7099 (N_7099,N_3839,N_3022);
or U7100 (N_7100,N_4619,N_1700);
and U7101 (N_7101,N_2712,N_4874);
nand U7102 (N_7102,N_2371,N_4792);
xor U7103 (N_7103,N_885,N_2211);
and U7104 (N_7104,N_4172,N_209);
and U7105 (N_7105,N_2043,N_3773);
or U7106 (N_7106,N_419,N_2119);
nor U7107 (N_7107,N_3082,N_2351);
xor U7108 (N_7108,N_4017,N_2430);
or U7109 (N_7109,N_3460,N_2599);
and U7110 (N_7110,N_2761,N_651);
and U7111 (N_7111,N_3415,N_4478);
nand U7112 (N_7112,N_1017,N_3308);
nor U7113 (N_7113,N_2848,N_4951);
and U7114 (N_7114,N_1126,N_2702);
nor U7115 (N_7115,N_2701,N_483);
nor U7116 (N_7116,N_4573,N_2422);
or U7117 (N_7117,N_4666,N_4105);
nor U7118 (N_7118,N_1,N_4862);
or U7119 (N_7119,N_2166,N_3854);
or U7120 (N_7120,N_4304,N_1200);
or U7121 (N_7121,N_494,N_115);
nand U7122 (N_7122,N_2058,N_3500);
or U7123 (N_7123,N_2085,N_3433);
nor U7124 (N_7124,N_2198,N_1900);
nor U7125 (N_7125,N_378,N_2592);
or U7126 (N_7126,N_1998,N_3332);
xor U7127 (N_7127,N_2557,N_1855);
xor U7128 (N_7128,N_3037,N_3688);
nor U7129 (N_7129,N_640,N_2336);
xnor U7130 (N_7130,N_641,N_803);
or U7131 (N_7131,N_2355,N_295);
nor U7132 (N_7132,N_523,N_4428);
or U7133 (N_7133,N_3489,N_1703);
nor U7134 (N_7134,N_1583,N_4306);
nor U7135 (N_7135,N_2806,N_4376);
nand U7136 (N_7136,N_905,N_4780);
nor U7137 (N_7137,N_1248,N_454);
and U7138 (N_7138,N_1545,N_2192);
and U7139 (N_7139,N_3242,N_1131);
nand U7140 (N_7140,N_3944,N_1398);
and U7141 (N_7141,N_3570,N_2561);
xnor U7142 (N_7142,N_358,N_4498);
nor U7143 (N_7143,N_2460,N_3441);
nor U7144 (N_7144,N_3496,N_2161);
and U7145 (N_7145,N_685,N_1264);
nand U7146 (N_7146,N_1315,N_2165);
or U7147 (N_7147,N_1801,N_4654);
and U7148 (N_7148,N_1992,N_4292);
and U7149 (N_7149,N_4630,N_4647);
nor U7150 (N_7150,N_1701,N_2563);
or U7151 (N_7151,N_4138,N_2427);
nor U7152 (N_7152,N_3637,N_429);
nor U7153 (N_7153,N_1423,N_4195);
nand U7154 (N_7154,N_4823,N_1533);
and U7155 (N_7155,N_2893,N_2424);
and U7156 (N_7156,N_79,N_4704);
or U7157 (N_7157,N_3292,N_1945);
nor U7158 (N_7158,N_4759,N_4046);
or U7159 (N_7159,N_1318,N_3097);
nor U7160 (N_7160,N_1882,N_836);
xnor U7161 (N_7161,N_4598,N_4873);
or U7162 (N_7162,N_1697,N_1291);
or U7163 (N_7163,N_2470,N_712);
or U7164 (N_7164,N_4609,N_2578);
nor U7165 (N_7165,N_3559,N_3652);
or U7166 (N_7166,N_4320,N_3173);
nand U7167 (N_7167,N_4807,N_349);
and U7168 (N_7168,N_3484,N_4067);
xnor U7169 (N_7169,N_2825,N_2088);
or U7170 (N_7170,N_3556,N_168);
xnor U7171 (N_7171,N_4980,N_984);
xor U7172 (N_7172,N_3136,N_3385);
nor U7173 (N_7173,N_1403,N_4291);
nor U7174 (N_7174,N_841,N_125);
xor U7175 (N_7175,N_2686,N_2457);
xnor U7176 (N_7176,N_4203,N_2357);
nor U7177 (N_7177,N_4626,N_2152);
nor U7178 (N_7178,N_325,N_545);
or U7179 (N_7179,N_2431,N_193);
nor U7180 (N_7180,N_2307,N_2388);
and U7181 (N_7181,N_2953,N_333);
nand U7182 (N_7182,N_554,N_1776);
xnor U7183 (N_7183,N_3248,N_692);
nor U7184 (N_7184,N_3286,N_1600);
and U7185 (N_7185,N_2410,N_3407);
and U7186 (N_7186,N_1580,N_2083);
xnor U7187 (N_7187,N_4090,N_4737);
and U7188 (N_7188,N_3016,N_2731);
nor U7189 (N_7189,N_1886,N_2891);
xnor U7190 (N_7190,N_4032,N_1572);
and U7191 (N_7191,N_2529,N_2479);
and U7192 (N_7192,N_889,N_714);
or U7193 (N_7193,N_3012,N_2871);
xnor U7194 (N_7194,N_1397,N_3062);
nand U7195 (N_7195,N_1694,N_1754);
or U7196 (N_7196,N_779,N_3425);
or U7197 (N_7197,N_2361,N_3340);
and U7198 (N_7198,N_4853,N_317);
nand U7199 (N_7199,N_1826,N_667);
xor U7200 (N_7200,N_3382,N_675);
and U7201 (N_7201,N_724,N_592);
and U7202 (N_7202,N_1159,N_1319);
nor U7203 (N_7203,N_3734,N_2757);
xor U7204 (N_7204,N_3577,N_99);
and U7205 (N_7205,N_1259,N_2956);
and U7206 (N_7206,N_894,N_191);
or U7207 (N_7207,N_2799,N_3128);
xor U7208 (N_7208,N_2134,N_3796);
or U7209 (N_7209,N_3886,N_3213);
xor U7210 (N_7210,N_4444,N_531);
and U7211 (N_7211,N_4696,N_1660);
xor U7212 (N_7212,N_4788,N_4485);
nand U7213 (N_7213,N_4091,N_2272);
nand U7214 (N_7214,N_4490,N_4025);
nor U7215 (N_7215,N_2347,N_4078);
and U7216 (N_7216,N_2933,N_1402);
nand U7217 (N_7217,N_4924,N_1556);
nand U7218 (N_7218,N_935,N_2787);
nor U7219 (N_7219,N_3660,N_3451);
or U7220 (N_7220,N_1559,N_2643);
and U7221 (N_7221,N_2425,N_746);
xnor U7222 (N_7222,N_2943,N_969);
nor U7223 (N_7223,N_2903,N_3619);
nor U7224 (N_7224,N_276,N_1023);
and U7225 (N_7225,N_4760,N_1311);
xnor U7226 (N_7226,N_843,N_2632);
xor U7227 (N_7227,N_4246,N_3005);
or U7228 (N_7228,N_799,N_3541);
and U7229 (N_7229,N_3748,N_4448);
xnor U7230 (N_7230,N_570,N_2414);
or U7231 (N_7231,N_4166,N_3323);
xor U7232 (N_7232,N_422,N_2975);
nor U7233 (N_7233,N_4648,N_278);
and U7234 (N_7234,N_4545,N_4927);
or U7235 (N_7235,N_3324,N_4662);
and U7236 (N_7236,N_4160,N_4858);
or U7237 (N_7237,N_1153,N_1593);
nand U7238 (N_7238,N_1863,N_3518);
nor U7239 (N_7239,N_702,N_827);
or U7240 (N_7240,N_766,N_3001);
nor U7241 (N_7241,N_2444,N_4744);
and U7242 (N_7242,N_3493,N_1894);
nand U7243 (N_7243,N_1718,N_1075);
and U7244 (N_7244,N_1458,N_172);
or U7245 (N_7245,N_3378,N_2308);
nor U7246 (N_7246,N_581,N_167);
nor U7247 (N_7247,N_285,N_3253);
or U7248 (N_7248,N_340,N_1548);
nor U7249 (N_7249,N_4122,N_4010);
and U7250 (N_7250,N_4821,N_4716);
or U7251 (N_7251,N_3283,N_998);
nand U7252 (N_7252,N_4033,N_759);
nand U7253 (N_7253,N_3755,N_2237);
nand U7254 (N_7254,N_2140,N_4466);
xor U7255 (N_7255,N_3494,N_4676);
nand U7256 (N_7256,N_1636,N_693);
and U7257 (N_7257,N_3805,N_1783);
xnor U7258 (N_7258,N_4717,N_576);
xnor U7259 (N_7259,N_1509,N_2120);
and U7260 (N_7260,N_2226,N_4424);
and U7261 (N_7261,N_4746,N_2626);
nand U7262 (N_7262,N_3606,N_4631);
nor U7263 (N_7263,N_1467,N_741);
xnor U7264 (N_7264,N_3031,N_1898);
nand U7265 (N_7265,N_390,N_2753);
and U7266 (N_7266,N_2535,N_3138);
nor U7267 (N_7267,N_710,N_1206);
and U7268 (N_7268,N_3210,N_2262);
nand U7269 (N_7269,N_1833,N_4947);
xnor U7270 (N_7270,N_733,N_1296);
nor U7271 (N_7271,N_2275,N_4523);
nand U7272 (N_7272,N_3523,N_561);
and U7273 (N_7273,N_1007,N_75);
xor U7274 (N_7274,N_1917,N_1346);
or U7275 (N_7275,N_2087,N_3712);
nor U7276 (N_7276,N_2337,N_2571);
xor U7277 (N_7277,N_610,N_726);
xor U7278 (N_7278,N_4357,N_1601);
xor U7279 (N_7279,N_3456,N_2363);
nor U7280 (N_7280,N_113,N_4467);
nand U7281 (N_7281,N_3623,N_2227);
nor U7282 (N_7282,N_1238,N_2314);
nor U7283 (N_7283,N_4866,N_2635);
and U7284 (N_7284,N_831,N_4501);
nor U7285 (N_7285,N_1797,N_660);
nand U7286 (N_7286,N_924,N_4982);
or U7287 (N_7287,N_832,N_3439);
xor U7288 (N_7288,N_4072,N_2469);
nor U7289 (N_7289,N_2023,N_3331);
xnor U7290 (N_7290,N_3599,N_4566);
nor U7291 (N_7291,N_2217,N_3422);
nor U7292 (N_7292,N_985,N_3546);
or U7293 (N_7293,N_518,N_4838);
nor U7294 (N_7294,N_1490,N_1962);
xor U7295 (N_7295,N_4723,N_176);
nor U7296 (N_7296,N_3543,N_2254);
nor U7297 (N_7297,N_400,N_3188);
nor U7298 (N_7298,N_1663,N_4938);
nand U7299 (N_7299,N_875,N_1092);
nor U7300 (N_7300,N_2411,N_4174);
xor U7301 (N_7301,N_572,N_1090);
or U7302 (N_7302,N_3704,N_2179);
or U7303 (N_7303,N_2552,N_1910);
nor U7304 (N_7304,N_3640,N_691);
nor U7305 (N_7305,N_2484,N_3024);
or U7306 (N_7306,N_4893,N_1446);
nand U7307 (N_7307,N_525,N_1298);
and U7308 (N_7308,N_1748,N_2006);
xnor U7309 (N_7309,N_3498,N_1113);
nand U7310 (N_7310,N_4040,N_420);
and U7311 (N_7311,N_4765,N_3045);
and U7312 (N_7312,N_462,N_4940);
nor U7313 (N_7313,N_3298,N_1067);
nor U7314 (N_7314,N_1914,N_2191);
nor U7315 (N_7315,N_1488,N_1868);
or U7316 (N_7316,N_3488,N_3239);
xnor U7317 (N_7317,N_719,N_195);
xnor U7318 (N_7318,N_492,N_2664);
and U7319 (N_7319,N_4775,N_2162);
xor U7320 (N_7320,N_3894,N_2840);
nor U7321 (N_7321,N_2066,N_1960);
xnor U7322 (N_7322,N_4063,N_2654);
xor U7323 (N_7323,N_3509,N_1343);
nor U7324 (N_7324,N_636,N_3684);
xor U7325 (N_7325,N_4123,N_3876);
nor U7326 (N_7326,N_2797,N_1274);
or U7327 (N_7327,N_2313,N_3573);
or U7328 (N_7328,N_2340,N_3504);
nor U7329 (N_7329,N_1231,N_1560);
xor U7330 (N_7330,N_962,N_2784);
nor U7331 (N_7331,N_3725,N_2074);
nor U7332 (N_7332,N_2398,N_1114);
and U7333 (N_7333,N_2458,N_698);
xnor U7334 (N_7334,N_4629,N_3968);
nor U7335 (N_7335,N_3205,N_3462);
nand U7336 (N_7336,N_1564,N_2584);
xnor U7337 (N_7337,N_2243,N_1563);
xnor U7338 (N_7338,N_558,N_386);
xnor U7339 (N_7339,N_2586,N_37);
or U7340 (N_7340,N_1890,N_266);
and U7341 (N_7341,N_1074,N_3369);
or U7342 (N_7342,N_2319,N_615);
and U7343 (N_7343,N_4181,N_1638);
xnor U7344 (N_7344,N_1422,N_1846);
nand U7345 (N_7345,N_2725,N_2921);
nor U7346 (N_7346,N_4682,N_1495);
xor U7347 (N_7347,N_2069,N_3885);
and U7348 (N_7348,N_481,N_3656);
and U7349 (N_7349,N_1165,N_3140);
xor U7350 (N_7350,N_4118,N_2719);
nor U7351 (N_7351,N_1184,N_3587);
nand U7352 (N_7352,N_4651,N_3154);
nand U7353 (N_7353,N_181,N_950);
nand U7354 (N_7354,N_3141,N_1265);
nor U7355 (N_7355,N_156,N_412);
nor U7356 (N_7356,N_341,N_3779);
nor U7357 (N_7357,N_3204,N_1907);
and U7358 (N_7358,N_4613,N_711);
and U7359 (N_7359,N_896,N_2962);
or U7360 (N_7360,N_3293,N_713);
and U7361 (N_7361,N_3258,N_1934);
nand U7362 (N_7362,N_2146,N_1145);
nor U7363 (N_7363,N_3179,N_1442);
or U7364 (N_7364,N_3350,N_4276);
and U7365 (N_7365,N_1166,N_2167);
nor U7366 (N_7366,N_3724,N_4437);
nand U7367 (N_7367,N_725,N_535);
xor U7368 (N_7368,N_4089,N_1901);
or U7369 (N_7369,N_2456,N_1086);
nor U7370 (N_7370,N_2017,N_4471);
xnor U7371 (N_7371,N_3054,N_144);
xor U7372 (N_7372,N_2874,N_1235);
nand U7373 (N_7373,N_3235,N_1789);
and U7374 (N_7374,N_304,N_677);
and U7375 (N_7375,N_4043,N_82);
nand U7376 (N_7376,N_2774,N_1696);
nand U7377 (N_7377,N_4062,N_1883);
or U7378 (N_7378,N_3255,N_2600);
and U7379 (N_7379,N_748,N_4178);
and U7380 (N_7380,N_1947,N_1046);
or U7381 (N_7381,N_786,N_2566);
nand U7382 (N_7382,N_1896,N_1525);
or U7383 (N_7383,N_175,N_1471);
xor U7384 (N_7384,N_2967,N_4109);
and U7385 (N_7385,N_3562,N_1735);
xor U7386 (N_7386,N_580,N_3320);
and U7387 (N_7387,N_4511,N_90);
nor U7388 (N_7388,N_3649,N_940);
or U7389 (N_7389,N_17,N_1295);
and U7390 (N_7390,N_2185,N_4602);
and U7391 (N_7391,N_380,N_4597);
xnor U7392 (N_7392,N_3480,N_4361);
or U7393 (N_7393,N_4305,N_4295);
and U7394 (N_7394,N_3848,N_277);
and U7395 (N_7395,N_2261,N_1710);
and U7396 (N_7396,N_190,N_3222);
nor U7397 (N_7397,N_2619,N_794);
nand U7398 (N_7398,N_2175,N_169);
nand U7399 (N_7399,N_1634,N_450);
and U7400 (N_7400,N_2299,N_1597);
nor U7401 (N_7401,N_9,N_4149);
nor U7402 (N_7402,N_4534,N_3404);
nor U7403 (N_7403,N_4531,N_2022);
nor U7404 (N_7404,N_1918,N_3815);
xnor U7405 (N_7405,N_3165,N_2762);
or U7406 (N_7406,N_2419,N_718);
or U7407 (N_7407,N_1887,N_4100);
xnor U7408 (N_7408,N_2263,N_2149);
xor U7409 (N_7409,N_4454,N_4645);
nor U7410 (N_7410,N_3048,N_1853);
or U7411 (N_7411,N_777,N_958);
nor U7412 (N_7412,N_3826,N_3387);
nor U7413 (N_7413,N_490,N_2830);
nand U7414 (N_7414,N_3737,N_2939);
nand U7415 (N_7415,N_2289,N_2200);
nor U7416 (N_7416,N_1550,N_4198);
or U7417 (N_7417,N_1585,N_3903);
nor U7418 (N_7418,N_4928,N_439);
nor U7419 (N_7419,N_1213,N_1246);
nor U7420 (N_7420,N_1157,N_1125);
xor U7421 (N_7421,N_3160,N_213);
and U7422 (N_7422,N_4910,N_2629);
xor U7423 (N_7423,N_3788,N_2201);
and U7424 (N_7424,N_1731,N_2482);
nor U7425 (N_7425,N_3247,N_4353);
and U7426 (N_7426,N_458,N_2029);
nor U7427 (N_7427,N_1581,N_4167);
or U7428 (N_7428,N_1790,N_391);
nand U7429 (N_7429,N_4635,N_2176);
or U7430 (N_7430,N_3478,N_3663);
nand U7431 (N_7431,N_3865,N_4343);
and U7432 (N_7432,N_4097,N_1537);
and U7433 (N_7433,N_2532,N_650);
and U7434 (N_7434,N_1734,N_4590);
nand U7435 (N_7435,N_2977,N_2911);
nor U7436 (N_7436,N_1650,N_3351);
xor U7437 (N_7437,N_3726,N_66);
and U7438 (N_7438,N_3842,N_3802);
and U7439 (N_7439,N_2413,N_486);
nor U7440 (N_7440,N_4839,N_2148);
xnor U7441 (N_7441,N_4013,N_3363);
and U7442 (N_7442,N_4959,N_1158);
xnor U7443 (N_7443,N_1306,N_707);
or U7444 (N_7444,N_3334,N_4503);
nand U7445 (N_7445,N_907,N_4407);
or U7446 (N_7446,N_4232,N_145);
nor U7447 (N_7447,N_1903,N_1470);
or U7448 (N_7448,N_2135,N_449);
nand U7449 (N_7449,N_3389,N_3776);
or U7450 (N_7450,N_441,N_666);
xnor U7451 (N_7451,N_1375,N_789);
or U7452 (N_7452,N_2317,N_1320);
and U7453 (N_7453,N_3396,N_3386);
and U7454 (N_7454,N_994,N_1974);
or U7455 (N_7455,N_345,N_3394);
or U7456 (N_7456,N_1469,N_740);
and U7457 (N_7457,N_2108,N_3440);
and U7458 (N_7458,N_298,N_4076);
xnor U7459 (N_7459,N_3414,N_1255);
or U7460 (N_7460,N_3731,N_612);
or U7461 (N_7461,N_4151,N_2033);
or U7462 (N_7462,N_487,N_3418);
or U7463 (N_7463,N_3413,N_1003);
xor U7464 (N_7464,N_4034,N_2883);
nand U7465 (N_7465,N_4494,N_1651);
nor U7466 (N_7466,N_1847,N_623);
nand U7467 (N_7467,N_136,N_353);
nand U7468 (N_7468,N_1949,N_4848);
xnor U7469 (N_7469,N_4715,N_2867);
and U7470 (N_7470,N_202,N_3395);
nand U7471 (N_7471,N_3050,N_1813);
xor U7472 (N_7472,N_1617,N_2837);
and U7473 (N_7473,N_3507,N_2803);
xnor U7474 (N_7474,N_1205,N_4958);
or U7475 (N_7475,N_4770,N_2310);
nor U7476 (N_7476,N_3859,N_41);
and U7477 (N_7477,N_3808,N_3740);
xor U7478 (N_7478,N_4753,N_3465);
nand U7479 (N_7479,N_3151,N_1996);
xnor U7480 (N_7480,N_335,N_1369);
or U7481 (N_7481,N_4008,N_575);
and U7482 (N_7482,N_2856,N_991);
xor U7483 (N_7483,N_366,N_2089);
and U7484 (N_7484,N_4382,N_625);
nand U7485 (N_7485,N_4771,N_1196);
nand U7486 (N_7486,N_2204,N_3371);
or U7487 (N_7487,N_3741,N_4260);
xnor U7488 (N_7488,N_3882,N_243);
and U7489 (N_7489,N_1822,N_2021);
and U7490 (N_7490,N_1885,N_4282);
or U7491 (N_7491,N_245,N_3534);
and U7492 (N_7492,N_1211,N_4859);
nand U7493 (N_7493,N_4229,N_1218);
nand U7494 (N_7494,N_2057,N_4593);
xnor U7495 (N_7495,N_221,N_149);
nor U7496 (N_7496,N_248,N_3036);
or U7497 (N_7497,N_534,N_1725);
xor U7498 (N_7498,N_1985,N_1762);
or U7499 (N_7499,N_1275,N_4055);
and U7500 (N_7500,N_1195,N_521);
nor U7501 (N_7501,N_644,N_4305);
nand U7502 (N_7502,N_2845,N_1753);
nand U7503 (N_7503,N_2429,N_1291);
or U7504 (N_7504,N_3292,N_3085);
nand U7505 (N_7505,N_3227,N_4665);
xnor U7506 (N_7506,N_3861,N_4207);
and U7507 (N_7507,N_1574,N_3828);
xor U7508 (N_7508,N_1100,N_681);
nand U7509 (N_7509,N_1587,N_1237);
and U7510 (N_7510,N_1400,N_4043);
or U7511 (N_7511,N_2491,N_4608);
and U7512 (N_7512,N_4011,N_4735);
nand U7513 (N_7513,N_4603,N_4926);
or U7514 (N_7514,N_4133,N_69);
and U7515 (N_7515,N_2105,N_682);
nand U7516 (N_7516,N_3366,N_3905);
nor U7517 (N_7517,N_3927,N_3599);
xnor U7518 (N_7518,N_4465,N_1041);
nand U7519 (N_7519,N_1345,N_2288);
xnor U7520 (N_7520,N_159,N_776);
nor U7521 (N_7521,N_1891,N_2153);
or U7522 (N_7522,N_4045,N_3546);
nor U7523 (N_7523,N_2023,N_3845);
nand U7524 (N_7524,N_4442,N_1654);
nand U7525 (N_7525,N_3345,N_1693);
and U7526 (N_7526,N_2126,N_1816);
and U7527 (N_7527,N_239,N_1439);
nor U7528 (N_7528,N_3566,N_2370);
or U7529 (N_7529,N_2164,N_118);
nand U7530 (N_7530,N_3261,N_933);
nor U7531 (N_7531,N_1004,N_3814);
xnor U7532 (N_7532,N_786,N_4675);
or U7533 (N_7533,N_731,N_885);
xor U7534 (N_7534,N_3766,N_2719);
or U7535 (N_7535,N_1420,N_328);
or U7536 (N_7536,N_945,N_4301);
nor U7537 (N_7537,N_3614,N_4567);
xor U7538 (N_7538,N_1929,N_4799);
and U7539 (N_7539,N_3297,N_2483);
and U7540 (N_7540,N_3245,N_2883);
xnor U7541 (N_7541,N_702,N_1821);
or U7542 (N_7542,N_3832,N_4721);
or U7543 (N_7543,N_958,N_2211);
xnor U7544 (N_7544,N_2448,N_1390);
and U7545 (N_7545,N_2435,N_3816);
or U7546 (N_7546,N_3544,N_2347);
and U7547 (N_7547,N_2106,N_3120);
nor U7548 (N_7548,N_1270,N_2351);
nor U7549 (N_7549,N_894,N_2092);
nor U7550 (N_7550,N_1,N_4366);
nand U7551 (N_7551,N_2037,N_4313);
nand U7552 (N_7552,N_2713,N_2984);
xor U7553 (N_7553,N_2955,N_124);
or U7554 (N_7554,N_4324,N_2938);
nor U7555 (N_7555,N_1873,N_2393);
nor U7556 (N_7556,N_2878,N_1240);
nand U7557 (N_7557,N_451,N_3645);
or U7558 (N_7558,N_1392,N_939);
nand U7559 (N_7559,N_3367,N_3210);
or U7560 (N_7560,N_3480,N_3983);
or U7561 (N_7561,N_2417,N_3880);
nand U7562 (N_7562,N_2392,N_1150);
nor U7563 (N_7563,N_279,N_4569);
and U7564 (N_7564,N_1291,N_4047);
nor U7565 (N_7565,N_2321,N_1997);
nand U7566 (N_7566,N_2799,N_3131);
nor U7567 (N_7567,N_4689,N_435);
nand U7568 (N_7568,N_3208,N_1168);
xnor U7569 (N_7569,N_1007,N_3718);
xnor U7570 (N_7570,N_4422,N_4319);
nor U7571 (N_7571,N_4873,N_4341);
nand U7572 (N_7572,N_389,N_284);
and U7573 (N_7573,N_3713,N_4590);
nand U7574 (N_7574,N_3793,N_4392);
and U7575 (N_7575,N_2549,N_1205);
nand U7576 (N_7576,N_89,N_3128);
nor U7577 (N_7577,N_4345,N_1528);
or U7578 (N_7578,N_250,N_4575);
nand U7579 (N_7579,N_4139,N_784);
nor U7580 (N_7580,N_4520,N_641);
and U7581 (N_7581,N_4767,N_4930);
or U7582 (N_7582,N_2245,N_3470);
xor U7583 (N_7583,N_3573,N_948);
xnor U7584 (N_7584,N_1016,N_1974);
nand U7585 (N_7585,N_4817,N_4369);
nand U7586 (N_7586,N_2298,N_1751);
and U7587 (N_7587,N_4731,N_4409);
xor U7588 (N_7588,N_1490,N_1807);
xor U7589 (N_7589,N_41,N_2278);
nor U7590 (N_7590,N_3573,N_3115);
or U7591 (N_7591,N_1924,N_2910);
and U7592 (N_7592,N_3776,N_474);
nand U7593 (N_7593,N_1936,N_2144);
xnor U7594 (N_7594,N_3730,N_2560);
xnor U7595 (N_7595,N_3279,N_134);
and U7596 (N_7596,N_2005,N_2821);
nand U7597 (N_7597,N_1199,N_2415);
nor U7598 (N_7598,N_1360,N_4615);
nor U7599 (N_7599,N_1175,N_168);
or U7600 (N_7600,N_789,N_2709);
nand U7601 (N_7601,N_1886,N_3888);
xor U7602 (N_7602,N_2077,N_2117);
or U7603 (N_7603,N_3187,N_1903);
nor U7604 (N_7604,N_1476,N_2302);
or U7605 (N_7605,N_4327,N_1683);
and U7606 (N_7606,N_4088,N_3800);
and U7607 (N_7607,N_4054,N_1505);
xnor U7608 (N_7608,N_4148,N_3191);
or U7609 (N_7609,N_1106,N_2019);
nor U7610 (N_7610,N_3959,N_2335);
nand U7611 (N_7611,N_953,N_2271);
or U7612 (N_7612,N_1316,N_1195);
or U7613 (N_7613,N_4295,N_4187);
nor U7614 (N_7614,N_2478,N_1848);
or U7615 (N_7615,N_3356,N_2143);
nor U7616 (N_7616,N_818,N_2034);
nand U7617 (N_7617,N_1154,N_4713);
nor U7618 (N_7618,N_4098,N_3209);
nand U7619 (N_7619,N_1793,N_4220);
nand U7620 (N_7620,N_2808,N_302);
or U7621 (N_7621,N_2385,N_2717);
nand U7622 (N_7622,N_4311,N_2027);
and U7623 (N_7623,N_157,N_2755);
nor U7624 (N_7624,N_2786,N_150);
nand U7625 (N_7625,N_2570,N_4347);
xor U7626 (N_7626,N_4973,N_3821);
nand U7627 (N_7627,N_555,N_3824);
nand U7628 (N_7628,N_4657,N_952);
nor U7629 (N_7629,N_649,N_1273);
or U7630 (N_7630,N_1717,N_3106);
nor U7631 (N_7631,N_4648,N_3787);
xor U7632 (N_7632,N_847,N_805);
nand U7633 (N_7633,N_1859,N_3498);
nor U7634 (N_7634,N_1624,N_4618);
nor U7635 (N_7635,N_2219,N_148);
and U7636 (N_7636,N_434,N_2021);
nor U7637 (N_7637,N_3216,N_3653);
xnor U7638 (N_7638,N_39,N_113);
nand U7639 (N_7639,N_219,N_3109);
nor U7640 (N_7640,N_3229,N_291);
xor U7641 (N_7641,N_3960,N_4292);
nand U7642 (N_7642,N_2613,N_3678);
or U7643 (N_7643,N_2978,N_1350);
or U7644 (N_7644,N_4174,N_381);
nand U7645 (N_7645,N_56,N_2570);
nand U7646 (N_7646,N_3028,N_2794);
nor U7647 (N_7647,N_4380,N_2865);
and U7648 (N_7648,N_901,N_120);
and U7649 (N_7649,N_1825,N_2643);
nor U7650 (N_7650,N_2254,N_1596);
or U7651 (N_7651,N_4670,N_1712);
nor U7652 (N_7652,N_3206,N_25);
or U7653 (N_7653,N_2773,N_1028);
xor U7654 (N_7654,N_1517,N_63);
nand U7655 (N_7655,N_4705,N_4558);
nor U7656 (N_7656,N_4670,N_966);
xnor U7657 (N_7657,N_3897,N_380);
or U7658 (N_7658,N_3993,N_1396);
nand U7659 (N_7659,N_4888,N_4090);
nor U7660 (N_7660,N_3844,N_4884);
xor U7661 (N_7661,N_4191,N_4649);
xor U7662 (N_7662,N_2904,N_2466);
and U7663 (N_7663,N_472,N_2905);
nand U7664 (N_7664,N_3137,N_985);
nand U7665 (N_7665,N_3562,N_3381);
and U7666 (N_7666,N_2123,N_1996);
or U7667 (N_7667,N_4378,N_1742);
nor U7668 (N_7668,N_1763,N_345);
xnor U7669 (N_7669,N_4137,N_4970);
and U7670 (N_7670,N_42,N_741);
nor U7671 (N_7671,N_1610,N_1878);
xor U7672 (N_7672,N_2140,N_384);
nor U7673 (N_7673,N_1679,N_2606);
nor U7674 (N_7674,N_2214,N_2624);
and U7675 (N_7675,N_1933,N_2160);
or U7676 (N_7676,N_1240,N_1009);
nor U7677 (N_7677,N_1518,N_2158);
and U7678 (N_7678,N_287,N_1818);
xor U7679 (N_7679,N_4587,N_1435);
nor U7680 (N_7680,N_1478,N_1663);
xnor U7681 (N_7681,N_738,N_1962);
nor U7682 (N_7682,N_2883,N_1597);
or U7683 (N_7683,N_4758,N_1465);
nor U7684 (N_7684,N_419,N_2801);
or U7685 (N_7685,N_1833,N_3152);
xor U7686 (N_7686,N_465,N_952);
xnor U7687 (N_7687,N_4954,N_1939);
nand U7688 (N_7688,N_2314,N_3313);
nand U7689 (N_7689,N_1487,N_4605);
and U7690 (N_7690,N_70,N_3218);
nand U7691 (N_7691,N_4661,N_3796);
or U7692 (N_7692,N_4482,N_3006);
xor U7693 (N_7693,N_786,N_953);
and U7694 (N_7694,N_4590,N_4768);
nand U7695 (N_7695,N_3112,N_624);
and U7696 (N_7696,N_4962,N_3644);
and U7697 (N_7697,N_4007,N_850);
xor U7698 (N_7698,N_1693,N_1785);
and U7699 (N_7699,N_2172,N_459);
and U7700 (N_7700,N_1353,N_4437);
nor U7701 (N_7701,N_6,N_573);
and U7702 (N_7702,N_3528,N_1248);
nor U7703 (N_7703,N_1359,N_806);
nor U7704 (N_7704,N_1553,N_2646);
or U7705 (N_7705,N_3366,N_1597);
nor U7706 (N_7706,N_1791,N_1698);
nand U7707 (N_7707,N_1612,N_2332);
or U7708 (N_7708,N_3792,N_2272);
nor U7709 (N_7709,N_4030,N_1917);
and U7710 (N_7710,N_2689,N_213);
xnor U7711 (N_7711,N_2858,N_2385);
xnor U7712 (N_7712,N_1628,N_4557);
and U7713 (N_7713,N_541,N_1217);
or U7714 (N_7714,N_3375,N_1170);
or U7715 (N_7715,N_4390,N_1821);
or U7716 (N_7716,N_3448,N_980);
and U7717 (N_7717,N_3473,N_267);
nand U7718 (N_7718,N_952,N_1171);
nand U7719 (N_7719,N_1569,N_2111);
nor U7720 (N_7720,N_1736,N_897);
xor U7721 (N_7721,N_712,N_4020);
or U7722 (N_7722,N_988,N_4416);
nand U7723 (N_7723,N_4605,N_2824);
nand U7724 (N_7724,N_2632,N_1719);
and U7725 (N_7725,N_4863,N_3542);
nand U7726 (N_7726,N_1952,N_2155);
nand U7727 (N_7727,N_3854,N_4542);
and U7728 (N_7728,N_2665,N_4717);
nor U7729 (N_7729,N_2157,N_519);
nor U7730 (N_7730,N_1074,N_3250);
and U7731 (N_7731,N_4392,N_1480);
nor U7732 (N_7732,N_1845,N_2857);
nor U7733 (N_7733,N_3248,N_3874);
xor U7734 (N_7734,N_2223,N_2416);
or U7735 (N_7735,N_444,N_4769);
nand U7736 (N_7736,N_3559,N_2327);
nand U7737 (N_7737,N_1483,N_3656);
xnor U7738 (N_7738,N_2275,N_4417);
xnor U7739 (N_7739,N_4455,N_2870);
or U7740 (N_7740,N_1555,N_4884);
or U7741 (N_7741,N_951,N_1224);
nor U7742 (N_7742,N_1390,N_2543);
nor U7743 (N_7743,N_1953,N_535);
nand U7744 (N_7744,N_1416,N_3269);
or U7745 (N_7745,N_4675,N_1024);
nand U7746 (N_7746,N_3887,N_450);
nand U7747 (N_7747,N_709,N_3115);
or U7748 (N_7748,N_1829,N_3777);
nor U7749 (N_7749,N_131,N_2614);
or U7750 (N_7750,N_3106,N_3664);
xor U7751 (N_7751,N_2494,N_834);
or U7752 (N_7752,N_3704,N_587);
or U7753 (N_7753,N_3522,N_31);
nor U7754 (N_7754,N_420,N_3324);
and U7755 (N_7755,N_1832,N_1239);
xor U7756 (N_7756,N_2070,N_3082);
nor U7757 (N_7757,N_2864,N_1747);
nand U7758 (N_7758,N_21,N_1461);
and U7759 (N_7759,N_1548,N_2553);
nor U7760 (N_7760,N_45,N_986);
nand U7761 (N_7761,N_2935,N_2828);
nor U7762 (N_7762,N_3223,N_1953);
and U7763 (N_7763,N_1055,N_2233);
xor U7764 (N_7764,N_329,N_3067);
and U7765 (N_7765,N_1483,N_2571);
nor U7766 (N_7766,N_4492,N_4851);
nor U7767 (N_7767,N_1228,N_1654);
and U7768 (N_7768,N_2491,N_4213);
xor U7769 (N_7769,N_3668,N_262);
and U7770 (N_7770,N_2625,N_641);
and U7771 (N_7771,N_988,N_2957);
and U7772 (N_7772,N_2486,N_3510);
xnor U7773 (N_7773,N_452,N_3656);
and U7774 (N_7774,N_3635,N_4113);
and U7775 (N_7775,N_3055,N_2557);
and U7776 (N_7776,N_3789,N_1505);
nor U7777 (N_7777,N_719,N_3263);
or U7778 (N_7778,N_3695,N_266);
nand U7779 (N_7779,N_2672,N_1563);
nor U7780 (N_7780,N_3528,N_1968);
nand U7781 (N_7781,N_475,N_2043);
xnor U7782 (N_7782,N_186,N_4022);
xnor U7783 (N_7783,N_3291,N_733);
or U7784 (N_7784,N_3513,N_1251);
xnor U7785 (N_7785,N_2657,N_2845);
xnor U7786 (N_7786,N_3140,N_4027);
and U7787 (N_7787,N_4862,N_537);
and U7788 (N_7788,N_420,N_2000);
and U7789 (N_7789,N_109,N_1638);
nand U7790 (N_7790,N_2371,N_1519);
and U7791 (N_7791,N_4921,N_2730);
or U7792 (N_7792,N_3580,N_4374);
and U7793 (N_7793,N_2352,N_1349);
nand U7794 (N_7794,N_4313,N_2885);
and U7795 (N_7795,N_77,N_4255);
nand U7796 (N_7796,N_480,N_2358);
or U7797 (N_7797,N_618,N_532);
xnor U7798 (N_7798,N_2055,N_48);
and U7799 (N_7799,N_2191,N_3827);
nor U7800 (N_7800,N_2360,N_1477);
and U7801 (N_7801,N_1755,N_1984);
and U7802 (N_7802,N_185,N_3991);
nand U7803 (N_7803,N_434,N_4402);
xnor U7804 (N_7804,N_1032,N_865);
nand U7805 (N_7805,N_1613,N_3563);
or U7806 (N_7806,N_1293,N_399);
and U7807 (N_7807,N_3991,N_4659);
nor U7808 (N_7808,N_4116,N_2792);
xnor U7809 (N_7809,N_594,N_3325);
nor U7810 (N_7810,N_1157,N_2300);
nand U7811 (N_7811,N_705,N_1149);
or U7812 (N_7812,N_2907,N_1625);
xor U7813 (N_7813,N_3750,N_3429);
or U7814 (N_7814,N_544,N_1127);
or U7815 (N_7815,N_4712,N_3771);
and U7816 (N_7816,N_2282,N_3248);
nor U7817 (N_7817,N_3749,N_4831);
nor U7818 (N_7818,N_4859,N_3321);
nor U7819 (N_7819,N_39,N_4093);
and U7820 (N_7820,N_2869,N_4026);
or U7821 (N_7821,N_4741,N_489);
xor U7822 (N_7822,N_109,N_3235);
nand U7823 (N_7823,N_1628,N_3242);
xor U7824 (N_7824,N_2042,N_1944);
xnor U7825 (N_7825,N_1759,N_122);
nor U7826 (N_7826,N_914,N_2690);
and U7827 (N_7827,N_4508,N_2695);
and U7828 (N_7828,N_3468,N_499);
and U7829 (N_7829,N_2645,N_4965);
nor U7830 (N_7830,N_2507,N_2180);
and U7831 (N_7831,N_2655,N_2898);
nand U7832 (N_7832,N_1448,N_3704);
and U7833 (N_7833,N_4,N_156);
and U7834 (N_7834,N_2710,N_4943);
and U7835 (N_7835,N_3361,N_3853);
and U7836 (N_7836,N_179,N_3007);
xor U7837 (N_7837,N_471,N_4949);
nand U7838 (N_7838,N_576,N_1322);
or U7839 (N_7839,N_203,N_1701);
nor U7840 (N_7840,N_4609,N_460);
or U7841 (N_7841,N_988,N_3919);
or U7842 (N_7842,N_2538,N_1528);
xor U7843 (N_7843,N_3739,N_4655);
nor U7844 (N_7844,N_1271,N_3713);
nand U7845 (N_7845,N_3734,N_1102);
and U7846 (N_7846,N_638,N_4495);
and U7847 (N_7847,N_311,N_4426);
and U7848 (N_7848,N_2152,N_3677);
nor U7849 (N_7849,N_4936,N_4477);
or U7850 (N_7850,N_2287,N_232);
nor U7851 (N_7851,N_4556,N_4583);
and U7852 (N_7852,N_3595,N_3798);
nand U7853 (N_7853,N_1182,N_825);
or U7854 (N_7854,N_4381,N_2199);
and U7855 (N_7855,N_2373,N_1611);
or U7856 (N_7856,N_347,N_4350);
xor U7857 (N_7857,N_1257,N_1682);
xnor U7858 (N_7858,N_3909,N_2956);
or U7859 (N_7859,N_2678,N_2743);
and U7860 (N_7860,N_1265,N_1850);
and U7861 (N_7861,N_1800,N_4289);
and U7862 (N_7862,N_4959,N_2036);
xor U7863 (N_7863,N_3868,N_4528);
nand U7864 (N_7864,N_2574,N_2891);
nor U7865 (N_7865,N_4775,N_1428);
nor U7866 (N_7866,N_2394,N_3546);
nand U7867 (N_7867,N_1701,N_3380);
or U7868 (N_7868,N_3989,N_3858);
or U7869 (N_7869,N_4270,N_1236);
nand U7870 (N_7870,N_1436,N_288);
nand U7871 (N_7871,N_4764,N_364);
nand U7872 (N_7872,N_3947,N_4116);
xnor U7873 (N_7873,N_4218,N_325);
or U7874 (N_7874,N_4360,N_3137);
nand U7875 (N_7875,N_3023,N_3567);
nand U7876 (N_7876,N_4980,N_3013);
and U7877 (N_7877,N_4423,N_4115);
xor U7878 (N_7878,N_297,N_4407);
nand U7879 (N_7879,N_2660,N_4779);
or U7880 (N_7880,N_3720,N_3641);
xnor U7881 (N_7881,N_243,N_3757);
or U7882 (N_7882,N_4198,N_4428);
and U7883 (N_7883,N_3745,N_3193);
nor U7884 (N_7884,N_3948,N_2480);
nand U7885 (N_7885,N_1983,N_3965);
and U7886 (N_7886,N_4065,N_4637);
nor U7887 (N_7887,N_65,N_4709);
or U7888 (N_7888,N_785,N_953);
xnor U7889 (N_7889,N_1792,N_4628);
nand U7890 (N_7890,N_3179,N_4803);
or U7891 (N_7891,N_546,N_4521);
nor U7892 (N_7892,N_1277,N_4389);
or U7893 (N_7893,N_1116,N_672);
nand U7894 (N_7894,N_1951,N_3315);
nor U7895 (N_7895,N_4740,N_1921);
xor U7896 (N_7896,N_155,N_562);
and U7897 (N_7897,N_2186,N_3094);
and U7898 (N_7898,N_2577,N_2806);
or U7899 (N_7899,N_4797,N_2484);
nand U7900 (N_7900,N_3395,N_4814);
or U7901 (N_7901,N_110,N_324);
and U7902 (N_7902,N_2304,N_1897);
and U7903 (N_7903,N_3547,N_2618);
nor U7904 (N_7904,N_322,N_2801);
nor U7905 (N_7905,N_4911,N_117);
and U7906 (N_7906,N_285,N_1655);
nor U7907 (N_7907,N_1332,N_2245);
and U7908 (N_7908,N_1916,N_903);
or U7909 (N_7909,N_334,N_1309);
nor U7910 (N_7910,N_2733,N_4793);
nand U7911 (N_7911,N_4569,N_2578);
nor U7912 (N_7912,N_2306,N_1745);
xnor U7913 (N_7913,N_2606,N_2616);
and U7914 (N_7914,N_2357,N_2650);
nor U7915 (N_7915,N_674,N_2708);
nor U7916 (N_7916,N_1065,N_1214);
or U7917 (N_7917,N_1585,N_958);
xnor U7918 (N_7918,N_4483,N_3544);
or U7919 (N_7919,N_770,N_680);
nand U7920 (N_7920,N_376,N_4472);
or U7921 (N_7921,N_215,N_3174);
or U7922 (N_7922,N_390,N_1606);
or U7923 (N_7923,N_2108,N_396);
xor U7924 (N_7924,N_2769,N_4253);
nand U7925 (N_7925,N_3920,N_2728);
nor U7926 (N_7926,N_2206,N_610);
and U7927 (N_7927,N_2828,N_840);
nor U7928 (N_7928,N_3180,N_2400);
nand U7929 (N_7929,N_635,N_3889);
xnor U7930 (N_7930,N_1924,N_622);
and U7931 (N_7931,N_3180,N_1785);
xnor U7932 (N_7932,N_1628,N_1976);
nor U7933 (N_7933,N_1706,N_1947);
xor U7934 (N_7934,N_405,N_3880);
nand U7935 (N_7935,N_2019,N_3488);
nand U7936 (N_7936,N_2797,N_3788);
and U7937 (N_7937,N_1188,N_2208);
or U7938 (N_7938,N_3142,N_2337);
nor U7939 (N_7939,N_2476,N_4501);
xnor U7940 (N_7940,N_2851,N_2009);
and U7941 (N_7941,N_1052,N_4014);
xor U7942 (N_7942,N_1798,N_1359);
nand U7943 (N_7943,N_1685,N_3293);
or U7944 (N_7944,N_585,N_2383);
or U7945 (N_7945,N_1548,N_3420);
and U7946 (N_7946,N_120,N_4367);
xor U7947 (N_7947,N_1538,N_3984);
nand U7948 (N_7948,N_2043,N_2919);
xnor U7949 (N_7949,N_3557,N_1051);
and U7950 (N_7950,N_1695,N_1245);
and U7951 (N_7951,N_4588,N_2007);
nand U7952 (N_7952,N_220,N_146);
or U7953 (N_7953,N_2522,N_450);
nor U7954 (N_7954,N_1078,N_2634);
xor U7955 (N_7955,N_4898,N_3728);
and U7956 (N_7956,N_1960,N_1042);
or U7957 (N_7957,N_3524,N_4615);
or U7958 (N_7958,N_1746,N_3637);
or U7959 (N_7959,N_1190,N_1663);
nand U7960 (N_7960,N_2691,N_4974);
xor U7961 (N_7961,N_2529,N_1114);
and U7962 (N_7962,N_3763,N_4593);
and U7963 (N_7963,N_3070,N_3618);
and U7964 (N_7964,N_2041,N_4282);
nand U7965 (N_7965,N_3261,N_2399);
or U7966 (N_7966,N_942,N_395);
and U7967 (N_7967,N_2576,N_2748);
xnor U7968 (N_7968,N_618,N_1278);
xnor U7969 (N_7969,N_340,N_2798);
nand U7970 (N_7970,N_98,N_2620);
nor U7971 (N_7971,N_2239,N_4495);
xnor U7972 (N_7972,N_3714,N_1479);
xnor U7973 (N_7973,N_3576,N_4562);
nand U7974 (N_7974,N_3379,N_1607);
xnor U7975 (N_7975,N_2228,N_3793);
nor U7976 (N_7976,N_4461,N_4901);
and U7977 (N_7977,N_4436,N_2805);
nor U7978 (N_7978,N_4625,N_773);
and U7979 (N_7979,N_2204,N_1446);
nor U7980 (N_7980,N_683,N_299);
nor U7981 (N_7981,N_3943,N_3200);
and U7982 (N_7982,N_4897,N_2259);
nor U7983 (N_7983,N_2057,N_1178);
and U7984 (N_7984,N_176,N_468);
or U7985 (N_7985,N_3540,N_914);
nand U7986 (N_7986,N_4778,N_1082);
nor U7987 (N_7987,N_808,N_4024);
nand U7988 (N_7988,N_4132,N_2900);
nor U7989 (N_7989,N_1142,N_1976);
nor U7990 (N_7990,N_331,N_1535);
nand U7991 (N_7991,N_3180,N_3536);
nor U7992 (N_7992,N_3659,N_1615);
or U7993 (N_7993,N_3843,N_4586);
and U7994 (N_7994,N_3407,N_3386);
or U7995 (N_7995,N_1481,N_3425);
xor U7996 (N_7996,N_2093,N_4461);
nand U7997 (N_7997,N_1395,N_818);
and U7998 (N_7998,N_1596,N_2093);
or U7999 (N_7999,N_185,N_4728);
nand U8000 (N_8000,N_583,N_4636);
nor U8001 (N_8001,N_1335,N_1262);
and U8002 (N_8002,N_2600,N_1968);
xnor U8003 (N_8003,N_2470,N_3966);
and U8004 (N_8004,N_4275,N_853);
nand U8005 (N_8005,N_3922,N_3607);
or U8006 (N_8006,N_2347,N_2053);
nor U8007 (N_8007,N_77,N_4284);
and U8008 (N_8008,N_2150,N_28);
nand U8009 (N_8009,N_3836,N_4410);
nand U8010 (N_8010,N_811,N_904);
nor U8011 (N_8011,N_3680,N_2710);
nor U8012 (N_8012,N_3617,N_4968);
and U8013 (N_8013,N_1217,N_918);
nand U8014 (N_8014,N_4895,N_3769);
or U8015 (N_8015,N_3730,N_4201);
xor U8016 (N_8016,N_4211,N_254);
nand U8017 (N_8017,N_998,N_2496);
xnor U8018 (N_8018,N_501,N_4375);
or U8019 (N_8019,N_1593,N_2758);
xnor U8020 (N_8020,N_669,N_1817);
nor U8021 (N_8021,N_2830,N_102);
or U8022 (N_8022,N_4433,N_3880);
nor U8023 (N_8023,N_1167,N_2320);
or U8024 (N_8024,N_4152,N_4758);
or U8025 (N_8025,N_828,N_493);
or U8026 (N_8026,N_419,N_1840);
or U8027 (N_8027,N_1895,N_4069);
nor U8028 (N_8028,N_1042,N_3863);
and U8029 (N_8029,N_2964,N_1323);
nand U8030 (N_8030,N_2749,N_1762);
and U8031 (N_8031,N_1603,N_3845);
nand U8032 (N_8032,N_3630,N_766);
and U8033 (N_8033,N_4830,N_3015);
nand U8034 (N_8034,N_750,N_3016);
or U8035 (N_8035,N_1289,N_2282);
and U8036 (N_8036,N_1253,N_3509);
and U8037 (N_8037,N_2520,N_940);
nor U8038 (N_8038,N_3666,N_352);
nor U8039 (N_8039,N_1976,N_1564);
nand U8040 (N_8040,N_4438,N_1764);
nand U8041 (N_8041,N_3615,N_3188);
xor U8042 (N_8042,N_1001,N_215);
and U8043 (N_8043,N_3054,N_876);
nor U8044 (N_8044,N_4729,N_3432);
or U8045 (N_8045,N_3665,N_4265);
nand U8046 (N_8046,N_3762,N_410);
nand U8047 (N_8047,N_4129,N_82);
nor U8048 (N_8048,N_2868,N_4020);
or U8049 (N_8049,N_4552,N_3643);
or U8050 (N_8050,N_3523,N_806);
xor U8051 (N_8051,N_3694,N_332);
xnor U8052 (N_8052,N_1335,N_627);
xor U8053 (N_8053,N_3742,N_1562);
or U8054 (N_8054,N_4416,N_1848);
nand U8055 (N_8055,N_104,N_3944);
and U8056 (N_8056,N_883,N_4735);
nand U8057 (N_8057,N_4828,N_1702);
nand U8058 (N_8058,N_4949,N_3370);
and U8059 (N_8059,N_2301,N_313);
and U8060 (N_8060,N_1183,N_1817);
or U8061 (N_8061,N_2971,N_4201);
and U8062 (N_8062,N_2718,N_519);
and U8063 (N_8063,N_4411,N_883);
and U8064 (N_8064,N_3989,N_2425);
xor U8065 (N_8065,N_1600,N_3317);
nand U8066 (N_8066,N_4729,N_534);
and U8067 (N_8067,N_3494,N_3812);
nor U8068 (N_8068,N_2641,N_2991);
nor U8069 (N_8069,N_2267,N_1409);
or U8070 (N_8070,N_3157,N_4063);
xor U8071 (N_8071,N_1416,N_293);
nand U8072 (N_8072,N_3340,N_1407);
nand U8073 (N_8073,N_578,N_4969);
xnor U8074 (N_8074,N_3472,N_3276);
nand U8075 (N_8075,N_1907,N_1614);
or U8076 (N_8076,N_3719,N_4686);
nor U8077 (N_8077,N_3210,N_2367);
and U8078 (N_8078,N_2684,N_734);
nand U8079 (N_8079,N_25,N_1602);
or U8080 (N_8080,N_4840,N_4728);
and U8081 (N_8081,N_4831,N_955);
and U8082 (N_8082,N_4492,N_327);
xnor U8083 (N_8083,N_1036,N_466);
nand U8084 (N_8084,N_903,N_12);
nand U8085 (N_8085,N_4813,N_1692);
or U8086 (N_8086,N_4888,N_2112);
or U8087 (N_8087,N_504,N_2427);
nand U8088 (N_8088,N_2174,N_1247);
nor U8089 (N_8089,N_1544,N_1205);
nor U8090 (N_8090,N_647,N_1699);
and U8091 (N_8091,N_2160,N_1434);
nor U8092 (N_8092,N_4040,N_1603);
nor U8093 (N_8093,N_3830,N_2078);
nor U8094 (N_8094,N_1875,N_4545);
or U8095 (N_8095,N_642,N_1900);
or U8096 (N_8096,N_3483,N_1260);
or U8097 (N_8097,N_228,N_976);
nand U8098 (N_8098,N_3849,N_489);
nor U8099 (N_8099,N_1667,N_996);
nand U8100 (N_8100,N_240,N_214);
nor U8101 (N_8101,N_1850,N_1690);
or U8102 (N_8102,N_910,N_383);
nor U8103 (N_8103,N_3925,N_3954);
nor U8104 (N_8104,N_1235,N_1311);
and U8105 (N_8105,N_398,N_1568);
xnor U8106 (N_8106,N_1273,N_4378);
nor U8107 (N_8107,N_900,N_3116);
or U8108 (N_8108,N_3297,N_915);
nand U8109 (N_8109,N_3561,N_1894);
xnor U8110 (N_8110,N_2822,N_1803);
or U8111 (N_8111,N_4583,N_3311);
and U8112 (N_8112,N_1096,N_407);
or U8113 (N_8113,N_521,N_2798);
and U8114 (N_8114,N_4280,N_312);
nor U8115 (N_8115,N_89,N_2262);
nor U8116 (N_8116,N_4543,N_2835);
or U8117 (N_8117,N_2788,N_613);
nand U8118 (N_8118,N_3428,N_606);
nor U8119 (N_8119,N_3823,N_3407);
nand U8120 (N_8120,N_2604,N_222);
and U8121 (N_8121,N_3022,N_1121);
and U8122 (N_8122,N_752,N_1339);
nor U8123 (N_8123,N_3589,N_3683);
nand U8124 (N_8124,N_2148,N_386);
nor U8125 (N_8125,N_4003,N_1476);
nand U8126 (N_8126,N_1944,N_2860);
nor U8127 (N_8127,N_3064,N_2188);
xor U8128 (N_8128,N_4043,N_4696);
or U8129 (N_8129,N_4945,N_3588);
or U8130 (N_8130,N_1127,N_1388);
nor U8131 (N_8131,N_4386,N_4442);
or U8132 (N_8132,N_2569,N_1578);
or U8133 (N_8133,N_2925,N_3119);
nor U8134 (N_8134,N_1864,N_3484);
xor U8135 (N_8135,N_3065,N_690);
nor U8136 (N_8136,N_4403,N_1788);
nor U8137 (N_8137,N_4352,N_1951);
or U8138 (N_8138,N_3144,N_4962);
or U8139 (N_8139,N_2918,N_157);
nand U8140 (N_8140,N_2571,N_1696);
nor U8141 (N_8141,N_1279,N_4955);
xor U8142 (N_8142,N_2019,N_1430);
or U8143 (N_8143,N_4032,N_4159);
xnor U8144 (N_8144,N_966,N_738);
or U8145 (N_8145,N_4194,N_3574);
xor U8146 (N_8146,N_667,N_2833);
and U8147 (N_8147,N_4820,N_2670);
nor U8148 (N_8148,N_279,N_3696);
and U8149 (N_8149,N_1314,N_255);
nand U8150 (N_8150,N_549,N_182);
or U8151 (N_8151,N_3737,N_399);
xor U8152 (N_8152,N_2260,N_3080);
or U8153 (N_8153,N_2223,N_3178);
nor U8154 (N_8154,N_403,N_2637);
and U8155 (N_8155,N_935,N_2492);
xnor U8156 (N_8156,N_3784,N_3273);
or U8157 (N_8157,N_2041,N_360);
and U8158 (N_8158,N_2369,N_3761);
xor U8159 (N_8159,N_3629,N_4561);
nor U8160 (N_8160,N_2489,N_3772);
or U8161 (N_8161,N_1808,N_1729);
nand U8162 (N_8162,N_2610,N_557);
or U8163 (N_8163,N_575,N_4755);
nor U8164 (N_8164,N_3909,N_163);
nand U8165 (N_8165,N_2175,N_3600);
nand U8166 (N_8166,N_2252,N_3013);
and U8167 (N_8167,N_3315,N_703);
or U8168 (N_8168,N_626,N_2161);
nor U8169 (N_8169,N_2128,N_4087);
or U8170 (N_8170,N_1986,N_484);
xor U8171 (N_8171,N_2607,N_1150);
or U8172 (N_8172,N_2357,N_4917);
nand U8173 (N_8173,N_3908,N_2250);
and U8174 (N_8174,N_1168,N_809);
or U8175 (N_8175,N_3619,N_991);
nand U8176 (N_8176,N_2195,N_4193);
nor U8177 (N_8177,N_3478,N_359);
xnor U8178 (N_8178,N_3115,N_612);
nor U8179 (N_8179,N_3240,N_735);
xnor U8180 (N_8180,N_4141,N_359);
xor U8181 (N_8181,N_2909,N_1901);
or U8182 (N_8182,N_3476,N_1161);
or U8183 (N_8183,N_1298,N_3730);
xor U8184 (N_8184,N_498,N_4619);
nand U8185 (N_8185,N_4944,N_4915);
and U8186 (N_8186,N_4444,N_2794);
and U8187 (N_8187,N_1934,N_1410);
nand U8188 (N_8188,N_2669,N_387);
nand U8189 (N_8189,N_3775,N_615);
xor U8190 (N_8190,N_4927,N_3487);
nor U8191 (N_8191,N_2112,N_3035);
nand U8192 (N_8192,N_3338,N_528);
and U8193 (N_8193,N_4742,N_2617);
and U8194 (N_8194,N_4095,N_1595);
and U8195 (N_8195,N_2792,N_4059);
nor U8196 (N_8196,N_4838,N_785);
or U8197 (N_8197,N_814,N_1732);
or U8198 (N_8198,N_3260,N_4734);
or U8199 (N_8199,N_2585,N_129);
nor U8200 (N_8200,N_1842,N_3935);
or U8201 (N_8201,N_216,N_2042);
or U8202 (N_8202,N_1790,N_2961);
nor U8203 (N_8203,N_4594,N_2365);
nor U8204 (N_8204,N_1460,N_2505);
or U8205 (N_8205,N_1180,N_436);
nor U8206 (N_8206,N_2503,N_3700);
xor U8207 (N_8207,N_3065,N_81);
and U8208 (N_8208,N_3794,N_4944);
and U8209 (N_8209,N_1667,N_3566);
or U8210 (N_8210,N_2029,N_768);
nand U8211 (N_8211,N_491,N_671);
nand U8212 (N_8212,N_1982,N_4378);
and U8213 (N_8213,N_1132,N_1449);
nand U8214 (N_8214,N_3528,N_3730);
nand U8215 (N_8215,N_1815,N_2184);
xnor U8216 (N_8216,N_3964,N_4099);
and U8217 (N_8217,N_4399,N_1959);
nor U8218 (N_8218,N_1122,N_2050);
or U8219 (N_8219,N_1388,N_2687);
or U8220 (N_8220,N_2552,N_2443);
nand U8221 (N_8221,N_167,N_1161);
and U8222 (N_8222,N_2453,N_1712);
or U8223 (N_8223,N_88,N_4743);
xor U8224 (N_8224,N_443,N_4780);
or U8225 (N_8225,N_2219,N_4138);
nor U8226 (N_8226,N_4836,N_4147);
and U8227 (N_8227,N_4600,N_2062);
xnor U8228 (N_8228,N_3194,N_3271);
and U8229 (N_8229,N_1685,N_2212);
or U8230 (N_8230,N_4218,N_1692);
nand U8231 (N_8231,N_4204,N_1881);
or U8232 (N_8232,N_331,N_1823);
or U8233 (N_8233,N_808,N_4483);
and U8234 (N_8234,N_3536,N_2401);
or U8235 (N_8235,N_4434,N_4038);
and U8236 (N_8236,N_4372,N_359);
xnor U8237 (N_8237,N_1072,N_4754);
xor U8238 (N_8238,N_2932,N_204);
xnor U8239 (N_8239,N_111,N_2344);
or U8240 (N_8240,N_3954,N_373);
or U8241 (N_8241,N_151,N_1559);
or U8242 (N_8242,N_2253,N_1923);
or U8243 (N_8243,N_348,N_3747);
nor U8244 (N_8244,N_2126,N_1032);
or U8245 (N_8245,N_1358,N_2022);
nand U8246 (N_8246,N_4475,N_3618);
and U8247 (N_8247,N_2867,N_1260);
and U8248 (N_8248,N_4141,N_4024);
xnor U8249 (N_8249,N_4042,N_3511);
and U8250 (N_8250,N_3312,N_1453);
or U8251 (N_8251,N_230,N_2261);
nor U8252 (N_8252,N_1795,N_4060);
nor U8253 (N_8253,N_3039,N_1257);
nor U8254 (N_8254,N_825,N_2940);
or U8255 (N_8255,N_2521,N_3814);
xor U8256 (N_8256,N_3670,N_3283);
or U8257 (N_8257,N_674,N_4740);
nand U8258 (N_8258,N_294,N_747);
or U8259 (N_8259,N_2598,N_149);
or U8260 (N_8260,N_3232,N_1212);
nand U8261 (N_8261,N_3115,N_1837);
nor U8262 (N_8262,N_2383,N_3743);
and U8263 (N_8263,N_4818,N_4048);
or U8264 (N_8264,N_660,N_1032);
and U8265 (N_8265,N_3608,N_1969);
or U8266 (N_8266,N_1937,N_2514);
xnor U8267 (N_8267,N_2538,N_1485);
and U8268 (N_8268,N_1733,N_2280);
or U8269 (N_8269,N_1820,N_1142);
nand U8270 (N_8270,N_3609,N_1742);
or U8271 (N_8271,N_4876,N_3566);
xor U8272 (N_8272,N_3595,N_2549);
xnor U8273 (N_8273,N_1496,N_3848);
and U8274 (N_8274,N_860,N_4487);
nand U8275 (N_8275,N_504,N_186);
nand U8276 (N_8276,N_3999,N_3931);
and U8277 (N_8277,N_1098,N_3407);
and U8278 (N_8278,N_4695,N_3509);
or U8279 (N_8279,N_1525,N_2072);
or U8280 (N_8280,N_2144,N_4836);
nor U8281 (N_8281,N_3533,N_1843);
nor U8282 (N_8282,N_3905,N_4852);
xor U8283 (N_8283,N_2754,N_120);
nand U8284 (N_8284,N_4713,N_278);
and U8285 (N_8285,N_4192,N_4198);
nor U8286 (N_8286,N_3914,N_4683);
nor U8287 (N_8287,N_1652,N_615);
xnor U8288 (N_8288,N_2098,N_608);
and U8289 (N_8289,N_359,N_513);
nand U8290 (N_8290,N_627,N_4192);
and U8291 (N_8291,N_374,N_1606);
and U8292 (N_8292,N_4439,N_170);
and U8293 (N_8293,N_143,N_1007);
nand U8294 (N_8294,N_1533,N_4214);
nand U8295 (N_8295,N_1842,N_3335);
xnor U8296 (N_8296,N_4337,N_2277);
nand U8297 (N_8297,N_982,N_3050);
and U8298 (N_8298,N_1018,N_3794);
or U8299 (N_8299,N_1448,N_2206);
nand U8300 (N_8300,N_1700,N_1877);
nor U8301 (N_8301,N_1618,N_1756);
or U8302 (N_8302,N_4705,N_1782);
and U8303 (N_8303,N_1715,N_2908);
or U8304 (N_8304,N_1554,N_4600);
or U8305 (N_8305,N_3162,N_4472);
xor U8306 (N_8306,N_2643,N_4065);
nand U8307 (N_8307,N_186,N_1108);
xnor U8308 (N_8308,N_3086,N_2054);
or U8309 (N_8309,N_1474,N_3397);
nor U8310 (N_8310,N_3519,N_1264);
and U8311 (N_8311,N_4368,N_4489);
xor U8312 (N_8312,N_4906,N_2748);
nand U8313 (N_8313,N_2119,N_1371);
nand U8314 (N_8314,N_2524,N_3800);
or U8315 (N_8315,N_841,N_3113);
and U8316 (N_8316,N_3768,N_408);
or U8317 (N_8317,N_360,N_990);
nand U8318 (N_8318,N_2531,N_2434);
and U8319 (N_8319,N_4392,N_1607);
or U8320 (N_8320,N_4217,N_4391);
or U8321 (N_8321,N_3289,N_1270);
and U8322 (N_8322,N_3826,N_3372);
or U8323 (N_8323,N_2379,N_3349);
nor U8324 (N_8324,N_4864,N_633);
nand U8325 (N_8325,N_1933,N_3597);
or U8326 (N_8326,N_313,N_4116);
nor U8327 (N_8327,N_168,N_1497);
or U8328 (N_8328,N_4058,N_1129);
or U8329 (N_8329,N_1528,N_2118);
nor U8330 (N_8330,N_1647,N_3653);
and U8331 (N_8331,N_816,N_3994);
nand U8332 (N_8332,N_662,N_163);
or U8333 (N_8333,N_2639,N_2028);
xor U8334 (N_8334,N_1855,N_4818);
nand U8335 (N_8335,N_2512,N_3215);
xnor U8336 (N_8336,N_194,N_972);
or U8337 (N_8337,N_2063,N_651);
nand U8338 (N_8338,N_3379,N_3613);
nor U8339 (N_8339,N_4886,N_4083);
and U8340 (N_8340,N_4717,N_4735);
nor U8341 (N_8341,N_3098,N_2381);
or U8342 (N_8342,N_3755,N_2215);
or U8343 (N_8343,N_4376,N_4154);
nand U8344 (N_8344,N_2310,N_959);
xnor U8345 (N_8345,N_151,N_3999);
nand U8346 (N_8346,N_4627,N_3989);
or U8347 (N_8347,N_2909,N_440);
xnor U8348 (N_8348,N_281,N_3592);
xor U8349 (N_8349,N_132,N_1776);
and U8350 (N_8350,N_4699,N_4888);
or U8351 (N_8351,N_2244,N_1195);
xnor U8352 (N_8352,N_158,N_3200);
xor U8353 (N_8353,N_2227,N_229);
and U8354 (N_8354,N_3554,N_3405);
or U8355 (N_8355,N_3376,N_802);
nor U8356 (N_8356,N_122,N_1983);
or U8357 (N_8357,N_3291,N_4941);
nand U8358 (N_8358,N_3571,N_4512);
xor U8359 (N_8359,N_170,N_1597);
or U8360 (N_8360,N_3898,N_576);
and U8361 (N_8361,N_4815,N_4543);
nand U8362 (N_8362,N_1966,N_2675);
nand U8363 (N_8363,N_2725,N_239);
and U8364 (N_8364,N_1037,N_410);
and U8365 (N_8365,N_808,N_1512);
and U8366 (N_8366,N_876,N_1668);
xor U8367 (N_8367,N_111,N_3724);
and U8368 (N_8368,N_1343,N_583);
nor U8369 (N_8369,N_4713,N_4595);
and U8370 (N_8370,N_2686,N_1431);
nand U8371 (N_8371,N_1990,N_4555);
nor U8372 (N_8372,N_3792,N_3135);
and U8373 (N_8373,N_2797,N_2672);
xor U8374 (N_8374,N_375,N_3148);
xor U8375 (N_8375,N_4731,N_844);
xor U8376 (N_8376,N_2448,N_3912);
or U8377 (N_8377,N_4254,N_1041);
or U8378 (N_8378,N_564,N_634);
and U8379 (N_8379,N_1653,N_551);
and U8380 (N_8380,N_1411,N_3908);
xnor U8381 (N_8381,N_3586,N_2811);
xor U8382 (N_8382,N_2101,N_408);
nor U8383 (N_8383,N_4195,N_4995);
nand U8384 (N_8384,N_633,N_2729);
or U8385 (N_8385,N_2321,N_1718);
nand U8386 (N_8386,N_3142,N_1042);
and U8387 (N_8387,N_3391,N_2336);
xnor U8388 (N_8388,N_3749,N_3156);
and U8389 (N_8389,N_1532,N_1567);
and U8390 (N_8390,N_1520,N_1160);
nor U8391 (N_8391,N_1661,N_4644);
nor U8392 (N_8392,N_3606,N_3462);
and U8393 (N_8393,N_4301,N_606);
or U8394 (N_8394,N_1640,N_3989);
nor U8395 (N_8395,N_4905,N_2712);
xnor U8396 (N_8396,N_4286,N_359);
nor U8397 (N_8397,N_1130,N_3547);
and U8398 (N_8398,N_3550,N_2309);
nor U8399 (N_8399,N_1727,N_1123);
and U8400 (N_8400,N_2753,N_3773);
and U8401 (N_8401,N_3403,N_513);
xor U8402 (N_8402,N_4718,N_4593);
xor U8403 (N_8403,N_4533,N_635);
nand U8404 (N_8404,N_3451,N_4036);
or U8405 (N_8405,N_3898,N_745);
nor U8406 (N_8406,N_3056,N_1958);
or U8407 (N_8407,N_251,N_2822);
and U8408 (N_8408,N_718,N_1542);
xor U8409 (N_8409,N_1195,N_4610);
nor U8410 (N_8410,N_1679,N_4272);
and U8411 (N_8411,N_4092,N_3752);
xnor U8412 (N_8412,N_4759,N_3435);
xor U8413 (N_8413,N_4639,N_128);
nor U8414 (N_8414,N_2921,N_1434);
nor U8415 (N_8415,N_4931,N_2549);
xor U8416 (N_8416,N_450,N_3464);
and U8417 (N_8417,N_2886,N_4664);
nand U8418 (N_8418,N_4326,N_1067);
xnor U8419 (N_8419,N_1891,N_4839);
xnor U8420 (N_8420,N_4079,N_3072);
nor U8421 (N_8421,N_635,N_2520);
nand U8422 (N_8422,N_783,N_3818);
nand U8423 (N_8423,N_2804,N_1502);
xnor U8424 (N_8424,N_3512,N_1511);
and U8425 (N_8425,N_372,N_3427);
xnor U8426 (N_8426,N_3554,N_146);
and U8427 (N_8427,N_2668,N_783);
and U8428 (N_8428,N_3984,N_2571);
nand U8429 (N_8429,N_4885,N_4691);
and U8430 (N_8430,N_1654,N_1016);
or U8431 (N_8431,N_4314,N_257);
xor U8432 (N_8432,N_2437,N_3655);
or U8433 (N_8433,N_4104,N_499);
nand U8434 (N_8434,N_4216,N_107);
xor U8435 (N_8435,N_1143,N_4265);
nand U8436 (N_8436,N_3406,N_1116);
nand U8437 (N_8437,N_4957,N_3040);
or U8438 (N_8438,N_2849,N_973);
nand U8439 (N_8439,N_4803,N_3185);
or U8440 (N_8440,N_353,N_3544);
or U8441 (N_8441,N_4336,N_2646);
nor U8442 (N_8442,N_2164,N_768);
xnor U8443 (N_8443,N_158,N_474);
xor U8444 (N_8444,N_906,N_3058);
or U8445 (N_8445,N_224,N_4763);
xor U8446 (N_8446,N_2015,N_161);
xor U8447 (N_8447,N_3493,N_2405);
nor U8448 (N_8448,N_3885,N_1750);
or U8449 (N_8449,N_676,N_2104);
nor U8450 (N_8450,N_517,N_4549);
or U8451 (N_8451,N_3510,N_2449);
nand U8452 (N_8452,N_2508,N_3159);
or U8453 (N_8453,N_4282,N_3555);
or U8454 (N_8454,N_145,N_2864);
xor U8455 (N_8455,N_1026,N_408);
xnor U8456 (N_8456,N_528,N_3504);
nor U8457 (N_8457,N_2453,N_4417);
or U8458 (N_8458,N_605,N_1645);
xor U8459 (N_8459,N_2629,N_1621);
or U8460 (N_8460,N_2974,N_3575);
or U8461 (N_8461,N_1593,N_2895);
and U8462 (N_8462,N_4397,N_3974);
xnor U8463 (N_8463,N_966,N_4954);
nor U8464 (N_8464,N_567,N_3504);
xnor U8465 (N_8465,N_3007,N_946);
xnor U8466 (N_8466,N_3228,N_2881);
and U8467 (N_8467,N_1147,N_2930);
nand U8468 (N_8468,N_528,N_3223);
and U8469 (N_8469,N_3026,N_2015);
or U8470 (N_8470,N_4866,N_4919);
and U8471 (N_8471,N_4047,N_1949);
nor U8472 (N_8472,N_3351,N_2618);
nand U8473 (N_8473,N_311,N_3757);
and U8474 (N_8474,N_364,N_837);
nand U8475 (N_8475,N_3898,N_778);
and U8476 (N_8476,N_1767,N_262);
and U8477 (N_8477,N_324,N_2080);
and U8478 (N_8478,N_763,N_1778);
or U8479 (N_8479,N_4381,N_530);
or U8480 (N_8480,N_3587,N_4977);
nor U8481 (N_8481,N_516,N_1489);
and U8482 (N_8482,N_3864,N_3356);
xor U8483 (N_8483,N_3143,N_3330);
or U8484 (N_8484,N_2016,N_3465);
xor U8485 (N_8485,N_2282,N_1722);
or U8486 (N_8486,N_2378,N_2653);
xor U8487 (N_8487,N_1559,N_1854);
nor U8488 (N_8488,N_554,N_4662);
nand U8489 (N_8489,N_2596,N_2242);
xnor U8490 (N_8490,N_2120,N_4195);
xor U8491 (N_8491,N_3019,N_1800);
and U8492 (N_8492,N_503,N_1782);
and U8493 (N_8493,N_1118,N_4721);
nor U8494 (N_8494,N_3355,N_2691);
nor U8495 (N_8495,N_1013,N_1827);
or U8496 (N_8496,N_4135,N_1268);
nand U8497 (N_8497,N_1674,N_596);
xnor U8498 (N_8498,N_4602,N_1596);
nor U8499 (N_8499,N_3559,N_4570);
nand U8500 (N_8500,N_1488,N_875);
and U8501 (N_8501,N_1340,N_3972);
or U8502 (N_8502,N_981,N_2245);
nand U8503 (N_8503,N_2239,N_3880);
or U8504 (N_8504,N_1391,N_1437);
nand U8505 (N_8505,N_4464,N_3148);
or U8506 (N_8506,N_3547,N_1096);
or U8507 (N_8507,N_682,N_4288);
and U8508 (N_8508,N_304,N_3150);
and U8509 (N_8509,N_3473,N_427);
nand U8510 (N_8510,N_207,N_4085);
and U8511 (N_8511,N_3886,N_3600);
or U8512 (N_8512,N_2373,N_1658);
and U8513 (N_8513,N_2638,N_4720);
nor U8514 (N_8514,N_223,N_3713);
or U8515 (N_8515,N_2843,N_1737);
nand U8516 (N_8516,N_2111,N_942);
nor U8517 (N_8517,N_4776,N_133);
and U8518 (N_8518,N_4733,N_3112);
nor U8519 (N_8519,N_2810,N_2940);
and U8520 (N_8520,N_2213,N_4345);
and U8521 (N_8521,N_143,N_3874);
and U8522 (N_8522,N_4499,N_636);
nor U8523 (N_8523,N_898,N_3041);
or U8524 (N_8524,N_3262,N_3539);
xor U8525 (N_8525,N_2406,N_4334);
xor U8526 (N_8526,N_1756,N_2432);
and U8527 (N_8527,N_1275,N_4662);
nor U8528 (N_8528,N_3759,N_3436);
nand U8529 (N_8529,N_4164,N_217);
nand U8530 (N_8530,N_752,N_1272);
xor U8531 (N_8531,N_459,N_4765);
xnor U8532 (N_8532,N_1039,N_4785);
nor U8533 (N_8533,N_878,N_3245);
and U8534 (N_8534,N_663,N_1069);
nor U8535 (N_8535,N_2931,N_4445);
nand U8536 (N_8536,N_2634,N_3177);
xnor U8537 (N_8537,N_3980,N_3312);
nor U8538 (N_8538,N_534,N_2583);
nand U8539 (N_8539,N_3013,N_223);
or U8540 (N_8540,N_1203,N_12);
or U8541 (N_8541,N_1460,N_3768);
xor U8542 (N_8542,N_4339,N_1731);
nand U8543 (N_8543,N_3590,N_2387);
xnor U8544 (N_8544,N_1958,N_2244);
and U8545 (N_8545,N_2864,N_1258);
nor U8546 (N_8546,N_1858,N_2130);
nand U8547 (N_8547,N_2182,N_3870);
xor U8548 (N_8548,N_1556,N_3909);
and U8549 (N_8549,N_3866,N_3728);
nor U8550 (N_8550,N_1722,N_2489);
nand U8551 (N_8551,N_3631,N_2261);
nor U8552 (N_8552,N_3829,N_3698);
and U8553 (N_8553,N_4052,N_911);
nand U8554 (N_8554,N_570,N_1168);
and U8555 (N_8555,N_4767,N_1664);
xnor U8556 (N_8556,N_2719,N_4280);
and U8557 (N_8557,N_4884,N_1784);
nand U8558 (N_8558,N_504,N_4977);
or U8559 (N_8559,N_897,N_4294);
and U8560 (N_8560,N_4773,N_17);
xnor U8561 (N_8561,N_3936,N_2723);
or U8562 (N_8562,N_2330,N_2234);
and U8563 (N_8563,N_3356,N_1267);
nand U8564 (N_8564,N_2790,N_3250);
nand U8565 (N_8565,N_3940,N_4233);
nor U8566 (N_8566,N_4556,N_3688);
xnor U8567 (N_8567,N_2567,N_2505);
xor U8568 (N_8568,N_4735,N_2222);
nor U8569 (N_8569,N_792,N_719);
or U8570 (N_8570,N_1800,N_4062);
nor U8571 (N_8571,N_775,N_795);
and U8572 (N_8572,N_3120,N_4471);
xnor U8573 (N_8573,N_244,N_1198);
xnor U8574 (N_8574,N_3996,N_2832);
nor U8575 (N_8575,N_3566,N_3768);
and U8576 (N_8576,N_992,N_4309);
xnor U8577 (N_8577,N_3255,N_4906);
and U8578 (N_8578,N_4123,N_1803);
or U8579 (N_8579,N_3567,N_3821);
or U8580 (N_8580,N_3074,N_4020);
nand U8581 (N_8581,N_2889,N_3480);
nor U8582 (N_8582,N_4146,N_3836);
nand U8583 (N_8583,N_490,N_4166);
or U8584 (N_8584,N_2283,N_1865);
nand U8585 (N_8585,N_2304,N_4148);
and U8586 (N_8586,N_3322,N_125);
nand U8587 (N_8587,N_3272,N_2051);
or U8588 (N_8588,N_1218,N_4987);
nor U8589 (N_8589,N_2872,N_4895);
and U8590 (N_8590,N_1067,N_3812);
or U8591 (N_8591,N_4402,N_4006);
and U8592 (N_8592,N_4930,N_2095);
nor U8593 (N_8593,N_3836,N_3949);
nand U8594 (N_8594,N_3140,N_1416);
and U8595 (N_8595,N_4662,N_2018);
or U8596 (N_8596,N_1247,N_1448);
nand U8597 (N_8597,N_984,N_4843);
nand U8598 (N_8598,N_4420,N_2658);
or U8599 (N_8599,N_1240,N_820);
and U8600 (N_8600,N_2899,N_3289);
nor U8601 (N_8601,N_3555,N_3736);
nand U8602 (N_8602,N_3159,N_379);
xor U8603 (N_8603,N_4791,N_1638);
nor U8604 (N_8604,N_995,N_4217);
xnor U8605 (N_8605,N_884,N_143);
and U8606 (N_8606,N_4388,N_1650);
and U8607 (N_8607,N_323,N_4584);
and U8608 (N_8608,N_1488,N_1121);
xor U8609 (N_8609,N_4725,N_588);
and U8610 (N_8610,N_3753,N_124);
nor U8611 (N_8611,N_1614,N_1235);
nand U8612 (N_8612,N_705,N_1508);
nand U8613 (N_8613,N_3649,N_4652);
nor U8614 (N_8614,N_2869,N_2989);
nand U8615 (N_8615,N_1016,N_3050);
xor U8616 (N_8616,N_1510,N_1380);
nor U8617 (N_8617,N_1412,N_2168);
nor U8618 (N_8618,N_2434,N_382);
xor U8619 (N_8619,N_845,N_645);
xnor U8620 (N_8620,N_2679,N_2435);
nand U8621 (N_8621,N_360,N_2604);
nor U8622 (N_8622,N_3121,N_1746);
nand U8623 (N_8623,N_4210,N_1820);
and U8624 (N_8624,N_2932,N_2073);
nor U8625 (N_8625,N_3102,N_6);
xnor U8626 (N_8626,N_858,N_4535);
and U8627 (N_8627,N_3260,N_1554);
and U8628 (N_8628,N_1354,N_1734);
and U8629 (N_8629,N_1962,N_4037);
or U8630 (N_8630,N_3404,N_557);
and U8631 (N_8631,N_3768,N_4513);
or U8632 (N_8632,N_2507,N_96);
nand U8633 (N_8633,N_3762,N_1513);
nor U8634 (N_8634,N_2043,N_432);
nor U8635 (N_8635,N_1093,N_2440);
xnor U8636 (N_8636,N_3845,N_2132);
nand U8637 (N_8637,N_3822,N_767);
xnor U8638 (N_8638,N_549,N_2040);
xnor U8639 (N_8639,N_1104,N_1730);
or U8640 (N_8640,N_4267,N_1560);
nor U8641 (N_8641,N_2041,N_87);
nor U8642 (N_8642,N_1442,N_263);
or U8643 (N_8643,N_536,N_1967);
xnor U8644 (N_8644,N_4100,N_4610);
nand U8645 (N_8645,N_3469,N_4461);
or U8646 (N_8646,N_269,N_4657);
and U8647 (N_8647,N_193,N_3357);
nor U8648 (N_8648,N_4665,N_2649);
nand U8649 (N_8649,N_3752,N_2420);
nor U8650 (N_8650,N_1143,N_3944);
and U8651 (N_8651,N_900,N_1150);
nand U8652 (N_8652,N_4328,N_2055);
xor U8653 (N_8653,N_4774,N_3534);
xnor U8654 (N_8654,N_2920,N_1695);
xnor U8655 (N_8655,N_4215,N_2575);
nand U8656 (N_8656,N_949,N_1555);
nor U8657 (N_8657,N_3829,N_2621);
nand U8658 (N_8658,N_2849,N_4301);
nor U8659 (N_8659,N_1908,N_4854);
or U8660 (N_8660,N_4582,N_1082);
xor U8661 (N_8661,N_2684,N_1455);
nand U8662 (N_8662,N_4754,N_536);
nand U8663 (N_8663,N_4268,N_1611);
xnor U8664 (N_8664,N_4417,N_1418);
nor U8665 (N_8665,N_2010,N_3507);
nand U8666 (N_8666,N_425,N_346);
or U8667 (N_8667,N_3612,N_3792);
nand U8668 (N_8668,N_2390,N_1520);
nor U8669 (N_8669,N_3398,N_1029);
nor U8670 (N_8670,N_887,N_4426);
nor U8671 (N_8671,N_419,N_311);
nor U8672 (N_8672,N_432,N_3463);
nand U8673 (N_8673,N_1457,N_4699);
or U8674 (N_8674,N_2630,N_4691);
nor U8675 (N_8675,N_2947,N_2505);
or U8676 (N_8676,N_3828,N_3386);
xnor U8677 (N_8677,N_2236,N_3509);
and U8678 (N_8678,N_1946,N_1756);
nand U8679 (N_8679,N_3517,N_4579);
xnor U8680 (N_8680,N_3157,N_2502);
xnor U8681 (N_8681,N_1678,N_2754);
xnor U8682 (N_8682,N_2028,N_3080);
nand U8683 (N_8683,N_4626,N_1862);
nand U8684 (N_8684,N_3768,N_3122);
xnor U8685 (N_8685,N_2105,N_1478);
and U8686 (N_8686,N_1582,N_3784);
and U8687 (N_8687,N_1596,N_2169);
nand U8688 (N_8688,N_189,N_3490);
nand U8689 (N_8689,N_206,N_4264);
xor U8690 (N_8690,N_598,N_1625);
and U8691 (N_8691,N_40,N_2935);
or U8692 (N_8692,N_4355,N_3758);
nand U8693 (N_8693,N_2270,N_4276);
or U8694 (N_8694,N_1759,N_3945);
and U8695 (N_8695,N_2729,N_1368);
and U8696 (N_8696,N_3118,N_3488);
nand U8697 (N_8697,N_1673,N_1211);
xor U8698 (N_8698,N_4688,N_659);
nand U8699 (N_8699,N_4733,N_4216);
xor U8700 (N_8700,N_2540,N_266);
nand U8701 (N_8701,N_744,N_3608);
xnor U8702 (N_8702,N_4813,N_578);
and U8703 (N_8703,N_3641,N_2780);
xnor U8704 (N_8704,N_4918,N_2332);
nand U8705 (N_8705,N_1159,N_893);
nor U8706 (N_8706,N_1211,N_4444);
nand U8707 (N_8707,N_27,N_3080);
and U8708 (N_8708,N_472,N_4548);
nand U8709 (N_8709,N_883,N_3586);
or U8710 (N_8710,N_1296,N_2709);
and U8711 (N_8711,N_700,N_4090);
nand U8712 (N_8712,N_1489,N_4635);
or U8713 (N_8713,N_1543,N_611);
nor U8714 (N_8714,N_1219,N_4709);
or U8715 (N_8715,N_2265,N_1409);
and U8716 (N_8716,N_1345,N_4121);
nor U8717 (N_8717,N_1935,N_2439);
nand U8718 (N_8718,N_4610,N_3604);
nor U8719 (N_8719,N_4413,N_3231);
xnor U8720 (N_8720,N_4387,N_906);
or U8721 (N_8721,N_4022,N_1180);
nand U8722 (N_8722,N_2681,N_3200);
nand U8723 (N_8723,N_438,N_3704);
and U8724 (N_8724,N_3999,N_1580);
xnor U8725 (N_8725,N_2262,N_2502);
nor U8726 (N_8726,N_2590,N_4864);
nor U8727 (N_8727,N_4913,N_2079);
and U8728 (N_8728,N_1800,N_2001);
nand U8729 (N_8729,N_949,N_3811);
and U8730 (N_8730,N_2146,N_1902);
xnor U8731 (N_8731,N_4679,N_3701);
or U8732 (N_8732,N_3817,N_3068);
and U8733 (N_8733,N_888,N_3258);
and U8734 (N_8734,N_3877,N_2805);
xnor U8735 (N_8735,N_50,N_3126);
and U8736 (N_8736,N_1957,N_1273);
xnor U8737 (N_8737,N_4707,N_95);
nand U8738 (N_8738,N_4702,N_1961);
and U8739 (N_8739,N_4124,N_4458);
or U8740 (N_8740,N_4347,N_4019);
or U8741 (N_8741,N_164,N_1354);
nand U8742 (N_8742,N_1585,N_28);
and U8743 (N_8743,N_134,N_2758);
or U8744 (N_8744,N_106,N_458);
or U8745 (N_8745,N_975,N_2982);
nand U8746 (N_8746,N_902,N_2633);
xnor U8747 (N_8747,N_4876,N_3352);
or U8748 (N_8748,N_3815,N_2811);
xnor U8749 (N_8749,N_2692,N_4780);
nor U8750 (N_8750,N_3860,N_49);
nand U8751 (N_8751,N_97,N_3736);
or U8752 (N_8752,N_1959,N_2853);
xnor U8753 (N_8753,N_108,N_4619);
xor U8754 (N_8754,N_4032,N_2737);
nand U8755 (N_8755,N_1211,N_1071);
and U8756 (N_8756,N_3980,N_1904);
and U8757 (N_8757,N_3447,N_4777);
or U8758 (N_8758,N_3338,N_334);
xor U8759 (N_8759,N_2672,N_3340);
nor U8760 (N_8760,N_1013,N_3249);
nand U8761 (N_8761,N_1793,N_3387);
nand U8762 (N_8762,N_1664,N_3411);
nor U8763 (N_8763,N_4247,N_410);
nor U8764 (N_8764,N_1913,N_497);
nor U8765 (N_8765,N_3275,N_4149);
and U8766 (N_8766,N_3079,N_4885);
nor U8767 (N_8767,N_3968,N_3488);
nor U8768 (N_8768,N_2358,N_4184);
or U8769 (N_8769,N_4213,N_473);
or U8770 (N_8770,N_2030,N_511);
nand U8771 (N_8771,N_816,N_1695);
xnor U8772 (N_8772,N_2274,N_1017);
nor U8773 (N_8773,N_1632,N_2529);
xnor U8774 (N_8774,N_1237,N_4047);
nor U8775 (N_8775,N_3518,N_4505);
nand U8776 (N_8776,N_3379,N_2276);
nor U8777 (N_8777,N_631,N_3584);
and U8778 (N_8778,N_1562,N_3185);
xor U8779 (N_8779,N_738,N_4082);
or U8780 (N_8780,N_1890,N_2155);
xnor U8781 (N_8781,N_2521,N_1392);
and U8782 (N_8782,N_4781,N_15);
or U8783 (N_8783,N_4560,N_3096);
or U8784 (N_8784,N_572,N_1984);
nor U8785 (N_8785,N_4584,N_3876);
and U8786 (N_8786,N_233,N_4190);
nand U8787 (N_8787,N_2144,N_3195);
and U8788 (N_8788,N_1187,N_1924);
nor U8789 (N_8789,N_468,N_3458);
and U8790 (N_8790,N_3381,N_2956);
nor U8791 (N_8791,N_4598,N_3180);
and U8792 (N_8792,N_833,N_4530);
nand U8793 (N_8793,N_1563,N_2263);
xnor U8794 (N_8794,N_775,N_974);
nor U8795 (N_8795,N_667,N_4650);
or U8796 (N_8796,N_631,N_4415);
nand U8797 (N_8797,N_1033,N_4160);
nor U8798 (N_8798,N_3386,N_2859);
nand U8799 (N_8799,N_1510,N_4933);
and U8800 (N_8800,N_1981,N_2382);
nand U8801 (N_8801,N_1881,N_4420);
nor U8802 (N_8802,N_876,N_2925);
or U8803 (N_8803,N_4532,N_1978);
nor U8804 (N_8804,N_3590,N_3099);
nor U8805 (N_8805,N_3490,N_3391);
nand U8806 (N_8806,N_1462,N_1611);
or U8807 (N_8807,N_4254,N_3683);
nor U8808 (N_8808,N_3149,N_3319);
xnor U8809 (N_8809,N_2535,N_2699);
xnor U8810 (N_8810,N_2522,N_1391);
or U8811 (N_8811,N_1621,N_618);
nor U8812 (N_8812,N_4811,N_3045);
nor U8813 (N_8813,N_1878,N_565);
or U8814 (N_8814,N_3899,N_199);
xor U8815 (N_8815,N_2403,N_2398);
or U8816 (N_8816,N_4991,N_1172);
nand U8817 (N_8817,N_3137,N_1106);
nand U8818 (N_8818,N_1058,N_2449);
or U8819 (N_8819,N_4804,N_4597);
nand U8820 (N_8820,N_1803,N_3862);
nand U8821 (N_8821,N_165,N_1406);
or U8822 (N_8822,N_1551,N_3902);
xor U8823 (N_8823,N_4485,N_974);
nand U8824 (N_8824,N_2522,N_3555);
nand U8825 (N_8825,N_100,N_575);
and U8826 (N_8826,N_4942,N_2547);
nor U8827 (N_8827,N_2438,N_2098);
and U8828 (N_8828,N_3932,N_3846);
xnor U8829 (N_8829,N_2894,N_4043);
xor U8830 (N_8830,N_3835,N_2090);
and U8831 (N_8831,N_2771,N_563);
and U8832 (N_8832,N_3761,N_3397);
xnor U8833 (N_8833,N_2080,N_2974);
xor U8834 (N_8834,N_4422,N_2183);
nand U8835 (N_8835,N_3262,N_616);
xor U8836 (N_8836,N_3274,N_3300);
nand U8837 (N_8837,N_1362,N_4044);
xor U8838 (N_8838,N_638,N_130);
xnor U8839 (N_8839,N_3348,N_2402);
and U8840 (N_8840,N_2389,N_3806);
nand U8841 (N_8841,N_1609,N_2212);
and U8842 (N_8842,N_96,N_3432);
nand U8843 (N_8843,N_2454,N_1684);
and U8844 (N_8844,N_4071,N_2080);
xnor U8845 (N_8845,N_4519,N_3851);
xnor U8846 (N_8846,N_1605,N_795);
nor U8847 (N_8847,N_2462,N_1340);
or U8848 (N_8848,N_3653,N_3483);
nand U8849 (N_8849,N_2338,N_605);
nand U8850 (N_8850,N_1293,N_2406);
nor U8851 (N_8851,N_468,N_2475);
nor U8852 (N_8852,N_782,N_2115);
or U8853 (N_8853,N_3860,N_1047);
xnor U8854 (N_8854,N_721,N_2045);
nand U8855 (N_8855,N_4908,N_2536);
or U8856 (N_8856,N_4933,N_3371);
xnor U8857 (N_8857,N_2060,N_1978);
and U8858 (N_8858,N_2906,N_1156);
nand U8859 (N_8859,N_805,N_4119);
nand U8860 (N_8860,N_4413,N_2763);
and U8861 (N_8861,N_1385,N_4900);
or U8862 (N_8862,N_4434,N_2851);
nand U8863 (N_8863,N_4476,N_4397);
nor U8864 (N_8864,N_116,N_4755);
nand U8865 (N_8865,N_4783,N_1844);
or U8866 (N_8866,N_1582,N_77);
nand U8867 (N_8867,N_2737,N_2517);
nand U8868 (N_8868,N_2863,N_4235);
or U8869 (N_8869,N_3561,N_1072);
and U8870 (N_8870,N_946,N_2851);
or U8871 (N_8871,N_1099,N_3773);
and U8872 (N_8872,N_4580,N_3998);
nand U8873 (N_8873,N_4428,N_4944);
xnor U8874 (N_8874,N_4413,N_1903);
or U8875 (N_8875,N_685,N_744);
and U8876 (N_8876,N_915,N_3034);
or U8877 (N_8877,N_123,N_3641);
nor U8878 (N_8878,N_3301,N_905);
nor U8879 (N_8879,N_375,N_407);
or U8880 (N_8880,N_4778,N_2330);
or U8881 (N_8881,N_3226,N_2083);
xnor U8882 (N_8882,N_2833,N_1410);
nand U8883 (N_8883,N_4736,N_395);
and U8884 (N_8884,N_3832,N_3050);
xnor U8885 (N_8885,N_3069,N_4381);
and U8886 (N_8886,N_3108,N_2617);
nand U8887 (N_8887,N_892,N_4174);
xor U8888 (N_8888,N_4648,N_2095);
or U8889 (N_8889,N_2197,N_4115);
nor U8890 (N_8890,N_1205,N_2613);
xor U8891 (N_8891,N_34,N_2155);
xor U8892 (N_8892,N_3134,N_3249);
and U8893 (N_8893,N_1978,N_859);
nor U8894 (N_8894,N_1570,N_1274);
nor U8895 (N_8895,N_4845,N_2585);
or U8896 (N_8896,N_4599,N_4858);
xnor U8897 (N_8897,N_594,N_724);
nor U8898 (N_8898,N_4647,N_65);
or U8899 (N_8899,N_2227,N_586);
or U8900 (N_8900,N_2469,N_3172);
xnor U8901 (N_8901,N_3217,N_2777);
or U8902 (N_8902,N_3847,N_4650);
nand U8903 (N_8903,N_1955,N_2586);
or U8904 (N_8904,N_4306,N_4641);
xnor U8905 (N_8905,N_4455,N_1688);
nand U8906 (N_8906,N_43,N_2700);
xor U8907 (N_8907,N_193,N_2824);
xnor U8908 (N_8908,N_4845,N_1629);
or U8909 (N_8909,N_2369,N_1013);
nand U8910 (N_8910,N_3920,N_1702);
or U8911 (N_8911,N_3556,N_3015);
nand U8912 (N_8912,N_4091,N_1159);
or U8913 (N_8913,N_792,N_4608);
nor U8914 (N_8914,N_2253,N_4809);
and U8915 (N_8915,N_770,N_2990);
xnor U8916 (N_8916,N_2355,N_4735);
xnor U8917 (N_8917,N_4799,N_3880);
nand U8918 (N_8918,N_3886,N_3354);
and U8919 (N_8919,N_2142,N_663);
xor U8920 (N_8920,N_3634,N_3856);
nor U8921 (N_8921,N_3186,N_1522);
nand U8922 (N_8922,N_1540,N_1678);
and U8923 (N_8923,N_3348,N_1916);
xor U8924 (N_8924,N_1001,N_2189);
nor U8925 (N_8925,N_1007,N_2686);
and U8926 (N_8926,N_4986,N_620);
nand U8927 (N_8927,N_2000,N_3973);
nor U8928 (N_8928,N_1506,N_4053);
nor U8929 (N_8929,N_625,N_2839);
and U8930 (N_8930,N_4368,N_4726);
or U8931 (N_8931,N_2902,N_4050);
xnor U8932 (N_8932,N_1202,N_526);
and U8933 (N_8933,N_3328,N_478);
nand U8934 (N_8934,N_3575,N_4223);
nand U8935 (N_8935,N_2385,N_3315);
or U8936 (N_8936,N_269,N_3748);
xor U8937 (N_8937,N_4293,N_4786);
and U8938 (N_8938,N_1020,N_2127);
xor U8939 (N_8939,N_4340,N_3534);
nand U8940 (N_8940,N_1305,N_3820);
nor U8941 (N_8941,N_495,N_4816);
and U8942 (N_8942,N_178,N_2986);
nand U8943 (N_8943,N_1224,N_3379);
nor U8944 (N_8944,N_2005,N_2112);
xnor U8945 (N_8945,N_3426,N_4201);
nand U8946 (N_8946,N_1920,N_3295);
or U8947 (N_8947,N_3331,N_4640);
and U8948 (N_8948,N_1281,N_4655);
or U8949 (N_8949,N_4155,N_2653);
nor U8950 (N_8950,N_3817,N_2462);
or U8951 (N_8951,N_1794,N_1629);
or U8952 (N_8952,N_3539,N_1434);
or U8953 (N_8953,N_3215,N_3395);
nor U8954 (N_8954,N_1883,N_2773);
xnor U8955 (N_8955,N_2860,N_792);
and U8956 (N_8956,N_1821,N_905);
nand U8957 (N_8957,N_761,N_4500);
nand U8958 (N_8958,N_2332,N_3565);
and U8959 (N_8959,N_4708,N_3675);
xnor U8960 (N_8960,N_905,N_4094);
nor U8961 (N_8961,N_4513,N_1097);
xor U8962 (N_8962,N_3352,N_1273);
or U8963 (N_8963,N_4743,N_684);
nand U8964 (N_8964,N_4469,N_199);
nand U8965 (N_8965,N_2697,N_689);
and U8966 (N_8966,N_3717,N_1709);
and U8967 (N_8967,N_4483,N_3706);
nand U8968 (N_8968,N_3454,N_1997);
nand U8969 (N_8969,N_4675,N_625);
nand U8970 (N_8970,N_512,N_168);
nor U8971 (N_8971,N_4753,N_4658);
nor U8972 (N_8972,N_3207,N_342);
or U8973 (N_8973,N_3117,N_4097);
nand U8974 (N_8974,N_1465,N_3792);
xor U8975 (N_8975,N_2220,N_69);
nand U8976 (N_8976,N_2439,N_3755);
or U8977 (N_8977,N_436,N_2580);
xnor U8978 (N_8978,N_4530,N_2331);
or U8979 (N_8979,N_4064,N_2087);
or U8980 (N_8980,N_3150,N_943);
and U8981 (N_8981,N_3503,N_3093);
nor U8982 (N_8982,N_339,N_2194);
nand U8983 (N_8983,N_1043,N_1465);
nor U8984 (N_8984,N_2497,N_2761);
nand U8985 (N_8985,N_3378,N_1652);
or U8986 (N_8986,N_4603,N_2274);
nor U8987 (N_8987,N_4522,N_2631);
and U8988 (N_8988,N_1084,N_4039);
nor U8989 (N_8989,N_984,N_2558);
nand U8990 (N_8990,N_1704,N_4096);
or U8991 (N_8991,N_4818,N_3424);
nand U8992 (N_8992,N_2464,N_2805);
xnor U8993 (N_8993,N_3496,N_4403);
or U8994 (N_8994,N_2603,N_1280);
nor U8995 (N_8995,N_3175,N_744);
xnor U8996 (N_8996,N_2539,N_4497);
xnor U8997 (N_8997,N_4449,N_1681);
xor U8998 (N_8998,N_3381,N_1218);
nand U8999 (N_8999,N_4526,N_326);
nand U9000 (N_9000,N_458,N_1723);
xor U9001 (N_9001,N_847,N_1525);
xor U9002 (N_9002,N_493,N_561);
nor U9003 (N_9003,N_760,N_475);
xor U9004 (N_9004,N_4079,N_3662);
and U9005 (N_9005,N_3422,N_3267);
nor U9006 (N_9006,N_2108,N_2223);
xor U9007 (N_9007,N_3429,N_4800);
nor U9008 (N_9008,N_4437,N_2923);
nor U9009 (N_9009,N_3286,N_477);
nor U9010 (N_9010,N_1184,N_4868);
nand U9011 (N_9011,N_4386,N_397);
nor U9012 (N_9012,N_2194,N_66);
nor U9013 (N_9013,N_1384,N_1188);
and U9014 (N_9014,N_1859,N_330);
xnor U9015 (N_9015,N_3609,N_3250);
xnor U9016 (N_9016,N_1238,N_4316);
and U9017 (N_9017,N_3965,N_2901);
nand U9018 (N_9018,N_4238,N_3118);
xor U9019 (N_9019,N_2260,N_3708);
and U9020 (N_9020,N_4070,N_442);
nand U9021 (N_9021,N_1206,N_846);
and U9022 (N_9022,N_2839,N_2015);
or U9023 (N_9023,N_1226,N_1044);
and U9024 (N_9024,N_3714,N_2973);
or U9025 (N_9025,N_1254,N_470);
nand U9026 (N_9026,N_2697,N_2629);
xor U9027 (N_9027,N_3404,N_3601);
nand U9028 (N_9028,N_4797,N_4382);
or U9029 (N_9029,N_4782,N_2611);
or U9030 (N_9030,N_3523,N_3758);
or U9031 (N_9031,N_3669,N_2128);
and U9032 (N_9032,N_920,N_1670);
and U9033 (N_9033,N_2591,N_4266);
nand U9034 (N_9034,N_1,N_4618);
or U9035 (N_9035,N_2669,N_3917);
nor U9036 (N_9036,N_1971,N_3793);
nor U9037 (N_9037,N_185,N_8);
and U9038 (N_9038,N_2101,N_2457);
and U9039 (N_9039,N_4294,N_4304);
or U9040 (N_9040,N_4962,N_2926);
nor U9041 (N_9041,N_2746,N_3212);
xnor U9042 (N_9042,N_3085,N_2039);
nand U9043 (N_9043,N_4296,N_3972);
nand U9044 (N_9044,N_1187,N_4556);
and U9045 (N_9045,N_4894,N_2368);
or U9046 (N_9046,N_4601,N_3544);
nor U9047 (N_9047,N_2836,N_2871);
nand U9048 (N_9048,N_3707,N_4247);
nand U9049 (N_9049,N_4279,N_977);
or U9050 (N_9050,N_4184,N_1115);
or U9051 (N_9051,N_2465,N_4405);
or U9052 (N_9052,N_2582,N_2387);
or U9053 (N_9053,N_2965,N_453);
and U9054 (N_9054,N_1546,N_3818);
and U9055 (N_9055,N_2422,N_1715);
nand U9056 (N_9056,N_1862,N_4723);
or U9057 (N_9057,N_2843,N_1227);
or U9058 (N_9058,N_2059,N_997);
or U9059 (N_9059,N_2751,N_2068);
and U9060 (N_9060,N_3417,N_1167);
nand U9061 (N_9061,N_2188,N_1785);
or U9062 (N_9062,N_3646,N_1128);
or U9063 (N_9063,N_1833,N_1193);
and U9064 (N_9064,N_1934,N_649);
nor U9065 (N_9065,N_2242,N_336);
nand U9066 (N_9066,N_4779,N_4525);
or U9067 (N_9067,N_4915,N_3614);
nand U9068 (N_9068,N_3113,N_2198);
xnor U9069 (N_9069,N_1412,N_3330);
or U9070 (N_9070,N_2157,N_1494);
xor U9071 (N_9071,N_3085,N_3372);
xor U9072 (N_9072,N_3461,N_89);
or U9073 (N_9073,N_3121,N_120);
nor U9074 (N_9074,N_2051,N_3985);
or U9075 (N_9075,N_4844,N_4485);
xor U9076 (N_9076,N_1480,N_1172);
nand U9077 (N_9077,N_4203,N_1858);
nor U9078 (N_9078,N_1111,N_2749);
nor U9079 (N_9079,N_94,N_3158);
and U9080 (N_9080,N_1281,N_2370);
or U9081 (N_9081,N_3621,N_1273);
or U9082 (N_9082,N_1730,N_3518);
or U9083 (N_9083,N_3719,N_3715);
xnor U9084 (N_9084,N_638,N_1804);
nand U9085 (N_9085,N_3883,N_1752);
xnor U9086 (N_9086,N_4217,N_4256);
or U9087 (N_9087,N_407,N_4207);
nor U9088 (N_9088,N_468,N_4792);
nor U9089 (N_9089,N_3202,N_2176);
nand U9090 (N_9090,N_3560,N_578);
and U9091 (N_9091,N_4882,N_4373);
nor U9092 (N_9092,N_1621,N_2531);
nor U9093 (N_9093,N_2587,N_3757);
nor U9094 (N_9094,N_860,N_1231);
xnor U9095 (N_9095,N_4957,N_3766);
or U9096 (N_9096,N_3149,N_753);
nand U9097 (N_9097,N_3854,N_4079);
nand U9098 (N_9098,N_4160,N_1452);
xnor U9099 (N_9099,N_2709,N_1845);
or U9100 (N_9100,N_4054,N_4828);
xnor U9101 (N_9101,N_3307,N_2111);
and U9102 (N_9102,N_260,N_496);
and U9103 (N_9103,N_2950,N_4748);
nor U9104 (N_9104,N_3935,N_2911);
nor U9105 (N_9105,N_4195,N_50);
nand U9106 (N_9106,N_4049,N_699);
or U9107 (N_9107,N_88,N_702);
nand U9108 (N_9108,N_2373,N_4222);
nand U9109 (N_9109,N_2021,N_584);
or U9110 (N_9110,N_4539,N_4784);
xor U9111 (N_9111,N_4139,N_4030);
or U9112 (N_9112,N_2929,N_1913);
and U9113 (N_9113,N_4825,N_225);
nand U9114 (N_9114,N_4263,N_1486);
xor U9115 (N_9115,N_2982,N_4860);
xor U9116 (N_9116,N_4772,N_3557);
and U9117 (N_9117,N_2816,N_4682);
nor U9118 (N_9118,N_4188,N_834);
xor U9119 (N_9119,N_1242,N_2899);
xnor U9120 (N_9120,N_248,N_3782);
nor U9121 (N_9121,N_412,N_3405);
or U9122 (N_9122,N_1173,N_3916);
xnor U9123 (N_9123,N_4774,N_2856);
and U9124 (N_9124,N_1237,N_2357);
xor U9125 (N_9125,N_2163,N_1911);
and U9126 (N_9126,N_1892,N_2982);
and U9127 (N_9127,N_3369,N_4460);
or U9128 (N_9128,N_3205,N_1613);
or U9129 (N_9129,N_550,N_1164);
xor U9130 (N_9130,N_4946,N_605);
xor U9131 (N_9131,N_3872,N_3989);
nor U9132 (N_9132,N_2338,N_1553);
xnor U9133 (N_9133,N_3000,N_3794);
nor U9134 (N_9134,N_160,N_2988);
xnor U9135 (N_9135,N_1836,N_4811);
or U9136 (N_9136,N_3456,N_4328);
and U9137 (N_9137,N_4098,N_4956);
xor U9138 (N_9138,N_1053,N_4264);
or U9139 (N_9139,N_4338,N_3834);
xnor U9140 (N_9140,N_1948,N_2043);
nand U9141 (N_9141,N_3194,N_1023);
nor U9142 (N_9142,N_3643,N_478);
nor U9143 (N_9143,N_3532,N_4719);
xor U9144 (N_9144,N_3609,N_4068);
nand U9145 (N_9145,N_202,N_4046);
nor U9146 (N_9146,N_2277,N_11);
nor U9147 (N_9147,N_4161,N_1132);
nand U9148 (N_9148,N_1645,N_293);
xnor U9149 (N_9149,N_105,N_158);
xnor U9150 (N_9150,N_2772,N_3457);
nand U9151 (N_9151,N_4346,N_1811);
xnor U9152 (N_9152,N_4022,N_2341);
nand U9153 (N_9153,N_3542,N_856);
and U9154 (N_9154,N_1842,N_3634);
or U9155 (N_9155,N_690,N_1855);
xor U9156 (N_9156,N_330,N_556);
or U9157 (N_9157,N_2483,N_3785);
xnor U9158 (N_9158,N_1399,N_2366);
nand U9159 (N_9159,N_2072,N_126);
nand U9160 (N_9160,N_2579,N_730);
or U9161 (N_9161,N_2564,N_3830);
nor U9162 (N_9162,N_980,N_3355);
xnor U9163 (N_9163,N_1571,N_204);
nor U9164 (N_9164,N_1118,N_4027);
nand U9165 (N_9165,N_1626,N_164);
xnor U9166 (N_9166,N_1274,N_4047);
and U9167 (N_9167,N_4895,N_2934);
nand U9168 (N_9168,N_2204,N_2000);
and U9169 (N_9169,N_1454,N_2650);
nor U9170 (N_9170,N_2588,N_3595);
xor U9171 (N_9171,N_4877,N_2905);
and U9172 (N_9172,N_1812,N_704);
nand U9173 (N_9173,N_4122,N_1172);
nand U9174 (N_9174,N_4307,N_1932);
nor U9175 (N_9175,N_4981,N_3595);
xnor U9176 (N_9176,N_2913,N_3625);
nor U9177 (N_9177,N_788,N_3612);
nand U9178 (N_9178,N_2384,N_1661);
xor U9179 (N_9179,N_1804,N_2988);
nor U9180 (N_9180,N_3839,N_59);
or U9181 (N_9181,N_4760,N_733);
or U9182 (N_9182,N_3450,N_4087);
and U9183 (N_9183,N_990,N_3401);
nor U9184 (N_9184,N_3057,N_1126);
nor U9185 (N_9185,N_10,N_1490);
xnor U9186 (N_9186,N_790,N_2554);
or U9187 (N_9187,N_1603,N_3305);
xnor U9188 (N_9188,N_344,N_2314);
xnor U9189 (N_9189,N_1703,N_2253);
xnor U9190 (N_9190,N_1296,N_1993);
or U9191 (N_9191,N_104,N_4860);
nand U9192 (N_9192,N_4465,N_4516);
nor U9193 (N_9193,N_3966,N_4199);
or U9194 (N_9194,N_3269,N_2053);
xnor U9195 (N_9195,N_4902,N_810);
and U9196 (N_9196,N_1280,N_4415);
nand U9197 (N_9197,N_3289,N_4274);
nand U9198 (N_9198,N_3907,N_405);
xnor U9199 (N_9199,N_2881,N_89);
nand U9200 (N_9200,N_2684,N_4141);
xnor U9201 (N_9201,N_197,N_4163);
xnor U9202 (N_9202,N_2770,N_3337);
nand U9203 (N_9203,N_2135,N_2472);
xnor U9204 (N_9204,N_448,N_2312);
nand U9205 (N_9205,N_4833,N_1030);
nor U9206 (N_9206,N_1125,N_3211);
and U9207 (N_9207,N_4306,N_4368);
nand U9208 (N_9208,N_4434,N_2842);
nor U9209 (N_9209,N_4402,N_2557);
and U9210 (N_9210,N_1118,N_3592);
xnor U9211 (N_9211,N_4216,N_10);
or U9212 (N_9212,N_772,N_3965);
xor U9213 (N_9213,N_1871,N_3172);
and U9214 (N_9214,N_3373,N_3372);
nor U9215 (N_9215,N_2385,N_1188);
xnor U9216 (N_9216,N_4446,N_4460);
and U9217 (N_9217,N_3585,N_1197);
xor U9218 (N_9218,N_1793,N_3508);
nor U9219 (N_9219,N_2813,N_1704);
or U9220 (N_9220,N_2922,N_4108);
nand U9221 (N_9221,N_2219,N_79);
xnor U9222 (N_9222,N_3835,N_2171);
nand U9223 (N_9223,N_1553,N_922);
nand U9224 (N_9224,N_3114,N_1305);
or U9225 (N_9225,N_1741,N_3126);
nor U9226 (N_9226,N_1181,N_484);
or U9227 (N_9227,N_914,N_2518);
nand U9228 (N_9228,N_2785,N_3968);
nor U9229 (N_9229,N_2392,N_4804);
xor U9230 (N_9230,N_1775,N_3121);
and U9231 (N_9231,N_574,N_899);
nor U9232 (N_9232,N_2431,N_1831);
or U9233 (N_9233,N_2512,N_2726);
nand U9234 (N_9234,N_3196,N_2960);
nor U9235 (N_9235,N_4206,N_4167);
and U9236 (N_9236,N_1818,N_2071);
xnor U9237 (N_9237,N_3961,N_2953);
xor U9238 (N_9238,N_2714,N_4579);
and U9239 (N_9239,N_4883,N_1772);
nor U9240 (N_9240,N_1673,N_3792);
or U9241 (N_9241,N_4655,N_1915);
and U9242 (N_9242,N_2852,N_1968);
nand U9243 (N_9243,N_4279,N_4712);
nor U9244 (N_9244,N_1936,N_4883);
or U9245 (N_9245,N_2451,N_1287);
or U9246 (N_9246,N_2713,N_2871);
or U9247 (N_9247,N_857,N_4677);
nor U9248 (N_9248,N_4866,N_4260);
nand U9249 (N_9249,N_4872,N_605);
and U9250 (N_9250,N_2439,N_549);
or U9251 (N_9251,N_805,N_4811);
and U9252 (N_9252,N_2706,N_4836);
nor U9253 (N_9253,N_2247,N_3317);
nand U9254 (N_9254,N_495,N_3602);
nand U9255 (N_9255,N_341,N_243);
nand U9256 (N_9256,N_400,N_3540);
nand U9257 (N_9257,N_1136,N_51);
and U9258 (N_9258,N_4801,N_3795);
and U9259 (N_9259,N_1742,N_1546);
and U9260 (N_9260,N_1379,N_475);
nor U9261 (N_9261,N_3486,N_1576);
or U9262 (N_9262,N_3789,N_1624);
and U9263 (N_9263,N_1597,N_1395);
xnor U9264 (N_9264,N_2186,N_4770);
nand U9265 (N_9265,N_2554,N_4107);
xnor U9266 (N_9266,N_373,N_3656);
nor U9267 (N_9267,N_2606,N_4062);
nor U9268 (N_9268,N_2605,N_2547);
nand U9269 (N_9269,N_3972,N_4440);
nor U9270 (N_9270,N_4429,N_3206);
nand U9271 (N_9271,N_1680,N_419);
or U9272 (N_9272,N_2390,N_1470);
xnor U9273 (N_9273,N_157,N_1292);
and U9274 (N_9274,N_1381,N_3423);
nor U9275 (N_9275,N_213,N_3801);
xnor U9276 (N_9276,N_3118,N_2727);
nor U9277 (N_9277,N_2961,N_4803);
or U9278 (N_9278,N_4652,N_2088);
and U9279 (N_9279,N_1863,N_296);
nand U9280 (N_9280,N_4842,N_223);
nor U9281 (N_9281,N_3310,N_1331);
nand U9282 (N_9282,N_521,N_2559);
nor U9283 (N_9283,N_1968,N_2459);
or U9284 (N_9284,N_3235,N_2942);
or U9285 (N_9285,N_4584,N_4929);
and U9286 (N_9286,N_4004,N_911);
or U9287 (N_9287,N_4597,N_4921);
nor U9288 (N_9288,N_2290,N_168);
nor U9289 (N_9289,N_2490,N_1541);
xnor U9290 (N_9290,N_2056,N_3563);
nor U9291 (N_9291,N_426,N_581);
xnor U9292 (N_9292,N_4119,N_3993);
nor U9293 (N_9293,N_2058,N_4580);
nor U9294 (N_9294,N_2528,N_1084);
and U9295 (N_9295,N_2851,N_576);
or U9296 (N_9296,N_4992,N_1171);
nor U9297 (N_9297,N_4663,N_2608);
and U9298 (N_9298,N_4616,N_1878);
or U9299 (N_9299,N_700,N_4365);
nand U9300 (N_9300,N_1105,N_1951);
nand U9301 (N_9301,N_2832,N_186);
nor U9302 (N_9302,N_1248,N_4931);
nor U9303 (N_9303,N_1712,N_319);
and U9304 (N_9304,N_4539,N_3168);
xor U9305 (N_9305,N_1509,N_475);
and U9306 (N_9306,N_533,N_4610);
nand U9307 (N_9307,N_1221,N_4401);
or U9308 (N_9308,N_808,N_4758);
nand U9309 (N_9309,N_3793,N_3607);
or U9310 (N_9310,N_1703,N_1194);
xnor U9311 (N_9311,N_1449,N_78);
xor U9312 (N_9312,N_282,N_4004);
or U9313 (N_9313,N_1620,N_4470);
xor U9314 (N_9314,N_2074,N_3989);
nand U9315 (N_9315,N_299,N_4724);
xor U9316 (N_9316,N_969,N_4844);
or U9317 (N_9317,N_2308,N_718);
nand U9318 (N_9318,N_1945,N_1324);
nor U9319 (N_9319,N_3563,N_1139);
xor U9320 (N_9320,N_4079,N_889);
or U9321 (N_9321,N_1529,N_4012);
and U9322 (N_9322,N_274,N_3214);
nor U9323 (N_9323,N_2311,N_3974);
and U9324 (N_9324,N_4825,N_80);
or U9325 (N_9325,N_4169,N_2296);
nand U9326 (N_9326,N_23,N_4290);
and U9327 (N_9327,N_711,N_1395);
or U9328 (N_9328,N_874,N_2564);
and U9329 (N_9329,N_441,N_1146);
and U9330 (N_9330,N_3519,N_400);
or U9331 (N_9331,N_3311,N_4961);
xnor U9332 (N_9332,N_3033,N_1592);
or U9333 (N_9333,N_1464,N_1320);
xnor U9334 (N_9334,N_4807,N_1674);
nor U9335 (N_9335,N_3244,N_3847);
xnor U9336 (N_9336,N_219,N_4961);
xnor U9337 (N_9337,N_1163,N_2239);
and U9338 (N_9338,N_3536,N_795);
and U9339 (N_9339,N_4793,N_4297);
and U9340 (N_9340,N_2813,N_2695);
or U9341 (N_9341,N_3802,N_334);
nor U9342 (N_9342,N_1417,N_2149);
xnor U9343 (N_9343,N_3063,N_178);
nor U9344 (N_9344,N_640,N_825);
nor U9345 (N_9345,N_1323,N_582);
or U9346 (N_9346,N_246,N_390);
and U9347 (N_9347,N_2369,N_663);
xnor U9348 (N_9348,N_2586,N_3913);
nand U9349 (N_9349,N_1254,N_1280);
and U9350 (N_9350,N_3630,N_3638);
and U9351 (N_9351,N_1269,N_603);
and U9352 (N_9352,N_1887,N_3881);
nand U9353 (N_9353,N_3212,N_1460);
nand U9354 (N_9354,N_896,N_2139);
nor U9355 (N_9355,N_579,N_818);
xor U9356 (N_9356,N_2751,N_3444);
and U9357 (N_9357,N_87,N_508);
nor U9358 (N_9358,N_2665,N_3421);
nor U9359 (N_9359,N_4131,N_4637);
nor U9360 (N_9360,N_2155,N_3303);
nand U9361 (N_9361,N_1793,N_581);
nor U9362 (N_9362,N_3545,N_1765);
and U9363 (N_9363,N_4469,N_2635);
or U9364 (N_9364,N_1730,N_964);
or U9365 (N_9365,N_1246,N_2453);
nand U9366 (N_9366,N_3214,N_934);
or U9367 (N_9367,N_652,N_1306);
and U9368 (N_9368,N_2780,N_1999);
xnor U9369 (N_9369,N_2318,N_796);
and U9370 (N_9370,N_3141,N_4931);
nor U9371 (N_9371,N_3377,N_1854);
nand U9372 (N_9372,N_1205,N_3829);
or U9373 (N_9373,N_2528,N_749);
nand U9374 (N_9374,N_3943,N_682);
xor U9375 (N_9375,N_1062,N_830);
xor U9376 (N_9376,N_4654,N_2700);
or U9377 (N_9377,N_3060,N_4701);
nand U9378 (N_9378,N_788,N_4567);
nor U9379 (N_9379,N_588,N_3023);
nand U9380 (N_9380,N_1158,N_3239);
or U9381 (N_9381,N_2810,N_2906);
xnor U9382 (N_9382,N_2888,N_465);
and U9383 (N_9383,N_3480,N_4425);
nand U9384 (N_9384,N_799,N_1580);
xnor U9385 (N_9385,N_1536,N_630);
or U9386 (N_9386,N_1584,N_1175);
nor U9387 (N_9387,N_2807,N_2233);
nand U9388 (N_9388,N_1176,N_2245);
nor U9389 (N_9389,N_2741,N_4002);
nand U9390 (N_9390,N_4782,N_2773);
or U9391 (N_9391,N_2548,N_3954);
xor U9392 (N_9392,N_531,N_2007);
or U9393 (N_9393,N_6,N_2247);
xnor U9394 (N_9394,N_2204,N_95);
or U9395 (N_9395,N_4556,N_1165);
nand U9396 (N_9396,N_4466,N_467);
xnor U9397 (N_9397,N_326,N_3332);
nand U9398 (N_9398,N_3664,N_983);
xnor U9399 (N_9399,N_2451,N_1258);
xor U9400 (N_9400,N_1033,N_4807);
xor U9401 (N_9401,N_3328,N_314);
nand U9402 (N_9402,N_442,N_474);
nand U9403 (N_9403,N_1470,N_4396);
xnor U9404 (N_9404,N_4249,N_3901);
xor U9405 (N_9405,N_4661,N_1878);
or U9406 (N_9406,N_4016,N_3690);
nor U9407 (N_9407,N_4666,N_4211);
and U9408 (N_9408,N_921,N_2190);
or U9409 (N_9409,N_2695,N_1338);
or U9410 (N_9410,N_2665,N_4081);
nand U9411 (N_9411,N_3708,N_4884);
nor U9412 (N_9412,N_3757,N_2267);
nand U9413 (N_9413,N_4214,N_3535);
nand U9414 (N_9414,N_4810,N_4489);
and U9415 (N_9415,N_3581,N_3420);
xor U9416 (N_9416,N_154,N_4924);
or U9417 (N_9417,N_3788,N_1770);
nor U9418 (N_9418,N_2446,N_3488);
or U9419 (N_9419,N_4370,N_2917);
xnor U9420 (N_9420,N_3187,N_2606);
and U9421 (N_9421,N_992,N_3454);
or U9422 (N_9422,N_1261,N_3809);
xnor U9423 (N_9423,N_1158,N_4669);
nor U9424 (N_9424,N_4017,N_956);
xor U9425 (N_9425,N_4515,N_2745);
or U9426 (N_9426,N_877,N_1517);
nor U9427 (N_9427,N_377,N_672);
nor U9428 (N_9428,N_2879,N_3978);
nor U9429 (N_9429,N_716,N_3831);
or U9430 (N_9430,N_4057,N_4468);
nand U9431 (N_9431,N_4278,N_4244);
or U9432 (N_9432,N_4065,N_1733);
nand U9433 (N_9433,N_2374,N_367);
nor U9434 (N_9434,N_631,N_4674);
or U9435 (N_9435,N_3739,N_359);
or U9436 (N_9436,N_4841,N_4101);
and U9437 (N_9437,N_4210,N_3890);
and U9438 (N_9438,N_1382,N_185);
and U9439 (N_9439,N_77,N_2388);
nand U9440 (N_9440,N_1569,N_3606);
and U9441 (N_9441,N_3878,N_4279);
nand U9442 (N_9442,N_2468,N_3570);
nand U9443 (N_9443,N_151,N_3375);
xnor U9444 (N_9444,N_4884,N_189);
xnor U9445 (N_9445,N_2429,N_2655);
xnor U9446 (N_9446,N_2782,N_2957);
or U9447 (N_9447,N_442,N_1334);
xor U9448 (N_9448,N_2631,N_36);
or U9449 (N_9449,N_1551,N_3364);
and U9450 (N_9450,N_4927,N_1544);
xnor U9451 (N_9451,N_4759,N_4403);
nor U9452 (N_9452,N_326,N_1324);
and U9453 (N_9453,N_1842,N_55);
nand U9454 (N_9454,N_931,N_827);
nand U9455 (N_9455,N_4801,N_947);
nand U9456 (N_9456,N_4125,N_4962);
and U9457 (N_9457,N_1387,N_2021);
xor U9458 (N_9458,N_737,N_2133);
and U9459 (N_9459,N_1278,N_44);
nor U9460 (N_9460,N_2031,N_42);
nor U9461 (N_9461,N_2006,N_3958);
and U9462 (N_9462,N_3204,N_2020);
or U9463 (N_9463,N_4935,N_2342);
nor U9464 (N_9464,N_2177,N_3375);
xnor U9465 (N_9465,N_1672,N_4613);
nor U9466 (N_9466,N_4296,N_815);
xor U9467 (N_9467,N_1184,N_4801);
nor U9468 (N_9468,N_4241,N_4487);
nor U9469 (N_9469,N_1350,N_4253);
and U9470 (N_9470,N_446,N_2060);
and U9471 (N_9471,N_4959,N_253);
nor U9472 (N_9472,N_2692,N_4972);
xor U9473 (N_9473,N_3408,N_3660);
nor U9474 (N_9474,N_3376,N_1473);
nor U9475 (N_9475,N_4752,N_266);
xnor U9476 (N_9476,N_1069,N_3144);
nor U9477 (N_9477,N_2705,N_3835);
nor U9478 (N_9478,N_817,N_4059);
or U9479 (N_9479,N_4059,N_3775);
and U9480 (N_9480,N_404,N_2648);
nor U9481 (N_9481,N_3777,N_1823);
nor U9482 (N_9482,N_846,N_4945);
xor U9483 (N_9483,N_705,N_4418);
nor U9484 (N_9484,N_2750,N_918);
or U9485 (N_9485,N_1959,N_4604);
nand U9486 (N_9486,N_4192,N_1026);
and U9487 (N_9487,N_3017,N_488);
or U9488 (N_9488,N_1842,N_3435);
xnor U9489 (N_9489,N_3562,N_2040);
and U9490 (N_9490,N_4857,N_3800);
nor U9491 (N_9491,N_3340,N_316);
and U9492 (N_9492,N_3311,N_523);
nand U9493 (N_9493,N_2053,N_1926);
and U9494 (N_9494,N_4328,N_4049);
or U9495 (N_9495,N_411,N_2467);
and U9496 (N_9496,N_1776,N_247);
nand U9497 (N_9497,N_189,N_259);
xnor U9498 (N_9498,N_100,N_1896);
or U9499 (N_9499,N_3687,N_1228);
and U9500 (N_9500,N_475,N_3598);
nand U9501 (N_9501,N_3265,N_1164);
nor U9502 (N_9502,N_3747,N_940);
xor U9503 (N_9503,N_4844,N_3819);
xnor U9504 (N_9504,N_2878,N_1393);
nand U9505 (N_9505,N_3390,N_3026);
and U9506 (N_9506,N_2491,N_1118);
and U9507 (N_9507,N_799,N_1681);
xnor U9508 (N_9508,N_203,N_1030);
and U9509 (N_9509,N_668,N_2430);
xnor U9510 (N_9510,N_4047,N_749);
xor U9511 (N_9511,N_3546,N_4705);
xnor U9512 (N_9512,N_674,N_3200);
nor U9513 (N_9513,N_4219,N_2431);
and U9514 (N_9514,N_2683,N_4385);
xnor U9515 (N_9515,N_2646,N_3750);
nand U9516 (N_9516,N_4279,N_1389);
and U9517 (N_9517,N_151,N_1906);
xnor U9518 (N_9518,N_3917,N_1971);
or U9519 (N_9519,N_4469,N_3242);
nor U9520 (N_9520,N_1709,N_2207);
xor U9521 (N_9521,N_4845,N_2990);
nand U9522 (N_9522,N_1947,N_370);
nor U9523 (N_9523,N_4951,N_1539);
xor U9524 (N_9524,N_300,N_568);
xnor U9525 (N_9525,N_2378,N_1199);
xor U9526 (N_9526,N_2619,N_249);
nand U9527 (N_9527,N_666,N_3642);
and U9528 (N_9528,N_4322,N_1109);
nor U9529 (N_9529,N_309,N_4579);
or U9530 (N_9530,N_3925,N_121);
and U9531 (N_9531,N_1573,N_1436);
nor U9532 (N_9532,N_1468,N_1224);
nand U9533 (N_9533,N_4408,N_4801);
nand U9534 (N_9534,N_2991,N_1919);
nor U9535 (N_9535,N_2586,N_476);
or U9536 (N_9536,N_826,N_4086);
xor U9537 (N_9537,N_4182,N_716);
nor U9538 (N_9538,N_680,N_2781);
xnor U9539 (N_9539,N_2079,N_2577);
nand U9540 (N_9540,N_4699,N_1862);
nand U9541 (N_9541,N_294,N_2420);
and U9542 (N_9542,N_3868,N_1593);
and U9543 (N_9543,N_1245,N_3122);
and U9544 (N_9544,N_3775,N_1316);
and U9545 (N_9545,N_9,N_409);
nor U9546 (N_9546,N_4791,N_392);
nor U9547 (N_9547,N_2990,N_419);
or U9548 (N_9548,N_2589,N_1904);
and U9549 (N_9549,N_3107,N_1866);
nor U9550 (N_9550,N_2231,N_3528);
or U9551 (N_9551,N_702,N_1727);
or U9552 (N_9552,N_376,N_57);
nand U9553 (N_9553,N_4740,N_2732);
xor U9554 (N_9554,N_32,N_9);
xnor U9555 (N_9555,N_2370,N_3661);
xnor U9556 (N_9556,N_1511,N_1305);
and U9557 (N_9557,N_4357,N_3259);
nand U9558 (N_9558,N_2008,N_3056);
xnor U9559 (N_9559,N_2869,N_57);
nand U9560 (N_9560,N_4108,N_770);
and U9561 (N_9561,N_1189,N_322);
xnor U9562 (N_9562,N_4516,N_2338);
nand U9563 (N_9563,N_2528,N_3478);
and U9564 (N_9564,N_4208,N_1850);
or U9565 (N_9565,N_4784,N_244);
nand U9566 (N_9566,N_4875,N_384);
and U9567 (N_9567,N_3839,N_240);
nor U9568 (N_9568,N_2703,N_2091);
and U9569 (N_9569,N_2049,N_4495);
xnor U9570 (N_9570,N_4323,N_1825);
xor U9571 (N_9571,N_1870,N_1140);
and U9572 (N_9572,N_4904,N_3111);
and U9573 (N_9573,N_4414,N_4919);
or U9574 (N_9574,N_3159,N_3512);
nand U9575 (N_9575,N_2749,N_684);
xor U9576 (N_9576,N_799,N_1411);
or U9577 (N_9577,N_3775,N_2494);
and U9578 (N_9578,N_3442,N_4252);
or U9579 (N_9579,N_2133,N_1572);
and U9580 (N_9580,N_131,N_2030);
and U9581 (N_9581,N_1919,N_403);
nand U9582 (N_9582,N_3858,N_3447);
and U9583 (N_9583,N_4176,N_119);
or U9584 (N_9584,N_3615,N_4681);
or U9585 (N_9585,N_3102,N_1348);
and U9586 (N_9586,N_4236,N_750);
nor U9587 (N_9587,N_1494,N_3749);
and U9588 (N_9588,N_1516,N_4893);
xnor U9589 (N_9589,N_4642,N_899);
or U9590 (N_9590,N_1527,N_1293);
xnor U9591 (N_9591,N_226,N_1199);
and U9592 (N_9592,N_4251,N_2425);
or U9593 (N_9593,N_900,N_4644);
or U9594 (N_9594,N_2132,N_3168);
and U9595 (N_9595,N_2957,N_3827);
and U9596 (N_9596,N_2380,N_1717);
nor U9597 (N_9597,N_3622,N_4876);
xnor U9598 (N_9598,N_4918,N_1668);
xor U9599 (N_9599,N_2432,N_3098);
xnor U9600 (N_9600,N_1936,N_2318);
nor U9601 (N_9601,N_2061,N_1232);
or U9602 (N_9602,N_4393,N_4101);
xnor U9603 (N_9603,N_688,N_832);
nand U9604 (N_9604,N_2921,N_3851);
and U9605 (N_9605,N_3976,N_1501);
xor U9606 (N_9606,N_728,N_65);
and U9607 (N_9607,N_4054,N_2484);
nand U9608 (N_9608,N_1993,N_4752);
xor U9609 (N_9609,N_2934,N_2181);
xor U9610 (N_9610,N_2935,N_1616);
nand U9611 (N_9611,N_3375,N_4428);
and U9612 (N_9612,N_2142,N_2887);
nand U9613 (N_9613,N_3352,N_1987);
and U9614 (N_9614,N_4666,N_1317);
nand U9615 (N_9615,N_2642,N_700);
nor U9616 (N_9616,N_3207,N_518);
xor U9617 (N_9617,N_1714,N_2556);
nand U9618 (N_9618,N_2508,N_387);
nor U9619 (N_9619,N_3669,N_2254);
and U9620 (N_9620,N_1552,N_3331);
nand U9621 (N_9621,N_398,N_2025);
or U9622 (N_9622,N_3372,N_3590);
nand U9623 (N_9623,N_4483,N_4845);
nor U9624 (N_9624,N_2454,N_2907);
xnor U9625 (N_9625,N_2400,N_3730);
nor U9626 (N_9626,N_4188,N_372);
nand U9627 (N_9627,N_2773,N_4834);
or U9628 (N_9628,N_651,N_2681);
nand U9629 (N_9629,N_734,N_3707);
xnor U9630 (N_9630,N_4702,N_4450);
nand U9631 (N_9631,N_3215,N_1883);
nand U9632 (N_9632,N_1750,N_908);
nand U9633 (N_9633,N_3949,N_1193);
or U9634 (N_9634,N_1816,N_3520);
nand U9635 (N_9635,N_1275,N_1291);
nor U9636 (N_9636,N_4115,N_1616);
or U9637 (N_9637,N_1109,N_28);
nand U9638 (N_9638,N_601,N_2122);
nor U9639 (N_9639,N_3423,N_2021);
and U9640 (N_9640,N_4883,N_3015);
nor U9641 (N_9641,N_1434,N_146);
nor U9642 (N_9642,N_471,N_2168);
xor U9643 (N_9643,N_4440,N_2925);
and U9644 (N_9644,N_545,N_3250);
nand U9645 (N_9645,N_375,N_1699);
xnor U9646 (N_9646,N_740,N_4611);
xnor U9647 (N_9647,N_4379,N_2904);
nor U9648 (N_9648,N_4784,N_2830);
and U9649 (N_9649,N_2605,N_2156);
nand U9650 (N_9650,N_1874,N_4954);
nand U9651 (N_9651,N_1522,N_2786);
xnor U9652 (N_9652,N_3583,N_318);
and U9653 (N_9653,N_1211,N_2466);
nand U9654 (N_9654,N_4885,N_691);
nand U9655 (N_9655,N_804,N_2779);
or U9656 (N_9656,N_4974,N_4823);
nand U9657 (N_9657,N_3643,N_3816);
nor U9658 (N_9658,N_4790,N_2195);
and U9659 (N_9659,N_2790,N_4673);
and U9660 (N_9660,N_3578,N_1586);
and U9661 (N_9661,N_4546,N_2197);
nand U9662 (N_9662,N_4588,N_2685);
xor U9663 (N_9663,N_1168,N_965);
xor U9664 (N_9664,N_2467,N_2050);
or U9665 (N_9665,N_229,N_1893);
nand U9666 (N_9666,N_4732,N_97);
nor U9667 (N_9667,N_1781,N_4214);
xor U9668 (N_9668,N_2296,N_2621);
xnor U9669 (N_9669,N_4201,N_1107);
and U9670 (N_9670,N_1374,N_1689);
xnor U9671 (N_9671,N_38,N_1920);
nand U9672 (N_9672,N_1566,N_1018);
and U9673 (N_9673,N_4696,N_2299);
xor U9674 (N_9674,N_229,N_4899);
and U9675 (N_9675,N_475,N_3526);
nand U9676 (N_9676,N_2617,N_2505);
nor U9677 (N_9677,N_4183,N_459);
xnor U9678 (N_9678,N_1249,N_1626);
nand U9679 (N_9679,N_4971,N_2840);
nor U9680 (N_9680,N_3064,N_4228);
nand U9681 (N_9681,N_3114,N_3272);
and U9682 (N_9682,N_4122,N_996);
xnor U9683 (N_9683,N_3644,N_1376);
and U9684 (N_9684,N_1597,N_4202);
and U9685 (N_9685,N_2500,N_253);
or U9686 (N_9686,N_3849,N_1177);
nand U9687 (N_9687,N_2436,N_1956);
or U9688 (N_9688,N_3253,N_1935);
xnor U9689 (N_9689,N_4596,N_2882);
xnor U9690 (N_9690,N_654,N_1819);
or U9691 (N_9691,N_1532,N_2251);
xor U9692 (N_9692,N_4592,N_1377);
or U9693 (N_9693,N_4387,N_3705);
or U9694 (N_9694,N_4285,N_1441);
or U9695 (N_9695,N_1104,N_630);
nor U9696 (N_9696,N_3146,N_3724);
nand U9697 (N_9697,N_320,N_447);
nand U9698 (N_9698,N_2827,N_2246);
xor U9699 (N_9699,N_4271,N_3029);
or U9700 (N_9700,N_1676,N_1243);
and U9701 (N_9701,N_1396,N_59);
nand U9702 (N_9702,N_1766,N_202);
and U9703 (N_9703,N_3483,N_1362);
nand U9704 (N_9704,N_4133,N_2288);
or U9705 (N_9705,N_337,N_3081);
nand U9706 (N_9706,N_2216,N_3229);
nor U9707 (N_9707,N_4810,N_3118);
nand U9708 (N_9708,N_2321,N_4783);
and U9709 (N_9709,N_3858,N_4423);
nor U9710 (N_9710,N_3098,N_1158);
and U9711 (N_9711,N_1708,N_2917);
and U9712 (N_9712,N_4491,N_2614);
nor U9713 (N_9713,N_3674,N_37);
and U9714 (N_9714,N_1403,N_1328);
nor U9715 (N_9715,N_15,N_3238);
and U9716 (N_9716,N_3631,N_2971);
and U9717 (N_9717,N_2329,N_588);
nor U9718 (N_9718,N_252,N_211);
and U9719 (N_9719,N_4154,N_2485);
nor U9720 (N_9720,N_1139,N_2721);
nor U9721 (N_9721,N_2519,N_4796);
nor U9722 (N_9722,N_291,N_4447);
xor U9723 (N_9723,N_4417,N_169);
or U9724 (N_9724,N_1235,N_3064);
or U9725 (N_9725,N_892,N_533);
or U9726 (N_9726,N_1008,N_3325);
xnor U9727 (N_9727,N_2889,N_3580);
xnor U9728 (N_9728,N_3577,N_728);
nand U9729 (N_9729,N_4786,N_2135);
nand U9730 (N_9730,N_4104,N_3535);
xnor U9731 (N_9731,N_4354,N_4818);
or U9732 (N_9732,N_3065,N_12);
and U9733 (N_9733,N_3081,N_4676);
or U9734 (N_9734,N_1161,N_3548);
nor U9735 (N_9735,N_1021,N_1683);
xor U9736 (N_9736,N_4190,N_674);
or U9737 (N_9737,N_807,N_4775);
nand U9738 (N_9738,N_2174,N_2931);
xnor U9739 (N_9739,N_1330,N_1209);
nand U9740 (N_9740,N_4571,N_1040);
and U9741 (N_9741,N_2300,N_2235);
nor U9742 (N_9742,N_492,N_971);
xnor U9743 (N_9743,N_2839,N_125);
xor U9744 (N_9744,N_1469,N_2250);
nor U9745 (N_9745,N_630,N_643);
and U9746 (N_9746,N_3252,N_3730);
or U9747 (N_9747,N_299,N_517);
or U9748 (N_9748,N_2569,N_602);
or U9749 (N_9749,N_1716,N_3522);
xnor U9750 (N_9750,N_2625,N_3952);
nor U9751 (N_9751,N_2239,N_3021);
and U9752 (N_9752,N_150,N_1923);
nor U9753 (N_9753,N_2286,N_3641);
xnor U9754 (N_9754,N_3237,N_2809);
or U9755 (N_9755,N_4701,N_1919);
nand U9756 (N_9756,N_4191,N_315);
and U9757 (N_9757,N_1865,N_4005);
or U9758 (N_9758,N_1032,N_2518);
nor U9759 (N_9759,N_3591,N_2600);
nor U9760 (N_9760,N_3648,N_2941);
nor U9761 (N_9761,N_185,N_4703);
xnor U9762 (N_9762,N_771,N_3288);
nand U9763 (N_9763,N_637,N_3046);
and U9764 (N_9764,N_2671,N_1034);
or U9765 (N_9765,N_1450,N_3720);
xnor U9766 (N_9766,N_3502,N_4879);
xnor U9767 (N_9767,N_802,N_4808);
xnor U9768 (N_9768,N_1824,N_3518);
xor U9769 (N_9769,N_3518,N_3543);
nand U9770 (N_9770,N_3557,N_4808);
or U9771 (N_9771,N_4992,N_3566);
or U9772 (N_9772,N_3467,N_545);
and U9773 (N_9773,N_591,N_3426);
and U9774 (N_9774,N_3172,N_1137);
nor U9775 (N_9775,N_747,N_1830);
nor U9776 (N_9776,N_152,N_2428);
nand U9777 (N_9777,N_1816,N_2792);
xnor U9778 (N_9778,N_4762,N_1940);
and U9779 (N_9779,N_1633,N_65);
xnor U9780 (N_9780,N_2898,N_3169);
or U9781 (N_9781,N_1225,N_4595);
and U9782 (N_9782,N_4587,N_4675);
and U9783 (N_9783,N_152,N_4054);
nor U9784 (N_9784,N_2199,N_1643);
or U9785 (N_9785,N_539,N_655);
or U9786 (N_9786,N_1850,N_1754);
and U9787 (N_9787,N_2671,N_2728);
nor U9788 (N_9788,N_3015,N_2982);
nand U9789 (N_9789,N_1779,N_4245);
xor U9790 (N_9790,N_1503,N_2597);
xnor U9791 (N_9791,N_1062,N_4109);
nor U9792 (N_9792,N_2375,N_2071);
nor U9793 (N_9793,N_3976,N_3171);
and U9794 (N_9794,N_3513,N_250);
xnor U9795 (N_9795,N_2793,N_1550);
or U9796 (N_9796,N_2050,N_4804);
and U9797 (N_9797,N_3107,N_1208);
xnor U9798 (N_9798,N_4754,N_1515);
xnor U9799 (N_9799,N_27,N_4968);
nand U9800 (N_9800,N_263,N_3761);
nor U9801 (N_9801,N_1244,N_4431);
xnor U9802 (N_9802,N_1914,N_4974);
xor U9803 (N_9803,N_2175,N_4056);
xor U9804 (N_9804,N_3129,N_4622);
or U9805 (N_9805,N_4190,N_581);
nand U9806 (N_9806,N_1629,N_4355);
xnor U9807 (N_9807,N_249,N_840);
nor U9808 (N_9808,N_3062,N_620);
and U9809 (N_9809,N_4136,N_4479);
xor U9810 (N_9810,N_1053,N_3001);
or U9811 (N_9811,N_4720,N_2174);
or U9812 (N_9812,N_1058,N_1613);
xor U9813 (N_9813,N_1015,N_2217);
and U9814 (N_9814,N_2207,N_1788);
and U9815 (N_9815,N_2133,N_4797);
nand U9816 (N_9816,N_224,N_3322);
or U9817 (N_9817,N_1386,N_356);
and U9818 (N_9818,N_3852,N_1920);
and U9819 (N_9819,N_1158,N_4060);
xnor U9820 (N_9820,N_1091,N_4174);
and U9821 (N_9821,N_723,N_1893);
and U9822 (N_9822,N_1386,N_588);
or U9823 (N_9823,N_3009,N_3358);
or U9824 (N_9824,N_359,N_891);
and U9825 (N_9825,N_3993,N_951);
or U9826 (N_9826,N_1711,N_4228);
nand U9827 (N_9827,N_2525,N_1906);
nor U9828 (N_9828,N_4159,N_2748);
xor U9829 (N_9829,N_4391,N_1798);
nand U9830 (N_9830,N_1717,N_4447);
xor U9831 (N_9831,N_3520,N_2914);
nand U9832 (N_9832,N_501,N_3794);
or U9833 (N_9833,N_288,N_3638);
xnor U9834 (N_9834,N_4216,N_4130);
and U9835 (N_9835,N_3852,N_4021);
nor U9836 (N_9836,N_244,N_3803);
nand U9837 (N_9837,N_1314,N_1947);
and U9838 (N_9838,N_2429,N_1431);
nor U9839 (N_9839,N_1621,N_3303);
or U9840 (N_9840,N_4844,N_428);
nand U9841 (N_9841,N_3464,N_4010);
and U9842 (N_9842,N_3487,N_4561);
or U9843 (N_9843,N_2074,N_2687);
nor U9844 (N_9844,N_3775,N_3967);
xnor U9845 (N_9845,N_2026,N_2371);
nor U9846 (N_9846,N_4274,N_2592);
nand U9847 (N_9847,N_2949,N_2385);
or U9848 (N_9848,N_2508,N_4838);
nand U9849 (N_9849,N_1476,N_4026);
xor U9850 (N_9850,N_2054,N_858);
or U9851 (N_9851,N_3604,N_1354);
or U9852 (N_9852,N_4888,N_4655);
nand U9853 (N_9853,N_2556,N_3442);
and U9854 (N_9854,N_85,N_4188);
or U9855 (N_9855,N_3846,N_587);
nand U9856 (N_9856,N_4248,N_2058);
xor U9857 (N_9857,N_3959,N_135);
or U9858 (N_9858,N_1693,N_4544);
nor U9859 (N_9859,N_38,N_236);
nor U9860 (N_9860,N_2779,N_878);
nand U9861 (N_9861,N_4211,N_1616);
nor U9862 (N_9862,N_4551,N_976);
xor U9863 (N_9863,N_2858,N_1628);
nor U9864 (N_9864,N_2290,N_2880);
xnor U9865 (N_9865,N_1798,N_1049);
and U9866 (N_9866,N_1445,N_1562);
or U9867 (N_9867,N_3706,N_570);
or U9868 (N_9868,N_3467,N_1893);
xor U9869 (N_9869,N_598,N_3904);
nor U9870 (N_9870,N_3973,N_4068);
xnor U9871 (N_9871,N_2036,N_2580);
nor U9872 (N_9872,N_2007,N_1705);
and U9873 (N_9873,N_391,N_2069);
and U9874 (N_9874,N_863,N_673);
xnor U9875 (N_9875,N_3728,N_1414);
nor U9876 (N_9876,N_1634,N_1726);
or U9877 (N_9877,N_194,N_1561);
nand U9878 (N_9878,N_235,N_4910);
or U9879 (N_9879,N_4278,N_4001);
nand U9880 (N_9880,N_1078,N_1004);
xnor U9881 (N_9881,N_2120,N_4249);
nor U9882 (N_9882,N_4650,N_4991);
or U9883 (N_9883,N_2977,N_1925);
nor U9884 (N_9884,N_1765,N_1297);
xnor U9885 (N_9885,N_718,N_1120);
or U9886 (N_9886,N_2170,N_4425);
or U9887 (N_9887,N_2429,N_1473);
nand U9888 (N_9888,N_4532,N_200);
or U9889 (N_9889,N_4276,N_1267);
or U9890 (N_9890,N_2729,N_1728);
nor U9891 (N_9891,N_284,N_1106);
nand U9892 (N_9892,N_1910,N_122);
and U9893 (N_9893,N_249,N_1018);
nor U9894 (N_9894,N_4166,N_1616);
xnor U9895 (N_9895,N_3829,N_3645);
and U9896 (N_9896,N_1202,N_1574);
or U9897 (N_9897,N_1545,N_2685);
and U9898 (N_9898,N_114,N_126);
or U9899 (N_9899,N_4388,N_2491);
nor U9900 (N_9900,N_4641,N_1578);
xor U9901 (N_9901,N_3905,N_1460);
nand U9902 (N_9902,N_2482,N_4608);
or U9903 (N_9903,N_3293,N_1397);
nor U9904 (N_9904,N_1600,N_3529);
xor U9905 (N_9905,N_2456,N_2410);
nand U9906 (N_9906,N_2197,N_4838);
or U9907 (N_9907,N_4023,N_795);
and U9908 (N_9908,N_2476,N_4333);
and U9909 (N_9909,N_2352,N_2345);
nor U9910 (N_9910,N_1688,N_3046);
nor U9911 (N_9911,N_2721,N_284);
xor U9912 (N_9912,N_1558,N_4233);
nand U9913 (N_9913,N_998,N_658);
nor U9914 (N_9914,N_4738,N_3566);
nand U9915 (N_9915,N_2159,N_4108);
nand U9916 (N_9916,N_1721,N_4452);
xnor U9917 (N_9917,N_409,N_4848);
and U9918 (N_9918,N_4888,N_4767);
nand U9919 (N_9919,N_3760,N_399);
and U9920 (N_9920,N_2463,N_278);
xor U9921 (N_9921,N_1,N_3449);
and U9922 (N_9922,N_4226,N_2149);
or U9923 (N_9923,N_2273,N_685);
or U9924 (N_9924,N_2805,N_3243);
and U9925 (N_9925,N_2470,N_3785);
and U9926 (N_9926,N_2182,N_4993);
nand U9927 (N_9927,N_4295,N_1342);
nor U9928 (N_9928,N_4283,N_2788);
nor U9929 (N_9929,N_375,N_2402);
nand U9930 (N_9930,N_2352,N_564);
nor U9931 (N_9931,N_1771,N_4270);
nor U9932 (N_9932,N_129,N_2112);
nand U9933 (N_9933,N_1855,N_1010);
nand U9934 (N_9934,N_4826,N_2250);
or U9935 (N_9935,N_4397,N_1955);
and U9936 (N_9936,N_4329,N_4731);
nor U9937 (N_9937,N_1866,N_2341);
nand U9938 (N_9938,N_4520,N_728);
xor U9939 (N_9939,N_4999,N_1057);
nor U9940 (N_9940,N_3723,N_1254);
nand U9941 (N_9941,N_877,N_669);
nor U9942 (N_9942,N_4883,N_2256);
and U9943 (N_9943,N_4838,N_2076);
or U9944 (N_9944,N_4308,N_742);
xor U9945 (N_9945,N_4200,N_2304);
or U9946 (N_9946,N_1873,N_4544);
nand U9947 (N_9947,N_252,N_3393);
nand U9948 (N_9948,N_1388,N_3735);
or U9949 (N_9949,N_3778,N_4118);
nand U9950 (N_9950,N_4148,N_818);
xor U9951 (N_9951,N_3424,N_3929);
xnor U9952 (N_9952,N_1164,N_2780);
xor U9953 (N_9953,N_2362,N_4278);
and U9954 (N_9954,N_2299,N_4580);
and U9955 (N_9955,N_3487,N_2589);
and U9956 (N_9956,N_4865,N_3828);
or U9957 (N_9957,N_2687,N_3272);
and U9958 (N_9958,N_3304,N_2555);
and U9959 (N_9959,N_3170,N_1513);
nor U9960 (N_9960,N_3464,N_3139);
nand U9961 (N_9961,N_4165,N_3769);
nor U9962 (N_9962,N_491,N_3135);
xor U9963 (N_9963,N_4162,N_3756);
nand U9964 (N_9964,N_3449,N_3451);
and U9965 (N_9965,N_4233,N_4490);
and U9966 (N_9966,N_2402,N_11);
or U9967 (N_9967,N_1361,N_2889);
nand U9968 (N_9968,N_309,N_4761);
and U9969 (N_9969,N_1023,N_4332);
and U9970 (N_9970,N_3857,N_4461);
nor U9971 (N_9971,N_2289,N_975);
xor U9972 (N_9972,N_2972,N_4935);
and U9973 (N_9973,N_2979,N_1721);
xnor U9974 (N_9974,N_241,N_338);
nor U9975 (N_9975,N_3451,N_3277);
nand U9976 (N_9976,N_1594,N_2705);
and U9977 (N_9977,N_1142,N_4232);
or U9978 (N_9978,N_2163,N_1360);
xnor U9979 (N_9979,N_2092,N_1459);
nand U9980 (N_9980,N_679,N_1712);
and U9981 (N_9981,N_3374,N_3794);
or U9982 (N_9982,N_3943,N_1719);
xnor U9983 (N_9983,N_3138,N_4952);
xnor U9984 (N_9984,N_3939,N_4764);
and U9985 (N_9985,N_1977,N_1045);
nor U9986 (N_9986,N_4707,N_422);
and U9987 (N_9987,N_1944,N_1004);
and U9988 (N_9988,N_666,N_551);
and U9989 (N_9989,N_3138,N_344);
nor U9990 (N_9990,N_2026,N_3952);
xnor U9991 (N_9991,N_875,N_3713);
nor U9992 (N_9992,N_1911,N_318);
xnor U9993 (N_9993,N_3405,N_2870);
nand U9994 (N_9994,N_3577,N_2333);
nor U9995 (N_9995,N_2916,N_375);
and U9996 (N_9996,N_4817,N_3071);
or U9997 (N_9997,N_4578,N_4568);
nand U9998 (N_9998,N_3154,N_2801);
nand U9999 (N_9999,N_883,N_423);
and U10000 (N_10000,N_7985,N_9151);
nand U10001 (N_10001,N_5221,N_6078);
nand U10002 (N_10002,N_8965,N_9583);
nand U10003 (N_10003,N_8624,N_6769);
and U10004 (N_10004,N_5954,N_6452);
and U10005 (N_10005,N_6791,N_7339);
nor U10006 (N_10006,N_6060,N_7751);
nand U10007 (N_10007,N_5302,N_5290);
and U10008 (N_10008,N_7872,N_9341);
nand U10009 (N_10009,N_9187,N_8815);
nand U10010 (N_10010,N_9765,N_5627);
nand U10011 (N_10011,N_8614,N_6351);
or U10012 (N_10012,N_8490,N_9854);
xnor U10013 (N_10013,N_8521,N_7785);
and U10014 (N_10014,N_5557,N_6873);
nor U10015 (N_10015,N_6957,N_8399);
and U10016 (N_10016,N_6359,N_9822);
xor U10017 (N_10017,N_6937,N_5875);
or U10018 (N_10018,N_6729,N_5502);
nor U10019 (N_10019,N_5842,N_7773);
nand U10020 (N_10020,N_9381,N_8658);
nor U10021 (N_10021,N_5069,N_7114);
and U10022 (N_10022,N_6991,N_7035);
and U10023 (N_10023,N_8685,N_6635);
or U10024 (N_10024,N_9928,N_5346);
nand U10025 (N_10025,N_5908,N_9336);
xor U10026 (N_10026,N_8319,N_6542);
or U10027 (N_10027,N_7240,N_6698);
and U10028 (N_10028,N_9374,N_8651);
xnor U10029 (N_10029,N_8394,N_9299);
xnor U10030 (N_10030,N_9937,N_5227);
nand U10031 (N_10031,N_8453,N_8713);
nor U10032 (N_10032,N_6165,N_6960);
nand U10033 (N_10033,N_6712,N_5930);
nor U10034 (N_10034,N_7253,N_8751);
nand U10035 (N_10035,N_5417,N_9490);
xnor U10036 (N_10036,N_8058,N_7653);
xor U10037 (N_10037,N_5085,N_7798);
or U10038 (N_10038,N_6963,N_6909);
nor U10039 (N_10039,N_8491,N_7198);
or U10040 (N_10040,N_6074,N_6915);
nand U10041 (N_10041,N_5402,N_5165);
xnor U10042 (N_10042,N_8725,N_5688);
nor U10043 (N_10043,N_5988,N_9392);
or U10044 (N_10044,N_8062,N_8020);
and U10045 (N_10045,N_7536,N_7405);
xor U10046 (N_10046,N_8832,N_9575);
and U10047 (N_10047,N_8083,N_8695);
xnor U10048 (N_10048,N_6996,N_5642);
xor U10049 (N_10049,N_5824,N_7953);
and U10050 (N_10050,N_5549,N_7584);
and U10051 (N_10051,N_7874,N_6867);
and U10052 (N_10052,N_6150,N_9723);
nor U10053 (N_10053,N_8530,N_5255);
and U10054 (N_10054,N_8137,N_7732);
nand U10055 (N_10055,N_5683,N_6715);
and U10056 (N_10056,N_5952,N_5163);
nand U10057 (N_10057,N_6825,N_7166);
xor U10058 (N_10058,N_9206,N_8424);
or U10059 (N_10059,N_7999,N_9538);
and U10060 (N_10060,N_9785,N_8865);
nand U10061 (N_10061,N_7682,N_9165);
nand U10062 (N_10062,N_7337,N_6953);
nand U10063 (N_10063,N_5127,N_6718);
nor U10064 (N_10064,N_9791,N_6749);
or U10065 (N_10065,N_5115,N_5919);
xnor U10066 (N_10066,N_5006,N_9088);
xor U10067 (N_10067,N_9640,N_8148);
and U10068 (N_10068,N_5041,N_7412);
nand U10069 (N_10069,N_8379,N_5641);
and U10070 (N_10070,N_5409,N_5825);
nor U10071 (N_10071,N_9933,N_8668);
xor U10072 (N_10072,N_6246,N_7576);
xnor U10073 (N_10073,N_9498,N_6231);
or U10074 (N_10074,N_5288,N_8561);
nor U10075 (N_10075,N_8580,N_6869);
nand U10076 (N_10076,N_8452,N_7467);
nand U10077 (N_10077,N_8056,N_8544);
and U10078 (N_10078,N_8267,N_8712);
nor U10079 (N_10079,N_9115,N_9186);
or U10080 (N_10080,N_9922,N_6018);
or U10081 (N_10081,N_6551,N_6198);
nor U10082 (N_10082,N_8134,N_9063);
and U10083 (N_10083,N_8364,N_5796);
and U10084 (N_10084,N_9805,N_7525);
nand U10085 (N_10085,N_5622,N_5379);
and U10086 (N_10086,N_6031,N_8564);
and U10087 (N_10087,N_9740,N_6586);
xor U10088 (N_10088,N_9462,N_9105);
and U10089 (N_10089,N_8735,N_7714);
nand U10090 (N_10090,N_8207,N_7028);
and U10091 (N_10091,N_5845,N_8920);
and U10092 (N_10092,N_5631,N_5092);
or U10093 (N_10093,N_8075,N_7251);
nor U10094 (N_10094,N_9830,N_7976);
xor U10095 (N_10095,N_9265,N_5084);
and U10096 (N_10096,N_8155,N_7709);
xor U10097 (N_10097,N_8680,N_7772);
and U10098 (N_10098,N_5305,N_7776);
nor U10099 (N_10099,N_5701,N_7876);
and U10100 (N_10100,N_6591,N_7054);
or U10101 (N_10101,N_8940,N_6990);
nand U10102 (N_10102,N_5687,N_8114);
xnor U10103 (N_10103,N_7242,N_6888);
xor U10104 (N_10104,N_5582,N_5510);
nor U10105 (N_10105,N_9434,N_9215);
or U10106 (N_10106,N_9935,N_5038);
and U10107 (N_10107,N_6977,N_9620);
xnor U10108 (N_10108,N_8604,N_6259);
xnor U10109 (N_10109,N_6904,N_5148);
nor U10110 (N_10110,N_7185,N_6041);
and U10111 (N_10111,N_9636,N_5174);
nor U10112 (N_10112,N_7688,N_7571);
and U10113 (N_10113,N_9261,N_5937);
or U10114 (N_10114,N_8791,N_8851);
and U10115 (N_10115,N_8605,N_9623);
and U10116 (N_10116,N_8288,N_6035);
or U10117 (N_10117,N_5414,N_9309);
nand U10118 (N_10118,N_8859,N_7851);
nor U10119 (N_10119,N_7012,N_7582);
nand U10120 (N_10120,N_7239,N_5061);
xor U10121 (N_10121,N_9222,N_9015);
nand U10122 (N_10122,N_9611,N_8444);
xnor U10123 (N_10123,N_7205,N_8099);
xor U10124 (N_10124,N_9470,N_6308);
nor U10125 (N_10125,N_7159,N_5261);
xnor U10126 (N_10126,N_5134,N_7015);
or U10127 (N_10127,N_6810,N_7188);
nor U10128 (N_10128,N_6249,N_8172);
nand U10129 (N_10129,N_9851,N_8887);
and U10130 (N_10130,N_5124,N_6085);
xnor U10131 (N_10131,N_9317,N_8100);
nor U10132 (N_10132,N_8138,N_9170);
or U10133 (N_10133,N_8807,N_5511);
xor U10134 (N_10134,N_8919,N_8915);
xnor U10135 (N_10135,N_7706,N_7244);
xnor U10136 (N_10136,N_7445,N_8958);
nand U10137 (N_10137,N_5287,N_6263);
or U10138 (N_10138,N_5435,N_6084);
and U10139 (N_10139,N_6483,N_9437);
nor U10140 (N_10140,N_7098,N_9752);
and U10141 (N_10141,N_8697,N_7712);
and U10142 (N_10142,N_8290,N_5434);
xor U10143 (N_10143,N_9993,N_6558);
and U10144 (N_10144,N_5050,N_7138);
nand U10145 (N_10145,N_6264,N_5334);
nand U10146 (N_10146,N_6874,N_9012);
xnor U10147 (N_10147,N_5349,N_8875);
nor U10148 (N_10148,N_6570,N_5877);
nor U10149 (N_10149,N_7115,N_9534);
xor U10150 (N_10150,N_8526,N_8672);
nand U10151 (N_10151,N_7025,N_7089);
nor U10152 (N_10152,N_8009,N_5487);
or U10153 (N_10153,N_6132,N_9913);
nand U10154 (N_10154,N_8086,N_8271);
nand U10155 (N_10155,N_7447,N_9714);
or U10156 (N_10156,N_5560,N_5230);
and U10157 (N_10157,N_5076,N_6242);
nor U10158 (N_10158,N_7270,N_6390);
and U10159 (N_10159,N_7905,N_6076);
nor U10160 (N_10160,N_7094,N_9986);
nor U10161 (N_10161,N_5772,N_5843);
and U10162 (N_10162,N_7863,N_8185);
or U10163 (N_10163,N_8700,N_5633);
and U10164 (N_10164,N_8819,N_5602);
nor U10165 (N_10165,N_9590,N_5141);
xnor U10166 (N_10166,N_8511,N_8592);
or U10167 (N_10167,N_6235,N_7116);
and U10168 (N_10168,N_5586,N_7379);
xor U10169 (N_10169,N_8142,N_9720);
xnor U10170 (N_10170,N_8397,N_8664);
nand U10171 (N_10171,N_7814,N_5566);
xor U10172 (N_10172,N_5516,N_5961);
and U10173 (N_10173,N_9258,N_6208);
and U10174 (N_10174,N_6890,N_8782);
or U10175 (N_10175,N_7972,N_8077);
nand U10176 (N_10176,N_6830,N_7321);
or U10177 (N_10177,N_7430,N_8659);
nor U10178 (N_10178,N_6329,N_5425);
and U10179 (N_10179,N_7333,N_9248);
and U10180 (N_10180,N_6152,N_6145);
nand U10181 (N_10181,N_9756,N_5581);
nor U10182 (N_10182,N_5430,N_7127);
xnor U10183 (N_10183,N_5292,N_7649);
and U10184 (N_10184,N_9333,N_8903);
xnor U10185 (N_10185,N_7520,N_6181);
and U10186 (N_10186,N_5541,N_7804);
or U10187 (N_10187,N_6632,N_7928);
and U10188 (N_10188,N_8494,N_9990);
xnor U10189 (N_10189,N_6357,N_8060);
nand U10190 (N_10190,N_6600,N_7501);
nand U10191 (N_10191,N_9728,N_7125);
xor U10192 (N_10192,N_7550,N_5972);
xnor U10193 (N_10193,N_5544,N_6614);
and U10194 (N_10194,N_5555,N_8006);
xnor U10195 (N_10195,N_9451,N_8415);
nand U10196 (N_10196,N_7671,N_5059);
nor U10197 (N_10197,N_5568,N_9008);
xor U10198 (N_10198,N_9754,N_5012);
nand U10199 (N_10199,N_5389,N_9069);
xor U10200 (N_10200,N_9262,N_9831);
and U10201 (N_10201,N_8677,N_7782);
xor U10202 (N_10202,N_6553,N_6330);
nor U10203 (N_10203,N_5691,N_9410);
or U10204 (N_10204,N_5597,N_8775);
and U10205 (N_10205,N_9995,N_8902);
nand U10206 (N_10206,N_5104,N_5486);
nor U10207 (N_10207,N_8322,N_9563);
and U10208 (N_10208,N_5337,N_6428);
and U10209 (N_10209,N_5032,N_8844);
xor U10210 (N_10210,N_8373,N_7858);
nor U10211 (N_10211,N_8046,N_5672);
nor U10212 (N_10212,N_8089,N_7900);
nand U10213 (N_10213,N_6244,N_8690);
nor U10214 (N_10214,N_6625,N_7055);
xnor U10215 (N_10215,N_7901,N_6640);
and U10216 (N_10216,N_9251,N_9887);
nor U10217 (N_10217,N_7859,N_5376);
and U10218 (N_10218,N_8302,N_8527);
or U10219 (N_10219,N_9766,N_6500);
or U10220 (N_10220,N_7064,N_8554);
nand U10221 (N_10221,N_6101,N_8079);
or U10222 (N_10222,N_7091,N_7764);
nand U10223 (N_10223,N_7439,N_7508);
or U10224 (N_10224,N_7606,N_6194);
xor U10225 (N_10225,N_7005,N_6803);
or U10226 (N_10226,N_7562,N_9607);
nand U10227 (N_10227,N_7493,N_5780);
nand U10228 (N_10228,N_6684,N_5956);
nor U10229 (N_10229,N_7314,N_5262);
xor U10230 (N_10230,N_9696,N_7986);
xnor U10231 (N_10231,N_6216,N_9874);
nor U10232 (N_10232,N_9709,N_5538);
and U10233 (N_10233,N_9896,N_7518);
and U10234 (N_10234,N_8929,N_6938);
nand U10235 (N_10235,N_9014,N_7462);
or U10236 (N_10236,N_6106,N_5917);
or U10237 (N_10237,N_7331,N_6462);
and U10238 (N_10238,N_8716,N_5596);
or U10239 (N_10239,N_7450,N_6849);
nor U10240 (N_10240,N_7301,N_7631);
or U10241 (N_10241,N_6276,N_6789);
and U10242 (N_10242,N_6405,N_8800);
xnor U10243 (N_10243,N_9485,N_7008);
or U10244 (N_10244,N_8626,N_9362);
nor U10245 (N_10245,N_9037,N_8538);
nand U10246 (N_10246,N_9814,N_8729);
nor U10247 (N_10247,N_9919,N_6742);
nor U10248 (N_10248,N_6136,N_8970);
nor U10249 (N_10249,N_7601,N_5240);
nand U10250 (N_10250,N_8771,N_8840);
nor U10251 (N_10251,N_8565,N_7715);
or U10252 (N_10252,N_6641,N_7415);
nand U10253 (N_10253,N_6782,N_9673);
nor U10254 (N_10254,N_9264,N_7200);
xor U10255 (N_10255,N_7963,N_9983);
nand U10256 (N_10256,N_6660,N_9132);
nand U10257 (N_10257,N_7130,N_8434);
nand U10258 (N_10258,N_7749,N_6797);
nor U10259 (N_10259,N_7598,N_9006);
nor U10260 (N_10260,N_7970,N_5542);
nor U10261 (N_10261,N_5997,N_9135);
or U10262 (N_10262,N_8125,N_8553);
and U10263 (N_10263,N_8124,N_8646);
and U10264 (N_10264,N_7647,N_7800);
xor U10265 (N_10265,N_9395,N_5836);
xor U10266 (N_10266,N_7592,N_7474);
nor U10267 (N_10267,N_8351,N_9904);
and U10268 (N_10268,N_6111,N_6653);
and U10269 (N_10269,N_8837,N_5680);
or U10270 (N_10270,N_6372,N_5439);
nand U10271 (N_10271,N_9349,N_9196);
nand U10272 (N_10272,N_7209,N_6627);
nor U10273 (N_10273,N_8590,N_7983);
nand U10274 (N_10274,N_5598,N_9554);
nor U10275 (N_10275,N_7787,N_7288);
or U10276 (N_10276,N_6439,N_8641);
or U10277 (N_10277,N_7622,N_6342);
xnor U10278 (N_10278,N_8978,N_8528);
or U10279 (N_10279,N_9188,N_9256);
nor U10280 (N_10280,N_6967,N_9301);
xnor U10281 (N_10281,N_5013,N_9096);
nor U10282 (N_10282,N_7716,N_6796);
and U10283 (N_10283,N_8231,N_7875);
and U10284 (N_10284,N_8779,N_7665);
xor U10285 (N_10285,N_7805,N_6793);
or U10286 (N_10286,N_5556,N_9059);
nor U10287 (N_10287,N_9289,N_7882);
and U10288 (N_10288,N_5120,N_5738);
nor U10289 (N_10289,N_6995,N_8310);
or U10290 (N_10290,N_5847,N_8756);
or U10291 (N_10291,N_7980,N_5018);
or U10292 (N_10292,N_5411,N_9963);
and U10293 (N_10293,N_7925,N_8248);
or U10294 (N_10294,N_9079,N_5767);
xor U10295 (N_10295,N_9284,N_7173);
or U10296 (N_10296,N_9227,N_7548);
and U10297 (N_10297,N_8684,N_6328);
nand U10298 (N_10298,N_7762,N_7401);
and U10299 (N_10299,N_7663,N_7384);
nand U10300 (N_10300,N_9394,N_6839);
xor U10301 (N_10301,N_9164,N_6391);
xnor U10302 (N_10302,N_6532,N_6549);
nand U10303 (N_10303,N_6057,N_6155);
or U10304 (N_10304,N_8295,N_9131);
nor U10305 (N_10305,N_5397,N_6817);
xnor U10306 (N_10306,N_8662,N_8213);
nand U10307 (N_10307,N_8469,N_8571);
or U10308 (N_10308,N_8010,N_9357);
nand U10309 (N_10309,N_8164,N_9544);
nand U10310 (N_10310,N_6138,N_8316);
nor U10311 (N_10311,N_9414,N_6190);
nand U10312 (N_10312,N_6788,N_9890);
nand U10313 (N_10313,N_9236,N_8132);
or U10314 (N_10314,N_7477,N_9587);
and U10315 (N_10315,N_7561,N_7616);
nand U10316 (N_10316,N_8067,N_5437);
nand U10317 (N_10317,N_5565,N_5388);
nor U10318 (N_10318,N_9457,N_9405);
nand U10319 (N_10319,N_7659,N_5238);
or U10320 (N_10320,N_8686,N_5294);
and U10321 (N_10321,N_9139,N_5746);
or U10322 (N_10322,N_7319,N_8917);
nand U10323 (N_10323,N_5870,N_9029);
or U10324 (N_10324,N_6802,N_7527);
nand U10325 (N_10325,N_9898,N_9824);
xor U10326 (N_10326,N_8471,N_6571);
and U10327 (N_10327,N_7388,N_7009);
xor U10328 (N_10328,N_9936,N_6153);
xnor U10329 (N_10329,N_9124,N_5995);
nor U10330 (N_10330,N_5599,N_6255);
or U10331 (N_10331,N_9199,N_5743);
nand U10332 (N_10332,N_9569,N_6747);
xnor U10333 (N_10333,N_7848,N_5123);
and U10334 (N_10334,N_7498,N_8273);
and U10335 (N_10335,N_7552,N_9427);
and U10336 (N_10336,N_7394,N_9578);
nand U10337 (N_10337,N_5193,N_7846);
nor U10338 (N_10338,N_5770,N_7074);
nand U10339 (N_10339,N_7190,N_8694);
and U10340 (N_10340,N_8476,N_7034);
and U10341 (N_10341,N_6238,N_9409);
xnor U10342 (N_10342,N_5694,N_5953);
or U10343 (N_10343,N_8082,N_9425);
or U10344 (N_10344,N_6936,N_7162);
nand U10345 (N_10345,N_7750,N_9297);
or U10346 (N_10346,N_8219,N_6082);
nand U10347 (N_10347,N_5206,N_8296);
or U10348 (N_10348,N_6576,N_8532);
or U10349 (N_10349,N_5635,N_7690);
xnor U10350 (N_10350,N_8904,N_8555);
or U10351 (N_10351,N_5257,N_8964);
nand U10352 (N_10352,N_6575,N_8894);
xnor U10353 (N_10353,N_5045,N_7057);
or U10354 (N_10354,N_6119,N_6232);
nor U10355 (N_10355,N_7014,N_6603);
nor U10356 (N_10356,N_5938,N_9126);
nor U10357 (N_10357,N_8939,N_5777);
xnor U10358 (N_10358,N_9158,N_5390);
xor U10359 (N_10359,N_6363,N_6606);
xor U10360 (N_10360,N_8161,N_9643);
or U10361 (N_10361,N_8938,N_7155);
nor U10362 (N_10362,N_6702,N_9651);
nand U10363 (N_10363,N_5501,N_7408);
or U10364 (N_10364,N_9504,N_8353);
xor U10365 (N_10365,N_9976,N_7457);
nor U10366 (N_10366,N_5518,N_9250);
nand U10367 (N_10367,N_8040,N_7791);
or U10368 (N_10368,N_9960,N_7026);
nand U10369 (N_10369,N_9351,N_9802);
nor U10370 (N_10370,N_5705,N_9171);
nor U10371 (N_10371,N_9924,N_8843);
nand U10372 (N_10372,N_5569,N_8933);
xnor U10373 (N_10373,N_7753,N_6827);
and U10374 (N_10374,N_6555,N_5601);
nor U10375 (N_10375,N_5293,N_9618);
xnor U10376 (N_10376,N_7304,N_6294);
and U10377 (N_10377,N_7556,N_9859);
nor U10378 (N_10378,N_6666,N_9323);
xnor U10379 (N_10379,N_5204,N_9827);
or U10380 (N_10380,N_9017,N_5583);
nand U10381 (N_10381,N_5177,N_9305);
or U10382 (N_10382,N_5657,N_9524);
or U10383 (N_10383,N_7358,N_5670);
nor U10384 (N_10384,N_9880,N_5656);
or U10385 (N_10385,N_8732,N_7469);
xnor U10386 (N_10386,N_5757,N_6271);
xnor U10387 (N_10387,N_9626,N_5030);
and U10388 (N_10388,N_8699,N_7360);
and U10389 (N_10389,N_8076,N_6456);
nand U10390 (N_10390,N_6086,N_6978);
and U10391 (N_10391,N_6805,N_6736);
and U10392 (N_10392,N_7542,N_5215);
and U10393 (N_10393,N_5244,N_5882);
or U10394 (N_10394,N_6489,N_9396);
or U10395 (N_10395,N_5716,N_5857);
nand U10396 (N_10396,N_9878,N_6507);
xor U10397 (N_10397,N_8906,N_9268);
nor U10398 (N_10398,N_7330,N_6593);
nor U10399 (N_10399,N_8611,N_8749);
and U10400 (N_10400,N_7563,N_6872);
xor U10401 (N_10401,N_8615,N_8632);
nor U10402 (N_10402,N_9843,N_8879);
nor U10403 (N_10403,N_9629,N_6319);
or U10404 (N_10404,N_9167,N_8849);
and U10405 (N_10405,N_7081,N_6433);
nor U10406 (N_10406,N_6902,N_5887);
or U10407 (N_10407,N_9459,N_7249);
or U10408 (N_10408,N_6044,N_7795);
nor U10409 (N_10409,N_5328,N_9781);
and U10410 (N_10410,N_7728,N_6882);
nand U10411 (N_10411,N_8459,N_5764);
nand U10412 (N_10412,N_6400,N_6040);
xnor U10413 (N_10413,N_5912,N_6427);
nor U10414 (N_10414,N_8678,N_7036);
or U10415 (N_10415,N_5609,N_6204);
nor U10416 (N_10416,N_8850,N_6757);
nand U10417 (N_10417,N_6160,N_9925);
nand U10418 (N_10418,N_6466,N_9550);
nand U10419 (N_10419,N_6442,N_9445);
or U10420 (N_10420,N_7271,N_5114);
and U10421 (N_10421,N_5101,N_5125);
nand U10422 (N_10422,N_5546,N_5179);
nor U10423 (N_10423,N_6804,N_5632);
xnor U10424 (N_10424,N_9208,N_5011);
nor U10425 (N_10425,N_8609,N_6856);
or U10426 (N_10426,N_8810,N_7618);
and U10427 (N_10427,N_7955,N_9180);
nor U10428 (N_10428,N_6761,N_5021);
nand U10429 (N_10429,N_9912,N_7084);
nand U10430 (N_10430,N_8584,N_5533);
xnor U10431 (N_10431,N_8261,N_6080);
or U10432 (N_10432,N_5572,N_8764);
or U10433 (N_10433,N_6886,N_8753);
and U10434 (N_10434,N_6203,N_9682);
xor U10435 (N_10435,N_7892,N_9685);
xnor U10436 (N_10436,N_9920,N_9853);
xor U10437 (N_10437,N_9693,N_9969);
xor U10438 (N_10438,N_8946,N_6800);
nor U10439 (N_10439,N_5078,N_7765);
or U10440 (N_10440,N_8736,N_8406);
and U10441 (N_10441,N_9971,N_5278);
xnor U10442 (N_10442,N_7284,N_8557);
xor U10443 (N_10443,N_7039,N_6048);
and U10444 (N_10444,N_7745,N_6646);
xnor U10445 (N_10445,N_9056,N_6855);
and U10446 (N_10446,N_7698,N_6730);
nor U10447 (N_10447,N_9282,N_5800);
xor U10448 (N_10448,N_9376,N_9038);
nor U10449 (N_10449,N_8622,N_7656);
and U10450 (N_10450,N_5667,N_6331);
nor U10451 (N_10451,N_6472,N_5806);
nand U10452 (N_10452,N_8827,N_8795);
or U10453 (N_10453,N_6421,N_6941);
xor U10454 (N_10454,N_7974,N_7815);
nor U10455 (N_10455,N_7224,N_6369);
nand U10456 (N_10456,N_6192,N_7769);
nor U10457 (N_10457,N_5304,N_5587);
nor U10458 (N_10458,N_6744,N_5155);
nor U10459 (N_10459,N_7357,N_5342);
or U10460 (N_10460,N_7723,N_5769);
xor U10461 (N_10461,N_7407,N_7334);
nand U10462 (N_10462,N_6877,N_9062);
nor U10463 (N_10463,N_6126,N_6598);
xor U10464 (N_10464,N_5385,N_9061);
or U10465 (N_10465,N_6465,N_5907);
and U10466 (N_10466,N_6110,N_5499);
xor U10467 (N_10467,N_9358,N_7816);
nand U10468 (N_10468,N_7417,N_8102);
nand U10469 (N_10469,N_8123,N_8518);
xor U10470 (N_10470,N_8330,N_9300);
and U10471 (N_10471,N_7218,N_9329);
nor U10472 (N_10472,N_5422,N_9892);
nand U10473 (N_10473,N_6674,N_7532);
nor U10474 (N_10474,N_5629,N_5802);
or U10475 (N_10475,N_7307,N_8000);
and U10476 (N_10476,N_6335,N_6128);
nor U10477 (N_10477,N_6753,N_8975);
nor U10478 (N_10478,N_6971,N_7423);
and U10479 (N_10479,N_8355,N_8154);
nand U10480 (N_10480,N_7860,N_5864);
nor U10481 (N_10481,N_6186,N_8466);
and U10482 (N_10482,N_5377,N_5354);
nor U10483 (N_10483,N_5016,N_9500);
nand U10484 (N_10484,N_8182,N_9999);
nand U10485 (N_10485,N_6824,N_7558);
and U10486 (N_10486,N_7965,N_7870);
xnor U10487 (N_10487,N_8473,N_5428);
xor U10488 (N_10488,N_8866,N_9953);
nor U10489 (N_10489,N_7950,N_7263);
and U10490 (N_10490,N_8465,N_6063);
or U10491 (N_10491,N_5024,N_5811);
or U10492 (N_10492,N_7944,N_8921);
nand U10493 (N_10493,N_8210,N_9681);
or U10494 (N_10494,N_8117,N_9852);
or U10495 (N_10495,N_6579,N_9129);
and U10496 (N_10496,N_8292,N_6197);
or U10497 (N_10497,N_7660,N_6950);
and U10498 (N_10498,N_7310,N_8242);
nand U10499 (N_10499,N_9375,N_8801);
nor U10500 (N_10500,N_9016,N_5088);
nor U10501 (N_10501,N_8703,N_9873);
nand U10502 (N_10502,N_8282,N_8926);
and U10503 (N_10503,N_5909,N_7272);
xnor U10504 (N_10504,N_9585,N_8914);
xor U10505 (N_10505,N_8952,N_9221);
and U10506 (N_10506,N_5093,N_5366);
or U10507 (N_10507,N_7017,N_8514);
and U10508 (N_10508,N_9562,N_9254);
nor U10509 (N_10509,N_7038,N_5979);
xor U10510 (N_10510,N_8141,N_7123);
xor U10511 (N_10511,N_9712,N_7623);
and U10512 (N_10512,N_7018,N_5270);
nor U10513 (N_10513,N_8166,N_7739);
and U10514 (N_10514,N_5263,N_7719);
nand U10515 (N_10515,N_8948,N_7831);
and U10516 (N_10516,N_6604,N_8240);
nand U10517 (N_10517,N_7144,N_8994);
xor U10518 (N_10518,N_6694,N_8812);
or U10519 (N_10519,N_9232,N_5009);
and U10520 (N_10520,N_8362,N_6697);
xnor U10521 (N_10521,N_5400,N_6103);
xnor U10522 (N_10522,N_9950,N_5678);
nand U10523 (N_10523,N_9371,N_9040);
and U10524 (N_10524,N_9918,N_7291);
nor U10525 (N_10525,N_5459,N_9768);
or U10526 (N_10526,N_7472,N_7538);
nor U10527 (N_10527,N_5528,N_6506);
xnor U10528 (N_10528,N_8644,N_6234);
nand U10529 (N_10529,N_7226,N_5898);
nand U10530 (N_10530,N_6146,N_8472);
xor U10531 (N_10531,N_9343,N_6360);
nand U10532 (N_10532,N_9087,N_8585);
and U10533 (N_10533,N_6017,N_6008);
nand U10534 (N_10534,N_5495,N_7575);
or U10535 (N_10535,N_6821,N_9255);
or U10536 (N_10536,N_9152,N_8597);
and U10537 (N_10537,N_8588,N_6179);
nor U10538 (N_10538,N_8693,N_5094);
or U10539 (N_10539,N_8392,N_8002);
or U10540 (N_10540,N_8577,N_7444);
xnor U10541 (N_10541,N_7657,N_5463);
xnor U10542 (N_10542,N_7266,N_6556);
and U10543 (N_10543,N_7943,N_6286);
or U10544 (N_10544,N_5464,N_7904);
and U10545 (N_10545,N_5398,N_5001);
nor U10546 (N_10546,N_7644,N_5308);
nor U10547 (N_10547,N_9168,N_7705);
xnor U10548 (N_10548,N_6813,N_8979);
xnor U10549 (N_10549,N_6636,N_8824);
nor U10550 (N_10550,N_8794,N_9642);
and U10551 (N_10551,N_7830,N_8358);
and U10552 (N_10552,N_7471,N_9706);
nor U10553 (N_10553,N_6564,N_8253);
nand U10554 (N_10554,N_6717,N_6218);
or U10555 (N_10555,N_9800,N_9540);
or U10556 (N_10556,N_5368,N_7513);
nor U10557 (N_10557,N_9803,N_7744);
nor U10558 (N_10558,N_8228,N_5485);
or U10559 (N_10559,N_5172,N_6583);
or U10560 (N_10560,N_8513,N_7473);
nand U10561 (N_10561,N_8515,N_6907);
nand U10562 (N_10562,N_6441,N_7346);
nand U10563 (N_10563,N_8549,N_7540);
nand U10564 (N_10564,N_5998,N_9591);
nor U10565 (N_10565,N_6274,N_5042);
and U10566 (N_10566,N_7329,N_8617);
nand U10567 (N_10567,N_7119,N_5474);
nand U10568 (N_10568,N_9116,N_7254);
or U10569 (N_10569,N_9879,N_9294);
nand U10570 (N_10570,N_9130,N_5208);
and U10571 (N_10571,N_5607,N_9869);
xnor U10572 (N_10572,N_7362,N_9197);
or U10573 (N_10573,N_9432,N_7779);
nor U10574 (N_10574,N_7877,N_7268);
nand U10575 (N_10575,N_7354,N_9387);
nand U10576 (N_10576,N_6443,N_6518);
xor U10577 (N_10577,N_8846,N_7680);
and U10578 (N_10578,N_8435,N_6906);
or U10579 (N_10579,N_9074,N_8037);
nand U10580 (N_10580,N_9400,N_5827);
nand U10581 (N_10581,N_6509,N_5372);
or U10582 (N_10582,N_8367,N_6602);
or U10583 (N_10583,N_8385,N_5455);
nor U10584 (N_10584,N_6536,N_8516);
nand U10585 (N_10585,N_5438,N_6131);
xor U10586 (N_10586,N_5833,N_5253);
nand U10587 (N_10587,N_7187,N_6946);
xnor U10588 (N_10588,N_6523,N_9911);
nand U10589 (N_10589,N_5154,N_7311);
and U10590 (N_10590,N_8439,N_6738);
and U10591 (N_10591,N_8839,N_6826);
or U10592 (N_10592,N_7255,N_6033);
nand U10593 (N_10593,N_8562,N_5838);
xor U10594 (N_10594,N_6247,N_5863);
and U10595 (N_10595,N_8545,N_6686);
nand U10596 (N_10596,N_5375,N_9865);
xor U10597 (N_10597,N_7495,N_8723);
nand U10598 (N_10598,N_9159,N_8637);
xnor U10599 (N_10599,N_5999,N_5496);
and U10600 (N_10600,N_7747,N_9089);
nor U10601 (N_10601,N_6845,N_5519);
and U10602 (N_10602,N_5614,N_7854);
xor U10603 (N_10603,N_7886,N_8499);
and U10604 (N_10604,N_6047,N_8556);
nand U10605 (N_10605,N_7013,N_5106);
xor U10606 (N_10606,N_7350,N_6794);
xor U10607 (N_10607,N_9699,N_9572);
or U10608 (N_10608,N_7593,N_7118);
and U10609 (N_10609,N_8165,N_5625);
or U10610 (N_10610,N_7786,N_5363);
or U10611 (N_10611,N_7808,N_9743);
nor U10612 (N_10612,N_9840,N_6942);
or U10613 (N_10613,N_8317,N_7126);
xnor U10614 (N_10614,N_6416,N_6444);
xor U10615 (N_10615,N_6268,N_7006);
xor U10616 (N_10616,N_6220,N_6083);
nand U10617 (N_10617,N_9820,N_8595);
and U10618 (N_10618,N_6681,N_9034);
xnor U10619 (N_10619,N_6550,N_7184);
and U10620 (N_10620,N_8291,N_5809);
xor U10621 (N_10621,N_8944,N_7315);
nor U10622 (N_10622,N_7398,N_6531);
and U10623 (N_10623,N_5064,N_9308);
xor U10624 (N_10624,N_8341,N_5826);
nand U10625 (N_10625,N_6120,N_9423);
nor U10626 (N_10626,N_7429,N_7988);
nor U10627 (N_10627,N_7676,N_8029);
or U10628 (N_10628,N_7341,N_7555);
xnor U10629 (N_10629,N_6988,N_7169);
nor U10630 (N_10630,N_5110,N_5079);
nand U10631 (N_10631,N_6482,N_5862);
nor U10632 (N_10632,N_8654,N_6121);
nor U10633 (N_10633,N_5489,N_6980);
or U10634 (N_10634,N_6376,N_5086);
or U10635 (N_10635,N_6172,N_5759);
xnor U10636 (N_10636,N_5832,N_5942);
xnor U10637 (N_10637,N_8455,N_8574);
xnor U10638 (N_10638,N_5822,N_6881);
nand U10639 (N_10639,N_5219,N_9850);
nor U10640 (N_10640,N_5630,N_5530);
or U10641 (N_10641,N_7422,N_5410);
xor U10642 (N_10642,N_7889,N_9379);
and U10643 (N_10643,N_8318,N_7406);
or U10644 (N_10644,N_8336,N_9273);
nand U10645 (N_10645,N_5234,N_7605);
xor U10646 (N_10646,N_9443,N_8024);
xnor U10647 (N_10647,N_8283,N_8540);
nor U10648 (N_10648,N_7933,N_8828);
and U10649 (N_10649,N_6240,N_5874);
nand U10650 (N_10650,N_8500,N_6201);
and U10651 (N_10651,N_8635,N_9465);
nor U10652 (N_10652,N_8489,N_8848);
nand U10653 (N_10653,N_5621,N_6774);
or U10654 (N_10654,N_8982,N_5526);
xor U10655 (N_10655,N_7506,N_8885);
and U10656 (N_10656,N_6127,N_6605);
and U10657 (N_10657,N_6910,N_6260);
nand U10658 (N_10658,N_5747,N_7774);
nor U10659 (N_10659,N_7864,N_9325);
nor U10660 (N_10660,N_7699,N_9242);
and U10661 (N_10661,N_5613,N_5146);
nor U10662 (N_10662,N_8451,N_7024);
nand U10663 (N_10663,N_5876,N_6102);
and U10664 (N_10664,N_8201,N_6370);
nand U10665 (N_10665,N_7646,N_8759);
nor U10666 (N_10666,N_5745,N_5739);
and U10667 (N_10667,N_8949,N_9370);
xor U10668 (N_10668,N_5250,N_8101);
nor U10669 (N_10669,N_9393,N_8419);
and U10670 (N_10670,N_6695,N_5886);
nor U10671 (N_10671,N_8531,N_9857);
or U10672 (N_10672,N_7823,N_6423);
and U10673 (N_10673,N_6823,N_7106);
and U10674 (N_10674,N_5117,N_8718);
xor U10675 (N_10675,N_7295,N_5896);
xor U10676 (N_10676,N_9296,N_9676);
xor U10677 (N_10677,N_5969,N_8209);
or U10678 (N_10678,N_5493,N_5212);
or U10679 (N_10679,N_5118,N_9057);
nor U10680 (N_10680,N_6009,N_6732);
nor U10681 (N_10681,N_8314,N_8872);
nand U10682 (N_10682,N_6289,N_7803);
nor U10683 (N_10683,N_7920,N_8842);
and U10684 (N_10684,N_5725,N_9828);
and U10685 (N_10685,N_7837,N_9944);
nor U10686 (N_10686,N_9224,N_9200);
nor U10687 (N_10687,N_6947,N_8087);
and U10688 (N_10688,N_5523,N_9792);
xor U10689 (N_10689,N_5279,N_5527);
xnor U10690 (N_10690,N_7308,N_5646);
nor U10691 (N_10691,N_8670,N_9252);
or U10692 (N_10692,N_8573,N_5033);
xor U10693 (N_10693,N_9775,N_5152);
or U10694 (N_10694,N_5503,N_6972);
nor U10695 (N_10695,N_9039,N_9270);
nor U10696 (N_10696,N_5242,N_5188);
xnor U10697 (N_10697,N_7645,N_8275);
or U10698 (N_10698,N_8023,N_8360);
or U10699 (N_10699,N_9471,N_5765);
nand U10700 (N_10700,N_6700,N_9450);
nor U10701 (N_10701,N_7637,N_7120);
and U10702 (N_10702,N_5577,N_9244);
xnor U10703 (N_10703,N_8893,N_9678);
and U10704 (N_10704,N_8643,N_6594);
nor U10705 (N_10705,N_7022,N_8506);
nand U10706 (N_10706,N_9749,N_9068);
nor U10707 (N_10707,N_5048,N_5470);
xnor U10708 (N_10708,N_6914,N_8599);
or U10709 (N_10709,N_9433,N_6637);
or U10710 (N_10710,N_7544,N_7629);
xor U10711 (N_10711,N_7215,N_9386);
nor U10712 (N_10712,N_6837,N_6621);
or U10713 (N_10713,N_6822,N_8696);
xnor U10714 (N_10714,N_7079,N_7994);
and U10715 (N_10715,N_5352,N_6865);
xnor U10716 (N_10716,N_5479,N_8607);
or U10717 (N_10717,N_8168,N_7806);
nor U10718 (N_10718,N_8667,N_5957);
xnor U10719 (N_10719,N_5962,N_8442);
nand U10720 (N_10720,N_8339,N_8104);
and U10721 (N_10721,N_6534,N_8313);
or U10722 (N_10722,N_5600,N_7227);
and U10723 (N_10723,N_5881,N_7259);
or U10724 (N_10724,N_8507,N_6256);
nor U10725 (N_10725,N_5243,N_5758);
xnor U10726 (N_10726,N_5481,N_8477);
xnor U10727 (N_10727,N_6292,N_6043);
xor U10728 (N_10728,N_8886,N_9045);
xnor U10729 (N_10729,N_9795,N_5792);
xor U10730 (N_10730,N_6038,N_7446);
xnor U10731 (N_10731,N_9664,N_6069);
and U10732 (N_10732,N_9028,N_9513);
nand U10733 (N_10733,N_7230,N_9290);
xnor U10734 (N_10734,N_7083,N_7730);
and U10735 (N_10735,N_8187,N_6763);
xor U10736 (N_10736,N_5766,N_8823);
and U10737 (N_10737,N_6969,N_8796);
xnor U10738 (N_10738,N_6818,N_7807);
xnor U10739 (N_10739,N_8642,N_9398);
xor U10740 (N_10740,N_7541,N_9518);
or U10741 (N_10741,N_6493,N_9514);
xor U10742 (N_10742,N_8052,N_5447);
and U10743 (N_10743,N_7684,N_8284);
nand U10744 (N_10744,N_9978,N_8613);
nor U10745 (N_10745,N_6199,N_6521);
nand U10746 (N_10746,N_8747,N_9140);
xnor U10747 (N_10747,N_6284,N_5167);
nor U10748 (N_10748,N_8698,N_6075);
xor U10749 (N_10749,N_9721,N_5925);
xnor U10750 (N_10750,N_6314,N_6365);
nor U10751 (N_10751,N_5504,N_6723);
xor U10752 (N_10752,N_9638,N_8320);
xnor U10753 (N_10753,N_7797,N_9903);
nor U10754 (N_10754,N_5984,N_9377);
and U10755 (N_10755,N_7977,N_7258);
nor U10756 (N_10756,N_7436,N_5955);
or U10757 (N_10757,N_6501,N_6795);
or U10758 (N_10758,N_5484,N_7557);
nand U10759 (N_10759,N_9223,N_8328);
nor U10760 (N_10760,N_5706,N_9189);
xor U10761 (N_10761,N_6422,N_6535);
nor U10762 (N_10762,N_7634,N_6394);
or U10763 (N_10763,N_9072,N_5073);
or U10764 (N_10764,N_9788,N_7403);
or U10765 (N_10765,N_5264,N_7277);
and U10766 (N_10766,N_7326,N_6058);
nor U10767 (N_10767,N_9688,N_5928);
or U10768 (N_10768,N_7679,N_5246);
xnor U10769 (N_10769,N_8226,N_7246);
and U10770 (N_10770,N_8357,N_6015);
or U10771 (N_10771,N_5752,N_8996);
nand U10772 (N_10772,N_9972,N_8563);
and U10773 (N_10773,N_9117,N_6176);
xor U10774 (N_10774,N_6714,N_8591);
nand U10775 (N_10775,N_7843,N_5319);
and U10776 (N_10776,N_8268,N_8691);
and U10777 (N_10777,N_9526,N_8927);
xor U10778 (N_10778,N_7007,N_9653);
xnor U10779 (N_10779,N_5697,N_7918);
nor U10780 (N_10780,N_9659,N_6623);
nand U10781 (N_10781,N_8934,N_6696);
xor U10782 (N_10782,N_9464,N_6711);
nand U10783 (N_10783,N_8943,N_6470);
and U10784 (N_10784,N_7998,N_5043);
and U10785 (N_10785,N_5612,N_8495);
nor U10786 (N_10786,N_7297,N_5537);
nor U10787 (N_10787,N_7946,N_8631);
xnor U10788 (N_10788,N_9689,N_5191);
nor U10789 (N_10789,N_5872,N_8370);
or U10790 (N_10790,N_6678,N_5072);
xor U10791 (N_10791,N_8247,N_7802);
xnor U10792 (N_10792,N_8945,N_7917);
nand U10793 (N_10793,N_9160,N_9002);
nand U10794 (N_10794,N_6469,N_5604);
and U10795 (N_10795,N_6526,N_9454);
or U10796 (N_10796,N_6538,N_7934);
and U10797 (N_10797,N_6277,N_7100);
nor U10798 (N_10798,N_6053,N_7651);
xor U10799 (N_10799,N_6776,N_9776);
xnor U10800 (N_10800,N_5793,N_9385);
and U10801 (N_10801,N_9818,N_6677);
or U10802 (N_10802,N_5090,N_9571);
xnor U10803 (N_10803,N_8014,N_9233);
and U10804 (N_10804,N_6072,N_7245);
xor U10805 (N_10805,N_8265,N_9331);
nand U10806 (N_10806,N_7612,N_5933);
or U10807 (N_10807,N_7072,N_7643);
nand U10808 (N_10808,N_9147,N_9101);
or U10809 (N_10809,N_7539,N_6280);
nor U10810 (N_10810,N_6829,N_6524);
and U10811 (N_10811,N_6647,N_9359);
or U10812 (N_10812,N_9939,N_9817);
nor U10813 (N_10813,N_5662,N_5080);
xnor U10814 (N_10814,N_9145,N_9099);
and U10815 (N_10815,N_8246,N_8505);
or U10816 (N_10816,N_9047,N_6853);
and U10817 (N_10817,N_5703,N_5112);
and U10818 (N_10818,N_5205,N_5650);
or U10819 (N_10819,N_9320,N_5638);
and U10820 (N_10820,N_6897,N_5283);
xor U10821 (N_10821,N_8003,N_8533);
nor U10822 (N_10822,N_6224,N_6122);
nor U10823 (N_10823,N_9010,N_9637);
nand U10824 (N_10824,N_5859,N_7839);
nor U10825 (N_10825,N_7280,N_9958);
nand U10826 (N_10826,N_9104,N_6683);
or U10827 (N_10827,N_6230,N_6693);
or U10828 (N_10828,N_8429,N_6177);
nor U10829 (N_10829,N_5445,N_9942);
nand U10830 (N_10830,N_7726,N_5531);
nand U10831 (N_10831,N_8403,N_6899);
nand U10832 (N_10832,N_6097,N_6373);
nand U10833 (N_10833,N_9286,N_9521);
and U10834 (N_10834,N_7099,N_7095);
nand U10835 (N_10835,N_9801,N_8808);
nor U10836 (N_10836,N_7894,N_8867);
and U10837 (N_10837,N_5145,N_8766);
or U10838 (N_10838,N_9730,N_8884);
nor U10839 (N_10839,N_6668,N_7932);
and U10840 (N_10840,N_5651,N_7743);
nand U10841 (N_10841,N_5466,N_6002);
and U10842 (N_10842,N_5854,N_8663);
xnor U10843 (N_10843,N_5039,N_9893);
and U10844 (N_10844,N_6525,N_9003);
or U10845 (N_10845,N_8636,N_9310);
or U10846 (N_10846,N_6006,N_6987);
or U10847 (N_10847,N_7603,N_9051);
or U10848 (N_10848,N_7484,N_6601);
and U10849 (N_10849,N_7574,N_7746);
xor U10850 (N_10850,N_9683,N_9901);
or U10851 (N_10851,N_9621,N_5306);
xor U10852 (N_10852,N_8928,N_5991);
nor U10853 (N_10853,N_9923,N_6733);
xnor U10854 (N_10854,N_9452,N_8493);
xor U10855 (N_10855,N_6323,N_6748);
or U10856 (N_10856,N_6411,N_6862);
and U10857 (N_10857,N_7479,N_9247);
nor U10858 (N_10858,N_8679,N_9401);
nor U10859 (N_10859,N_6654,N_7936);
nor U10860 (N_10860,N_5296,N_8390);
nor U10861 (N_10861,N_9679,N_5616);
nor U10862 (N_10862,N_7111,N_8041);
and U10863 (N_10863,N_7468,N_6554);
nor U10864 (N_10864,N_5545,N_5807);
nand U10865 (N_10865,N_8737,N_5648);
and U10866 (N_10866,N_8266,N_7794);
nand U10867 (N_10867,N_5130,N_9622);
or U10868 (N_10868,N_9416,N_7678);
and U10869 (N_10869,N_5681,N_5008);
and U10870 (N_10870,N_6773,N_9226);
xor U10871 (N_10871,N_6461,N_8687);
nand U10872 (N_10872,N_6092,N_5636);
or U10873 (N_10873,N_9510,N_6381);
nand U10874 (N_10874,N_5543,N_7849);
and U10875 (N_10875,N_9773,N_7046);
and U10876 (N_10876,N_7619,N_5338);
xor U10877 (N_10877,N_9832,N_9380);
and U10878 (N_10878,N_7440,N_6316);
xnor U10879 (N_10879,N_5178,N_9304);
xor U10880 (N_10880,N_6724,N_8671);
xor U10881 (N_10881,N_5429,N_5761);
nand U10882 (N_10882,N_9697,N_7566);
and U10883 (N_10883,N_5702,N_6171);
or U10884 (N_10884,N_5029,N_8153);
or U10885 (N_10885,N_8702,N_5514);
nor U10886 (N_10886,N_7186,N_6861);
xor U10887 (N_10887,N_7948,N_8033);
xnor U10888 (N_10888,N_5737,N_6566);
or U10889 (N_10889,N_7916,N_9532);
nor U10890 (N_10890,N_6999,N_8474);
xor U10891 (N_10891,N_9847,N_8862);
and U10892 (N_10892,N_9715,N_9066);
xor U10893 (N_10893,N_6740,N_5788);
nor U10894 (N_10894,N_8484,N_5348);
nand U10895 (N_10895,N_5332,N_8443);
and U10896 (N_10896,N_6315,N_6913);
xnor U10897 (N_10897,N_9081,N_8826);
nand U10898 (N_10898,N_6333,N_8405);
nand U10899 (N_10899,N_5245,N_5480);
nand U10900 (N_10900,N_9734,N_5258);
and U10901 (N_10901,N_6468,N_5097);
nor U10902 (N_10902,N_5968,N_6345);
xnor U10903 (N_10903,N_9334,N_7045);
nor U10904 (N_10904,N_8501,N_5615);
and U10905 (N_10905,N_9512,N_9759);
and U10906 (N_10906,N_8993,N_8529);
xor U10907 (N_10907,N_7336,N_7182);
nor U10908 (N_10908,N_7170,N_5214);
nand U10909 (N_10909,N_6760,N_7510);
nor U10910 (N_10910,N_8576,N_9143);
xor U10911 (N_10911,N_5482,N_7770);
and U10912 (N_10912,N_7511,N_8510);
nor U10913 (N_10913,N_7279,N_9141);
nand U10914 (N_10914,N_5552,N_7710);
or U10915 (N_10915,N_5548,N_7004);
nand U10916 (N_10916,N_9174,N_7500);
xnor U10917 (N_10917,N_9644,N_7108);
and U10918 (N_10918,N_9352,N_9365);
xor U10919 (N_10919,N_7391,N_8196);
or U10920 (N_10920,N_8787,N_5149);
nor U10921 (N_10921,N_5883,N_8178);
nor U10922 (N_10922,N_6173,N_9531);
and U10923 (N_10923,N_8570,N_9763);
nand U10924 (N_10924,N_9656,N_8259);
or U10925 (N_10925,N_8963,N_8129);
or U10926 (N_10926,N_5333,N_5330);
nand U10927 (N_10927,N_5755,N_9819);
xnor U10928 (N_10928,N_5844,N_8380);
nand U10929 (N_10929,N_7281,N_9489);
xor U10930 (N_10930,N_8143,N_6311);
xor U10931 (N_10931,N_5444,N_8192);
nor U10932 (N_10932,N_5931,N_8793);
and U10933 (N_10933,N_7993,N_5558);
or U10934 (N_10934,N_7136,N_6690);
xnor U10935 (N_10935,N_5922,N_7577);
xnor U10936 (N_10936,N_8423,N_7919);
nand U10937 (N_10937,N_8647,N_6615);
nand U10938 (N_10938,N_5562,N_6491);
nor U10939 (N_10939,N_8363,N_9767);
xor U10940 (N_10940,N_9778,N_8194);
or U10941 (N_10941,N_7068,N_7610);
and U10942 (N_10942,N_5935,N_5233);
and U10943 (N_10943,N_6251,N_8359);
xnor U10944 (N_10944,N_8375,N_8618);
nand U10945 (N_10945,N_9602,N_7122);
xor U10946 (N_10946,N_6061,N_6239);
nor U10947 (N_10947,N_6864,N_9613);
nor U10948 (N_10948,N_5506,N_6065);
and U10949 (N_10949,N_8772,N_7367);
or U10950 (N_10950,N_7547,N_6004);
or U10951 (N_10951,N_7771,N_7565);
nor U10952 (N_10952,N_8950,N_8822);
nand U10953 (N_10953,N_8263,N_6341);
and U10954 (N_10954,N_8480,N_6355);
xnor U10955 (N_10955,N_9382,N_7264);
nand U10956 (N_10956,N_9361,N_7995);
and U10957 (N_10957,N_5958,N_6852);
nand U10958 (N_10958,N_7296,N_8610);
and U10959 (N_10959,N_9934,N_6573);
nand U10960 (N_10960,N_7788,N_6380);
or U10961 (N_10961,N_8983,N_5966);
nand U10962 (N_10962,N_6109,N_5307);
nor U10963 (N_10963,N_6113,N_6124);
or U10964 (N_10964,N_7596,N_5272);
xor U10965 (N_10965,N_9708,N_7411);
nor U10966 (N_10966,N_9144,N_9872);
or U10967 (N_10967,N_7842,N_6094);
or U10968 (N_10968,N_7838,N_8881);
xor U10969 (N_10969,N_5664,N_7058);
xnor U10970 (N_10970,N_5190,N_5858);
nor U10971 (N_10971,N_9724,N_7826);
xnor U10972 (N_10972,N_6918,N_8190);
nor U10973 (N_10973,N_6948,N_6458);
or U10974 (N_10974,N_6490,N_7560);
and U10975 (N_10975,N_8356,N_8871);
nor U10976 (N_10976,N_5126,N_7175);
nand U10977 (N_10977,N_8193,N_8157);
nand U10978 (N_10978,N_8323,N_6282);
xnor U10979 (N_10979,N_5137,N_8279);
nand U10980 (N_10980,N_6764,N_9315);
nand U10981 (N_10981,N_5990,N_8987);
xor U10982 (N_10982,N_6281,N_6982);
xor U10983 (N_10983,N_8321,N_7352);
nand U10984 (N_10984,N_9455,N_5223);
and U10985 (N_10985,N_7737,N_7229);
nor U10986 (N_10986,N_6213,N_9411);
and U10987 (N_10987,N_5164,N_7010);
xor U10988 (N_10988,N_5468,N_6036);
xnor U10989 (N_10989,N_8203,N_9582);
and U10990 (N_10990,N_5652,N_6561);
nor U10991 (N_10991,N_8144,N_6159);
xor U10992 (N_10992,N_7413,N_8757);
or U10993 (N_10993,N_7694,N_6651);
nor U10994 (N_10994,N_8870,N_5729);
xor U10995 (N_10995,N_8214,N_9771);
xor U10996 (N_10996,N_9065,N_6474);
or U10997 (N_10997,N_7978,N_6919);
xnor U10998 (N_10998,N_5395,N_7432);
nor U10999 (N_10999,N_7594,N_6059);
nor U11000 (N_11000,N_8704,N_9480);
or U11001 (N_11001,N_7335,N_7759);
nand U11002 (N_11002,N_8324,N_6505);
xor U11003 (N_11003,N_6261,N_7982);
nor U11004 (N_11004,N_8239,N_7591);
and U11005 (N_11005,N_7427,N_8289);
nand U11006 (N_11006,N_8044,N_5199);
nand U11007 (N_11007,N_8391,N_9291);
nand U11008 (N_11008,N_9109,N_6814);
nor U11009 (N_11009,N_7731,N_5696);
or U11010 (N_11010,N_8551,N_6403);
and U11011 (N_11011,N_7361,N_9338);
or U11012 (N_11012,N_9444,N_5741);
nor U11013 (N_11013,N_8951,N_7628);
nor U11014 (N_11014,N_7438,N_9897);
nor U11015 (N_11015,N_5535,N_8028);
nor U11016 (N_11016,N_7453,N_7210);
nand U11017 (N_11017,N_6847,N_9533);
nand U11018 (N_11018,N_8280,N_9342);
or U11019 (N_11019,N_8589,N_9150);
xnor U11020 (N_11020,N_6639,N_7041);
and U11021 (N_11021,N_7466,N_9671);
nand U11022 (N_11022,N_8783,N_6620);
or U11023 (N_11023,N_9502,N_5129);
nor U11024 (N_11024,N_9311,N_8216);
or U11025 (N_11025,N_6854,N_7583);
or U11026 (N_11026,N_7778,N_6701);
or U11027 (N_11027,N_8728,N_5731);
and U11028 (N_11028,N_5201,N_8930);
and U11029 (N_11029,N_7509,N_7689);
and U11030 (N_11030,N_6457,N_9545);
nand U11031 (N_11031,N_8621,N_7049);
and U11032 (N_11032,N_8743,N_6994);
xnor U11033 (N_11033,N_7177,N_5423);
xor U11034 (N_11034,N_5364,N_9835);
nor U11035 (N_11035,N_8820,N_5815);
nand U11036 (N_11036,N_8401,N_6229);
xnor U11037 (N_11037,N_5071,N_7533);
xor U11038 (N_11038,N_9246,N_7303);
and U11039 (N_11039,N_6545,N_9605);
nor U11040 (N_11040,N_8620,N_5839);
and U11041 (N_11041,N_5229,N_6767);
nor U11042 (N_11042,N_8381,N_6288);
xnor U11043 (N_11043,N_5259,N_7590);
nor U11044 (N_11044,N_5019,N_8208);
or U11045 (N_11045,N_8593,N_9625);
and U11046 (N_11046,N_9473,N_6049);
nand U11047 (N_11047,N_8043,N_7383);
nor U11048 (N_11048,N_6859,N_5623);
or U11049 (N_11049,N_6392,N_8249);
and U11050 (N_11050,N_5911,N_8411);
nor U11051 (N_11051,N_5798,N_6816);
xnor U11052 (N_11052,N_5040,N_7370);
or U11053 (N_11053,N_5074,N_9790);
nand U11054 (N_11054,N_9249,N_9440);
and U11055 (N_11055,N_7109,N_7630);
nand U11056 (N_11056,N_8250,N_6166);
nor U11057 (N_11057,N_8682,N_9020);
nand U11058 (N_11058,N_9700,N_5345);
nor U11059 (N_11059,N_5109,N_8986);
or U11060 (N_11060,N_6413,N_8596);
or U11061 (N_11061,N_7581,N_5441);
nor U11062 (N_11062,N_8335,N_9492);
xor U11063 (N_11063,N_6975,N_7664);
xnor U11064 (N_11064,N_7216,N_8426);
xnor U11065 (N_11065,N_7183,N_7766);
nor U11066 (N_11066,N_9193,N_8955);
or U11067 (N_11067,N_9067,N_5268);
and U11068 (N_11068,N_7638,N_7958);
nor U11069 (N_11069,N_8382,N_6366);
nand U11070 (N_11070,N_9478,N_9568);
xor U11071 (N_11071,N_6860,N_6332);
or U11072 (N_11072,N_5036,N_7292);
nand U11073 (N_11073,N_7225,N_6569);
nor U11074 (N_11074,N_8776,N_8969);
and U11075 (N_11075,N_6189,N_9054);
and U11076 (N_11076,N_9799,N_9970);
nor U11077 (N_11077,N_6045,N_8175);
or U11078 (N_11078,N_9272,N_5005);
and U11079 (N_11079,N_7027,N_5378);
nor U11080 (N_11080,N_8184,N_9684);
xor U11081 (N_11081,N_6156,N_9940);
nand U11082 (N_11082,N_9906,N_5471);
nor U11083 (N_11083,N_8299,N_9855);
or U11084 (N_11084,N_6675,N_8898);
nand U11085 (N_11085,N_7302,N_7624);
xor U11086 (N_11086,N_5628,N_5744);
nand U11087 (N_11087,N_9142,N_9690);
or U11088 (N_11088,N_9399,N_9076);
nand U11089 (N_11089,N_8285,N_9589);
nand U11090 (N_11090,N_5710,N_6956);
nor U11091 (N_11091,N_8485,N_6618);
nor U11092 (N_11092,N_7792,N_8508);
and U11093 (N_11093,N_7717,N_9549);
nor U11094 (N_11094,N_5698,N_8340);
and U11095 (N_11095,N_5819,N_6338);
or U11096 (N_11096,N_5297,N_8937);
xnor U11097 (N_11097,N_5595,N_5669);
nor U11098 (N_11098,N_7654,N_8568);
nor U11099 (N_11099,N_7071,N_9213);
nand U11100 (N_11100,N_8088,N_7193);
nand U11101 (N_11101,N_9516,N_8206);
or U11102 (N_11102,N_7171,N_6178);
xnor U11103 (N_11103,N_8854,N_6137);
or U11104 (N_11104,N_5063,N_5932);
xor U11105 (N_11105,N_8084,N_6848);
and U11106 (N_11106,N_5453,N_6562);
and U11107 (N_11107,N_5787,N_8073);
nand U11108 (N_11108,N_8170,N_5273);
nand U11109 (N_11109,N_8876,N_7419);
nand U11110 (N_11110,N_5158,N_7910);
or U11111 (N_11111,N_5753,N_7881);
nor U11112 (N_11112,N_7996,N_7219);
nand U11113 (N_11113,N_8069,N_6459);
and U11114 (N_11114,N_6300,N_8133);
nor U11115 (N_11115,N_5914,N_6685);
and U11116 (N_11116,N_7414,N_6502);
xnor U11117 (N_11117,N_5878,N_6527);
nor U11118 (N_11118,N_5892,N_7784);
nor U11119 (N_11119,N_6850,N_9018);
and U11120 (N_11120,N_5418,N_9654);
nand U11121 (N_11121,N_6205,N_9169);
nor U11122 (N_11122,N_6768,N_5782);
nand U11123 (N_11123,N_7282,N_5353);
xor U11124 (N_11124,N_5442,N_6887);
or U11125 (N_11125,N_5866,N_8105);
xnor U11126 (N_11126,N_5014,N_8064);
or U11127 (N_11127,N_7492,N_6935);
nor U11128 (N_11128,N_8177,N_7260);
or U11129 (N_11129,N_6368,N_5736);
nand U11130 (N_11130,N_5150,N_7478);
nor U11131 (N_11131,N_5773,N_5974);
nand U11132 (N_11132,N_8080,N_7322);
nand U11133 (N_11133,N_5760,N_6920);
xnor U11134 (N_11134,N_5404,N_6609);
nand U11135 (N_11135,N_7911,N_9764);
and U11136 (N_11136,N_6529,N_8070);
xnor U11137 (N_11137,N_9639,N_9930);
or U11138 (N_11138,N_6077,N_8183);
and U11139 (N_11139,N_8223,N_7290);
xor U11140 (N_11140,N_8947,N_6090);
and U11141 (N_11141,N_9389,N_9523);
nor U11142 (N_11142,N_6777,N_5684);
xnor U11143 (N_11143,N_7668,N_5817);
nor U11144 (N_11144,N_8583,N_8007);
nor U11145 (N_11145,N_9420,N_8853);
and U11146 (N_11146,N_5637,N_6834);
or U11147 (N_11147,N_9783,N_8912);
nor U11148 (N_11148,N_9106,N_6959);
nand U11149 (N_11149,N_6302,N_8750);
or U11150 (N_11150,N_5852,N_7211);
nor U11151 (N_11151,N_8121,N_8816);
or U11152 (N_11152,N_6014,N_7695);
nor U11153 (N_11153,N_8569,N_9599);
xnor U11154 (N_11154,N_5977,N_6892);
and U11155 (N_11155,N_9866,N_7056);
or U11156 (N_11156,N_5640,N_7921);
nor U11157 (N_11157,N_9154,N_6223);
xor U11158 (N_11158,N_5477,N_8901);
nand U11159 (N_11159,N_7365,N_7608);
and U11160 (N_11160,N_9102,N_7648);
or U11161 (N_11161,N_6032,N_8019);
nand U11162 (N_11162,N_6515,N_8337);
xnor U11163 (N_11163,N_6974,N_6170);
or U11164 (N_11164,N_8278,N_9032);
nand U11165 (N_11165,N_8197,N_9529);
nand U11166 (N_11166,N_5812,N_5406);
nor U11167 (N_11167,N_5458,N_8600);
nor U11168 (N_11168,N_5360,N_7879);
xnor U11169 (N_11169,N_7001,N_5983);
nor U11170 (N_11170,N_5903,N_5055);
and U11171 (N_11171,N_8425,N_6436);
xnor U11172 (N_11172,N_5256,N_7729);
xor U11173 (N_11173,N_8860,N_5066);
nor U11174 (N_11174,N_6612,N_9293);
or U11175 (N_11175,N_9535,N_5797);
or U11176 (N_11176,N_5303,N_7107);
xnor U11177 (N_11177,N_5313,N_8119);
xor U11178 (N_11178,N_9527,N_5239);
xnor U11179 (N_11179,N_5665,N_8956);
and U11180 (N_11180,N_6114,N_7891);
nand U11181 (N_11181,N_6046,N_5947);
and U11182 (N_11182,N_8049,N_6624);
and U11183 (N_11183,N_9956,N_9112);
xor U11184 (N_11184,N_9520,N_5704);
and U11185 (N_11185,N_9479,N_8967);
or U11186 (N_11186,N_8660,N_7476);
nand U11187 (N_11187,N_5712,N_9974);
xor U11188 (N_11188,N_9397,N_7143);
xnor U11189 (N_11189,N_8396,N_8777);
or U11190 (N_11190,N_6900,N_9646);
and U11191 (N_11191,N_6001,N_8754);
nand U11192 (N_11192,N_6151,N_7516);
and U11193 (N_11193,N_9804,N_6831);
nor U11194 (N_11194,N_9467,N_9424);
xor U11195 (N_11195,N_7080,N_5454);
or U11196 (N_11196,N_8954,N_8821);
and U11197 (N_11197,N_6350,N_6512);
xor U11198 (N_11198,N_5643,N_7040);
and U11199 (N_11199,N_9053,N_8925);
xor U11200 (N_11200,N_9522,N_9686);
xor U11201 (N_11201,N_8145,N_6547);
nor U11202 (N_11202,N_5525,N_7528);
nand U11203 (N_11203,N_9161,N_5981);
and U11204 (N_11204,N_8140,N_5095);
nand U11205 (N_11205,N_7588,N_9468);
or U11206 (N_11206,N_8188,N_7293);
and U11207 (N_11207,N_9220,N_9711);
or U11208 (N_11208,N_8481,N_5198);
nand U11209 (N_11209,N_9439,N_9780);
nor U11210 (N_11210,N_5369,N_5567);
nand U11211 (N_11211,N_5890,N_6480);
nand U11212 (N_11212,N_7283,N_7754);
and U11213 (N_11213,N_9558,N_8388);
or U11214 (N_11214,N_5762,N_9777);
or U11215 (N_11215,N_6093,N_7066);
nor U11216 (N_11216,N_8778,N_9560);
xor U11217 (N_11217,N_7238,N_9108);
or U11218 (N_11218,N_7866,N_8984);
xor U11219 (N_11219,N_7221,N_7852);
nor U11220 (N_11220,N_5456,N_5799);
nand U11221 (N_11221,N_6375,N_6471);
xor U11222 (N_11222,N_8673,N_8792);
xnor U11223 (N_11223,N_7275,N_8537);
nand U11224 (N_11224,N_6775,N_6340);
or U11225 (N_11225,N_9806,N_9022);
nor U11226 (N_11226,N_8652,N_5025);
xor U11227 (N_11227,N_5508,N_6037);
nor U11228 (N_11228,N_6254,N_5661);
or U11229 (N_11229,N_9049,N_8705);
and U11230 (N_11230,N_9344,N_8719);
nor U11231 (N_11231,N_9146,N_6565);
and U11232 (N_11232,N_6164,N_7376);
nand U11233 (N_11233,N_7470,N_5915);
nor U11234 (N_11234,N_9456,N_6530);
and U11235 (N_11235,N_8496,N_6728);
and U11236 (N_11236,N_9448,N_7893);
or U11237 (N_11237,N_8211,N_5194);
or U11238 (N_11238,N_7112,N_6118);
and U11239 (N_11239,N_6784,N_8110);
and U11240 (N_11240,N_8281,N_7809);
or U11241 (N_11241,N_7424,N_9929);
nor U11242 (N_11242,N_8799,N_8755);
and U11243 (N_11243,N_8093,N_6716);
nor U11244 (N_11244,N_9722,N_7862);
nor U11245 (N_11245,N_9787,N_7133);
nand U11246 (N_11246,N_7871,N_8575);
or U11247 (N_11247,N_8868,N_8189);
nor U11248 (N_11248,N_6898,N_8486);
nor U11249 (N_11249,N_5170,N_6656);
and U11250 (N_11250,N_7325,N_5715);
nand U11251 (N_11251,N_9307,N_7232);
nand U11252 (N_11252,N_5945,N_8733);
nor U11253 (N_11253,N_9276,N_7856);
nor U11254 (N_11254,N_6266,N_7344);
nor U11255 (N_11255,N_8338,N_8464);
xnor U11256 (N_11256,N_7780,N_8081);
or U11257 (N_11257,N_9692,N_5017);
and U11258 (N_11258,N_7220,N_9732);
and U11259 (N_11259,N_7063,N_9298);
nor U11260 (N_11260,N_7425,N_9111);
nand U11261 (N_11261,N_9318,N_8413);
or U11262 (N_11262,N_7032,N_6642);
and U11263 (N_11263,N_5451,N_8838);
nor U11264 (N_11264,N_8995,N_7392);
or U11265 (N_11265,N_8365,N_5440);
or U11266 (N_11266,N_6087,N_5060);
and U11267 (N_11267,N_9973,N_7206);
or U11268 (N_11268,N_6487,N_6019);
xor U11269 (N_11269,N_6344,N_9867);
nor U11270 (N_11270,N_8309,N_7793);
xor U11271 (N_11271,N_6557,N_6945);
or U11272 (N_11272,N_9353,N_7214);
nand U11273 (N_11273,N_7903,N_5594);
nand U11274 (N_11274,N_7824,N_8387);
xor U11275 (N_11275,N_8524,N_6511);
nor U11276 (N_11276,N_5271,N_9082);
and U11277 (N_11277,N_5049,N_5197);
nor U11278 (N_11278,N_8606,N_7945);
nor U11279 (N_11279,N_6202,N_6495);
nor U11280 (N_11280,N_7821,N_7975);
xnor U11281 (N_11281,N_8306,N_7768);
and U11282 (N_11282,N_8858,N_5161);
nor U11283 (N_11283,N_5051,N_9661);
nand U11284 (N_11284,N_6022,N_9645);
xor U11285 (N_11285,N_7387,N_5563);
or U11286 (N_11286,N_7704,N_5895);
or U11287 (N_11287,N_9205,N_6770);
xnor U11288 (N_11288,N_5965,N_5023);
nor U11289 (N_11289,N_8786,N_5603);
or U11290 (N_11290,N_6206,N_8151);
or U11291 (N_11291,N_6437,N_6098);
and U11292 (N_11292,N_8616,N_8998);
nor U11293 (N_11293,N_8427,N_5044);
or U11294 (N_11294,N_6771,N_8941);
and U11295 (N_11295,N_8191,N_5654);
nand U11296 (N_11296,N_5671,N_8433);
and U11297 (N_11297,N_7142,N_7070);
or U11298 (N_11298,N_6783,N_7475);
nor U11299 (N_11299,N_7961,N_9368);
xnor U11300 (N_11300,N_5142,N_6626);
xor U11301 (N_11301,N_9493,N_7267);
xnor U11302 (N_11302,N_6619,N_8298);
or U11303 (N_11303,N_6307,N_8260);
or U11304 (N_11304,N_7929,N_5867);
and U11305 (N_11305,N_6448,N_8997);
and U11306 (N_11306,N_6962,N_7675);
nor U11307 (N_11307,N_7902,N_5475);
or U11308 (N_11308,N_9027,N_9458);
and U11309 (N_11309,N_5810,N_7235);
xnor U11310 (N_11310,N_6011,N_8091);
or U11311 (N_11311,N_7252,N_6508);
xor U11312 (N_11312,N_9030,N_9153);
and U11313 (N_11313,N_8763,N_7720);
nand U11314 (N_11314,N_9641,N_5588);
nor U11315 (N_11315,N_7373,N_5949);
and U11316 (N_11316,N_8026,N_6589);
nor U11317 (N_11317,N_7523,N_8803);
xnor U11318 (N_11318,N_9162,N_8431);
xor U11319 (N_11319,N_8608,N_8398);
or U11320 (N_11320,N_6981,N_7247);
or U11321 (N_11321,N_6806,N_8045);
nand U11322 (N_11322,N_8788,N_6397);
nor U11323 (N_11323,N_9760,N_9536);
and U11324 (N_11324,N_9909,N_7131);
nor U11325 (N_11325,N_7937,N_8836);
or U11326 (N_11326,N_9815,N_6269);
and U11327 (N_11327,N_5785,N_6099);
nand U11328 (N_11328,N_6680,N_7526);
or U11329 (N_11329,N_7611,N_8707);
nand U11330 (N_11330,N_7381,N_9992);
xor U11331 (N_11331,N_9354,N_9364);
and U11332 (N_11332,N_6650,N_6485);
xnor U11333 (N_11333,N_8769,N_7140);
nand U11334 (N_11334,N_9231,N_9324);
nor U11335 (N_11335,N_9657,N_5100);
nand U11336 (N_11336,N_5326,N_8173);
nand U11337 (N_11337,N_6320,N_5031);
or U11338 (N_11338,N_8402,N_8724);
or U11339 (N_11339,N_9996,N_9881);
nand U11340 (N_11340,N_9991,N_6079);
nand U11341 (N_11341,N_9474,N_7174);
nor U11342 (N_11342,N_9366,N_5089);
nand U11343 (N_11343,N_6258,N_9113);
xor U11344 (N_11344,N_7160,N_8350);
and U11345 (N_11345,N_5314,N_8294);
nand U11346 (N_11346,N_5320,N_9738);
nor U11347 (N_11347,N_9886,N_7451);
or U11348 (N_11348,N_5564,N_8942);
or U11349 (N_11349,N_7855,N_9704);
or U11350 (N_11350,N_5730,N_5419);
nor U11351 (N_11351,N_6180,N_8586);
and U11352 (N_11352,N_8630,N_5107);
xor U11353 (N_11353,N_5868,N_7990);
xor U11354 (N_11354,N_7686,N_5180);
and U11355 (N_11355,N_5131,N_7517);
nand U11356 (N_11356,N_6309,N_8421);
xnor U11357 (N_11357,N_9278,N_6548);
and U11358 (N_11358,N_7269,N_6613);
xor U11359 (N_11359,N_8907,N_6195);
nor U11360 (N_11360,N_7305,N_6479);
and U11361 (N_11361,N_6584,N_9941);
nor U11362 (N_11362,N_5322,N_5476);
and U11363 (N_11363,N_8012,N_6066);
nand U11364 (N_11364,N_5224,N_7228);
nand U11365 (N_11365,N_6901,N_9718);
nor U11366 (N_11366,N_9280,N_9807);
xor U11367 (N_11367,N_5020,N_6798);
nor U11368 (N_11368,N_7234,N_7885);
nor U11369 (N_11369,N_6003,N_7927);
and U11370 (N_11370,N_9418,N_8504);
and U11371 (N_11371,N_6973,N_5606);
nand U11372 (N_11372,N_5216,N_6429);
nand U11373 (N_11373,N_7763,N_8841);
nor U11374 (N_11374,N_5673,N_6851);
or U11375 (N_11375,N_5446,N_8414);
nor U11376 (N_11376,N_9769,N_7051);
nor U11377 (N_11377,N_5323,N_9209);
and U11378 (N_11378,N_6759,N_6820);
and U11379 (N_11379,N_5449,N_7519);
nor U11380 (N_11380,N_6384,N_9979);
nand U11381 (N_11381,N_9195,N_6361);
and U11382 (N_11382,N_9553,N_6389);
or U11383 (N_11383,N_8311,N_7061);
xnor U11384 (N_11384,N_9316,N_5963);
nand U11385 (N_11385,N_9449,N_7163);
nand U11386 (N_11386,N_8333,N_9598);
nor U11387 (N_11387,N_5873,N_7564);
or U11388 (N_11388,N_9968,N_6142);
nand U11389 (N_11389,N_5301,N_9488);
xor U11390 (N_11390,N_5469,N_5818);
or U11391 (N_11391,N_6708,N_8619);
nand U11392 (N_11392,N_9279,N_8103);
nand U11393 (N_11393,N_6364,N_9319);
nor U11394 (N_11394,N_9517,N_9023);
nand U11395 (N_11395,N_6610,N_6544);
xor U11396 (N_11396,N_8768,N_8139);
and U11397 (N_11397,N_7207,N_9772);
xnor U11398 (N_11398,N_5720,N_8218);
nand U11399 (N_11399,N_9330,N_5321);
and U11400 (N_11400,N_8498,N_7922);
and U11401 (N_11401,N_9367,N_9052);
and U11402 (N_11402,N_5433,N_9606);
xnor U11403 (N_11403,N_6552,N_7410);
and U11404 (N_11404,N_7708,N_7149);
nand U11405 (N_11405,N_6227,N_9604);
or U11406 (N_11406,N_9770,N_9218);
or U11407 (N_11407,N_8122,N_9194);
nor U11408 (N_11408,N_7371,N_8478);
nand U11409 (N_11409,N_5707,N_9412);
nand U11410 (N_11410,N_9491,N_9716);
nor U11411 (N_11411,N_5171,N_9383);
nand U11412 (N_11412,N_5808,N_9134);
and U11413 (N_11413,N_7052,N_7529);
nand U11414 (N_11414,N_6541,N_8960);
or U11415 (N_11415,N_9951,N_5571);
and U11416 (N_11416,N_6064,N_7016);
nor U11417 (N_11417,N_7428,N_9601);
or U11418 (N_11418,N_7707,N_7869);
nand U11419 (N_11419,N_5365,N_8727);
nand U11420 (N_11420,N_8953,N_6293);
nand U11421 (N_11421,N_5573,N_6638);
and U11422 (N_11422,N_7158,N_9487);
nor U11423 (N_11423,N_7165,N_6582);
xnor U11424 (N_11424,N_5783,N_8011);
or U11425 (N_11425,N_8255,N_5473);
xor U11426 (N_11426,N_7683,N_6756);
nand U11427 (N_11427,N_9155,N_7967);
xnor U11428 (N_11428,N_6455,N_6187);
or U11429 (N_11429,N_6928,N_5182);
nor U11430 (N_11430,N_7176,N_9292);
or U11431 (N_11431,N_8287,N_6754);
xnor U11432 (N_11432,N_9812,N_6563);
xor U11433 (N_11433,N_9565,N_5392);
or U11434 (N_11434,N_7167,N_6979);
or U11435 (N_11435,N_6762,N_6424);
nor U11436 (N_11436,N_8456,N_5056);
or U11437 (N_11437,N_9163,N_9476);
and U11438 (N_11438,N_9848,N_8027);
nor U11439 (N_11439,N_6866,N_6986);
and U11440 (N_11440,N_8109,N_9907);
nand U11441 (N_11441,N_6212,N_7549);
nor U11442 (N_11442,N_9981,N_7604);
nand U11443 (N_11443,N_5740,N_8262);
xnor U11444 (N_11444,N_8740,N_5399);
xnor U11445 (N_11445,N_9507,N_7661);
nand U11446 (N_11446,N_8864,N_8057);
and U11447 (N_11447,N_9580,N_5951);
or U11448 (N_11448,N_6819,N_9019);
or U11449 (N_11449,N_7356,N_8855);
xor U11450 (N_11450,N_7161,N_8441);
nor U11451 (N_11451,N_5976,N_5855);
xnor U11452 (N_11452,N_7890,N_8277);
or U11453 (N_11453,N_8369,N_5382);
xnor U11454 (N_11454,N_7752,N_9959);
nor U11455 (N_11455,N_9337,N_7942);
nand U11456 (N_11456,N_6587,N_6895);
and U11457 (N_11457,N_6052,N_8730);
and U11458 (N_11458,N_8883,N_9808);
or U11459 (N_11459,N_9809,N_6347);
and U11460 (N_11460,N_9042,N_9539);
nor U11461 (N_11461,N_9668,N_6628);
or U11462 (N_11462,N_9340,N_6460);
nand U11463 (N_11463,N_9429,N_7767);
and U11464 (N_11464,N_5347,N_8882);
or U11465 (N_11465,N_9234,N_5884);
and U11466 (N_11466,N_8156,N_8780);
nand U11467 (N_11467,N_8892,N_7850);
nor U11468 (N_11468,N_7069,N_8657);
and U11469 (N_11469,N_9543,N_5222);
xor U11470 (N_11470,N_7691,N_8233);
xnor U11471 (N_11471,N_6408,N_6399);
and U11472 (N_11472,N_7585,N_7502);
nor U11473 (N_11473,N_9314,N_7906);
nand U11474 (N_11474,N_8221,N_5249);
nor U11475 (N_11475,N_8634,N_6779);
xor U11476 (N_11476,N_8293,N_5904);
nor U11477 (N_11477,N_5325,N_6513);
or U11478 (N_11478,N_9183,N_7073);
or U11479 (N_11479,N_8097,N_9883);
or U11480 (N_11480,N_9332,N_5871);
nor U11481 (N_11481,N_9864,N_8270);
nor U11482 (N_11482,N_8479,N_7363);
xnor U11483 (N_11483,N_7758,N_9041);
nand U11484 (N_11484,N_6214,N_6325);
and U11485 (N_11485,N_7812,N_6722);
nand U11486 (N_11486,N_8436,N_7202);
xnor U11487 (N_11487,N_7813,N_8417);
or U11488 (N_11488,N_7148,N_5894);
nand U11489 (N_11489,N_8675,N_5467);
and U11490 (N_11490,N_5717,N_8205);
nor U11491 (N_11491,N_5848,N_5058);
and U11492 (N_11492,N_8059,N_7572);
nand U11493 (N_11493,N_7711,N_5841);
nor U11494 (N_11494,N_9407,N_5111);
nand U11495 (N_11495,N_8199,N_9703);
xor U11496 (N_11496,N_6143,N_8633);
nor U11497 (N_11497,N_9813,N_7151);
nand U11498 (N_11498,N_7775,N_9009);
nand U11499 (N_11499,N_5727,N_8202);
and U11500 (N_11500,N_6596,N_9216);
and U11501 (N_11501,N_7734,N_8048);
xor U11502 (N_11502,N_5081,N_9184);
and U11503 (N_11503,N_6175,N_7482);
and U11504 (N_11504,N_6875,N_6270);
nor U11505 (N_11505,N_9080,N_9877);
nor U11506 (N_11506,N_9987,N_7309);
nor U11507 (N_11507,N_6516,N_6183);
and U11508 (N_11508,N_5734,N_8162);
or U11509 (N_11509,N_5143,N_5693);
or U11510 (N_11510,N_7345,N_9905);
xor U11511 (N_11511,N_7755,N_5462);
nor U11512 (N_11512,N_6665,N_5869);
and U11513 (N_11513,N_6401,N_8804);
and U11514 (N_11514,N_5207,N_5065);
or U11515 (N_11515,N_5786,N_5113);
nor U11516 (N_11516,N_5959,N_9508);
nand U11517 (N_11517,N_9312,N_8856);
and U11518 (N_11518,N_8241,N_7243);
or U11519 (N_11519,N_8985,N_8639);
and U11520 (N_11520,N_6704,N_7524);
nor U11521 (N_11521,N_6354,N_9339);
and U11522 (N_11522,N_5122,N_9647);
xnor U11523 (N_11523,N_7454,N_7443);
nor U11524 (N_11524,N_9994,N_7031);
or U11525 (N_11525,N_5254,N_7029);
nor U11526 (N_11526,N_8008,N_9632);
nand U11527 (N_11527,N_6670,N_9388);
nor U11528 (N_11528,N_5805,N_6543);
nand U11529 (N_11529,N_9608,N_6780);
nand U11530 (N_11530,N_5529,N_7908);
nor U11531 (N_11531,N_5512,N_7377);
xnor U11532 (N_11532,N_9497,N_5497);
nor U11533 (N_11533,N_9998,N_9313);
nor U11534 (N_11534,N_7274,N_6245);
nor U11535 (N_11535,N_9701,N_9302);
nor U11536 (N_11536,N_6778,N_6168);
or U11537 (N_11537,N_8598,N_7197);
or U11538 (N_11538,N_9574,N_7047);
or U11539 (N_11539,N_5719,N_7867);
xor U11540 (N_11540,N_6922,N_6157);
and U11541 (N_11541,N_8650,N_7514);
nand U11542 (N_11542,N_8015,N_9086);
xnor U11543 (N_11543,N_7369,N_6144);
and U11544 (N_11544,N_9044,N_9710);
nand U11545 (N_11545,N_6425,N_7740);
xnor U11546 (N_11546,N_8186,N_8745);
nand U11547 (N_11547,N_6026,N_6054);
and U11548 (N_11548,N_7992,N_8301);
and U11549 (N_11549,N_7313,N_5010);
or U11550 (N_11550,N_6222,N_8980);
nor U11551 (N_11551,N_6925,N_9655);
nor U11552 (N_11552,N_7261,N_9917);
or U11553 (N_11553,N_6705,N_7102);
nand U11554 (N_11554,N_7132,N_8502);
nor U11555 (N_11555,N_5660,N_9875);
and U11556 (N_11556,N_6578,N_7515);
nand U11557 (N_11557,N_5132,N_6599);
or U11558 (N_11558,N_6929,N_8582);
nand U11559 (N_11559,N_9177,N_5046);
and U11560 (N_11560,N_8974,N_8349);
and U11561 (N_11561,N_8900,N_9046);
nor U11562 (N_11562,N_6211,N_6440);
nand U11563 (N_11563,N_9870,N_9499);
xnor U11564 (N_11564,N_8971,N_8236);
or U11565 (N_11565,N_7448,N_8234);
nand U11566 (N_11566,N_5905,N_7725);
nand U11567 (N_11567,N_5750,N_8112);
nor U11568 (N_11568,N_6970,N_5575);
nand U11569 (N_11569,N_5116,N_7062);
nand U11570 (N_11570,N_7386,N_5196);
nand U11571 (N_11571,N_7602,N_8683);
and U11572 (N_11572,N_6863,N_9149);
xor U11573 (N_11573,N_5457,N_5483);
xnor U11574 (N_11574,N_9071,N_8552);
nor U11575 (N_11575,N_5970,N_8258);
and U11576 (N_11576,N_7213,N_8809);
and U11577 (N_11577,N_8708,N_5655);
nor U11578 (N_11578,N_6944,N_7733);
and U11579 (N_11579,N_6463,N_5658);
nor U11580 (N_11580,N_7494,N_7485);
or U11581 (N_11581,N_5978,N_8149);
nor U11582 (N_11582,N_5711,N_9283);
or U11583 (N_11583,N_5357,N_8916);
or U11584 (N_11584,N_6622,N_6799);
nand U11585 (N_11585,N_5103,N_8220);
nand U11586 (N_11586,N_8013,N_6257);
and U11587 (N_11587,N_9561,N_9078);
nand U11588 (N_11588,N_8061,N_6200);
nand U11589 (N_11589,N_8558,N_7053);
or U11590 (N_11590,N_9122,N_7597);
nand U11591 (N_11591,N_8966,N_5620);
or U11592 (N_11592,N_5559,N_9931);
nor U11593 (N_11593,N_9793,N_7382);
nor U11594 (N_11594,N_5989,N_8344);
xor U11595 (N_11595,N_5003,N_8989);
or U11596 (N_11596,N_7742,N_8594);
nand U11597 (N_11597,N_8661,N_7396);
nand U11598 (N_11598,N_8503,N_9083);
and U11599 (N_11599,N_9026,N_9902);
or U11600 (N_11600,N_8638,N_9833);
and U11601 (N_11601,N_8446,N_9288);
or U11602 (N_11602,N_5534,N_6398);
nand U11603 (N_11603,N_7931,N_9175);
nor U11604 (N_11604,N_6367,N_8746);
and U11605 (N_11605,N_6420,N_7607);
xor U11606 (N_11606,N_5682,N_7145);
nand U11607 (N_11607,N_8579,N_5791);
nand U11608 (N_11608,N_7065,N_7545);
nand U11609 (N_11609,N_9725,N_9137);
or U11610 (N_11610,N_8817,N_9627);
or U11611 (N_11611,N_9839,N_8918);
nand U11612 (N_11612,N_5814,N_5675);
xnor U11613 (N_11613,N_9001,N_5732);
nand U11614 (N_11614,N_6336,N_7353);
nor U11615 (N_11615,N_7402,N_7456);
nor U11616 (N_11616,N_8039,N_9680);
nand U11617 (N_11617,N_7727,N_8308);
nor U11618 (N_11618,N_5768,N_7626);
xor U11619 (N_11619,N_6484,N_6498);
nand U11620 (N_11620,N_9955,N_6504);
nor U11621 (N_11621,N_7236,N_9356);
nand U11622 (N_11622,N_9013,N_6720);
or U11623 (N_11623,N_5885,N_8825);
and U11624 (N_11624,N_9239,N_8332);
and U11625 (N_11625,N_8022,N_9570);
or U11626 (N_11626,N_5920,N_7139);
and U11627 (N_11627,N_9271,N_5169);
and U11628 (N_11628,N_5828,N_5971);
and U11629 (N_11629,N_5465,N_6147);
nor U11630 (N_11630,N_6580,N_9097);
xor U11631 (N_11631,N_5075,N_8230);
xnor U11632 (N_11632,N_8829,N_9810);
nand U11633 (N_11633,N_7483,N_9635);
nand U11634 (N_11634,N_9750,N_6488);
nor U11635 (N_11635,N_5424,N_8150);
xor U11636 (N_11636,N_5461,N_7179);
or U11637 (N_11637,N_8017,N_7129);
nor U11638 (N_11638,N_6020,N_8710);
and U11639 (N_11639,N_8462,N_8376);
nor U11640 (N_11640,N_9675,N_9031);
nand U11641 (N_11641,N_8450,N_6117);
or U11642 (N_11642,N_6746,N_6734);
nor U11643 (N_11643,N_7196,N_5225);
nor U11644 (N_11644,N_6989,N_6857);
and U11645 (N_11645,N_7662,N_5589);
or U11646 (N_11646,N_5052,N_6432);
xnor U11647 (N_11647,N_9584,N_7673);
xor U11648 (N_11648,N_9914,N_8863);
nand U11649 (N_11649,N_7298,N_5275);
and U11650 (N_11650,N_6494,N_7461);
xnor U11651 (N_11651,N_8286,N_6410);
nand U11652 (N_11652,N_8629,N_7873);
nand U11653 (N_11653,N_6445,N_5096);
xor U11654 (N_11654,N_9156,N_7060);
and U11655 (N_11655,N_8601,N_8536);
and U11656 (N_11656,N_6926,N_5505);
and U11657 (N_11657,N_6905,N_5804);
xor U11658 (N_11658,N_5751,N_6932);
and U11659 (N_11659,N_8158,N_9669);
nand U11660 (N_11660,N_7825,N_5394);
or U11661 (N_11661,N_8159,N_7503);
xor U11662 (N_11662,N_6467,N_6517);
xnor U11663 (N_11663,N_5708,N_8160);
xnor U11664 (N_11664,N_9846,N_8078);
nand U11665 (N_11665,N_8818,N_6707);
and U11666 (N_11666,N_8877,N_6196);
nor U11667 (N_11667,N_5986,N_8245);
and U11668 (N_11668,N_9698,N_8047);
xnor U11669 (N_11669,N_6955,N_6228);
or U11670 (N_11670,N_9245,N_7938);
and U11671 (N_11671,N_7781,N_5547);
nand U11672 (N_11672,N_5286,N_8254);
and U11673 (N_11673,N_7181,N_7121);
xor U11674 (N_11674,N_7000,N_5359);
xnor U11675 (N_11675,N_6917,N_9005);
or U11676 (N_11676,N_9390,N_7499);
and U11677 (N_11677,N_6191,N_7372);
and U11678 (N_11678,N_6464,N_8761);
xnor U11679 (N_11679,N_5992,N_5709);
xor U11680 (N_11680,N_7951,N_8774);
nor U11681 (N_11681,N_8430,N_8566);
xnor U11682 (N_11682,N_8176,N_7434);
and U11683 (N_11683,N_9266,N_6248);
or U11684 (N_11684,N_7375,N_5000);
nand U11685 (N_11685,N_8329,N_5900);
and U11686 (N_11686,N_5362,N_7351);
or U11687 (N_11687,N_9595,N_8878);
nor U11688 (N_11688,N_7530,N_6051);
and U11689 (N_11689,N_5285,N_6657);
nor U11690 (N_11690,N_7666,N_7761);
or U11691 (N_11691,N_6633,N_6528);
and U11692 (N_11692,N_8748,N_6993);
nand U11693 (N_11693,N_5408,N_6070);
nor U11694 (N_11694,N_8758,N_7857);
nor U11695 (N_11695,N_7256,N_7465);
nand U11696 (N_11696,N_6891,N_5415);
nor U11697 (N_11697,N_7724,N_9552);
xnor U11698 (N_11698,N_5593,N_6537);
or U11699 (N_11699,N_6476,N_6283);
nor U11700 (N_11700,N_8437,N_7573);
and U11701 (N_11701,N_5724,N_6412);
nor U11702 (N_11702,N_9123,N_9496);
and U11703 (N_11703,N_5396,N_8957);
or U11704 (N_11704,N_5982,N_7050);
xor U11705 (N_11705,N_9025,N_8408);
nor U11706 (N_11706,N_5611,N_5507);
and U11707 (N_11707,N_7658,N_7672);
or U11708 (N_11708,N_9322,N_5329);
xor U11709 (N_11709,N_9747,N_8666);
xor U11710 (N_11710,N_5077,N_6689);
and U11711 (N_11711,N_6630,N_8701);
and U11712 (N_11712,N_5317,N_5893);
and U11713 (N_11713,N_6992,N_7718);
and U11714 (N_11714,N_5289,N_5173);
xnor U11715 (N_11715,N_8315,N_9624);
nor U11716 (N_11716,N_5187,N_5312);
and U11717 (N_11717,N_9369,N_6210);
xor U11718 (N_11718,N_6298,N_7930);
and U11719 (N_11719,N_8167,N_8909);
xnor U11720 (N_11720,N_9181,N_5610);
xor U11721 (N_11721,N_7044,N_9821);
and U11722 (N_11722,N_9267,N_9967);
xor U11723 (N_11723,N_6012,N_5639);
nor U11724 (N_11724,N_6406,N_6743);
and U11725 (N_11725,N_8977,N_5421);
nor U11726 (N_11726,N_7393,N_9927);
xor U11727 (N_11727,N_6174,N_7790);
or U11728 (N_11728,N_7320,N_9786);
or U11729 (N_11729,N_7146,N_5228);
xnor U11730 (N_11730,N_6808,N_5336);
or U11731 (N_11731,N_7332,N_5248);
nand U11732 (N_11732,N_8307,N_5189);
nor U11733 (N_11733,N_8243,N_6750);
xnor U11734 (N_11734,N_6726,N_8676);
or U11735 (N_11735,N_5053,N_8567);
xor U11736 (N_11736,N_8085,N_5584);
nand U11737 (N_11737,N_5099,N_9274);
nand U11738 (N_11738,N_7327,N_9077);
and U11739 (N_11739,N_9430,N_9509);
and U11740 (N_11740,N_9977,N_5448);
nor U11741 (N_11741,N_6034,N_9551);
and U11742 (N_11742,N_8372,N_5192);
xor U11743 (N_11743,N_7865,N_8744);
nand U11744 (N_11744,N_5144,N_8706);
and U11745 (N_11745,N_5478,N_5339);
nand U11746 (N_11746,N_5834,N_6652);
nor U11747 (N_11747,N_5247,N_8386);
xnor U11748 (N_11748,N_6383,N_7059);
or U11749 (N_11749,N_6574,N_9798);
xnor U11750 (N_11750,N_7971,N_6396);
nor U11751 (N_11751,N_6634,N_9148);
nor U11752 (N_11752,N_5906,N_9229);
nand U11753 (N_11753,N_7586,N_5147);
nor U11754 (N_11754,N_8627,N_9948);
nor U11755 (N_11755,N_8251,N_8409);
and U11756 (N_11756,N_7568,N_7037);
and U11757 (N_11757,N_6871,N_8232);
or U11758 (N_11758,N_7935,N_5274);
or U11759 (N_11759,N_6434,N_8343);
nand U11760 (N_11760,N_6262,N_5624);
nand U11761 (N_11761,N_5265,N_9741);
nand U11762 (N_11762,N_6546,N_5913);
or U11763 (N_11763,N_7991,N_9630);
nand U11764 (N_11764,N_6703,N_6838);
xor U11765 (N_11765,N_5119,N_6940);
xor U11766 (N_11766,N_9090,N_5781);
xor U11767 (N_11767,N_5370,N_9347);
and U11768 (N_11768,N_5160,N_9211);
nor U11769 (N_11769,N_7366,N_7030);
nor U11770 (N_11770,N_8767,N_7735);
and U11771 (N_11771,N_7033,N_5054);
or U11772 (N_11772,N_8130,N_7531);
and U11773 (N_11773,N_7912,N_6870);
nand U11774 (N_11774,N_7655,N_8888);
or U11775 (N_11775,N_8348,N_6727);
and U11776 (N_11776,N_8297,N_6807);
or U11777 (N_11777,N_9729,N_9748);
and U11778 (N_11778,N_5108,N_8988);
nor U11779 (N_11779,N_7452,N_6908);
nor U11780 (N_11780,N_5570,N_6951);
xnor U11781 (N_11781,N_5220,N_5281);
xnor U11782 (N_11782,N_5934,N_7966);
nand U11783 (N_11783,N_7960,N_6135);
xnor U11784 (N_11784,N_6577,N_8874);
and U11785 (N_11785,N_9666,N_6911);
nor U11786 (N_11786,N_6984,N_9612);
and U11787 (N_11787,N_5384,N_8448);
nor U11788 (N_11788,N_8422,N_6435);
xnor U11789 (N_11789,N_6964,N_8715);
and U11790 (N_11790,N_7435,N_7841);
and U11791 (N_11791,N_5674,N_6349);
or U11792 (N_11792,N_6607,N_6386);
or U11793 (N_11793,N_6949,N_6741);
nand U11794 (N_11794,N_6894,N_6140);
nand U11795 (N_11795,N_9631,N_6010);
or U11796 (N_11796,N_7048,N_7609);
and U11797 (N_11797,N_7685,N_6617);
and U11798 (N_11798,N_9737,N_7599);
and U11799 (N_11799,N_8115,N_5846);
nor U11800 (N_11800,N_9417,N_6130);
and U11801 (N_11801,N_8244,N_6042);
and U11802 (N_11802,N_5578,N_8669);
nor U11803 (N_11803,N_6801,N_5028);
nor U11804 (N_11804,N_8389,N_8068);
xnor U11805 (N_11805,N_8001,N_7300);
nor U11806 (N_11806,N_7640,N_7223);
nor U11807 (N_11807,N_8550,N_7913);
nor U11808 (N_11808,N_6025,N_7203);
nand U11809 (N_11809,N_5831,N_8523);
nor U11810 (N_11810,N_7822,N_7567);
nor U11811 (N_11811,N_7011,N_6322);
and U11812 (N_11812,N_9745,N_5027);
and U11813 (N_11813,N_8959,N_8305);
and U11814 (N_11814,N_5299,N_6809);
or U11815 (N_11815,N_6752,N_7964);
and U11816 (N_11816,N_9838,N_7543);
nor U11817 (N_11817,N_9784,N_8264);
xnor U11818 (N_11818,N_7459,N_8342);
and U11819 (N_11819,N_7947,N_7949);
xnor U11820 (N_11820,N_6812,N_9281);
or U11821 (N_11821,N_5923,N_9609);
nor U11822 (N_11822,N_5948,N_5889);
or U11823 (N_11823,N_5070,N_7979);
and U11824 (N_11824,N_9762,N_5939);
nor U11825 (N_11825,N_9926,N_9303);
xnor U11826 (N_11826,N_7888,N_8852);
nand U11827 (N_11827,N_9687,N_7087);
xnor U11828 (N_11828,N_7318,N_8195);
xnor U11829 (N_11829,N_6572,N_7374);
nor U11830 (N_11830,N_6133,N_9378);
xor U11831 (N_11831,N_9757,N_8304);
and U11832 (N_11832,N_6682,N_9202);
xor U11833 (N_11833,N_5351,N_7312);
and U11834 (N_11834,N_8217,N_7019);
and U11835 (N_11835,N_6792,N_7278);
nor U11836 (N_11836,N_5500,N_7490);
and U11837 (N_11837,N_5902,N_9975);
or U11838 (N_11838,N_7043,N_7397);
nor U11839 (N_11839,N_6182,N_8603);
nand U11840 (N_11840,N_7323,N_5200);
nand U11841 (N_11841,N_5685,N_8790);
and U11842 (N_11842,N_8352,N_5776);
xor U11843 (N_11843,N_7627,N_7199);
nor U11844 (N_11844,N_9628,N_9556);
xnor U11845 (N_11845,N_8470,N_5853);
nand U11846 (N_11846,N_6692,N_7674);
xor U11847 (N_11847,N_7389,N_9726);
or U11848 (N_11848,N_8488,N_8257);
and U11849 (N_11849,N_6299,N_9285);
nand U11850 (N_11850,N_5929,N_6585);
or U11851 (N_11851,N_6560,N_8548);
or U11852 (N_11852,N_9823,N_8922);
and U11853 (N_11853,N_5821,N_9742);
xor U11854 (N_11854,N_5432,N_6426);
and U11855 (N_11855,N_6691,N_5861);
xnor U11856 (N_11856,N_8107,N_9103);
xor U11857 (N_11857,N_8276,N_7789);
xnor U11858 (N_11858,N_5102,N_8931);
and U11859 (N_11859,N_9235,N_5269);
and U11860 (N_11860,N_6958,N_6379);
nor U11861 (N_11861,N_9460,N_6492);
nor U11862 (N_11862,N_9482,N_9120);
nor U11863 (N_11863,N_7395,N_8520);
nor U11864 (N_11864,N_6735,N_8334);
and U11865 (N_11865,N_6687,N_5987);
nand U11866 (N_11866,N_8802,N_9707);
xnor U11867 (N_11867,N_8896,N_6943);
xnor U11868 (N_11868,N_6473,N_6236);
and U11869 (N_11869,N_8653,N_7426);
nand U11870 (N_11870,N_6339,N_8325);
or U11871 (N_11871,N_7952,N_8830);
nand U11872 (N_11872,N_6725,N_8021);
or U11873 (N_11873,N_6134,N_9178);
xnor U11874 (N_11874,N_9566,N_5211);
or U11875 (N_11875,N_5295,N_5994);
nor U11876 (N_11876,N_9345,N_5926);
and U11877 (N_11877,N_9058,N_9836);
and U11878 (N_11878,N_6673,N_9910);
or U11879 (N_11879,N_8131,N_6148);
nor U11880 (N_11880,N_7110,N_7385);
nand U11881 (N_11881,N_9616,N_9739);
or U11882 (N_11882,N_9036,N_9557);
nand U11883 (N_11883,N_6739,N_7907);
and U11884 (N_11884,N_5950,N_7505);
nor U11885 (N_11885,N_5068,N_8354);
and U11886 (N_11886,N_9989,N_6889);
and U11887 (N_11887,N_8378,N_9461);
nor U11888 (N_11888,N_5367,N_5217);
xnor U11889 (N_11889,N_9997,N_7748);
or U11890 (N_11890,N_9118,N_5996);
or U11891 (N_11891,N_9849,N_9882);
nand U11892 (N_11892,N_6430,N_8645);
nand U11893 (N_11893,N_5742,N_9243);
nand U11894 (N_11894,N_5340,N_8910);
and U11895 (N_11895,N_7101,N_8272);
nor U11896 (N_11896,N_6273,N_7276);
nor U11897 (N_11897,N_8416,N_6104);
nor U11898 (N_11898,N_9173,N_7703);
and U11899 (N_11899,N_5226,N_7420);
or U11900 (N_11900,N_8833,N_6496);
nand U11901 (N_11901,N_7124,N_9858);
and U11902 (N_11902,N_6608,N_7250);
and U11903 (N_11903,N_6362,N_9179);
nand U11904 (N_11904,N_7847,N_5472);
nand U11905 (N_11905,N_9419,N_7722);
nand U11906 (N_11906,N_7957,N_8447);
xor U11907 (N_11907,N_8897,N_5209);
or U11908 (N_11908,N_6007,N_6842);
xor U11909 (N_11909,N_9541,N_5960);
nand U11910 (N_11910,N_6671,N_5062);
and U11911 (N_11911,N_5520,N_5897);
nand U11912 (N_11912,N_6313,N_6241);
and U11913 (N_11913,N_8113,N_9899);
nand U11914 (N_11914,N_9436,N_8487);
xnor U11915 (N_11915,N_6021,N_5157);
xor U11916 (N_11916,N_8237,N_9962);
xor U11917 (N_11917,N_6611,N_5183);
nor U11918 (N_11918,N_6659,N_6499);
xor U11919 (N_11919,N_5579,N_9945);
or U11920 (N_11920,N_8813,N_5026);
or U11921 (N_11921,N_6275,N_7820);
nand U11922 (N_11922,N_6841,N_5585);
xnor U11923 (N_11923,N_6005,N_6934);
xnor U11924 (N_11924,N_7178,N_5260);
nand U11925 (N_11925,N_5034,N_9011);
or U11926 (N_11926,N_6438,N_7194);
or U11927 (N_11927,N_5723,N_9796);
nand U11928 (N_11928,N_7799,N_6279);
nand U11929 (N_11929,N_5091,N_9916);
nand U11930 (N_11930,N_6243,N_6667);
nand U11931 (N_11931,N_5159,N_9055);
nand U11932 (N_11932,N_7355,N_5605);
or U11933 (N_11933,N_9753,N_5835);
or U11934 (N_11934,N_8457,N_6409);
and U11935 (N_11935,N_8869,N_7416);
or U11936 (N_11936,N_7316,N_8371);
or U11937 (N_11937,N_9447,N_7677);
xnor U11938 (N_11938,N_6207,N_6129);
nor U11939 (N_11939,N_8163,N_6961);
and U11940 (N_11940,N_6158,N_6737);
xnor U11941 (N_11941,N_6931,N_9441);
and U11942 (N_11942,N_5936,N_5901);
and U11943 (N_11943,N_5355,N_8269);
or U11944 (N_11944,N_7736,N_6843);
nand U11945 (N_11945,N_9567,N_9438);
xor U11946 (N_11946,N_6304,N_9210);
xor U11947 (N_11947,N_5393,N_6884);
and U11948 (N_11948,N_9938,N_8458);
or U11949 (N_11949,N_9477,N_5087);
nor U11950 (N_11950,N_7614,N_9672);
nor U11951 (N_11951,N_8072,N_7117);
nor U11952 (N_11952,N_5754,N_5733);
nor U11953 (N_11953,N_5436,N_9603);
or U11954 (N_11954,N_5700,N_8992);
nand U11955 (N_11955,N_7551,N_7914);
nor U11956 (N_11956,N_6356,N_8492);
nor U11957 (N_11957,N_6382,N_6318);
and U11958 (N_11958,N_7625,N_9125);
nor U11959 (N_11959,N_6287,N_9665);
xnor U11960 (N_11960,N_8393,N_5677);
xor U11961 (N_11961,N_5361,N_7442);
and U11962 (N_11962,N_7342,N_7537);
nand U11963 (N_11963,N_6581,N_8377);
nand U11964 (N_11964,N_5784,N_7721);
xor U11965 (N_11965,N_6540,N_5195);
nor U11966 (N_11966,N_5801,N_6305);
nor U11967 (N_11967,N_8517,N_7827);
or U11968 (N_11968,N_5644,N_7328);
and U11969 (N_11969,N_9402,N_7880);
xor U11970 (N_11970,N_8873,N_8200);
and U11971 (N_11971,N_9731,N_6663);
nor U11972 (N_11972,N_7496,N_8179);
nand U11973 (N_11973,N_7954,N_9050);
xor U11974 (N_11974,N_7534,N_6139);
and U11975 (N_11975,N_8798,N_8227);
nand U11976 (N_11976,N_5136,N_6306);
nand U11977 (N_11977,N_5592,N_9573);
xor U11978 (N_11978,N_9501,N_8689);
xor U11979 (N_11979,N_5940,N_7884);
and U11980 (N_11980,N_7507,N_5659);
and U11981 (N_11981,N_9007,N_6921);
and U11982 (N_11982,N_8990,N_8981);
and U11983 (N_11983,N_6056,N_8741);
and U11984 (N_11984,N_7090,N_8482);
nand U11985 (N_11985,N_6291,N_9844);
and U11986 (N_11986,N_8936,N_6116);
xor U11987 (N_11987,N_5324,N_9915);
nor U11988 (N_11988,N_8806,N_8765);
and U11989 (N_11989,N_9596,N_9511);
nand U11990 (N_11990,N_7364,N_7639);
and U11991 (N_11991,N_9837,N_8432);
xor U11992 (N_11992,N_7201,N_5553);
xnor U11993 (N_11993,N_7343,N_9980);
or U11994 (N_11994,N_6669,N_9190);
nand U11995 (N_11995,N_8438,N_8734);
nor U11996 (N_11996,N_5383,N_7204);
xor U11997 (N_11997,N_6785,N_8215);
nor U11998 (N_11998,N_7828,N_9908);
or U11999 (N_11999,N_5634,N_9713);
nand U12000 (N_12000,N_7962,N_7923);
xnor U12001 (N_12001,N_6123,N_8018);
and U12002 (N_12002,N_7134,N_7940);
nor U12003 (N_12003,N_6327,N_8890);
or U12004 (N_12004,N_6141,N_6976);
nand U12005 (N_12005,N_7845,N_9581);
nand U12006 (N_12006,N_9207,N_9212);
and U12007 (N_12007,N_6334,N_7615);
nor U12008 (N_12008,N_6188,N_7168);
or U12009 (N_12009,N_9494,N_5373);
xnor U12010 (N_12010,N_5450,N_9845);
xor U12011 (N_12011,N_9481,N_5918);
and U12012 (N_12012,N_8738,N_6923);
nor U12013 (N_12013,N_6590,N_8560);
nor U12014 (N_12014,N_9060,N_8460);
or U12015 (N_12015,N_9988,N_9650);
xnor U12016 (N_12016,N_6326,N_7212);
and U12017 (N_12017,N_6568,N_9469);
and U12018 (N_12018,N_8760,N_5403);
and U12019 (N_12019,N_6939,N_9964);
or U12020 (N_12020,N_5344,N_8797);
nor U12021 (N_12021,N_9691,N_8742);
nand U12022 (N_12022,N_5645,N_9021);
xnor U12023 (N_12023,N_6393,N_6533);
and U12024 (N_12024,N_9744,N_6385);
nand U12025 (N_12025,N_8127,N_5252);
or U12026 (N_12026,N_8721,N_8235);
nor U12027 (N_12027,N_7801,N_8913);
and U12028 (N_12028,N_6781,N_7285);
nand U12029 (N_12029,N_7020,N_5619);
nor U12030 (N_12030,N_6514,N_8534);
and U12031 (N_12031,N_6916,N_9466);
nand U12032 (N_12032,N_6447,N_6209);
or U12033 (N_12033,N_9422,N_9428);
xor U12034 (N_12034,N_6402,N_8224);
or U12035 (N_12035,N_6418,N_8454);
and U12036 (N_12036,N_5837,N_9408);
nor U12037 (N_12037,N_6321,N_6751);
and U12038 (N_12038,N_7097,N_7273);
nor U12039 (N_12039,N_7898,N_9327);
nand U12040 (N_12040,N_9228,N_9746);
nand U12041 (N_12041,N_7915,N_6374);
nor U12042 (N_12042,N_6616,N_8880);
xor U12043 (N_12043,N_8546,N_5037);
or U12044 (N_12044,N_5748,N_9093);
xnor U12045 (N_12045,N_7135,N_6301);
and U12046 (N_12046,N_8032,N_7969);
nor U12047 (N_12047,N_9705,N_6828);
nand U12048 (N_12048,N_9841,N_9542);
nand U12049 (N_12049,N_5300,N_7687);
xor U12050 (N_12050,N_9597,N_9348);
or U12051 (N_12051,N_7939,N_6840);
and U12052 (N_12052,N_6643,N_9860);
nor U12053 (N_12053,N_6713,N_7959);
and U12054 (N_12054,N_6215,N_9085);
nor U12055 (N_12055,N_9610,N_7463);
nor U12056 (N_12056,N_5166,N_9321);
or U12057 (N_12057,N_5910,N_5690);
xor U12058 (N_12058,N_7497,N_7340);
xor U12059 (N_12059,N_7521,N_7853);
or U12060 (N_12060,N_5241,N_7153);
xnor U12061 (N_12061,N_7150,N_6903);
nor U12062 (N_12062,N_5973,N_6731);
xor U12063 (N_12063,N_9119,N_9674);
or U12064 (N_12064,N_7559,N_6592);
nand U12065 (N_12065,N_9727,N_8628);
nor U12066 (N_12066,N_8005,N_9295);
nor U12067 (N_12067,N_6721,N_6844);
or U12068 (N_12068,N_8108,N_6068);
xnor U12069 (N_12069,N_7458,N_7156);
or U12070 (N_12070,N_5576,N_7317);
xnor U12071 (N_12071,N_7868,N_6089);
nand U12072 (N_12072,N_8096,N_8300);
nand U12073 (N_12073,N_7486,N_8050);
or U12074 (N_12074,N_6107,N_6395);
nor U12075 (N_12075,N_9797,N_6073);
or U12076 (N_12076,N_9406,N_7883);
and U12077 (N_12077,N_5924,N_8445);
nor U12078 (N_12078,N_8038,N_5532);
and U12079 (N_12079,N_8968,N_7489);
nor U12080 (N_12080,N_5856,N_8665);
xor U12081 (N_12081,N_8400,N_5692);
nand U12082 (N_12082,N_6661,N_9372);
or U12083 (N_12083,N_5251,N_5413);
or U12084 (N_12084,N_5405,N_8368);
and U12085 (N_12085,N_8174,N_6649);
and U12086 (N_12086,N_6745,N_7418);
or U12087 (N_12087,N_7579,N_8648);
nor U12088 (N_12088,N_6431,N_7652);
nand U12089 (N_12089,N_7760,N_8623);
and U12090 (N_12090,N_9547,N_5536);
nor U12091 (N_12091,N_9128,N_5509);
nor U12092 (N_12092,N_6451,N_8924);
or U12093 (N_12093,N_7286,N_6772);
xnor U12094 (N_12094,N_8512,N_5327);
and U12095 (N_12095,N_9328,N_6404);
xor U12096 (N_12096,N_5380,N_6835);
or U12097 (N_12097,N_7819,N_7620);
or U12098 (N_12098,N_8303,N_5276);
nand U12099 (N_12099,N_5865,N_8412);
and U12100 (N_12100,N_8483,N_9214);
or U12101 (N_12101,N_8095,N_5460);
nand U12102 (N_12102,N_6378,N_9736);
nand U12103 (N_12103,N_8094,N_9191);
nand U12104 (N_12104,N_9564,N_7003);
nand U12105 (N_12105,N_8861,N_7399);
nand U12106 (N_12106,N_8857,N_8036);
xor U12107 (N_12107,N_7464,N_6050);
or U12108 (N_12108,N_8118,N_9660);
or U12109 (N_12109,N_9546,N_5778);
and U12110 (N_12110,N_8972,N_5829);
nand U12111 (N_12111,N_6983,N_7441);
nand U12112 (N_12112,N_9733,N_5236);
nand U12113 (N_12113,N_5561,N_9306);
xor U12114 (N_12114,N_6324,N_9384);
and U12115 (N_12115,N_9404,N_5310);
xor U12116 (N_12116,N_8449,N_9947);
nor U12117 (N_12117,N_9201,N_5128);
and U12118 (N_12118,N_6629,N_9826);
and U12119 (N_12119,N_9885,N_7587);
or U12120 (N_12120,N_8034,N_8497);
nor U12121 (N_12121,N_5916,N_8805);
or U12122 (N_12122,N_7433,N_9326);
and U12123 (N_12123,N_6348,N_9182);
xnor U12124 (N_12124,N_8326,N_7113);
or U12125 (N_12125,N_7840,N_6030);
xnor U12126 (N_12126,N_6252,N_7103);
and U12127 (N_12127,N_6868,N_9098);
nor U12128 (N_12128,N_7306,N_6112);
xnor U12129 (N_12129,N_7347,N_7693);
and U12130 (N_12130,N_5426,N_5098);
nor U12131 (N_12131,N_8720,N_8066);
nand U12132 (N_12132,N_8781,N_7741);
nor U12133 (N_12133,N_7023,N_8016);
nor U12134 (N_12134,N_7621,N_9192);
or U12135 (N_12135,N_9185,N_8395);
nor U12136 (N_12136,N_6272,N_5790);
or U12137 (N_12137,N_6876,N_5316);
nor U12138 (N_12138,N_8146,N_8692);
xnor U12139 (N_12139,N_9391,N_9751);
nor U12140 (N_12140,N_8905,N_8071);
or U12141 (N_12141,N_9048,N_5626);
or U12142 (N_12142,N_9663,N_8428);
nor U12143 (N_12143,N_5291,N_5663);
nor U12144 (N_12144,N_8345,N_6162);
xor U12145 (N_12145,N_6353,N_6071);
and U12146 (N_12146,N_9586,N_8063);
xor U12147 (N_12147,N_5714,N_5713);
or U12148 (N_12148,N_5431,N_9453);
or U12149 (N_12149,N_7522,N_5985);
or U12150 (N_12150,N_9633,N_6815);
nor U12151 (N_12151,N_9530,N_5202);
nor U12152 (N_12152,N_6450,N_5590);
nand U12153 (N_12153,N_8111,N_5803);
and U12154 (N_12154,N_5235,N_8547);
nor U12155 (N_12155,N_9505,N_7701);
or U12156 (N_12156,N_6265,N_7085);
nor U12157 (N_12157,N_8789,N_9107);
and U12158 (N_12158,N_8640,N_7078);
xor U12159 (N_12159,N_9403,N_9475);
and U12160 (N_12160,N_7697,N_7082);
and U12161 (N_12161,N_5374,N_8726);
and U12162 (N_12162,N_7105,N_6419);
and U12163 (N_12163,N_6417,N_9237);
or U12164 (N_12164,N_7504,N_9528);
nor U12165 (N_12165,N_6095,N_8895);
and U12166 (N_12166,N_7431,N_8074);
nor U12167 (N_12167,N_9133,N_8847);
xnor U12168 (N_12168,N_9588,N_5699);
nand U12169 (N_12169,N_9863,N_7349);
xor U12170 (N_12170,N_9946,N_9652);
or U12171 (N_12171,N_5284,N_5647);
xnor U12172 (N_12172,N_7633,N_9702);
or U12173 (N_12173,N_7696,N_8420);
or U12174 (N_12174,N_8198,N_6846);
nor U12175 (N_12175,N_7535,N_9811);
or U12176 (N_12176,N_8578,N_6346);
or U12177 (N_12177,N_9084,N_7796);
nor U12178 (N_12178,N_7076,N_5676);
nand U12179 (N_12179,N_5851,N_7613);
and U12180 (N_12180,N_7844,N_5550);
and U12181 (N_12181,N_6303,N_7096);
and U12182 (N_12182,N_8065,N_5007);
and U12183 (N_12183,N_8674,N_9884);
xnor U12184 (N_12184,N_8731,N_9895);
and U12185 (N_12185,N_6233,N_5574);
xnor U12186 (N_12186,N_7222,N_6631);
xnor U12187 (N_12187,N_5391,N_9579);
or U12188 (N_12188,N_7400,N_5133);
and U12189 (N_12189,N_6644,N_8128);
nor U12190 (N_12190,N_6296,N_9506);
and U12191 (N_12191,N_7141,N_6672);
nand U12192 (N_12192,N_5427,N_9114);
nand U12193 (N_12193,N_8681,N_7713);
nor U12194 (N_12194,N_6965,N_7093);
nand U12195 (N_12195,N_5083,N_6250);
nand U12196 (N_12196,N_9862,N_7926);
nand U12197 (N_12197,N_6415,N_8845);
and U12198 (N_12198,N_8717,N_6766);
or U12199 (N_12199,N_9092,N_8042);
xor U12200 (N_12200,N_8366,N_8098);
or U12201 (N_12201,N_8559,N_5015);
xnor U12202 (N_12202,N_9070,N_5830);
or U12203 (N_12203,N_7172,N_7077);
or U12204 (N_12204,N_6285,N_6664);
nor U12205 (N_12205,N_7997,N_9355);
nor U12206 (N_12206,N_8581,N_7834);
xnor U12207 (N_12207,N_9876,N_9888);
and U12208 (N_12208,N_7667,N_9842);
or U12209 (N_12209,N_7650,N_7600);
xnor U12210 (N_12210,N_9346,N_9677);
nand U12211 (N_12211,N_6952,N_6039);
xor U12212 (N_12212,N_5176,N_9782);
nand U12213 (N_12213,N_6595,N_5618);
nor U12214 (N_12214,N_5749,N_6219);
and U12215 (N_12215,N_9577,N_5666);
and U12216 (N_12216,N_9525,N_8212);
or U12217 (N_12217,N_6081,N_9127);
and U12218 (N_12218,N_8785,N_7897);
nand U12219 (N_12219,N_9415,N_5794);
nor U12220 (N_12220,N_6655,N_6125);
nor U12221 (N_12221,N_8347,N_7968);
nor U12222 (N_12222,N_5311,N_6108);
or U12223 (N_12223,N_8962,N_7390);
xor U12224 (N_12224,N_7075,N_7810);
nor U12225 (N_12225,N_5267,N_7895);
nor U12226 (N_12226,N_7368,N_9033);
nand U12227 (N_12227,N_5689,N_9779);
nand U12228 (N_12228,N_9761,N_5135);
nand U12229 (N_12229,N_7833,N_6790);
nor U12230 (N_12230,N_8180,N_6154);
nor U12231 (N_12231,N_5210,N_6968);
nand U12232 (N_12232,N_5175,N_6371);
nand U12233 (N_12233,N_8814,N_7578);
or U12234 (N_12234,N_5771,N_7580);
and U12235 (N_12235,N_9110,N_5140);
and U12236 (N_12236,N_7289,N_5343);
or U12237 (N_12237,N_5356,N_6317);
nand U12238 (N_12238,N_5539,N_5728);
xor U12239 (N_12239,N_5181,N_6387);
and U12240 (N_12240,N_7287,N_9435);
or U12241 (N_12241,N_9240,N_8238);
and U12242 (N_12242,N_9495,N_6954);
xnor U12243 (N_12243,N_6337,N_6100);
nor U12244 (N_12244,N_5941,N_5860);
or U12245 (N_12245,N_6267,N_9463);
nor U12246 (N_12246,N_9024,N_5186);
nor U12247 (N_12247,N_7553,N_5891);
or U12248 (N_12248,N_6597,N_5121);
nor U12249 (N_12249,N_6149,N_5318);
and U12250 (N_12250,N_8418,N_9442);
xnor U12251 (N_12251,N_9825,N_9735);
nor U12252 (N_12252,N_6503,N_5524);
or U12253 (N_12253,N_7636,N_6237);
and U12254 (N_12254,N_9662,N_5452);
or U12255 (N_12255,N_5358,N_6481);
xor U12256 (N_12256,N_5491,N_8911);
nor U12257 (N_12257,N_9555,N_9949);
nor U12258 (N_12258,N_9075,N_9957);
or U12259 (N_12259,N_8908,N_6912);
nor U12260 (N_12260,N_6883,N_6567);
and U12261 (N_12261,N_9966,N_6927);
xor U12262 (N_12262,N_7669,N_5551);
xnor U12263 (N_12263,N_6414,N_7818);
xnor U12264 (N_12264,N_9932,N_8467);
or U12265 (N_12265,N_8136,N_9576);
nor U12266 (N_12266,N_8120,N_5718);
nand U12267 (N_12267,N_6833,N_6679);
and U12268 (N_12268,N_8773,N_5002);
xnor U12269 (N_12269,N_5993,N_7491);
nor U12270 (N_12270,N_9095,N_9472);
or U12271 (N_12271,N_9593,N_7570);
nor U12272 (N_12272,N_7241,N_5756);
xor U12273 (N_12273,N_7481,N_8312);
or U12274 (N_12274,N_5162,N_5067);
nand U12275 (N_12275,N_7231,N_8899);
xor U12276 (N_12276,N_6449,N_5280);
xor U12277 (N_12277,N_5350,N_7887);
xor U12278 (N_12278,N_5282,N_6067);
nor U12279 (N_12279,N_5944,N_9816);
nor U12280 (N_12280,N_9943,N_9515);
and U12281 (N_12281,N_5823,N_5185);
and U12282 (N_12282,N_6169,N_5381);
xor U12283 (N_12283,N_5443,N_9373);
and U12284 (N_12284,N_5490,N_6016);
and U12285 (N_12285,N_9413,N_5789);
and U12286 (N_12286,N_9961,N_9594);
xor U12287 (N_12287,N_7569,N_6184);
nand U12288 (N_12288,N_5964,N_9091);
nor U12289 (N_12289,N_9891,N_8889);
xor U12290 (N_12290,N_5513,N_9176);
nor U12291 (N_12291,N_6278,N_5735);
or U12292 (N_12292,N_7757,N_6519);
or U12293 (N_12293,N_6765,N_9335);
xor U12294 (N_12294,N_6676,N_9259);
nand U12295 (N_12295,N_9834,N_9138);
xor U12296 (N_12296,N_6832,N_9548);
nor U12297 (N_12297,N_6096,N_8891);
xnor U12298 (N_12298,N_9965,N_6024);
xor U12299 (N_12299,N_9241,N_5298);
xor U12300 (N_12300,N_5686,N_5591);
xor U12301 (N_12301,N_6297,N_5151);
or U12302 (N_12302,N_6453,N_9667);
and U12303 (N_12303,N_6000,N_6290);
nor U12304 (N_12304,N_6879,N_7380);
nand U12305 (N_12305,N_9043,N_6217);
nor U12306 (N_12306,N_8587,N_8204);
nor U12307 (N_12307,N_7700,N_5774);
nand U12308 (N_12308,N_7777,N_7984);
xnor U12309 (N_12309,N_6885,N_5494);
and U12310 (N_12310,N_6225,N_7783);
nand U12311 (N_12311,N_8256,N_8722);
or U12312 (N_12312,N_6312,N_8374);
and U12313 (N_12313,N_7512,N_9719);
nor U12314 (N_12314,N_7154,N_5899);
nor U12315 (N_12315,N_6710,N_6388);
xor U12316 (N_12316,N_8346,N_6588);
or U12317 (N_12317,N_8147,N_8714);
or U12318 (N_12318,N_9004,N_8572);
or U12319 (N_12319,N_8739,N_6645);
nand U12320 (N_12320,N_5138,N_6896);
and U12321 (N_12321,N_8932,N_8688);
xnor U12322 (N_12322,N_5515,N_9717);
xnor U12323 (N_12323,N_5608,N_6811);
xnor U12324 (N_12324,N_6161,N_9363);
or U12325 (N_12325,N_6055,N_8752);
and U12326 (N_12326,N_9204,N_7617);
or U12327 (N_12327,N_7180,N_9985);
nand U12328 (N_12328,N_6658,N_6163);
nor U12329 (N_12329,N_5168,N_8004);
nor U12330 (N_12330,N_8055,N_6352);
and U12331 (N_12331,N_9198,N_5218);
nand U12332 (N_12332,N_7981,N_9649);
xor U12333 (N_12333,N_8999,N_8327);
and U12334 (N_12334,N_5266,N_5156);
or U12335 (N_12335,N_5980,N_5668);
and U12336 (N_12336,N_5335,N_7192);
nand U12337 (N_12337,N_9871,N_7973);
xnor U12338 (N_12338,N_6787,N_7480);
nor U12339 (N_12339,N_5315,N_6559);
nand U12340 (N_12340,N_6105,N_5387);
and U12341 (N_12341,N_9426,N_8602);
nor U12342 (N_12342,N_9217,N_5203);
xnor U12343 (N_12343,N_7670,N_7554);
or U12344 (N_12344,N_6221,N_7021);
or U12345 (N_12345,N_6699,N_6454);
nor U12346 (N_12346,N_8535,N_5850);
and U12347 (N_12347,N_8407,N_8762);
or U12348 (N_12348,N_5653,N_9035);
or U12349 (N_12349,N_9982,N_9225);
and U12350 (N_12350,N_7299,N_9360);
or U12351 (N_12351,N_6510,N_9219);
nand U12352 (N_12352,N_9503,N_5331);
xnor U12353 (N_12353,N_7941,N_7404);
and U12354 (N_12354,N_8976,N_8025);
xnor U12355 (N_12355,N_9253,N_9166);
xor U12356 (N_12356,N_6688,N_5231);
nand U12357 (N_12357,N_8656,N_8539);
and U12358 (N_12358,N_7002,N_7956);
and U12359 (N_12359,N_7189,N_7164);
nand U12360 (N_12360,N_5105,N_6028);
or U12361 (N_12361,N_8468,N_6924);
nor U12362 (N_12362,N_5927,N_9136);
nand U12363 (N_12363,N_8126,N_9064);
nand U12364 (N_12364,N_9789,N_9856);
xnor U12365 (N_12365,N_9952,N_7217);
xor U12366 (N_12366,N_8135,N_8383);
xor U12367 (N_12367,N_9658,N_5967);
nor U12368 (N_12368,N_7042,N_8519);
nor U12369 (N_12369,N_9868,N_8509);
and U12370 (N_12370,N_9774,N_6091);
nand U12371 (N_12371,N_7449,N_5035);
nand U12372 (N_12372,N_8543,N_8612);
or U12373 (N_12373,N_7896,N_8229);
and U12374 (N_12374,N_6295,N_5849);
nor U12375 (N_12375,N_7157,N_9619);
nor U12376 (N_12376,N_5779,N_9350);
or U12377 (N_12377,N_9829,N_9559);
or U12378 (N_12378,N_8116,N_6786);
xnor U12379 (N_12379,N_5492,N_6998);
and U12380 (N_12380,N_9238,N_5386);
nand U12381 (N_12381,N_5488,N_7589);
xor U12382 (N_12382,N_7642,N_5420);
nor U12383 (N_12383,N_6226,N_7294);
nand U12384 (N_12384,N_9157,N_5498);
or U12385 (N_12385,N_6836,N_8923);
nor U12386 (N_12386,N_7487,N_5184);
and U12387 (N_12387,N_7324,N_7836);
nand U12388 (N_12388,N_8035,N_5695);
and U12389 (N_12389,N_9230,N_8542);
and U12390 (N_12390,N_7811,N_7989);
nand U12391 (N_12391,N_6966,N_5416);
nand U12392 (N_12392,N_8030,N_5840);
or U12393 (N_12393,N_9617,N_8709);
or U12394 (N_12394,N_7092,N_9954);
xnor U12395 (N_12395,N_7924,N_8935);
nor U12396 (N_12396,N_9446,N_7067);
xor U12397 (N_12397,N_7233,N_7265);
or U12398 (N_12398,N_5139,N_7152);
and U12399 (N_12399,N_9100,N_5721);
and U12400 (N_12400,N_8274,N_9263);
nor U12401 (N_12401,N_6486,N_8461);
nand U12402 (N_12402,N_6755,N_6062);
xor U12403 (N_12403,N_7104,N_6358);
or U12404 (N_12404,N_9121,N_9889);
and U12405 (N_12405,N_9257,N_6985);
or U12406 (N_12406,N_5521,N_6709);
or U12407 (N_12407,N_7359,N_7835);
nor U12408 (N_12408,N_7248,N_9073);
xor U12409 (N_12409,N_9287,N_8152);
nand U12410 (N_12410,N_7632,N_8525);
nor U12411 (N_12411,N_9794,N_8090);
and U12412 (N_12412,N_8463,N_6522);
nor U12413 (N_12413,N_8169,N_9894);
nand U12414 (N_12414,N_9592,N_5237);
xnor U12415 (N_12415,N_6343,N_8092);
nor U12416 (N_12416,N_7088,N_9260);
and U12417 (N_12417,N_8770,N_7460);
nand U12418 (N_12418,N_9648,N_5022);
and U12419 (N_12419,N_7455,N_7878);
and U12420 (N_12420,N_7128,N_9000);
xor U12421 (N_12421,N_6310,N_8410);
nor U12422 (N_12422,N_6029,N_8625);
xnor U12423 (N_12423,N_6115,N_9277);
xor U12424 (N_12424,N_8522,N_7987);
xor U12425 (N_12425,N_5795,N_7086);
and U12426 (N_12426,N_7861,N_5921);
xor U12427 (N_12427,N_7338,N_6167);
nand U12428 (N_12428,N_9670,N_8811);
or U12429 (N_12429,N_7692,N_6933);
or U12430 (N_12430,N_5888,N_5580);
nor U12431 (N_12431,N_9421,N_6539);
and U12432 (N_12432,N_5004,N_8475);
and U12433 (N_12433,N_7702,N_5880);
or U12434 (N_12434,N_5277,N_5309);
xor U12435 (N_12435,N_6193,N_9600);
or U12436 (N_12436,N_9519,N_9861);
and U12437 (N_12437,N_5232,N_7829);
or U12438 (N_12438,N_5816,N_7257);
xnor U12439 (N_12439,N_8961,N_5047);
and U12440 (N_12440,N_8991,N_6185);
nor U12441 (N_12441,N_5775,N_6027);
and U12442 (N_12442,N_6662,N_8331);
and U12443 (N_12443,N_8834,N_6893);
nand U12444 (N_12444,N_6497,N_5407);
nor U12445 (N_12445,N_8031,N_5341);
nand U12446 (N_12446,N_5554,N_9203);
xnor U12447 (N_12447,N_6878,N_7595);
nor U12448 (N_12448,N_9486,N_6253);
or U12449 (N_12449,N_5763,N_7409);
xor U12450 (N_12450,N_8051,N_8649);
nand U12451 (N_12451,N_5371,N_9431);
or U12452 (N_12452,N_8831,N_9275);
xor U12453 (N_12453,N_5975,N_5879);
nor U12454 (N_12454,N_5726,N_5153);
nor U12455 (N_12455,N_9615,N_7208);
or U12456 (N_12456,N_5943,N_9900);
nor U12457 (N_12457,N_5522,N_8225);
xnor U12458 (N_12458,N_6520,N_5540);
nand U12459 (N_12459,N_5082,N_6088);
or U12460 (N_12460,N_5722,N_8784);
and U12461 (N_12461,N_6377,N_6478);
nand U12462 (N_12462,N_5412,N_6013);
or U12463 (N_12463,N_7262,N_5679);
and U12464 (N_12464,N_7137,N_6407);
xnor U12465 (N_12465,N_6997,N_7437);
and U12466 (N_12466,N_6758,N_7421);
or U12467 (N_12467,N_5946,N_8440);
xnor U12468 (N_12468,N_8711,N_7641);
nor U12469 (N_12469,N_7237,N_7738);
nand U12470 (N_12470,N_6858,N_9634);
xnor U12471 (N_12471,N_7635,N_8384);
xor U12472 (N_12472,N_8361,N_8655);
xor U12473 (N_12473,N_9537,N_5813);
xor U12474 (N_12474,N_8106,N_5617);
xor U12475 (N_12475,N_6023,N_7378);
and U12476 (N_12476,N_9758,N_8973);
and U12477 (N_12477,N_7147,N_7348);
nor U12478 (N_12478,N_8404,N_8054);
and U12479 (N_12479,N_5057,N_6880);
nand U12480 (N_12480,N_7546,N_8222);
and U12481 (N_12481,N_6446,N_5649);
and U12482 (N_12482,N_9483,N_6719);
or U12483 (N_12483,N_9984,N_9695);
and U12484 (N_12484,N_8835,N_8252);
xor U12485 (N_12485,N_9755,N_9094);
nor U12486 (N_12486,N_5820,N_5517);
or U12487 (N_12487,N_6477,N_7756);
and U12488 (N_12488,N_9614,N_5401);
nand U12489 (N_12489,N_6475,N_5213);
and U12490 (N_12490,N_7195,N_7832);
xor U12491 (N_12491,N_8181,N_6930);
nor U12492 (N_12492,N_7817,N_6706);
nor U12493 (N_12493,N_9694,N_7191);
nand U12494 (N_12494,N_8171,N_6648);
nor U12495 (N_12495,N_7899,N_8541);
xor U12496 (N_12496,N_7488,N_7909);
xnor U12497 (N_12497,N_9484,N_9921);
nor U12498 (N_12498,N_8053,N_9172);
nor U12499 (N_12499,N_9269,N_7681);
xor U12500 (N_12500,N_8782,N_9108);
xor U12501 (N_12501,N_5045,N_9004);
xnor U12502 (N_12502,N_6078,N_8046);
xor U12503 (N_12503,N_9717,N_6183);
and U12504 (N_12504,N_8331,N_7936);
nand U12505 (N_12505,N_6797,N_8135);
or U12506 (N_12506,N_7035,N_5983);
or U12507 (N_12507,N_6330,N_8472);
and U12508 (N_12508,N_5930,N_6006);
and U12509 (N_12509,N_8104,N_6542);
xor U12510 (N_12510,N_7981,N_5712);
and U12511 (N_12511,N_6501,N_6259);
or U12512 (N_12512,N_5026,N_9855);
xnor U12513 (N_12513,N_6869,N_5918);
nand U12514 (N_12514,N_6561,N_7623);
nand U12515 (N_12515,N_7872,N_6783);
nand U12516 (N_12516,N_6842,N_9745);
xor U12517 (N_12517,N_8508,N_8702);
and U12518 (N_12518,N_5930,N_5624);
nand U12519 (N_12519,N_7098,N_5259);
or U12520 (N_12520,N_8519,N_9095);
xor U12521 (N_12521,N_8767,N_7577);
and U12522 (N_12522,N_9854,N_7334);
nor U12523 (N_12523,N_8036,N_5833);
nor U12524 (N_12524,N_8740,N_5822);
or U12525 (N_12525,N_5820,N_6652);
nand U12526 (N_12526,N_7668,N_6058);
nand U12527 (N_12527,N_5629,N_9713);
xnor U12528 (N_12528,N_6314,N_7926);
or U12529 (N_12529,N_5451,N_8000);
and U12530 (N_12530,N_7046,N_5812);
xor U12531 (N_12531,N_6434,N_8730);
or U12532 (N_12532,N_8123,N_8005);
or U12533 (N_12533,N_5180,N_5815);
and U12534 (N_12534,N_5331,N_5686);
and U12535 (N_12535,N_6187,N_5919);
and U12536 (N_12536,N_9790,N_5487);
nor U12537 (N_12537,N_5629,N_8118);
and U12538 (N_12538,N_5078,N_5893);
xnor U12539 (N_12539,N_6326,N_6789);
or U12540 (N_12540,N_5308,N_7334);
nand U12541 (N_12541,N_8987,N_6120);
and U12542 (N_12542,N_5259,N_6463);
or U12543 (N_12543,N_9929,N_9053);
and U12544 (N_12544,N_7215,N_6806);
xnor U12545 (N_12545,N_7213,N_9251);
or U12546 (N_12546,N_7334,N_6978);
nand U12547 (N_12547,N_5657,N_5784);
nor U12548 (N_12548,N_7984,N_6162);
and U12549 (N_12549,N_8995,N_8966);
and U12550 (N_12550,N_7206,N_9125);
nor U12551 (N_12551,N_5718,N_6560);
and U12552 (N_12552,N_9805,N_7049);
xor U12553 (N_12553,N_9084,N_7499);
or U12554 (N_12554,N_8204,N_5549);
nand U12555 (N_12555,N_5003,N_8259);
nand U12556 (N_12556,N_8415,N_8246);
or U12557 (N_12557,N_9863,N_8313);
nor U12558 (N_12558,N_8653,N_6821);
nand U12559 (N_12559,N_5125,N_6981);
nand U12560 (N_12560,N_9322,N_5158);
or U12561 (N_12561,N_7061,N_9362);
nand U12562 (N_12562,N_9949,N_8249);
xor U12563 (N_12563,N_9231,N_9001);
and U12564 (N_12564,N_7116,N_8394);
or U12565 (N_12565,N_8232,N_6841);
xor U12566 (N_12566,N_7425,N_7523);
and U12567 (N_12567,N_6768,N_5825);
or U12568 (N_12568,N_5468,N_7336);
or U12569 (N_12569,N_6504,N_9336);
and U12570 (N_12570,N_8889,N_8230);
xor U12571 (N_12571,N_9712,N_9096);
nor U12572 (N_12572,N_8699,N_7875);
and U12573 (N_12573,N_7227,N_7946);
or U12574 (N_12574,N_9833,N_6737);
and U12575 (N_12575,N_7150,N_7773);
xnor U12576 (N_12576,N_5333,N_5709);
nand U12577 (N_12577,N_5615,N_8583);
xnor U12578 (N_12578,N_9372,N_5573);
nand U12579 (N_12579,N_7193,N_8414);
nand U12580 (N_12580,N_9779,N_7225);
nand U12581 (N_12581,N_5329,N_7895);
or U12582 (N_12582,N_8088,N_8602);
nor U12583 (N_12583,N_7654,N_8315);
and U12584 (N_12584,N_6308,N_5211);
and U12585 (N_12585,N_8475,N_8307);
xnor U12586 (N_12586,N_8678,N_9331);
or U12587 (N_12587,N_6783,N_9785);
nor U12588 (N_12588,N_8008,N_7401);
nor U12589 (N_12589,N_5201,N_8196);
nor U12590 (N_12590,N_8564,N_6711);
or U12591 (N_12591,N_7421,N_9761);
xnor U12592 (N_12592,N_9828,N_8037);
and U12593 (N_12593,N_9938,N_7623);
nor U12594 (N_12594,N_6918,N_7240);
nand U12595 (N_12595,N_7610,N_7050);
nand U12596 (N_12596,N_8158,N_5734);
and U12597 (N_12597,N_8946,N_6091);
nor U12598 (N_12598,N_8825,N_8593);
and U12599 (N_12599,N_8067,N_9292);
or U12600 (N_12600,N_9380,N_6842);
nand U12601 (N_12601,N_8110,N_6754);
nand U12602 (N_12602,N_5151,N_9077);
and U12603 (N_12603,N_5515,N_5536);
nand U12604 (N_12604,N_5775,N_6687);
xnor U12605 (N_12605,N_5609,N_8164);
xor U12606 (N_12606,N_7580,N_7441);
nand U12607 (N_12607,N_7644,N_5854);
and U12608 (N_12608,N_6260,N_9056);
nor U12609 (N_12609,N_6403,N_8096);
and U12610 (N_12610,N_8587,N_9435);
or U12611 (N_12611,N_8532,N_9210);
nand U12612 (N_12612,N_5551,N_8278);
nand U12613 (N_12613,N_9563,N_8149);
and U12614 (N_12614,N_8492,N_9128);
and U12615 (N_12615,N_6496,N_9735);
and U12616 (N_12616,N_7826,N_8171);
and U12617 (N_12617,N_6000,N_8744);
nand U12618 (N_12618,N_9937,N_5028);
and U12619 (N_12619,N_6260,N_9727);
and U12620 (N_12620,N_6490,N_7693);
and U12621 (N_12621,N_5206,N_7421);
nor U12622 (N_12622,N_6154,N_8990);
nand U12623 (N_12623,N_8827,N_9494);
and U12624 (N_12624,N_6557,N_6895);
and U12625 (N_12625,N_5560,N_8932);
and U12626 (N_12626,N_5878,N_5677);
and U12627 (N_12627,N_8427,N_9640);
and U12628 (N_12628,N_7181,N_7499);
or U12629 (N_12629,N_6747,N_9681);
xnor U12630 (N_12630,N_8295,N_6312);
and U12631 (N_12631,N_5448,N_5874);
or U12632 (N_12632,N_5185,N_9898);
nor U12633 (N_12633,N_9677,N_9574);
and U12634 (N_12634,N_9092,N_8064);
nor U12635 (N_12635,N_7371,N_6136);
xor U12636 (N_12636,N_8560,N_5237);
and U12637 (N_12637,N_6674,N_9082);
nand U12638 (N_12638,N_8895,N_8595);
nand U12639 (N_12639,N_6238,N_5174);
xnor U12640 (N_12640,N_8922,N_9260);
nor U12641 (N_12641,N_7805,N_7186);
nor U12642 (N_12642,N_8459,N_9707);
nor U12643 (N_12643,N_6343,N_8963);
nand U12644 (N_12644,N_9973,N_9837);
nor U12645 (N_12645,N_8170,N_7368);
nor U12646 (N_12646,N_7022,N_7249);
and U12647 (N_12647,N_9725,N_8228);
and U12648 (N_12648,N_5950,N_8865);
nor U12649 (N_12649,N_7908,N_8375);
and U12650 (N_12650,N_7708,N_6762);
and U12651 (N_12651,N_7569,N_8731);
nand U12652 (N_12652,N_8268,N_7573);
xor U12653 (N_12653,N_9422,N_5796);
and U12654 (N_12654,N_8955,N_6701);
or U12655 (N_12655,N_8327,N_8859);
xnor U12656 (N_12656,N_5606,N_9315);
nor U12657 (N_12657,N_5192,N_7229);
nand U12658 (N_12658,N_7899,N_7773);
xor U12659 (N_12659,N_6692,N_9423);
nor U12660 (N_12660,N_9603,N_7349);
and U12661 (N_12661,N_5589,N_6488);
or U12662 (N_12662,N_5887,N_7027);
nor U12663 (N_12663,N_6415,N_9835);
nand U12664 (N_12664,N_5870,N_6179);
nand U12665 (N_12665,N_9704,N_7706);
and U12666 (N_12666,N_9061,N_8741);
or U12667 (N_12667,N_7412,N_8552);
or U12668 (N_12668,N_5727,N_7176);
or U12669 (N_12669,N_5333,N_5460);
nor U12670 (N_12670,N_5543,N_8083);
or U12671 (N_12671,N_6990,N_6930);
nor U12672 (N_12672,N_7328,N_9306);
nand U12673 (N_12673,N_6149,N_9689);
xor U12674 (N_12674,N_8475,N_5857);
and U12675 (N_12675,N_6927,N_7312);
nand U12676 (N_12676,N_5882,N_8113);
nor U12677 (N_12677,N_9984,N_6006);
and U12678 (N_12678,N_5575,N_6056);
or U12679 (N_12679,N_6281,N_7616);
nand U12680 (N_12680,N_6788,N_6487);
nor U12681 (N_12681,N_6675,N_9958);
or U12682 (N_12682,N_7061,N_7136);
nor U12683 (N_12683,N_9187,N_5735);
xnor U12684 (N_12684,N_7483,N_8589);
nor U12685 (N_12685,N_7777,N_7497);
nor U12686 (N_12686,N_9116,N_7268);
nand U12687 (N_12687,N_9105,N_9172);
or U12688 (N_12688,N_6273,N_9548);
xor U12689 (N_12689,N_8073,N_5447);
and U12690 (N_12690,N_8818,N_5358);
nor U12691 (N_12691,N_7142,N_9998);
nand U12692 (N_12692,N_7762,N_8410);
nor U12693 (N_12693,N_9355,N_9694);
and U12694 (N_12694,N_6160,N_5106);
nor U12695 (N_12695,N_6754,N_8246);
and U12696 (N_12696,N_6741,N_7189);
xor U12697 (N_12697,N_9304,N_8283);
xnor U12698 (N_12698,N_9615,N_6295);
and U12699 (N_12699,N_6761,N_9977);
nor U12700 (N_12700,N_7849,N_7524);
xor U12701 (N_12701,N_8667,N_5963);
xnor U12702 (N_12702,N_5793,N_6702);
nor U12703 (N_12703,N_9783,N_6877);
or U12704 (N_12704,N_8508,N_8235);
nand U12705 (N_12705,N_6921,N_9483);
or U12706 (N_12706,N_7965,N_5696);
xnor U12707 (N_12707,N_6879,N_5348);
or U12708 (N_12708,N_7147,N_5927);
or U12709 (N_12709,N_8692,N_9864);
nand U12710 (N_12710,N_6393,N_5264);
nand U12711 (N_12711,N_6170,N_8777);
and U12712 (N_12712,N_8843,N_6848);
nor U12713 (N_12713,N_7035,N_8971);
nand U12714 (N_12714,N_5737,N_9139);
nor U12715 (N_12715,N_9023,N_7136);
and U12716 (N_12716,N_5574,N_9152);
nand U12717 (N_12717,N_6619,N_8740);
or U12718 (N_12718,N_7038,N_9345);
and U12719 (N_12719,N_7038,N_7908);
nand U12720 (N_12720,N_7824,N_9403);
nor U12721 (N_12721,N_5464,N_6228);
and U12722 (N_12722,N_5354,N_6200);
or U12723 (N_12723,N_6140,N_8203);
nor U12724 (N_12724,N_9032,N_6828);
or U12725 (N_12725,N_7533,N_7769);
or U12726 (N_12726,N_6706,N_6564);
or U12727 (N_12727,N_8255,N_9922);
xnor U12728 (N_12728,N_9089,N_7602);
xnor U12729 (N_12729,N_8003,N_9746);
nand U12730 (N_12730,N_9122,N_8073);
or U12731 (N_12731,N_5493,N_9629);
nor U12732 (N_12732,N_5695,N_8446);
or U12733 (N_12733,N_6847,N_9470);
nor U12734 (N_12734,N_9702,N_6181);
or U12735 (N_12735,N_5606,N_5209);
nor U12736 (N_12736,N_8067,N_5744);
and U12737 (N_12737,N_5561,N_5076);
and U12738 (N_12738,N_8131,N_9220);
nand U12739 (N_12739,N_7182,N_8040);
nor U12740 (N_12740,N_5162,N_7686);
or U12741 (N_12741,N_6083,N_8154);
or U12742 (N_12742,N_9491,N_9320);
nor U12743 (N_12743,N_8554,N_7076);
xor U12744 (N_12744,N_7418,N_6354);
nand U12745 (N_12745,N_5094,N_5986);
nand U12746 (N_12746,N_7697,N_8251);
and U12747 (N_12747,N_8099,N_9437);
nor U12748 (N_12748,N_7590,N_6298);
xor U12749 (N_12749,N_9097,N_7401);
nor U12750 (N_12750,N_5830,N_5689);
and U12751 (N_12751,N_8072,N_9715);
nor U12752 (N_12752,N_5315,N_5388);
or U12753 (N_12753,N_9982,N_9097);
nor U12754 (N_12754,N_9232,N_9020);
or U12755 (N_12755,N_9956,N_9062);
nand U12756 (N_12756,N_9092,N_7570);
xnor U12757 (N_12757,N_6141,N_9407);
and U12758 (N_12758,N_8863,N_9401);
xnor U12759 (N_12759,N_8542,N_8200);
nand U12760 (N_12760,N_5888,N_8277);
nand U12761 (N_12761,N_7938,N_7806);
nand U12762 (N_12762,N_7598,N_9324);
nor U12763 (N_12763,N_8084,N_7965);
nor U12764 (N_12764,N_8546,N_6880);
xor U12765 (N_12765,N_6187,N_8902);
nor U12766 (N_12766,N_7486,N_6680);
nor U12767 (N_12767,N_5989,N_6224);
xnor U12768 (N_12768,N_7388,N_9956);
xnor U12769 (N_12769,N_7906,N_8157);
nor U12770 (N_12770,N_9818,N_6704);
nor U12771 (N_12771,N_8379,N_7416);
nand U12772 (N_12772,N_5537,N_9660);
nand U12773 (N_12773,N_6062,N_9402);
nor U12774 (N_12774,N_5613,N_5685);
and U12775 (N_12775,N_6789,N_5250);
nand U12776 (N_12776,N_6443,N_5669);
xor U12777 (N_12777,N_5999,N_9802);
nand U12778 (N_12778,N_7459,N_6440);
xnor U12779 (N_12779,N_6531,N_8079);
and U12780 (N_12780,N_7271,N_5391);
and U12781 (N_12781,N_8617,N_5820);
nor U12782 (N_12782,N_5374,N_7083);
and U12783 (N_12783,N_5290,N_9973);
nor U12784 (N_12784,N_7514,N_9065);
nand U12785 (N_12785,N_5756,N_8971);
and U12786 (N_12786,N_6011,N_5056);
nand U12787 (N_12787,N_8234,N_8105);
or U12788 (N_12788,N_6114,N_8970);
and U12789 (N_12789,N_7239,N_5711);
and U12790 (N_12790,N_5740,N_8325);
and U12791 (N_12791,N_5146,N_8747);
or U12792 (N_12792,N_5106,N_6008);
xnor U12793 (N_12793,N_9997,N_9627);
or U12794 (N_12794,N_9246,N_7562);
xor U12795 (N_12795,N_8108,N_8204);
xnor U12796 (N_12796,N_7964,N_7497);
xnor U12797 (N_12797,N_7907,N_8063);
and U12798 (N_12798,N_5836,N_6671);
nand U12799 (N_12799,N_6645,N_9500);
and U12800 (N_12800,N_9699,N_5973);
and U12801 (N_12801,N_8209,N_7311);
xnor U12802 (N_12802,N_6320,N_5376);
nor U12803 (N_12803,N_6431,N_6850);
nor U12804 (N_12804,N_9629,N_8462);
and U12805 (N_12805,N_8507,N_8347);
or U12806 (N_12806,N_5867,N_7198);
xor U12807 (N_12807,N_9920,N_6469);
and U12808 (N_12808,N_7193,N_9326);
xor U12809 (N_12809,N_6995,N_8791);
xnor U12810 (N_12810,N_5175,N_5097);
or U12811 (N_12811,N_5864,N_8851);
nor U12812 (N_12812,N_6514,N_7988);
xnor U12813 (N_12813,N_5167,N_5380);
xnor U12814 (N_12814,N_5665,N_5325);
and U12815 (N_12815,N_8515,N_7907);
or U12816 (N_12816,N_6563,N_7322);
nor U12817 (N_12817,N_6497,N_5458);
xnor U12818 (N_12818,N_7771,N_6596);
nand U12819 (N_12819,N_8050,N_7802);
and U12820 (N_12820,N_9029,N_5557);
nand U12821 (N_12821,N_5775,N_9814);
and U12822 (N_12822,N_5274,N_9993);
nand U12823 (N_12823,N_9576,N_8544);
xnor U12824 (N_12824,N_6891,N_7210);
and U12825 (N_12825,N_7112,N_9763);
and U12826 (N_12826,N_6853,N_9692);
xor U12827 (N_12827,N_9909,N_6975);
xor U12828 (N_12828,N_7510,N_6352);
xor U12829 (N_12829,N_5746,N_7729);
nor U12830 (N_12830,N_8837,N_9509);
nor U12831 (N_12831,N_8759,N_6132);
or U12832 (N_12832,N_5566,N_5138);
nor U12833 (N_12833,N_6505,N_5516);
nand U12834 (N_12834,N_5821,N_8705);
and U12835 (N_12835,N_9382,N_5857);
or U12836 (N_12836,N_8953,N_9712);
nor U12837 (N_12837,N_5248,N_9269);
or U12838 (N_12838,N_8329,N_8807);
and U12839 (N_12839,N_9485,N_9621);
and U12840 (N_12840,N_8111,N_6595);
or U12841 (N_12841,N_6903,N_6568);
and U12842 (N_12842,N_5413,N_9801);
and U12843 (N_12843,N_8349,N_5926);
or U12844 (N_12844,N_9140,N_8168);
or U12845 (N_12845,N_9293,N_6361);
or U12846 (N_12846,N_8629,N_8469);
and U12847 (N_12847,N_6776,N_5886);
nand U12848 (N_12848,N_9826,N_5180);
nand U12849 (N_12849,N_5209,N_6364);
xor U12850 (N_12850,N_8864,N_9564);
or U12851 (N_12851,N_6822,N_7512);
nor U12852 (N_12852,N_5308,N_6063);
nand U12853 (N_12853,N_5074,N_8192);
xnor U12854 (N_12854,N_7153,N_9087);
xnor U12855 (N_12855,N_6541,N_5891);
xnor U12856 (N_12856,N_7026,N_9643);
xor U12857 (N_12857,N_6845,N_7606);
nand U12858 (N_12858,N_5524,N_7396);
nand U12859 (N_12859,N_8372,N_7267);
and U12860 (N_12860,N_5531,N_9115);
nor U12861 (N_12861,N_8996,N_9770);
xor U12862 (N_12862,N_8314,N_5697);
xor U12863 (N_12863,N_7861,N_8901);
or U12864 (N_12864,N_9919,N_6368);
and U12865 (N_12865,N_6175,N_7607);
xor U12866 (N_12866,N_7430,N_9483);
nand U12867 (N_12867,N_8837,N_6836);
nor U12868 (N_12868,N_8305,N_7458);
nor U12869 (N_12869,N_8276,N_9398);
nand U12870 (N_12870,N_9759,N_7095);
and U12871 (N_12871,N_5990,N_5610);
nor U12872 (N_12872,N_7824,N_7775);
nor U12873 (N_12873,N_7132,N_5595);
xnor U12874 (N_12874,N_7705,N_6440);
xor U12875 (N_12875,N_6200,N_5118);
and U12876 (N_12876,N_7719,N_8556);
or U12877 (N_12877,N_5301,N_6478);
or U12878 (N_12878,N_6631,N_9851);
nor U12879 (N_12879,N_5147,N_6356);
nand U12880 (N_12880,N_6010,N_8124);
xnor U12881 (N_12881,N_9194,N_6015);
and U12882 (N_12882,N_5812,N_6351);
and U12883 (N_12883,N_5529,N_6883);
nor U12884 (N_12884,N_5229,N_9549);
or U12885 (N_12885,N_7382,N_8752);
and U12886 (N_12886,N_7062,N_6586);
nor U12887 (N_12887,N_7721,N_5101);
nor U12888 (N_12888,N_7510,N_5973);
and U12889 (N_12889,N_7545,N_6273);
nand U12890 (N_12890,N_6959,N_8928);
nand U12891 (N_12891,N_6881,N_5063);
or U12892 (N_12892,N_7062,N_7732);
nor U12893 (N_12893,N_9885,N_9335);
xor U12894 (N_12894,N_6895,N_5819);
or U12895 (N_12895,N_8823,N_7008);
xor U12896 (N_12896,N_5176,N_5737);
xor U12897 (N_12897,N_8204,N_6151);
or U12898 (N_12898,N_9092,N_6669);
xnor U12899 (N_12899,N_7037,N_7750);
or U12900 (N_12900,N_8182,N_5171);
or U12901 (N_12901,N_8195,N_5827);
xnor U12902 (N_12902,N_8328,N_9897);
or U12903 (N_12903,N_7318,N_7981);
xnor U12904 (N_12904,N_6920,N_9986);
and U12905 (N_12905,N_5608,N_7863);
nor U12906 (N_12906,N_5210,N_8499);
xnor U12907 (N_12907,N_9151,N_6881);
xnor U12908 (N_12908,N_8450,N_6497);
nand U12909 (N_12909,N_5161,N_6579);
xor U12910 (N_12910,N_5128,N_8657);
xor U12911 (N_12911,N_6784,N_9941);
or U12912 (N_12912,N_6862,N_5053);
nand U12913 (N_12913,N_8130,N_8565);
nand U12914 (N_12914,N_6878,N_5953);
nor U12915 (N_12915,N_8249,N_8682);
or U12916 (N_12916,N_7487,N_9113);
or U12917 (N_12917,N_9649,N_8922);
nor U12918 (N_12918,N_8227,N_9809);
or U12919 (N_12919,N_7692,N_5444);
nand U12920 (N_12920,N_7759,N_7841);
and U12921 (N_12921,N_5482,N_8560);
nand U12922 (N_12922,N_6403,N_7965);
or U12923 (N_12923,N_8358,N_6571);
nand U12924 (N_12924,N_5076,N_6689);
nor U12925 (N_12925,N_8342,N_5934);
and U12926 (N_12926,N_5726,N_9588);
and U12927 (N_12927,N_6089,N_6466);
nor U12928 (N_12928,N_6086,N_5089);
and U12929 (N_12929,N_9714,N_8756);
nor U12930 (N_12930,N_6638,N_5035);
xnor U12931 (N_12931,N_7065,N_5670);
or U12932 (N_12932,N_5555,N_5031);
nor U12933 (N_12933,N_5491,N_8819);
or U12934 (N_12934,N_9915,N_5712);
nor U12935 (N_12935,N_6422,N_5069);
xor U12936 (N_12936,N_5273,N_7375);
xor U12937 (N_12937,N_7198,N_9712);
or U12938 (N_12938,N_8232,N_7140);
xnor U12939 (N_12939,N_7759,N_6525);
nor U12940 (N_12940,N_8291,N_6201);
and U12941 (N_12941,N_8553,N_6698);
and U12942 (N_12942,N_7040,N_5751);
or U12943 (N_12943,N_5335,N_6019);
nor U12944 (N_12944,N_6683,N_5816);
xnor U12945 (N_12945,N_8740,N_8334);
nor U12946 (N_12946,N_9028,N_9090);
and U12947 (N_12947,N_5954,N_5243);
nand U12948 (N_12948,N_9990,N_6604);
or U12949 (N_12949,N_8542,N_6317);
or U12950 (N_12950,N_5911,N_8623);
nor U12951 (N_12951,N_9787,N_6141);
nor U12952 (N_12952,N_8591,N_7691);
and U12953 (N_12953,N_9569,N_7353);
or U12954 (N_12954,N_6412,N_6608);
xor U12955 (N_12955,N_6947,N_6369);
nor U12956 (N_12956,N_6607,N_8953);
xnor U12957 (N_12957,N_6372,N_7585);
and U12958 (N_12958,N_7970,N_8951);
and U12959 (N_12959,N_9911,N_6533);
xor U12960 (N_12960,N_5133,N_7411);
nand U12961 (N_12961,N_8717,N_9263);
and U12962 (N_12962,N_7072,N_7605);
xor U12963 (N_12963,N_5172,N_5313);
nor U12964 (N_12964,N_8503,N_7453);
xnor U12965 (N_12965,N_6498,N_8721);
or U12966 (N_12966,N_9262,N_6387);
or U12967 (N_12967,N_6978,N_6351);
and U12968 (N_12968,N_6062,N_7025);
xor U12969 (N_12969,N_5306,N_6399);
and U12970 (N_12970,N_8902,N_6638);
xnor U12971 (N_12971,N_9029,N_6593);
and U12972 (N_12972,N_8355,N_6833);
nand U12973 (N_12973,N_9340,N_7895);
nand U12974 (N_12974,N_6575,N_9108);
and U12975 (N_12975,N_6643,N_8231);
nand U12976 (N_12976,N_6513,N_5114);
nor U12977 (N_12977,N_7316,N_8953);
nand U12978 (N_12978,N_9062,N_6340);
nor U12979 (N_12979,N_7460,N_9856);
nor U12980 (N_12980,N_9725,N_5298);
xor U12981 (N_12981,N_9381,N_6475);
and U12982 (N_12982,N_7522,N_6053);
and U12983 (N_12983,N_7019,N_9380);
xnor U12984 (N_12984,N_9292,N_7770);
nand U12985 (N_12985,N_6638,N_5189);
xnor U12986 (N_12986,N_5455,N_7913);
nand U12987 (N_12987,N_7652,N_5998);
and U12988 (N_12988,N_9624,N_6298);
and U12989 (N_12989,N_5936,N_5627);
or U12990 (N_12990,N_7635,N_8738);
nor U12991 (N_12991,N_9889,N_9785);
or U12992 (N_12992,N_5486,N_8046);
nand U12993 (N_12993,N_7220,N_8774);
nor U12994 (N_12994,N_8638,N_7293);
or U12995 (N_12995,N_5345,N_7668);
nor U12996 (N_12996,N_6205,N_5571);
nor U12997 (N_12997,N_9039,N_8429);
and U12998 (N_12998,N_6734,N_6149);
or U12999 (N_12999,N_6965,N_6968);
or U13000 (N_13000,N_6205,N_8363);
and U13001 (N_13001,N_5169,N_5098);
nand U13002 (N_13002,N_8534,N_9853);
xnor U13003 (N_13003,N_9293,N_9736);
nor U13004 (N_13004,N_7774,N_8647);
xnor U13005 (N_13005,N_6501,N_5915);
nor U13006 (N_13006,N_6073,N_7284);
nand U13007 (N_13007,N_7066,N_7577);
or U13008 (N_13008,N_6718,N_8574);
xnor U13009 (N_13009,N_7263,N_5435);
xnor U13010 (N_13010,N_7143,N_5576);
or U13011 (N_13011,N_6565,N_8624);
nand U13012 (N_13012,N_7369,N_9165);
xnor U13013 (N_13013,N_8798,N_9091);
nor U13014 (N_13014,N_5827,N_9741);
and U13015 (N_13015,N_6310,N_8441);
or U13016 (N_13016,N_8576,N_7985);
xnor U13017 (N_13017,N_9177,N_7440);
nand U13018 (N_13018,N_6192,N_7877);
nor U13019 (N_13019,N_8747,N_5701);
nand U13020 (N_13020,N_5055,N_7938);
or U13021 (N_13021,N_7359,N_7632);
or U13022 (N_13022,N_5164,N_5151);
and U13023 (N_13023,N_8867,N_9171);
nor U13024 (N_13024,N_5259,N_9940);
and U13025 (N_13025,N_5522,N_6613);
or U13026 (N_13026,N_9553,N_8973);
and U13027 (N_13027,N_7940,N_9048);
xor U13028 (N_13028,N_7488,N_9295);
nand U13029 (N_13029,N_7772,N_6131);
xnor U13030 (N_13030,N_6007,N_6862);
nor U13031 (N_13031,N_8241,N_5296);
xor U13032 (N_13032,N_6380,N_6946);
xnor U13033 (N_13033,N_9681,N_8704);
or U13034 (N_13034,N_8816,N_7788);
nor U13035 (N_13035,N_6236,N_8997);
nand U13036 (N_13036,N_9704,N_9763);
nand U13037 (N_13037,N_7483,N_9999);
nand U13038 (N_13038,N_8562,N_5347);
nand U13039 (N_13039,N_7567,N_9493);
or U13040 (N_13040,N_7809,N_5337);
nand U13041 (N_13041,N_7472,N_6463);
and U13042 (N_13042,N_7986,N_7443);
xnor U13043 (N_13043,N_6494,N_7258);
and U13044 (N_13044,N_5393,N_8612);
nor U13045 (N_13045,N_9642,N_6313);
xnor U13046 (N_13046,N_7346,N_9653);
nor U13047 (N_13047,N_9167,N_9856);
and U13048 (N_13048,N_8438,N_8926);
nor U13049 (N_13049,N_6198,N_9046);
xor U13050 (N_13050,N_9362,N_7702);
and U13051 (N_13051,N_7777,N_8609);
nand U13052 (N_13052,N_8279,N_5819);
nor U13053 (N_13053,N_8657,N_7601);
xnor U13054 (N_13054,N_7324,N_7665);
nand U13055 (N_13055,N_8215,N_5751);
xnor U13056 (N_13056,N_8733,N_5662);
nor U13057 (N_13057,N_6188,N_6207);
and U13058 (N_13058,N_8582,N_6509);
nand U13059 (N_13059,N_8405,N_6526);
nor U13060 (N_13060,N_8066,N_6431);
xor U13061 (N_13061,N_9973,N_6246);
nand U13062 (N_13062,N_5540,N_6891);
nor U13063 (N_13063,N_7474,N_6223);
xor U13064 (N_13064,N_6664,N_5074);
nor U13065 (N_13065,N_7138,N_8377);
nor U13066 (N_13066,N_9325,N_9314);
nor U13067 (N_13067,N_9313,N_5572);
nor U13068 (N_13068,N_8603,N_9543);
nor U13069 (N_13069,N_8542,N_9052);
or U13070 (N_13070,N_9837,N_7412);
and U13071 (N_13071,N_6107,N_7692);
or U13072 (N_13072,N_9746,N_6840);
nor U13073 (N_13073,N_9149,N_7823);
xor U13074 (N_13074,N_9242,N_5895);
xor U13075 (N_13075,N_7715,N_8633);
and U13076 (N_13076,N_8766,N_7965);
xor U13077 (N_13077,N_9870,N_9001);
nand U13078 (N_13078,N_7798,N_5835);
nor U13079 (N_13079,N_7182,N_6766);
xor U13080 (N_13080,N_8764,N_9393);
and U13081 (N_13081,N_9584,N_9258);
nand U13082 (N_13082,N_9166,N_9729);
xor U13083 (N_13083,N_6303,N_6655);
or U13084 (N_13084,N_6829,N_9437);
and U13085 (N_13085,N_8632,N_5453);
xnor U13086 (N_13086,N_7014,N_9344);
xor U13087 (N_13087,N_6108,N_9125);
nand U13088 (N_13088,N_5585,N_7948);
nand U13089 (N_13089,N_5733,N_5520);
xor U13090 (N_13090,N_7753,N_8648);
or U13091 (N_13091,N_9138,N_5397);
or U13092 (N_13092,N_6222,N_5491);
nor U13093 (N_13093,N_8232,N_8052);
and U13094 (N_13094,N_7874,N_9462);
or U13095 (N_13095,N_8336,N_5972);
nand U13096 (N_13096,N_8409,N_5881);
nor U13097 (N_13097,N_7322,N_9707);
nand U13098 (N_13098,N_9977,N_5501);
nor U13099 (N_13099,N_7209,N_6653);
xnor U13100 (N_13100,N_5309,N_8287);
nor U13101 (N_13101,N_6990,N_8847);
nor U13102 (N_13102,N_6035,N_8450);
nand U13103 (N_13103,N_7093,N_9647);
nand U13104 (N_13104,N_9788,N_6934);
and U13105 (N_13105,N_9838,N_7653);
nor U13106 (N_13106,N_5694,N_8157);
xor U13107 (N_13107,N_8384,N_9411);
or U13108 (N_13108,N_6692,N_5558);
nand U13109 (N_13109,N_9181,N_8756);
nand U13110 (N_13110,N_9254,N_9586);
and U13111 (N_13111,N_8565,N_5902);
nand U13112 (N_13112,N_6649,N_5010);
xor U13113 (N_13113,N_9610,N_7019);
and U13114 (N_13114,N_6857,N_8486);
nor U13115 (N_13115,N_6380,N_6584);
nor U13116 (N_13116,N_9602,N_6691);
nor U13117 (N_13117,N_5305,N_9656);
xnor U13118 (N_13118,N_5492,N_7161);
xor U13119 (N_13119,N_6879,N_8787);
nand U13120 (N_13120,N_7693,N_5354);
and U13121 (N_13121,N_5724,N_5168);
or U13122 (N_13122,N_6176,N_9156);
nand U13123 (N_13123,N_9918,N_6760);
nor U13124 (N_13124,N_8268,N_9542);
nor U13125 (N_13125,N_8371,N_6067);
nand U13126 (N_13126,N_9034,N_9400);
nor U13127 (N_13127,N_9442,N_6507);
and U13128 (N_13128,N_7405,N_9808);
or U13129 (N_13129,N_7940,N_5112);
nor U13130 (N_13130,N_6234,N_6425);
or U13131 (N_13131,N_5447,N_9406);
or U13132 (N_13132,N_9006,N_7678);
and U13133 (N_13133,N_6359,N_7678);
xnor U13134 (N_13134,N_5703,N_5233);
or U13135 (N_13135,N_8485,N_5229);
and U13136 (N_13136,N_5633,N_7931);
or U13137 (N_13137,N_5430,N_8296);
nand U13138 (N_13138,N_6296,N_5674);
nor U13139 (N_13139,N_5991,N_9319);
xnor U13140 (N_13140,N_9986,N_7973);
and U13141 (N_13141,N_6020,N_6024);
nand U13142 (N_13142,N_5649,N_5388);
nand U13143 (N_13143,N_9369,N_6839);
and U13144 (N_13144,N_6783,N_6263);
xor U13145 (N_13145,N_7493,N_6334);
or U13146 (N_13146,N_8069,N_6051);
and U13147 (N_13147,N_7743,N_7187);
nand U13148 (N_13148,N_7002,N_8868);
and U13149 (N_13149,N_7473,N_9581);
and U13150 (N_13150,N_5556,N_8782);
xnor U13151 (N_13151,N_7978,N_5635);
nand U13152 (N_13152,N_5905,N_6328);
and U13153 (N_13153,N_6922,N_9170);
xor U13154 (N_13154,N_6930,N_6784);
or U13155 (N_13155,N_8409,N_5576);
nand U13156 (N_13156,N_6483,N_7711);
nor U13157 (N_13157,N_7798,N_6984);
nand U13158 (N_13158,N_6829,N_7738);
xor U13159 (N_13159,N_9991,N_8260);
nand U13160 (N_13160,N_5999,N_8779);
and U13161 (N_13161,N_7912,N_7608);
nor U13162 (N_13162,N_9345,N_8726);
nand U13163 (N_13163,N_9753,N_6402);
or U13164 (N_13164,N_9723,N_5088);
and U13165 (N_13165,N_9696,N_5505);
or U13166 (N_13166,N_7820,N_7129);
and U13167 (N_13167,N_6143,N_8301);
nand U13168 (N_13168,N_9821,N_5737);
nand U13169 (N_13169,N_9777,N_5760);
nand U13170 (N_13170,N_9913,N_8314);
xnor U13171 (N_13171,N_7143,N_6958);
nor U13172 (N_13172,N_5980,N_9469);
and U13173 (N_13173,N_9111,N_7152);
nor U13174 (N_13174,N_6520,N_8601);
or U13175 (N_13175,N_7028,N_6944);
nand U13176 (N_13176,N_6257,N_8371);
and U13177 (N_13177,N_8987,N_9212);
or U13178 (N_13178,N_5955,N_7724);
xor U13179 (N_13179,N_9451,N_9701);
xor U13180 (N_13180,N_6704,N_5653);
nor U13181 (N_13181,N_7564,N_9272);
and U13182 (N_13182,N_7493,N_8351);
and U13183 (N_13183,N_8310,N_7716);
nor U13184 (N_13184,N_8736,N_9470);
xor U13185 (N_13185,N_9595,N_9901);
xnor U13186 (N_13186,N_7787,N_6527);
or U13187 (N_13187,N_5121,N_8647);
or U13188 (N_13188,N_8372,N_5430);
and U13189 (N_13189,N_7720,N_9895);
xor U13190 (N_13190,N_6784,N_7372);
and U13191 (N_13191,N_8694,N_8641);
xnor U13192 (N_13192,N_9462,N_7147);
nand U13193 (N_13193,N_6006,N_5475);
or U13194 (N_13194,N_7751,N_9712);
and U13195 (N_13195,N_5330,N_5303);
nand U13196 (N_13196,N_7569,N_8925);
xor U13197 (N_13197,N_5771,N_5352);
or U13198 (N_13198,N_5065,N_7426);
or U13199 (N_13199,N_5629,N_7127);
nand U13200 (N_13200,N_7081,N_5522);
nor U13201 (N_13201,N_9545,N_5689);
nand U13202 (N_13202,N_5646,N_6371);
and U13203 (N_13203,N_9420,N_7207);
nor U13204 (N_13204,N_9731,N_9321);
or U13205 (N_13205,N_5329,N_6412);
xnor U13206 (N_13206,N_7760,N_7138);
xnor U13207 (N_13207,N_6422,N_6765);
nand U13208 (N_13208,N_5056,N_9902);
and U13209 (N_13209,N_7725,N_9824);
and U13210 (N_13210,N_6710,N_9927);
xor U13211 (N_13211,N_7445,N_8928);
xnor U13212 (N_13212,N_9300,N_8881);
xnor U13213 (N_13213,N_6390,N_6303);
xnor U13214 (N_13214,N_8504,N_8054);
and U13215 (N_13215,N_5168,N_5985);
and U13216 (N_13216,N_7708,N_6969);
xnor U13217 (N_13217,N_9421,N_6464);
nand U13218 (N_13218,N_5594,N_7771);
nand U13219 (N_13219,N_5449,N_9019);
or U13220 (N_13220,N_9429,N_9587);
and U13221 (N_13221,N_7112,N_7470);
and U13222 (N_13222,N_5754,N_6162);
and U13223 (N_13223,N_8407,N_7280);
nor U13224 (N_13224,N_7813,N_5679);
and U13225 (N_13225,N_6961,N_7915);
nand U13226 (N_13226,N_8534,N_6180);
nor U13227 (N_13227,N_6104,N_7199);
or U13228 (N_13228,N_5793,N_7211);
nand U13229 (N_13229,N_5952,N_6346);
or U13230 (N_13230,N_7352,N_5901);
nor U13231 (N_13231,N_9956,N_8245);
and U13232 (N_13232,N_6196,N_5069);
nand U13233 (N_13233,N_6571,N_5043);
nor U13234 (N_13234,N_8194,N_6243);
xnor U13235 (N_13235,N_6645,N_8872);
and U13236 (N_13236,N_8059,N_7385);
or U13237 (N_13237,N_9255,N_7975);
nor U13238 (N_13238,N_8646,N_6814);
xor U13239 (N_13239,N_8820,N_9622);
or U13240 (N_13240,N_9616,N_5892);
or U13241 (N_13241,N_5096,N_9920);
or U13242 (N_13242,N_7205,N_5980);
nor U13243 (N_13243,N_5116,N_5932);
or U13244 (N_13244,N_8334,N_6086);
nor U13245 (N_13245,N_6371,N_6768);
nand U13246 (N_13246,N_6260,N_5101);
and U13247 (N_13247,N_9343,N_7984);
xor U13248 (N_13248,N_7653,N_5245);
xor U13249 (N_13249,N_8560,N_7360);
or U13250 (N_13250,N_7392,N_6599);
nand U13251 (N_13251,N_9694,N_7570);
nand U13252 (N_13252,N_6155,N_6836);
nand U13253 (N_13253,N_7351,N_9066);
nand U13254 (N_13254,N_8252,N_5732);
xnor U13255 (N_13255,N_5660,N_6848);
xnor U13256 (N_13256,N_5046,N_7647);
nand U13257 (N_13257,N_6758,N_5507);
nand U13258 (N_13258,N_9221,N_5989);
xnor U13259 (N_13259,N_8788,N_7634);
nand U13260 (N_13260,N_6413,N_5328);
nand U13261 (N_13261,N_7039,N_6801);
xnor U13262 (N_13262,N_6085,N_8532);
xor U13263 (N_13263,N_9345,N_7379);
nor U13264 (N_13264,N_7036,N_8934);
nor U13265 (N_13265,N_8334,N_5187);
or U13266 (N_13266,N_6791,N_6758);
xnor U13267 (N_13267,N_9629,N_7408);
nand U13268 (N_13268,N_6429,N_9025);
nor U13269 (N_13269,N_5971,N_8085);
nor U13270 (N_13270,N_7834,N_9142);
xor U13271 (N_13271,N_6881,N_9241);
nand U13272 (N_13272,N_6772,N_8431);
nor U13273 (N_13273,N_6507,N_8475);
nor U13274 (N_13274,N_9667,N_6558);
and U13275 (N_13275,N_7772,N_9016);
and U13276 (N_13276,N_6701,N_6876);
or U13277 (N_13277,N_5229,N_6704);
and U13278 (N_13278,N_5636,N_9506);
xor U13279 (N_13279,N_6484,N_6179);
nor U13280 (N_13280,N_5765,N_9040);
and U13281 (N_13281,N_6714,N_6974);
nor U13282 (N_13282,N_6133,N_9204);
xor U13283 (N_13283,N_6787,N_8820);
xnor U13284 (N_13284,N_7486,N_8681);
and U13285 (N_13285,N_5649,N_6178);
nor U13286 (N_13286,N_7688,N_7812);
nand U13287 (N_13287,N_9152,N_5255);
xnor U13288 (N_13288,N_8450,N_8638);
and U13289 (N_13289,N_7523,N_6229);
xnor U13290 (N_13290,N_6734,N_5913);
xor U13291 (N_13291,N_7709,N_5855);
nand U13292 (N_13292,N_8805,N_6532);
xnor U13293 (N_13293,N_8152,N_5795);
xnor U13294 (N_13294,N_9472,N_5719);
or U13295 (N_13295,N_6082,N_9984);
or U13296 (N_13296,N_7559,N_5613);
and U13297 (N_13297,N_7544,N_5616);
nor U13298 (N_13298,N_7238,N_7399);
nand U13299 (N_13299,N_7256,N_8026);
nor U13300 (N_13300,N_9314,N_6578);
xor U13301 (N_13301,N_7419,N_6323);
and U13302 (N_13302,N_8821,N_8555);
nor U13303 (N_13303,N_9889,N_9065);
and U13304 (N_13304,N_5139,N_6943);
nand U13305 (N_13305,N_7678,N_9478);
nand U13306 (N_13306,N_7954,N_5119);
xnor U13307 (N_13307,N_8075,N_5464);
nor U13308 (N_13308,N_7029,N_8178);
nor U13309 (N_13309,N_7575,N_9874);
nand U13310 (N_13310,N_6584,N_7254);
xnor U13311 (N_13311,N_9523,N_6391);
nand U13312 (N_13312,N_5177,N_9755);
nand U13313 (N_13313,N_8863,N_9722);
xnor U13314 (N_13314,N_7713,N_9699);
and U13315 (N_13315,N_5934,N_9068);
and U13316 (N_13316,N_9696,N_5855);
xor U13317 (N_13317,N_7923,N_6156);
or U13318 (N_13318,N_6374,N_8283);
xnor U13319 (N_13319,N_6111,N_8394);
nor U13320 (N_13320,N_5393,N_8826);
nand U13321 (N_13321,N_8514,N_7730);
nand U13322 (N_13322,N_5540,N_9558);
or U13323 (N_13323,N_7628,N_7017);
xnor U13324 (N_13324,N_8633,N_8503);
xor U13325 (N_13325,N_7370,N_6719);
or U13326 (N_13326,N_5722,N_8920);
xnor U13327 (N_13327,N_6557,N_9042);
nor U13328 (N_13328,N_8277,N_9145);
and U13329 (N_13329,N_9830,N_8588);
and U13330 (N_13330,N_8066,N_5209);
nand U13331 (N_13331,N_9991,N_8818);
nor U13332 (N_13332,N_9184,N_7652);
nand U13333 (N_13333,N_5500,N_8428);
nor U13334 (N_13334,N_8864,N_6615);
xor U13335 (N_13335,N_6441,N_8985);
xor U13336 (N_13336,N_6072,N_7587);
or U13337 (N_13337,N_5274,N_5028);
xor U13338 (N_13338,N_8963,N_8274);
nor U13339 (N_13339,N_6456,N_6017);
nand U13340 (N_13340,N_7782,N_9380);
and U13341 (N_13341,N_6414,N_6591);
and U13342 (N_13342,N_6372,N_7951);
xor U13343 (N_13343,N_5774,N_9220);
nor U13344 (N_13344,N_8576,N_9314);
xor U13345 (N_13345,N_6012,N_8562);
xnor U13346 (N_13346,N_7708,N_5811);
and U13347 (N_13347,N_8520,N_5395);
or U13348 (N_13348,N_6816,N_6082);
nand U13349 (N_13349,N_8083,N_6253);
and U13350 (N_13350,N_9196,N_9494);
nand U13351 (N_13351,N_8051,N_8086);
nor U13352 (N_13352,N_6384,N_5158);
nand U13353 (N_13353,N_9388,N_6715);
or U13354 (N_13354,N_6890,N_8955);
or U13355 (N_13355,N_7164,N_5411);
or U13356 (N_13356,N_9148,N_7567);
nand U13357 (N_13357,N_5985,N_6790);
xor U13358 (N_13358,N_7044,N_7164);
or U13359 (N_13359,N_5823,N_9865);
nor U13360 (N_13360,N_6282,N_8498);
xnor U13361 (N_13361,N_6716,N_6821);
xor U13362 (N_13362,N_9849,N_6295);
or U13363 (N_13363,N_6128,N_5563);
nor U13364 (N_13364,N_9320,N_5910);
nand U13365 (N_13365,N_7584,N_8630);
and U13366 (N_13366,N_8892,N_9659);
and U13367 (N_13367,N_6864,N_5891);
and U13368 (N_13368,N_6758,N_8162);
and U13369 (N_13369,N_9026,N_7170);
or U13370 (N_13370,N_8447,N_6873);
xor U13371 (N_13371,N_8964,N_6200);
xor U13372 (N_13372,N_5702,N_8616);
xnor U13373 (N_13373,N_6306,N_8093);
or U13374 (N_13374,N_5635,N_5016);
or U13375 (N_13375,N_7256,N_7644);
xor U13376 (N_13376,N_9135,N_5359);
nand U13377 (N_13377,N_5311,N_6416);
nand U13378 (N_13378,N_9852,N_8413);
or U13379 (N_13379,N_6846,N_7318);
nor U13380 (N_13380,N_9689,N_8329);
and U13381 (N_13381,N_9927,N_8328);
nor U13382 (N_13382,N_7941,N_9159);
nor U13383 (N_13383,N_9492,N_5761);
or U13384 (N_13384,N_6555,N_6194);
nor U13385 (N_13385,N_5728,N_6911);
and U13386 (N_13386,N_9433,N_5969);
xor U13387 (N_13387,N_8698,N_9193);
xnor U13388 (N_13388,N_8500,N_8438);
and U13389 (N_13389,N_8651,N_9772);
and U13390 (N_13390,N_7745,N_6677);
xnor U13391 (N_13391,N_8874,N_8935);
and U13392 (N_13392,N_9297,N_8024);
and U13393 (N_13393,N_8491,N_9953);
or U13394 (N_13394,N_9779,N_8436);
xor U13395 (N_13395,N_6055,N_7359);
or U13396 (N_13396,N_7593,N_9003);
or U13397 (N_13397,N_7711,N_8677);
xor U13398 (N_13398,N_6371,N_8320);
xor U13399 (N_13399,N_8359,N_6010);
nor U13400 (N_13400,N_9182,N_5163);
or U13401 (N_13401,N_6644,N_8750);
nor U13402 (N_13402,N_6718,N_6488);
xnor U13403 (N_13403,N_8017,N_6929);
and U13404 (N_13404,N_7269,N_7811);
and U13405 (N_13405,N_8550,N_7922);
and U13406 (N_13406,N_7778,N_5366);
nor U13407 (N_13407,N_6261,N_7956);
and U13408 (N_13408,N_6714,N_5205);
nor U13409 (N_13409,N_5049,N_7086);
xor U13410 (N_13410,N_9693,N_6117);
and U13411 (N_13411,N_6195,N_8388);
nor U13412 (N_13412,N_6302,N_7912);
nand U13413 (N_13413,N_8919,N_8824);
or U13414 (N_13414,N_8952,N_5143);
or U13415 (N_13415,N_9316,N_5871);
or U13416 (N_13416,N_9603,N_7741);
and U13417 (N_13417,N_9268,N_8959);
xor U13418 (N_13418,N_5155,N_7727);
and U13419 (N_13419,N_5214,N_5979);
and U13420 (N_13420,N_5756,N_8700);
xnor U13421 (N_13421,N_5848,N_7574);
or U13422 (N_13422,N_8425,N_7124);
nand U13423 (N_13423,N_7072,N_9383);
nor U13424 (N_13424,N_5738,N_6054);
nand U13425 (N_13425,N_9943,N_9692);
xnor U13426 (N_13426,N_8013,N_5191);
and U13427 (N_13427,N_5507,N_7118);
or U13428 (N_13428,N_5743,N_7237);
nand U13429 (N_13429,N_7609,N_8860);
and U13430 (N_13430,N_6713,N_5864);
or U13431 (N_13431,N_9992,N_5044);
and U13432 (N_13432,N_9683,N_8894);
nor U13433 (N_13433,N_7569,N_7493);
and U13434 (N_13434,N_8088,N_8489);
or U13435 (N_13435,N_7534,N_6367);
or U13436 (N_13436,N_5097,N_5784);
nand U13437 (N_13437,N_6349,N_9845);
and U13438 (N_13438,N_6820,N_8030);
or U13439 (N_13439,N_8657,N_7519);
and U13440 (N_13440,N_7842,N_7987);
nor U13441 (N_13441,N_5929,N_7735);
nand U13442 (N_13442,N_9878,N_8825);
and U13443 (N_13443,N_8594,N_6748);
or U13444 (N_13444,N_8388,N_9126);
nand U13445 (N_13445,N_5487,N_6798);
nand U13446 (N_13446,N_9918,N_7229);
nor U13447 (N_13447,N_8439,N_7087);
and U13448 (N_13448,N_8248,N_6572);
nor U13449 (N_13449,N_5874,N_6003);
nand U13450 (N_13450,N_8118,N_6268);
and U13451 (N_13451,N_6977,N_7621);
and U13452 (N_13452,N_9312,N_8173);
or U13453 (N_13453,N_9508,N_5637);
xnor U13454 (N_13454,N_6047,N_6541);
xor U13455 (N_13455,N_9270,N_7260);
and U13456 (N_13456,N_6655,N_6562);
xor U13457 (N_13457,N_6881,N_8716);
or U13458 (N_13458,N_6420,N_6279);
nor U13459 (N_13459,N_5866,N_7854);
and U13460 (N_13460,N_7699,N_6135);
nor U13461 (N_13461,N_9259,N_8619);
or U13462 (N_13462,N_7818,N_5881);
nor U13463 (N_13463,N_5772,N_5854);
nand U13464 (N_13464,N_7766,N_7081);
nor U13465 (N_13465,N_6949,N_6488);
nand U13466 (N_13466,N_9705,N_6174);
and U13467 (N_13467,N_8599,N_5622);
xor U13468 (N_13468,N_5950,N_7610);
or U13469 (N_13469,N_9527,N_7732);
xnor U13470 (N_13470,N_7975,N_9200);
xor U13471 (N_13471,N_5692,N_7985);
or U13472 (N_13472,N_5727,N_5286);
and U13473 (N_13473,N_9621,N_8236);
nor U13474 (N_13474,N_8293,N_6406);
nand U13475 (N_13475,N_8883,N_9059);
or U13476 (N_13476,N_7414,N_9846);
and U13477 (N_13477,N_6855,N_6698);
or U13478 (N_13478,N_6094,N_9004);
or U13479 (N_13479,N_6455,N_8601);
nand U13480 (N_13480,N_7595,N_9098);
or U13481 (N_13481,N_9169,N_6897);
and U13482 (N_13482,N_9718,N_9443);
xnor U13483 (N_13483,N_5521,N_7556);
nor U13484 (N_13484,N_6255,N_6769);
nor U13485 (N_13485,N_9732,N_6304);
nand U13486 (N_13486,N_9372,N_7817);
and U13487 (N_13487,N_6727,N_6660);
xnor U13488 (N_13488,N_8264,N_8547);
and U13489 (N_13489,N_8368,N_9318);
xnor U13490 (N_13490,N_8997,N_9074);
or U13491 (N_13491,N_5624,N_6919);
and U13492 (N_13492,N_9735,N_5649);
xor U13493 (N_13493,N_5526,N_8789);
nand U13494 (N_13494,N_7130,N_6112);
and U13495 (N_13495,N_5397,N_7547);
nand U13496 (N_13496,N_8269,N_9170);
xor U13497 (N_13497,N_6042,N_8222);
and U13498 (N_13498,N_9860,N_6364);
nor U13499 (N_13499,N_7488,N_8802);
xnor U13500 (N_13500,N_7498,N_7466);
nand U13501 (N_13501,N_8007,N_8371);
and U13502 (N_13502,N_6770,N_6327);
and U13503 (N_13503,N_9062,N_8127);
xnor U13504 (N_13504,N_5665,N_6172);
nor U13505 (N_13505,N_9750,N_6586);
xnor U13506 (N_13506,N_9901,N_6227);
and U13507 (N_13507,N_6140,N_8553);
nor U13508 (N_13508,N_6611,N_9366);
and U13509 (N_13509,N_5955,N_6384);
and U13510 (N_13510,N_6219,N_6173);
nand U13511 (N_13511,N_9066,N_8818);
nor U13512 (N_13512,N_7350,N_9668);
or U13513 (N_13513,N_9909,N_7260);
xnor U13514 (N_13514,N_6294,N_9957);
and U13515 (N_13515,N_9808,N_9740);
and U13516 (N_13516,N_6246,N_9869);
nand U13517 (N_13517,N_5465,N_6127);
nor U13518 (N_13518,N_8457,N_5052);
xnor U13519 (N_13519,N_6699,N_7923);
and U13520 (N_13520,N_5313,N_8497);
xor U13521 (N_13521,N_5717,N_7661);
and U13522 (N_13522,N_8035,N_5911);
nor U13523 (N_13523,N_6586,N_7338);
or U13524 (N_13524,N_7016,N_7766);
and U13525 (N_13525,N_8429,N_8161);
xnor U13526 (N_13526,N_5805,N_8488);
or U13527 (N_13527,N_5714,N_5562);
or U13528 (N_13528,N_5557,N_7545);
xor U13529 (N_13529,N_9885,N_9500);
nor U13530 (N_13530,N_8716,N_6423);
nor U13531 (N_13531,N_6551,N_8739);
or U13532 (N_13532,N_5684,N_6378);
and U13533 (N_13533,N_8997,N_7497);
or U13534 (N_13534,N_5285,N_8376);
or U13535 (N_13535,N_8804,N_5483);
nand U13536 (N_13536,N_6206,N_9259);
nor U13537 (N_13537,N_6252,N_8760);
or U13538 (N_13538,N_6026,N_5201);
and U13539 (N_13539,N_7875,N_9884);
xnor U13540 (N_13540,N_5756,N_9871);
and U13541 (N_13541,N_8013,N_7813);
and U13542 (N_13542,N_6497,N_7626);
and U13543 (N_13543,N_9948,N_9539);
and U13544 (N_13544,N_9103,N_7887);
nand U13545 (N_13545,N_9100,N_6997);
xor U13546 (N_13546,N_9574,N_6055);
and U13547 (N_13547,N_7500,N_8961);
and U13548 (N_13548,N_5966,N_6560);
and U13549 (N_13549,N_6663,N_7965);
or U13550 (N_13550,N_8455,N_5742);
nand U13551 (N_13551,N_8736,N_5982);
xnor U13552 (N_13552,N_5859,N_5155);
nor U13553 (N_13553,N_8788,N_6444);
and U13554 (N_13554,N_9668,N_5491);
nor U13555 (N_13555,N_5095,N_8536);
or U13556 (N_13556,N_6954,N_5441);
xor U13557 (N_13557,N_7013,N_7970);
nor U13558 (N_13558,N_8132,N_8528);
nand U13559 (N_13559,N_8328,N_6621);
or U13560 (N_13560,N_7679,N_9763);
nand U13561 (N_13561,N_5714,N_7718);
xnor U13562 (N_13562,N_8552,N_6596);
or U13563 (N_13563,N_6226,N_8164);
and U13564 (N_13564,N_8583,N_6091);
or U13565 (N_13565,N_8396,N_9367);
xnor U13566 (N_13566,N_5400,N_5182);
nand U13567 (N_13567,N_6198,N_7992);
xor U13568 (N_13568,N_7690,N_6319);
and U13569 (N_13569,N_8788,N_5073);
nand U13570 (N_13570,N_8544,N_8796);
nor U13571 (N_13571,N_9797,N_9230);
nor U13572 (N_13572,N_6999,N_5288);
xor U13573 (N_13573,N_8319,N_7953);
nand U13574 (N_13574,N_5582,N_9792);
nor U13575 (N_13575,N_8574,N_9151);
nand U13576 (N_13576,N_6215,N_5527);
and U13577 (N_13577,N_7510,N_8747);
nor U13578 (N_13578,N_7564,N_9963);
xnor U13579 (N_13579,N_8905,N_7685);
or U13580 (N_13580,N_6445,N_9817);
and U13581 (N_13581,N_9958,N_5228);
xor U13582 (N_13582,N_8410,N_6263);
and U13583 (N_13583,N_8728,N_6513);
and U13584 (N_13584,N_8404,N_8731);
and U13585 (N_13585,N_6090,N_6835);
or U13586 (N_13586,N_6230,N_6024);
xor U13587 (N_13587,N_9154,N_7897);
nand U13588 (N_13588,N_7322,N_5400);
nor U13589 (N_13589,N_9914,N_6378);
or U13590 (N_13590,N_8518,N_5468);
xnor U13591 (N_13591,N_6711,N_7802);
nand U13592 (N_13592,N_9258,N_6543);
and U13593 (N_13593,N_7290,N_7932);
and U13594 (N_13594,N_6172,N_8176);
nor U13595 (N_13595,N_6660,N_7191);
or U13596 (N_13596,N_8655,N_7990);
or U13597 (N_13597,N_9430,N_9589);
xor U13598 (N_13598,N_9377,N_6290);
nand U13599 (N_13599,N_5160,N_9683);
xnor U13600 (N_13600,N_5985,N_5068);
nand U13601 (N_13601,N_8689,N_6425);
xor U13602 (N_13602,N_7997,N_6602);
xor U13603 (N_13603,N_6675,N_8551);
or U13604 (N_13604,N_7606,N_7049);
and U13605 (N_13605,N_5763,N_5330);
xor U13606 (N_13606,N_9459,N_8236);
xor U13607 (N_13607,N_7340,N_6180);
and U13608 (N_13608,N_8169,N_9238);
and U13609 (N_13609,N_5204,N_8303);
nor U13610 (N_13610,N_7454,N_8061);
or U13611 (N_13611,N_7791,N_5582);
and U13612 (N_13612,N_9546,N_6912);
xor U13613 (N_13613,N_7568,N_5244);
xnor U13614 (N_13614,N_9640,N_8619);
nor U13615 (N_13615,N_5257,N_6470);
and U13616 (N_13616,N_5635,N_5427);
nand U13617 (N_13617,N_6741,N_6074);
xor U13618 (N_13618,N_8759,N_7626);
nand U13619 (N_13619,N_9929,N_8470);
or U13620 (N_13620,N_7798,N_7849);
nand U13621 (N_13621,N_7412,N_8799);
or U13622 (N_13622,N_5816,N_5423);
nand U13623 (N_13623,N_7850,N_6696);
nand U13624 (N_13624,N_5357,N_6833);
xor U13625 (N_13625,N_9439,N_7667);
nand U13626 (N_13626,N_8212,N_9292);
or U13627 (N_13627,N_9565,N_8335);
nand U13628 (N_13628,N_6966,N_6880);
nor U13629 (N_13629,N_7441,N_6272);
and U13630 (N_13630,N_8731,N_7204);
xor U13631 (N_13631,N_5816,N_7177);
and U13632 (N_13632,N_9431,N_6067);
and U13633 (N_13633,N_9998,N_8397);
or U13634 (N_13634,N_5233,N_9840);
nand U13635 (N_13635,N_5556,N_9880);
nor U13636 (N_13636,N_5424,N_5312);
nand U13637 (N_13637,N_9791,N_7341);
nand U13638 (N_13638,N_8865,N_7123);
and U13639 (N_13639,N_5018,N_9651);
xnor U13640 (N_13640,N_5503,N_6436);
nor U13641 (N_13641,N_7244,N_7085);
and U13642 (N_13642,N_5157,N_9196);
nand U13643 (N_13643,N_7249,N_7852);
and U13644 (N_13644,N_7510,N_7278);
nand U13645 (N_13645,N_7991,N_8420);
or U13646 (N_13646,N_8923,N_8086);
nand U13647 (N_13647,N_7535,N_5592);
or U13648 (N_13648,N_9539,N_9303);
and U13649 (N_13649,N_8834,N_9256);
nor U13650 (N_13650,N_8510,N_9450);
or U13651 (N_13651,N_9103,N_8412);
nor U13652 (N_13652,N_9514,N_7717);
and U13653 (N_13653,N_7945,N_6772);
nor U13654 (N_13654,N_8224,N_8605);
or U13655 (N_13655,N_8900,N_6031);
and U13656 (N_13656,N_9329,N_7843);
and U13657 (N_13657,N_9352,N_7230);
nand U13658 (N_13658,N_7519,N_8177);
and U13659 (N_13659,N_8034,N_7327);
nand U13660 (N_13660,N_6578,N_7484);
nand U13661 (N_13661,N_8730,N_8225);
nor U13662 (N_13662,N_9224,N_8708);
nor U13663 (N_13663,N_5690,N_6224);
nand U13664 (N_13664,N_9965,N_7994);
nand U13665 (N_13665,N_9333,N_5281);
nor U13666 (N_13666,N_7826,N_8855);
nand U13667 (N_13667,N_7619,N_7691);
or U13668 (N_13668,N_6827,N_9345);
and U13669 (N_13669,N_5608,N_6392);
or U13670 (N_13670,N_5052,N_6304);
nor U13671 (N_13671,N_7371,N_9010);
nand U13672 (N_13672,N_5545,N_8801);
xnor U13673 (N_13673,N_8059,N_7606);
nand U13674 (N_13674,N_6866,N_7029);
and U13675 (N_13675,N_6594,N_6224);
or U13676 (N_13676,N_8631,N_5195);
nand U13677 (N_13677,N_5255,N_8413);
nor U13678 (N_13678,N_6927,N_5510);
or U13679 (N_13679,N_8106,N_8700);
or U13680 (N_13680,N_8136,N_9638);
nor U13681 (N_13681,N_7981,N_9028);
xor U13682 (N_13682,N_8515,N_6366);
xnor U13683 (N_13683,N_6770,N_5490);
xor U13684 (N_13684,N_5676,N_9340);
nor U13685 (N_13685,N_9552,N_8382);
xnor U13686 (N_13686,N_6068,N_5921);
nand U13687 (N_13687,N_7056,N_6003);
nand U13688 (N_13688,N_9831,N_8324);
nand U13689 (N_13689,N_8046,N_8188);
and U13690 (N_13690,N_7709,N_6508);
xor U13691 (N_13691,N_9197,N_9814);
nor U13692 (N_13692,N_5145,N_9850);
xnor U13693 (N_13693,N_5540,N_9924);
nand U13694 (N_13694,N_5664,N_5961);
xor U13695 (N_13695,N_6120,N_9675);
xor U13696 (N_13696,N_5892,N_5952);
or U13697 (N_13697,N_8864,N_6129);
nor U13698 (N_13698,N_7462,N_8838);
nor U13699 (N_13699,N_8749,N_9429);
nor U13700 (N_13700,N_6655,N_8033);
and U13701 (N_13701,N_9407,N_9855);
nor U13702 (N_13702,N_5089,N_9114);
xnor U13703 (N_13703,N_6198,N_8877);
xor U13704 (N_13704,N_8599,N_9074);
and U13705 (N_13705,N_7028,N_7230);
nor U13706 (N_13706,N_9330,N_7656);
xnor U13707 (N_13707,N_8606,N_9115);
and U13708 (N_13708,N_7004,N_8253);
nand U13709 (N_13709,N_6972,N_9069);
and U13710 (N_13710,N_8199,N_5470);
nand U13711 (N_13711,N_9782,N_5633);
xor U13712 (N_13712,N_6076,N_6714);
xor U13713 (N_13713,N_9627,N_9634);
nand U13714 (N_13714,N_6170,N_7805);
nor U13715 (N_13715,N_8397,N_6577);
xnor U13716 (N_13716,N_8649,N_5215);
nor U13717 (N_13717,N_5048,N_8029);
and U13718 (N_13718,N_8658,N_8885);
nand U13719 (N_13719,N_7832,N_7340);
or U13720 (N_13720,N_6934,N_7417);
or U13721 (N_13721,N_6627,N_9764);
nor U13722 (N_13722,N_6892,N_5953);
xnor U13723 (N_13723,N_8422,N_5620);
and U13724 (N_13724,N_9323,N_7226);
and U13725 (N_13725,N_5878,N_5020);
or U13726 (N_13726,N_7379,N_6280);
and U13727 (N_13727,N_6013,N_5174);
or U13728 (N_13728,N_6284,N_6713);
and U13729 (N_13729,N_9442,N_6041);
nor U13730 (N_13730,N_7933,N_6548);
or U13731 (N_13731,N_8613,N_8099);
or U13732 (N_13732,N_7111,N_9552);
xnor U13733 (N_13733,N_9076,N_8622);
nand U13734 (N_13734,N_5704,N_6173);
nand U13735 (N_13735,N_9804,N_7797);
and U13736 (N_13736,N_8955,N_5614);
nor U13737 (N_13737,N_6727,N_5995);
and U13738 (N_13738,N_5377,N_6162);
and U13739 (N_13739,N_9386,N_8134);
nor U13740 (N_13740,N_6100,N_5685);
or U13741 (N_13741,N_9273,N_7143);
nor U13742 (N_13742,N_8367,N_6755);
nand U13743 (N_13743,N_6129,N_6485);
xor U13744 (N_13744,N_8698,N_7374);
nand U13745 (N_13745,N_9290,N_8014);
nand U13746 (N_13746,N_9118,N_8342);
or U13747 (N_13747,N_5157,N_6530);
or U13748 (N_13748,N_8198,N_5241);
or U13749 (N_13749,N_5220,N_8780);
and U13750 (N_13750,N_5625,N_8162);
nand U13751 (N_13751,N_6238,N_9615);
nand U13752 (N_13752,N_6909,N_7757);
and U13753 (N_13753,N_7148,N_5231);
or U13754 (N_13754,N_8787,N_9147);
nor U13755 (N_13755,N_6271,N_6287);
nand U13756 (N_13756,N_8218,N_8073);
xnor U13757 (N_13757,N_5143,N_7991);
xnor U13758 (N_13758,N_8382,N_7111);
nor U13759 (N_13759,N_6996,N_6178);
nand U13760 (N_13760,N_5476,N_8560);
and U13761 (N_13761,N_7796,N_7038);
nand U13762 (N_13762,N_9095,N_9819);
nand U13763 (N_13763,N_7508,N_8950);
nand U13764 (N_13764,N_8031,N_7433);
nand U13765 (N_13765,N_5198,N_7427);
xor U13766 (N_13766,N_6073,N_7709);
nand U13767 (N_13767,N_7111,N_5569);
nand U13768 (N_13768,N_7827,N_6221);
or U13769 (N_13769,N_5082,N_9809);
xnor U13770 (N_13770,N_6876,N_5746);
xnor U13771 (N_13771,N_9746,N_5831);
nor U13772 (N_13772,N_5079,N_6122);
xnor U13773 (N_13773,N_9738,N_8140);
xor U13774 (N_13774,N_9076,N_5090);
xor U13775 (N_13775,N_9340,N_7162);
nand U13776 (N_13776,N_9450,N_6523);
xnor U13777 (N_13777,N_8372,N_6812);
nand U13778 (N_13778,N_6812,N_5389);
nor U13779 (N_13779,N_6256,N_5223);
or U13780 (N_13780,N_7307,N_9371);
nor U13781 (N_13781,N_5926,N_6891);
xnor U13782 (N_13782,N_5427,N_9514);
nand U13783 (N_13783,N_6874,N_8643);
nand U13784 (N_13784,N_8078,N_8191);
nand U13785 (N_13785,N_6775,N_9344);
or U13786 (N_13786,N_8005,N_5625);
nand U13787 (N_13787,N_7417,N_5985);
nand U13788 (N_13788,N_6550,N_5549);
nand U13789 (N_13789,N_6374,N_6769);
nand U13790 (N_13790,N_9050,N_8289);
xnor U13791 (N_13791,N_7539,N_9883);
and U13792 (N_13792,N_8074,N_5291);
and U13793 (N_13793,N_8079,N_7319);
and U13794 (N_13794,N_8815,N_6145);
or U13795 (N_13795,N_9429,N_8509);
xnor U13796 (N_13796,N_7291,N_5807);
nand U13797 (N_13797,N_7608,N_7035);
and U13798 (N_13798,N_5230,N_5614);
nor U13799 (N_13799,N_9563,N_5236);
nand U13800 (N_13800,N_8452,N_8547);
xor U13801 (N_13801,N_8157,N_9061);
and U13802 (N_13802,N_9790,N_9891);
nand U13803 (N_13803,N_6489,N_5976);
xnor U13804 (N_13804,N_7429,N_8424);
nand U13805 (N_13805,N_7889,N_7207);
nor U13806 (N_13806,N_8820,N_5070);
nor U13807 (N_13807,N_5973,N_8391);
nand U13808 (N_13808,N_5879,N_8880);
nor U13809 (N_13809,N_6819,N_9818);
or U13810 (N_13810,N_5745,N_7615);
nand U13811 (N_13811,N_6774,N_8851);
nor U13812 (N_13812,N_9582,N_9533);
xnor U13813 (N_13813,N_8970,N_6408);
xor U13814 (N_13814,N_7212,N_8744);
nor U13815 (N_13815,N_5688,N_9303);
or U13816 (N_13816,N_9413,N_9033);
nand U13817 (N_13817,N_6675,N_5333);
and U13818 (N_13818,N_7443,N_7644);
and U13819 (N_13819,N_6528,N_9766);
nor U13820 (N_13820,N_8982,N_8356);
or U13821 (N_13821,N_8515,N_6243);
and U13822 (N_13822,N_8022,N_9036);
or U13823 (N_13823,N_5451,N_8827);
xnor U13824 (N_13824,N_6376,N_8121);
xor U13825 (N_13825,N_8495,N_6063);
nor U13826 (N_13826,N_6929,N_6249);
xnor U13827 (N_13827,N_9515,N_5884);
xnor U13828 (N_13828,N_5132,N_7347);
nand U13829 (N_13829,N_8125,N_5295);
and U13830 (N_13830,N_6075,N_8848);
nand U13831 (N_13831,N_9599,N_9769);
or U13832 (N_13832,N_8853,N_6508);
nor U13833 (N_13833,N_9216,N_7231);
nand U13834 (N_13834,N_8046,N_8303);
nor U13835 (N_13835,N_5366,N_7483);
or U13836 (N_13836,N_8859,N_5436);
and U13837 (N_13837,N_7797,N_7568);
xnor U13838 (N_13838,N_9643,N_7745);
xnor U13839 (N_13839,N_7235,N_8884);
xor U13840 (N_13840,N_8301,N_5222);
and U13841 (N_13841,N_8365,N_7331);
or U13842 (N_13842,N_8584,N_7723);
nand U13843 (N_13843,N_7205,N_6164);
or U13844 (N_13844,N_6913,N_5513);
or U13845 (N_13845,N_5463,N_6272);
xnor U13846 (N_13846,N_5840,N_6048);
nand U13847 (N_13847,N_7352,N_9937);
or U13848 (N_13848,N_5735,N_7953);
nand U13849 (N_13849,N_5347,N_6968);
nand U13850 (N_13850,N_5740,N_8707);
or U13851 (N_13851,N_5316,N_7192);
xnor U13852 (N_13852,N_8989,N_9905);
nor U13853 (N_13853,N_9568,N_9281);
nor U13854 (N_13854,N_8074,N_7504);
nand U13855 (N_13855,N_6274,N_7340);
or U13856 (N_13856,N_7318,N_9110);
nand U13857 (N_13857,N_5623,N_5316);
and U13858 (N_13858,N_7968,N_5281);
nor U13859 (N_13859,N_7764,N_8907);
and U13860 (N_13860,N_5463,N_7050);
nor U13861 (N_13861,N_7736,N_8025);
xnor U13862 (N_13862,N_8495,N_7845);
xor U13863 (N_13863,N_7815,N_8222);
xnor U13864 (N_13864,N_6370,N_7831);
or U13865 (N_13865,N_6376,N_5079);
xor U13866 (N_13866,N_7431,N_5195);
and U13867 (N_13867,N_8132,N_7754);
nor U13868 (N_13868,N_5973,N_8124);
and U13869 (N_13869,N_9908,N_9525);
and U13870 (N_13870,N_5059,N_7649);
xnor U13871 (N_13871,N_9189,N_7353);
nand U13872 (N_13872,N_8648,N_5628);
and U13873 (N_13873,N_9982,N_9289);
or U13874 (N_13874,N_9414,N_5178);
or U13875 (N_13875,N_9640,N_5006);
nor U13876 (N_13876,N_5768,N_5810);
nor U13877 (N_13877,N_6770,N_9552);
or U13878 (N_13878,N_8576,N_9681);
or U13879 (N_13879,N_6303,N_5503);
xnor U13880 (N_13880,N_8287,N_7347);
or U13881 (N_13881,N_9443,N_6518);
or U13882 (N_13882,N_5654,N_7482);
nand U13883 (N_13883,N_5660,N_7691);
or U13884 (N_13884,N_5211,N_8117);
and U13885 (N_13885,N_8717,N_6685);
xnor U13886 (N_13886,N_8803,N_7327);
xnor U13887 (N_13887,N_6462,N_5913);
nor U13888 (N_13888,N_6747,N_8783);
and U13889 (N_13889,N_7380,N_7912);
xnor U13890 (N_13890,N_9912,N_6971);
xnor U13891 (N_13891,N_6283,N_7274);
nand U13892 (N_13892,N_9298,N_7138);
and U13893 (N_13893,N_7177,N_8997);
and U13894 (N_13894,N_9245,N_7825);
xnor U13895 (N_13895,N_7974,N_8709);
or U13896 (N_13896,N_7156,N_6066);
nor U13897 (N_13897,N_8296,N_9658);
xor U13898 (N_13898,N_6850,N_7068);
nor U13899 (N_13899,N_7484,N_9194);
or U13900 (N_13900,N_7888,N_8102);
nand U13901 (N_13901,N_5060,N_6638);
nand U13902 (N_13902,N_8835,N_9965);
xnor U13903 (N_13903,N_5081,N_5909);
or U13904 (N_13904,N_8214,N_5756);
nor U13905 (N_13905,N_5894,N_8257);
or U13906 (N_13906,N_5214,N_8825);
or U13907 (N_13907,N_5135,N_6060);
or U13908 (N_13908,N_7806,N_7296);
xor U13909 (N_13909,N_7007,N_5243);
nand U13910 (N_13910,N_9732,N_8031);
nand U13911 (N_13911,N_6753,N_7681);
nand U13912 (N_13912,N_6389,N_7580);
or U13913 (N_13913,N_7632,N_6985);
nand U13914 (N_13914,N_7081,N_5541);
nand U13915 (N_13915,N_7454,N_6132);
nor U13916 (N_13916,N_6703,N_7055);
nand U13917 (N_13917,N_8221,N_6985);
nor U13918 (N_13918,N_6140,N_6318);
xnor U13919 (N_13919,N_8905,N_5064);
and U13920 (N_13920,N_6231,N_5133);
or U13921 (N_13921,N_6348,N_6808);
nor U13922 (N_13922,N_7174,N_7080);
nand U13923 (N_13923,N_8534,N_9546);
and U13924 (N_13924,N_8059,N_8988);
and U13925 (N_13925,N_5156,N_8450);
nand U13926 (N_13926,N_7011,N_5522);
or U13927 (N_13927,N_6156,N_5734);
nor U13928 (N_13928,N_6640,N_6625);
nor U13929 (N_13929,N_5913,N_5038);
or U13930 (N_13930,N_9920,N_5202);
or U13931 (N_13931,N_7351,N_6671);
or U13932 (N_13932,N_9379,N_8897);
nand U13933 (N_13933,N_7261,N_9400);
or U13934 (N_13934,N_5727,N_7538);
or U13935 (N_13935,N_9861,N_5898);
xor U13936 (N_13936,N_5841,N_7269);
or U13937 (N_13937,N_5402,N_6367);
or U13938 (N_13938,N_9362,N_6153);
xor U13939 (N_13939,N_8777,N_5194);
or U13940 (N_13940,N_6384,N_9998);
xnor U13941 (N_13941,N_7526,N_6436);
or U13942 (N_13942,N_9403,N_6557);
xnor U13943 (N_13943,N_6476,N_7491);
or U13944 (N_13944,N_7226,N_7201);
and U13945 (N_13945,N_6672,N_7350);
nand U13946 (N_13946,N_7517,N_5651);
nor U13947 (N_13947,N_9419,N_7155);
nand U13948 (N_13948,N_9988,N_7215);
nand U13949 (N_13949,N_8085,N_7252);
and U13950 (N_13950,N_7083,N_6983);
xor U13951 (N_13951,N_5423,N_8487);
and U13952 (N_13952,N_9728,N_7900);
or U13953 (N_13953,N_7439,N_8386);
xnor U13954 (N_13954,N_7848,N_9210);
xnor U13955 (N_13955,N_5282,N_9471);
nand U13956 (N_13956,N_9832,N_8027);
or U13957 (N_13957,N_9692,N_7853);
xor U13958 (N_13958,N_8433,N_7814);
nor U13959 (N_13959,N_8742,N_7992);
nand U13960 (N_13960,N_5053,N_5761);
nor U13961 (N_13961,N_8277,N_5953);
or U13962 (N_13962,N_7244,N_7142);
or U13963 (N_13963,N_6979,N_9602);
and U13964 (N_13964,N_6311,N_8321);
nand U13965 (N_13965,N_5182,N_7557);
and U13966 (N_13966,N_8125,N_6915);
or U13967 (N_13967,N_7242,N_8979);
nand U13968 (N_13968,N_9249,N_5207);
nor U13969 (N_13969,N_5201,N_6024);
nand U13970 (N_13970,N_9224,N_7090);
nor U13971 (N_13971,N_7002,N_9703);
xor U13972 (N_13972,N_8732,N_6051);
and U13973 (N_13973,N_5153,N_5911);
nand U13974 (N_13974,N_5090,N_8168);
xnor U13975 (N_13975,N_5788,N_5224);
nand U13976 (N_13976,N_5294,N_9830);
and U13977 (N_13977,N_8802,N_6203);
or U13978 (N_13978,N_7429,N_6214);
xnor U13979 (N_13979,N_5692,N_6372);
nor U13980 (N_13980,N_9344,N_7666);
or U13981 (N_13981,N_7998,N_6373);
xnor U13982 (N_13982,N_9015,N_9280);
xor U13983 (N_13983,N_9125,N_7911);
nand U13984 (N_13984,N_6478,N_8381);
or U13985 (N_13985,N_8743,N_9821);
and U13986 (N_13986,N_9095,N_6525);
nand U13987 (N_13987,N_8199,N_7793);
xor U13988 (N_13988,N_7757,N_7239);
and U13989 (N_13989,N_9207,N_9948);
xor U13990 (N_13990,N_5756,N_9488);
nand U13991 (N_13991,N_9051,N_8611);
and U13992 (N_13992,N_6494,N_5901);
and U13993 (N_13993,N_6501,N_7412);
nand U13994 (N_13994,N_5671,N_9954);
nor U13995 (N_13995,N_6266,N_6453);
xnor U13996 (N_13996,N_7056,N_8833);
nor U13997 (N_13997,N_5262,N_5252);
or U13998 (N_13998,N_6679,N_7011);
nor U13999 (N_13999,N_9301,N_7227);
xnor U14000 (N_14000,N_8537,N_5267);
or U14001 (N_14001,N_9149,N_7177);
nor U14002 (N_14002,N_8137,N_9974);
nand U14003 (N_14003,N_7635,N_6032);
nand U14004 (N_14004,N_6719,N_6966);
or U14005 (N_14005,N_7818,N_9585);
nand U14006 (N_14006,N_6039,N_8094);
and U14007 (N_14007,N_9864,N_8998);
and U14008 (N_14008,N_7060,N_6674);
xor U14009 (N_14009,N_9626,N_6562);
xor U14010 (N_14010,N_9680,N_5112);
xnor U14011 (N_14011,N_6122,N_5406);
or U14012 (N_14012,N_9002,N_9651);
nand U14013 (N_14013,N_5643,N_6927);
and U14014 (N_14014,N_7960,N_9862);
nand U14015 (N_14015,N_9385,N_8654);
xor U14016 (N_14016,N_8587,N_6416);
nand U14017 (N_14017,N_5812,N_7247);
and U14018 (N_14018,N_5530,N_7744);
nand U14019 (N_14019,N_9741,N_6695);
nand U14020 (N_14020,N_9225,N_8649);
xnor U14021 (N_14021,N_6923,N_8811);
and U14022 (N_14022,N_5493,N_6652);
and U14023 (N_14023,N_5360,N_5488);
or U14024 (N_14024,N_7210,N_7778);
nor U14025 (N_14025,N_8960,N_6391);
xor U14026 (N_14026,N_7602,N_9964);
or U14027 (N_14027,N_6515,N_5596);
and U14028 (N_14028,N_5374,N_5540);
xnor U14029 (N_14029,N_9595,N_6852);
and U14030 (N_14030,N_8293,N_6121);
nor U14031 (N_14031,N_8136,N_9959);
xnor U14032 (N_14032,N_8674,N_7671);
or U14033 (N_14033,N_7645,N_5507);
and U14034 (N_14034,N_6355,N_6318);
and U14035 (N_14035,N_8863,N_9286);
or U14036 (N_14036,N_5363,N_8910);
nor U14037 (N_14037,N_8652,N_6212);
xor U14038 (N_14038,N_8998,N_7127);
and U14039 (N_14039,N_9320,N_7609);
or U14040 (N_14040,N_9675,N_8906);
and U14041 (N_14041,N_9079,N_6924);
nand U14042 (N_14042,N_6950,N_9995);
xor U14043 (N_14043,N_8423,N_9291);
and U14044 (N_14044,N_9519,N_6487);
nand U14045 (N_14045,N_6374,N_8037);
nand U14046 (N_14046,N_9769,N_9915);
xor U14047 (N_14047,N_6759,N_5681);
and U14048 (N_14048,N_8967,N_6683);
and U14049 (N_14049,N_8889,N_5552);
nor U14050 (N_14050,N_5799,N_6880);
xnor U14051 (N_14051,N_8785,N_5392);
or U14052 (N_14052,N_6475,N_6314);
xor U14053 (N_14053,N_7343,N_8467);
or U14054 (N_14054,N_8771,N_8569);
nor U14055 (N_14055,N_5763,N_6702);
and U14056 (N_14056,N_5543,N_9600);
and U14057 (N_14057,N_6331,N_8170);
nand U14058 (N_14058,N_6914,N_5470);
or U14059 (N_14059,N_9715,N_6952);
nor U14060 (N_14060,N_6361,N_7966);
xor U14061 (N_14061,N_8160,N_8223);
nor U14062 (N_14062,N_6474,N_8418);
nor U14063 (N_14063,N_5277,N_5611);
and U14064 (N_14064,N_5334,N_6846);
xnor U14065 (N_14065,N_7762,N_5145);
nand U14066 (N_14066,N_9540,N_7705);
and U14067 (N_14067,N_6126,N_5214);
or U14068 (N_14068,N_6851,N_9974);
nand U14069 (N_14069,N_6589,N_7882);
nor U14070 (N_14070,N_9055,N_6906);
xor U14071 (N_14071,N_7792,N_7916);
and U14072 (N_14072,N_7130,N_5250);
nand U14073 (N_14073,N_7488,N_6945);
nand U14074 (N_14074,N_6130,N_7759);
nor U14075 (N_14075,N_6300,N_7583);
xor U14076 (N_14076,N_9764,N_7028);
or U14077 (N_14077,N_5740,N_6325);
and U14078 (N_14078,N_8762,N_9221);
or U14079 (N_14079,N_6746,N_6035);
xnor U14080 (N_14080,N_9748,N_5631);
and U14081 (N_14081,N_5413,N_8852);
nor U14082 (N_14082,N_6497,N_6271);
or U14083 (N_14083,N_7724,N_9329);
xnor U14084 (N_14084,N_9138,N_9280);
xnor U14085 (N_14085,N_8043,N_7353);
nand U14086 (N_14086,N_9689,N_6443);
nor U14087 (N_14087,N_7075,N_9986);
or U14088 (N_14088,N_8301,N_7798);
nor U14089 (N_14089,N_6756,N_6762);
or U14090 (N_14090,N_8608,N_8556);
and U14091 (N_14091,N_8051,N_6200);
and U14092 (N_14092,N_7607,N_8840);
and U14093 (N_14093,N_6708,N_9465);
nor U14094 (N_14094,N_9545,N_5062);
nor U14095 (N_14095,N_8144,N_7874);
or U14096 (N_14096,N_8240,N_7635);
and U14097 (N_14097,N_8101,N_6127);
or U14098 (N_14098,N_8940,N_5721);
nand U14099 (N_14099,N_9596,N_8905);
or U14100 (N_14100,N_7327,N_7956);
nor U14101 (N_14101,N_9329,N_5206);
nor U14102 (N_14102,N_9765,N_8382);
or U14103 (N_14103,N_9641,N_5154);
nand U14104 (N_14104,N_8188,N_7946);
or U14105 (N_14105,N_9977,N_9108);
and U14106 (N_14106,N_9194,N_8290);
xor U14107 (N_14107,N_8138,N_5726);
or U14108 (N_14108,N_5587,N_5995);
xor U14109 (N_14109,N_9943,N_6869);
nor U14110 (N_14110,N_7546,N_5398);
or U14111 (N_14111,N_9001,N_8696);
xnor U14112 (N_14112,N_9700,N_9735);
xnor U14113 (N_14113,N_6346,N_8152);
or U14114 (N_14114,N_9723,N_6499);
nand U14115 (N_14115,N_9118,N_9582);
nor U14116 (N_14116,N_9616,N_6756);
or U14117 (N_14117,N_5280,N_8203);
nand U14118 (N_14118,N_8246,N_5638);
xnor U14119 (N_14119,N_6818,N_9209);
or U14120 (N_14120,N_6266,N_7657);
nor U14121 (N_14121,N_8430,N_5945);
nand U14122 (N_14122,N_9149,N_8169);
nor U14123 (N_14123,N_9918,N_9451);
nor U14124 (N_14124,N_9391,N_5323);
nand U14125 (N_14125,N_6534,N_5688);
nand U14126 (N_14126,N_7244,N_6922);
nand U14127 (N_14127,N_8739,N_9083);
and U14128 (N_14128,N_7315,N_9175);
and U14129 (N_14129,N_5333,N_8092);
or U14130 (N_14130,N_5586,N_8651);
or U14131 (N_14131,N_6508,N_7540);
nor U14132 (N_14132,N_6438,N_7343);
and U14133 (N_14133,N_5098,N_7680);
nor U14134 (N_14134,N_9896,N_8045);
nor U14135 (N_14135,N_9497,N_5987);
nand U14136 (N_14136,N_9799,N_5364);
and U14137 (N_14137,N_9936,N_7199);
nand U14138 (N_14138,N_5064,N_5344);
xnor U14139 (N_14139,N_7544,N_5816);
nand U14140 (N_14140,N_9235,N_8561);
nor U14141 (N_14141,N_9372,N_8488);
or U14142 (N_14142,N_6315,N_8158);
nand U14143 (N_14143,N_9420,N_7578);
or U14144 (N_14144,N_8569,N_7621);
nor U14145 (N_14145,N_9614,N_6891);
or U14146 (N_14146,N_7231,N_5692);
or U14147 (N_14147,N_8035,N_9030);
or U14148 (N_14148,N_5591,N_6459);
and U14149 (N_14149,N_6474,N_9536);
nand U14150 (N_14150,N_8747,N_6634);
nand U14151 (N_14151,N_8513,N_7013);
nand U14152 (N_14152,N_7566,N_9514);
or U14153 (N_14153,N_9911,N_7045);
and U14154 (N_14154,N_9428,N_7041);
nand U14155 (N_14155,N_7572,N_5446);
or U14156 (N_14156,N_7588,N_8968);
nor U14157 (N_14157,N_5301,N_9201);
and U14158 (N_14158,N_6471,N_6914);
nand U14159 (N_14159,N_5085,N_6988);
xnor U14160 (N_14160,N_8458,N_5821);
nor U14161 (N_14161,N_5316,N_6875);
xnor U14162 (N_14162,N_8440,N_7795);
nor U14163 (N_14163,N_7457,N_8493);
nor U14164 (N_14164,N_8503,N_6169);
nor U14165 (N_14165,N_5975,N_8057);
or U14166 (N_14166,N_7045,N_6664);
xor U14167 (N_14167,N_9910,N_5563);
nand U14168 (N_14168,N_6503,N_5328);
nor U14169 (N_14169,N_7842,N_8612);
nor U14170 (N_14170,N_9284,N_5243);
nand U14171 (N_14171,N_9550,N_7002);
nor U14172 (N_14172,N_8586,N_5292);
and U14173 (N_14173,N_8493,N_5057);
and U14174 (N_14174,N_7491,N_9377);
nand U14175 (N_14175,N_8168,N_7064);
nor U14176 (N_14176,N_7493,N_8515);
xor U14177 (N_14177,N_9297,N_5946);
nand U14178 (N_14178,N_6179,N_5770);
nand U14179 (N_14179,N_6439,N_5869);
nand U14180 (N_14180,N_7546,N_5124);
nor U14181 (N_14181,N_9818,N_5417);
xor U14182 (N_14182,N_9865,N_9294);
and U14183 (N_14183,N_9063,N_5818);
nor U14184 (N_14184,N_9918,N_9990);
nand U14185 (N_14185,N_8301,N_5306);
or U14186 (N_14186,N_5545,N_6949);
nor U14187 (N_14187,N_5392,N_5467);
nand U14188 (N_14188,N_6742,N_6662);
nor U14189 (N_14189,N_7791,N_7591);
and U14190 (N_14190,N_7813,N_8737);
nand U14191 (N_14191,N_6460,N_7648);
or U14192 (N_14192,N_6648,N_8319);
and U14193 (N_14193,N_8087,N_6242);
nand U14194 (N_14194,N_9579,N_7572);
xor U14195 (N_14195,N_8829,N_6935);
nand U14196 (N_14196,N_7739,N_6078);
xor U14197 (N_14197,N_9130,N_9104);
xor U14198 (N_14198,N_7314,N_9046);
or U14199 (N_14199,N_9949,N_9671);
xor U14200 (N_14200,N_8628,N_8369);
or U14201 (N_14201,N_5354,N_7345);
nor U14202 (N_14202,N_5531,N_6357);
xor U14203 (N_14203,N_6344,N_7984);
nor U14204 (N_14204,N_9709,N_5305);
or U14205 (N_14205,N_8006,N_6356);
and U14206 (N_14206,N_9649,N_7612);
xnor U14207 (N_14207,N_5415,N_5620);
nand U14208 (N_14208,N_9318,N_9823);
or U14209 (N_14209,N_7998,N_5584);
nor U14210 (N_14210,N_7849,N_9252);
xnor U14211 (N_14211,N_6249,N_9357);
xnor U14212 (N_14212,N_6709,N_7741);
xnor U14213 (N_14213,N_8963,N_5664);
and U14214 (N_14214,N_5625,N_9909);
nor U14215 (N_14215,N_7183,N_8037);
and U14216 (N_14216,N_6099,N_5320);
or U14217 (N_14217,N_8541,N_9792);
nor U14218 (N_14218,N_5526,N_7162);
nor U14219 (N_14219,N_7515,N_8698);
nand U14220 (N_14220,N_5174,N_5462);
and U14221 (N_14221,N_6356,N_6888);
and U14222 (N_14222,N_9701,N_7421);
xnor U14223 (N_14223,N_6416,N_5807);
xor U14224 (N_14224,N_5772,N_6582);
or U14225 (N_14225,N_8486,N_9831);
xnor U14226 (N_14226,N_9282,N_9189);
nor U14227 (N_14227,N_8347,N_8647);
nor U14228 (N_14228,N_7864,N_6813);
nor U14229 (N_14229,N_8134,N_9486);
and U14230 (N_14230,N_9094,N_8782);
or U14231 (N_14231,N_9622,N_7416);
and U14232 (N_14232,N_6728,N_5354);
xor U14233 (N_14233,N_5541,N_7057);
and U14234 (N_14234,N_6406,N_6089);
and U14235 (N_14235,N_5942,N_7243);
xor U14236 (N_14236,N_9778,N_7770);
nand U14237 (N_14237,N_6641,N_9148);
and U14238 (N_14238,N_5573,N_9787);
nand U14239 (N_14239,N_5168,N_7115);
nor U14240 (N_14240,N_5612,N_7227);
nor U14241 (N_14241,N_5547,N_8953);
and U14242 (N_14242,N_7852,N_9523);
nand U14243 (N_14243,N_9614,N_6904);
and U14244 (N_14244,N_6399,N_7309);
nor U14245 (N_14245,N_8285,N_5428);
and U14246 (N_14246,N_9925,N_7829);
xnor U14247 (N_14247,N_9243,N_9249);
or U14248 (N_14248,N_9117,N_5996);
nand U14249 (N_14249,N_6984,N_8086);
nand U14250 (N_14250,N_7521,N_6059);
nand U14251 (N_14251,N_5051,N_8952);
nand U14252 (N_14252,N_8926,N_5536);
and U14253 (N_14253,N_9210,N_8313);
nor U14254 (N_14254,N_8532,N_7993);
or U14255 (N_14255,N_8448,N_7140);
xnor U14256 (N_14256,N_9421,N_5709);
xnor U14257 (N_14257,N_6378,N_8217);
nand U14258 (N_14258,N_7627,N_8784);
nor U14259 (N_14259,N_8489,N_8192);
nand U14260 (N_14260,N_8538,N_7866);
or U14261 (N_14261,N_6608,N_5834);
nand U14262 (N_14262,N_9902,N_8288);
or U14263 (N_14263,N_7307,N_7800);
or U14264 (N_14264,N_5068,N_9642);
nor U14265 (N_14265,N_5938,N_6742);
or U14266 (N_14266,N_7010,N_7650);
nand U14267 (N_14267,N_8978,N_7724);
nand U14268 (N_14268,N_6930,N_5206);
and U14269 (N_14269,N_5638,N_8580);
nand U14270 (N_14270,N_5644,N_5687);
nor U14271 (N_14271,N_5968,N_6800);
nor U14272 (N_14272,N_8076,N_8611);
xor U14273 (N_14273,N_9071,N_9870);
or U14274 (N_14274,N_5422,N_7339);
xor U14275 (N_14275,N_9002,N_8875);
and U14276 (N_14276,N_6266,N_8904);
or U14277 (N_14277,N_6664,N_7032);
nor U14278 (N_14278,N_9162,N_8486);
and U14279 (N_14279,N_5234,N_9564);
xor U14280 (N_14280,N_9098,N_7845);
xor U14281 (N_14281,N_8493,N_7700);
and U14282 (N_14282,N_7391,N_9139);
xor U14283 (N_14283,N_9749,N_7124);
or U14284 (N_14284,N_7049,N_7331);
nor U14285 (N_14285,N_9698,N_6458);
or U14286 (N_14286,N_8069,N_8796);
or U14287 (N_14287,N_8361,N_7980);
xnor U14288 (N_14288,N_7064,N_9549);
and U14289 (N_14289,N_7376,N_6105);
and U14290 (N_14290,N_5980,N_7774);
and U14291 (N_14291,N_8698,N_7669);
and U14292 (N_14292,N_6135,N_9241);
xor U14293 (N_14293,N_7432,N_5094);
nand U14294 (N_14294,N_6844,N_8692);
nor U14295 (N_14295,N_6564,N_6707);
nor U14296 (N_14296,N_5080,N_5900);
nor U14297 (N_14297,N_5737,N_7797);
and U14298 (N_14298,N_8870,N_6103);
nor U14299 (N_14299,N_6518,N_7985);
nand U14300 (N_14300,N_6391,N_5815);
and U14301 (N_14301,N_7483,N_9835);
xor U14302 (N_14302,N_7283,N_8691);
nor U14303 (N_14303,N_5576,N_9977);
nor U14304 (N_14304,N_6361,N_7816);
and U14305 (N_14305,N_7055,N_7735);
xnor U14306 (N_14306,N_6266,N_5209);
xnor U14307 (N_14307,N_8389,N_8748);
or U14308 (N_14308,N_9750,N_6411);
nand U14309 (N_14309,N_8905,N_7823);
nand U14310 (N_14310,N_7197,N_6261);
and U14311 (N_14311,N_9108,N_5796);
nand U14312 (N_14312,N_9533,N_6996);
or U14313 (N_14313,N_9829,N_8358);
nor U14314 (N_14314,N_8363,N_8231);
and U14315 (N_14315,N_8824,N_5805);
nor U14316 (N_14316,N_8094,N_9469);
nor U14317 (N_14317,N_9976,N_9026);
nor U14318 (N_14318,N_8480,N_7022);
or U14319 (N_14319,N_7656,N_7331);
or U14320 (N_14320,N_5219,N_6320);
nor U14321 (N_14321,N_9326,N_7034);
nand U14322 (N_14322,N_5540,N_8068);
nor U14323 (N_14323,N_8882,N_9996);
and U14324 (N_14324,N_6467,N_5613);
nor U14325 (N_14325,N_8881,N_7743);
or U14326 (N_14326,N_5375,N_7020);
or U14327 (N_14327,N_7262,N_5710);
or U14328 (N_14328,N_9413,N_8957);
and U14329 (N_14329,N_6753,N_8468);
or U14330 (N_14330,N_9070,N_5664);
nor U14331 (N_14331,N_5616,N_5763);
or U14332 (N_14332,N_8270,N_8391);
or U14333 (N_14333,N_5147,N_5353);
and U14334 (N_14334,N_6789,N_5318);
xor U14335 (N_14335,N_7381,N_6508);
nor U14336 (N_14336,N_7674,N_7266);
and U14337 (N_14337,N_5774,N_7891);
nand U14338 (N_14338,N_7808,N_8266);
xnor U14339 (N_14339,N_8094,N_9336);
or U14340 (N_14340,N_7242,N_6419);
nand U14341 (N_14341,N_8242,N_5668);
and U14342 (N_14342,N_9368,N_5080);
xnor U14343 (N_14343,N_9955,N_5539);
xor U14344 (N_14344,N_7692,N_7211);
or U14345 (N_14345,N_5101,N_5286);
and U14346 (N_14346,N_5428,N_7708);
xnor U14347 (N_14347,N_9526,N_6899);
nor U14348 (N_14348,N_9074,N_5952);
nor U14349 (N_14349,N_9980,N_8484);
xnor U14350 (N_14350,N_8618,N_5314);
nand U14351 (N_14351,N_9515,N_6911);
or U14352 (N_14352,N_8858,N_5024);
and U14353 (N_14353,N_9534,N_7478);
xor U14354 (N_14354,N_5814,N_5762);
nand U14355 (N_14355,N_5067,N_9391);
or U14356 (N_14356,N_9036,N_6703);
and U14357 (N_14357,N_7130,N_5324);
or U14358 (N_14358,N_9246,N_6248);
nor U14359 (N_14359,N_6576,N_9024);
and U14360 (N_14360,N_5277,N_6925);
or U14361 (N_14361,N_6945,N_7709);
or U14362 (N_14362,N_8202,N_5973);
or U14363 (N_14363,N_6019,N_5916);
nor U14364 (N_14364,N_7714,N_5407);
xor U14365 (N_14365,N_8201,N_6700);
or U14366 (N_14366,N_5796,N_8342);
or U14367 (N_14367,N_5561,N_5173);
and U14368 (N_14368,N_8128,N_8620);
or U14369 (N_14369,N_8590,N_9718);
or U14370 (N_14370,N_9234,N_9534);
and U14371 (N_14371,N_6198,N_7712);
xnor U14372 (N_14372,N_5020,N_6761);
or U14373 (N_14373,N_8730,N_9084);
and U14374 (N_14374,N_8816,N_6744);
nor U14375 (N_14375,N_5604,N_9467);
xnor U14376 (N_14376,N_5184,N_6102);
xnor U14377 (N_14377,N_8793,N_5685);
nor U14378 (N_14378,N_6433,N_6354);
or U14379 (N_14379,N_9724,N_6445);
xnor U14380 (N_14380,N_9164,N_8129);
and U14381 (N_14381,N_6547,N_6581);
or U14382 (N_14382,N_6024,N_6394);
nor U14383 (N_14383,N_5801,N_8454);
or U14384 (N_14384,N_7353,N_8157);
xnor U14385 (N_14385,N_8743,N_8927);
and U14386 (N_14386,N_6378,N_6196);
and U14387 (N_14387,N_6513,N_5012);
nand U14388 (N_14388,N_9976,N_7337);
and U14389 (N_14389,N_8095,N_9568);
nor U14390 (N_14390,N_6367,N_9043);
nor U14391 (N_14391,N_5089,N_9167);
nor U14392 (N_14392,N_5710,N_7715);
or U14393 (N_14393,N_5625,N_5451);
nor U14394 (N_14394,N_7255,N_5267);
and U14395 (N_14395,N_9482,N_5336);
xor U14396 (N_14396,N_7448,N_7366);
and U14397 (N_14397,N_5922,N_8986);
and U14398 (N_14398,N_6166,N_8121);
nand U14399 (N_14399,N_7127,N_8162);
and U14400 (N_14400,N_9751,N_8319);
or U14401 (N_14401,N_6774,N_7283);
or U14402 (N_14402,N_6556,N_8873);
nand U14403 (N_14403,N_7713,N_5557);
or U14404 (N_14404,N_6964,N_5532);
nor U14405 (N_14405,N_5141,N_5940);
nand U14406 (N_14406,N_5446,N_5805);
nand U14407 (N_14407,N_9043,N_5639);
nor U14408 (N_14408,N_9777,N_7427);
nand U14409 (N_14409,N_6342,N_9171);
and U14410 (N_14410,N_9581,N_7645);
and U14411 (N_14411,N_7372,N_7317);
or U14412 (N_14412,N_5109,N_5588);
and U14413 (N_14413,N_6246,N_8489);
nor U14414 (N_14414,N_7132,N_8680);
xor U14415 (N_14415,N_5339,N_8414);
nor U14416 (N_14416,N_8355,N_5306);
or U14417 (N_14417,N_6400,N_6765);
xnor U14418 (N_14418,N_7942,N_5241);
nand U14419 (N_14419,N_8518,N_7003);
and U14420 (N_14420,N_8616,N_5219);
nor U14421 (N_14421,N_7528,N_7458);
xor U14422 (N_14422,N_5016,N_6393);
nand U14423 (N_14423,N_6717,N_7742);
nor U14424 (N_14424,N_5516,N_7368);
xor U14425 (N_14425,N_7566,N_6310);
nand U14426 (N_14426,N_8146,N_6892);
nor U14427 (N_14427,N_8684,N_8059);
nor U14428 (N_14428,N_5231,N_7676);
nand U14429 (N_14429,N_5171,N_9815);
nand U14430 (N_14430,N_8545,N_8926);
xnor U14431 (N_14431,N_8229,N_8144);
and U14432 (N_14432,N_5288,N_9791);
nand U14433 (N_14433,N_9749,N_9067);
and U14434 (N_14434,N_9232,N_8814);
nor U14435 (N_14435,N_7639,N_5467);
or U14436 (N_14436,N_7150,N_8533);
nand U14437 (N_14437,N_7857,N_6733);
or U14438 (N_14438,N_6190,N_8615);
xnor U14439 (N_14439,N_9579,N_6207);
or U14440 (N_14440,N_5612,N_6140);
and U14441 (N_14441,N_9516,N_6073);
nand U14442 (N_14442,N_8538,N_8311);
and U14443 (N_14443,N_6086,N_9431);
and U14444 (N_14444,N_5451,N_9384);
or U14445 (N_14445,N_6202,N_5024);
and U14446 (N_14446,N_9484,N_6906);
xor U14447 (N_14447,N_5024,N_8582);
or U14448 (N_14448,N_6889,N_7748);
nor U14449 (N_14449,N_6671,N_7637);
nand U14450 (N_14450,N_6274,N_6124);
or U14451 (N_14451,N_7777,N_9668);
xnor U14452 (N_14452,N_7331,N_8888);
and U14453 (N_14453,N_9906,N_7679);
xor U14454 (N_14454,N_9532,N_8201);
nor U14455 (N_14455,N_5167,N_5812);
and U14456 (N_14456,N_9773,N_6641);
or U14457 (N_14457,N_6306,N_9191);
xnor U14458 (N_14458,N_7481,N_6217);
and U14459 (N_14459,N_8430,N_5793);
xor U14460 (N_14460,N_7159,N_6140);
nand U14461 (N_14461,N_6635,N_8637);
and U14462 (N_14462,N_7941,N_9902);
xnor U14463 (N_14463,N_8101,N_6240);
and U14464 (N_14464,N_7275,N_7004);
nor U14465 (N_14465,N_5022,N_8495);
xor U14466 (N_14466,N_8911,N_8658);
nor U14467 (N_14467,N_7480,N_5384);
nor U14468 (N_14468,N_7987,N_6613);
and U14469 (N_14469,N_9370,N_7835);
nand U14470 (N_14470,N_9632,N_5412);
nor U14471 (N_14471,N_6542,N_9531);
or U14472 (N_14472,N_5837,N_7296);
or U14473 (N_14473,N_8890,N_8792);
xor U14474 (N_14474,N_7824,N_6274);
xnor U14475 (N_14475,N_7065,N_9657);
nand U14476 (N_14476,N_9463,N_7849);
xor U14477 (N_14477,N_6600,N_5307);
nor U14478 (N_14478,N_7573,N_5014);
nand U14479 (N_14479,N_5278,N_7191);
nor U14480 (N_14480,N_5392,N_6881);
or U14481 (N_14481,N_9296,N_7426);
or U14482 (N_14482,N_5022,N_8101);
xnor U14483 (N_14483,N_9143,N_7295);
nor U14484 (N_14484,N_6634,N_8493);
nor U14485 (N_14485,N_9322,N_6770);
and U14486 (N_14486,N_5090,N_9883);
nor U14487 (N_14487,N_6954,N_8081);
nor U14488 (N_14488,N_6650,N_6892);
nand U14489 (N_14489,N_5870,N_8001);
nor U14490 (N_14490,N_8849,N_7458);
nand U14491 (N_14491,N_9230,N_8970);
and U14492 (N_14492,N_8493,N_8325);
and U14493 (N_14493,N_9703,N_6621);
and U14494 (N_14494,N_5162,N_9920);
nand U14495 (N_14495,N_9591,N_6158);
nand U14496 (N_14496,N_5168,N_7549);
and U14497 (N_14497,N_7721,N_5505);
nand U14498 (N_14498,N_7369,N_9479);
xnor U14499 (N_14499,N_6503,N_8221);
and U14500 (N_14500,N_8826,N_9114);
nor U14501 (N_14501,N_5001,N_9801);
or U14502 (N_14502,N_8270,N_7985);
nor U14503 (N_14503,N_8798,N_9901);
nor U14504 (N_14504,N_7988,N_6672);
and U14505 (N_14505,N_9184,N_8337);
nand U14506 (N_14506,N_9466,N_6722);
xnor U14507 (N_14507,N_9511,N_8593);
or U14508 (N_14508,N_5334,N_7649);
nor U14509 (N_14509,N_9042,N_7556);
nand U14510 (N_14510,N_8841,N_5173);
nor U14511 (N_14511,N_6206,N_7570);
and U14512 (N_14512,N_5090,N_9239);
and U14513 (N_14513,N_6344,N_7709);
nand U14514 (N_14514,N_5378,N_5676);
and U14515 (N_14515,N_8125,N_7099);
nand U14516 (N_14516,N_5899,N_8999);
and U14517 (N_14517,N_9348,N_8334);
nand U14518 (N_14518,N_7899,N_8148);
and U14519 (N_14519,N_5432,N_8907);
nand U14520 (N_14520,N_5161,N_8066);
nand U14521 (N_14521,N_9034,N_6669);
nor U14522 (N_14522,N_5794,N_7586);
nor U14523 (N_14523,N_5351,N_9068);
xnor U14524 (N_14524,N_6801,N_8705);
and U14525 (N_14525,N_5016,N_9530);
nand U14526 (N_14526,N_8681,N_6265);
or U14527 (N_14527,N_8569,N_7036);
nor U14528 (N_14528,N_8265,N_6396);
and U14529 (N_14529,N_8890,N_9747);
and U14530 (N_14530,N_8953,N_5204);
nand U14531 (N_14531,N_5718,N_5142);
nand U14532 (N_14532,N_6906,N_6931);
nor U14533 (N_14533,N_8191,N_9618);
xnor U14534 (N_14534,N_8514,N_9142);
or U14535 (N_14535,N_9333,N_5406);
xor U14536 (N_14536,N_9842,N_8633);
nor U14537 (N_14537,N_7320,N_7885);
xnor U14538 (N_14538,N_6356,N_9173);
or U14539 (N_14539,N_7275,N_5023);
and U14540 (N_14540,N_6677,N_7517);
and U14541 (N_14541,N_6447,N_8804);
or U14542 (N_14542,N_5424,N_9507);
nand U14543 (N_14543,N_5333,N_9606);
and U14544 (N_14544,N_5249,N_8133);
nand U14545 (N_14545,N_7387,N_7548);
or U14546 (N_14546,N_6467,N_9804);
or U14547 (N_14547,N_5894,N_9654);
nor U14548 (N_14548,N_8216,N_5406);
nor U14549 (N_14549,N_7033,N_9337);
or U14550 (N_14550,N_9518,N_6051);
and U14551 (N_14551,N_7228,N_8847);
and U14552 (N_14552,N_9873,N_9766);
or U14553 (N_14553,N_9313,N_7980);
and U14554 (N_14554,N_6665,N_6597);
nand U14555 (N_14555,N_6496,N_5603);
nor U14556 (N_14556,N_9623,N_5701);
nor U14557 (N_14557,N_7575,N_9984);
nor U14558 (N_14558,N_6551,N_9638);
xor U14559 (N_14559,N_6323,N_5623);
or U14560 (N_14560,N_7026,N_6142);
and U14561 (N_14561,N_9347,N_6645);
nor U14562 (N_14562,N_5109,N_9147);
and U14563 (N_14563,N_6399,N_9077);
and U14564 (N_14564,N_8437,N_8984);
and U14565 (N_14565,N_5747,N_8451);
nand U14566 (N_14566,N_9169,N_9467);
or U14567 (N_14567,N_6075,N_9807);
nand U14568 (N_14568,N_6022,N_9957);
xor U14569 (N_14569,N_8345,N_5967);
and U14570 (N_14570,N_5404,N_8648);
xnor U14571 (N_14571,N_8533,N_8618);
xor U14572 (N_14572,N_8930,N_6320);
nor U14573 (N_14573,N_6433,N_7629);
and U14574 (N_14574,N_9531,N_8638);
or U14575 (N_14575,N_8527,N_8245);
and U14576 (N_14576,N_8678,N_7632);
or U14577 (N_14577,N_6928,N_7403);
nand U14578 (N_14578,N_5436,N_8523);
and U14579 (N_14579,N_7303,N_8149);
nand U14580 (N_14580,N_6443,N_6961);
nor U14581 (N_14581,N_6901,N_7786);
and U14582 (N_14582,N_6557,N_6570);
nand U14583 (N_14583,N_7969,N_9193);
and U14584 (N_14584,N_7013,N_6929);
nand U14585 (N_14585,N_8321,N_6517);
or U14586 (N_14586,N_6788,N_9451);
or U14587 (N_14587,N_9621,N_7870);
xor U14588 (N_14588,N_5267,N_7643);
or U14589 (N_14589,N_7449,N_9439);
nor U14590 (N_14590,N_6083,N_5499);
nor U14591 (N_14591,N_5151,N_9826);
or U14592 (N_14592,N_5196,N_9429);
nor U14593 (N_14593,N_9022,N_6961);
nand U14594 (N_14594,N_9107,N_5896);
xor U14595 (N_14595,N_8323,N_6957);
xnor U14596 (N_14596,N_6336,N_5249);
xor U14597 (N_14597,N_6011,N_6458);
nand U14598 (N_14598,N_6288,N_6723);
or U14599 (N_14599,N_9594,N_6870);
and U14600 (N_14600,N_8102,N_5053);
xor U14601 (N_14601,N_7135,N_8093);
and U14602 (N_14602,N_7895,N_6804);
xor U14603 (N_14603,N_9449,N_9712);
and U14604 (N_14604,N_9224,N_8047);
nand U14605 (N_14605,N_7245,N_7046);
nand U14606 (N_14606,N_7703,N_9600);
nand U14607 (N_14607,N_6786,N_8477);
xnor U14608 (N_14608,N_6083,N_9769);
nor U14609 (N_14609,N_7569,N_7921);
or U14610 (N_14610,N_7087,N_5211);
and U14611 (N_14611,N_9609,N_6245);
nor U14612 (N_14612,N_5792,N_6877);
nor U14613 (N_14613,N_9170,N_6025);
xnor U14614 (N_14614,N_8770,N_6227);
nor U14615 (N_14615,N_6103,N_8748);
nand U14616 (N_14616,N_6518,N_8513);
nor U14617 (N_14617,N_8765,N_6921);
nor U14618 (N_14618,N_7703,N_6880);
and U14619 (N_14619,N_9538,N_5273);
nand U14620 (N_14620,N_8537,N_6350);
nand U14621 (N_14621,N_7595,N_5998);
or U14622 (N_14622,N_5083,N_7261);
or U14623 (N_14623,N_5230,N_6429);
or U14624 (N_14624,N_5199,N_6663);
nor U14625 (N_14625,N_7874,N_7204);
nand U14626 (N_14626,N_7292,N_6270);
nor U14627 (N_14627,N_8389,N_9411);
nand U14628 (N_14628,N_7337,N_8766);
nor U14629 (N_14629,N_7063,N_9989);
and U14630 (N_14630,N_9898,N_7956);
and U14631 (N_14631,N_6607,N_9340);
and U14632 (N_14632,N_9360,N_8845);
nor U14633 (N_14633,N_9085,N_5661);
nor U14634 (N_14634,N_6676,N_9341);
or U14635 (N_14635,N_6395,N_9646);
nor U14636 (N_14636,N_5693,N_5296);
nor U14637 (N_14637,N_8695,N_8236);
or U14638 (N_14638,N_8996,N_6627);
nand U14639 (N_14639,N_7615,N_6738);
and U14640 (N_14640,N_9273,N_7421);
and U14641 (N_14641,N_9836,N_7780);
nor U14642 (N_14642,N_9582,N_9925);
nor U14643 (N_14643,N_6239,N_7347);
and U14644 (N_14644,N_9539,N_9278);
xnor U14645 (N_14645,N_6292,N_7188);
or U14646 (N_14646,N_8140,N_5169);
nand U14647 (N_14647,N_6884,N_6603);
nor U14648 (N_14648,N_7300,N_5331);
xor U14649 (N_14649,N_7379,N_6591);
nor U14650 (N_14650,N_6980,N_9579);
or U14651 (N_14651,N_5504,N_5344);
xnor U14652 (N_14652,N_7301,N_8212);
and U14653 (N_14653,N_5888,N_7195);
or U14654 (N_14654,N_8455,N_7141);
or U14655 (N_14655,N_6975,N_5799);
and U14656 (N_14656,N_9975,N_6878);
nand U14657 (N_14657,N_8848,N_5724);
nor U14658 (N_14658,N_5471,N_7572);
and U14659 (N_14659,N_9017,N_6657);
and U14660 (N_14660,N_5642,N_8468);
or U14661 (N_14661,N_7742,N_9179);
nand U14662 (N_14662,N_9700,N_5469);
and U14663 (N_14663,N_7666,N_5780);
nor U14664 (N_14664,N_7255,N_7682);
or U14665 (N_14665,N_9457,N_8481);
nor U14666 (N_14666,N_8311,N_6567);
xor U14667 (N_14667,N_7573,N_7586);
or U14668 (N_14668,N_5395,N_9826);
nor U14669 (N_14669,N_5305,N_8552);
or U14670 (N_14670,N_9748,N_6260);
nor U14671 (N_14671,N_6252,N_7476);
and U14672 (N_14672,N_8506,N_9418);
nand U14673 (N_14673,N_5429,N_9110);
or U14674 (N_14674,N_7009,N_9300);
xnor U14675 (N_14675,N_9082,N_5404);
xnor U14676 (N_14676,N_5355,N_6223);
and U14677 (N_14677,N_7625,N_9146);
nor U14678 (N_14678,N_8265,N_7147);
and U14679 (N_14679,N_6883,N_8676);
nand U14680 (N_14680,N_6382,N_9493);
xnor U14681 (N_14681,N_5573,N_8795);
nor U14682 (N_14682,N_7070,N_9524);
nand U14683 (N_14683,N_8288,N_7004);
nor U14684 (N_14684,N_7427,N_7590);
and U14685 (N_14685,N_8536,N_5433);
nand U14686 (N_14686,N_6489,N_5987);
nand U14687 (N_14687,N_8073,N_5230);
nand U14688 (N_14688,N_7658,N_6778);
xnor U14689 (N_14689,N_5801,N_7312);
nor U14690 (N_14690,N_9197,N_7155);
xor U14691 (N_14691,N_7067,N_8328);
nand U14692 (N_14692,N_7872,N_5070);
xor U14693 (N_14693,N_5031,N_6880);
nand U14694 (N_14694,N_6299,N_9233);
nor U14695 (N_14695,N_7236,N_7643);
nor U14696 (N_14696,N_8977,N_9382);
xnor U14697 (N_14697,N_6825,N_7356);
nor U14698 (N_14698,N_8421,N_8011);
nand U14699 (N_14699,N_8296,N_5456);
xor U14700 (N_14700,N_9959,N_8260);
xnor U14701 (N_14701,N_7176,N_6771);
nor U14702 (N_14702,N_5542,N_5702);
nand U14703 (N_14703,N_5652,N_9456);
or U14704 (N_14704,N_8105,N_8176);
nor U14705 (N_14705,N_7598,N_7040);
and U14706 (N_14706,N_9810,N_5219);
xor U14707 (N_14707,N_5810,N_7695);
nand U14708 (N_14708,N_9291,N_5555);
xnor U14709 (N_14709,N_9536,N_9022);
nor U14710 (N_14710,N_9593,N_7498);
xor U14711 (N_14711,N_6377,N_7448);
and U14712 (N_14712,N_9884,N_9593);
xor U14713 (N_14713,N_8405,N_5964);
or U14714 (N_14714,N_9724,N_9434);
nor U14715 (N_14715,N_8384,N_8740);
or U14716 (N_14716,N_9318,N_8010);
nand U14717 (N_14717,N_6986,N_9420);
and U14718 (N_14718,N_7979,N_9949);
and U14719 (N_14719,N_7258,N_8499);
xor U14720 (N_14720,N_6502,N_7761);
nand U14721 (N_14721,N_5863,N_9194);
nand U14722 (N_14722,N_6060,N_9215);
and U14723 (N_14723,N_9872,N_6691);
nand U14724 (N_14724,N_6995,N_9574);
nor U14725 (N_14725,N_5575,N_5465);
or U14726 (N_14726,N_5352,N_7317);
xnor U14727 (N_14727,N_9767,N_6209);
nand U14728 (N_14728,N_6268,N_9443);
or U14729 (N_14729,N_5845,N_9485);
nand U14730 (N_14730,N_8390,N_7698);
nor U14731 (N_14731,N_6600,N_7074);
and U14732 (N_14732,N_6293,N_8030);
and U14733 (N_14733,N_7720,N_6507);
xnor U14734 (N_14734,N_7923,N_6767);
xor U14735 (N_14735,N_7946,N_8872);
nand U14736 (N_14736,N_8593,N_9533);
and U14737 (N_14737,N_8872,N_7556);
nand U14738 (N_14738,N_9031,N_9833);
or U14739 (N_14739,N_7785,N_9319);
xor U14740 (N_14740,N_8875,N_7364);
and U14741 (N_14741,N_7294,N_9526);
and U14742 (N_14742,N_8514,N_5071);
or U14743 (N_14743,N_5930,N_6023);
nand U14744 (N_14744,N_6882,N_9888);
and U14745 (N_14745,N_7369,N_5904);
xor U14746 (N_14746,N_8652,N_5545);
or U14747 (N_14747,N_5477,N_5859);
xnor U14748 (N_14748,N_9129,N_8910);
nand U14749 (N_14749,N_5579,N_5465);
xor U14750 (N_14750,N_5799,N_5727);
nor U14751 (N_14751,N_9012,N_9634);
or U14752 (N_14752,N_7981,N_7090);
nand U14753 (N_14753,N_9700,N_5445);
and U14754 (N_14754,N_5143,N_7250);
or U14755 (N_14755,N_6197,N_9555);
and U14756 (N_14756,N_7991,N_9873);
xor U14757 (N_14757,N_8510,N_8770);
nor U14758 (N_14758,N_8096,N_5187);
nand U14759 (N_14759,N_7598,N_7070);
or U14760 (N_14760,N_7909,N_5262);
xor U14761 (N_14761,N_8066,N_7530);
nor U14762 (N_14762,N_7859,N_9798);
and U14763 (N_14763,N_5632,N_9683);
or U14764 (N_14764,N_6122,N_5237);
nand U14765 (N_14765,N_8765,N_7813);
or U14766 (N_14766,N_5052,N_8775);
or U14767 (N_14767,N_6879,N_9699);
and U14768 (N_14768,N_6501,N_8232);
nor U14769 (N_14769,N_7805,N_7415);
nor U14770 (N_14770,N_6169,N_8270);
nor U14771 (N_14771,N_5482,N_8954);
xor U14772 (N_14772,N_5802,N_6316);
or U14773 (N_14773,N_6717,N_9724);
and U14774 (N_14774,N_7866,N_5320);
or U14775 (N_14775,N_5979,N_6220);
xnor U14776 (N_14776,N_9425,N_5280);
nand U14777 (N_14777,N_8620,N_9031);
nor U14778 (N_14778,N_9363,N_9116);
xor U14779 (N_14779,N_9261,N_8771);
and U14780 (N_14780,N_8395,N_6228);
xnor U14781 (N_14781,N_5485,N_8333);
nand U14782 (N_14782,N_8113,N_9302);
xor U14783 (N_14783,N_6748,N_5427);
and U14784 (N_14784,N_5041,N_8019);
nand U14785 (N_14785,N_5918,N_9266);
or U14786 (N_14786,N_6879,N_7210);
nor U14787 (N_14787,N_5548,N_9828);
and U14788 (N_14788,N_5825,N_8157);
nor U14789 (N_14789,N_9603,N_6283);
and U14790 (N_14790,N_7969,N_6259);
xor U14791 (N_14791,N_9197,N_7345);
or U14792 (N_14792,N_6143,N_9668);
or U14793 (N_14793,N_6666,N_5313);
xnor U14794 (N_14794,N_5603,N_8716);
nand U14795 (N_14795,N_8404,N_9077);
nor U14796 (N_14796,N_9730,N_8894);
or U14797 (N_14797,N_6128,N_6209);
nand U14798 (N_14798,N_7930,N_5454);
nand U14799 (N_14799,N_8597,N_7092);
xor U14800 (N_14800,N_9947,N_6352);
or U14801 (N_14801,N_5571,N_5162);
nand U14802 (N_14802,N_9199,N_5754);
xor U14803 (N_14803,N_5686,N_7139);
nand U14804 (N_14804,N_7797,N_9194);
and U14805 (N_14805,N_6765,N_5007);
or U14806 (N_14806,N_8243,N_8329);
and U14807 (N_14807,N_7703,N_5572);
nor U14808 (N_14808,N_8584,N_9497);
or U14809 (N_14809,N_7808,N_8383);
or U14810 (N_14810,N_6463,N_8155);
nor U14811 (N_14811,N_8779,N_7194);
and U14812 (N_14812,N_8292,N_6879);
xor U14813 (N_14813,N_5850,N_6764);
nor U14814 (N_14814,N_9955,N_5265);
xor U14815 (N_14815,N_8601,N_6000);
nor U14816 (N_14816,N_5666,N_5588);
or U14817 (N_14817,N_6044,N_7421);
nor U14818 (N_14818,N_8909,N_8253);
nand U14819 (N_14819,N_7076,N_5182);
xnor U14820 (N_14820,N_7966,N_8755);
and U14821 (N_14821,N_9106,N_5010);
nand U14822 (N_14822,N_8935,N_7485);
xnor U14823 (N_14823,N_5688,N_8810);
or U14824 (N_14824,N_5128,N_6316);
and U14825 (N_14825,N_7665,N_6790);
and U14826 (N_14826,N_8094,N_7659);
xnor U14827 (N_14827,N_5683,N_9096);
and U14828 (N_14828,N_6597,N_9200);
nor U14829 (N_14829,N_5427,N_8769);
or U14830 (N_14830,N_7314,N_6538);
nor U14831 (N_14831,N_9520,N_7205);
and U14832 (N_14832,N_6347,N_8230);
and U14833 (N_14833,N_5019,N_7863);
and U14834 (N_14834,N_7064,N_8852);
nor U14835 (N_14835,N_8508,N_9129);
or U14836 (N_14836,N_7472,N_5934);
and U14837 (N_14837,N_5398,N_6884);
xnor U14838 (N_14838,N_7849,N_7580);
xnor U14839 (N_14839,N_9505,N_5840);
nand U14840 (N_14840,N_5200,N_9583);
and U14841 (N_14841,N_6524,N_5001);
nand U14842 (N_14842,N_7470,N_6684);
nor U14843 (N_14843,N_9460,N_9978);
nand U14844 (N_14844,N_5761,N_9372);
or U14845 (N_14845,N_5338,N_9001);
nor U14846 (N_14846,N_8044,N_6201);
and U14847 (N_14847,N_6004,N_9904);
or U14848 (N_14848,N_5187,N_6464);
or U14849 (N_14849,N_7249,N_9045);
nand U14850 (N_14850,N_8657,N_8231);
xor U14851 (N_14851,N_9386,N_6383);
nand U14852 (N_14852,N_6230,N_9096);
nor U14853 (N_14853,N_7901,N_7122);
and U14854 (N_14854,N_7809,N_7028);
or U14855 (N_14855,N_5796,N_7289);
nor U14856 (N_14856,N_8331,N_9522);
xor U14857 (N_14857,N_5610,N_9487);
and U14858 (N_14858,N_9737,N_6542);
nor U14859 (N_14859,N_9132,N_8234);
nor U14860 (N_14860,N_9953,N_7584);
or U14861 (N_14861,N_7561,N_8840);
nor U14862 (N_14862,N_5112,N_6222);
and U14863 (N_14863,N_6468,N_7701);
or U14864 (N_14864,N_9158,N_5400);
nand U14865 (N_14865,N_8790,N_6558);
nor U14866 (N_14866,N_7865,N_7445);
nand U14867 (N_14867,N_5391,N_8193);
or U14868 (N_14868,N_9712,N_8362);
and U14869 (N_14869,N_8317,N_9624);
xnor U14870 (N_14870,N_9901,N_7074);
xnor U14871 (N_14871,N_6363,N_9128);
nor U14872 (N_14872,N_7148,N_8739);
nor U14873 (N_14873,N_8914,N_6271);
or U14874 (N_14874,N_8437,N_8691);
xor U14875 (N_14875,N_9313,N_5806);
or U14876 (N_14876,N_5863,N_6009);
or U14877 (N_14877,N_7893,N_9519);
and U14878 (N_14878,N_9973,N_5033);
xor U14879 (N_14879,N_5690,N_9358);
or U14880 (N_14880,N_6606,N_9547);
xor U14881 (N_14881,N_5849,N_7249);
and U14882 (N_14882,N_6238,N_7167);
nor U14883 (N_14883,N_6990,N_5445);
nor U14884 (N_14884,N_7850,N_8046);
nand U14885 (N_14885,N_6857,N_6913);
or U14886 (N_14886,N_6386,N_8071);
nor U14887 (N_14887,N_6512,N_9053);
or U14888 (N_14888,N_7622,N_8564);
nand U14889 (N_14889,N_7539,N_9195);
nand U14890 (N_14890,N_7496,N_8803);
nand U14891 (N_14891,N_6215,N_8901);
and U14892 (N_14892,N_8498,N_8207);
or U14893 (N_14893,N_8078,N_7564);
nand U14894 (N_14894,N_7208,N_5731);
and U14895 (N_14895,N_7321,N_5435);
xor U14896 (N_14896,N_8698,N_7242);
or U14897 (N_14897,N_7198,N_9147);
nor U14898 (N_14898,N_5424,N_9787);
and U14899 (N_14899,N_7758,N_7666);
nand U14900 (N_14900,N_9104,N_7974);
or U14901 (N_14901,N_8380,N_7839);
and U14902 (N_14902,N_8920,N_8335);
and U14903 (N_14903,N_5309,N_6884);
nor U14904 (N_14904,N_5102,N_5059);
or U14905 (N_14905,N_5030,N_9123);
nand U14906 (N_14906,N_9862,N_9555);
nand U14907 (N_14907,N_7671,N_6288);
and U14908 (N_14908,N_5166,N_8292);
xnor U14909 (N_14909,N_5381,N_8790);
nor U14910 (N_14910,N_5332,N_5316);
xor U14911 (N_14911,N_8175,N_7460);
or U14912 (N_14912,N_6173,N_6061);
xor U14913 (N_14913,N_9871,N_5740);
and U14914 (N_14914,N_7425,N_7123);
or U14915 (N_14915,N_5303,N_5974);
nor U14916 (N_14916,N_5092,N_8266);
xnor U14917 (N_14917,N_9550,N_8475);
nand U14918 (N_14918,N_6984,N_5314);
and U14919 (N_14919,N_9400,N_5894);
and U14920 (N_14920,N_6325,N_8304);
and U14921 (N_14921,N_6391,N_7501);
xnor U14922 (N_14922,N_9505,N_6055);
nor U14923 (N_14923,N_8155,N_6636);
or U14924 (N_14924,N_9668,N_9601);
nand U14925 (N_14925,N_8381,N_5154);
or U14926 (N_14926,N_6294,N_5409);
nor U14927 (N_14927,N_5327,N_6825);
or U14928 (N_14928,N_8847,N_5436);
nor U14929 (N_14929,N_9017,N_7591);
or U14930 (N_14930,N_8110,N_9197);
xor U14931 (N_14931,N_5110,N_9347);
or U14932 (N_14932,N_7686,N_7250);
nand U14933 (N_14933,N_6112,N_6599);
xnor U14934 (N_14934,N_5082,N_6370);
nand U14935 (N_14935,N_5989,N_5740);
or U14936 (N_14936,N_9862,N_7147);
nor U14937 (N_14937,N_9763,N_5475);
or U14938 (N_14938,N_5207,N_5928);
or U14939 (N_14939,N_9686,N_8679);
nand U14940 (N_14940,N_8487,N_7310);
nor U14941 (N_14941,N_7505,N_7643);
or U14942 (N_14942,N_8827,N_5245);
nand U14943 (N_14943,N_5875,N_5238);
nand U14944 (N_14944,N_8096,N_7634);
or U14945 (N_14945,N_7124,N_5011);
or U14946 (N_14946,N_8797,N_5363);
nand U14947 (N_14947,N_6800,N_9988);
nor U14948 (N_14948,N_7715,N_9506);
nand U14949 (N_14949,N_8019,N_5139);
nor U14950 (N_14950,N_9975,N_9695);
or U14951 (N_14951,N_9494,N_8274);
or U14952 (N_14952,N_9746,N_8221);
and U14953 (N_14953,N_9053,N_9421);
xor U14954 (N_14954,N_6442,N_8474);
or U14955 (N_14955,N_8411,N_7073);
nand U14956 (N_14956,N_9296,N_5727);
or U14957 (N_14957,N_7590,N_9491);
xnor U14958 (N_14958,N_6369,N_8211);
or U14959 (N_14959,N_6974,N_7473);
and U14960 (N_14960,N_6574,N_7289);
or U14961 (N_14961,N_5281,N_9981);
nor U14962 (N_14962,N_9665,N_8494);
and U14963 (N_14963,N_6315,N_5588);
and U14964 (N_14964,N_7408,N_8528);
nor U14965 (N_14965,N_7748,N_7615);
or U14966 (N_14966,N_5059,N_6801);
and U14967 (N_14967,N_6158,N_6005);
and U14968 (N_14968,N_7480,N_5338);
xor U14969 (N_14969,N_9175,N_8028);
and U14970 (N_14970,N_5514,N_5510);
or U14971 (N_14971,N_7571,N_5729);
nor U14972 (N_14972,N_6541,N_9816);
nand U14973 (N_14973,N_7254,N_6223);
nand U14974 (N_14974,N_5551,N_9852);
nand U14975 (N_14975,N_9969,N_6386);
and U14976 (N_14976,N_6390,N_9180);
nand U14977 (N_14977,N_7086,N_8345);
nand U14978 (N_14978,N_8057,N_8261);
nand U14979 (N_14979,N_9580,N_8175);
and U14980 (N_14980,N_6583,N_8739);
and U14981 (N_14981,N_5254,N_6212);
and U14982 (N_14982,N_7418,N_7524);
and U14983 (N_14983,N_7891,N_8768);
and U14984 (N_14984,N_6381,N_8272);
xor U14985 (N_14985,N_9749,N_9666);
xnor U14986 (N_14986,N_7271,N_6228);
nand U14987 (N_14987,N_5557,N_8612);
or U14988 (N_14988,N_5124,N_5042);
and U14989 (N_14989,N_8153,N_9297);
and U14990 (N_14990,N_5214,N_9411);
xnor U14991 (N_14991,N_8449,N_5191);
and U14992 (N_14992,N_9134,N_8544);
and U14993 (N_14993,N_9774,N_5757);
nor U14994 (N_14994,N_6763,N_5380);
xnor U14995 (N_14995,N_8548,N_8853);
and U14996 (N_14996,N_5984,N_8292);
or U14997 (N_14997,N_5025,N_6915);
xor U14998 (N_14998,N_6993,N_5522);
nand U14999 (N_14999,N_7466,N_7909);
nor U15000 (N_15000,N_11598,N_14752);
and U15001 (N_15001,N_12340,N_13802);
nor U15002 (N_15002,N_11159,N_11651);
nor U15003 (N_15003,N_12150,N_10491);
xnor U15004 (N_15004,N_12321,N_14700);
or U15005 (N_15005,N_10326,N_10955);
xnor U15006 (N_15006,N_13780,N_11989);
or U15007 (N_15007,N_10696,N_10007);
or U15008 (N_15008,N_12147,N_13675);
nor U15009 (N_15009,N_12322,N_12248);
and U15010 (N_15010,N_11256,N_12880);
nand U15011 (N_15011,N_12582,N_12157);
nor U15012 (N_15012,N_11603,N_10868);
and U15013 (N_15013,N_10161,N_12085);
nor U15014 (N_15014,N_11125,N_12726);
nand U15015 (N_15015,N_12914,N_10486);
nor U15016 (N_15016,N_13018,N_14532);
nand U15017 (N_15017,N_12634,N_14530);
nor U15018 (N_15018,N_13432,N_10543);
and U15019 (N_15019,N_14090,N_10873);
and U15020 (N_15020,N_14824,N_14765);
or U15021 (N_15021,N_13824,N_10946);
nand U15022 (N_15022,N_14014,N_10714);
or U15023 (N_15023,N_11414,N_10431);
nand U15024 (N_15024,N_10321,N_14629);
nor U15025 (N_15025,N_11253,N_13427);
xnor U15026 (N_15026,N_14266,N_14357);
xor U15027 (N_15027,N_14243,N_14725);
or U15028 (N_15028,N_13852,N_11747);
and U15029 (N_15029,N_13647,N_11756);
and U15030 (N_15030,N_14408,N_13561);
and U15031 (N_15031,N_12264,N_10823);
nor U15032 (N_15032,N_10464,N_13634);
nor U15033 (N_15033,N_14662,N_10273);
or U15034 (N_15034,N_13810,N_14773);
or U15035 (N_15035,N_12204,N_10647);
nor U15036 (N_15036,N_11086,N_10481);
nand U15037 (N_15037,N_12183,N_13145);
or U15038 (N_15038,N_12168,N_13407);
or U15039 (N_15039,N_10104,N_10318);
nor U15040 (N_15040,N_10772,N_14779);
xnor U15041 (N_15041,N_12612,N_14488);
nand U15042 (N_15042,N_13158,N_12754);
nor U15043 (N_15043,N_14802,N_14427);
nor U15044 (N_15044,N_12929,N_14068);
nand U15045 (N_15045,N_11996,N_14180);
and U15046 (N_15046,N_12367,N_13028);
xnor U15047 (N_15047,N_12934,N_13701);
and U15048 (N_15048,N_12959,N_11302);
nor U15049 (N_15049,N_14064,N_14193);
or U15050 (N_15050,N_14581,N_13200);
and U15051 (N_15051,N_10448,N_11542);
and U15052 (N_15052,N_10409,N_12283);
nor U15053 (N_15053,N_14609,N_10537);
or U15054 (N_15054,N_13431,N_13651);
nor U15055 (N_15055,N_11047,N_12190);
or U15056 (N_15056,N_12558,N_14447);
and U15057 (N_15057,N_12678,N_14424);
and U15058 (N_15058,N_11306,N_10351);
nor U15059 (N_15059,N_14350,N_11232);
nand U15060 (N_15060,N_12623,N_14345);
or U15061 (N_15061,N_12456,N_12108);
xor U15062 (N_15062,N_12775,N_12960);
xor U15063 (N_15063,N_11568,N_14285);
and U15064 (N_15064,N_10971,N_10003);
nand U15065 (N_15065,N_14711,N_11399);
nand U15066 (N_15066,N_11121,N_10432);
nand U15067 (N_15067,N_13104,N_12566);
xnor U15068 (N_15068,N_14258,N_13749);
nand U15069 (N_15069,N_14928,N_13392);
or U15070 (N_15070,N_14132,N_12382);
nor U15071 (N_15071,N_13494,N_11553);
or U15072 (N_15072,N_12691,N_12557);
and U15073 (N_15073,N_12835,N_10836);
xor U15074 (N_15074,N_13899,N_11498);
xnor U15075 (N_15075,N_12770,N_13015);
nor U15076 (N_15076,N_10757,N_14944);
or U15077 (N_15077,N_10586,N_11029);
xor U15078 (N_15078,N_10435,N_10992);
xnor U15079 (N_15079,N_12496,N_13667);
and U15080 (N_15080,N_10081,N_11055);
and U15081 (N_15081,N_13459,N_14709);
xor U15082 (N_15082,N_11693,N_14081);
xor U15083 (N_15083,N_11641,N_11026);
nor U15084 (N_15084,N_14766,N_12832);
nand U15085 (N_15085,N_11209,N_10581);
and U15086 (N_15086,N_11290,N_11742);
and U15087 (N_15087,N_12453,N_12102);
and U15088 (N_15088,N_11751,N_12621);
nand U15089 (N_15089,N_13702,N_14087);
or U15090 (N_15090,N_10952,N_13763);
or U15091 (N_15091,N_13272,N_13411);
nand U15092 (N_15092,N_14103,N_13574);
nand U15093 (N_15093,N_11995,N_14411);
or U15094 (N_15094,N_12261,N_13515);
nor U15095 (N_15095,N_12166,N_12945);
xnor U15096 (N_15096,N_13744,N_11176);
nand U15097 (N_15097,N_13951,N_14888);
or U15098 (N_15098,N_12710,N_13241);
nand U15099 (N_15099,N_11769,N_12984);
xnor U15100 (N_15100,N_11350,N_14853);
xnor U15101 (N_15101,N_12266,N_12611);
or U15102 (N_15102,N_12796,N_14994);
nor U15103 (N_15103,N_12311,N_12620);
xnor U15104 (N_15104,N_13134,N_11247);
nor U15105 (N_15105,N_12193,N_13090);
and U15106 (N_15106,N_14204,N_11223);
and U15107 (N_15107,N_14242,N_13179);
and U15108 (N_15108,N_11636,N_10482);
nor U15109 (N_15109,N_12257,N_12199);
xor U15110 (N_15110,N_13017,N_12830);
xnor U15111 (N_15111,N_11975,N_10433);
or U15112 (N_15112,N_13854,N_14474);
or U15113 (N_15113,N_10341,N_11738);
and U15114 (N_15114,N_11311,N_11065);
or U15115 (N_15115,N_11936,N_13990);
nor U15116 (N_15116,N_14328,N_10426);
nand U15117 (N_15117,N_12990,N_11168);
or U15118 (N_15118,N_10562,N_12347);
xnor U15119 (N_15119,N_10851,N_11563);
xnor U15120 (N_15120,N_11551,N_14030);
xnor U15121 (N_15121,N_14852,N_11073);
nor U15122 (N_15122,N_14987,N_12731);
and U15123 (N_15123,N_12436,N_12454);
and U15124 (N_15124,N_11405,N_10191);
or U15125 (N_15125,N_11803,N_11666);
nand U15126 (N_15126,N_14714,N_10393);
nand U15127 (N_15127,N_11404,N_13299);
or U15128 (N_15128,N_11415,N_13313);
nor U15129 (N_15129,N_10792,N_13855);
xor U15130 (N_15130,N_13528,N_11074);
and U15131 (N_15131,N_11658,N_12250);
nand U15132 (N_15132,N_13929,N_13026);
or U15133 (N_15133,N_14848,N_11943);
and U15134 (N_15134,N_13805,N_12317);
nor U15135 (N_15135,N_13013,N_12702);
nor U15136 (N_15136,N_14673,N_11338);
nor U15137 (N_15137,N_11972,N_14572);
xor U15138 (N_15138,N_12887,N_13493);
nor U15139 (N_15139,N_14067,N_10347);
or U15140 (N_15140,N_13434,N_14120);
or U15141 (N_15141,N_13117,N_12227);
and U15142 (N_15142,N_13745,N_11200);
nand U15143 (N_15143,N_14943,N_11783);
and U15144 (N_15144,N_12536,N_12253);
nand U15145 (N_15145,N_10332,N_14906);
nor U15146 (N_15146,N_11204,N_12053);
nand U15147 (N_15147,N_12370,N_14229);
xor U15148 (N_15148,N_10374,N_14294);
and U15149 (N_15149,N_10826,N_11565);
nand U15150 (N_15150,N_11499,N_11011);
and U15151 (N_15151,N_14201,N_11827);
and U15152 (N_15152,N_10532,N_11661);
and U15153 (N_15153,N_12735,N_10678);
and U15154 (N_15154,N_12553,N_10730);
nor U15155 (N_15155,N_12782,N_14797);
nor U15156 (N_15156,N_14835,N_11013);
xnor U15157 (N_15157,N_11591,N_13441);
xnor U15158 (N_15158,N_12290,N_11562);
or U15159 (N_15159,N_10066,N_12245);
or U15160 (N_15160,N_13338,N_11838);
xor U15161 (N_15161,N_12416,N_14856);
nand U15162 (N_15162,N_14825,N_11703);
nand U15163 (N_15163,N_11508,N_11167);
or U15164 (N_15164,N_13361,N_11805);
xor U15165 (N_15165,N_11813,N_10812);
nor U15166 (N_15166,N_12368,N_10376);
nand U15167 (N_15167,N_14384,N_10014);
or U15168 (N_15168,N_11123,N_13303);
nor U15169 (N_15169,N_12985,N_14615);
nand U15170 (N_15170,N_11888,N_13778);
or U15171 (N_15171,N_13624,N_13697);
and U15172 (N_15172,N_11667,N_10858);
nor U15173 (N_15173,N_10020,N_13927);
or U15174 (N_15174,N_10369,N_13497);
xnor U15175 (N_15175,N_13022,N_14753);
nor U15176 (N_15176,N_14050,N_13753);
and U15177 (N_15177,N_11673,N_12997);
and U15178 (N_15178,N_10987,N_13069);
and U15179 (N_15179,N_14860,N_11211);
and U15180 (N_15180,N_13189,N_10650);
and U15181 (N_15181,N_13663,N_14513);
and U15182 (N_15182,N_14890,N_10886);
nand U15183 (N_15183,N_14054,N_14181);
or U15184 (N_15184,N_11064,N_12451);
xnor U15185 (N_15185,N_13264,N_14227);
and U15186 (N_15186,N_12084,N_14101);
xnor U15187 (N_15187,N_13857,N_12588);
xnor U15188 (N_15188,N_12259,N_13447);
nor U15189 (N_15189,N_13061,N_13840);
or U15190 (N_15190,N_11949,N_11412);
xnor U15191 (N_15191,N_14106,N_13830);
nor U15192 (N_15192,N_12174,N_14024);
and U15193 (N_15193,N_13049,N_10303);
nor U15194 (N_15194,N_11434,N_11057);
nor U15195 (N_15195,N_14263,N_10563);
or U15196 (N_15196,N_14051,N_14857);
or U15197 (N_15197,N_11303,N_10060);
nand U15198 (N_15198,N_12720,N_13308);
and U15199 (N_15199,N_11076,N_14781);
xnor U15200 (N_15200,N_13558,N_10785);
or U15201 (N_15201,N_12222,N_12424);
nand U15202 (N_15202,N_12391,N_11774);
nand U15203 (N_15203,N_12412,N_13812);
nor U15204 (N_15204,N_11318,N_12342);
or U15205 (N_15205,N_11725,N_14800);
nor U15206 (N_15206,N_14078,N_13596);
xnor U15207 (N_15207,N_11767,N_10447);
nand U15208 (N_15208,N_11590,N_10598);
xor U15209 (N_15209,N_13381,N_13288);
and U15210 (N_15210,N_10291,N_14139);
and U15211 (N_15211,N_10266,N_10371);
nand U15212 (N_15212,N_12477,N_11336);
and U15213 (N_15213,N_13928,N_14331);
xnor U15214 (N_15214,N_11850,N_12527);
nand U15215 (N_15215,N_11371,N_10015);
or U15216 (N_15216,N_10407,N_10993);
and U15217 (N_15217,N_14272,N_14275);
nand U15218 (N_15218,N_14321,N_12766);
or U15219 (N_15219,N_11569,N_11018);
and U15220 (N_15220,N_14869,N_10986);
xnor U15221 (N_15221,N_11115,N_10139);
or U15222 (N_15222,N_13395,N_10203);
nand U15223 (N_15223,N_12410,N_11698);
and U15224 (N_15224,N_11595,N_13671);
nor U15225 (N_15225,N_13607,N_10441);
or U15226 (N_15226,N_13404,N_12507);
or U15227 (N_15227,N_13362,N_10824);
nand U15228 (N_15228,N_12211,N_12121);
xnor U15229 (N_15229,N_10931,N_11328);
xnor U15230 (N_15230,N_12661,N_13642);
nor U15231 (N_15231,N_11879,N_10402);
and U15232 (N_15232,N_13746,N_11707);
nor U15233 (N_15233,N_14032,N_10592);
nand U15234 (N_15234,N_12255,N_13364);
nor U15235 (N_15235,N_10395,N_13032);
nor U15236 (N_15236,N_12695,N_11552);
nor U15237 (N_15237,N_10373,N_10743);
and U15238 (N_15238,N_10880,N_11281);
and U15239 (N_15239,N_13977,N_12337);
and U15240 (N_15240,N_13110,N_14141);
xnor U15241 (N_15241,N_10058,N_14584);
nor U15242 (N_15242,N_14144,N_14940);
and U15243 (N_15243,N_11951,N_12119);
xor U15244 (N_15244,N_14085,N_12913);
and U15245 (N_15245,N_14630,N_11748);
or U15246 (N_15246,N_10192,N_10666);
or U15247 (N_15247,N_11981,N_10603);
nand U15248 (N_15248,N_12508,N_14186);
xor U15249 (N_15249,N_14373,N_11155);
xor U15250 (N_15250,N_11687,N_14205);
xnor U15251 (N_15251,N_14963,N_10553);
or U15252 (N_15252,N_11749,N_10041);
and U15253 (N_15253,N_14597,N_13124);
nor U15254 (N_15254,N_11726,N_14933);
or U15255 (N_15255,N_14654,N_12971);
or U15256 (N_15256,N_10504,N_14596);
nand U15257 (N_15257,N_12564,N_13961);
nand U15258 (N_15258,N_14587,N_12897);
and U15259 (N_15259,N_13730,N_10011);
and U15260 (N_15260,N_11034,N_10908);
nand U15261 (N_15261,N_12196,N_10244);
nor U15262 (N_15262,N_11017,N_11557);
or U15263 (N_15263,N_11825,N_12677);
nor U15264 (N_15264,N_11697,N_10084);
and U15265 (N_15265,N_12002,N_10424);
and U15266 (N_15266,N_10815,N_14412);
or U15267 (N_15267,N_11614,N_10789);
xnor U15268 (N_15268,N_12671,N_12906);
xor U15269 (N_15269,N_13819,N_13628);
or U15270 (N_15270,N_13781,N_14312);
nand U15271 (N_15271,N_13185,N_11453);
or U15272 (N_15272,N_13326,N_13403);
or U15273 (N_15273,N_11461,N_12907);
and U15274 (N_15274,N_13556,N_10089);
nor U15275 (N_15275,N_10818,N_11704);
and U15276 (N_15276,N_14276,N_14501);
nor U15277 (N_15277,N_10388,N_12239);
nand U15278 (N_15278,N_11846,N_12954);
nand U15279 (N_15279,N_10198,N_14589);
and U15280 (N_15280,N_10633,N_13563);
nand U15281 (N_15281,N_10867,N_10252);
nor U15282 (N_15282,N_13945,N_11583);
and U15283 (N_15283,N_10056,N_10710);
and U15284 (N_15284,N_11108,N_10363);
nand U15285 (N_15285,N_13236,N_13256);
nor U15286 (N_15286,N_12585,N_13051);
xor U15287 (N_15287,N_12938,N_12519);
or U15288 (N_15288,N_11067,N_12855);
nand U15289 (N_15289,N_13794,N_12867);
xor U15290 (N_15290,N_12663,N_10063);
xnor U15291 (N_15291,N_12610,N_10655);
nor U15292 (N_15292,N_14478,N_10087);
or U15293 (N_15293,N_14196,N_12212);
nand U15294 (N_15294,N_14375,N_14052);
and U15295 (N_15295,N_11037,N_11676);
and U15296 (N_15296,N_11628,N_13354);
or U15297 (N_15297,N_12176,N_14209);
xnor U15298 (N_15298,N_12666,N_12806);
nor U15299 (N_15299,N_13925,N_12891);
nand U15300 (N_15300,N_11023,N_12371);
and U15301 (N_15301,N_14889,N_14649);
or U15302 (N_15302,N_11114,N_12698);
nor U15303 (N_15303,N_13983,N_10194);
nand U15304 (N_15304,N_12706,N_12177);
or U15305 (N_15305,N_10293,N_13578);
nand U15306 (N_15306,N_13294,N_13889);
xor U15307 (N_15307,N_12968,N_14667);
nor U15308 (N_15308,N_13631,N_14096);
nand U15309 (N_15309,N_10861,N_11528);
nor U15310 (N_15310,N_14819,N_13712);
or U15311 (N_15311,N_14685,N_10495);
and U15312 (N_15312,N_12750,N_10392);
nand U15313 (N_15313,N_11844,N_14417);
or U15314 (N_15314,N_11680,N_11624);
xnor U15315 (N_15315,N_12426,N_11548);
nand U15316 (N_15316,N_11225,N_12859);
nor U15317 (N_15317,N_11814,N_10680);
nand U15318 (N_15318,N_11181,N_12597);
xor U15319 (N_15319,N_13458,N_14945);
nor U15320 (N_15320,N_12873,N_14539);
or U15321 (N_15321,N_10800,N_11798);
xnor U15322 (N_15322,N_13552,N_13152);
xnor U15323 (N_15323,N_10183,N_14033);
nor U15324 (N_15324,N_11104,N_12852);
nand U15325 (N_15325,N_10966,N_13460);
nand U15326 (N_15326,N_10217,N_14962);
and U15327 (N_15327,N_12447,N_12417);
nand U15328 (N_15328,N_13621,N_10002);
or U15329 (N_15329,N_14999,N_14398);
nor U15330 (N_15330,N_14082,N_13973);
nor U15331 (N_15331,N_11255,N_13228);
and U15332 (N_15332,N_14924,N_13793);
nor U15333 (N_15333,N_11983,N_11745);
nor U15334 (N_15334,N_14524,N_13918);
and U15335 (N_15335,N_10488,N_13325);
nor U15336 (N_15336,N_11020,N_11918);
and U15337 (N_15337,N_14682,N_14562);
nor U15338 (N_15338,N_12935,N_14152);
nor U15339 (N_15339,N_11884,N_14200);
and U15340 (N_15340,N_12438,N_12643);
and U15341 (N_15341,N_14475,N_10439);
xor U15342 (N_15342,N_11470,N_14011);
xnor U15343 (N_15343,N_10485,N_12330);
nand U15344 (N_15344,N_12348,N_10930);
xnor U15345 (N_15345,N_12413,N_10956);
or U15346 (N_15346,N_11619,N_12814);
nor U15347 (N_15347,N_14606,N_10640);
or U15348 (N_15348,N_12601,N_12433);
xnor U15349 (N_15349,N_13987,N_11711);
or U15350 (N_15350,N_14592,N_11607);
nand U15351 (N_15351,N_13917,N_14750);
nor U15352 (N_15352,N_10847,N_14843);
or U15353 (N_15353,N_13620,N_10333);
or U15354 (N_15354,N_11664,N_10571);
or U15355 (N_15355,N_14703,N_11644);
and U15356 (N_15356,N_11764,N_14167);
or U15357 (N_15357,N_13969,N_12472);
nand U15358 (N_15358,N_13766,N_13290);
nor U15359 (N_15359,N_13449,N_10699);
and U15360 (N_15360,N_10994,N_13510);
xnor U15361 (N_15361,N_12983,N_11300);
nor U15362 (N_15362,N_11893,N_10250);
nand U15363 (N_15363,N_14639,N_10314);
or U15364 (N_15364,N_14493,N_11183);
xor U15365 (N_15365,N_12141,N_10325);
or U15366 (N_15366,N_13275,N_14916);
nand U15367 (N_15367,N_11510,N_10635);
nor U15368 (N_15368,N_12219,N_12995);
xnor U15369 (N_15369,N_11297,N_11625);
or U15370 (N_15370,N_11663,N_11642);
nand U15371 (N_15371,N_13891,N_10996);
or U15372 (N_15372,N_11695,N_12288);
xor U15373 (N_15373,N_13503,N_13747);
and U15374 (N_15374,N_14128,N_14971);
xor U15375 (N_15375,N_11330,N_13739);
nand U15376 (N_15376,N_13711,N_12635);
nand U15377 (N_15377,N_12058,N_13949);
xor U15378 (N_15378,N_13379,N_12045);
nand U15379 (N_15379,N_12403,N_14370);
or U15380 (N_15380,N_12461,N_14953);
nand U15381 (N_15381,N_11111,N_13959);
xor U15382 (N_15382,N_10806,N_10386);
or U15383 (N_15383,N_10362,N_11939);
nand U15384 (N_15384,N_11275,N_11103);
nand U15385 (N_15385,N_14519,N_11276);
nor U15386 (N_15386,N_14433,N_10367);
xor U15387 (N_15387,N_11238,N_13005);
xnor U15388 (N_15388,N_10646,N_14019);
nand U15389 (N_15389,N_12341,N_14241);
or U15390 (N_15390,N_10339,N_10416);
nor U15391 (N_15391,N_12460,N_14998);
and U15392 (N_15392,N_14731,N_11196);
or U15393 (N_15393,N_12310,N_10617);
xor U15394 (N_15394,N_14541,N_14428);
nor U15395 (N_15395,N_13516,N_14577);
and U15396 (N_15396,N_14449,N_10057);
nand U15397 (N_15397,N_12182,N_13813);
nand U15398 (N_15398,N_10974,N_10403);
nor U15399 (N_15399,N_11438,N_10619);
and U15400 (N_15400,N_14362,N_11826);
nor U15401 (N_15401,N_10828,N_14912);
and U15402 (N_15402,N_11776,N_14135);
or U15403 (N_15403,N_11611,N_14363);
nand U15404 (N_15404,N_10255,N_10809);
nor U15405 (N_15405,N_11616,N_14670);
xnor U15406 (N_15406,N_10644,N_10983);
and U15407 (N_15407,N_11481,N_13869);
nand U15408 (N_15408,N_10807,N_13215);
and U15409 (N_15409,N_14844,N_11659);
or U15410 (N_15410,N_14365,N_14013);
xnor U15411 (N_15411,N_11050,N_12686);
xor U15412 (N_15412,N_14970,N_13052);
or U15413 (N_15413,N_10421,N_13317);
and U15414 (N_15414,N_12493,N_13014);
nand U15415 (N_15415,N_11770,N_13077);
xnor U15416 (N_15416,N_13223,N_12503);
and U15417 (N_15417,N_14724,N_13811);
nand U15418 (N_15418,N_12618,N_11736);
nand U15419 (N_15419,N_12818,N_10896);
xnor U15420 (N_15420,N_11357,N_14304);
and U15421 (N_15421,N_14107,N_14394);
nand U15422 (N_15422,N_11237,N_14183);
xor U15423 (N_15423,N_13547,N_13496);
and U15424 (N_15424,N_10688,N_12052);
and U15425 (N_15425,N_11224,N_11402);
nor U15426 (N_15426,N_12145,N_13971);
or U15427 (N_15427,N_10205,N_12861);
xor U15428 (N_15428,N_13323,N_11771);
nand U15429 (N_15429,N_11380,N_14619);
or U15430 (N_15430,N_13226,N_11561);
or U15431 (N_15431,N_11420,N_14418);
nor U15432 (N_15432,N_13260,N_14638);
nand U15433 (N_15433,N_10559,N_13491);
or U15434 (N_15434,N_12151,N_10628);
nor U15435 (N_15435,N_11335,N_12027);
or U15436 (N_15436,N_10385,N_14406);
nor U15437 (N_15437,N_10538,N_13074);
xor U15438 (N_15438,N_13357,N_11033);
and U15439 (N_15439,N_10202,N_12860);
or U15440 (N_15440,N_14671,N_11922);
and U15441 (N_15441,N_11264,N_12969);
nor U15442 (N_15442,N_12580,N_14862);
or U15443 (N_15443,N_12827,N_14621);
nor U15444 (N_15444,N_14911,N_10687);
nand U15445 (N_15445,N_12172,N_12037);
nand U15446 (N_15446,N_12180,N_11973);
nor U15447 (N_15447,N_13687,N_10418);
xnor U15448 (N_15448,N_10595,N_13425);
nor U15449 (N_15449,N_12918,N_13219);
nand U15450 (N_15450,N_13542,N_11874);
and U15451 (N_15451,N_10112,N_11855);
and U15452 (N_15452,N_13314,N_14546);
nor U15453 (N_15453,N_13581,N_14663);
xor U15454 (N_15454,N_11991,N_14691);
and U15455 (N_15455,N_13285,N_12820);
or U15456 (N_15456,N_12425,N_12292);
nand U15457 (N_15457,N_11165,N_11559);
or U15458 (N_15458,N_13776,N_13967);
xnor U15459 (N_15459,N_12506,N_12070);
xnor U15460 (N_15460,N_13553,N_10004);
and U15461 (N_15461,N_10232,N_11282);
and U15462 (N_15462,N_12771,N_14341);
and U15463 (N_15463,N_12896,N_13016);
xor U15464 (N_15464,N_14774,N_13849);
and U15465 (N_15465,N_14993,N_12135);
nor U15466 (N_15466,N_12889,N_11424);
nor U15467 (N_15467,N_12134,N_13346);
or U15468 (N_15468,N_12912,N_13437);
nand U15469 (N_15469,N_11821,N_13393);
and U15470 (N_15470,N_11483,N_11920);
or U15471 (N_15471,N_12846,N_13420);
nor U15472 (N_15472,N_13768,N_13019);
xor U15473 (N_15473,N_11078,N_14219);
nand U15474 (N_15474,N_12946,N_10375);
or U15475 (N_15475,N_12615,N_10256);
nor U15476 (N_15476,N_13640,N_14435);
xnor U15477 (N_15477,N_14512,N_11604);
nand U15478 (N_15478,N_10415,N_14870);
or U15479 (N_15479,N_14823,N_11645);
or U15480 (N_15480,N_13380,N_12834);
nor U15481 (N_15481,N_14594,N_10988);
xor U15482 (N_15482,N_11164,N_11556);
or U15483 (N_15483,N_14111,N_11314);
or U15484 (N_15484,N_10870,N_10948);
nand U15485 (N_15485,N_10214,N_14628);
xnor U15486 (N_15486,N_12287,N_12687);
or U15487 (N_15487,N_12017,N_13755);
or U15488 (N_15488,N_10659,N_14874);
nor U15489 (N_15489,N_10282,N_14378);
xor U15490 (N_15490,N_13820,N_10304);
or U15491 (N_15491,N_12389,N_14784);
and U15492 (N_15492,N_12802,N_12073);
or U15493 (N_15493,N_11720,N_10156);
nor U15494 (N_15494,N_12046,N_13057);
or U15495 (N_15495,N_11700,N_13141);
or U15496 (N_15496,N_10759,N_10959);
xnor U15497 (N_15497,N_12289,N_13970);
nand U15498 (N_15498,N_11101,N_14029);
nor U15499 (N_15499,N_13907,N_11811);
nor U15500 (N_15500,N_10505,N_13184);
or U15501 (N_15501,N_14877,N_10267);
or U15502 (N_15502,N_11494,N_14009);
xnor U15503 (N_15503,N_13086,N_12800);
nor U15504 (N_15504,N_13650,N_13166);
nor U15505 (N_15505,N_11016,N_12584);
and U15506 (N_15506,N_14980,N_10061);
and U15507 (N_15507,N_10077,N_13044);
nand U15508 (N_15508,N_14496,N_14846);
and U15509 (N_15509,N_10927,N_11897);
xor U15510 (N_15510,N_14093,N_12483);
and U15511 (N_15511,N_13097,N_13706);
xnor U15512 (N_15512,N_14640,N_13790);
or U15513 (N_15513,N_13374,N_10940);
or U15514 (N_15514,N_12518,N_10511);
nor U15515 (N_15515,N_14668,N_11935);
or U15516 (N_15516,N_14212,N_11780);
nand U15517 (N_15517,N_12680,N_14776);
and U15518 (N_15518,N_11889,N_13344);
or U15519 (N_15519,N_14469,N_14875);
and U15520 (N_15520,N_11536,N_10379);
or U15521 (N_15521,N_12777,N_12263);
xor U15522 (N_15522,N_13451,N_11654);
nor U15523 (N_15523,N_12363,N_12238);
xor U15524 (N_15524,N_10290,N_11677);
nor U15525 (N_15525,N_11287,N_11866);
xnor U15526 (N_15526,N_13950,N_11252);
nor U15527 (N_15527,N_13733,N_11274);
and U15528 (N_15528,N_12092,N_14919);
or U15529 (N_15529,N_13067,N_11772);
and U15530 (N_15530,N_12197,N_12361);
or U15531 (N_15531,N_11191,N_12077);
or U15532 (N_15532,N_13641,N_14956);
or U15533 (N_15533,N_14377,N_14145);
nor U15534 (N_15534,N_13988,N_12679);
nand U15535 (N_15535,N_12010,N_11532);
nand U15536 (N_15536,N_12949,N_11222);
or U15537 (N_15537,N_11059,N_10279);
nand U15538 (N_15538,N_11601,N_11491);
and U15539 (N_15539,N_12243,N_10158);
nor U15540 (N_15540,N_10735,N_10074);
or U15541 (N_15541,N_10091,N_11570);
nor U15542 (N_15542,N_13302,N_11195);
xor U15543 (N_15543,N_11286,N_12103);
xnor U15544 (N_15544,N_11503,N_12542);
nor U15545 (N_15545,N_13784,N_14320);
or U15546 (N_15546,N_14837,N_11000);
xor U15547 (N_15547,N_11820,N_12051);
nand U15548 (N_15548,N_12991,N_14886);
nor U15549 (N_15549,N_12704,N_11597);
and U15550 (N_15550,N_10837,N_13131);
and U15551 (N_15551,N_14191,N_12162);
nand U15552 (N_15552,N_12474,N_13605);
nor U15553 (N_15553,N_11130,N_11212);
or U15554 (N_15554,N_11002,N_11221);
or U15555 (N_15555,N_14359,N_14388);
nand U15556 (N_15556,N_12025,N_12992);
xnor U15557 (N_15557,N_14876,N_12439);
xnor U15558 (N_15558,N_10457,N_13715);
xnor U15559 (N_15559,N_11395,N_13157);
or U15560 (N_15560,N_10776,N_12594);
xor U15561 (N_15561,N_13267,N_14441);
nor U15562 (N_15562,N_14251,N_12517);
xor U15563 (N_15563,N_14689,N_13532);
xnor U15564 (N_15564,N_11518,N_14404);
nor U15565 (N_15565,N_11834,N_14273);
and U15566 (N_15566,N_11670,N_12786);
xor U15567 (N_15567,N_12345,N_13705);
xnor U15568 (N_15568,N_12062,N_14070);
and U15569 (N_15569,N_12655,N_14299);
and U15570 (N_15570,N_11727,N_11440);
nor U15571 (N_15571,N_11848,N_11009);
and U15572 (N_15572,N_14353,N_14583);
or U15573 (N_15573,N_12996,N_13965);
xnor U15574 (N_15574,N_10247,N_10131);
nor U15575 (N_15575,N_11381,N_12563);
or U15576 (N_15576,N_11427,N_13149);
or U15577 (N_15577,N_13271,N_12898);
and U15578 (N_15578,N_12631,N_10187);
nor U15579 (N_15579,N_10005,N_12606);
or U15580 (N_15580,N_14931,N_12790);
and U15581 (N_15581,N_14470,N_14647);
nor U15582 (N_15582,N_10857,N_13888);
xnor U15583 (N_15583,N_12231,N_12252);
nand U15584 (N_15584,N_14437,N_12552);
xnor U15585 (N_15585,N_12902,N_10240);
and U15586 (N_15586,N_10967,N_13713);
and U15587 (N_15587,N_13808,N_11393);
and U15588 (N_15588,N_10564,N_13782);
nor U15589 (N_15589,N_13534,N_13893);
and U15590 (N_15590,N_14486,N_11250);
and U15591 (N_15591,N_11959,N_13111);
nand U15592 (N_15592,N_11269,N_11416);
or U15593 (N_15593,N_10763,N_14045);
or U15594 (N_15594,N_11647,N_14737);
and U15595 (N_15595,N_14678,N_14195);
xnor U15596 (N_15596,N_14792,N_11131);
nor U15597 (N_15597,N_12423,N_13011);
or U15598 (N_15598,N_11378,N_12957);
and U15599 (N_15599,N_14799,N_11126);
and U15600 (N_15600,N_13492,N_10287);
or U15601 (N_15601,N_11149,N_14785);
or U15602 (N_15602,N_12753,N_11053);
nor U15603 (N_15603,N_10981,N_14762);
and U15604 (N_15604,N_14559,N_13735);
nor U15605 (N_15605,N_12161,N_13197);
xnor U15606 (N_15606,N_13192,N_11849);
or U15607 (N_15607,N_11744,N_11558);
nand U15608 (N_15608,N_10229,N_13391);
and U15609 (N_15609,N_12920,N_10508);
nor U15610 (N_15610,N_13307,N_12384);
or U15611 (N_15611,N_14845,N_12942);
nand U15612 (N_15612,N_13428,N_13541);
nor U15613 (N_15613,N_12649,N_10315);
xor U15614 (N_15614,N_14458,N_13406);
and U15615 (N_15615,N_10631,N_13585);
xor U15616 (N_15616,N_13389,N_14807);
or U15617 (N_15617,N_12724,N_13001);
or U15618 (N_15618,N_13283,N_14560);
or U15619 (N_15619,N_12764,N_14250);
nand U15620 (N_15620,N_12240,N_12739);
nand U15621 (N_15621,N_12525,N_11243);
or U15622 (N_15622,N_13758,N_11313);
and U15623 (N_15623,N_13280,N_10346);
xnor U15624 (N_15624,N_10608,N_12273);
nand U15625 (N_15625,N_10579,N_14462);
xor U15626 (N_15626,N_11904,N_14965);
nor U15627 (N_15627,N_10045,N_11072);
and U15628 (N_15628,N_11626,N_13583);
xor U15629 (N_15629,N_10109,N_10258);
or U15630 (N_15630,N_10937,N_10612);
and U15631 (N_15631,N_10459,N_14509);
nand U15632 (N_15632,N_14355,N_11137);
and U15633 (N_15633,N_13539,N_11289);
xor U15634 (N_15634,N_12711,N_14232);
nor U15635 (N_15635,N_11010,N_11220);
xnor U15636 (N_15636,N_12851,N_10299);
xnor U15637 (N_15637,N_13194,N_12016);
xnor U15638 (N_15638,N_12574,N_10906);
nand U15639 (N_15639,N_12230,N_14892);
nand U15640 (N_15640,N_10228,N_11588);
nor U15641 (N_15641,N_10753,N_12798);
nand U15642 (N_15642,N_11379,N_12961);
nand U15643 (N_15643,N_13140,N_11474);
or U15644 (N_15644,N_12988,N_11102);
or U15645 (N_15645,N_10831,N_11334);
and U15646 (N_15646,N_11785,N_13176);
xor U15647 (N_15647,N_10895,N_11691);
or U15648 (N_15648,N_13088,N_12903);
and U15649 (N_15649,N_12179,N_14740);
nor U15650 (N_15650,N_13587,N_13944);
or U15651 (N_15651,N_11260,N_13257);
and U15652 (N_15652,N_11227,N_13931);
nand U15653 (N_15653,N_10035,N_11043);
or U15654 (N_15654,N_13293,N_10692);
xnor U15655 (N_15655,N_11817,N_12843);
and U15656 (N_15656,N_12297,N_14571);
nor U15657 (N_15657,N_10535,N_11809);
nor U15658 (N_15658,N_14847,N_14256);
nor U15659 (N_15659,N_12619,N_11305);
or U15660 (N_15660,N_12571,N_14783);
and U15661 (N_15661,N_13372,N_10193);
nand U15662 (N_15662,N_12778,N_13481);
xnor U15663 (N_15663,N_11279,N_13172);
nor U15664 (N_15664,N_12220,N_14815);
and U15665 (N_15665,N_13512,N_10611);
nor U15666 (N_15666,N_14696,N_12130);
nor U15667 (N_15667,N_12186,N_12106);
and U15668 (N_15668,N_14554,N_12950);
nor U15669 (N_15669,N_13957,N_11081);
or U15670 (N_15670,N_13439,N_11506);
xor U15671 (N_15671,N_11974,N_13356);
or U15672 (N_15672,N_10330,N_13292);
nand U15673 (N_15673,N_14573,N_10207);
or U15674 (N_15674,N_14641,N_13743);
and U15675 (N_15675,N_13181,N_11840);
nand U15676 (N_15676,N_11448,N_12888);
nand U15677 (N_15677,N_10584,N_13010);
nor U15678 (N_15678,N_13102,N_11549);
xor U15679 (N_15679,N_14248,N_12908);
nor U15680 (N_15680,N_13818,N_11019);
nand U15681 (N_15681,N_14210,N_10059);
nor U15682 (N_15682,N_10254,N_10149);
and U15683 (N_15683,N_14116,N_10737);
or U15684 (N_15684,N_11319,N_14281);
or U15685 (N_15685,N_14545,N_10230);
or U15686 (N_15686,N_12401,N_14599);
or U15687 (N_15687,N_12668,N_11618);
nand U15688 (N_15688,N_14984,N_12156);
nor U15689 (N_15689,N_13905,N_12065);
xor U15690 (N_15690,N_12762,N_14058);
or U15691 (N_15691,N_12776,N_10277);
nor U15692 (N_15692,N_10024,N_10411);
and U15693 (N_15693,N_11574,N_13203);
nand U15694 (N_15694,N_14508,N_11109);
xor U15695 (N_15695,N_10739,N_11655);
and U15696 (N_15696,N_14957,N_13366);
nand U15697 (N_15697,N_10810,N_12603);
nor U15698 (N_15698,N_14839,N_14616);
or U15699 (N_15699,N_13572,N_14286);
nand U15700 (N_15700,N_14658,N_14692);
and U15701 (N_15701,N_14787,N_11163);
nand U15702 (N_15702,N_12465,N_13985);
or U15703 (N_15703,N_13672,N_10917);
and U15704 (N_15704,N_11801,N_10297);
nor U15705 (N_15705,N_10349,N_12707);
and U15706 (N_15706,N_10756,N_12627);
and U15707 (N_15707,N_10813,N_12921);
nor U15708 (N_15708,N_14436,N_10577);
nor U15709 (N_15709,N_12286,N_12791);
nand U15710 (N_15710,N_11429,N_11882);
nand U15711 (N_15711,N_14927,N_10524);
nor U15712 (N_15712,N_10984,N_13807);
nand U15713 (N_15713,N_13360,N_10306);
and U15714 (N_15714,N_10055,N_10030);
nor U15715 (N_15715,N_10071,N_13213);
nand U15716 (N_15716,N_12757,N_14650);
and U15717 (N_15717,N_13703,N_14208);
xnor U15718 (N_15718,N_13932,N_11714);
nand U15719 (N_15719,N_11577,N_13021);
xnor U15720 (N_15720,N_14164,N_11462);
xnor U15721 (N_15721,N_12756,N_12142);
and U15722 (N_15722,N_11712,N_13029);
nand U15723 (N_15723,N_10947,N_12931);
xnor U15724 (N_15724,N_11630,N_13760);
nor U15725 (N_15725,N_11251,N_11580);
and U15726 (N_15726,N_12719,N_12158);
or U15727 (N_15727,N_10625,N_10814);
or U15728 (N_15728,N_14495,N_12458);
or U15729 (N_15729,N_14347,N_11071);
nand U15730 (N_15730,N_14561,N_14467);
xor U15731 (N_15731,N_12015,N_11993);
xnor U15732 (N_15732,N_13771,N_12194);
and U15733 (N_15733,N_14072,N_11863);
and U15734 (N_15734,N_10399,N_10483);
and U15735 (N_15735,N_12799,N_11021);
xnor U15736 (N_15736,N_10175,N_11873);
and U15737 (N_15737,N_11403,N_12041);
or U15738 (N_15738,N_13602,N_13643);
and U15739 (N_15739,N_14410,N_14095);
xor U15740 (N_15740,N_10090,N_10642);
nor U15741 (N_15741,N_14878,N_14409);
and U15742 (N_15742,N_14939,N_11366);
and U15743 (N_15743,N_10549,N_14105);
or U15744 (N_15744,N_13936,N_12359);
xor U15745 (N_15745,N_12842,N_13479);
and U15746 (N_15746,N_12788,N_13259);
or U15747 (N_15747,N_14812,N_13277);
and U15748 (N_15748,N_13661,N_13373);
nand U15749 (N_15749,N_13489,N_13146);
nand U15750 (N_15750,N_10168,N_12459);
or U15751 (N_15751,N_11288,N_11489);
or U15752 (N_15752,N_14483,N_13923);
nor U15753 (N_15753,N_14790,N_12492);
nand U15754 (N_15754,N_12296,N_13130);
and U15755 (N_15755,N_12055,N_11129);
and U15756 (N_15756,N_13615,N_14617);
and U15757 (N_15757,N_12748,N_14025);
xnor U15758 (N_15758,N_13644,N_10248);
xnor U15759 (N_15759,N_13958,N_11589);
or U15760 (N_15760,N_14788,N_14897);
xnor U15761 (N_15761,N_14659,N_14502);
and U15762 (N_15762,N_13846,N_13886);
nor U15763 (N_15763,N_14598,N_11970);
nor U15764 (N_15764,N_10741,N_13098);
nor U15765 (N_15765,N_10370,N_10241);
xnor U15766 (N_15766,N_13519,N_11348);
or U15767 (N_15767,N_10038,N_14187);
or U15768 (N_15768,N_12464,N_10629);
xor U15769 (N_15769,N_14684,N_13588);
nor U15770 (N_15770,N_13065,N_14610);
nor U15771 (N_15771,N_12315,N_12982);
nand U15772 (N_15772,N_10838,N_14552);
or U15773 (N_15773,N_13665,N_14131);
nand U15774 (N_15774,N_13142,N_14147);
xnor U15775 (N_15775,N_12350,N_11890);
and U15776 (N_15776,N_14871,N_10470);
and U15777 (N_15777,N_11858,N_12431);
nand U15778 (N_15778,N_13269,N_12937);
and U15779 (N_15779,N_10478,N_13402);
xnor U15780 (N_15780,N_12358,N_12225);
xnor U15781 (N_15781,N_13440,N_14543);
xnor U15782 (N_15782,N_11953,N_14637);
or U15783 (N_15783,N_10727,N_10271);
or U15784 (N_15784,N_14687,N_12874);
and U15785 (N_15785,N_14379,N_14907);
xor U15786 (N_15786,N_14683,N_14289);
xnor U15787 (N_15787,N_13649,N_10151);
nand U15788 (N_15788,N_10260,N_13879);
nand U15789 (N_15789,N_10869,N_14591);
nand U15790 (N_15790,N_11529,N_13463);
nor U15791 (N_15791,N_10316,N_11413);
and U15792 (N_15792,N_10844,N_13876);
xnor U15793 (N_15793,N_13848,N_12626);
nor U15794 (N_15794,N_11242,N_10997);
nor U15795 (N_15795,N_12554,N_11746);
nor U15796 (N_15796,N_13276,N_11509);
or U15797 (N_15797,N_14936,N_12882);
nand U15798 (N_15798,N_12269,N_10272);
nor U15799 (N_15799,N_11301,N_13080);
nand U15800 (N_15800,N_13386,N_13405);
or U15801 (N_15801,N_10493,N_14099);
and U15802 (N_15802,N_13694,N_11899);
nor U15803 (N_15803,N_14834,N_14608);
nand U15804 (N_15804,N_12608,N_10461);
nor U15805 (N_15805,N_11807,N_10977);
or U15806 (N_15806,N_11054,N_11715);
nand U15807 (N_15807,N_11777,N_11587);
xor U15808 (N_15808,N_13874,N_11660);
and U15809 (N_15809,N_13686,N_10671);
xnor U15810 (N_15810,N_14882,N_11594);
nand U15811 (N_15811,N_10872,N_11579);
and U15812 (N_15812,N_11716,N_10133);
xnor U15813 (N_15813,N_13199,N_13870);
nor U15814 (N_15814,N_14828,N_13984);
and U15815 (N_15815,N_10305,N_10408);
or U15816 (N_15816,N_13068,N_11432);
xnor U15817 (N_15817,N_14743,N_13234);
nor U15818 (N_15818,N_10920,N_11463);
nand U15819 (N_15819,N_14636,N_14556);
or U15820 (N_15820,N_10322,N_11169);
or U15821 (N_15821,N_13495,N_10173);
or U15822 (N_15822,N_12716,N_14672);
xnor U15823 (N_15823,N_10679,N_13630);
or U15824 (N_15824,N_13498,N_13000);
and U15825 (N_15825,N_10758,N_12980);
nand U15826 (N_15826,N_14430,N_14914);
nor U15827 (N_15827,N_10361,N_13894);
or U15828 (N_15828,N_12038,N_14036);
nand U15829 (N_15829,N_14213,N_12466);
nor U15830 (N_15830,N_10695,N_14407);
nor U15831 (N_15831,N_13873,N_10164);
and U15832 (N_15832,N_14380,N_14228);
and U15833 (N_15833,N_14117,N_14926);
nor U15834 (N_15834,N_14134,N_10668);
xor U15835 (N_15835,N_12986,N_10853);
xor U15836 (N_15836,N_11359,N_14569);
nor U15837 (N_15837,N_11442,N_13904);
nand U15838 (N_15838,N_12427,N_12976);
nand U15839 (N_15839,N_14959,N_11354);
and U15840 (N_15840,N_13205,N_11940);
nand U15841 (N_15841,N_13633,N_11263);
and U15842 (N_15842,N_10879,N_12640);
xor U15843 (N_15843,N_14061,N_14961);
and U15844 (N_15844,N_10476,N_13670);
nor U15845 (N_15845,N_11244,N_14118);
nor U15846 (N_15846,N_11806,N_13580);
or U15847 (N_15847,N_11272,N_14817);
nand U15848 (N_15848,N_14982,N_10166);
nand U15849 (N_15849,N_10462,N_12265);
and U15850 (N_15850,N_14290,N_13487);
nand U15851 (N_15851,N_11585,N_10049);
xnor U15852 (N_15852,N_14252,N_12114);
nor U15853 (N_15853,N_10817,N_12555);
and U15854 (N_15854,N_13864,N_12781);
nor U15855 (N_15855,N_13397,N_11353);
or U15856 (N_15856,N_13244,N_12648);
xnor U15857 (N_15857,N_10075,N_14613);
nor U15858 (N_15858,N_13454,N_14827);
xor U15859 (N_15859,N_10661,N_10430);
xor U15860 (N_15860,N_10958,N_14570);
xnor U15861 (N_15861,N_13196,N_14607);
nand U15862 (N_15862,N_14310,N_14126);
xnor U15863 (N_15863,N_10179,N_14727);
xnor U15864 (N_15864,N_10884,N_12729);
and U15865 (N_15865,N_10894,N_11478);
xor U15866 (N_15866,N_10269,N_13589);
nand U15867 (N_15867,N_12381,N_11804);
and U15868 (N_15868,N_11485,N_13953);
nor U15869 (N_15869,N_12013,N_14977);
and U15870 (N_15870,N_12349,N_10404);
xnor U15871 (N_15871,N_10526,N_12303);
nor U15872 (N_15872,N_12462,N_12515);
xor U15873 (N_15873,N_10552,N_10106);
nor U15874 (N_15874,N_14679,N_14995);
or U15875 (N_15875,N_14611,N_14972);
xor U15876 (N_15876,N_14255,N_10380);
or U15877 (N_15877,N_13384,N_12964);
nand U15878 (N_15878,N_14510,N_14459);
nand U15879 (N_15879,N_13571,N_10468);
or U15880 (N_15880,N_13270,N_14329);
nand U15881 (N_15881,N_11584,N_12737);
xor U15882 (N_15882,N_13474,N_13003);
or U15883 (N_15883,N_11791,N_14764);
and U15884 (N_15884,N_12100,N_11198);
xor U15885 (N_15885,N_11271,N_13568);
nand U15886 (N_15886,N_10593,N_10064);
nor U15887 (N_15887,N_10963,N_11219);
and U15888 (N_15888,N_11352,N_14309);
nand U15889 (N_15889,N_14421,N_13348);
nand U15890 (N_15890,N_12241,N_11069);
and U15891 (N_15891,N_11246,N_11835);
nor U15892 (N_15892,N_10523,N_11332);
nand U15893 (N_15893,N_11231,N_10188);
or U15894 (N_15894,N_14754,N_12810);
nor U15895 (N_15895,N_12352,N_14274);
nor U15896 (N_15896,N_12333,N_12808);
or U15897 (N_15897,N_14590,N_13898);
xnor U15898 (N_15898,N_14160,N_11280);
xor U15899 (N_15899,N_12409,N_12546);
nand U15900 (N_15900,N_13311,N_13043);
or U15901 (N_15901,N_10410,N_13375);
xnor U15902 (N_15902,N_10979,N_13304);
xnor U15903 (N_15903,N_10137,N_14660);
nor U15904 (N_15904,N_13321,N_12646);
or U15905 (N_15905,N_11754,N_14487);
nor U15906 (N_15906,N_14133,N_12690);
or U15907 (N_15907,N_14801,N_11267);
nor U15908 (N_15908,N_10775,N_10171);
xor U15909 (N_15909,N_11460,N_11458);
nor U15910 (N_15910,N_11960,N_14517);
or U15911 (N_15911,N_14461,N_10167);
and U15912 (N_15912,N_11439,N_14777);
or U15913 (N_15913,N_10893,N_10390);
and U15914 (N_15914,N_10718,N_12871);
nand U15915 (N_15915,N_14076,N_13858);
or U15916 (N_15916,N_10700,N_10442);
nor U15917 (N_15917,N_11789,N_13107);
and U15918 (N_15918,N_11862,N_11477);
and U15919 (N_15919,N_12633,N_11741);
and U15920 (N_15920,N_13177,N_11768);
nor U15921 (N_15921,N_12693,N_14217);
nand U15922 (N_15922,N_13443,N_11234);
and U15923 (N_15923,N_13822,N_14527);
nand U15924 (N_15924,N_11156,N_13531);
and U15925 (N_15925,N_13121,N_14021);
or U15926 (N_15926,N_12267,N_12069);
and U15927 (N_15927,N_10622,N_10046);
and U15928 (N_15928,N_14680,N_10583);
and U15929 (N_15929,N_14722,N_13901);
or U15930 (N_15930,N_12327,N_13218);
nor U15931 (N_15931,N_14426,N_13333);
xor U15932 (N_15932,N_13725,N_12708);
or U15933 (N_15933,N_12063,N_12792);
or U15934 (N_15934,N_12308,N_11475);
xor U15935 (N_15935,N_11120,N_10618);
nand U15936 (N_15936,N_11467,N_10420);
and U15937 (N_15937,N_11218,N_11638);
or U15938 (N_15938,N_11705,N_14600);
or U15939 (N_15939,N_13690,N_10799);
nor U15940 (N_15940,N_12281,N_10876);
and U15941 (N_15941,N_10698,N_11599);
xnor U15942 (N_15942,N_10405,N_10652);
nand U15943 (N_15943,N_11740,N_14444);
or U15944 (N_15944,N_11365,N_14464);
nand U15945 (N_15945,N_13761,N_10709);
xor U15946 (N_15946,N_10039,N_10597);
nand U15947 (N_15947,N_14922,N_12978);
or U15948 (N_15948,N_10261,N_10567);
nand U15949 (N_15949,N_11830,N_13956);
nand U15950 (N_15950,N_10850,N_10547);
nand U15951 (N_15951,N_13084,N_13897);
or U15952 (N_15952,N_10712,N_11087);
or U15953 (N_15953,N_10599,N_12207);
nand U15954 (N_15954,N_11887,N_14075);
and U15955 (N_15955,N_11933,N_10043);
and U15956 (N_15956,N_13033,N_12206);
nor U15957 (N_15957,N_11684,N_10531);
or U15958 (N_15958,N_12828,N_12494);
or U15959 (N_15959,N_10760,N_14108);
nand U15960 (N_15960,N_14482,N_10443);
nor U15961 (N_15961,N_10270,N_13533);
or U15962 (N_15962,N_11154,N_10051);
xor U15963 (N_15963,N_10406,N_11916);
nand U15964 (N_15964,N_14655,N_12535);
and U15965 (N_15965,N_10916,N_14485);
and U15966 (N_15966,N_12332,N_12490);
nand U15967 (N_15967,N_13736,N_14749);
and U15968 (N_15968,N_11351,N_14393);
or U15969 (N_15969,N_10653,N_14516);
nand U15970 (N_15970,N_12478,N_13683);
xnor U15971 (N_15971,N_11653,N_14376);
nor U15972 (N_15972,N_11581,N_10474);
xnor U15973 (N_15973,N_14346,N_12549);
xor U15974 (N_15974,N_11089,N_13841);
nand U15975 (N_15975,N_14746,N_11763);
and U15976 (N_15976,N_12133,N_13318);
or U15977 (N_15977,N_12396,N_10440);
xor U15978 (N_15978,N_10342,N_13573);
or U15979 (N_15979,N_13594,N_10053);
or U15980 (N_15980,N_11138,N_10515);
and U15981 (N_15981,N_10394,N_14012);
or U15982 (N_15982,N_10724,N_10849);
nor U15983 (N_15983,N_14307,N_14935);
nor U15984 (N_15984,N_13843,N_11028);
or U15985 (N_15985,N_12159,N_12074);
xnor U15986 (N_15986,N_13127,N_10144);
nand U15987 (N_15987,N_11385,N_11333);
xor U15988 (N_15988,N_10129,N_10110);
and U15989 (N_15989,N_10337,N_11182);
or U15990 (N_15990,N_11859,N_14718);
xnor U15991 (N_15991,N_11472,N_12387);
nand U15992 (N_15992,N_12972,N_12981);
and U15993 (N_15993,N_11637,N_12632);
and U15994 (N_15994,N_13383,N_14941);
and U15995 (N_15995,N_10525,N_12300);
nor U15996 (N_15996,N_14456,N_12355);
and U15997 (N_15997,N_14908,N_13499);
nor U15998 (N_15998,N_13770,N_11501);
nor U15999 (N_15999,N_10381,N_13610);
xor U16000 (N_16000,N_12374,N_11007);
nand U16001 (N_16001,N_10285,N_13839);
nand U16002 (N_16002,N_12021,N_13966);
nand U16003 (N_16003,N_10794,N_11493);
nor U16004 (N_16004,N_14371,N_13688);
and U16005 (N_16005,N_14511,N_13501);
nand U16006 (N_16006,N_14382,N_10209);
or U16007 (N_16007,N_12489,N_14681);
and U16008 (N_16008,N_10866,N_13312);
or U16009 (N_16009,N_12139,N_12674);
xnor U16010 (N_16010,N_10662,N_11958);
nor U16011 (N_16011,N_11185,N_11482);
xnor U16012 (N_16012,N_12388,N_12028);
nand U16013 (N_16013,N_12862,N_14451);
and U16014 (N_16014,N_13732,N_11646);
and U16015 (N_16015,N_11990,N_14896);
xor U16016 (N_16016,N_11110,N_11502);
nor U16017 (N_16017,N_14284,N_12155);
nor U16018 (N_16018,N_14405,N_13438);
and U16019 (N_16019,N_11228,N_11546);
xor U16020 (N_16020,N_11988,N_14016);
nand U16021 (N_16021,N_10236,N_14368);
nand U16022 (N_16022,N_13566,N_10280);
or U16023 (N_16023,N_10037,N_11175);
nor U16024 (N_16024,N_14288,N_12833);
xor U16025 (N_16025,N_12900,N_13225);
nand U16026 (N_16026,N_14214,N_11784);
or U16027 (N_16027,N_13227,N_11883);
or U16028 (N_16028,N_13845,N_13787);
and U16029 (N_16029,N_11408,N_13716);
xnor U16030 (N_16030,N_10082,N_10487);
and U16031 (N_16031,N_12850,N_11425);
and U16032 (N_16032,N_12963,N_11046);
or U16033 (N_16033,N_14973,N_11063);
nor U16034 (N_16034,N_10308,N_14580);
nor U16035 (N_16035,N_10676,N_13803);
nor U16036 (N_16036,N_13062,N_11957);
or U16037 (N_16037,N_12917,N_10591);
nand U16038 (N_16038,N_11900,N_12967);
xor U16039 (N_16039,N_14073,N_13656);
xor U16040 (N_16040,N_10023,N_13880);
xnor U16041 (N_16041,N_12364,N_11298);
and U16042 (N_16042,N_14431,N_10494);
and U16043 (N_16043,N_10897,N_13597);
nor U16044 (N_16044,N_11146,N_14262);
nor U16045 (N_16045,N_12817,N_11934);
nor U16046 (N_16046,N_14748,N_10761);
or U16047 (N_16047,N_13470,N_10919);
or U16048 (N_16048,N_13128,N_13968);
xor U16049 (N_16049,N_13429,N_14761);
and U16050 (N_16050,N_14989,N_10336);
nor U16051 (N_16051,N_13101,N_11189);
or U16052 (N_16052,N_12970,N_10120);
nand U16053 (N_16053,N_12595,N_11823);
xor U16054 (N_16054,N_14489,N_12744);
and U16055 (N_16055,N_14542,N_10123);
xor U16056 (N_16056,N_12624,N_14233);
nor U16057 (N_16057,N_12112,N_12299);
xnor U16058 (N_16058,N_14526,N_10821);
nor U16059 (N_16059,N_11919,N_12759);
or U16060 (N_16060,N_12941,N_14521);
nand U16061 (N_16061,N_10784,N_11151);
xor U16062 (N_16062,N_12302,N_10068);
nor U16063 (N_16063,N_11370,N_14605);
and U16064 (N_16064,N_12395,N_14189);
xor U16065 (N_16065,N_12313,N_10517);
nand U16066 (N_16066,N_12115,N_10779);
or U16067 (N_16067,N_11141,N_14402);
xnor U16068 (N_16068,N_12520,N_11391);
and U16069 (N_16069,N_13779,N_13895);
xnor U16070 (N_16070,N_10738,N_14121);
or U16071 (N_16071,N_11479,N_12958);
nor U16072 (N_16072,N_12301,N_14349);
nand U16073 (N_16073,N_14300,N_14389);
nor U16074 (N_16074,N_14071,N_12488);
nand U16075 (N_16075,N_11652,N_10576);
xor U16076 (N_16076,N_14419,N_12188);
xnor U16077 (N_16077,N_11531,N_13232);
and U16078 (N_16078,N_13992,N_10031);
and U16079 (N_16079,N_11230,N_12794);
or U16080 (N_16080,N_13993,N_13159);
nor U16081 (N_16081,N_12268,N_10519);
nor U16082 (N_16082,N_10596,N_14803);
xnor U16083 (N_16083,N_12872,N_10726);
and U16084 (N_16084,N_12064,N_13334);
xnor U16085 (N_16085,N_14909,N_11788);
nor U16086 (N_16086,N_11793,N_10086);
or U16087 (N_16087,N_11187,N_12547);
xnor U16088 (N_16088,N_12717,N_10001);
or U16089 (N_16089,N_14062,N_10274);
nand U16090 (N_16090,N_13306,N_11377);
and U16091 (N_16091,N_11527,N_12398);
or U16092 (N_16092,N_13448,N_12026);
xor U16093 (N_16093,N_12625,N_11567);
nor U16094 (N_16094,N_11397,N_11610);
and U16095 (N_16095,N_12249,N_13263);
nor U16096 (N_16096,N_13167,N_13986);
nand U16097 (N_16097,N_14893,N_10899);
and U16098 (N_16098,N_12540,N_14699);
nand U16099 (N_16099,N_13638,N_12170);
nor U16100 (N_16100,N_13409,N_11615);
nand U16101 (N_16101,N_12475,N_10437);
nor U16102 (N_16102,N_13295,N_14125);
nor U16103 (N_16103,N_10298,N_11537);
nand U16104 (N_16104,N_11851,N_11085);
nand U16105 (N_16105,N_12714,N_12675);
nor U16106 (N_16106,N_14579,N_10132);
and U16107 (N_16107,N_10533,N_11112);
nor U16108 (N_16108,N_10197,N_12316);
nor U16109 (N_16109,N_12353,N_13369);
or U16110 (N_16110,N_12372,N_10259);
and U16111 (N_16111,N_11719,N_12164);
xor U16112 (N_16112,N_10883,N_12404);
xor U16113 (N_16113,N_14522,N_14983);
or U16114 (N_16114,N_12169,N_10711);
xnor U16115 (N_16115,N_12819,N_13093);
nor U16116 (N_16116,N_10951,N_12665);
xor U16117 (N_16117,N_11199,N_14423);
nor U16118 (N_16118,N_14574,N_11547);
and U16119 (N_16119,N_12048,N_12233);
nor U16120 (N_16120,N_10764,N_11235);
nand U16121 (N_16121,N_13550,N_10026);
xor U16122 (N_16122,N_11127,N_12463);
or U16123 (N_16123,N_13297,N_14741);
and U16124 (N_16124,N_13261,N_12000);
and U16125 (N_16125,N_12804,N_14136);
and U16126 (N_16126,N_14414,N_10052);
nand U16127 (N_16127,N_13560,N_10972);
or U16128 (N_16128,N_13833,N_10887);
and U16129 (N_16129,N_13139,N_13071);
nand U16130 (N_16130,N_13731,N_10450);
or U16131 (N_16131,N_13180,N_10569);
nor U16132 (N_16132,N_13774,N_13193);
xnor U16133 (N_16133,N_14159,N_13548);
xnor U16134 (N_16134,N_13300,N_11049);
and U16135 (N_16135,N_13681,N_14841);
nor U16136 (N_16136,N_10099,N_12848);
and U16137 (N_16137,N_11456,N_11775);
nand U16138 (N_16138,N_12405,N_10530);
or U16139 (N_16139,N_11722,N_12831);
nor U16140 (N_16140,N_14805,N_13981);
and U16141 (N_16141,N_13695,N_13305);
or U16142 (N_16142,N_12007,N_12559);
or U16143 (N_16143,N_10970,N_11430);
nand U16144 (N_16144,N_13798,N_14083);
xor U16145 (N_16145,N_14756,N_14775);
or U16146 (N_16146,N_10985,N_10127);
nor U16147 (N_16147,N_12386,N_11982);
nor U16148 (N_16148,N_11052,N_13942);
nand U16149 (N_16149,N_12192,N_11902);
xnor U16150 (N_16150,N_10073,N_13785);
nor U16151 (N_16151,N_12271,N_12732);
xor U16152 (N_16152,N_13821,N_12008);
nor U16153 (N_16153,N_10121,N_13345);
and U16154 (N_16154,N_12556,N_13727);
xor U16155 (N_16155,N_10939,N_10962);
nand U16156 (N_16156,N_11291,N_10539);
nand U16157 (N_16157,N_14829,N_14988);
xnor U16158 (N_16158,N_10196,N_14981);
nand U16159 (N_16159,N_11968,N_14318);
and U16160 (N_16160,N_13835,N_11320);
or U16161 (N_16161,N_11766,N_10143);
and U16162 (N_16162,N_10928,N_10943);
nand U16163 (N_16163,N_10320,N_14162);
xnor U16164 (N_16164,N_13230,N_10798);
xor U16165 (N_16165,N_10521,N_10231);
nor U16166 (N_16166,N_11376,N_14002);
nand U16167 (N_16167,N_11436,N_10636);
or U16168 (N_16168,N_10148,N_12779);
nor U16169 (N_16169,N_13209,N_11465);
nand U16170 (N_16170,N_11133,N_14712);
or U16171 (N_16171,N_14400,N_10615);
or U16172 (N_16172,N_11987,N_13377);
xnor U16173 (N_16173,N_12125,N_12437);
xor U16174 (N_16174,N_14930,N_12435);
or U16175 (N_16175,N_10343,N_14330);
and U16176 (N_16176,N_13229,N_11349);
and U16177 (N_16177,N_14020,N_10383);
or U16178 (N_16178,N_14976,N_12399);
nor U16179 (N_16179,N_14015,N_10728);
and U16180 (N_16180,N_11202,N_12999);
xnor U16181 (N_16181,N_14325,N_12513);
xnor U16182 (N_16182,N_10990,N_13551);
nor U16183 (N_16183,N_11285,N_10871);
xnor U16184 (N_16184,N_10545,N_10160);
xor U16185 (N_16185,N_12132,N_12692);
or U16186 (N_16186,N_14237,N_13814);
nand U16187 (N_16187,N_14367,N_11294);
or U16188 (N_16188,N_10725,N_11520);
nor U16189 (N_16189,N_13791,N_12081);
xnor U16190 (N_16190,N_14974,N_12278);
nor U16191 (N_16191,N_11881,N_14150);
nor U16192 (N_16192,N_13767,N_12043);
xor U16193 (N_16193,N_13991,N_14460);
nor U16194 (N_16194,N_12524,N_10412);
nand U16195 (N_16195,N_10456,N_10875);
and U16196 (N_16196,N_13002,N_11315);
xor U16197 (N_16197,N_13445,N_11696);
and U16198 (N_16198,N_12940,N_12004);
xor U16199 (N_16199,N_11382,N_14767);
and U16200 (N_16200,N_10312,N_12126);
nand U16201 (N_16201,N_13696,N_14216);
or U16202 (N_16202,N_12450,N_11941);
nand U16203 (N_16203,N_10580,N_11679);
xnor U16204 (N_16204,N_10968,N_10528);
nor U16205 (N_16205,N_14153,N_10169);
or U16206 (N_16206,N_10094,N_11639);
nand U16207 (N_16207,N_13376,N_14005);
and U16208 (N_16208,N_12276,N_11686);
and U16209 (N_16209,N_12275,N_13653);
nand U16210 (N_16210,N_11490,N_13919);
or U16211 (N_16211,N_12548,N_13544);
and U16212 (N_16212,N_10098,N_11511);
or U16213 (N_16213,N_11066,N_10136);
nand U16214 (N_16214,N_12932,N_13371);
nor U16215 (N_16215,N_13635,N_10097);
or U16216 (N_16216,N_12380,N_11540);
xnor U16217 (N_16217,N_10783,N_12319);
nand U16218 (N_16218,N_11406,N_13116);
or U16219 (N_16219,N_13309,N_13039);
nand U16220 (N_16220,N_11535,N_10472);
xnor U16221 (N_16221,N_11113,N_11572);
or U16222 (N_16222,N_11488,N_12651);
or U16223 (N_16223,N_12356,N_10162);
and U16224 (N_16224,N_12858,N_12003);
or U16225 (N_16225,N_13217,N_11640);
and U16226 (N_16226,N_14717,N_11454);
or U16227 (N_16227,N_11925,N_13444);
nand U16228 (N_16228,N_10107,N_12928);
nand U16229 (N_16229,N_12590,N_12277);
nand U16230 (N_16230,N_10289,N_12050);
and U16231 (N_16231,N_12733,N_14239);
or U16232 (N_16232,N_10145,N_13046);
nand U16233 (N_16233,N_14301,N_10557);
nand U16234 (N_16234,N_13135,N_11369);
nand U16235 (N_16235,N_14383,N_13220);
nor U16236 (N_16236,N_14697,N_10354);
and U16237 (N_16237,N_10224,N_14042);
nor U16238 (N_16238,N_13545,N_10338);
nor U16239 (N_16239,N_13488,N_14403);
or U16240 (N_16240,N_13350,N_11143);
and U16241 (N_16241,N_10154,N_12682);
or U16242 (N_16242,N_11045,N_10703);
or U16243 (N_16243,N_10781,N_13645);
xor U16244 (N_16244,N_14060,N_14343);
or U16245 (N_16245,N_10945,N_11522);
nand U16246 (N_16246,N_13948,N_10675);
xnor U16247 (N_16247,N_10276,N_10734);
nor U16248 (N_16248,N_14246,N_13151);
or U16249 (N_16249,N_12541,N_12244);
nor U16250 (N_16250,N_11012,N_14796);
and U16251 (N_16251,N_11965,N_13600);
nand U16252 (N_16252,N_11273,N_10892);
nor U16253 (N_16253,N_14381,N_12153);
or U16254 (N_16254,N_13999,N_12098);
or U16255 (N_16255,N_14602,N_14578);
nand U16256 (N_16256,N_13549,N_14694);
nor U16257 (N_16257,N_11950,N_13710);
xor U16258 (N_16258,N_12080,N_10740);
and U16259 (N_16259,N_13279,N_13885);
and U16260 (N_16260,N_13358,N_11419);
nor U16261 (N_16261,N_13521,N_11689);
nor U16262 (N_16262,N_12516,N_10932);
and U16263 (N_16263,N_14657,N_13637);
xnor U16264 (N_16264,N_11400,N_14833);
nor U16265 (N_16265,N_13722,N_13245);
or U16266 (N_16266,N_13530,N_11596);
xnor U16267 (N_16267,N_10832,N_13466);
nand U16268 (N_16268,N_13680,N_10473);
or U16269 (N_16269,N_13797,N_11759);
nor U16270 (N_16270,N_12024,N_11732);
xor U16271 (N_16271,N_11634,N_12534);
xor U16272 (N_16272,N_13543,N_10575);
xor U16273 (N_16273,N_12205,N_14707);
nor U16274 (N_16274,N_14634,N_10497);
xnor U16275 (N_16275,N_13890,N_11692);
nand U16276 (N_16276,N_10924,N_13118);
and U16277 (N_16277,N_14261,N_12774);
nor U16278 (N_16278,N_11880,N_12109);
or U16279 (N_16279,N_12532,N_11118);
nand U16280 (N_16280,N_11822,N_13692);
or U16281 (N_16281,N_14564,N_10649);
or U16282 (N_16282,N_11152,N_13201);
nor U16283 (N_16283,N_14119,N_12087);
nand U16284 (N_16284,N_14514,N_11913);
nand U16285 (N_16285,N_11672,N_10042);
nor U16286 (N_16286,N_11048,N_10935);
and U16287 (N_16287,N_14260,N_11885);
nor U16288 (N_16288,N_10300,N_10694);
or U16289 (N_16289,N_12228,N_13025);
or U16290 (N_16290,N_10656,N_10353);
nor U16291 (N_16291,N_13616,N_13978);
nor U16292 (N_16292,N_13332,N_12683);
or U16293 (N_16293,N_13960,N_10980);
nand U16294 (N_16294,N_11469,N_11967);
and U16295 (N_16295,N_12673,N_12647);
and U16296 (N_16296,N_11507,N_14934);
or U16297 (N_16297,N_11752,N_13728);
nor U16298 (N_16298,N_14185,N_10957);
nand U16299 (N_16299,N_11853,N_12237);
xor U16300 (N_16300,N_14690,N_14089);
nand U16301 (N_16301,N_11254,N_14612);
xor U16302 (N_16302,N_11060,N_12936);
or U16303 (N_16303,N_10054,N_13868);
or U16304 (N_16304,N_12154,N_10859);
or U16305 (N_16305,N_13399,N_10686);
nor U16306 (N_16306,N_13036,N_13198);
xnor U16307 (N_16307,N_11808,N_11343);
xnor U16308 (N_16308,N_14317,N_12029);
nand U16309 (N_16309,N_11144,N_13896);
nand U16310 (N_16310,N_12501,N_13660);
or U16311 (N_16311,N_10754,N_13913);
and U16312 (N_16312,N_11265,N_11364);
nand U16313 (N_16313,N_11781,N_14158);
xnor U16314 (N_16314,N_10902,N_12336);
nand U16315 (N_16315,N_10391,N_13914);
xnor U16316 (N_16316,N_13007,N_12669);
or U16317 (N_16317,N_10973,N_13939);
xor U16318 (N_16318,N_11912,N_10331);
nor U16319 (N_16319,N_12977,N_12393);
nor U16320 (N_16320,N_11495,N_13729);
or U16321 (N_16321,N_14921,N_11106);
nand U16322 (N_16322,N_12293,N_12840);
nor U16323 (N_16323,N_10544,N_14868);
xnor U16324 (N_16324,N_14997,N_11457);
and U16325 (N_16325,N_14397,N_14477);
nand U16326 (N_16326,N_12826,N_11906);
or U16327 (N_16327,N_10681,N_11008);
or U16328 (N_16328,N_12242,N_13085);
and U16329 (N_16329,N_13513,N_14832);
and U16330 (N_16330,N_10296,N_13717);
xor U16331 (N_16331,N_10246,N_12845);
nand U16332 (N_16332,N_14455,N_11710);
and U16333 (N_16333,N_13989,N_13457);
and U16334 (N_16334,N_12613,N_11875);
nand U16335 (N_16335,N_11466,N_10995);
and U16336 (N_16336,N_11139,N_12198);
and U16337 (N_16337,N_10795,N_13757);
nor U16338 (N_16338,N_11980,N_13253);
xor U16339 (N_16339,N_11092,N_11088);
nand U16340 (N_16340,N_14917,N_12522);
nand U16341 (N_16341,N_10529,N_10614);
nand U16342 (N_16342,N_13699,N_13401);
and U16343 (N_16343,N_13570,N_11292);
and U16344 (N_16344,N_11932,N_14401);
and U16345 (N_16345,N_12120,N_14296);
and U16346 (N_16346,N_10542,N_12944);
nand U16347 (N_16347,N_13937,N_14282);
xnor U16348 (N_16348,N_13806,N_11153);
nor U16349 (N_16349,N_13693,N_11843);
nor U16350 (N_16350,N_10400,N_12083);
and U16351 (N_16351,N_11923,N_12645);
and U16352 (N_16352,N_14698,N_13476);
or U16353 (N_16353,N_11188,N_10122);
nor U16354 (N_16354,N_14808,N_12740);
or U16355 (N_16355,N_11193,N_14215);
nand U16356 (N_16356,N_13020,N_13082);
xor U16357 (N_16357,N_12113,N_11864);
or U16358 (N_16358,N_11387,N_13851);
and U16359 (N_16359,N_10114,N_10434);
nor U16360 (N_16360,N_11955,N_12001);
and U16361 (N_16361,N_12101,N_14326);
nor U16362 (N_16362,N_14850,N_14759);
nor U16363 (N_16363,N_13915,N_14948);
nor U16364 (N_16364,N_12059,N_11892);
and U16365 (N_16365,N_14166,N_11373);
and U16366 (N_16366,N_13143,N_11657);
or U16367 (N_16367,N_12746,N_13446);
nand U16368 (N_16368,N_12599,N_13483);
nand U16369 (N_16369,N_12075,N_10397);
or U16370 (N_16370,N_14197,N_13281);
or U16371 (N_16371,N_13947,N_14504);
and U16372 (N_16372,N_13450,N_11857);
and U16373 (N_16373,N_14450,N_13769);
or U16374 (N_16374,N_11617,N_13627);
xor U16375 (N_16375,N_11339,N_13617);
xor U16376 (N_16376,N_10626,N_14066);
nor U16377 (N_16377,N_12927,N_14757);
nor U16378 (N_16378,N_14726,N_11787);
nand U16379 (N_16379,N_13674,N_10914);
nand U16380 (N_16380,N_12569,N_13860);
nand U16381 (N_16381,N_13247,N_13619);
nand U16382 (N_16382,N_11476,N_10190);
or U16383 (N_16383,N_11799,N_14646);
nand U16384 (N_16384,N_10889,N_12226);
or U16385 (N_16385,N_12586,N_10118);
xnor U16386 (N_16386,N_14873,N_11179);
or U16387 (N_16387,N_12210,N_13456);
nand U16388 (N_16388,N_11132,N_10801);
or U16389 (N_16389,N_14446,N_13210);
nand U16390 (N_16390,N_14038,N_12952);
or U16391 (N_16391,N_13604,N_11203);
or U16392 (N_16392,N_10660,N_12630);
nand U16393 (N_16393,N_13595,N_14298);
and U16394 (N_16394,N_14360,N_11383);
or U16395 (N_16395,N_14558,N_13390);
and U16396 (N_16396,N_11927,N_12803);
or U16397 (N_16397,N_11782,N_10101);
and U16398 (N_16398,N_10820,N_11091);
xnor U16399 (N_16399,N_12730,N_13935);
nand U16400 (N_16400,N_14172,N_11984);
nand U16401 (N_16401,N_13611,N_11166);
or U16402 (N_16402,N_14127,N_14069);
nand U16403 (N_16403,N_10991,N_12919);
and U16404 (N_16404,N_10693,N_10105);
nor U16405 (N_16405,N_10585,N_13714);
and U16406 (N_16406,N_14354,N_11718);
nor U16407 (N_16407,N_13484,N_12443);
xor U16408 (N_16408,N_12636,N_14336);
nand U16409 (N_16409,N_14768,N_14533);
and U16410 (N_16410,N_10350,N_12446);
and U16411 (N_16411,N_14429,N_11035);
nor U16412 (N_16412,N_14547,N_11326);
nand U16413 (N_16413,N_12221,N_12165);
xor U16414 (N_16414,N_12284,N_13535);
xnor U16415 (N_16415,N_12741,N_14735);
xor U16416 (N_16416,N_12486,N_14500);
xnor U16417 (N_16417,N_10458,N_11790);
xor U16418 (N_16418,N_14674,N_12989);
or U16419 (N_16419,N_11538,N_10413);
xnor U16420 (N_16420,N_14859,N_13004);
and U16421 (N_16421,N_10140,N_12377);
and U16422 (N_16422,N_11845,N_12979);
or U16423 (N_16423,N_11917,N_10527);
and U16424 (N_16424,N_12143,N_13737);
nand U16425 (N_16425,N_13471,N_13106);
and U16426 (N_16426,N_13659,N_10213);
nand U16427 (N_16427,N_14492,N_12329);
nor U16428 (N_16428,N_12167,N_10275);
nor U16429 (N_16429,N_13599,N_14471);
and U16430 (N_16430,N_10142,N_14969);
xnor U16431 (N_16431,N_12939,N_13208);
xor U16432 (N_16432,N_10092,N_12884);
nor U16433 (N_16433,N_11344,N_12747);
xor U16434 (N_16434,N_12452,N_11685);
xor U16435 (N_16435,N_13340,N_13040);
nand U16436 (N_16436,N_10309,N_12344);
and U16437 (N_16437,N_13316,N_12054);
nand U16438 (N_16438,N_10165,N_12531);
nor U16439 (N_16439,N_12721,N_10335);
nand U16440 (N_16440,N_13059,N_14721);
and U16441 (N_16441,N_13796,N_12712);
xor U16442 (N_16442,N_12079,N_10467);
or U16443 (N_16443,N_14955,N_14565);
or U16444 (N_16444,N_11307,N_11031);
or U16445 (N_16445,N_10804,N_11312);
nand U16446 (N_16446,N_10226,N_14240);
nand U16447 (N_16447,N_11190,N_13331);
or U16448 (N_16448,N_13654,N_11929);
and U16449 (N_16449,N_14269,N_12644);
xnor U16450 (N_16450,N_13394,N_10833);
or U16451 (N_16451,N_10177,N_14593);
and U16452 (N_16452,N_10842,N_11762);
nand U16453 (N_16453,N_12562,N_10317);
nand U16454 (N_16454,N_14476,N_10766);
or U16455 (N_16455,N_14149,N_12578);
and U16456 (N_16456,N_10141,N_14811);
or U16457 (N_16457,N_12502,N_14138);
nand U16458 (N_16458,N_11384,N_14813);
nand U16459 (N_16459,N_10513,N_13636);
or U16460 (N_16460,N_14311,N_13526);
and U16461 (N_16461,N_10721,N_14968);
nand U16462 (N_16462,N_13031,N_11869);
and U16463 (N_16463,N_14340,N_14736);
nor U16464 (N_16464,N_10324,N_12662);
nand U16465 (N_16465,N_11171,N_10490);
nor U16466 (N_16466,N_11192,N_12868);
nand U16467 (N_16467,N_12420,N_13339);
and U16468 (N_16468,N_13941,N_11961);
xor U16469 (N_16469,N_13060,N_10926);
xnor U16470 (N_16470,N_11459,N_14978);
xnor U16471 (N_16471,N_12915,N_12894);
xnor U16472 (N_16472,N_14170,N_13884);
or U16473 (N_16473,N_12853,N_12334);
nand U16474 (N_16474,N_13035,N_14173);
nand U16475 (N_16475,N_11831,N_12816);
xnor U16476 (N_16476,N_13473,N_12408);
nand U16477 (N_16477,N_13861,N_11755);
or U16478 (N_16478,N_10210,N_11550);
xnor U16479 (N_16479,N_10683,N_11277);
or U16480 (N_16480,N_10170,N_13590);
nor U16481 (N_16481,N_11778,N_13614);
nand U16482 (N_16482,N_12572,N_13224);
nor U16483 (N_16483,N_10822,N_12497);
or U16484 (N_16484,N_13349,N_14863);
nor U16485 (N_16485,N_14086,N_11058);
and U16486 (N_16486,N_12592,N_10839);
nor U16487 (N_16487,N_11877,N_14950);
nor U16488 (N_16488,N_10201,N_11942);
xnor U16489 (N_16489,N_13160,N_10085);
or U16490 (N_16490,N_10605,N_12709);
xnor U16491 (N_16491,N_11907,N_13310);
nor U16492 (N_16492,N_12821,N_11833);
or U16493 (N_16493,N_14023,N_11099);
or U16494 (N_16494,N_11201,N_10913);
xnor U16495 (N_16495,N_10040,N_12005);
xnor U16496 (N_16496,N_12338,N_14523);
and U16497 (N_16497,N_10707,N_11368);
and U16498 (N_16498,N_14614,N_10172);
nor U16499 (N_16499,N_11447,N_10890);
nor U16500 (N_16500,N_13273,N_10860);
nand U16501 (N_16501,N_13995,N_13974);
xnor U16502 (N_16502,N_11903,N_11194);
nor U16503 (N_16503,N_10796,N_10072);
and U16504 (N_16504,N_10113,N_14235);
and U16505 (N_16505,N_13169,N_13799);
nand U16506 (N_16506,N_11390,N_14549);
or U16507 (N_16507,N_12406,N_14017);
nor U16508 (N_16508,N_13582,N_13242);
nor U16509 (N_16509,N_14494,N_10243);
nand U16510 (N_16510,N_13221,N_10454);
nor U16511 (N_16511,N_14505,N_13161);
nor U16512 (N_16512,N_12071,N_11445);
nand U16513 (N_16513,N_10863,N_13579);
and U16514 (N_16514,N_14910,N_10262);
or U16515 (N_16515,N_13475,N_12694);
nand U16516 (N_16516,N_13887,N_10745);
and U16517 (N_16517,N_11543,N_10637);
xnor U16518 (N_16518,N_10574,N_12262);
nor U16519 (N_16519,N_12432,N_11608);
nor U16520 (N_16520,N_14854,N_12745);
and U16521 (N_16521,N_10627,N_14960);
nor U16522 (N_16522,N_13099,N_13435);
xnor U16523 (N_16523,N_11360,N_13742);
or U16524 (N_16524,N_14899,N_10216);
xnor U16525 (N_16525,N_11977,N_12295);
and U16526 (N_16526,N_10028,N_14361);
xor U16527 (N_16527,N_12543,N_11908);
nand U16528 (N_16528,N_13368,N_14313);
and U16529 (N_16529,N_10329,N_10791);
nor U16530 (N_16530,N_11015,N_11986);
nand U16531 (N_16531,N_14283,N_10453);
or U16532 (N_16532,N_11444,N_14695);
and U16533 (N_16533,N_10782,N_10805);
or U16534 (N_16534,N_11240,N_12943);
or U16535 (N_16535,N_12849,N_11633);
nor U16536 (N_16536,N_12441,N_10360);
nand U16537 (N_16537,N_12751,N_12418);
and U16538 (N_16538,N_12209,N_12657);
nand U16539 (N_16539,N_12660,N_10128);
and U16540 (N_16540,N_10717,N_12670);
xnor U16541 (N_16541,N_14840,N_13883);
and U16542 (N_16542,N_10111,N_11080);
or U16543 (N_16543,N_13115,N_11606);
or U16544 (N_16544,N_10648,N_14163);
and U16545 (N_16545,N_13287,N_10221);
and U16546 (N_16546,N_12844,N_13485);
nand U16547 (N_16547,N_12148,N_10638);
or U16548 (N_16548,N_12568,N_12560);
nand U16549 (N_16549,N_10572,N_13055);
or U16550 (N_16550,N_14490,N_13801);
and U16551 (N_16551,N_10594,N_10307);
xnor U16552 (N_16552,N_14385,N_10062);
or U16553 (N_16553,N_14864,N_13330);
nor U16554 (N_16554,N_12339,N_11090);
and U16555 (N_16555,N_13618,N_14932);
and U16556 (N_16556,N_11832,N_11656);
nand U16557 (N_16557,N_11107,N_13765);
nor U16558 (N_16558,N_14898,N_11356);
and U16559 (N_16559,N_13685,N_14084);
and U16560 (N_16560,N_11841,N_12616);
or U16561 (N_16561,N_12487,N_14958);
xor U16562 (N_16562,N_11027,N_10787);
or U16563 (N_16563,N_12899,N_10752);
nand U16564 (N_16564,N_14575,N_14279);
or U16565 (N_16565,N_14442,N_13878);
nand U16566 (N_16566,N_13507,N_13518);
and U16567 (N_16567,N_14356,N_10153);
xor U16568 (N_16568,N_12607,N_12813);
nand U16569 (N_16569,N_14751,N_14861);
or U16570 (N_16570,N_14676,N_10189);
xnor U16571 (N_16571,N_10746,N_13240);
and U16572 (N_16572,N_10976,N_10903);
nand U16573 (N_16573,N_13183,N_14026);
nand U16574 (N_16574,N_12933,N_10742);
nor U16575 (N_16575,N_11952,N_12893);
xor U16576 (N_16576,N_13976,N_14669);
or U16577 (N_16577,N_12602,N_13700);
and U16578 (N_16578,N_13691,N_11620);
nand U16579 (N_16579,N_14744,N_14902);
nand U16580 (N_16580,N_13461,N_12688);
and U16581 (N_16581,N_11226,N_12789);
nor U16582 (N_16582,N_12504,N_12272);
nor U16583 (N_16583,N_12082,N_12511);
xnor U16584 (N_16584,N_10222,N_11730);
xnor U16585 (N_16585,N_12036,N_14794);
and U16586 (N_16586,N_12658,N_13994);
xor U16587 (N_16587,N_10723,N_12749);
and U16588 (N_16588,N_14245,N_11411);
nand U16589 (N_16589,N_12622,N_13078);
or U16590 (N_16590,N_12703,N_10249);
xor U16591 (N_16591,N_11632,N_14010);
xor U16592 (N_16592,N_10874,N_14918);
and U16593 (N_16593,N_14238,N_11337);
or U16594 (N_16594,N_13657,N_12628);
nand U16595 (N_16595,N_10155,N_12600);
or U16596 (N_16596,N_13322,N_10589);
nor U16597 (N_16597,N_12086,N_11157);
nand U16598 (N_16598,N_11605,N_11750);
or U16599 (N_16599,N_11361,N_14031);
xor U16600 (N_16600,N_14867,N_13741);
xor U16601 (N_16601,N_10446,N_12251);
and U16602 (N_16602,N_13511,N_10816);
xor U16603 (N_16603,N_12394,N_10401);
xnor U16604 (N_16604,N_13576,N_11145);
or U16605 (N_16605,N_11468,N_10389);
nand U16606 (N_16606,N_14525,N_12993);
nor U16607 (N_16607,N_11216,N_11136);
and U16608 (N_16608,N_14479,N_13926);
xor U16609 (N_16609,N_13012,N_11948);
nand U16610 (N_16610,N_13249,N_10208);
or U16611 (N_16611,N_13422,N_11388);
nor U16612 (N_16612,N_11084,N_11876);
and U16613 (N_16613,N_12414,N_11070);
or U16614 (N_16614,N_14836,N_12530);
nor U16615 (N_16615,N_12234,N_11779);
and U16616 (N_16616,N_12298,N_12057);
nor U16617 (N_16617,N_13206,N_10429);
xor U16618 (N_16618,N_14432,N_10942);
nor U16619 (N_16619,N_14979,N_14986);
xor U16620 (N_16620,N_10147,N_11815);
and U16621 (N_16621,N_13075,N_11158);
nor U16622 (N_16622,N_11178,N_11870);
nor U16623 (N_16623,N_14314,N_12829);
xor U16624 (N_16624,N_11573,N_12911);
xor U16625 (N_16625,N_10263,N_12545);
xnor U16626 (N_16626,N_14925,N_11341);
and U16627 (N_16627,N_12526,N_10949);
nor U16628 (N_16628,N_12354,N_10301);
xor U16629 (N_16629,N_11117,N_12699);
or U16630 (N_16630,N_14702,N_13486);
nor U16631 (N_16631,N_13109,N_11512);
nand U16632 (N_16632,N_12565,N_13921);
or U16633 (N_16633,N_11937,N_14816);
xor U16634 (N_16634,N_10852,N_12593);
xor U16635 (N_16635,N_12324,N_13555);
and U16636 (N_16636,N_13347,N_10283);
or U16637 (N_16637,N_10377,N_14795);
and U16638 (N_16638,N_12090,N_10215);
or U16639 (N_16639,N_10268,N_14198);
xor U16640 (N_16640,N_11340,N_14151);
xnor U16641 (N_16641,N_11392,N_14595);
nand U16642 (N_16642,N_14568,N_13909);
nor U16643 (N_16643,N_13423,N_12144);
and U16644 (N_16644,N_14728,N_11539);
nor U16645 (N_16645,N_12128,N_11629);
nand U16646 (N_16646,N_12012,N_13792);
xor U16647 (N_16647,N_14633,N_14333);
or U16648 (N_16648,N_10602,N_12056);
xnor U16649 (N_16649,N_11249,N_11627);
nand U16650 (N_16650,N_13522,N_11363);
and U16651 (N_16651,N_14202,N_10313);
and U16652 (N_16652,N_14094,N_14772);
or U16653 (N_16653,N_13964,N_12881);
xnor U16654 (N_16654,N_14259,N_14291);
xnor U16655 (N_16655,N_13982,N_10685);
xor U16656 (N_16656,N_13623,N_11773);
xnor U16657 (N_16657,N_11119,N_14177);
xnor U16658 (N_16658,N_10664,N_12973);
or U16659 (N_16659,N_14079,N_13298);
and U16660 (N_16660,N_10465,N_14322);
xnor U16661 (N_16661,N_14366,N_11966);
nand U16662 (N_16662,N_12392,N_14327);
nor U16663 (N_16663,N_14814,N_12533);
nand U16664 (N_16664,N_10654,N_12357);
nand U16665 (N_16665,N_10083,N_10573);
and U16666 (N_16666,N_10006,N_14146);
and U16667 (N_16667,N_10663,N_12755);
or U16668 (N_16668,N_12718,N_10771);
or U16669 (N_16669,N_10518,N_10484);
nand U16670 (N_16670,N_14653,N_12116);
and U16671 (N_16671,N_13091,N_11795);
nor U16672 (N_16672,N_11517,N_10536);
xor U16673 (N_16673,N_12104,N_12173);
nand U16674 (N_16674,N_14452,N_11001);
or U16675 (N_16675,N_13094,N_14563);
or U16676 (N_16676,N_11699,N_11174);
nand U16677 (N_16677,N_10690,N_10242);
and U16678 (N_16678,N_12514,N_11743);
and U16679 (N_16679,N_14080,N_11417);
nand U16680 (N_16680,N_14463,N_11513);
nand U16681 (N_16681,N_14207,N_10311);
nand U16682 (N_16682,N_10176,N_12023);
xor U16683 (N_16683,N_12031,N_14041);
xor U16684 (N_16684,N_13418,N_10808);
and U16685 (N_16685,N_11734,N_12282);
xnor U16686 (N_16686,N_14305,N_13353);
nor U16687 (N_16687,N_14157,N_13759);
and U16688 (N_16688,N_14520,N_14445);
xor U16689 (N_16689,N_10047,N_10384);
nor U16690 (N_16690,N_14037,N_13881);
and U16691 (N_16691,N_13826,N_13289);
nand U16692 (N_16692,N_12841,N_12505);
nor U16693 (N_16693,N_14782,N_14625);
and U16694 (N_16694,N_10206,N_11650);
or U16695 (N_16695,N_12854,N_14632);
nand U16696 (N_16696,N_10019,N_10033);
and U16697 (N_16697,N_12343,N_11096);
or U16698 (N_16698,N_12140,N_12605);
or U16699 (N_16699,N_12877,N_14369);
nand U16700 (N_16700,N_14534,N_12096);
nor U16701 (N_16701,N_13972,N_10159);
nor U16702 (N_16702,N_10496,N_14601);
nand U16703 (N_16703,N_10684,N_12965);
nor U16704 (N_16704,N_12175,N_14439);
or U16705 (N_16705,N_11038,N_12078);
nor U16706 (N_16706,N_11041,N_10819);
or U16707 (N_16707,N_13207,N_13529);
nand U16708 (N_16708,N_13436,N_12047);
and U16709 (N_16709,N_12216,N_13154);
xnor U16710 (N_16710,N_12956,N_14065);
nand U16711 (N_16711,N_10509,N_14644);
nand U16712 (N_16712,N_10921,N_10877);
nor U16713 (N_16713,N_14557,N_11061);
and U16714 (N_16714,N_14387,N_11068);
xor U16715 (N_16715,N_11819,N_11796);
and U16716 (N_16716,N_13592,N_10964);
and U16717 (N_16717,N_10978,N_13598);
nor U16718 (N_16718,N_10185,N_13930);
and U16719 (N_16719,N_12032,N_14048);
and U16720 (N_16720,N_11083,N_13162);
or U16721 (N_16721,N_14007,N_10777);
and U16722 (N_16722,N_13072,N_12824);
nand U16723 (N_16723,N_14937,N_11560);
or U16724 (N_16724,N_14716,N_14791);
or U16725 (N_16725,N_12576,N_13537);
nand U16726 (N_16726,N_13343,N_13048);
xor U16727 (N_16727,N_13278,N_14830);
and U16728 (N_16728,N_13455,N_10609);
xnor U16729 (N_16729,N_10891,N_13174);
nand U16730 (N_16730,N_12875,N_14686);
or U16731 (N_16731,N_12551,N_12060);
xnor U16732 (N_16732,N_12376,N_10731);
nand U16733 (N_16733,N_12362,N_13975);
nand U16734 (N_16734,N_11308,N_14097);
and U16735 (N_16735,N_14000,N_13027);
or U16736 (N_16736,N_14008,N_14466);
nand U16737 (N_16737,N_10669,N_12346);
nand U16738 (N_16738,N_10327,N_14901);
and U16739 (N_16739,N_11674,N_12589);
nand U16740 (N_16740,N_13112,N_11426);
and U16741 (N_16741,N_10607,N_10218);
nor U16742 (N_16742,N_10234,N_14964);
nor U16743 (N_16743,N_11450,N_12495);
nor U16744 (N_16744,N_12201,N_10182);
nor U16745 (N_16745,N_11757,N_14053);
and U16746 (N_16746,N_14206,N_12009);
nand U16747 (N_16747,N_11324,N_14739);
and U16748 (N_16748,N_13041,N_10767);
or U16749 (N_16749,N_10134,N_11954);
xnor U16750 (N_16750,N_10503,N_12236);
and U16751 (N_16751,N_11487,N_14952);
nor U16752 (N_16752,N_13239,N_12095);
or U16753 (N_16753,N_10044,N_12752);
nand U16754 (N_16754,N_14422,N_13678);
xnor U16755 (N_16755,N_14129,N_10769);
and U16756 (N_16756,N_14623,N_12291);
xnor U16757 (N_16757,N_12617,N_12883);
nor U16758 (N_16758,N_10452,N_14887);
xor U16759 (N_16759,N_13188,N_10095);
nand U16760 (N_16760,N_13235,N_12129);
xor U16761 (N_16761,N_10489,N_14268);
or U16762 (N_16762,N_12879,N_12538);
or U16763 (N_16763,N_10009,N_14996);
and U16764 (N_16764,N_12847,N_10125);
or U16765 (N_16765,N_12768,N_10878);
or U16766 (N_16766,N_12419,N_10466);
xor U16767 (N_16767,N_13564,N_12922);
or U16768 (N_16768,N_12030,N_12122);
nand U16769 (N_16769,N_12039,N_11978);
xor U16770 (N_16770,N_11541,N_11431);
and U16771 (N_16771,N_11005,N_14497);
or U16772 (N_16772,N_12449,N_11971);
and U16773 (N_16773,N_12076,N_13202);
or U16774 (N_16774,N_13073,N_13536);
xor U16775 (N_16775,N_13823,N_10278);
or U16776 (N_16776,N_10702,N_11945);
or U16777 (N_16777,N_10027,N_10423);
xor U16778 (N_16778,N_11963,N_10427);
xor U16779 (N_16779,N_11504,N_12246);
or U16780 (N_16780,N_11786,N_14001);
nor U16781 (N_16781,N_14582,N_13707);
or U16782 (N_16782,N_11505,N_10630);
nand U16783 (N_16783,N_14720,N_13669);
nor U16784 (N_16784,N_10419,N_11215);
or U16785 (N_16785,N_12638,N_12773);
xor U16786 (N_16786,N_14278,N_14114);
and U16787 (N_16787,N_13920,N_11492);
and U16788 (N_16788,N_10378,N_10352);
nand U16789 (N_16789,N_10372,N_13122);
and U16790 (N_16790,N_11032,N_11396);
or U16791 (N_16791,N_13153,N_11451);
or U16792 (N_16792,N_14540,N_12801);
and U16793 (N_16793,N_12587,N_10502);
or U16794 (N_16794,N_10768,N_13070);
and U16795 (N_16795,N_12328,N_13113);
xnor U16796 (N_16796,N_11284,N_12110);
xnor U16797 (N_16797,N_13464,N_14203);
nand U16798 (N_16798,N_10288,N_14004);
and U16799 (N_16799,N_14247,N_14194);
nor U16800 (N_16800,N_12019,N_10124);
or U16801 (N_16801,N_14804,N_10512);
or U16802 (N_16802,N_12285,N_14553);
xnor U16803 (N_16803,N_11455,N_12200);
and U16804 (N_16804,N_12836,N_11262);
nand U16805 (N_16805,N_10829,N_10856);
and U16806 (N_16806,N_13751,N_10510);
xor U16807 (N_16807,N_12876,N_10251);
xor U16808 (N_16808,N_11449,N_14438);
xor U16809 (N_16809,N_10834,N_13795);
nand U16810 (N_16810,N_10428,N_12033);
and U16811 (N_16811,N_13296,N_14723);
and U16812 (N_16812,N_11731,N_14627);
nand U16813 (N_16813,N_14891,N_14538);
xnor U16814 (N_16814,N_11208,N_11259);
xnor U16815 (N_16815,N_11800,N_11905);
nor U16816 (N_16816,N_13557,N_10245);
nand U16817 (N_16817,N_12491,N_13291);
or U16818 (N_16818,N_13063,N_12274);
and U16819 (N_16819,N_11409,N_10910);
and U16820 (N_16820,N_10588,N_10825);
or U16821 (N_16821,N_10357,N_13170);
nor U16822 (N_16822,N_12195,N_11854);
and U16823 (N_16823,N_10888,N_14306);
nor U16824 (N_16824,N_13467,N_13023);
nor U16825 (N_16825,N_11514,N_14842);
or U16826 (N_16826,N_12127,N_11347);
or U16827 (N_16827,N_12093,N_10954);
xnor U16828 (N_16828,N_13009,N_14161);
and U16829 (N_16829,N_12235,N_13355);
nor U16830 (N_16830,N_13282,N_14894);
nand U16831 (N_16831,N_12213,N_14507);
and U16832 (N_16832,N_14913,N_14230);
nand U16833 (N_16833,N_11128,N_12473);
or U16834 (N_16834,N_13419,N_11147);
nor U16835 (N_16835,N_10982,N_10302);
nor U16836 (N_16836,N_13480,N_12375);
nor U16837 (N_16837,N_14218,N_13414);
xnor U16838 (N_16838,N_10455,N_12575);
or U16839 (N_16839,N_11717,N_12772);
or U16840 (N_16840,N_10667,N_12306);
nor U16841 (N_16841,N_12784,N_10665);
xnor U16842 (N_16842,N_10000,N_13416);
xnor U16843 (N_16843,N_12742,N_12734);
nand U16844 (N_16844,N_12335,N_12326);
xnor U16845 (N_16845,N_13477,N_12415);
or U16846 (N_16846,N_13666,N_10778);
or U16847 (N_16847,N_10904,N_10744);
nor U16848 (N_16848,N_12484,N_13684);
nand U16849 (N_16849,N_12421,N_14954);
nand U16850 (N_16850,N_14055,N_12856);
or U16851 (N_16851,N_14225,N_13212);
nor U16852 (N_16852,N_11386,N_12948);
nor U16853 (N_16853,N_10780,N_11186);
nand U16854 (N_16854,N_14043,N_13569);
or U16855 (N_16855,N_11293,N_14234);
nor U16856 (N_16856,N_14211,N_11998);
xor U16857 (N_16857,N_13125,N_12793);
xor U16858 (N_16858,N_11309,N_13652);
and U16859 (N_16859,N_11150,N_12573);
xor U16860 (N_16860,N_14100,N_12325);
xnor U16861 (N_16861,N_12510,N_13726);
xor U16862 (N_16862,N_12604,N_14221);
nand U16863 (N_16863,N_14603,N_11210);
nor U16864 (N_16864,N_12124,N_14178);
or U16865 (N_16865,N_14123,N_14789);
and U16866 (N_16866,N_10590,N_10941);
xor U16867 (N_16867,N_11582,N_11910);
nand U16868 (N_16868,N_13505,N_10540);
nor U16869 (N_16869,N_12728,N_12215);
or U16870 (N_16870,N_14865,N_13100);
nand U16871 (N_16871,N_13144,N_10382);
nand U16872 (N_16872,N_11056,N_13024);
xor U16873 (N_16873,N_14991,N_13214);
xnor U16874 (N_16874,N_10722,N_12975);
nor U16875 (N_16875,N_12763,N_13829);
nor U16876 (N_16876,N_10238,N_14323);
and U16877 (N_16877,N_13465,N_11760);
xor U16878 (N_16878,N_12676,N_11713);
xnor U16879 (N_16879,N_13008,N_13336);
nor U16880 (N_16880,N_13577,N_11394);
and U16881 (N_16881,N_12761,N_13625);
nor U16882 (N_16882,N_14664,N_13963);
and U16883 (N_16883,N_11317,N_11374);
xnor U16884 (N_16884,N_13996,N_11162);
nand U16885 (N_16885,N_12149,N_14551);
and U16886 (N_16886,N_11304,N_10225);
and U16887 (N_16887,N_12765,N_14503);
or U16888 (N_16888,N_11871,N_14140);
and U16889 (N_16889,N_14109,N_12467);
xor U16890 (N_16890,N_14518,N_14124);
xnor U16891 (N_16891,N_11042,N_13632);
nand U16892 (N_16892,N_11735,N_14544);
xor U16893 (N_16893,N_12904,N_14831);
and U16894 (N_16894,N_12581,N_14315);
and U16895 (N_16895,N_10882,N_10195);
and U16896 (N_16896,N_10253,N_14156);
and U16897 (N_16897,N_13723,N_11236);
nand U16898 (N_16898,N_11030,N_10323);
nor U16899 (N_16899,N_10975,N_11690);
nand U16900 (N_16900,N_14947,N_11484);
xnor U16901 (N_16901,N_10012,N_14693);
xnor U16902 (N_16902,N_11586,N_13734);
nand U16903 (N_16903,N_14915,N_14302);
or U16904 (N_16904,N_11575,N_12839);
nand U16905 (N_16905,N_14184,N_14652);
nor U16906 (N_16906,N_11701,N_14351);
nand U16907 (N_16907,N_12429,N_14175);
nand U16908 (N_16908,N_12509,N_12107);
nand U16909 (N_16909,N_10715,N_11909);
xnor U16910 (N_16910,N_14550,N_12440);
and U16911 (N_16911,N_11245,N_11239);
nand U16912 (N_16912,N_14226,N_10793);
xnor U16913 (N_16913,N_10934,N_11901);
nand U16914 (N_16914,N_12229,N_10616);
nand U16915 (N_16915,N_10239,N_14588);
or U16916 (N_16916,N_12697,N_13037);
nor U16917 (N_16917,N_10658,N_11524);
nor U16918 (N_16918,N_10130,N_13646);
and U16919 (N_16919,N_11600,N_14413);
xor U16920 (N_16920,N_13698,N_13255);
xor U16921 (N_16921,N_11612,N_13246);
and U16922 (N_16922,N_13412,N_13777);
xnor U16923 (N_16923,N_10830,N_14112);
xor U16924 (N_16924,N_14809,N_11268);
and U16925 (N_16925,N_10864,N_12270);
and U16926 (N_16926,N_11323,N_12561);
nor U16927 (N_16927,N_10220,N_10460);
xnor U16928 (N_16928,N_14006,N_13248);
nand U16929 (N_16929,N_14758,N_11898);
or U16930 (N_16930,N_11792,N_10750);
xnor U16931 (N_16931,N_13764,N_13442);
and U16932 (N_16932,N_13525,N_11097);
xor U16933 (N_16933,N_11322,N_11327);
or U16934 (N_16934,N_12117,N_10108);
and U16935 (N_16935,N_13593,N_13517);
nor U16936 (N_16936,N_14249,N_10212);
and U16937 (N_16937,N_10556,N_13946);
nor U16938 (N_16938,N_12656,N_10475);
nand U16939 (N_16939,N_10907,N_11702);
nor U16940 (N_16940,N_14092,N_10855);
or U16941 (N_16941,N_11895,N_11631);
xnor U16942 (N_16942,N_13912,N_11564);
and U16943 (N_16943,N_10548,N_11593);
xor U16944 (N_16944,N_14620,N_11095);
nand U16945 (N_16945,N_13998,N_13867);
and U16946 (N_16946,N_12184,N_10451);
nand U16947 (N_16947,N_13502,N_14287);
nor U16948 (N_16948,N_10463,N_14244);
and U16949 (N_16949,N_12878,N_12407);
nor U16950 (N_16950,N_10017,N_11172);
xnor U16951 (N_16951,N_13591,N_10076);
nor U16952 (N_16952,N_11643,N_11648);
nor U16953 (N_16953,N_10762,N_13872);
or U16954 (N_16954,N_13738,N_14319);
and U16955 (N_16955,N_11530,N_14280);
and U16956 (N_16956,N_12203,N_13834);
or U16957 (N_16957,N_10732,N_11206);
and U16958 (N_16958,N_14022,N_12044);
nor U16959 (N_16959,N_12930,N_13933);
nor U16960 (N_16960,N_11497,N_13047);
or U16961 (N_16961,N_13105,N_13058);
nor U16962 (N_16962,N_10264,N_11515);
nor U16963 (N_16963,N_14473,N_14555);
and U16964 (N_16964,N_13922,N_13430);
xnor U16965 (N_16965,N_10281,N_13762);
and U16966 (N_16966,N_12736,N_10965);
or U16967 (N_16967,N_11398,N_12785);
and U16968 (N_16968,N_12187,N_10211);
xnor U16969 (N_16969,N_13216,N_10933);
nor U16970 (N_16970,N_13251,N_13053);
nor U16971 (N_16971,N_12138,N_13155);
nand U16972 (N_16972,N_13056,N_14113);
nand U16973 (N_16973,N_14826,N_12018);
nand U16974 (N_16974,N_10116,N_14499);
nand U16975 (N_16975,N_11856,N_11401);
xnor U16976 (N_16976,N_13704,N_10348);
nand U16977 (N_16977,N_12760,N_12725);
or U16978 (N_16978,N_11924,N_14484);
nand U16979 (N_16979,N_14872,N_13083);
or U16980 (N_16980,N_11372,N_12385);
or U16981 (N_16981,N_10797,N_14738);
nor U16982 (N_16982,N_14895,N_10634);
nor U16983 (N_16983,N_12758,N_14905);
nand U16984 (N_16984,N_14148,N_12202);
nand U16985 (N_16985,N_13238,N_11173);
and U16986 (N_16986,N_14528,N_13955);
nor U16987 (N_16987,N_12279,N_10029);
nand U16988 (N_16988,N_14923,N_11148);
or U16989 (N_16989,N_11161,N_14179);
xor U16990 (N_16990,N_13038,N_14903);
xor U16991 (N_16991,N_13034,N_11082);
or U16992 (N_16992,N_11708,N_13266);
nand U16993 (N_16993,N_11075,N_14745);
nor U16994 (N_16994,N_10235,N_14324);
nor U16995 (N_16995,N_14018,N_14763);
xnor U16996 (N_16996,N_10841,N_10265);
xor U16997 (N_16997,N_12397,N_10929);
or U16998 (N_16998,N_13527,N_12471);
or U16999 (N_16999,N_11257,N_10366);
xnor U17000 (N_17000,N_13165,N_13837);
xor U17001 (N_17001,N_12469,N_14472);
and U17002 (N_17002,N_12689,N_10286);
nand U17003 (N_17003,N_12955,N_10854);
xnor U17004 (N_17004,N_10514,N_12383);
nand U17005 (N_17005,N_11142,N_11681);
nand U17006 (N_17006,N_14537,N_10747);
xor U17007 (N_17007,N_10751,N_11729);
or U17008 (N_17008,N_12111,N_14645);
nor U17009 (N_17009,N_11999,N_12294);
nand U17010 (N_17010,N_12974,N_11733);
and U17011 (N_17011,N_13908,N_10706);
nor U17012 (N_17012,N_11345,N_13842);
and U17013 (N_17013,N_14793,N_13342);
nor U17014 (N_17014,N_13750,N_14091);
or U17015 (N_17015,N_10480,N_11728);
xor U17016 (N_17016,N_10898,N_14264);
xor U17017 (N_17017,N_11229,N_14904);
nand U17018 (N_17018,N_12152,N_14171);
nor U17019 (N_17019,N_13327,N_13676);
nor U17020 (N_17020,N_11051,N_14448);
xor U17021 (N_17021,N_14742,N_13006);
xnor U17022 (N_17022,N_14137,N_14056);
xnor U17023 (N_17023,N_12905,N_12550);
nor U17024 (N_17024,N_14174,N_10755);
and U17025 (N_17025,N_10840,N_14946);
nor U17026 (N_17026,N_13655,N_12812);
or U17027 (N_17027,N_12006,N_13156);
nor U17028 (N_17028,N_14780,N_11135);
or U17029 (N_17029,N_13462,N_12825);
xor U17030 (N_17030,N_13934,N_12579);
or U17031 (N_17031,N_11100,N_11428);
xor U17032 (N_17032,N_10174,N_11931);
and U17033 (N_17033,N_11443,N_13095);
nor U17034 (N_17034,N_11321,N_13523);
xnor U17035 (N_17035,N_13335,N_13546);
and U17036 (N_17036,N_10422,N_12428);
and U17037 (N_17037,N_12811,N_14165);
nor U17038 (N_17038,N_11094,N_14088);
xnor U17039 (N_17039,N_12998,N_12641);
nand U17040 (N_17040,N_11886,N_14855);
or U17041 (N_17041,N_11464,N_13664);
nor U17042 (N_17042,N_10770,N_11894);
and U17043 (N_17043,N_11921,N_13076);
xor U17044 (N_17044,N_11342,N_12304);
or U17045 (N_17045,N_14348,N_14951);
nand U17046 (N_17046,N_12823,N_12567);
and U17047 (N_17047,N_11299,N_11105);
nor U17048 (N_17048,N_11688,N_12208);
nor U17049 (N_17049,N_11521,N_14344);
nand U17050 (N_17050,N_13562,N_12351);
xor U17051 (N_17051,N_10471,N_13337);
nor U17052 (N_17052,N_13622,N_11329);
and U17053 (N_17053,N_12146,N_12378);
and U17054 (N_17054,N_13721,N_11828);
or U17055 (N_17055,N_14039,N_13938);
nor U17056 (N_17056,N_13222,N_12870);
nor U17057 (N_17057,N_13286,N_14883);
xor U17058 (N_17058,N_10938,N_11233);
nor U17059 (N_17059,N_12885,N_10163);
or U17060 (N_17060,N_14337,N_14949);
and U17061 (N_17061,N_10018,N_10469);
nor U17062 (N_17062,N_10677,N_11682);
and U17063 (N_17063,N_10719,N_12123);
or U17064 (N_17064,N_12365,N_11170);
nand U17065 (N_17065,N_14810,N_13832);
and U17066 (N_17066,N_13178,N_12639);
or U17067 (N_17067,N_12020,N_13092);
nand U17068 (N_17068,N_14390,N_10295);
and U17069 (N_17069,N_12797,N_10233);
nor U17070 (N_17070,N_14358,N_10546);
nor U17071 (N_17071,N_10501,N_12947);
and U17072 (N_17072,N_12521,N_11545);
nand U17073 (N_17073,N_10969,N_11992);
xnor U17074 (N_17074,N_12539,N_12366);
nand U17075 (N_17075,N_10355,N_11480);
nand U17076 (N_17076,N_13087,N_11471);
nor U17077 (N_17077,N_11310,N_14386);
nand U17078 (N_17078,N_14705,N_13815);
xor U17079 (N_17079,N_12191,N_11810);
nor U17080 (N_17080,N_14254,N_13828);
and U17081 (N_17081,N_12953,N_13163);
nor U17082 (N_17082,N_13775,N_10989);
nand U17083 (N_17083,N_14335,N_14838);
nand U17084 (N_17084,N_12320,N_14938);
nor U17085 (N_17085,N_13831,N_11040);
or U17086 (N_17086,N_14769,N_14566);
or U17087 (N_17087,N_13114,N_11435);
nor U17088 (N_17088,N_11555,N_13413);
or U17089 (N_17089,N_14236,N_13398);
or U17090 (N_17090,N_12869,N_12136);
and U17091 (N_17091,N_12701,N_10368);
xnor U17092 (N_17092,N_13469,N_12629);
and U17093 (N_17093,N_11938,N_13853);
nand U17094 (N_17094,N_14498,N_13301);
nand U17095 (N_17095,N_10516,N_12088);
xnor U17096 (N_17096,N_12715,N_12455);
and U17097 (N_17097,N_14732,N_10008);
nor U17098 (N_17098,N_10774,N_12258);
nor U17099 (N_17099,N_14798,N_10284);
xor U17100 (N_17100,N_10069,N_14929);
xnor U17101 (N_17101,N_12094,N_12066);
or U17102 (N_17102,N_12609,N_13385);
or U17103 (N_17103,N_11683,N_13565);
nand U17104 (N_17104,N_10568,N_10204);
nand U17105 (N_17105,N_13175,N_12857);
nand U17106 (N_17106,N_14990,N_11571);
nor U17107 (N_17107,N_11446,N_10021);
nor U17108 (N_17108,N_10050,N_13575);
xnor U17109 (N_17109,N_12312,N_10096);
or U17110 (N_17110,N_14220,N_11533);
nor U17111 (N_17111,N_11036,N_14708);
and U17112 (N_17112,N_12256,N_12890);
nor U17113 (N_17113,N_14548,N_14342);
nand U17114 (N_17114,N_10100,N_12909);
and U17115 (N_17115,N_12685,N_13662);
nor U17116 (N_17116,N_12614,N_11721);
nor U17117 (N_17117,N_13400,N_10881);
and U17118 (N_17118,N_14585,N_12962);
nand U17119 (N_17119,N_11205,N_11944);
or U17120 (N_17120,N_13612,N_13424);
and U17121 (N_17121,N_11184,N_10790);
or U17122 (N_17122,N_14316,N_13387);
nand U17123 (N_17123,N_13274,N_14567);
nand U17124 (N_17124,N_10032,N_14293);
nor U17125 (N_17125,N_14457,N_10705);
xnor U17126 (N_17126,N_13952,N_12767);
xor U17127 (N_17127,N_10950,N_13911);
nor U17128 (N_17128,N_14154,N_12529);
xor U17129 (N_17129,N_11847,N_11867);
and U17130 (N_17130,N_13906,N_14985);
xor U17131 (N_17131,N_13538,N_10672);
or U17132 (N_17132,N_14622,N_10065);
or U17133 (N_17133,N_14648,N_12014);
nand U17134 (N_17134,N_11946,N_13877);
and U17135 (N_17135,N_12780,N_14057);
nand U17136 (N_17136,N_14416,N_14415);
xnor U17137 (N_17137,N_12189,N_12476);
or U17138 (N_17138,N_12035,N_13748);
and U17139 (N_17139,N_13586,N_10720);
nor U17140 (N_17140,N_12837,N_11837);
and U17141 (N_17141,N_12653,N_12822);
and U17142 (N_17142,N_10150,N_14604);
or U17143 (N_17143,N_10364,N_11039);
nor U17144 (N_17144,N_11842,N_10555);
nor U17145 (N_17145,N_12042,N_13081);
nand U17146 (N_17146,N_12318,N_14028);
nor U17147 (N_17147,N_10953,N_14786);
xnor U17148 (N_17148,N_10016,N_14047);
or U17149 (N_17149,N_13133,N_11723);
nor U17150 (N_17150,N_13789,N_12667);
and U17151 (N_17151,N_13567,N_12468);
nor U17152 (N_17152,N_13045,N_11872);
and U17153 (N_17153,N_10565,N_13030);
and U17154 (N_17154,N_12637,N_10340);
and U17155 (N_17155,N_11346,N_14975);
or U17156 (N_17156,N_13171,N_12809);
xor U17157 (N_17157,N_10620,N_13865);
nand U17158 (N_17158,N_10013,N_12537);
or U17159 (N_17159,N_14059,N_10103);
nor U17160 (N_17160,N_11829,N_13892);
xor U17161 (N_17161,N_13639,N_11213);
or U17162 (N_17162,N_13800,N_14003);
and U17163 (N_17163,N_12987,N_11915);
nor U17164 (N_17164,N_11248,N_11214);
nor U17165 (N_17165,N_10909,N_12217);
and U17166 (N_17166,N_14270,N_12067);
nor U17167 (N_17167,N_12485,N_11665);
nand U17168 (N_17168,N_10425,N_13708);
nand U17169 (N_17169,N_12118,N_13426);
nand U17170 (N_17170,N_13103,N_14192);
or U17171 (N_17171,N_12596,N_14624);
nor U17172 (N_17172,N_10541,N_11362);
and U17173 (N_17173,N_11421,N_10199);
nand U17174 (N_17174,N_12787,N_13168);
and U17175 (N_17175,N_11836,N_12700);
nand U17176 (N_17176,N_14168,N_13120);
and U17177 (N_17177,N_11802,N_10673);
nand U17178 (N_17178,N_13679,N_12091);
nor U17179 (N_17179,N_11389,N_10449);
nand U17180 (N_17180,N_10359,N_10078);
and U17181 (N_17181,N_13150,N_14506);
and U17182 (N_17182,N_11635,N_13816);
or U17183 (N_17183,N_11914,N_13129);
nor U17184 (N_17184,N_11077,N_13788);
or U17185 (N_17185,N_14334,N_14453);
or U17186 (N_17186,N_12681,N_14277);
nor U17187 (N_17187,N_13689,N_12434);
xor U17188 (N_17188,N_14443,N_13847);
or U17189 (N_17189,N_11441,N_10310);
nor U17190 (N_17190,N_14618,N_14399);
nor U17191 (N_17191,N_13320,N_11669);
or U17192 (N_17192,N_12131,N_12863);
or U17193 (N_17193,N_11671,N_14849);
nand U17194 (N_17194,N_13119,N_13137);
xor U17195 (N_17195,N_11926,N_12379);
xor U17196 (N_17196,N_10865,N_13265);
or U17197 (N_17197,N_13415,N_11160);
xnor U17198 (N_17198,N_12722,N_13506);
xnor U17199 (N_17199,N_11765,N_14651);
nand U17200 (N_17200,N_14481,N_11739);
xor U17201 (N_17201,N_12223,N_12654);
and U17202 (N_17202,N_10848,N_13954);
and U17203 (N_17203,N_11122,N_10294);
or U17204 (N_17204,N_12068,N_10802);
nand U17205 (N_17205,N_14027,N_12040);
xnor U17206 (N_17206,N_13123,N_14576);
xor U17207 (N_17207,N_10689,N_12247);
xor U17208 (N_17208,N_13490,N_12769);
xor U17209 (N_17209,N_14635,N_12743);
or U17210 (N_17210,N_13648,N_13096);
nor U17211 (N_17211,N_10578,N_12650);
xnor U17212 (N_17212,N_14392,N_13452);
xor U17213 (N_17213,N_13190,N_13186);
nand U17214 (N_17214,N_14143,N_12672);
or U17215 (N_17215,N_10657,N_10520);
nor U17216 (N_17216,N_13054,N_12305);
or U17217 (N_17217,N_13138,N_11044);
or U17218 (N_17218,N_12544,N_11140);
and U17219 (N_17219,N_14535,N_10998);
and U17220 (N_17220,N_14822,N_10345);
or U17221 (N_17221,N_11865,N_10227);
or U17222 (N_17222,N_13382,N_11678);
or U17223 (N_17223,N_10765,N_11241);
nor U17224 (N_17224,N_12171,N_14942);
or U17225 (N_17225,N_13524,N_11979);
or U17226 (N_17226,N_11662,N_14760);
xnor U17227 (N_17227,N_12470,N_13388);
and U17228 (N_17228,N_12373,N_12865);
xnor U17229 (N_17229,N_10414,N_14115);
or U17230 (N_17230,N_11956,N_12713);
nor U17231 (N_17231,N_11623,N_13066);
nor U17232 (N_17232,N_11325,N_14885);
or U17233 (N_17233,N_14755,N_13243);
or U17234 (N_17234,N_11947,N_11024);
and U17235 (N_17235,N_14364,N_10641);
or U17236 (N_17236,N_10550,N_10999);
or U17237 (N_17237,N_13191,N_14688);
or U17238 (N_17238,N_10570,N_11675);
or U17239 (N_17239,N_13609,N_14778);
nand U17240 (N_17240,N_14223,N_12178);
nor U17241 (N_17241,N_13608,N_12214);
and U17242 (N_17242,N_10961,N_10960);
and U17243 (N_17243,N_13254,N_10292);
nand U17244 (N_17244,N_13916,N_11724);
xor U17245 (N_17245,N_14176,N_10736);
nor U17246 (N_17246,N_14465,N_14851);
or U17247 (N_17247,N_13132,N_10632);
or U17248 (N_17248,N_13252,N_14253);
and U17249 (N_17249,N_12430,N_11976);
and U17250 (N_17250,N_13182,N_13352);
and U17251 (N_17251,N_13417,N_11794);
nand U17252 (N_17252,N_14967,N_14531);
and U17253 (N_17253,N_14920,N_10356);
xor U17254 (N_17254,N_11609,N_13509);
or U17255 (N_17255,N_10922,N_10606);
nand U17256 (N_17256,N_14900,N_10912);
or U17257 (N_17257,N_13719,N_14770);
xnor U17258 (N_17258,N_13268,N_11824);
nor U17259 (N_17259,N_14295,N_10436);
or U17260 (N_17260,N_10773,N_12011);
nand U17261 (N_17261,N_10219,N_13514);
nor U17262 (N_17262,N_11003,N_12260);
and U17263 (N_17263,N_13258,N_11525);
xnor U17264 (N_17264,N_13804,N_11177);
nand U17265 (N_17265,N_10328,N_10749);
or U17266 (N_17266,N_13943,N_10708);
nor U17267 (N_17267,N_13827,N_13359);
and U17268 (N_17268,N_12696,N_10697);
xnor U17269 (N_17269,N_10223,N_10093);
or U17270 (N_17270,N_13408,N_12181);
nor U17271 (N_17271,N_13613,N_10835);
nand U17272 (N_17272,N_11180,N_11278);
xor U17273 (N_17273,N_12815,N_13601);
nand U17274 (N_17274,N_14440,N_14352);
or U17275 (N_17275,N_12910,N_13284);
and U17276 (N_17276,N_14292,N_11852);
or U17277 (N_17277,N_11709,N_11523);
or U17278 (N_17278,N_12137,N_10558);
and U17279 (N_17279,N_12528,N_13756);
nor U17280 (N_17280,N_14586,N_10587);
nand U17281 (N_17281,N_14666,N_10080);
xor U17282 (N_17282,N_13042,N_12448);
and U17283 (N_17283,N_10643,N_14675);
nor U17284 (N_17284,N_11839,N_14656);
and U17285 (N_17285,N_13363,N_11022);
or U17286 (N_17286,N_13682,N_10036);
and U17287 (N_17287,N_10900,N_13164);
or U17288 (N_17288,N_11197,N_12795);
nor U17289 (N_17289,N_13980,N_13341);
nand U17290 (N_17290,N_11613,N_13844);
and U17291 (N_17291,N_12280,N_10918);
nor U17292 (N_17292,N_13315,N_10344);
nor U17293 (N_17293,N_14338,N_12160);
nand U17294 (N_17294,N_13859,N_14231);
or U17295 (N_17295,N_14710,N_11014);
xnor U17296 (N_17296,N_13838,N_14434);
xnor U17297 (N_17297,N_11797,N_12652);
nor U17298 (N_17298,N_10319,N_10477);
and U17299 (N_17299,N_11422,N_10396);
and U17300 (N_17300,N_14661,N_11375);
or U17301 (N_17301,N_14677,N_10704);
or U17302 (N_17302,N_10554,N_11576);
or U17303 (N_17303,N_13520,N_11098);
and U17304 (N_17304,N_11093,N_11964);
xnor U17305 (N_17305,N_10507,N_13187);
xnor U17306 (N_17306,N_11860,N_14222);
nor U17307 (N_17307,N_10651,N_11812);
and U17308 (N_17308,N_13817,N_11500);
and U17309 (N_17309,N_12360,N_13478);
nor U17310 (N_17310,N_13540,N_10788);
and U17311 (N_17311,N_10184,N_13089);
or U17312 (N_17312,N_10901,N_11578);
or U17313 (N_17313,N_13050,N_10925);
xnor U17314 (N_17314,N_10560,N_12402);
and U17315 (N_17315,N_11410,N_14529);
xor U17316 (N_17316,N_11649,N_11316);
and U17317 (N_17317,N_12642,N_11816);
or U17318 (N_17318,N_12512,N_12481);
xnor U17319 (N_17319,N_11079,N_14110);
or U17320 (N_17320,N_11116,N_13126);
nor U17321 (N_17321,N_10674,N_13365);
and U17322 (N_17322,N_10862,N_12445);
nor U17323 (N_17323,N_10200,N_14395);
and U17324 (N_17324,N_14102,N_12916);
or U17325 (N_17325,N_13786,N_11753);
nand U17326 (N_17326,N_14515,N_13836);
nor U17327 (N_17327,N_14626,N_12577);
or U17328 (N_17328,N_10827,N_10135);
and U17329 (N_17329,N_14049,N_14643);
and U17330 (N_17330,N_14715,N_10117);
nor U17331 (N_17331,N_14297,N_10911);
and U17332 (N_17332,N_10733,N_14104);
or U17333 (N_17333,N_14631,N_11217);
xnor U17334 (N_17334,N_10334,N_11962);
xnor U17335 (N_17335,N_12598,N_12723);
xnor U17336 (N_17336,N_13237,N_10604);
or U17337 (N_17337,N_13328,N_11134);
xor U17338 (N_17338,N_11878,N_11544);
nand U17339 (N_17339,N_10119,N_14866);
and U17340 (N_17340,N_13940,N_13626);
or U17341 (N_17341,N_13468,N_14142);
or U17342 (N_17342,N_13962,N_11818);
and U17343 (N_17343,N_12442,N_13979);
and U17344 (N_17344,N_13329,N_13754);
nand U17345 (N_17345,N_13882,N_13064);
and U17346 (N_17346,N_14396,N_11519);
or U17347 (N_17347,N_13378,N_14884);
and U17348 (N_17348,N_14332,N_14665);
nor U17349 (N_17349,N_12924,N_11004);
or U17350 (N_17350,N_13673,N_12072);
or U17351 (N_17351,N_12331,N_14199);
or U17352 (N_17352,N_12232,N_10905);
nand U17353 (N_17353,N_12966,N_11025);
nor U17354 (N_17354,N_12479,N_11367);
nand U17355 (N_17355,N_12925,N_12498);
xor U17356 (N_17356,N_10923,N_10701);
xnor U17357 (N_17357,N_14372,N_12254);
nor U17358 (N_17358,N_12499,N_12314);
and U17359 (N_17359,N_14420,N_13433);
and U17360 (N_17360,N_14730,N_14098);
and U17361 (N_17361,N_10498,N_13410);
xnor U17362 (N_17362,N_13584,N_11622);
xnor U17363 (N_17363,N_13262,N_10398);
or U17364 (N_17364,N_13871,N_13396);
or U17365 (N_17365,N_10600,N_11418);
or U17366 (N_17366,N_10803,N_11261);
nand U17367 (N_17367,N_13773,N_13250);
or U17368 (N_17368,N_10811,N_10566);
nand U17369 (N_17369,N_10445,N_10582);
and U17370 (N_17370,N_12684,N_10843);
and U17371 (N_17371,N_12895,N_11694);
nand U17372 (N_17372,N_10181,N_13910);
or U17373 (N_17373,N_14040,N_12886);
nand U17374 (N_17374,N_14729,N_12105);
and U17375 (N_17375,N_14992,N_11266);
nor U17376 (N_17376,N_14044,N_13136);
nor U17377 (N_17377,N_14425,N_12411);
xor U17378 (N_17378,N_14169,N_14491);
and U17379 (N_17379,N_11911,N_14734);
and U17380 (N_17380,N_11668,N_12866);
nand U17381 (N_17381,N_11331,N_13997);
nor U17382 (N_17382,N_10492,N_10010);
or U17383 (N_17383,N_11516,N_11437);
or U17384 (N_17384,N_13233,N_11526);
nor U17385 (N_17385,N_10034,N_14257);
or U17386 (N_17386,N_11062,N_14713);
or U17387 (N_17387,N_14771,N_12864);
nand U17388 (N_17388,N_10748,N_13606);
or U17389 (N_17389,N_14339,N_11296);
nand U17390 (N_17390,N_11534,N_14374);
xor U17391 (N_17391,N_12457,N_14046);
or U17392 (N_17392,N_10845,N_14303);
nand U17393 (N_17393,N_12901,N_10610);
or U17394 (N_17394,N_11969,N_12224);
or U17395 (N_17395,N_13629,N_14881);
or U17396 (N_17396,N_13453,N_12422);
nand U17397 (N_17397,N_11207,N_10237);
or U17398 (N_17398,N_10025,N_11423);
or U17399 (N_17399,N_13319,N_12727);
nor U17400 (N_17400,N_12307,N_10645);
xnor U17401 (N_17401,N_10561,N_13902);
nand U17402 (N_17402,N_13825,N_14806);
nand U17403 (N_17403,N_12705,N_13367);
and U17404 (N_17404,N_11928,N_14879);
or U17405 (N_17405,N_12738,N_10257);
nand U17406 (N_17406,N_10438,N_12926);
nor U17407 (N_17407,N_11758,N_12951);
nor U17408 (N_17408,N_10479,N_14820);
or U17409 (N_17409,N_10885,N_11930);
and U17410 (N_17410,N_12838,N_14182);
nor U17411 (N_17411,N_14880,N_13370);
xor U17412 (N_17412,N_11486,N_10178);
xnor U17413 (N_17413,N_14271,N_10358);
nand U17414 (N_17414,N_12783,N_10088);
and U17415 (N_17415,N_14224,N_13866);
and U17416 (N_17416,N_11621,N_13740);
and U17417 (N_17417,N_12807,N_12099);
nor U17418 (N_17418,N_10102,N_13724);
and U17419 (N_17419,N_10786,N_11994);
nand U17420 (N_17420,N_14468,N_13752);
nand U17421 (N_17421,N_10126,N_11891);
nand U17422 (N_17422,N_13351,N_14074);
or U17423 (N_17423,N_10534,N_14821);
or U17424 (N_17424,N_10417,N_12664);
nand U17425 (N_17425,N_10729,N_13875);
or U17426 (N_17426,N_13559,N_10022);
xor U17427 (N_17427,N_11737,N_10138);
or U17428 (N_17428,N_12805,N_14701);
or U17429 (N_17429,N_12480,N_10601);
nand U17430 (N_17430,N_10444,N_13709);
nor U17431 (N_17431,N_13204,N_13900);
nand U17432 (N_17432,N_11554,N_13903);
nor U17433 (N_17433,N_12022,N_11896);
and U17434 (N_17434,N_13108,N_12482);
or U17435 (N_17435,N_12583,N_13324);
nor U17436 (N_17436,N_10506,N_14063);
nor U17437 (N_17437,N_10522,N_13508);
nor U17438 (N_17438,N_10152,N_14818);
or U17439 (N_17439,N_11997,N_11433);
xor U17440 (N_17440,N_10670,N_11496);
nor U17441 (N_17441,N_12061,N_12923);
xnor U17442 (N_17442,N_10713,N_13850);
nand U17443 (N_17443,N_14130,N_10499);
xor U17444 (N_17444,N_12163,N_12994);
nor U17445 (N_17445,N_13148,N_12591);
and U17446 (N_17446,N_10623,N_13554);
nor U17447 (N_17447,N_10944,N_14454);
nor U17448 (N_17448,N_10365,N_12185);
nor U17449 (N_17449,N_14704,N_10915);
nor U17450 (N_17450,N_11985,N_14536);
or U17451 (N_17451,N_12034,N_10157);
and U17452 (N_17452,N_14265,N_14155);
xor U17453 (N_17453,N_14480,N_14733);
and U17454 (N_17454,N_11270,N_13421);
nand U17455 (N_17455,N_14190,N_10691);
or U17456 (N_17456,N_12323,N_10067);
or U17457 (N_17457,N_14122,N_12390);
nor U17458 (N_17458,N_12659,N_13500);
xnor U17459 (N_17459,N_13718,N_14308);
nor U17460 (N_17460,N_11124,N_14188);
nor U17461 (N_17461,N_13231,N_11473);
xor U17462 (N_17462,N_11355,N_13211);
nand U17463 (N_17463,N_11258,N_13079);
nand U17464 (N_17464,N_12369,N_12089);
nor U17465 (N_17465,N_10079,N_11861);
or U17466 (N_17466,N_14267,N_14747);
and U17467 (N_17467,N_14706,N_12892);
nor U17468 (N_17468,N_10682,N_13783);
or U17469 (N_17469,N_13603,N_14719);
nand U17470 (N_17470,N_10624,N_11407);
nor U17471 (N_17471,N_13173,N_13658);
xor U17472 (N_17472,N_10846,N_12400);
nor U17473 (N_17473,N_11283,N_10936);
xor U17474 (N_17474,N_10115,N_10146);
xor U17475 (N_17475,N_13472,N_13720);
xnor U17476 (N_17476,N_12570,N_10186);
nand U17477 (N_17477,N_14035,N_13677);
xor U17478 (N_17478,N_13147,N_12444);
nor U17479 (N_17479,N_13482,N_10613);
or U17480 (N_17480,N_11706,N_11602);
and U17481 (N_17481,N_11868,N_13504);
nand U17482 (N_17482,N_13924,N_10639);
nor U17483 (N_17483,N_11006,N_10551);
nand U17484 (N_17484,N_10500,N_13772);
nor U17485 (N_17485,N_14034,N_12309);
xor U17486 (N_17486,N_13195,N_14966);
nor U17487 (N_17487,N_10387,N_13856);
nand U17488 (N_17488,N_10180,N_11761);
xor U17489 (N_17489,N_11358,N_14858);
xnor U17490 (N_17490,N_14642,N_12500);
nand U17491 (N_17491,N_14077,N_10716);
nand U17492 (N_17492,N_10621,N_10048);
xor U17493 (N_17493,N_12049,N_11295);
xor U17494 (N_17494,N_14391,N_10070);
or U17495 (N_17495,N_13809,N_13863);
or U17496 (N_17496,N_12218,N_11452);
xnor U17497 (N_17497,N_11592,N_13862);
or U17498 (N_17498,N_12523,N_12097);
nor U17499 (N_17499,N_11566,N_13668);
nor U17500 (N_17500,N_13115,N_10402);
nor U17501 (N_17501,N_13460,N_11018);
and U17502 (N_17502,N_14893,N_10526);
or U17503 (N_17503,N_13387,N_11579);
xnor U17504 (N_17504,N_12737,N_13391);
or U17505 (N_17505,N_11158,N_11391);
xnor U17506 (N_17506,N_10399,N_12257);
or U17507 (N_17507,N_11562,N_12457);
nand U17508 (N_17508,N_13651,N_12638);
and U17509 (N_17509,N_14688,N_10504);
and U17510 (N_17510,N_13216,N_12482);
and U17511 (N_17511,N_10835,N_13445);
nand U17512 (N_17512,N_11601,N_10368);
or U17513 (N_17513,N_12405,N_12319);
nand U17514 (N_17514,N_12743,N_12873);
xor U17515 (N_17515,N_14138,N_13502);
nor U17516 (N_17516,N_10684,N_10819);
and U17517 (N_17517,N_12771,N_10352);
and U17518 (N_17518,N_12419,N_10192);
or U17519 (N_17519,N_11832,N_10298);
nand U17520 (N_17520,N_14049,N_10510);
xor U17521 (N_17521,N_13355,N_11753);
and U17522 (N_17522,N_10179,N_12628);
xor U17523 (N_17523,N_10706,N_10111);
or U17524 (N_17524,N_13024,N_14883);
or U17525 (N_17525,N_11698,N_12869);
nand U17526 (N_17526,N_10492,N_10636);
xor U17527 (N_17527,N_10845,N_13405);
nor U17528 (N_17528,N_14938,N_14621);
and U17529 (N_17529,N_11392,N_12514);
xor U17530 (N_17530,N_12923,N_14116);
nor U17531 (N_17531,N_10199,N_13770);
xnor U17532 (N_17532,N_12001,N_11112);
xnor U17533 (N_17533,N_11606,N_12113);
nor U17534 (N_17534,N_11485,N_13773);
or U17535 (N_17535,N_14945,N_13107);
xor U17536 (N_17536,N_10419,N_10246);
nor U17537 (N_17537,N_10224,N_13104);
and U17538 (N_17538,N_10381,N_11166);
nor U17539 (N_17539,N_14737,N_14040);
and U17540 (N_17540,N_11663,N_10568);
nand U17541 (N_17541,N_11546,N_11575);
or U17542 (N_17542,N_10323,N_11457);
nor U17543 (N_17543,N_12998,N_12704);
and U17544 (N_17544,N_12805,N_13808);
and U17545 (N_17545,N_13779,N_13760);
xor U17546 (N_17546,N_11521,N_14223);
xor U17547 (N_17547,N_10819,N_14285);
and U17548 (N_17548,N_14358,N_12337);
or U17549 (N_17549,N_12070,N_10178);
and U17550 (N_17550,N_13253,N_11677);
nand U17551 (N_17551,N_13349,N_13773);
and U17552 (N_17552,N_10987,N_14814);
or U17553 (N_17553,N_13291,N_12055);
xnor U17554 (N_17554,N_11340,N_13171);
or U17555 (N_17555,N_11406,N_12611);
nand U17556 (N_17556,N_11558,N_13279);
xor U17557 (N_17557,N_12049,N_11763);
nor U17558 (N_17558,N_11468,N_13029);
or U17559 (N_17559,N_12791,N_10138);
xor U17560 (N_17560,N_14605,N_10876);
or U17561 (N_17561,N_12018,N_11505);
and U17562 (N_17562,N_14854,N_14217);
nor U17563 (N_17563,N_12838,N_13349);
nor U17564 (N_17564,N_14584,N_11238);
xor U17565 (N_17565,N_12988,N_14240);
nand U17566 (N_17566,N_11832,N_14167);
nor U17567 (N_17567,N_14707,N_11433);
or U17568 (N_17568,N_11971,N_14354);
xor U17569 (N_17569,N_10934,N_11803);
nor U17570 (N_17570,N_14201,N_12146);
and U17571 (N_17571,N_13684,N_10393);
or U17572 (N_17572,N_14781,N_11750);
nor U17573 (N_17573,N_11090,N_10079);
xnor U17574 (N_17574,N_13917,N_13166);
or U17575 (N_17575,N_13435,N_14785);
and U17576 (N_17576,N_12032,N_11012);
or U17577 (N_17577,N_10221,N_11431);
xnor U17578 (N_17578,N_14844,N_14514);
nor U17579 (N_17579,N_11253,N_14072);
nand U17580 (N_17580,N_11990,N_12606);
and U17581 (N_17581,N_13663,N_13175);
nor U17582 (N_17582,N_11546,N_10630);
nor U17583 (N_17583,N_11846,N_11686);
and U17584 (N_17584,N_10024,N_12459);
nand U17585 (N_17585,N_14128,N_12257);
and U17586 (N_17586,N_12159,N_11899);
and U17587 (N_17587,N_10068,N_13860);
and U17588 (N_17588,N_14639,N_14287);
nor U17589 (N_17589,N_12621,N_12588);
nor U17590 (N_17590,N_14796,N_14371);
xnor U17591 (N_17591,N_13622,N_11292);
nor U17592 (N_17592,N_10891,N_12223);
or U17593 (N_17593,N_10450,N_13250);
xor U17594 (N_17594,N_13580,N_14091);
nand U17595 (N_17595,N_14228,N_11392);
nand U17596 (N_17596,N_13941,N_14790);
and U17597 (N_17597,N_12434,N_14073);
and U17598 (N_17598,N_12305,N_11770);
nor U17599 (N_17599,N_14218,N_10044);
and U17600 (N_17600,N_13098,N_12992);
nor U17601 (N_17601,N_11035,N_11100);
or U17602 (N_17602,N_10152,N_13825);
nor U17603 (N_17603,N_13189,N_11258);
nor U17604 (N_17604,N_10789,N_12645);
and U17605 (N_17605,N_13274,N_11608);
xor U17606 (N_17606,N_12693,N_11565);
nand U17607 (N_17607,N_10246,N_13917);
xnor U17608 (N_17608,N_10526,N_10432);
nor U17609 (N_17609,N_13006,N_10375);
xnor U17610 (N_17610,N_11687,N_12289);
or U17611 (N_17611,N_13151,N_11317);
nor U17612 (N_17612,N_14369,N_11205);
xnor U17613 (N_17613,N_14189,N_12153);
and U17614 (N_17614,N_14441,N_11780);
or U17615 (N_17615,N_10161,N_10210);
nor U17616 (N_17616,N_14215,N_14241);
and U17617 (N_17617,N_10484,N_13029);
nand U17618 (N_17618,N_13463,N_10265);
xnor U17619 (N_17619,N_11991,N_10435);
nor U17620 (N_17620,N_11752,N_11155);
or U17621 (N_17621,N_14844,N_12044);
nor U17622 (N_17622,N_14231,N_13457);
and U17623 (N_17623,N_12120,N_10268);
xnor U17624 (N_17624,N_10868,N_13278);
or U17625 (N_17625,N_12370,N_11340);
nor U17626 (N_17626,N_10499,N_12563);
xor U17627 (N_17627,N_14592,N_13266);
nor U17628 (N_17628,N_14261,N_14417);
xnor U17629 (N_17629,N_12780,N_12560);
or U17630 (N_17630,N_13646,N_11346);
and U17631 (N_17631,N_11347,N_11370);
or U17632 (N_17632,N_13009,N_11084);
xor U17633 (N_17633,N_14583,N_10503);
nor U17634 (N_17634,N_11915,N_11236);
or U17635 (N_17635,N_11111,N_13718);
nor U17636 (N_17636,N_10889,N_10668);
or U17637 (N_17637,N_13802,N_11363);
and U17638 (N_17638,N_13388,N_11219);
and U17639 (N_17639,N_11694,N_10856);
or U17640 (N_17640,N_11900,N_10592);
or U17641 (N_17641,N_11693,N_13918);
or U17642 (N_17642,N_12468,N_10151);
or U17643 (N_17643,N_10698,N_12253);
xor U17644 (N_17644,N_11192,N_14870);
nand U17645 (N_17645,N_14725,N_12258);
or U17646 (N_17646,N_13008,N_10879);
and U17647 (N_17647,N_10209,N_12434);
nor U17648 (N_17648,N_12873,N_14914);
xnor U17649 (N_17649,N_14510,N_11785);
nand U17650 (N_17650,N_14054,N_11185);
nor U17651 (N_17651,N_12125,N_10437);
xor U17652 (N_17652,N_12315,N_11041);
nor U17653 (N_17653,N_14306,N_14403);
nor U17654 (N_17654,N_10002,N_12544);
and U17655 (N_17655,N_11194,N_10633);
xor U17656 (N_17656,N_11478,N_11502);
nor U17657 (N_17657,N_10742,N_13699);
nand U17658 (N_17658,N_13448,N_13009);
and U17659 (N_17659,N_10202,N_11752);
nand U17660 (N_17660,N_12836,N_10071);
nand U17661 (N_17661,N_10062,N_13973);
or U17662 (N_17662,N_10954,N_13125);
xnor U17663 (N_17663,N_12540,N_11120);
or U17664 (N_17664,N_14626,N_10740);
nor U17665 (N_17665,N_14908,N_13146);
nand U17666 (N_17666,N_14900,N_10945);
xnor U17667 (N_17667,N_12991,N_13853);
nor U17668 (N_17668,N_14262,N_10856);
and U17669 (N_17669,N_11886,N_10740);
or U17670 (N_17670,N_14493,N_12832);
or U17671 (N_17671,N_13698,N_12495);
nand U17672 (N_17672,N_13059,N_10070);
and U17673 (N_17673,N_10632,N_14707);
or U17674 (N_17674,N_14951,N_11155);
xor U17675 (N_17675,N_11571,N_14140);
and U17676 (N_17676,N_12326,N_12637);
or U17677 (N_17677,N_11869,N_13768);
or U17678 (N_17678,N_12821,N_14233);
xor U17679 (N_17679,N_10210,N_13949);
and U17680 (N_17680,N_11052,N_13104);
nand U17681 (N_17681,N_11670,N_13360);
xor U17682 (N_17682,N_11542,N_14956);
nand U17683 (N_17683,N_13650,N_12762);
and U17684 (N_17684,N_10211,N_14494);
nor U17685 (N_17685,N_10309,N_11904);
nand U17686 (N_17686,N_11761,N_10363);
nand U17687 (N_17687,N_10614,N_12765);
xnor U17688 (N_17688,N_12387,N_10278);
nand U17689 (N_17689,N_13195,N_10418);
nand U17690 (N_17690,N_11907,N_10686);
xor U17691 (N_17691,N_11343,N_14723);
nand U17692 (N_17692,N_14642,N_12960);
nor U17693 (N_17693,N_14899,N_10096);
nor U17694 (N_17694,N_13870,N_10043);
or U17695 (N_17695,N_14683,N_12554);
or U17696 (N_17696,N_11559,N_10496);
nand U17697 (N_17697,N_10921,N_12839);
and U17698 (N_17698,N_13819,N_11883);
xor U17699 (N_17699,N_11311,N_12586);
or U17700 (N_17700,N_12237,N_11178);
or U17701 (N_17701,N_14106,N_14718);
xor U17702 (N_17702,N_14390,N_12414);
and U17703 (N_17703,N_13357,N_13255);
or U17704 (N_17704,N_14940,N_14658);
and U17705 (N_17705,N_10489,N_14020);
or U17706 (N_17706,N_13535,N_11652);
or U17707 (N_17707,N_14658,N_10424);
xor U17708 (N_17708,N_10237,N_10223);
nand U17709 (N_17709,N_14605,N_10888);
nor U17710 (N_17710,N_13854,N_14597);
xor U17711 (N_17711,N_14071,N_13215);
and U17712 (N_17712,N_12235,N_13437);
and U17713 (N_17713,N_11600,N_10557);
xnor U17714 (N_17714,N_10565,N_10237);
xnor U17715 (N_17715,N_10902,N_14932);
nand U17716 (N_17716,N_14513,N_11677);
and U17717 (N_17717,N_10998,N_10272);
or U17718 (N_17718,N_14941,N_10284);
nor U17719 (N_17719,N_12199,N_12121);
nand U17720 (N_17720,N_14366,N_11326);
nand U17721 (N_17721,N_10891,N_14599);
and U17722 (N_17722,N_14216,N_14008);
and U17723 (N_17723,N_11910,N_12483);
and U17724 (N_17724,N_14151,N_12105);
or U17725 (N_17725,N_12233,N_14998);
nand U17726 (N_17726,N_10398,N_12306);
and U17727 (N_17727,N_14768,N_11310);
nor U17728 (N_17728,N_11263,N_11041);
and U17729 (N_17729,N_14997,N_10255);
nand U17730 (N_17730,N_10978,N_11845);
and U17731 (N_17731,N_13589,N_11494);
or U17732 (N_17732,N_13412,N_10790);
xor U17733 (N_17733,N_11062,N_12757);
nor U17734 (N_17734,N_13868,N_12518);
or U17735 (N_17735,N_10022,N_14601);
and U17736 (N_17736,N_12219,N_12964);
or U17737 (N_17737,N_14119,N_12581);
nor U17738 (N_17738,N_13669,N_11532);
xnor U17739 (N_17739,N_11440,N_10445);
nor U17740 (N_17740,N_11482,N_12765);
nand U17741 (N_17741,N_14353,N_14413);
or U17742 (N_17742,N_10298,N_10667);
nor U17743 (N_17743,N_10097,N_12531);
xnor U17744 (N_17744,N_11617,N_10011);
xnor U17745 (N_17745,N_14986,N_11651);
nor U17746 (N_17746,N_13932,N_11599);
xnor U17747 (N_17747,N_11887,N_14825);
nand U17748 (N_17748,N_13973,N_13717);
xnor U17749 (N_17749,N_10878,N_13799);
nand U17750 (N_17750,N_11225,N_12824);
and U17751 (N_17751,N_12076,N_11260);
nand U17752 (N_17752,N_13896,N_13973);
xor U17753 (N_17753,N_10970,N_11825);
xor U17754 (N_17754,N_11765,N_11921);
xnor U17755 (N_17755,N_10551,N_11510);
nand U17756 (N_17756,N_10366,N_13349);
nand U17757 (N_17757,N_11829,N_10520);
nor U17758 (N_17758,N_14309,N_12269);
or U17759 (N_17759,N_11370,N_12112);
nand U17760 (N_17760,N_12442,N_10080);
xnor U17761 (N_17761,N_10764,N_13027);
nand U17762 (N_17762,N_10414,N_11495);
or U17763 (N_17763,N_14310,N_10180);
nand U17764 (N_17764,N_13109,N_11467);
nor U17765 (N_17765,N_12397,N_10626);
nand U17766 (N_17766,N_12639,N_12467);
nor U17767 (N_17767,N_12004,N_11100);
and U17768 (N_17768,N_14050,N_10575);
and U17769 (N_17769,N_14798,N_11032);
nor U17770 (N_17770,N_13357,N_13825);
nand U17771 (N_17771,N_14208,N_14403);
xor U17772 (N_17772,N_12167,N_11463);
xor U17773 (N_17773,N_11833,N_13800);
xnor U17774 (N_17774,N_10157,N_13853);
xor U17775 (N_17775,N_10861,N_14949);
or U17776 (N_17776,N_10103,N_12841);
xor U17777 (N_17777,N_12484,N_12843);
and U17778 (N_17778,N_13072,N_14637);
nor U17779 (N_17779,N_12543,N_10041);
and U17780 (N_17780,N_12789,N_12078);
or U17781 (N_17781,N_13473,N_11784);
xnor U17782 (N_17782,N_10850,N_10169);
or U17783 (N_17783,N_11699,N_10968);
or U17784 (N_17784,N_13436,N_13625);
nand U17785 (N_17785,N_14797,N_10658);
nand U17786 (N_17786,N_10333,N_14921);
nand U17787 (N_17787,N_11424,N_13393);
nand U17788 (N_17788,N_14210,N_12993);
or U17789 (N_17789,N_11867,N_14121);
or U17790 (N_17790,N_14277,N_14457);
nand U17791 (N_17791,N_10176,N_11456);
nor U17792 (N_17792,N_11997,N_10366);
nand U17793 (N_17793,N_14125,N_14461);
nor U17794 (N_17794,N_11111,N_14371);
nor U17795 (N_17795,N_12766,N_13769);
nand U17796 (N_17796,N_12071,N_12900);
or U17797 (N_17797,N_12730,N_13013);
nor U17798 (N_17798,N_10594,N_12578);
or U17799 (N_17799,N_14338,N_11084);
and U17800 (N_17800,N_10945,N_12946);
and U17801 (N_17801,N_11194,N_10465);
nor U17802 (N_17802,N_11514,N_11407);
and U17803 (N_17803,N_11922,N_14352);
xnor U17804 (N_17804,N_10274,N_12849);
and U17805 (N_17805,N_10998,N_13547);
xnor U17806 (N_17806,N_11907,N_12771);
and U17807 (N_17807,N_14072,N_12288);
or U17808 (N_17808,N_11308,N_11524);
and U17809 (N_17809,N_14281,N_10058);
or U17810 (N_17810,N_14148,N_13722);
xnor U17811 (N_17811,N_12183,N_12942);
nor U17812 (N_17812,N_11691,N_12991);
xor U17813 (N_17813,N_13666,N_14574);
and U17814 (N_17814,N_13317,N_11806);
nand U17815 (N_17815,N_11376,N_14821);
xor U17816 (N_17816,N_11840,N_13695);
and U17817 (N_17817,N_13293,N_12613);
xnor U17818 (N_17818,N_14174,N_10390);
and U17819 (N_17819,N_11940,N_10018);
nor U17820 (N_17820,N_11436,N_12300);
nand U17821 (N_17821,N_13842,N_11958);
nand U17822 (N_17822,N_11090,N_11594);
xor U17823 (N_17823,N_14390,N_10326);
and U17824 (N_17824,N_12550,N_13274);
nor U17825 (N_17825,N_11628,N_11007);
and U17826 (N_17826,N_12517,N_10877);
nand U17827 (N_17827,N_13019,N_14471);
nor U17828 (N_17828,N_11752,N_11182);
and U17829 (N_17829,N_11072,N_14202);
xnor U17830 (N_17830,N_12412,N_13655);
xnor U17831 (N_17831,N_10190,N_13161);
nor U17832 (N_17832,N_12706,N_10121);
or U17833 (N_17833,N_12785,N_14083);
or U17834 (N_17834,N_14579,N_14509);
nor U17835 (N_17835,N_11607,N_12920);
xor U17836 (N_17836,N_11369,N_10365);
nand U17837 (N_17837,N_11155,N_10227);
or U17838 (N_17838,N_13287,N_10607);
and U17839 (N_17839,N_10776,N_10421);
or U17840 (N_17840,N_13245,N_13096);
nand U17841 (N_17841,N_14435,N_12743);
nand U17842 (N_17842,N_11780,N_14312);
nand U17843 (N_17843,N_13196,N_11214);
nand U17844 (N_17844,N_14211,N_11372);
or U17845 (N_17845,N_12852,N_13799);
xnor U17846 (N_17846,N_14283,N_10124);
xnor U17847 (N_17847,N_14601,N_10130);
nand U17848 (N_17848,N_14560,N_10075);
nand U17849 (N_17849,N_13840,N_11878);
nand U17850 (N_17850,N_11152,N_12154);
nand U17851 (N_17851,N_14400,N_12889);
nor U17852 (N_17852,N_12996,N_12434);
xnor U17853 (N_17853,N_12210,N_14597);
or U17854 (N_17854,N_10090,N_14532);
or U17855 (N_17855,N_10121,N_10606);
nand U17856 (N_17856,N_10176,N_11015);
or U17857 (N_17857,N_14993,N_11153);
nand U17858 (N_17858,N_12752,N_11202);
nand U17859 (N_17859,N_12728,N_13847);
xor U17860 (N_17860,N_11194,N_14732);
nor U17861 (N_17861,N_14302,N_11942);
nand U17862 (N_17862,N_10800,N_11647);
nor U17863 (N_17863,N_10798,N_12688);
and U17864 (N_17864,N_10206,N_11294);
and U17865 (N_17865,N_12938,N_12627);
nand U17866 (N_17866,N_12281,N_13565);
nand U17867 (N_17867,N_10851,N_11071);
and U17868 (N_17868,N_14560,N_10246);
and U17869 (N_17869,N_10484,N_11852);
nand U17870 (N_17870,N_14191,N_10443);
xnor U17871 (N_17871,N_11688,N_10051);
nand U17872 (N_17872,N_13122,N_14081);
and U17873 (N_17873,N_14838,N_13398);
xnor U17874 (N_17874,N_12944,N_13576);
and U17875 (N_17875,N_12401,N_11809);
nand U17876 (N_17876,N_11692,N_10493);
or U17877 (N_17877,N_14869,N_12443);
or U17878 (N_17878,N_14551,N_13569);
nor U17879 (N_17879,N_13536,N_10490);
nor U17880 (N_17880,N_11440,N_14732);
nor U17881 (N_17881,N_10396,N_14331);
or U17882 (N_17882,N_13980,N_10370);
and U17883 (N_17883,N_13568,N_10730);
nor U17884 (N_17884,N_14227,N_14946);
or U17885 (N_17885,N_12136,N_12519);
nor U17886 (N_17886,N_12807,N_11706);
and U17887 (N_17887,N_12916,N_13480);
nor U17888 (N_17888,N_14859,N_14468);
nand U17889 (N_17889,N_10634,N_10455);
or U17890 (N_17890,N_14709,N_12942);
xor U17891 (N_17891,N_11025,N_13895);
or U17892 (N_17892,N_11624,N_11924);
nand U17893 (N_17893,N_10841,N_13933);
nand U17894 (N_17894,N_11077,N_13583);
nand U17895 (N_17895,N_10363,N_13398);
or U17896 (N_17896,N_12586,N_11892);
nor U17897 (N_17897,N_12607,N_10183);
nand U17898 (N_17898,N_14377,N_13944);
nand U17899 (N_17899,N_13611,N_14780);
nand U17900 (N_17900,N_11505,N_10617);
and U17901 (N_17901,N_11716,N_11798);
nor U17902 (N_17902,N_13643,N_13943);
xor U17903 (N_17903,N_11806,N_10238);
and U17904 (N_17904,N_13516,N_14786);
or U17905 (N_17905,N_13990,N_11618);
and U17906 (N_17906,N_11675,N_10956);
nor U17907 (N_17907,N_12665,N_13928);
xor U17908 (N_17908,N_12064,N_11444);
nand U17909 (N_17909,N_14630,N_11751);
nor U17910 (N_17910,N_13791,N_12132);
or U17911 (N_17911,N_14609,N_14305);
nor U17912 (N_17912,N_12623,N_14996);
and U17913 (N_17913,N_12237,N_12268);
nand U17914 (N_17914,N_13958,N_14131);
xor U17915 (N_17915,N_11121,N_11879);
nand U17916 (N_17916,N_11159,N_12410);
xor U17917 (N_17917,N_10300,N_14360);
xor U17918 (N_17918,N_12698,N_14816);
nand U17919 (N_17919,N_13403,N_11561);
nand U17920 (N_17920,N_10680,N_12143);
nor U17921 (N_17921,N_10470,N_14687);
nor U17922 (N_17922,N_10122,N_11585);
nor U17923 (N_17923,N_14429,N_11161);
xnor U17924 (N_17924,N_14629,N_13583);
xnor U17925 (N_17925,N_14513,N_11476);
nand U17926 (N_17926,N_12965,N_12997);
xnor U17927 (N_17927,N_13046,N_10762);
and U17928 (N_17928,N_13852,N_13721);
nand U17929 (N_17929,N_13719,N_11853);
nand U17930 (N_17930,N_11401,N_10531);
xnor U17931 (N_17931,N_10442,N_11452);
or U17932 (N_17932,N_12383,N_12501);
nand U17933 (N_17933,N_14827,N_12700);
and U17934 (N_17934,N_10770,N_13407);
or U17935 (N_17935,N_12699,N_13358);
xnor U17936 (N_17936,N_12930,N_13631);
nor U17937 (N_17937,N_14066,N_12762);
or U17938 (N_17938,N_11862,N_11356);
and U17939 (N_17939,N_14712,N_11816);
or U17940 (N_17940,N_11634,N_11190);
and U17941 (N_17941,N_14721,N_12191);
and U17942 (N_17942,N_12508,N_10039);
nand U17943 (N_17943,N_11922,N_10941);
nand U17944 (N_17944,N_10779,N_10334);
nor U17945 (N_17945,N_14166,N_14806);
nor U17946 (N_17946,N_12445,N_11295);
and U17947 (N_17947,N_10492,N_12872);
nand U17948 (N_17948,N_10603,N_13435);
nor U17949 (N_17949,N_11675,N_12961);
or U17950 (N_17950,N_10390,N_12962);
and U17951 (N_17951,N_12283,N_11925);
nor U17952 (N_17952,N_11379,N_11072);
xor U17953 (N_17953,N_14664,N_11237);
nand U17954 (N_17954,N_14650,N_11001);
or U17955 (N_17955,N_13403,N_14244);
xor U17956 (N_17956,N_11425,N_10758);
or U17957 (N_17957,N_12194,N_12974);
nor U17958 (N_17958,N_14895,N_13598);
or U17959 (N_17959,N_13452,N_14001);
nor U17960 (N_17960,N_10223,N_14045);
nand U17961 (N_17961,N_10955,N_11057);
nor U17962 (N_17962,N_10481,N_12606);
and U17963 (N_17963,N_14522,N_14817);
nor U17964 (N_17964,N_11574,N_12396);
nor U17965 (N_17965,N_13680,N_10270);
nand U17966 (N_17966,N_14292,N_14142);
nand U17967 (N_17967,N_12677,N_10943);
xnor U17968 (N_17968,N_11063,N_12701);
nand U17969 (N_17969,N_13364,N_14557);
xor U17970 (N_17970,N_13797,N_11108);
nor U17971 (N_17971,N_14174,N_10916);
or U17972 (N_17972,N_11639,N_11476);
nor U17973 (N_17973,N_13346,N_11059);
and U17974 (N_17974,N_13802,N_14846);
or U17975 (N_17975,N_12341,N_11802);
xor U17976 (N_17976,N_10220,N_13013);
nor U17977 (N_17977,N_13896,N_11373);
nor U17978 (N_17978,N_11287,N_13098);
xor U17979 (N_17979,N_13114,N_13507);
and U17980 (N_17980,N_12641,N_11785);
and U17981 (N_17981,N_12833,N_10615);
or U17982 (N_17982,N_13835,N_11991);
xor U17983 (N_17983,N_10131,N_13420);
xnor U17984 (N_17984,N_10178,N_11623);
nand U17985 (N_17985,N_14634,N_12865);
nor U17986 (N_17986,N_11977,N_10498);
nand U17987 (N_17987,N_13838,N_12169);
nand U17988 (N_17988,N_10456,N_13639);
or U17989 (N_17989,N_11958,N_11714);
nor U17990 (N_17990,N_12557,N_13080);
and U17991 (N_17991,N_12236,N_11949);
nand U17992 (N_17992,N_13038,N_11639);
nand U17993 (N_17993,N_11323,N_13932);
nor U17994 (N_17994,N_11532,N_13204);
and U17995 (N_17995,N_13384,N_10421);
xnor U17996 (N_17996,N_14841,N_14787);
nor U17997 (N_17997,N_11307,N_12961);
nand U17998 (N_17998,N_11394,N_10704);
xnor U17999 (N_17999,N_14153,N_10935);
xnor U18000 (N_18000,N_13401,N_11835);
xor U18001 (N_18001,N_11863,N_13286);
xor U18002 (N_18002,N_11872,N_12274);
or U18003 (N_18003,N_11375,N_14133);
xor U18004 (N_18004,N_10124,N_14189);
nand U18005 (N_18005,N_14351,N_13290);
and U18006 (N_18006,N_12502,N_10414);
nand U18007 (N_18007,N_13293,N_10733);
or U18008 (N_18008,N_14705,N_14064);
nor U18009 (N_18009,N_11804,N_14608);
or U18010 (N_18010,N_13084,N_11646);
nand U18011 (N_18011,N_11548,N_12604);
or U18012 (N_18012,N_11622,N_13055);
and U18013 (N_18013,N_14598,N_11637);
nor U18014 (N_18014,N_13648,N_14437);
and U18015 (N_18015,N_10018,N_12569);
or U18016 (N_18016,N_14214,N_14274);
xnor U18017 (N_18017,N_11777,N_12693);
nand U18018 (N_18018,N_11971,N_13376);
nor U18019 (N_18019,N_11787,N_13505);
nor U18020 (N_18020,N_13946,N_13275);
nor U18021 (N_18021,N_11493,N_12154);
nor U18022 (N_18022,N_14060,N_12024);
and U18023 (N_18023,N_12514,N_13335);
nand U18024 (N_18024,N_13404,N_11548);
and U18025 (N_18025,N_14724,N_10056);
nand U18026 (N_18026,N_10691,N_10238);
and U18027 (N_18027,N_12071,N_14090);
nor U18028 (N_18028,N_11110,N_10207);
nand U18029 (N_18029,N_14192,N_14644);
or U18030 (N_18030,N_11177,N_13748);
or U18031 (N_18031,N_10837,N_14401);
nor U18032 (N_18032,N_14860,N_10292);
nand U18033 (N_18033,N_10939,N_13829);
and U18034 (N_18034,N_12742,N_14099);
and U18035 (N_18035,N_11380,N_14087);
nand U18036 (N_18036,N_13378,N_13657);
nor U18037 (N_18037,N_10505,N_10523);
and U18038 (N_18038,N_10844,N_12554);
nand U18039 (N_18039,N_10821,N_14391);
and U18040 (N_18040,N_14004,N_13628);
and U18041 (N_18041,N_10383,N_12577);
nand U18042 (N_18042,N_10058,N_11737);
xnor U18043 (N_18043,N_14251,N_13447);
xor U18044 (N_18044,N_12170,N_13815);
nor U18045 (N_18045,N_12915,N_12653);
xnor U18046 (N_18046,N_13533,N_13944);
xor U18047 (N_18047,N_10076,N_12406);
and U18048 (N_18048,N_14812,N_10465);
nand U18049 (N_18049,N_11241,N_12904);
nand U18050 (N_18050,N_10901,N_12033);
xnor U18051 (N_18051,N_13832,N_13514);
nand U18052 (N_18052,N_12555,N_10631);
nand U18053 (N_18053,N_10512,N_14109);
nor U18054 (N_18054,N_12146,N_13116);
nor U18055 (N_18055,N_14982,N_11599);
or U18056 (N_18056,N_14128,N_13871);
xnor U18057 (N_18057,N_14570,N_11766);
nor U18058 (N_18058,N_13057,N_10459);
and U18059 (N_18059,N_14451,N_13353);
and U18060 (N_18060,N_10965,N_14743);
or U18061 (N_18061,N_12603,N_14742);
nor U18062 (N_18062,N_14224,N_10605);
and U18063 (N_18063,N_14375,N_14630);
or U18064 (N_18064,N_14577,N_14231);
or U18065 (N_18065,N_11580,N_10472);
nor U18066 (N_18066,N_14981,N_11194);
nor U18067 (N_18067,N_13847,N_12684);
nand U18068 (N_18068,N_11160,N_13069);
xnor U18069 (N_18069,N_10279,N_12297);
and U18070 (N_18070,N_12820,N_12935);
nand U18071 (N_18071,N_11597,N_12839);
nor U18072 (N_18072,N_14052,N_14709);
or U18073 (N_18073,N_13674,N_11907);
xor U18074 (N_18074,N_13052,N_11160);
and U18075 (N_18075,N_11085,N_12475);
xor U18076 (N_18076,N_13965,N_14336);
xor U18077 (N_18077,N_12928,N_13166);
xor U18078 (N_18078,N_10196,N_10414);
or U18079 (N_18079,N_13911,N_11821);
nand U18080 (N_18080,N_12041,N_10486);
nand U18081 (N_18081,N_13217,N_14084);
nor U18082 (N_18082,N_14633,N_10337);
and U18083 (N_18083,N_14538,N_11139);
xor U18084 (N_18084,N_11535,N_10707);
nor U18085 (N_18085,N_14398,N_14476);
nor U18086 (N_18086,N_14175,N_11841);
or U18087 (N_18087,N_10169,N_10560);
or U18088 (N_18088,N_13756,N_14151);
xor U18089 (N_18089,N_12178,N_13474);
and U18090 (N_18090,N_10249,N_12062);
nor U18091 (N_18091,N_11616,N_10196);
xnor U18092 (N_18092,N_11825,N_14885);
xnor U18093 (N_18093,N_12129,N_11054);
or U18094 (N_18094,N_12005,N_12654);
or U18095 (N_18095,N_13810,N_12050);
xor U18096 (N_18096,N_11002,N_11282);
nor U18097 (N_18097,N_12542,N_13166);
xor U18098 (N_18098,N_11039,N_11999);
or U18099 (N_18099,N_11197,N_10398);
nor U18100 (N_18100,N_13524,N_11897);
and U18101 (N_18101,N_12035,N_13551);
and U18102 (N_18102,N_14971,N_13341);
or U18103 (N_18103,N_12140,N_10776);
and U18104 (N_18104,N_14235,N_12246);
nor U18105 (N_18105,N_12727,N_12068);
or U18106 (N_18106,N_12701,N_13452);
or U18107 (N_18107,N_14375,N_14215);
nand U18108 (N_18108,N_10783,N_10729);
and U18109 (N_18109,N_11337,N_11670);
nand U18110 (N_18110,N_10771,N_13788);
and U18111 (N_18111,N_11327,N_10441);
xor U18112 (N_18112,N_11630,N_12456);
xnor U18113 (N_18113,N_14473,N_12151);
xor U18114 (N_18114,N_13419,N_14901);
xor U18115 (N_18115,N_13016,N_12170);
and U18116 (N_18116,N_14983,N_14241);
nor U18117 (N_18117,N_10310,N_13526);
nor U18118 (N_18118,N_13560,N_13756);
xor U18119 (N_18119,N_12189,N_11975);
or U18120 (N_18120,N_12601,N_11186);
nor U18121 (N_18121,N_14686,N_13512);
xor U18122 (N_18122,N_10757,N_11759);
nor U18123 (N_18123,N_11244,N_10849);
nor U18124 (N_18124,N_10509,N_11508);
and U18125 (N_18125,N_10713,N_13442);
nand U18126 (N_18126,N_14740,N_12894);
and U18127 (N_18127,N_11239,N_14973);
nor U18128 (N_18128,N_13429,N_14550);
xor U18129 (N_18129,N_13550,N_12155);
and U18130 (N_18130,N_13036,N_14387);
and U18131 (N_18131,N_14786,N_14622);
and U18132 (N_18132,N_13217,N_12439);
xor U18133 (N_18133,N_11373,N_14262);
or U18134 (N_18134,N_10026,N_10106);
or U18135 (N_18135,N_12291,N_13859);
and U18136 (N_18136,N_14060,N_14529);
nand U18137 (N_18137,N_11924,N_12267);
nand U18138 (N_18138,N_14019,N_11672);
nor U18139 (N_18139,N_12401,N_10320);
and U18140 (N_18140,N_12468,N_14948);
or U18141 (N_18141,N_13686,N_11056);
or U18142 (N_18142,N_13187,N_13410);
nand U18143 (N_18143,N_12289,N_12870);
xnor U18144 (N_18144,N_10162,N_13580);
and U18145 (N_18145,N_10138,N_12435);
nand U18146 (N_18146,N_11608,N_10104);
and U18147 (N_18147,N_12203,N_13628);
xnor U18148 (N_18148,N_10598,N_14041);
nor U18149 (N_18149,N_10942,N_11098);
nor U18150 (N_18150,N_14476,N_10955);
or U18151 (N_18151,N_13086,N_10190);
and U18152 (N_18152,N_11900,N_13086);
nand U18153 (N_18153,N_11974,N_12988);
nor U18154 (N_18154,N_10739,N_11273);
nand U18155 (N_18155,N_13981,N_12478);
nor U18156 (N_18156,N_11416,N_11196);
xor U18157 (N_18157,N_14055,N_12125);
xor U18158 (N_18158,N_11972,N_10916);
xor U18159 (N_18159,N_13714,N_10743);
or U18160 (N_18160,N_14739,N_13506);
nand U18161 (N_18161,N_10978,N_12241);
and U18162 (N_18162,N_14143,N_13859);
xnor U18163 (N_18163,N_11135,N_10317);
nand U18164 (N_18164,N_13828,N_13111);
nand U18165 (N_18165,N_10680,N_12902);
xor U18166 (N_18166,N_14430,N_12426);
nor U18167 (N_18167,N_11011,N_10660);
nor U18168 (N_18168,N_13560,N_10268);
or U18169 (N_18169,N_12453,N_13923);
xor U18170 (N_18170,N_10815,N_11508);
and U18171 (N_18171,N_13797,N_14113);
nand U18172 (N_18172,N_10796,N_13502);
xnor U18173 (N_18173,N_12976,N_11194);
xor U18174 (N_18174,N_13430,N_10793);
or U18175 (N_18175,N_11079,N_13011);
or U18176 (N_18176,N_14581,N_10407);
xnor U18177 (N_18177,N_13055,N_11613);
nor U18178 (N_18178,N_11444,N_12339);
or U18179 (N_18179,N_14900,N_10873);
nor U18180 (N_18180,N_10734,N_13382);
or U18181 (N_18181,N_12824,N_13241);
or U18182 (N_18182,N_13994,N_13298);
nor U18183 (N_18183,N_10149,N_10592);
nand U18184 (N_18184,N_14021,N_11031);
nand U18185 (N_18185,N_13879,N_12447);
and U18186 (N_18186,N_12739,N_13468);
nand U18187 (N_18187,N_11072,N_12215);
and U18188 (N_18188,N_14928,N_10224);
and U18189 (N_18189,N_14463,N_11262);
xnor U18190 (N_18190,N_12101,N_12603);
xor U18191 (N_18191,N_12991,N_11206);
nor U18192 (N_18192,N_13894,N_12073);
and U18193 (N_18193,N_12236,N_10104);
nand U18194 (N_18194,N_12331,N_11943);
xor U18195 (N_18195,N_13294,N_11122);
or U18196 (N_18196,N_14752,N_14877);
or U18197 (N_18197,N_13135,N_14017);
xnor U18198 (N_18198,N_13396,N_14013);
xor U18199 (N_18199,N_10386,N_11138);
nand U18200 (N_18200,N_14652,N_13526);
and U18201 (N_18201,N_10093,N_10794);
nand U18202 (N_18202,N_12599,N_11486);
nand U18203 (N_18203,N_12597,N_11807);
nand U18204 (N_18204,N_14058,N_14755);
nor U18205 (N_18205,N_13057,N_11507);
nand U18206 (N_18206,N_13945,N_11876);
or U18207 (N_18207,N_12864,N_11179);
or U18208 (N_18208,N_14947,N_10310);
or U18209 (N_18209,N_11452,N_11640);
nand U18210 (N_18210,N_14364,N_14628);
nand U18211 (N_18211,N_10384,N_12306);
and U18212 (N_18212,N_12521,N_13625);
nor U18213 (N_18213,N_14940,N_12829);
nor U18214 (N_18214,N_13598,N_14657);
nor U18215 (N_18215,N_14489,N_10190);
nor U18216 (N_18216,N_13815,N_14024);
nand U18217 (N_18217,N_13599,N_11430);
nor U18218 (N_18218,N_11094,N_13992);
nand U18219 (N_18219,N_11042,N_12374);
or U18220 (N_18220,N_13024,N_12412);
xnor U18221 (N_18221,N_14083,N_14460);
or U18222 (N_18222,N_13961,N_10910);
and U18223 (N_18223,N_14279,N_11032);
nand U18224 (N_18224,N_12302,N_14209);
nand U18225 (N_18225,N_11680,N_10523);
and U18226 (N_18226,N_13793,N_13771);
nand U18227 (N_18227,N_13491,N_13055);
nor U18228 (N_18228,N_11102,N_13094);
or U18229 (N_18229,N_14410,N_11391);
nand U18230 (N_18230,N_10616,N_14285);
nor U18231 (N_18231,N_13000,N_14642);
and U18232 (N_18232,N_11983,N_14251);
or U18233 (N_18233,N_10264,N_13825);
nor U18234 (N_18234,N_11673,N_14701);
or U18235 (N_18235,N_13059,N_10409);
or U18236 (N_18236,N_14607,N_10196);
nor U18237 (N_18237,N_10283,N_10172);
nand U18238 (N_18238,N_11019,N_10897);
xor U18239 (N_18239,N_12951,N_11766);
xor U18240 (N_18240,N_10957,N_10595);
or U18241 (N_18241,N_13359,N_11978);
nor U18242 (N_18242,N_10575,N_12862);
nor U18243 (N_18243,N_14925,N_13253);
xnor U18244 (N_18244,N_10644,N_14329);
nor U18245 (N_18245,N_13515,N_13858);
nand U18246 (N_18246,N_14087,N_10486);
and U18247 (N_18247,N_10588,N_10685);
or U18248 (N_18248,N_11156,N_14049);
nor U18249 (N_18249,N_13620,N_13192);
nand U18250 (N_18250,N_13587,N_12604);
nor U18251 (N_18251,N_13795,N_10691);
nor U18252 (N_18252,N_11359,N_11136);
xor U18253 (N_18253,N_11765,N_10847);
xnor U18254 (N_18254,N_10883,N_12740);
and U18255 (N_18255,N_10561,N_10790);
nand U18256 (N_18256,N_14237,N_10306);
nand U18257 (N_18257,N_11926,N_13804);
nand U18258 (N_18258,N_11195,N_11780);
or U18259 (N_18259,N_12341,N_14771);
nand U18260 (N_18260,N_12098,N_13958);
nand U18261 (N_18261,N_12060,N_10489);
and U18262 (N_18262,N_11589,N_11032);
or U18263 (N_18263,N_13553,N_13340);
nand U18264 (N_18264,N_14287,N_11984);
or U18265 (N_18265,N_11857,N_11293);
nor U18266 (N_18266,N_12743,N_14044);
nor U18267 (N_18267,N_14917,N_11796);
xnor U18268 (N_18268,N_14867,N_11939);
or U18269 (N_18269,N_14026,N_13615);
nand U18270 (N_18270,N_11258,N_10987);
nand U18271 (N_18271,N_12189,N_12115);
or U18272 (N_18272,N_12784,N_11372);
nand U18273 (N_18273,N_14416,N_13740);
nor U18274 (N_18274,N_10405,N_11827);
xor U18275 (N_18275,N_14640,N_10904);
or U18276 (N_18276,N_10447,N_14945);
xnor U18277 (N_18277,N_14162,N_10713);
nor U18278 (N_18278,N_14481,N_14691);
xor U18279 (N_18279,N_11742,N_11590);
nand U18280 (N_18280,N_13074,N_14355);
nand U18281 (N_18281,N_13715,N_10371);
nor U18282 (N_18282,N_13987,N_12015);
and U18283 (N_18283,N_12434,N_10233);
nand U18284 (N_18284,N_12119,N_13461);
or U18285 (N_18285,N_10668,N_14691);
or U18286 (N_18286,N_11286,N_11468);
or U18287 (N_18287,N_10559,N_12156);
nand U18288 (N_18288,N_10521,N_10144);
nand U18289 (N_18289,N_14487,N_10801);
or U18290 (N_18290,N_14037,N_10504);
xnor U18291 (N_18291,N_11716,N_14291);
nand U18292 (N_18292,N_14345,N_11713);
and U18293 (N_18293,N_12205,N_14548);
nor U18294 (N_18294,N_14460,N_11660);
nor U18295 (N_18295,N_13277,N_12944);
and U18296 (N_18296,N_10100,N_12161);
nand U18297 (N_18297,N_12980,N_11999);
or U18298 (N_18298,N_13800,N_14405);
xor U18299 (N_18299,N_13723,N_12715);
or U18300 (N_18300,N_12644,N_14275);
and U18301 (N_18301,N_11273,N_12640);
or U18302 (N_18302,N_13087,N_12476);
or U18303 (N_18303,N_13311,N_10405);
xor U18304 (N_18304,N_12111,N_13923);
nand U18305 (N_18305,N_11625,N_11685);
nand U18306 (N_18306,N_12680,N_14006);
xor U18307 (N_18307,N_11078,N_13899);
xor U18308 (N_18308,N_13623,N_13633);
or U18309 (N_18309,N_12522,N_12885);
nand U18310 (N_18310,N_14206,N_12731);
nand U18311 (N_18311,N_11074,N_13087);
nor U18312 (N_18312,N_13103,N_10305);
nand U18313 (N_18313,N_13894,N_12957);
and U18314 (N_18314,N_12909,N_13208);
or U18315 (N_18315,N_12747,N_10223);
nand U18316 (N_18316,N_13238,N_13381);
nand U18317 (N_18317,N_10138,N_11819);
and U18318 (N_18318,N_13733,N_11493);
nand U18319 (N_18319,N_11813,N_14754);
and U18320 (N_18320,N_11123,N_10415);
nand U18321 (N_18321,N_14574,N_12873);
xor U18322 (N_18322,N_10300,N_11951);
nand U18323 (N_18323,N_14295,N_10524);
xor U18324 (N_18324,N_14190,N_14472);
and U18325 (N_18325,N_14927,N_10678);
nor U18326 (N_18326,N_10252,N_12404);
and U18327 (N_18327,N_11050,N_13951);
or U18328 (N_18328,N_14342,N_14978);
nor U18329 (N_18329,N_10563,N_11628);
nand U18330 (N_18330,N_13936,N_11287);
or U18331 (N_18331,N_12843,N_11766);
and U18332 (N_18332,N_14722,N_11884);
nand U18333 (N_18333,N_10146,N_14621);
and U18334 (N_18334,N_11323,N_11896);
nand U18335 (N_18335,N_14278,N_14706);
and U18336 (N_18336,N_14984,N_10375);
or U18337 (N_18337,N_11619,N_14646);
and U18338 (N_18338,N_10318,N_12780);
or U18339 (N_18339,N_10719,N_13574);
or U18340 (N_18340,N_12422,N_12770);
nor U18341 (N_18341,N_13846,N_10730);
nand U18342 (N_18342,N_13766,N_12384);
nand U18343 (N_18343,N_10190,N_11424);
xnor U18344 (N_18344,N_10507,N_11915);
nand U18345 (N_18345,N_10936,N_12747);
or U18346 (N_18346,N_14389,N_13873);
or U18347 (N_18347,N_12289,N_13115);
nand U18348 (N_18348,N_11348,N_14621);
xnor U18349 (N_18349,N_14391,N_14773);
or U18350 (N_18350,N_12442,N_11835);
or U18351 (N_18351,N_10726,N_11961);
or U18352 (N_18352,N_12931,N_10269);
xor U18353 (N_18353,N_12514,N_13186);
and U18354 (N_18354,N_13016,N_12656);
and U18355 (N_18355,N_11130,N_13330);
nor U18356 (N_18356,N_14151,N_11148);
or U18357 (N_18357,N_12828,N_10684);
xnor U18358 (N_18358,N_10984,N_10430);
nand U18359 (N_18359,N_11571,N_14993);
nor U18360 (N_18360,N_13509,N_14968);
nand U18361 (N_18361,N_13326,N_12645);
or U18362 (N_18362,N_11015,N_10096);
or U18363 (N_18363,N_13622,N_12724);
and U18364 (N_18364,N_11183,N_13774);
nand U18365 (N_18365,N_11159,N_10144);
xnor U18366 (N_18366,N_14596,N_13407);
xor U18367 (N_18367,N_10397,N_10607);
xor U18368 (N_18368,N_11080,N_10668);
nor U18369 (N_18369,N_12190,N_11909);
nor U18370 (N_18370,N_14718,N_11908);
nand U18371 (N_18371,N_12778,N_13699);
xor U18372 (N_18372,N_14681,N_10391);
xnor U18373 (N_18373,N_14247,N_14943);
and U18374 (N_18374,N_14853,N_10268);
xor U18375 (N_18375,N_12367,N_10343);
xnor U18376 (N_18376,N_14501,N_10522);
and U18377 (N_18377,N_10147,N_14001);
and U18378 (N_18378,N_11630,N_12081);
and U18379 (N_18379,N_10257,N_12210);
or U18380 (N_18380,N_11830,N_13194);
and U18381 (N_18381,N_13625,N_13286);
and U18382 (N_18382,N_11184,N_14346);
or U18383 (N_18383,N_11700,N_12363);
or U18384 (N_18384,N_12796,N_12608);
nand U18385 (N_18385,N_13429,N_10567);
and U18386 (N_18386,N_14360,N_11499);
xor U18387 (N_18387,N_13473,N_10927);
or U18388 (N_18388,N_14571,N_11633);
or U18389 (N_18389,N_14458,N_10282);
nor U18390 (N_18390,N_14224,N_11373);
and U18391 (N_18391,N_10517,N_12863);
nor U18392 (N_18392,N_10334,N_11555);
xnor U18393 (N_18393,N_13071,N_14259);
nor U18394 (N_18394,N_10031,N_13030);
or U18395 (N_18395,N_10399,N_14191);
or U18396 (N_18396,N_12902,N_10088);
or U18397 (N_18397,N_13237,N_12988);
xor U18398 (N_18398,N_12916,N_10680);
nand U18399 (N_18399,N_10082,N_13938);
xor U18400 (N_18400,N_10584,N_10774);
nor U18401 (N_18401,N_11968,N_10693);
xnor U18402 (N_18402,N_14587,N_12148);
nor U18403 (N_18403,N_14370,N_12278);
or U18404 (N_18404,N_12447,N_14143);
and U18405 (N_18405,N_11492,N_13284);
nand U18406 (N_18406,N_11370,N_13208);
or U18407 (N_18407,N_10607,N_10220);
nand U18408 (N_18408,N_10398,N_14891);
or U18409 (N_18409,N_13646,N_12399);
and U18410 (N_18410,N_10661,N_10564);
nor U18411 (N_18411,N_14136,N_12524);
xnor U18412 (N_18412,N_13356,N_14056);
and U18413 (N_18413,N_11018,N_11644);
xnor U18414 (N_18414,N_10182,N_14252);
nor U18415 (N_18415,N_10697,N_11166);
and U18416 (N_18416,N_10032,N_10648);
xnor U18417 (N_18417,N_12065,N_13863);
xor U18418 (N_18418,N_13468,N_10998);
and U18419 (N_18419,N_13232,N_13662);
nor U18420 (N_18420,N_14469,N_11475);
nor U18421 (N_18421,N_12549,N_11146);
or U18422 (N_18422,N_13178,N_10767);
or U18423 (N_18423,N_10581,N_11167);
nor U18424 (N_18424,N_14656,N_10664);
xnor U18425 (N_18425,N_14272,N_13344);
or U18426 (N_18426,N_12043,N_12207);
or U18427 (N_18427,N_10799,N_14722);
xnor U18428 (N_18428,N_11198,N_14899);
nand U18429 (N_18429,N_13541,N_13548);
and U18430 (N_18430,N_14480,N_14526);
or U18431 (N_18431,N_10760,N_14954);
nand U18432 (N_18432,N_10081,N_10801);
nand U18433 (N_18433,N_13474,N_13157);
nor U18434 (N_18434,N_10661,N_12528);
nand U18435 (N_18435,N_12950,N_12385);
and U18436 (N_18436,N_10947,N_11796);
nand U18437 (N_18437,N_11979,N_10166);
nor U18438 (N_18438,N_13640,N_14739);
nand U18439 (N_18439,N_10164,N_14591);
xor U18440 (N_18440,N_13950,N_14428);
nor U18441 (N_18441,N_10852,N_11095);
nand U18442 (N_18442,N_12181,N_11061);
and U18443 (N_18443,N_12121,N_12348);
and U18444 (N_18444,N_10009,N_12839);
or U18445 (N_18445,N_14941,N_12662);
and U18446 (N_18446,N_14471,N_12411);
nor U18447 (N_18447,N_14556,N_12918);
and U18448 (N_18448,N_14281,N_10661);
xor U18449 (N_18449,N_13137,N_12295);
nor U18450 (N_18450,N_13677,N_14518);
nand U18451 (N_18451,N_11684,N_12696);
or U18452 (N_18452,N_12317,N_14510);
xor U18453 (N_18453,N_13062,N_12184);
nor U18454 (N_18454,N_14870,N_14639);
nor U18455 (N_18455,N_14025,N_13929);
nor U18456 (N_18456,N_11797,N_14424);
xnor U18457 (N_18457,N_12135,N_11162);
or U18458 (N_18458,N_12734,N_10264);
nand U18459 (N_18459,N_12461,N_10467);
xnor U18460 (N_18460,N_14437,N_12475);
nor U18461 (N_18461,N_11960,N_12493);
or U18462 (N_18462,N_12017,N_10545);
and U18463 (N_18463,N_10836,N_11833);
nor U18464 (N_18464,N_10039,N_14085);
nor U18465 (N_18465,N_10208,N_13860);
xor U18466 (N_18466,N_13355,N_12454);
and U18467 (N_18467,N_14607,N_11748);
nand U18468 (N_18468,N_10403,N_14121);
or U18469 (N_18469,N_12704,N_10859);
nand U18470 (N_18470,N_12917,N_10347);
and U18471 (N_18471,N_11659,N_14683);
xnor U18472 (N_18472,N_13298,N_14514);
xnor U18473 (N_18473,N_13963,N_14493);
nand U18474 (N_18474,N_14625,N_10752);
nor U18475 (N_18475,N_12841,N_10404);
xnor U18476 (N_18476,N_13815,N_13509);
nand U18477 (N_18477,N_14252,N_13333);
nand U18478 (N_18478,N_10964,N_10188);
nor U18479 (N_18479,N_12834,N_12102);
nand U18480 (N_18480,N_14369,N_10984);
nand U18481 (N_18481,N_14018,N_14858);
xor U18482 (N_18482,N_10210,N_13530);
and U18483 (N_18483,N_11342,N_12721);
and U18484 (N_18484,N_10512,N_11802);
or U18485 (N_18485,N_12290,N_10791);
nand U18486 (N_18486,N_10096,N_11037);
nand U18487 (N_18487,N_14177,N_14884);
and U18488 (N_18488,N_11733,N_11108);
or U18489 (N_18489,N_12330,N_10293);
nand U18490 (N_18490,N_12129,N_13227);
xor U18491 (N_18491,N_13863,N_14494);
nor U18492 (N_18492,N_10362,N_11564);
or U18493 (N_18493,N_13225,N_12883);
nand U18494 (N_18494,N_11844,N_10948);
or U18495 (N_18495,N_12482,N_14022);
nor U18496 (N_18496,N_14508,N_10412);
or U18497 (N_18497,N_11218,N_11866);
and U18498 (N_18498,N_10173,N_11918);
and U18499 (N_18499,N_10556,N_12851);
xor U18500 (N_18500,N_14660,N_10069);
xor U18501 (N_18501,N_11147,N_12400);
nor U18502 (N_18502,N_12336,N_11847);
and U18503 (N_18503,N_12831,N_12079);
xnor U18504 (N_18504,N_11006,N_11524);
nand U18505 (N_18505,N_10020,N_13656);
and U18506 (N_18506,N_11600,N_11812);
or U18507 (N_18507,N_11713,N_13484);
nor U18508 (N_18508,N_12716,N_13983);
nor U18509 (N_18509,N_13748,N_11761);
xnor U18510 (N_18510,N_11234,N_10813);
nor U18511 (N_18511,N_13361,N_10698);
or U18512 (N_18512,N_13719,N_11212);
xnor U18513 (N_18513,N_12532,N_11793);
and U18514 (N_18514,N_11009,N_11944);
nand U18515 (N_18515,N_12150,N_13632);
nor U18516 (N_18516,N_10306,N_14518);
xor U18517 (N_18517,N_10137,N_12163);
nand U18518 (N_18518,N_12758,N_13362);
nand U18519 (N_18519,N_14097,N_13002);
nor U18520 (N_18520,N_14540,N_12809);
xnor U18521 (N_18521,N_11993,N_13641);
and U18522 (N_18522,N_11718,N_14065);
nand U18523 (N_18523,N_14286,N_10357);
nand U18524 (N_18524,N_10526,N_12375);
and U18525 (N_18525,N_13908,N_12358);
xnor U18526 (N_18526,N_12986,N_11918);
nor U18527 (N_18527,N_10031,N_13644);
or U18528 (N_18528,N_14244,N_11186);
or U18529 (N_18529,N_13297,N_12383);
or U18530 (N_18530,N_10098,N_10052);
xnor U18531 (N_18531,N_11910,N_14107);
nor U18532 (N_18532,N_12226,N_13388);
and U18533 (N_18533,N_11367,N_11421);
nand U18534 (N_18534,N_13315,N_10056);
or U18535 (N_18535,N_10524,N_11024);
xor U18536 (N_18536,N_14397,N_11966);
xnor U18537 (N_18537,N_11356,N_13350);
or U18538 (N_18538,N_10079,N_14920);
or U18539 (N_18539,N_10301,N_14914);
and U18540 (N_18540,N_13794,N_10633);
and U18541 (N_18541,N_12431,N_14650);
and U18542 (N_18542,N_11092,N_13405);
or U18543 (N_18543,N_13405,N_10763);
and U18544 (N_18544,N_13816,N_11604);
nand U18545 (N_18545,N_14636,N_11640);
xnor U18546 (N_18546,N_14427,N_11551);
and U18547 (N_18547,N_13198,N_11187);
xor U18548 (N_18548,N_11760,N_11582);
nand U18549 (N_18549,N_14190,N_13286);
nor U18550 (N_18550,N_13040,N_14221);
or U18551 (N_18551,N_14646,N_12637);
nor U18552 (N_18552,N_14486,N_12465);
nor U18553 (N_18553,N_13481,N_10753);
nand U18554 (N_18554,N_12922,N_10320);
nand U18555 (N_18555,N_13706,N_12454);
xor U18556 (N_18556,N_12193,N_10066);
xor U18557 (N_18557,N_11958,N_12388);
and U18558 (N_18558,N_13741,N_12060);
nand U18559 (N_18559,N_13205,N_12822);
nor U18560 (N_18560,N_11032,N_14968);
xnor U18561 (N_18561,N_10193,N_12193);
or U18562 (N_18562,N_14590,N_13270);
nand U18563 (N_18563,N_12466,N_10581);
or U18564 (N_18564,N_13445,N_13931);
xnor U18565 (N_18565,N_13646,N_10560);
nand U18566 (N_18566,N_10682,N_12880);
and U18567 (N_18567,N_12553,N_12971);
nand U18568 (N_18568,N_11140,N_12211);
nor U18569 (N_18569,N_14137,N_12331);
xnor U18570 (N_18570,N_12167,N_11329);
and U18571 (N_18571,N_10373,N_13735);
or U18572 (N_18572,N_12695,N_13117);
xor U18573 (N_18573,N_11535,N_14188);
and U18574 (N_18574,N_10756,N_12911);
nor U18575 (N_18575,N_14300,N_11863);
or U18576 (N_18576,N_13932,N_13474);
nor U18577 (N_18577,N_13053,N_14763);
and U18578 (N_18578,N_10517,N_13487);
or U18579 (N_18579,N_14643,N_11302);
nand U18580 (N_18580,N_14540,N_13854);
nand U18581 (N_18581,N_12901,N_13651);
and U18582 (N_18582,N_12605,N_11029);
xor U18583 (N_18583,N_13741,N_11110);
nor U18584 (N_18584,N_14042,N_14214);
and U18585 (N_18585,N_13243,N_11248);
or U18586 (N_18586,N_14303,N_11719);
xnor U18587 (N_18587,N_13377,N_12212);
and U18588 (N_18588,N_13757,N_11596);
nor U18589 (N_18589,N_14023,N_11147);
or U18590 (N_18590,N_14749,N_10163);
nand U18591 (N_18591,N_12110,N_12937);
nand U18592 (N_18592,N_13525,N_12462);
nand U18593 (N_18593,N_13514,N_12077);
nand U18594 (N_18594,N_14563,N_13323);
nand U18595 (N_18595,N_10201,N_10989);
or U18596 (N_18596,N_10586,N_11133);
and U18597 (N_18597,N_11419,N_12818);
nand U18598 (N_18598,N_12833,N_13850);
or U18599 (N_18599,N_14090,N_14457);
nor U18600 (N_18600,N_13537,N_10286);
xor U18601 (N_18601,N_14553,N_11517);
xnor U18602 (N_18602,N_11091,N_14530);
nand U18603 (N_18603,N_13586,N_11318);
xnor U18604 (N_18604,N_10671,N_13644);
nor U18605 (N_18605,N_10410,N_14359);
xnor U18606 (N_18606,N_13059,N_10489);
nor U18607 (N_18607,N_10736,N_11716);
xnor U18608 (N_18608,N_13800,N_12706);
xnor U18609 (N_18609,N_14313,N_12032);
nor U18610 (N_18610,N_11492,N_13130);
nor U18611 (N_18611,N_11569,N_11152);
and U18612 (N_18612,N_11580,N_13053);
xor U18613 (N_18613,N_11931,N_12651);
and U18614 (N_18614,N_11288,N_13947);
or U18615 (N_18615,N_13339,N_12015);
nor U18616 (N_18616,N_13852,N_11043);
nand U18617 (N_18617,N_12598,N_10878);
xnor U18618 (N_18618,N_11163,N_10517);
or U18619 (N_18619,N_14375,N_12580);
nand U18620 (N_18620,N_12299,N_11121);
or U18621 (N_18621,N_12314,N_13547);
xor U18622 (N_18622,N_14249,N_10154);
nand U18623 (N_18623,N_11850,N_12807);
and U18624 (N_18624,N_11312,N_13240);
nor U18625 (N_18625,N_10132,N_14549);
nor U18626 (N_18626,N_11324,N_14214);
xnor U18627 (N_18627,N_12763,N_14328);
nor U18628 (N_18628,N_10307,N_11658);
and U18629 (N_18629,N_10596,N_14811);
and U18630 (N_18630,N_12878,N_13304);
nand U18631 (N_18631,N_13612,N_12034);
or U18632 (N_18632,N_14393,N_14655);
or U18633 (N_18633,N_13637,N_11062);
and U18634 (N_18634,N_11142,N_10217);
xnor U18635 (N_18635,N_11185,N_11409);
nor U18636 (N_18636,N_10953,N_11349);
nand U18637 (N_18637,N_13539,N_12096);
or U18638 (N_18638,N_11065,N_11775);
or U18639 (N_18639,N_10341,N_10483);
nor U18640 (N_18640,N_10628,N_12226);
xnor U18641 (N_18641,N_13469,N_11158);
nor U18642 (N_18642,N_12734,N_14763);
or U18643 (N_18643,N_13294,N_13833);
xnor U18644 (N_18644,N_11910,N_14154);
and U18645 (N_18645,N_11712,N_11672);
nor U18646 (N_18646,N_14241,N_14550);
and U18647 (N_18647,N_14720,N_14604);
or U18648 (N_18648,N_12234,N_14615);
or U18649 (N_18649,N_10092,N_12558);
nor U18650 (N_18650,N_13139,N_11823);
nand U18651 (N_18651,N_14630,N_13846);
xnor U18652 (N_18652,N_14065,N_10824);
xnor U18653 (N_18653,N_11189,N_12396);
nor U18654 (N_18654,N_11865,N_11545);
or U18655 (N_18655,N_12239,N_12106);
xnor U18656 (N_18656,N_10227,N_11216);
and U18657 (N_18657,N_11370,N_14210);
nand U18658 (N_18658,N_10880,N_14958);
nand U18659 (N_18659,N_10033,N_14571);
or U18660 (N_18660,N_11585,N_14095);
nand U18661 (N_18661,N_13874,N_14587);
and U18662 (N_18662,N_10194,N_14172);
or U18663 (N_18663,N_13264,N_14413);
or U18664 (N_18664,N_13871,N_10207);
xnor U18665 (N_18665,N_12607,N_11171);
and U18666 (N_18666,N_12618,N_14667);
xor U18667 (N_18667,N_10844,N_13881);
nand U18668 (N_18668,N_10123,N_13974);
and U18669 (N_18669,N_12632,N_13092);
and U18670 (N_18670,N_14149,N_10887);
xor U18671 (N_18671,N_14387,N_11064);
nor U18672 (N_18672,N_11323,N_13269);
and U18673 (N_18673,N_11100,N_11836);
nand U18674 (N_18674,N_13348,N_13680);
nor U18675 (N_18675,N_11930,N_11132);
nor U18676 (N_18676,N_12515,N_11559);
and U18677 (N_18677,N_10697,N_12926);
or U18678 (N_18678,N_12246,N_12915);
xor U18679 (N_18679,N_11978,N_11428);
nor U18680 (N_18680,N_11265,N_12475);
nand U18681 (N_18681,N_10989,N_11348);
or U18682 (N_18682,N_11387,N_12905);
or U18683 (N_18683,N_11312,N_13138);
xnor U18684 (N_18684,N_11596,N_10200);
xor U18685 (N_18685,N_14869,N_14647);
xnor U18686 (N_18686,N_11399,N_10798);
nor U18687 (N_18687,N_14351,N_13833);
nand U18688 (N_18688,N_14036,N_12652);
nand U18689 (N_18689,N_11443,N_13269);
or U18690 (N_18690,N_14284,N_11667);
nand U18691 (N_18691,N_14930,N_11181);
nand U18692 (N_18692,N_13857,N_12226);
nand U18693 (N_18693,N_11877,N_10057);
xnor U18694 (N_18694,N_12243,N_11418);
nor U18695 (N_18695,N_11434,N_11112);
xor U18696 (N_18696,N_12686,N_10995);
nand U18697 (N_18697,N_10230,N_11618);
and U18698 (N_18698,N_10107,N_12857);
nand U18699 (N_18699,N_13015,N_14708);
and U18700 (N_18700,N_13621,N_10183);
nand U18701 (N_18701,N_13875,N_14903);
nor U18702 (N_18702,N_12568,N_10810);
or U18703 (N_18703,N_12833,N_13365);
and U18704 (N_18704,N_11507,N_14076);
or U18705 (N_18705,N_12348,N_11937);
nor U18706 (N_18706,N_13661,N_11266);
and U18707 (N_18707,N_11473,N_14652);
xor U18708 (N_18708,N_10680,N_10933);
and U18709 (N_18709,N_10451,N_14629);
nand U18710 (N_18710,N_13765,N_12030);
or U18711 (N_18711,N_11016,N_10079);
nor U18712 (N_18712,N_11792,N_11615);
nand U18713 (N_18713,N_14084,N_11827);
nand U18714 (N_18714,N_13256,N_11182);
xor U18715 (N_18715,N_14794,N_10641);
xnor U18716 (N_18716,N_11413,N_11551);
nand U18717 (N_18717,N_12824,N_10124);
and U18718 (N_18718,N_14627,N_10336);
and U18719 (N_18719,N_13775,N_11529);
or U18720 (N_18720,N_12455,N_14883);
nor U18721 (N_18721,N_13473,N_13388);
xor U18722 (N_18722,N_12869,N_14450);
or U18723 (N_18723,N_11805,N_14266);
or U18724 (N_18724,N_10447,N_10965);
or U18725 (N_18725,N_10717,N_13718);
or U18726 (N_18726,N_10652,N_12116);
xnor U18727 (N_18727,N_13579,N_11806);
or U18728 (N_18728,N_14229,N_11638);
nor U18729 (N_18729,N_11688,N_14885);
nand U18730 (N_18730,N_12345,N_13793);
nand U18731 (N_18731,N_14830,N_11417);
nor U18732 (N_18732,N_14970,N_11372);
and U18733 (N_18733,N_12224,N_10835);
or U18734 (N_18734,N_13179,N_10153);
and U18735 (N_18735,N_13735,N_11094);
nand U18736 (N_18736,N_13010,N_10379);
xnor U18737 (N_18737,N_13817,N_12660);
xor U18738 (N_18738,N_14345,N_12950);
or U18739 (N_18739,N_11743,N_10014);
nor U18740 (N_18740,N_13478,N_10279);
or U18741 (N_18741,N_12815,N_10418);
nor U18742 (N_18742,N_13355,N_12084);
nand U18743 (N_18743,N_12949,N_14675);
and U18744 (N_18744,N_12424,N_14351);
or U18745 (N_18745,N_12958,N_13784);
or U18746 (N_18746,N_14292,N_11162);
xnor U18747 (N_18747,N_13156,N_10890);
or U18748 (N_18748,N_13185,N_13072);
or U18749 (N_18749,N_14107,N_10041);
or U18750 (N_18750,N_10694,N_11853);
nand U18751 (N_18751,N_13180,N_12241);
xnor U18752 (N_18752,N_11606,N_14581);
nand U18753 (N_18753,N_10007,N_14486);
nor U18754 (N_18754,N_11839,N_12070);
and U18755 (N_18755,N_13369,N_11316);
nor U18756 (N_18756,N_11087,N_10614);
xor U18757 (N_18757,N_10509,N_13654);
or U18758 (N_18758,N_10699,N_10837);
and U18759 (N_18759,N_11287,N_12378);
and U18760 (N_18760,N_14680,N_11470);
xor U18761 (N_18761,N_11542,N_13863);
nor U18762 (N_18762,N_11077,N_14236);
or U18763 (N_18763,N_14010,N_12605);
xnor U18764 (N_18764,N_11974,N_14587);
nand U18765 (N_18765,N_11014,N_10008);
xnor U18766 (N_18766,N_11770,N_10069);
nand U18767 (N_18767,N_12327,N_11846);
xnor U18768 (N_18768,N_14838,N_10596);
xnor U18769 (N_18769,N_10126,N_12100);
xnor U18770 (N_18770,N_11490,N_10162);
xnor U18771 (N_18771,N_12717,N_13207);
xor U18772 (N_18772,N_13871,N_13242);
or U18773 (N_18773,N_13728,N_13138);
nor U18774 (N_18774,N_14455,N_11918);
nand U18775 (N_18775,N_12524,N_13090);
and U18776 (N_18776,N_10216,N_10506);
xor U18777 (N_18777,N_13183,N_14904);
and U18778 (N_18778,N_12419,N_12237);
or U18779 (N_18779,N_13701,N_12202);
nor U18780 (N_18780,N_10767,N_14068);
xnor U18781 (N_18781,N_11646,N_10612);
or U18782 (N_18782,N_12584,N_10074);
nor U18783 (N_18783,N_10904,N_11707);
nor U18784 (N_18784,N_10539,N_12125);
nor U18785 (N_18785,N_10193,N_12899);
or U18786 (N_18786,N_11950,N_13932);
xor U18787 (N_18787,N_12734,N_11644);
or U18788 (N_18788,N_12521,N_12488);
xor U18789 (N_18789,N_14154,N_10909);
nand U18790 (N_18790,N_13250,N_12468);
nand U18791 (N_18791,N_14977,N_12797);
nor U18792 (N_18792,N_11982,N_10951);
or U18793 (N_18793,N_11011,N_13005);
xnor U18794 (N_18794,N_14324,N_13397);
nand U18795 (N_18795,N_10842,N_14655);
or U18796 (N_18796,N_10746,N_10148);
nand U18797 (N_18797,N_10152,N_13647);
or U18798 (N_18798,N_12859,N_13660);
or U18799 (N_18799,N_10219,N_13271);
xor U18800 (N_18800,N_10148,N_10580);
nand U18801 (N_18801,N_14311,N_11706);
nand U18802 (N_18802,N_12601,N_14651);
nand U18803 (N_18803,N_10111,N_13268);
nor U18804 (N_18804,N_12612,N_13695);
nand U18805 (N_18805,N_14257,N_11176);
nor U18806 (N_18806,N_12219,N_14156);
xor U18807 (N_18807,N_14820,N_11493);
and U18808 (N_18808,N_13858,N_10101);
nand U18809 (N_18809,N_14616,N_12683);
xnor U18810 (N_18810,N_12978,N_14064);
nor U18811 (N_18811,N_14357,N_13069);
xor U18812 (N_18812,N_11039,N_10733);
and U18813 (N_18813,N_13242,N_13511);
nand U18814 (N_18814,N_11013,N_10297);
and U18815 (N_18815,N_12534,N_11933);
xnor U18816 (N_18816,N_12905,N_10258);
and U18817 (N_18817,N_13177,N_14306);
nor U18818 (N_18818,N_11013,N_13161);
and U18819 (N_18819,N_14795,N_14382);
xnor U18820 (N_18820,N_10658,N_12274);
xnor U18821 (N_18821,N_12010,N_11276);
xor U18822 (N_18822,N_10507,N_13451);
nor U18823 (N_18823,N_10027,N_13233);
and U18824 (N_18824,N_11840,N_14003);
nand U18825 (N_18825,N_12413,N_10905);
or U18826 (N_18826,N_11183,N_14064);
nor U18827 (N_18827,N_10840,N_12375);
and U18828 (N_18828,N_10278,N_12257);
xnor U18829 (N_18829,N_11001,N_11821);
or U18830 (N_18830,N_12077,N_11634);
nor U18831 (N_18831,N_10866,N_12838);
xor U18832 (N_18832,N_11453,N_11673);
and U18833 (N_18833,N_11343,N_12579);
and U18834 (N_18834,N_11341,N_10537);
xnor U18835 (N_18835,N_14648,N_13501);
or U18836 (N_18836,N_12645,N_14714);
and U18837 (N_18837,N_10073,N_10413);
nor U18838 (N_18838,N_14088,N_14930);
or U18839 (N_18839,N_14126,N_10144);
xnor U18840 (N_18840,N_13892,N_13229);
xnor U18841 (N_18841,N_11701,N_11599);
and U18842 (N_18842,N_12597,N_13514);
nor U18843 (N_18843,N_14688,N_14605);
nand U18844 (N_18844,N_12285,N_14813);
or U18845 (N_18845,N_13816,N_10741);
nand U18846 (N_18846,N_12782,N_11144);
or U18847 (N_18847,N_13405,N_12657);
and U18848 (N_18848,N_14530,N_13641);
xnor U18849 (N_18849,N_12261,N_11691);
xnor U18850 (N_18850,N_12890,N_10622);
nand U18851 (N_18851,N_14260,N_10606);
nand U18852 (N_18852,N_13282,N_13632);
xor U18853 (N_18853,N_12942,N_14173);
xor U18854 (N_18854,N_10424,N_11218);
or U18855 (N_18855,N_11093,N_12740);
and U18856 (N_18856,N_13198,N_11829);
and U18857 (N_18857,N_13173,N_11275);
xnor U18858 (N_18858,N_12301,N_11410);
nor U18859 (N_18859,N_14218,N_13291);
and U18860 (N_18860,N_14892,N_13011);
or U18861 (N_18861,N_12592,N_14292);
and U18862 (N_18862,N_12729,N_11956);
or U18863 (N_18863,N_14070,N_12189);
or U18864 (N_18864,N_10454,N_13749);
or U18865 (N_18865,N_10101,N_11469);
and U18866 (N_18866,N_10066,N_11206);
nand U18867 (N_18867,N_12830,N_14531);
nor U18868 (N_18868,N_11770,N_13724);
nand U18869 (N_18869,N_14870,N_12346);
or U18870 (N_18870,N_11209,N_11352);
xor U18871 (N_18871,N_11510,N_10019);
or U18872 (N_18872,N_11212,N_11969);
or U18873 (N_18873,N_14330,N_10686);
nand U18874 (N_18874,N_12777,N_14004);
and U18875 (N_18875,N_12161,N_11371);
xnor U18876 (N_18876,N_12125,N_11526);
nand U18877 (N_18877,N_14679,N_11529);
nor U18878 (N_18878,N_12500,N_10493);
nand U18879 (N_18879,N_11341,N_12135);
xor U18880 (N_18880,N_10324,N_12591);
or U18881 (N_18881,N_10723,N_13875);
nand U18882 (N_18882,N_13769,N_14838);
xor U18883 (N_18883,N_13838,N_14328);
or U18884 (N_18884,N_11307,N_10223);
xnor U18885 (N_18885,N_14334,N_11754);
nor U18886 (N_18886,N_14920,N_13299);
nand U18887 (N_18887,N_11794,N_12173);
nand U18888 (N_18888,N_10514,N_11272);
and U18889 (N_18889,N_11553,N_11097);
nor U18890 (N_18890,N_13893,N_12251);
nor U18891 (N_18891,N_14035,N_10336);
and U18892 (N_18892,N_10250,N_14521);
nand U18893 (N_18893,N_11999,N_11851);
and U18894 (N_18894,N_13391,N_11724);
nand U18895 (N_18895,N_11616,N_10108);
and U18896 (N_18896,N_12302,N_10703);
and U18897 (N_18897,N_11209,N_14543);
or U18898 (N_18898,N_10093,N_14232);
xnor U18899 (N_18899,N_14955,N_10169);
xnor U18900 (N_18900,N_14897,N_10722);
nor U18901 (N_18901,N_12578,N_13899);
nand U18902 (N_18902,N_11638,N_13979);
nor U18903 (N_18903,N_12474,N_10033);
nand U18904 (N_18904,N_14225,N_12858);
nor U18905 (N_18905,N_12892,N_13066);
or U18906 (N_18906,N_12761,N_11885);
and U18907 (N_18907,N_11595,N_12328);
xnor U18908 (N_18908,N_14789,N_12465);
and U18909 (N_18909,N_11360,N_12436);
nor U18910 (N_18910,N_13535,N_11628);
and U18911 (N_18911,N_14332,N_12314);
nand U18912 (N_18912,N_12037,N_14159);
or U18913 (N_18913,N_12894,N_13380);
and U18914 (N_18914,N_12346,N_11981);
and U18915 (N_18915,N_14955,N_13552);
or U18916 (N_18916,N_11948,N_14181);
xor U18917 (N_18917,N_11901,N_12895);
xor U18918 (N_18918,N_10483,N_14840);
and U18919 (N_18919,N_13787,N_14999);
or U18920 (N_18920,N_12215,N_12966);
and U18921 (N_18921,N_12599,N_14062);
or U18922 (N_18922,N_13544,N_12569);
nand U18923 (N_18923,N_11002,N_13264);
and U18924 (N_18924,N_12442,N_13195);
nand U18925 (N_18925,N_13795,N_10471);
xnor U18926 (N_18926,N_14596,N_10047);
or U18927 (N_18927,N_13906,N_10029);
xnor U18928 (N_18928,N_12538,N_14775);
nor U18929 (N_18929,N_12828,N_12010);
and U18930 (N_18930,N_13673,N_14781);
nand U18931 (N_18931,N_12830,N_11692);
xnor U18932 (N_18932,N_14948,N_13456);
xor U18933 (N_18933,N_13951,N_11727);
nor U18934 (N_18934,N_11768,N_10954);
and U18935 (N_18935,N_12198,N_10044);
xnor U18936 (N_18936,N_10158,N_10630);
xor U18937 (N_18937,N_14022,N_12847);
xnor U18938 (N_18938,N_14240,N_13893);
nand U18939 (N_18939,N_11889,N_12925);
xnor U18940 (N_18940,N_14737,N_11627);
or U18941 (N_18941,N_11701,N_13941);
nor U18942 (N_18942,N_14438,N_14409);
nand U18943 (N_18943,N_13690,N_13764);
nor U18944 (N_18944,N_11288,N_13054);
or U18945 (N_18945,N_14647,N_13929);
nor U18946 (N_18946,N_13165,N_10837);
nor U18947 (N_18947,N_13452,N_13615);
xor U18948 (N_18948,N_14346,N_13716);
or U18949 (N_18949,N_11364,N_10681);
xor U18950 (N_18950,N_14930,N_10293);
and U18951 (N_18951,N_14715,N_14323);
nor U18952 (N_18952,N_12815,N_10456);
and U18953 (N_18953,N_13766,N_10851);
nor U18954 (N_18954,N_11859,N_11645);
nor U18955 (N_18955,N_14272,N_11959);
xnor U18956 (N_18956,N_14360,N_14416);
xnor U18957 (N_18957,N_13965,N_12035);
or U18958 (N_18958,N_10359,N_12189);
and U18959 (N_18959,N_13196,N_12286);
or U18960 (N_18960,N_10102,N_13363);
nor U18961 (N_18961,N_10784,N_14458);
nand U18962 (N_18962,N_14888,N_14816);
nand U18963 (N_18963,N_10993,N_14308);
or U18964 (N_18964,N_11159,N_11360);
and U18965 (N_18965,N_11917,N_14857);
nor U18966 (N_18966,N_10224,N_14936);
or U18967 (N_18967,N_14484,N_12546);
nand U18968 (N_18968,N_12142,N_14346);
xor U18969 (N_18969,N_13006,N_12031);
nand U18970 (N_18970,N_12033,N_12330);
and U18971 (N_18971,N_12730,N_10966);
xnor U18972 (N_18972,N_12076,N_14575);
or U18973 (N_18973,N_14510,N_10747);
nor U18974 (N_18974,N_13273,N_10817);
xnor U18975 (N_18975,N_11781,N_13185);
nor U18976 (N_18976,N_10962,N_11584);
nor U18977 (N_18977,N_13729,N_12123);
or U18978 (N_18978,N_11647,N_10390);
and U18979 (N_18979,N_13147,N_14156);
or U18980 (N_18980,N_14964,N_10842);
nand U18981 (N_18981,N_13581,N_14801);
nor U18982 (N_18982,N_11192,N_10255);
or U18983 (N_18983,N_14891,N_12599);
xor U18984 (N_18984,N_12862,N_12107);
and U18985 (N_18985,N_10896,N_13720);
nand U18986 (N_18986,N_11859,N_14031);
nor U18987 (N_18987,N_12584,N_11842);
nor U18988 (N_18988,N_11965,N_10274);
nand U18989 (N_18989,N_13281,N_12575);
nand U18990 (N_18990,N_14551,N_10925);
or U18991 (N_18991,N_13603,N_13412);
and U18992 (N_18992,N_12123,N_12898);
or U18993 (N_18993,N_10720,N_12662);
xnor U18994 (N_18994,N_11666,N_10660);
and U18995 (N_18995,N_11523,N_14469);
nand U18996 (N_18996,N_13438,N_14076);
and U18997 (N_18997,N_14732,N_12103);
nand U18998 (N_18998,N_13739,N_11029);
nor U18999 (N_18999,N_14199,N_14818);
nor U19000 (N_19000,N_12890,N_14051);
or U19001 (N_19001,N_12749,N_11660);
and U19002 (N_19002,N_10865,N_10585);
nor U19003 (N_19003,N_11450,N_11667);
nor U19004 (N_19004,N_14676,N_13973);
xnor U19005 (N_19005,N_13098,N_14753);
nand U19006 (N_19006,N_12118,N_14324);
or U19007 (N_19007,N_12870,N_12636);
or U19008 (N_19008,N_14072,N_14593);
nand U19009 (N_19009,N_14053,N_13448);
and U19010 (N_19010,N_10732,N_11880);
nor U19011 (N_19011,N_14320,N_12031);
xor U19012 (N_19012,N_14960,N_12932);
xor U19013 (N_19013,N_12032,N_14070);
nand U19014 (N_19014,N_13100,N_14870);
and U19015 (N_19015,N_12356,N_14648);
and U19016 (N_19016,N_13204,N_11107);
and U19017 (N_19017,N_14443,N_10896);
nor U19018 (N_19018,N_13190,N_14055);
and U19019 (N_19019,N_12742,N_11116);
or U19020 (N_19020,N_13106,N_11170);
and U19021 (N_19021,N_12210,N_10728);
or U19022 (N_19022,N_12039,N_13929);
or U19023 (N_19023,N_14050,N_13678);
and U19024 (N_19024,N_14575,N_13298);
xor U19025 (N_19025,N_10399,N_12616);
nor U19026 (N_19026,N_14446,N_14396);
and U19027 (N_19027,N_12134,N_14843);
xnor U19028 (N_19028,N_13313,N_10003);
nand U19029 (N_19029,N_14095,N_10402);
or U19030 (N_19030,N_12663,N_13654);
nand U19031 (N_19031,N_13039,N_11506);
nand U19032 (N_19032,N_12467,N_10262);
and U19033 (N_19033,N_14590,N_14322);
and U19034 (N_19034,N_14475,N_14776);
nand U19035 (N_19035,N_14753,N_10670);
or U19036 (N_19036,N_13907,N_11002);
nor U19037 (N_19037,N_10591,N_13443);
nand U19038 (N_19038,N_13285,N_14277);
and U19039 (N_19039,N_13948,N_11239);
xor U19040 (N_19040,N_10383,N_12534);
xor U19041 (N_19041,N_13164,N_10139);
or U19042 (N_19042,N_13267,N_10735);
or U19043 (N_19043,N_12838,N_14915);
and U19044 (N_19044,N_12268,N_12814);
and U19045 (N_19045,N_10683,N_11845);
xnor U19046 (N_19046,N_11979,N_13952);
nor U19047 (N_19047,N_11154,N_10143);
nand U19048 (N_19048,N_10121,N_14039);
nand U19049 (N_19049,N_11808,N_12982);
xnor U19050 (N_19050,N_14785,N_12601);
or U19051 (N_19051,N_10630,N_13086);
nor U19052 (N_19052,N_12042,N_12153);
nand U19053 (N_19053,N_12256,N_10435);
nand U19054 (N_19054,N_10977,N_14844);
nor U19055 (N_19055,N_13328,N_14932);
nor U19056 (N_19056,N_11717,N_14382);
nor U19057 (N_19057,N_12175,N_10346);
or U19058 (N_19058,N_12243,N_11877);
or U19059 (N_19059,N_11640,N_11084);
nand U19060 (N_19060,N_13802,N_11408);
nand U19061 (N_19061,N_11840,N_13107);
nand U19062 (N_19062,N_14406,N_11822);
xnor U19063 (N_19063,N_11386,N_14008);
or U19064 (N_19064,N_10861,N_12450);
nand U19065 (N_19065,N_12961,N_14967);
nor U19066 (N_19066,N_13710,N_13156);
or U19067 (N_19067,N_11407,N_13008);
xor U19068 (N_19068,N_12841,N_14975);
nand U19069 (N_19069,N_13857,N_13056);
and U19070 (N_19070,N_10754,N_11450);
nor U19071 (N_19071,N_12509,N_14079);
and U19072 (N_19072,N_13566,N_11255);
nand U19073 (N_19073,N_11029,N_12341);
nor U19074 (N_19074,N_12698,N_11421);
nor U19075 (N_19075,N_13855,N_14547);
nor U19076 (N_19076,N_14080,N_14858);
and U19077 (N_19077,N_10003,N_14370);
xor U19078 (N_19078,N_12755,N_13010);
xor U19079 (N_19079,N_11936,N_12616);
or U19080 (N_19080,N_12621,N_14878);
nand U19081 (N_19081,N_14370,N_12910);
nor U19082 (N_19082,N_10998,N_13016);
or U19083 (N_19083,N_14604,N_11764);
or U19084 (N_19084,N_14778,N_10231);
or U19085 (N_19085,N_10804,N_13284);
or U19086 (N_19086,N_14490,N_12765);
and U19087 (N_19087,N_14667,N_13360);
and U19088 (N_19088,N_14665,N_14265);
and U19089 (N_19089,N_12564,N_14590);
and U19090 (N_19090,N_13183,N_10161);
and U19091 (N_19091,N_12404,N_10561);
nand U19092 (N_19092,N_14049,N_12338);
nand U19093 (N_19093,N_14339,N_12771);
and U19094 (N_19094,N_13242,N_10355);
nand U19095 (N_19095,N_11787,N_13943);
and U19096 (N_19096,N_13746,N_13066);
nor U19097 (N_19097,N_14081,N_14774);
and U19098 (N_19098,N_12386,N_11014);
or U19099 (N_19099,N_14135,N_14318);
nor U19100 (N_19100,N_11429,N_13091);
nand U19101 (N_19101,N_11458,N_11861);
nor U19102 (N_19102,N_11557,N_13679);
nor U19103 (N_19103,N_12419,N_11704);
xnor U19104 (N_19104,N_14822,N_13902);
nor U19105 (N_19105,N_10009,N_13845);
xor U19106 (N_19106,N_13773,N_10232);
xnor U19107 (N_19107,N_14873,N_11142);
or U19108 (N_19108,N_14947,N_11475);
xnor U19109 (N_19109,N_14522,N_11705);
xnor U19110 (N_19110,N_10554,N_13188);
nor U19111 (N_19111,N_13938,N_14140);
or U19112 (N_19112,N_11630,N_12239);
nand U19113 (N_19113,N_13089,N_14580);
nor U19114 (N_19114,N_10845,N_13966);
or U19115 (N_19115,N_10631,N_13774);
xor U19116 (N_19116,N_13658,N_14534);
nor U19117 (N_19117,N_10934,N_12519);
nand U19118 (N_19118,N_13172,N_10774);
nand U19119 (N_19119,N_14776,N_14780);
xnor U19120 (N_19120,N_12279,N_12336);
xnor U19121 (N_19121,N_13138,N_13715);
nor U19122 (N_19122,N_10480,N_12936);
nand U19123 (N_19123,N_14603,N_12936);
xor U19124 (N_19124,N_12622,N_14836);
and U19125 (N_19125,N_14226,N_11388);
nand U19126 (N_19126,N_14562,N_12871);
and U19127 (N_19127,N_10399,N_10260);
or U19128 (N_19128,N_13343,N_11554);
nand U19129 (N_19129,N_10825,N_11911);
or U19130 (N_19130,N_10741,N_13708);
and U19131 (N_19131,N_14487,N_14468);
nor U19132 (N_19132,N_11610,N_11253);
nand U19133 (N_19133,N_14900,N_14944);
nand U19134 (N_19134,N_12411,N_12537);
nor U19135 (N_19135,N_12992,N_11514);
nand U19136 (N_19136,N_10700,N_10795);
xnor U19137 (N_19137,N_11728,N_11005);
or U19138 (N_19138,N_13985,N_10575);
or U19139 (N_19139,N_13567,N_12954);
or U19140 (N_19140,N_13033,N_14214);
xor U19141 (N_19141,N_12422,N_10407);
and U19142 (N_19142,N_10398,N_14206);
and U19143 (N_19143,N_14400,N_12049);
xnor U19144 (N_19144,N_11698,N_11225);
nand U19145 (N_19145,N_12701,N_12733);
or U19146 (N_19146,N_13921,N_10223);
nor U19147 (N_19147,N_11654,N_14059);
nand U19148 (N_19148,N_12467,N_12775);
nor U19149 (N_19149,N_13551,N_14088);
or U19150 (N_19150,N_10194,N_12020);
and U19151 (N_19151,N_14903,N_13084);
nor U19152 (N_19152,N_11460,N_14351);
xnor U19153 (N_19153,N_11089,N_13269);
nor U19154 (N_19154,N_13053,N_12078);
or U19155 (N_19155,N_10416,N_10150);
or U19156 (N_19156,N_10138,N_13286);
or U19157 (N_19157,N_14337,N_11120);
nand U19158 (N_19158,N_14409,N_12259);
xnor U19159 (N_19159,N_11006,N_14729);
and U19160 (N_19160,N_13164,N_11179);
and U19161 (N_19161,N_11403,N_11366);
and U19162 (N_19162,N_11522,N_13056);
and U19163 (N_19163,N_12537,N_11083);
nand U19164 (N_19164,N_12340,N_11542);
nand U19165 (N_19165,N_10040,N_10462);
nor U19166 (N_19166,N_13105,N_10808);
nand U19167 (N_19167,N_14987,N_12600);
nand U19168 (N_19168,N_14024,N_10265);
nand U19169 (N_19169,N_14351,N_13600);
nand U19170 (N_19170,N_11616,N_11411);
xnor U19171 (N_19171,N_11210,N_13251);
and U19172 (N_19172,N_10629,N_12259);
and U19173 (N_19173,N_10466,N_11332);
and U19174 (N_19174,N_11313,N_10604);
nand U19175 (N_19175,N_14426,N_14115);
and U19176 (N_19176,N_14811,N_10261);
and U19177 (N_19177,N_14724,N_12704);
nor U19178 (N_19178,N_13536,N_11066);
or U19179 (N_19179,N_13321,N_14398);
nand U19180 (N_19180,N_10891,N_14270);
nand U19181 (N_19181,N_13688,N_11982);
and U19182 (N_19182,N_13603,N_11412);
xnor U19183 (N_19183,N_10599,N_11521);
or U19184 (N_19184,N_14601,N_12311);
nor U19185 (N_19185,N_12507,N_11220);
nand U19186 (N_19186,N_10846,N_14579);
and U19187 (N_19187,N_12674,N_13613);
or U19188 (N_19188,N_11895,N_13332);
and U19189 (N_19189,N_12753,N_11571);
nand U19190 (N_19190,N_14458,N_11077);
or U19191 (N_19191,N_11398,N_10630);
xnor U19192 (N_19192,N_10460,N_12501);
xnor U19193 (N_19193,N_11450,N_14659);
xor U19194 (N_19194,N_13200,N_11745);
or U19195 (N_19195,N_12162,N_14678);
xnor U19196 (N_19196,N_13260,N_14569);
and U19197 (N_19197,N_11963,N_11862);
and U19198 (N_19198,N_11402,N_10937);
and U19199 (N_19199,N_10804,N_10772);
or U19200 (N_19200,N_13850,N_11340);
or U19201 (N_19201,N_12603,N_11035);
nor U19202 (N_19202,N_13356,N_10381);
nand U19203 (N_19203,N_11376,N_12018);
and U19204 (N_19204,N_14512,N_11224);
or U19205 (N_19205,N_12363,N_12799);
or U19206 (N_19206,N_13975,N_12224);
nand U19207 (N_19207,N_12621,N_12344);
or U19208 (N_19208,N_12698,N_12489);
nor U19209 (N_19209,N_11798,N_12016);
or U19210 (N_19210,N_11747,N_12224);
xnor U19211 (N_19211,N_14157,N_11130);
and U19212 (N_19212,N_14143,N_11216);
xor U19213 (N_19213,N_13276,N_14785);
and U19214 (N_19214,N_10798,N_10149);
nand U19215 (N_19215,N_13749,N_14248);
or U19216 (N_19216,N_14581,N_10669);
and U19217 (N_19217,N_12527,N_13356);
xnor U19218 (N_19218,N_14039,N_10047);
nand U19219 (N_19219,N_12723,N_14303);
and U19220 (N_19220,N_12487,N_10830);
nand U19221 (N_19221,N_13688,N_11324);
nor U19222 (N_19222,N_13459,N_14141);
xnor U19223 (N_19223,N_11559,N_12631);
nor U19224 (N_19224,N_14795,N_11600);
xnor U19225 (N_19225,N_14471,N_14965);
or U19226 (N_19226,N_12887,N_13362);
nor U19227 (N_19227,N_12950,N_10686);
and U19228 (N_19228,N_11451,N_12508);
nand U19229 (N_19229,N_12830,N_13112);
nand U19230 (N_19230,N_11763,N_11905);
xor U19231 (N_19231,N_13647,N_12355);
or U19232 (N_19232,N_11377,N_14217);
nor U19233 (N_19233,N_14620,N_14468);
nand U19234 (N_19234,N_12990,N_13712);
or U19235 (N_19235,N_14847,N_13251);
and U19236 (N_19236,N_10192,N_14178);
xnor U19237 (N_19237,N_10963,N_11752);
nand U19238 (N_19238,N_12633,N_14414);
nand U19239 (N_19239,N_13664,N_11633);
xor U19240 (N_19240,N_11153,N_11207);
xnor U19241 (N_19241,N_11079,N_11433);
or U19242 (N_19242,N_13284,N_14474);
or U19243 (N_19243,N_14229,N_14712);
nor U19244 (N_19244,N_11900,N_13368);
nand U19245 (N_19245,N_11074,N_12150);
nand U19246 (N_19246,N_12963,N_14045);
nand U19247 (N_19247,N_14373,N_11902);
nand U19248 (N_19248,N_13394,N_14831);
or U19249 (N_19249,N_10562,N_12648);
xor U19250 (N_19250,N_13002,N_10628);
nor U19251 (N_19251,N_10277,N_10171);
nor U19252 (N_19252,N_14793,N_11357);
and U19253 (N_19253,N_12050,N_14028);
nand U19254 (N_19254,N_14676,N_14054);
or U19255 (N_19255,N_12295,N_14517);
or U19256 (N_19256,N_13592,N_12469);
and U19257 (N_19257,N_11208,N_10628);
nor U19258 (N_19258,N_13631,N_14057);
nor U19259 (N_19259,N_14358,N_13564);
nor U19260 (N_19260,N_13286,N_13490);
nand U19261 (N_19261,N_10941,N_13619);
and U19262 (N_19262,N_13295,N_12024);
and U19263 (N_19263,N_11058,N_12062);
nand U19264 (N_19264,N_13844,N_13424);
or U19265 (N_19265,N_14381,N_11696);
or U19266 (N_19266,N_12533,N_12980);
or U19267 (N_19267,N_12455,N_10047);
nand U19268 (N_19268,N_13503,N_11341);
nand U19269 (N_19269,N_12871,N_14511);
or U19270 (N_19270,N_14926,N_13704);
and U19271 (N_19271,N_13021,N_12610);
or U19272 (N_19272,N_11708,N_10235);
nand U19273 (N_19273,N_11284,N_11572);
or U19274 (N_19274,N_12087,N_11682);
xor U19275 (N_19275,N_12041,N_13360);
xor U19276 (N_19276,N_12007,N_12725);
or U19277 (N_19277,N_13579,N_14998);
nand U19278 (N_19278,N_14811,N_12092);
xor U19279 (N_19279,N_11514,N_13106);
and U19280 (N_19280,N_10486,N_10100);
nand U19281 (N_19281,N_10516,N_10861);
and U19282 (N_19282,N_14510,N_11996);
nor U19283 (N_19283,N_11733,N_12117);
xnor U19284 (N_19284,N_11091,N_13205);
and U19285 (N_19285,N_13824,N_13146);
or U19286 (N_19286,N_10170,N_14977);
nor U19287 (N_19287,N_11954,N_10880);
xnor U19288 (N_19288,N_12248,N_13695);
xor U19289 (N_19289,N_14040,N_12848);
nor U19290 (N_19290,N_13801,N_10123);
or U19291 (N_19291,N_11772,N_10644);
xor U19292 (N_19292,N_11849,N_14938);
nand U19293 (N_19293,N_13199,N_10950);
nand U19294 (N_19294,N_13878,N_10102);
nand U19295 (N_19295,N_10445,N_12479);
or U19296 (N_19296,N_10414,N_10785);
nand U19297 (N_19297,N_10965,N_14227);
or U19298 (N_19298,N_10576,N_13329);
or U19299 (N_19299,N_14735,N_10334);
nor U19300 (N_19300,N_12469,N_11712);
xor U19301 (N_19301,N_14634,N_12327);
nor U19302 (N_19302,N_13459,N_10207);
and U19303 (N_19303,N_13554,N_13096);
nor U19304 (N_19304,N_12149,N_14493);
or U19305 (N_19305,N_13591,N_11160);
and U19306 (N_19306,N_12322,N_14932);
nand U19307 (N_19307,N_11943,N_14496);
and U19308 (N_19308,N_14770,N_11015);
nand U19309 (N_19309,N_14763,N_13276);
xnor U19310 (N_19310,N_12143,N_13897);
xnor U19311 (N_19311,N_14034,N_13687);
xnor U19312 (N_19312,N_12849,N_14291);
xnor U19313 (N_19313,N_12357,N_14833);
nor U19314 (N_19314,N_12756,N_13519);
or U19315 (N_19315,N_11567,N_11373);
nand U19316 (N_19316,N_11552,N_10013);
or U19317 (N_19317,N_10020,N_13451);
nor U19318 (N_19318,N_10824,N_12057);
xnor U19319 (N_19319,N_13384,N_12947);
or U19320 (N_19320,N_14532,N_13323);
nand U19321 (N_19321,N_12283,N_10142);
xnor U19322 (N_19322,N_10278,N_13807);
and U19323 (N_19323,N_13127,N_14593);
nand U19324 (N_19324,N_11444,N_10163);
nor U19325 (N_19325,N_12477,N_11197);
xor U19326 (N_19326,N_10860,N_14837);
and U19327 (N_19327,N_14064,N_13300);
xor U19328 (N_19328,N_11973,N_13807);
or U19329 (N_19329,N_10637,N_14198);
nand U19330 (N_19330,N_14062,N_12330);
xor U19331 (N_19331,N_11940,N_10327);
or U19332 (N_19332,N_10581,N_10945);
nand U19333 (N_19333,N_12060,N_12788);
nand U19334 (N_19334,N_13830,N_13452);
nor U19335 (N_19335,N_10890,N_10322);
nand U19336 (N_19336,N_14676,N_12438);
xor U19337 (N_19337,N_13382,N_10431);
nand U19338 (N_19338,N_10295,N_10594);
nor U19339 (N_19339,N_10481,N_10708);
nand U19340 (N_19340,N_10387,N_12342);
nor U19341 (N_19341,N_13809,N_14251);
and U19342 (N_19342,N_12638,N_11700);
or U19343 (N_19343,N_14697,N_14863);
nor U19344 (N_19344,N_11444,N_13065);
and U19345 (N_19345,N_11262,N_12203);
and U19346 (N_19346,N_13925,N_11017);
or U19347 (N_19347,N_14115,N_11761);
xnor U19348 (N_19348,N_11967,N_14372);
xor U19349 (N_19349,N_10114,N_11984);
nor U19350 (N_19350,N_10430,N_13994);
xor U19351 (N_19351,N_11976,N_11172);
nor U19352 (N_19352,N_10931,N_10507);
and U19353 (N_19353,N_14207,N_12072);
nor U19354 (N_19354,N_13882,N_14841);
nor U19355 (N_19355,N_10688,N_10999);
and U19356 (N_19356,N_11839,N_11537);
or U19357 (N_19357,N_14972,N_13847);
or U19358 (N_19358,N_11565,N_13611);
or U19359 (N_19359,N_13779,N_10276);
nor U19360 (N_19360,N_14185,N_14218);
and U19361 (N_19361,N_12266,N_14783);
and U19362 (N_19362,N_13322,N_10342);
and U19363 (N_19363,N_11686,N_10338);
and U19364 (N_19364,N_12458,N_11249);
or U19365 (N_19365,N_10562,N_10485);
nor U19366 (N_19366,N_14445,N_13996);
or U19367 (N_19367,N_14293,N_11705);
nor U19368 (N_19368,N_13284,N_13168);
nor U19369 (N_19369,N_14020,N_11252);
nand U19370 (N_19370,N_14902,N_13697);
nor U19371 (N_19371,N_12380,N_10995);
and U19372 (N_19372,N_13540,N_13284);
nand U19373 (N_19373,N_14530,N_10625);
and U19374 (N_19374,N_13155,N_10864);
or U19375 (N_19375,N_10610,N_10780);
xor U19376 (N_19376,N_11876,N_11230);
or U19377 (N_19377,N_14642,N_13700);
or U19378 (N_19378,N_10778,N_14088);
or U19379 (N_19379,N_14595,N_10915);
nand U19380 (N_19380,N_14738,N_10329);
or U19381 (N_19381,N_12029,N_11093);
and U19382 (N_19382,N_10053,N_12588);
xnor U19383 (N_19383,N_10131,N_12286);
or U19384 (N_19384,N_13525,N_11679);
nand U19385 (N_19385,N_12235,N_11519);
or U19386 (N_19386,N_14038,N_12907);
nor U19387 (N_19387,N_14993,N_12372);
nor U19388 (N_19388,N_14617,N_12114);
nor U19389 (N_19389,N_12838,N_10346);
nor U19390 (N_19390,N_13332,N_12203);
xor U19391 (N_19391,N_11209,N_14074);
and U19392 (N_19392,N_12722,N_13723);
nor U19393 (N_19393,N_11510,N_11170);
nand U19394 (N_19394,N_13360,N_13350);
or U19395 (N_19395,N_14061,N_14790);
and U19396 (N_19396,N_14171,N_13058);
xor U19397 (N_19397,N_11232,N_10319);
or U19398 (N_19398,N_11245,N_10727);
xnor U19399 (N_19399,N_14205,N_13217);
nand U19400 (N_19400,N_13419,N_12804);
nor U19401 (N_19401,N_10542,N_13573);
nand U19402 (N_19402,N_12006,N_11130);
nand U19403 (N_19403,N_14333,N_12788);
nand U19404 (N_19404,N_13434,N_13491);
nor U19405 (N_19405,N_14850,N_12740);
nor U19406 (N_19406,N_13429,N_12122);
nand U19407 (N_19407,N_13989,N_13519);
and U19408 (N_19408,N_12203,N_10524);
nand U19409 (N_19409,N_13963,N_13452);
or U19410 (N_19410,N_12875,N_13973);
xor U19411 (N_19411,N_11435,N_13965);
nand U19412 (N_19412,N_12050,N_13578);
nor U19413 (N_19413,N_14431,N_10438);
nor U19414 (N_19414,N_14982,N_10302);
or U19415 (N_19415,N_13735,N_14302);
and U19416 (N_19416,N_12031,N_13485);
or U19417 (N_19417,N_13721,N_11200);
or U19418 (N_19418,N_12421,N_12614);
and U19419 (N_19419,N_13762,N_13377);
xnor U19420 (N_19420,N_12038,N_10446);
nor U19421 (N_19421,N_10516,N_12085);
xnor U19422 (N_19422,N_12647,N_14052);
nor U19423 (N_19423,N_11977,N_10070);
or U19424 (N_19424,N_14745,N_10101);
nor U19425 (N_19425,N_10679,N_14516);
xor U19426 (N_19426,N_10368,N_11057);
or U19427 (N_19427,N_10434,N_10006);
or U19428 (N_19428,N_12078,N_13159);
and U19429 (N_19429,N_13747,N_13303);
nor U19430 (N_19430,N_10543,N_10658);
nand U19431 (N_19431,N_14921,N_13588);
nor U19432 (N_19432,N_11124,N_10785);
xor U19433 (N_19433,N_12811,N_13936);
nor U19434 (N_19434,N_12771,N_10112);
nand U19435 (N_19435,N_12569,N_11278);
xnor U19436 (N_19436,N_12025,N_14498);
xor U19437 (N_19437,N_11332,N_11192);
nand U19438 (N_19438,N_12489,N_13957);
and U19439 (N_19439,N_11375,N_13599);
xnor U19440 (N_19440,N_11802,N_14763);
or U19441 (N_19441,N_12701,N_13361);
nand U19442 (N_19442,N_13024,N_12483);
and U19443 (N_19443,N_14220,N_14039);
nand U19444 (N_19444,N_13286,N_10782);
nand U19445 (N_19445,N_12196,N_14119);
and U19446 (N_19446,N_14150,N_11164);
nand U19447 (N_19447,N_11514,N_10570);
or U19448 (N_19448,N_10958,N_14366);
xnor U19449 (N_19449,N_10065,N_11150);
nor U19450 (N_19450,N_11507,N_11670);
nor U19451 (N_19451,N_13960,N_11294);
nor U19452 (N_19452,N_14028,N_11386);
nor U19453 (N_19453,N_13472,N_12657);
nand U19454 (N_19454,N_13904,N_10242);
nand U19455 (N_19455,N_14349,N_13338);
and U19456 (N_19456,N_14942,N_11390);
xor U19457 (N_19457,N_12171,N_11385);
and U19458 (N_19458,N_14382,N_13787);
nor U19459 (N_19459,N_13468,N_14634);
nor U19460 (N_19460,N_12117,N_12662);
xnor U19461 (N_19461,N_14845,N_10331);
xor U19462 (N_19462,N_14477,N_14565);
or U19463 (N_19463,N_13780,N_12418);
xnor U19464 (N_19464,N_12429,N_11471);
nor U19465 (N_19465,N_10556,N_14461);
xor U19466 (N_19466,N_10893,N_11641);
xor U19467 (N_19467,N_14906,N_13742);
xor U19468 (N_19468,N_12184,N_11512);
nand U19469 (N_19469,N_13514,N_14643);
xor U19470 (N_19470,N_11482,N_12764);
nand U19471 (N_19471,N_11579,N_12146);
xor U19472 (N_19472,N_11222,N_14247);
and U19473 (N_19473,N_13403,N_13115);
nand U19474 (N_19474,N_12764,N_12220);
and U19475 (N_19475,N_13863,N_10143);
nand U19476 (N_19476,N_14877,N_14198);
nand U19477 (N_19477,N_14794,N_12594);
and U19478 (N_19478,N_12483,N_10575);
and U19479 (N_19479,N_13798,N_10755);
xnor U19480 (N_19480,N_13623,N_13492);
nor U19481 (N_19481,N_14931,N_13153);
xnor U19482 (N_19482,N_14420,N_11598);
nand U19483 (N_19483,N_12999,N_11601);
xnor U19484 (N_19484,N_10020,N_10003);
nor U19485 (N_19485,N_14406,N_10597);
nand U19486 (N_19486,N_12558,N_14200);
xor U19487 (N_19487,N_12947,N_14810);
or U19488 (N_19488,N_12744,N_13378);
and U19489 (N_19489,N_12053,N_13892);
xnor U19490 (N_19490,N_14265,N_10265);
nor U19491 (N_19491,N_14348,N_13908);
xor U19492 (N_19492,N_11920,N_14304);
nor U19493 (N_19493,N_12790,N_10356);
and U19494 (N_19494,N_12026,N_14337);
nand U19495 (N_19495,N_11883,N_12917);
xor U19496 (N_19496,N_12601,N_14004);
and U19497 (N_19497,N_12246,N_13847);
and U19498 (N_19498,N_11068,N_13697);
and U19499 (N_19499,N_11716,N_13990);
xor U19500 (N_19500,N_14675,N_12341);
xnor U19501 (N_19501,N_14766,N_10799);
and U19502 (N_19502,N_13569,N_10118);
xnor U19503 (N_19503,N_12533,N_10813);
xnor U19504 (N_19504,N_13224,N_13849);
nor U19505 (N_19505,N_11491,N_11684);
nand U19506 (N_19506,N_12802,N_10677);
nand U19507 (N_19507,N_14093,N_11467);
xnor U19508 (N_19508,N_14591,N_12974);
nor U19509 (N_19509,N_10565,N_10166);
xnor U19510 (N_19510,N_13989,N_12066);
and U19511 (N_19511,N_12719,N_11729);
nor U19512 (N_19512,N_14992,N_14864);
nand U19513 (N_19513,N_11716,N_13104);
nor U19514 (N_19514,N_12844,N_12994);
nor U19515 (N_19515,N_10472,N_11981);
nand U19516 (N_19516,N_10430,N_13755);
xor U19517 (N_19517,N_14844,N_12869);
or U19518 (N_19518,N_12183,N_12639);
or U19519 (N_19519,N_10487,N_13312);
and U19520 (N_19520,N_13019,N_14261);
and U19521 (N_19521,N_12439,N_13957);
and U19522 (N_19522,N_10884,N_14912);
and U19523 (N_19523,N_11167,N_10495);
or U19524 (N_19524,N_10655,N_11216);
xor U19525 (N_19525,N_13511,N_11421);
and U19526 (N_19526,N_14566,N_11867);
nor U19527 (N_19527,N_10170,N_10229);
xor U19528 (N_19528,N_11194,N_14320);
nand U19529 (N_19529,N_12866,N_11753);
nor U19530 (N_19530,N_10355,N_14634);
nand U19531 (N_19531,N_11491,N_11313);
or U19532 (N_19532,N_10140,N_10156);
and U19533 (N_19533,N_11346,N_12071);
xnor U19534 (N_19534,N_11743,N_12885);
nand U19535 (N_19535,N_13967,N_14395);
xor U19536 (N_19536,N_13009,N_11274);
nand U19537 (N_19537,N_12283,N_10212);
nand U19538 (N_19538,N_13398,N_11260);
nand U19539 (N_19539,N_14180,N_14144);
nand U19540 (N_19540,N_13253,N_14420);
xor U19541 (N_19541,N_11693,N_11071);
nor U19542 (N_19542,N_13440,N_13760);
nand U19543 (N_19543,N_10230,N_11333);
xor U19544 (N_19544,N_13367,N_11140);
and U19545 (N_19545,N_14446,N_13330);
and U19546 (N_19546,N_12481,N_10290);
nand U19547 (N_19547,N_14157,N_13244);
or U19548 (N_19548,N_12371,N_10522);
or U19549 (N_19549,N_11955,N_14334);
and U19550 (N_19550,N_12025,N_14647);
or U19551 (N_19551,N_11826,N_12485);
and U19552 (N_19552,N_12481,N_13057);
or U19553 (N_19553,N_14408,N_14943);
and U19554 (N_19554,N_14813,N_11507);
nand U19555 (N_19555,N_14021,N_12336);
and U19556 (N_19556,N_10049,N_14658);
and U19557 (N_19557,N_14312,N_13228);
nor U19558 (N_19558,N_13218,N_10542);
nand U19559 (N_19559,N_12547,N_14250);
and U19560 (N_19560,N_14848,N_14317);
and U19561 (N_19561,N_13382,N_10741);
nor U19562 (N_19562,N_12773,N_14426);
nor U19563 (N_19563,N_11776,N_10822);
or U19564 (N_19564,N_10151,N_12116);
nor U19565 (N_19565,N_12617,N_14253);
and U19566 (N_19566,N_10189,N_11148);
or U19567 (N_19567,N_12145,N_11481);
nand U19568 (N_19568,N_14492,N_12372);
nor U19569 (N_19569,N_11807,N_11511);
and U19570 (N_19570,N_11278,N_12638);
xnor U19571 (N_19571,N_12850,N_12864);
or U19572 (N_19572,N_11219,N_10000);
or U19573 (N_19573,N_14204,N_10809);
nand U19574 (N_19574,N_14754,N_13901);
nor U19575 (N_19575,N_11368,N_12586);
xnor U19576 (N_19576,N_11456,N_14895);
nand U19577 (N_19577,N_12133,N_13146);
xor U19578 (N_19578,N_13167,N_10487);
xor U19579 (N_19579,N_12421,N_11961);
and U19580 (N_19580,N_14333,N_10525);
and U19581 (N_19581,N_11734,N_11274);
nand U19582 (N_19582,N_12392,N_13081);
nand U19583 (N_19583,N_13202,N_12505);
xnor U19584 (N_19584,N_10281,N_11741);
nor U19585 (N_19585,N_13312,N_10012);
xor U19586 (N_19586,N_12051,N_11425);
nand U19587 (N_19587,N_12949,N_13458);
nor U19588 (N_19588,N_11515,N_11513);
nand U19589 (N_19589,N_11590,N_10990);
nand U19590 (N_19590,N_10884,N_14622);
nor U19591 (N_19591,N_10745,N_12766);
or U19592 (N_19592,N_10283,N_14494);
or U19593 (N_19593,N_13746,N_11661);
and U19594 (N_19594,N_10054,N_11272);
nand U19595 (N_19595,N_10898,N_10271);
nand U19596 (N_19596,N_14406,N_10529);
nor U19597 (N_19597,N_12750,N_11003);
and U19598 (N_19598,N_12899,N_13494);
xor U19599 (N_19599,N_14142,N_13739);
or U19600 (N_19600,N_13707,N_10913);
and U19601 (N_19601,N_12096,N_14952);
and U19602 (N_19602,N_14634,N_12758);
nor U19603 (N_19603,N_13952,N_14715);
nand U19604 (N_19604,N_14731,N_12848);
xnor U19605 (N_19605,N_11444,N_14427);
and U19606 (N_19606,N_10906,N_10282);
or U19607 (N_19607,N_13449,N_13253);
nor U19608 (N_19608,N_10462,N_12756);
and U19609 (N_19609,N_14596,N_12715);
and U19610 (N_19610,N_10095,N_10883);
xor U19611 (N_19611,N_10646,N_11839);
nor U19612 (N_19612,N_10736,N_13333);
or U19613 (N_19613,N_12858,N_14319);
and U19614 (N_19614,N_14708,N_11137);
nand U19615 (N_19615,N_11820,N_14507);
or U19616 (N_19616,N_10349,N_12049);
nor U19617 (N_19617,N_13205,N_10508);
nor U19618 (N_19618,N_13608,N_13700);
nand U19619 (N_19619,N_12915,N_13702);
xnor U19620 (N_19620,N_10248,N_14651);
nor U19621 (N_19621,N_11567,N_11907);
nand U19622 (N_19622,N_11942,N_10569);
nand U19623 (N_19623,N_10743,N_11455);
or U19624 (N_19624,N_12662,N_11667);
nand U19625 (N_19625,N_10367,N_12174);
or U19626 (N_19626,N_11099,N_10755);
nand U19627 (N_19627,N_14585,N_14505);
nand U19628 (N_19628,N_11737,N_12309);
xnor U19629 (N_19629,N_10356,N_11041);
nand U19630 (N_19630,N_10841,N_11011);
or U19631 (N_19631,N_13648,N_13100);
xor U19632 (N_19632,N_13937,N_11163);
or U19633 (N_19633,N_13540,N_10864);
or U19634 (N_19634,N_14986,N_12543);
or U19635 (N_19635,N_13060,N_12188);
or U19636 (N_19636,N_13487,N_14477);
or U19637 (N_19637,N_12007,N_14746);
or U19638 (N_19638,N_11287,N_12174);
xor U19639 (N_19639,N_12345,N_12887);
nor U19640 (N_19640,N_10584,N_13243);
xnor U19641 (N_19641,N_14182,N_12180);
or U19642 (N_19642,N_11957,N_12512);
nand U19643 (N_19643,N_14916,N_12939);
xor U19644 (N_19644,N_11035,N_14727);
nor U19645 (N_19645,N_11484,N_10013);
xnor U19646 (N_19646,N_12310,N_12169);
nor U19647 (N_19647,N_10804,N_10439);
nand U19648 (N_19648,N_12656,N_10044);
xnor U19649 (N_19649,N_12149,N_12964);
nand U19650 (N_19650,N_12273,N_12518);
or U19651 (N_19651,N_12589,N_10709);
or U19652 (N_19652,N_10025,N_11738);
xnor U19653 (N_19653,N_11235,N_11040);
nand U19654 (N_19654,N_12551,N_10967);
or U19655 (N_19655,N_12392,N_14099);
nand U19656 (N_19656,N_14093,N_12209);
or U19657 (N_19657,N_12118,N_13904);
nand U19658 (N_19658,N_12819,N_11343);
xnor U19659 (N_19659,N_14802,N_12610);
or U19660 (N_19660,N_13865,N_14445);
nor U19661 (N_19661,N_10554,N_14446);
or U19662 (N_19662,N_13388,N_12989);
and U19663 (N_19663,N_11284,N_13728);
nor U19664 (N_19664,N_13324,N_10372);
nor U19665 (N_19665,N_11965,N_12202);
and U19666 (N_19666,N_13079,N_11337);
and U19667 (N_19667,N_10743,N_13116);
or U19668 (N_19668,N_12269,N_11660);
or U19669 (N_19669,N_10647,N_11541);
nand U19670 (N_19670,N_12610,N_13227);
nand U19671 (N_19671,N_11035,N_14177);
nor U19672 (N_19672,N_13198,N_10053);
and U19673 (N_19673,N_11722,N_12076);
and U19674 (N_19674,N_12243,N_11895);
nand U19675 (N_19675,N_10757,N_12953);
and U19676 (N_19676,N_11846,N_13628);
xor U19677 (N_19677,N_12232,N_13063);
nor U19678 (N_19678,N_11362,N_12326);
xor U19679 (N_19679,N_11057,N_11249);
and U19680 (N_19680,N_13754,N_14992);
or U19681 (N_19681,N_11433,N_12053);
or U19682 (N_19682,N_10230,N_11296);
xor U19683 (N_19683,N_14399,N_14998);
nand U19684 (N_19684,N_10184,N_10587);
or U19685 (N_19685,N_13359,N_11623);
and U19686 (N_19686,N_14430,N_12106);
nand U19687 (N_19687,N_13600,N_10908);
nor U19688 (N_19688,N_14619,N_12063);
and U19689 (N_19689,N_14940,N_10760);
nor U19690 (N_19690,N_12684,N_14760);
xnor U19691 (N_19691,N_14447,N_11785);
or U19692 (N_19692,N_11300,N_13691);
and U19693 (N_19693,N_10982,N_12764);
and U19694 (N_19694,N_10969,N_11995);
xnor U19695 (N_19695,N_11302,N_13022);
nor U19696 (N_19696,N_13936,N_12075);
nand U19697 (N_19697,N_13835,N_13592);
or U19698 (N_19698,N_14153,N_14918);
nand U19699 (N_19699,N_12018,N_12173);
and U19700 (N_19700,N_14802,N_10655);
nor U19701 (N_19701,N_10733,N_10901);
and U19702 (N_19702,N_10559,N_12748);
or U19703 (N_19703,N_10238,N_10122);
and U19704 (N_19704,N_14977,N_11187);
and U19705 (N_19705,N_10959,N_11387);
xnor U19706 (N_19706,N_14833,N_13902);
nand U19707 (N_19707,N_12147,N_12967);
and U19708 (N_19708,N_11727,N_10166);
or U19709 (N_19709,N_14952,N_14720);
nor U19710 (N_19710,N_13508,N_11853);
xor U19711 (N_19711,N_10196,N_14810);
nand U19712 (N_19712,N_10997,N_14075);
and U19713 (N_19713,N_11463,N_13624);
nor U19714 (N_19714,N_14641,N_11767);
xnor U19715 (N_19715,N_14008,N_14874);
or U19716 (N_19716,N_10093,N_12751);
or U19717 (N_19717,N_10330,N_10620);
and U19718 (N_19718,N_13050,N_13831);
and U19719 (N_19719,N_11014,N_11563);
nor U19720 (N_19720,N_10055,N_13120);
xor U19721 (N_19721,N_12760,N_12409);
nand U19722 (N_19722,N_12994,N_14885);
and U19723 (N_19723,N_10979,N_13588);
xnor U19724 (N_19724,N_11884,N_12137);
and U19725 (N_19725,N_14382,N_11651);
nand U19726 (N_19726,N_12304,N_13135);
and U19727 (N_19727,N_12418,N_11812);
xor U19728 (N_19728,N_11839,N_11303);
and U19729 (N_19729,N_10437,N_12938);
xnor U19730 (N_19730,N_14523,N_14818);
xnor U19731 (N_19731,N_13469,N_10338);
nand U19732 (N_19732,N_14838,N_12329);
nor U19733 (N_19733,N_14886,N_12584);
nand U19734 (N_19734,N_12759,N_14139);
xor U19735 (N_19735,N_11820,N_14924);
nand U19736 (N_19736,N_10748,N_13474);
or U19737 (N_19737,N_14490,N_14010);
xor U19738 (N_19738,N_13343,N_12273);
and U19739 (N_19739,N_12515,N_12592);
nor U19740 (N_19740,N_14074,N_14304);
xnor U19741 (N_19741,N_13403,N_14440);
and U19742 (N_19742,N_14470,N_13200);
nor U19743 (N_19743,N_14716,N_13858);
and U19744 (N_19744,N_10875,N_13096);
nor U19745 (N_19745,N_14981,N_13661);
nor U19746 (N_19746,N_11508,N_14233);
and U19747 (N_19747,N_13970,N_10070);
nand U19748 (N_19748,N_10024,N_14526);
nor U19749 (N_19749,N_13112,N_13405);
nand U19750 (N_19750,N_14013,N_12959);
nor U19751 (N_19751,N_14393,N_12913);
or U19752 (N_19752,N_14231,N_14771);
xor U19753 (N_19753,N_11309,N_11823);
or U19754 (N_19754,N_13686,N_11454);
and U19755 (N_19755,N_10425,N_12561);
and U19756 (N_19756,N_12734,N_10630);
or U19757 (N_19757,N_11251,N_14122);
or U19758 (N_19758,N_12203,N_14762);
or U19759 (N_19759,N_14822,N_14359);
nand U19760 (N_19760,N_11783,N_10870);
or U19761 (N_19761,N_12995,N_12887);
nand U19762 (N_19762,N_11229,N_10343);
xnor U19763 (N_19763,N_11914,N_14019);
nand U19764 (N_19764,N_10151,N_13680);
and U19765 (N_19765,N_13100,N_11474);
or U19766 (N_19766,N_14630,N_10917);
nand U19767 (N_19767,N_13460,N_14341);
xor U19768 (N_19768,N_14809,N_14193);
xnor U19769 (N_19769,N_10137,N_10929);
xor U19770 (N_19770,N_13892,N_13885);
and U19771 (N_19771,N_14148,N_12876);
nor U19772 (N_19772,N_11678,N_10308);
xnor U19773 (N_19773,N_10150,N_14871);
nor U19774 (N_19774,N_14392,N_14908);
xnor U19775 (N_19775,N_11301,N_12353);
xor U19776 (N_19776,N_10753,N_13367);
or U19777 (N_19777,N_12801,N_14098);
nor U19778 (N_19778,N_10063,N_11792);
or U19779 (N_19779,N_10541,N_10213);
xnor U19780 (N_19780,N_11871,N_10181);
or U19781 (N_19781,N_11190,N_13529);
or U19782 (N_19782,N_12611,N_10789);
nand U19783 (N_19783,N_14910,N_11403);
nand U19784 (N_19784,N_14380,N_14391);
nor U19785 (N_19785,N_12022,N_14492);
nor U19786 (N_19786,N_12909,N_10854);
xnor U19787 (N_19787,N_13917,N_11850);
nand U19788 (N_19788,N_13612,N_14273);
nor U19789 (N_19789,N_11413,N_13692);
or U19790 (N_19790,N_11565,N_13289);
nand U19791 (N_19791,N_12023,N_10553);
or U19792 (N_19792,N_12087,N_10494);
or U19793 (N_19793,N_14064,N_13569);
xnor U19794 (N_19794,N_13096,N_11898);
and U19795 (N_19795,N_12304,N_14977);
xnor U19796 (N_19796,N_11749,N_14766);
nand U19797 (N_19797,N_14163,N_11907);
and U19798 (N_19798,N_14609,N_13486);
xnor U19799 (N_19799,N_13858,N_13968);
nor U19800 (N_19800,N_13878,N_14414);
nor U19801 (N_19801,N_10923,N_10453);
nand U19802 (N_19802,N_11504,N_11832);
nand U19803 (N_19803,N_13960,N_11833);
and U19804 (N_19804,N_12103,N_10582);
xnor U19805 (N_19805,N_10922,N_10241);
nand U19806 (N_19806,N_13944,N_11095);
xor U19807 (N_19807,N_14289,N_13370);
or U19808 (N_19808,N_11936,N_12500);
nand U19809 (N_19809,N_14151,N_12890);
nor U19810 (N_19810,N_11966,N_10586);
and U19811 (N_19811,N_13807,N_11731);
xor U19812 (N_19812,N_10624,N_14881);
nor U19813 (N_19813,N_13657,N_11435);
nor U19814 (N_19814,N_12954,N_14645);
xor U19815 (N_19815,N_12185,N_12088);
or U19816 (N_19816,N_12065,N_12961);
nand U19817 (N_19817,N_11095,N_11239);
nand U19818 (N_19818,N_12271,N_14083);
nand U19819 (N_19819,N_11151,N_12476);
nand U19820 (N_19820,N_12579,N_11810);
xor U19821 (N_19821,N_11592,N_14514);
and U19822 (N_19822,N_14577,N_13896);
nand U19823 (N_19823,N_14997,N_11672);
nand U19824 (N_19824,N_10225,N_11875);
and U19825 (N_19825,N_12129,N_13474);
nor U19826 (N_19826,N_14699,N_13384);
and U19827 (N_19827,N_10154,N_13240);
and U19828 (N_19828,N_14539,N_11706);
and U19829 (N_19829,N_12019,N_13015);
or U19830 (N_19830,N_13835,N_13483);
nand U19831 (N_19831,N_12016,N_14355);
or U19832 (N_19832,N_13686,N_11888);
xnor U19833 (N_19833,N_10604,N_11144);
or U19834 (N_19834,N_13060,N_11039);
xnor U19835 (N_19835,N_10469,N_13327);
or U19836 (N_19836,N_14791,N_11083);
xor U19837 (N_19837,N_14644,N_13437);
or U19838 (N_19838,N_13668,N_13770);
and U19839 (N_19839,N_13007,N_11952);
xor U19840 (N_19840,N_11294,N_14220);
and U19841 (N_19841,N_12625,N_11577);
or U19842 (N_19842,N_12598,N_13283);
xnor U19843 (N_19843,N_11297,N_14818);
or U19844 (N_19844,N_12433,N_14953);
and U19845 (N_19845,N_10448,N_14600);
xor U19846 (N_19846,N_10872,N_14957);
nand U19847 (N_19847,N_10271,N_14114);
nor U19848 (N_19848,N_10115,N_14721);
xnor U19849 (N_19849,N_13350,N_13790);
or U19850 (N_19850,N_14708,N_13088);
nand U19851 (N_19851,N_14721,N_14239);
nor U19852 (N_19852,N_10965,N_11638);
or U19853 (N_19853,N_14702,N_12582);
xor U19854 (N_19854,N_14336,N_13445);
xor U19855 (N_19855,N_10900,N_14035);
and U19856 (N_19856,N_14659,N_10290);
nand U19857 (N_19857,N_10241,N_14376);
or U19858 (N_19858,N_11587,N_14529);
nand U19859 (N_19859,N_14764,N_14027);
nand U19860 (N_19860,N_11323,N_14909);
nor U19861 (N_19861,N_14316,N_12145);
xor U19862 (N_19862,N_11211,N_14678);
xor U19863 (N_19863,N_12007,N_11033);
or U19864 (N_19864,N_14000,N_11820);
or U19865 (N_19865,N_14593,N_12015);
nand U19866 (N_19866,N_10121,N_11112);
xor U19867 (N_19867,N_10068,N_14128);
or U19868 (N_19868,N_13999,N_10421);
nor U19869 (N_19869,N_13233,N_13815);
and U19870 (N_19870,N_12938,N_13799);
xnor U19871 (N_19871,N_14987,N_12921);
nor U19872 (N_19872,N_13514,N_11581);
or U19873 (N_19873,N_13776,N_12795);
or U19874 (N_19874,N_12307,N_12152);
and U19875 (N_19875,N_11971,N_11368);
xnor U19876 (N_19876,N_11799,N_12726);
nand U19877 (N_19877,N_14076,N_14969);
and U19878 (N_19878,N_11928,N_11930);
or U19879 (N_19879,N_11714,N_14796);
or U19880 (N_19880,N_14617,N_14121);
or U19881 (N_19881,N_11856,N_10698);
nor U19882 (N_19882,N_14011,N_10505);
nor U19883 (N_19883,N_10195,N_12882);
nand U19884 (N_19884,N_11204,N_14075);
and U19885 (N_19885,N_13411,N_14241);
and U19886 (N_19886,N_10150,N_14140);
nand U19887 (N_19887,N_14743,N_12447);
and U19888 (N_19888,N_10450,N_12348);
or U19889 (N_19889,N_14454,N_12214);
or U19890 (N_19890,N_14689,N_12849);
nand U19891 (N_19891,N_10459,N_14650);
nand U19892 (N_19892,N_13030,N_13741);
nand U19893 (N_19893,N_14000,N_11671);
or U19894 (N_19894,N_12662,N_10948);
or U19895 (N_19895,N_10821,N_11327);
and U19896 (N_19896,N_11954,N_13486);
or U19897 (N_19897,N_10379,N_13413);
nand U19898 (N_19898,N_11320,N_14373);
nor U19899 (N_19899,N_13721,N_10729);
nor U19900 (N_19900,N_10907,N_12499);
nand U19901 (N_19901,N_12698,N_13360);
and U19902 (N_19902,N_14424,N_10231);
or U19903 (N_19903,N_13893,N_11071);
nor U19904 (N_19904,N_10306,N_14739);
xnor U19905 (N_19905,N_11010,N_13125);
xnor U19906 (N_19906,N_13287,N_10896);
nand U19907 (N_19907,N_14152,N_11985);
xnor U19908 (N_19908,N_10341,N_13835);
nor U19909 (N_19909,N_13108,N_14109);
xor U19910 (N_19910,N_11913,N_14834);
nand U19911 (N_19911,N_13997,N_14323);
nand U19912 (N_19912,N_11527,N_10556);
nand U19913 (N_19913,N_10985,N_14329);
nand U19914 (N_19914,N_13940,N_10852);
nor U19915 (N_19915,N_13868,N_10146);
nand U19916 (N_19916,N_11170,N_10793);
and U19917 (N_19917,N_12996,N_12812);
or U19918 (N_19918,N_12100,N_14809);
xnor U19919 (N_19919,N_10047,N_13537);
nor U19920 (N_19920,N_14524,N_13913);
and U19921 (N_19921,N_11694,N_13659);
or U19922 (N_19922,N_10750,N_14004);
and U19923 (N_19923,N_10355,N_10560);
and U19924 (N_19924,N_13070,N_10859);
and U19925 (N_19925,N_12297,N_11090);
nand U19926 (N_19926,N_11516,N_12156);
and U19927 (N_19927,N_10179,N_12579);
and U19928 (N_19928,N_10324,N_11087);
or U19929 (N_19929,N_14224,N_14473);
or U19930 (N_19930,N_11548,N_11419);
or U19931 (N_19931,N_12383,N_12323);
nor U19932 (N_19932,N_14579,N_14637);
nand U19933 (N_19933,N_13154,N_14834);
or U19934 (N_19934,N_13922,N_10798);
and U19935 (N_19935,N_11287,N_14294);
nand U19936 (N_19936,N_14528,N_14005);
nor U19937 (N_19937,N_13469,N_10678);
nand U19938 (N_19938,N_10314,N_11114);
nand U19939 (N_19939,N_13159,N_13686);
or U19940 (N_19940,N_11318,N_10049);
xnor U19941 (N_19941,N_13343,N_13543);
and U19942 (N_19942,N_10105,N_14105);
or U19943 (N_19943,N_13954,N_10319);
xor U19944 (N_19944,N_13634,N_12832);
or U19945 (N_19945,N_13915,N_11963);
nand U19946 (N_19946,N_10583,N_13787);
or U19947 (N_19947,N_14212,N_12647);
nor U19948 (N_19948,N_10723,N_12632);
nand U19949 (N_19949,N_13216,N_14398);
xor U19950 (N_19950,N_10199,N_11728);
nand U19951 (N_19951,N_14584,N_14204);
and U19952 (N_19952,N_11361,N_12176);
xnor U19953 (N_19953,N_12942,N_12979);
xnor U19954 (N_19954,N_10679,N_13685);
or U19955 (N_19955,N_13835,N_10434);
nor U19956 (N_19956,N_12928,N_10841);
or U19957 (N_19957,N_13593,N_12233);
nor U19958 (N_19958,N_10418,N_11508);
xor U19959 (N_19959,N_11468,N_11668);
xor U19960 (N_19960,N_12181,N_11065);
or U19961 (N_19961,N_13855,N_13259);
and U19962 (N_19962,N_10006,N_11724);
nor U19963 (N_19963,N_14735,N_13878);
nor U19964 (N_19964,N_10801,N_11611);
and U19965 (N_19965,N_13051,N_14771);
and U19966 (N_19966,N_12989,N_12848);
nand U19967 (N_19967,N_12567,N_13393);
and U19968 (N_19968,N_10932,N_13219);
xnor U19969 (N_19969,N_12894,N_12658);
or U19970 (N_19970,N_14269,N_13583);
xnor U19971 (N_19971,N_10545,N_12665);
nand U19972 (N_19972,N_11668,N_13424);
or U19973 (N_19973,N_11112,N_10017);
xnor U19974 (N_19974,N_10809,N_14639);
and U19975 (N_19975,N_14644,N_13083);
xor U19976 (N_19976,N_13369,N_11913);
nand U19977 (N_19977,N_10087,N_14462);
nand U19978 (N_19978,N_11750,N_10639);
xor U19979 (N_19979,N_13748,N_14075);
xor U19980 (N_19980,N_11229,N_14254);
nand U19981 (N_19981,N_11258,N_14195);
nand U19982 (N_19982,N_11897,N_11564);
nor U19983 (N_19983,N_13428,N_11739);
or U19984 (N_19984,N_12823,N_14426);
nand U19985 (N_19985,N_12371,N_14763);
and U19986 (N_19986,N_10008,N_11747);
and U19987 (N_19987,N_10552,N_13578);
xor U19988 (N_19988,N_10830,N_10046);
or U19989 (N_19989,N_14987,N_14041);
nand U19990 (N_19990,N_14531,N_12459);
or U19991 (N_19991,N_13531,N_14576);
nand U19992 (N_19992,N_14862,N_14788);
or U19993 (N_19993,N_14492,N_11342);
nand U19994 (N_19994,N_13387,N_14199);
nor U19995 (N_19995,N_14084,N_12427);
or U19996 (N_19996,N_11219,N_10660);
or U19997 (N_19997,N_10753,N_14738);
xnor U19998 (N_19998,N_13942,N_10922);
nor U19999 (N_19999,N_10977,N_10218);
or U20000 (N_20000,N_16264,N_16334);
xor U20001 (N_20001,N_19374,N_18303);
or U20002 (N_20002,N_17019,N_16959);
or U20003 (N_20003,N_19140,N_19036);
xor U20004 (N_20004,N_16246,N_16466);
xnor U20005 (N_20005,N_17364,N_18278);
or U20006 (N_20006,N_16924,N_15736);
or U20007 (N_20007,N_15630,N_19984);
xor U20008 (N_20008,N_17874,N_16773);
xnor U20009 (N_20009,N_19006,N_18141);
nor U20010 (N_20010,N_17685,N_18922);
nor U20011 (N_20011,N_15345,N_16428);
xnor U20012 (N_20012,N_19137,N_15330);
xor U20013 (N_20013,N_16446,N_18232);
and U20014 (N_20014,N_19531,N_16853);
or U20015 (N_20015,N_16197,N_19479);
nor U20016 (N_20016,N_18847,N_18364);
or U20017 (N_20017,N_19507,N_16970);
xor U20018 (N_20018,N_18085,N_15378);
nand U20019 (N_20019,N_15390,N_15071);
nand U20020 (N_20020,N_17181,N_18376);
nor U20021 (N_20021,N_19571,N_19841);
and U20022 (N_20022,N_18222,N_18848);
or U20023 (N_20023,N_18290,N_15875);
or U20024 (N_20024,N_19541,N_17054);
nor U20025 (N_20025,N_17039,N_16700);
nand U20026 (N_20026,N_19964,N_16673);
or U20027 (N_20027,N_15165,N_15117);
nand U20028 (N_20028,N_17182,N_16597);
nor U20029 (N_20029,N_18521,N_19183);
xnor U20030 (N_20030,N_15313,N_19121);
xor U20031 (N_20031,N_19124,N_19520);
or U20032 (N_20032,N_15701,N_16003);
nand U20033 (N_20033,N_16694,N_16435);
nand U20034 (N_20034,N_16289,N_17522);
nand U20035 (N_20035,N_19126,N_18515);
nor U20036 (N_20036,N_17286,N_15749);
nor U20037 (N_20037,N_15148,N_15564);
and U20038 (N_20038,N_19999,N_15341);
or U20039 (N_20039,N_19175,N_15191);
nand U20040 (N_20040,N_16838,N_18583);
and U20041 (N_20041,N_17816,N_17305);
nand U20042 (N_20042,N_17830,N_15509);
nor U20043 (N_20043,N_16943,N_17367);
nor U20044 (N_20044,N_19113,N_16769);
and U20045 (N_20045,N_15628,N_18807);
nor U20046 (N_20046,N_16434,N_18211);
nand U20047 (N_20047,N_18787,N_19159);
or U20048 (N_20048,N_17570,N_17701);
xnor U20049 (N_20049,N_18569,N_19280);
or U20050 (N_20050,N_17975,N_15867);
and U20051 (N_20051,N_17949,N_19998);
and U20052 (N_20052,N_15863,N_19264);
or U20053 (N_20053,N_19332,N_19330);
nor U20054 (N_20054,N_15816,N_15942);
or U20055 (N_20055,N_18084,N_18086);
nand U20056 (N_20056,N_16922,N_18946);
nand U20057 (N_20057,N_19189,N_18094);
or U20058 (N_20058,N_17354,N_18355);
xnor U20059 (N_20059,N_16124,N_18554);
nand U20060 (N_20060,N_17130,N_15194);
xnor U20061 (N_20061,N_18872,N_19125);
and U20062 (N_20062,N_18185,N_16307);
and U20063 (N_20063,N_16297,N_16355);
xor U20064 (N_20064,N_15810,N_17251);
and U20065 (N_20065,N_17932,N_18213);
and U20066 (N_20066,N_16699,N_16559);
nand U20067 (N_20067,N_18129,N_18498);
xnor U20068 (N_20068,N_18256,N_17222);
and U20069 (N_20069,N_16238,N_19186);
xnor U20070 (N_20070,N_19007,N_19439);
nor U20071 (N_20071,N_16103,N_15304);
nor U20072 (N_20072,N_15461,N_18941);
nand U20073 (N_20073,N_16114,N_19556);
nor U20074 (N_20074,N_17422,N_15505);
or U20075 (N_20075,N_17024,N_19564);
and U20076 (N_20076,N_19549,N_18754);
xor U20077 (N_20077,N_15203,N_19798);
and U20078 (N_20078,N_17155,N_19711);
and U20079 (N_20079,N_19372,N_15357);
nand U20080 (N_20080,N_15112,N_15529);
nor U20081 (N_20081,N_15394,N_18984);
xor U20082 (N_20082,N_18121,N_19933);
nor U20083 (N_20083,N_17591,N_19995);
nand U20084 (N_20084,N_17191,N_18375);
or U20085 (N_20085,N_16230,N_18448);
or U20086 (N_20086,N_18451,N_17238);
nor U20087 (N_20087,N_16551,N_15737);
nor U20088 (N_20088,N_16933,N_15484);
or U20089 (N_20089,N_17533,N_18683);
xor U20090 (N_20090,N_15488,N_17760);
xor U20091 (N_20091,N_15368,N_18217);
or U20092 (N_20092,N_19793,N_18779);
xor U20093 (N_20093,N_18694,N_16011);
or U20094 (N_20094,N_16634,N_18423);
or U20095 (N_20095,N_17645,N_15985);
xor U20096 (N_20096,N_18116,N_17669);
nand U20097 (N_20097,N_17855,N_19055);
nor U20098 (N_20098,N_18652,N_15632);
xnor U20099 (N_20099,N_19572,N_18926);
nand U20100 (N_20100,N_18408,N_18748);
and U20101 (N_20101,N_19114,N_19821);
nor U20102 (N_20102,N_15075,N_15822);
nor U20103 (N_20103,N_19177,N_18192);
nand U20104 (N_20104,N_18488,N_19211);
xnor U20105 (N_20105,N_17921,N_18876);
or U20106 (N_20106,N_16851,N_15426);
and U20107 (N_20107,N_16412,N_15897);
xnor U20108 (N_20108,N_15236,N_16060);
xnor U20109 (N_20109,N_18246,N_15691);
xor U20110 (N_20110,N_16629,N_16852);
nor U20111 (N_20111,N_17886,N_19757);
nor U20112 (N_20112,N_18273,N_18069);
and U20113 (N_20113,N_15577,N_18861);
xor U20114 (N_20114,N_15472,N_18630);
nor U20115 (N_20115,N_19284,N_16367);
xnor U20116 (N_20116,N_16558,N_18102);
and U20117 (N_20117,N_15901,N_19134);
xor U20118 (N_20118,N_19593,N_17120);
and U20119 (N_20119,N_16732,N_19944);
or U20120 (N_20120,N_17271,N_19528);
xnor U20121 (N_20121,N_17609,N_19018);
nor U20122 (N_20122,N_15387,N_18743);
nor U20123 (N_20123,N_17909,N_18746);
and U20124 (N_20124,N_17508,N_15570);
or U20125 (N_20125,N_15351,N_17982);
nor U20126 (N_20126,N_19804,N_17708);
and U20127 (N_20127,N_17798,N_15187);
xnor U20128 (N_20128,N_18932,N_19930);
nor U20129 (N_20129,N_18467,N_15083);
and U20130 (N_20130,N_18877,N_19890);
or U20131 (N_20131,N_18082,N_16928);
nand U20132 (N_20132,N_15474,N_19288);
xnor U20133 (N_20133,N_17135,N_19588);
xnor U20134 (N_20134,N_16477,N_15731);
nor U20135 (N_20135,N_19973,N_19747);
nand U20136 (N_20136,N_15259,N_15371);
nand U20137 (N_20137,N_16473,N_18471);
nand U20138 (N_20138,N_16479,N_17449);
xnor U20139 (N_20139,N_15693,N_18601);
xnor U20140 (N_20140,N_19468,N_18429);
xnor U20141 (N_20141,N_15413,N_15896);
nand U20142 (N_20142,N_19581,N_18054);
xor U20143 (N_20143,N_15950,N_15626);
and U20144 (N_20144,N_17753,N_17608);
or U20145 (N_20145,N_18764,N_19809);
and U20146 (N_20146,N_17067,N_19522);
xor U20147 (N_20147,N_18666,N_19965);
xor U20148 (N_20148,N_16945,N_16319);
nor U20149 (N_20149,N_19112,N_17193);
nand U20150 (N_20150,N_15802,N_15040);
xor U20151 (N_20151,N_19215,N_19799);
and U20152 (N_20152,N_18130,N_18282);
nor U20153 (N_20153,N_16249,N_19024);
xnor U20154 (N_20154,N_15074,N_15515);
or U20155 (N_20155,N_19828,N_18534);
nand U20156 (N_20156,N_19253,N_15848);
or U20157 (N_20157,N_18917,N_18504);
xnor U20158 (N_20158,N_16211,N_19610);
xor U20159 (N_20159,N_18535,N_16512);
nand U20160 (N_20160,N_15927,N_18188);
nand U20161 (N_20161,N_15066,N_17379);
and U20162 (N_20162,N_16930,N_19101);
xor U20163 (N_20163,N_17291,N_17653);
and U20164 (N_20164,N_18019,N_17820);
xor U20165 (N_20165,N_19393,N_15358);
xnor U20166 (N_20166,N_18600,N_19636);
nand U20167 (N_20167,N_16219,N_15027);
or U20168 (N_20168,N_18604,N_18506);
and U20169 (N_20169,N_15336,N_19153);
nor U20170 (N_20170,N_15121,N_17705);
and U20171 (N_20171,N_16994,N_15939);
xnor U20172 (N_20172,N_15249,N_18293);
and U20173 (N_20173,N_16552,N_18038);
xnor U20174 (N_20174,N_19176,N_15072);
nor U20175 (N_20175,N_17868,N_19248);
nand U20176 (N_20176,N_16887,N_15321);
or U20177 (N_20177,N_16286,N_19945);
or U20178 (N_20178,N_15779,N_17944);
xor U20179 (N_20179,N_16734,N_19081);
or U20180 (N_20180,N_16121,N_17228);
nor U20181 (N_20181,N_16421,N_18938);
or U20182 (N_20182,N_15933,N_17863);
xnor U20183 (N_20183,N_16202,N_18418);
and U20184 (N_20184,N_15686,N_19763);
nor U20185 (N_20185,N_19245,N_16353);
xor U20186 (N_20186,N_16619,N_18551);
nor U20187 (N_20187,N_17757,N_17687);
xnor U20188 (N_20188,N_16173,N_15787);
xor U20189 (N_20189,N_19768,N_19819);
nor U20190 (N_20190,N_15512,N_19040);
nor U20191 (N_20191,N_15712,N_18720);
and U20192 (N_20192,N_18677,N_19260);
or U20193 (N_20193,N_15879,N_17343);
and U20194 (N_20194,N_18316,N_18829);
or U20195 (N_20195,N_16805,N_15553);
nor U20196 (N_20196,N_18356,N_17224);
or U20197 (N_20197,N_17233,N_15924);
nand U20198 (N_20198,N_17761,N_18147);
xor U20199 (N_20199,N_18400,N_17548);
xor U20200 (N_20200,N_18598,N_18280);
or U20201 (N_20201,N_19411,N_18459);
nor U20202 (N_20202,N_19442,N_17903);
xnor U20203 (N_20203,N_18585,N_15354);
and U20204 (N_20204,N_15937,N_16910);
and U20205 (N_20205,N_19139,N_19766);
nand U20206 (N_20206,N_17527,N_18603);
and U20207 (N_20207,N_15962,N_16997);
xor U20208 (N_20208,N_17123,N_16217);
or U20209 (N_20209,N_15852,N_15935);
nand U20210 (N_20210,N_16444,N_16453);
nor U20211 (N_20211,N_18939,N_19613);
and U20212 (N_20212,N_18647,N_15899);
nand U20213 (N_20213,N_16388,N_19417);
nand U20214 (N_20214,N_19046,N_18717);
and U20215 (N_20215,N_18258,N_16074);
nand U20216 (N_20216,N_15297,N_16799);
or U20217 (N_20217,N_17107,N_16102);
and U20218 (N_20218,N_15205,N_17558);
xnor U20219 (N_20219,N_18398,N_18638);
nor U20220 (N_20220,N_17457,N_16413);
xor U20221 (N_20221,N_15756,N_19584);
xor U20222 (N_20222,N_18699,N_15383);
nand U20223 (N_20223,N_16490,N_18715);
nand U20224 (N_20224,N_15558,N_18370);
nor U20225 (N_20225,N_17973,N_17606);
xnor U20226 (N_20226,N_16318,N_18099);
nor U20227 (N_20227,N_18242,N_15380);
nor U20228 (N_20228,N_17817,N_18317);
xor U20229 (N_20229,N_17843,N_16362);
xnor U20230 (N_20230,N_15098,N_18812);
or U20231 (N_20231,N_16979,N_16422);
or U20232 (N_20232,N_17128,N_15680);
xor U20233 (N_20233,N_17235,N_16497);
nand U20234 (N_20234,N_15776,N_17453);
nand U20235 (N_20235,N_15428,N_15561);
xor U20236 (N_20236,N_15716,N_18653);
and U20237 (N_20237,N_18179,N_16361);
nand U20238 (N_20238,N_17276,N_15653);
or U20239 (N_20239,N_15443,N_18046);
nand U20240 (N_20240,N_16690,N_16194);
and U20241 (N_20241,N_16300,N_18049);
or U20242 (N_20242,N_18842,N_19122);
nor U20243 (N_20243,N_17632,N_17226);
xor U20244 (N_20244,N_17517,N_17382);
nand U20245 (N_20245,N_18457,N_17890);
or U20246 (N_20246,N_19827,N_15821);
xnor U20247 (N_20247,N_16092,N_17152);
or U20248 (N_20248,N_17080,N_15690);
or U20249 (N_20249,N_18331,N_19585);
nor U20250 (N_20250,N_17378,N_19906);
and U20251 (N_20251,N_18184,N_17331);
and U20252 (N_20252,N_16235,N_18923);
xnor U20253 (N_20253,N_18750,N_18399);
xor U20254 (N_20254,N_17961,N_18912);
or U20255 (N_20255,N_17742,N_17244);
and U20256 (N_20256,N_18505,N_18070);
or U20257 (N_20257,N_15466,N_15087);
nand U20258 (N_20258,N_19661,N_17802);
and U20259 (N_20259,N_19707,N_19291);
nand U20260 (N_20260,N_15245,N_17791);
and U20261 (N_20261,N_16695,N_18072);
or U20262 (N_20262,N_15140,N_18824);
and U20263 (N_20263,N_15941,N_17582);
and U20264 (N_20264,N_19035,N_19366);
and U20265 (N_20265,N_15439,N_19235);
and U20266 (N_20266,N_19386,N_16964);
xor U20267 (N_20267,N_15361,N_17710);
or U20268 (N_20268,N_17161,N_18416);
nor U20269 (N_20269,N_19348,N_18533);
and U20270 (N_20270,N_15007,N_16956);
or U20271 (N_20271,N_19563,N_16187);
nor U20272 (N_20272,N_15284,N_17002);
nand U20273 (N_20273,N_16200,N_16213);
xor U20274 (N_20274,N_15227,N_17037);
and U20275 (N_20275,N_16332,N_15751);
and U20276 (N_20276,N_15009,N_15433);
xnor U20277 (N_20277,N_16154,N_15328);
xor U20278 (N_20278,N_19912,N_15678);
or U20279 (N_20279,N_16555,N_18560);
nand U20280 (N_20280,N_18675,N_18125);
or U20281 (N_20281,N_15274,N_16643);
xnor U20282 (N_20282,N_17333,N_17147);
nand U20283 (N_20283,N_18987,N_18587);
or U20284 (N_20284,N_15084,N_18319);
nor U20285 (N_20285,N_15424,N_17576);
nand U20286 (N_20286,N_15811,N_15531);
or U20287 (N_20287,N_15835,N_19084);
nand U20288 (N_20288,N_15667,N_19684);
nand U20289 (N_20289,N_17185,N_18526);
xor U20290 (N_20290,N_19025,N_19509);
and U20291 (N_20291,N_15928,N_18367);
and U20292 (N_20292,N_17918,N_18670);
and U20293 (N_20293,N_16537,N_16819);
nand U20294 (N_20294,N_19879,N_15155);
nand U20295 (N_20295,N_18615,N_16188);
xor U20296 (N_20296,N_17316,N_18344);
xor U20297 (N_20297,N_16637,N_18436);
xor U20298 (N_20298,N_19255,N_15959);
xor U20299 (N_20299,N_17882,N_19445);
or U20300 (N_20300,N_16091,N_19013);
nor U20301 (N_20301,N_16886,N_17295);
xnor U20302 (N_20302,N_16609,N_16195);
or U20303 (N_20303,N_16193,N_15535);
xnor U20304 (N_20304,N_19806,N_19225);
nand U20305 (N_20305,N_16645,N_18181);
xnor U20306 (N_20306,N_19170,N_18335);
nand U20307 (N_20307,N_18597,N_17636);
or U20308 (N_20308,N_17599,N_18577);
nand U20309 (N_20309,N_17528,N_16004);
nor U20310 (N_20310,N_16070,N_19166);
nand U20311 (N_20311,N_15992,N_15487);
or U20312 (N_20312,N_19005,N_15499);
nor U20313 (N_20313,N_16765,N_18542);
nor U20314 (N_20314,N_16644,N_18171);
and U20315 (N_20315,N_15715,N_17213);
xnor U20316 (N_20316,N_18480,N_17776);
nand U20317 (N_20317,N_19773,N_15763);
nor U20318 (N_20318,N_19418,N_19862);
nor U20319 (N_20319,N_15683,N_18678);
and U20320 (N_20320,N_15814,N_17472);
xnor U20321 (N_20321,N_17696,N_16939);
xor U20322 (N_20322,N_16849,N_18929);
or U20323 (N_20323,N_15877,N_15685);
nand U20324 (N_20324,N_17952,N_16142);
or U20325 (N_20325,N_16850,N_18351);
nand U20326 (N_20326,N_18701,N_16724);
nand U20327 (N_20327,N_19657,N_15762);
and U20328 (N_20328,N_19491,N_19412);
xnor U20329 (N_20329,N_19835,N_19554);
and U20330 (N_20330,N_19327,N_17427);
nand U20331 (N_20331,N_16824,N_15033);
xnor U20332 (N_20332,N_16082,N_17977);
nand U20333 (N_20333,N_18898,N_19882);
xor U20334 (N_20334,N_15905,N_16271);
and U20335 (N_20335,N_16798,N_19008);
nand U20336 (N_20336,N_19064,N_15659);
nand U20337 (N_20337,N_17160,N_18549);
and U20338 (N_20338,N_15981,N_18101);
or U20339 (N_20339,N_18374,N_17845);
nand U20340 (N_20340,N_15185,N_16483);
or U20341 (N_20341,N_18466,N_18794);
xnor U20342 (N_20342,N_16386,N_18993);
xnor U20343 (N_20343,N_19703,N_15677);
xnor U20344 (N_20344,N_15109,N_16665);
nand U20345 (N_20345,N_19550,N_15807);
or U20346 (N_20346,N_17467,N_16384);
xor U20347 (N_20347,N_17145,N_15291);
nand U20348 (N_20348,N_16547,N_16500);
xor U20349 (N_20349,N_15201,N_15961);
nand U20350 (N_20350,N_17063,N_17461);
nor U20351 (N_20351,N_16076,N_15847);
or U20352 (N_20352,N_16391,N_17571);
xor U20353 (N_20353,N_19041,N_17674);
nor U20354 (N_20354,N_16390,N_15022);
and U20355 (N_20355,N_16302,N_17664);
nand U20356 (N_20356,N_18301,N_17122);
nor U20357 (N_20357,N_19380,N_16430);
nand U20358 (N_20358,N_16431,N_16843);
and U20359 (N_20359,N_18999,N_19343);
or U20360 (N_20360,N_15524,N_17248);
nand U20361 (N_20361,N_18614,N_18059);
nand U20362 (N_20362,N_19487,N_15836);
and U20363 (N_20363,N_19996,N_18500);
or U20364 (N_20364,N_15932,N_18196);
or U20365 (N_20365,N_16398,N_15517);
xnor U20366 (N_20366,N_17389,N_17446);
nand U20367 (N_20367,N_15674,N_15809);
nand U20368 (N_20368,N_15335,N_18636);
nor U20369 (N_20369,N_17311,N_18065);
or U20370 (N_20370,N_16742,N_15419);
or U20371 (N_20371,N_17822,N_19003);
or U20372 (N_20372,N_16977,N_15514);
nand U20373 (N_20373,N_16018,N_18078);
xnor U20374 (N_20374,N_17428,N_17848);
or U20375 (N_20375,N_18843,N_18294);
nand U20376 (N_20376,N_16451,N_15100);
nor U20377 (N_20377,N_18381,N_16941);
or U20378 (N_20378,N_17730,N_18426);
and U20379 (N_20379,N_16298,N_19504);
and U20380 (N_20380,N_19472,N_17081);
or U20381 (N_20381,N_17484,N_18661);
nor U20382 (N_20382,N_16341,N_16876);
nand U20383 (N_20383,N_18163,N_19609);
xor U20384 (N_20384,N_18985,N_17951);
nor U20385 (N_20385,N_17747,N_16782);
and U20386 (N_20386,N_17876,N_18774);
and U20387 (N_20387,N_17448,N_19688);
or U20388 (N_20388,N_18363,N_18570);
or U20389 (N_20389,N_15592,N_16863);
nand U20390 (N_20390,N_16617,N_18839);
nand U20391 (N_20391,N_18863,N_19474);
nand U20392 (N_20392,N_16871,N_19622);
or U20393 (N_20393,N_15469,N_19807);
nor U20394 (N_20394,N_17277,N_15389);
and U20395 (N_20395,N_16581,N_19888);
xnor U20396 (N_20396,N_16761,N_15177);
nor U20397 (N_20397,N_15020,N_18279);
and U20398 (N_20398,N_16972,N_17313);
nand U20399 (N_20399,N_18479,N_17098);
nor U20400 (N_20400,N_17804,N_15833);
nor U20401 (N_20401,N_19246,N_19484);
nor U20402 (N_20402,N_18312,N_19043);
nand U20403 (N_20403,N_15002,N_19949);
or U20404 (N_20404,N_19234,N_16345);
nor U20405 (N_20405,N_16130,N_15161);
nor U20406 (N_20406,N_19130,N_19350);
and U20407 (N_20407,N_19524,N_18803);
and U20408 (N_20408,N_19953,N_19406);
nor U20409 (N_20409,N_19631,N_16952);
nand U20410 (N_20410,N_19664,N_17770);
nand U20411 (N_20411,N_16667,N_17901);
and U20412 (N_20412,N_19252,N_16315);
nand U20413 (N_20413,N_18413,N_18545);
nand U20414 (N_20414,N_19481,N_19325);
xor U20415 (N_20415,N_17841,N_16305);
nand U20416 (N_20416,N_15010,N_15127);
and U20417 (N_20417,N_19494,N_19203);
xnor U20418 (N_20418,N_18739,N_15416);
and U20419 (N_20419,N_15123,N_15591);
nand U20420 (N_20420,N_17989,N_18231);
xor U20421 (N_20421,N_16424,N_16840);
or U20422 (N_20422,N_16086,N_16225);
xor U20423 (N_20423,N_18040,N_17869);
nand U20424 (N_20424,N_16740,N_16636);
or U20425 (N_20425,N_19154,N_17631);
nor U20426 (N_20426,N_19150,N_16073);
nand U20427 (N_20427,N_15050,N_15583);
or U20428 (N_20428,N_19185,N_15507);
nor U20429 (N_20429,N_19922,N_19977);
or U20430 (N_20430,N_17920,N_17082);
nor U20431 (N_20431,N_15983,N_17199);
and U20432 (N_20432,N_18887,N_17041);
or U20433 (N_20433,N_17366,N_19562);
xor U20434 (N_20434,N_17934,N_16990);
nor U20435 (N_20435,N_15889,N_15266);
xnor U20436 (N_20436,N_16632,N_16804);
nor U20437 (N_20437,N_17229,N_19647);
xor U20438 (N_20438,N_18635,N_18024);
and U20439 (N_20439,N_18858,N_15569);
or U20440 (N_20440,N_18618,N_16836);
nor U20441 (N_20441,N_17061,N_19072);
nand U20442 (N_20442,N_18062,N_18202);
xor U20443 (N_20443,N_18673,N_16531);
or U20444 (N_20444,N_16296,N_15502);
xor U20445 (N_20445,N_18080,N_16801);
xnor U20446 (N_20446,N_17117,N_19874);
and U20447 (N_20447,N_15644,N_15940);
nor U20448 (N_20448,N_15790,N_16869);
or U20449 (N_20449,N_18891,N_19143);
nor U20450 (N_20450,N_18414,N_18128);
xnor U20451 (N_20451,N_17959,N_18913);
or U20452 (N_20452,N_17479,N_15202);
nand U20453 (N_20453,N_18836,N_18753);
and U20454 (N_20454,N_16001,N_17698);
nor U20455 (N_20455,N_16671,N_15135);
xnor U20456 (N_20456,N_15228,N_19698);
and U20457 (N_20457,N_17555,N_15042);
xnor U20458 (N_20458,N_18725,N_18291);
or U20459 (N_20459,N_18057,N_19924);
xnor U20460 (N_20460,N_19986,N_15708);
xnor U20461 (N_20461,N_18323,N_16050);
and U20462 (N_20462,N_19270,N_17994);
xnor U20463 (N_20463,N_16656,N_15610);
nand U20464 (N_20464,N_18287,N_18721);
nor U20465 (N_20465,N_18902,N_18266);
nand U20466 (N_20466,N_16462,N_19865);
xnor U20467 (N_20467,N_17827,N_18352);
nand U20468 (N_20468,N_15660,N_19056);
and U20469 (N_20469,N_17772,N_17397);
nand U20470 (N_20470,N_15545,N_17426);
and U20471 (N_20471,N_19453,N_17756);
or U20472 (N_20472,N_16168,N_19093);
and U20473 (N_20473,N_19034,N_16697);
nor U20474 (N_20474,N_19983,N_19843);
nor U20475 (N_20475,N_18048,N_18620);
xor U20476 (N_20476,N_18543,N_17781);
xor U20477 (N_20477,N_16321,N_16115);
nor U20478 (N_20478,N_15543,N_16164);
xnor U20479 (N_20479,N_19508,N_15733);
nand U20480 (N_20480,N_15921,N_16382);
xnor U20481 (N_20481,N_18110,N_18226);
and U20482 (N_20482,N_15520,N_17626);
nor U20483 (N_20483,N_18797,N_16865);
nor U20484 (N_20484,N_17356,N_19221);
or U20485 (N_20485,N_15318,N_19690);
and U20486 (N_20486,N_19920,N_16709);
nand U20487 (N_20487,N_18825,N_16456);
and U20488 (N_20488,N_17391,N_19641);
nor U20489 (N_20489,N_18579,N_15803);
xor U20490 (N_20490,N_16916,N_17071);
nand U20491 (N_20491,N_18074,N_17195);
or U20492 (N_20492,N_15971,N_17168);
or U20493 (N_20493,N_16165,N_16494);
and U20494 (N_20494,N_15021,N_17171);
or U20495 (N_20495,N_15510,N_19050);
nand U20496 (N_20496,N_17394,N_15876);
and U20497 (N_20497,N_16148,N_19178);
nor U20498 (N_20498,N_19765,N_16287);
xor U20499 (N_20499,N_17315,N_15622);
nand U20500 (N_20500,N_17040,N_17588);
or U20501 (N_20501,N_17691,N_15338);
xnor U20502 (N_20502,N_17859,N_17553);
xor U20503 (N_20503,N_15893,N_19846);
nor U20504 (N_20504,N_19448,N_18853);
nand U20505 (N_20505,N_17895,N_18557);
xnor U20506 (N_20506,N_18700,N_19449);
nor U20507 (N_20507,N_15724,N_15056);
xor U20508 (N_20508,N_17690,N_17451);
nor U20509 (N_20509,N_15844,N_17212);
or U20510 (N_20510,N_15748,N_17113);
and U20511 (N_20511,N_18852,N_16602);
nor U20512 (N_20512,N_17287,N_19469);
xor U20513 (N_20513,N_16360,N_18013);
nor U20514 (N_20514,N_17851,N_15222);
and U20515 (N_20515,N_18394,N_15743);
nand U20516 (N_20516,N_16035,N_15976);
nor U20517 (N_20517,N_18210,N_18173);
nor U20518 (N_20518,N_19669,N_19627);
or U20519 (N_20519,N_16088,N_17068);
or U20520 (N_20520,N_19377,N_18894);
or U20521 (N_20521,N_17794,N_17006);
nor U20522 (N_20522,N_17864,N_16816);
nor U20523 (N_20523,N_17188,N_16461);
nor U20524 (N_20524,N_16266,N_17501);
or U20525 (N_20525,N_15679,N_17175);
or U20526 (N_20526,N_18716,N_19937);
nand U20527 (N_20527,N_16504,N_16525);
nand U20528 (N_20528,N_16870,N_19629);
xor U20529 (N_20529,N_19667,N_19870);
nand U20530 (N_20530,N_18237,N_17779);
nand U20531 (N_20531,N_17639,N_15604);
and U20532 (N_20532,N_19340,N_15868);
xor U20533 (N_20533,N_15753,N_17953);
nand U20534 (N_20534,N_18719,N_16338);
xnor U20535 (N_20535,N_16192,N_16855);
nor U20536 (N_20536,N_15996,N_16794);
or U20537 (N_20537,N_15442,N_15200);
and U20538 (N_20538,N_17174,N_15485);
xor U20539 (N_20539,N_19336,N_18711);
and U20540 (N_20540,N_19891,N_15556);
nor U20541 (N_20541,N_18325,N_18823);
nor U20542 (N_20542,N_17675,N_15815);
nor U20543 (N_20543,N_15540,N_17726);
nand U20544 (N_20544,N_16582,N_16470);
xnor U20545 (N_20545,N_19422,N_19743);
xor U20546 (N_20546,N_18248,N_15392);
nor U20547 (N_20547,N_16079,N_17294);
and U20548 (N_20548,N_16839,N_17807);
xor U20549 (N_20549,N_17272,N_18737);
nand U20550 (N_20550,N_18854,N_17624);
nand U20551 (N_20551,N_16628,N_19637);
xnor U20552 (N_20552,N_15858,N_15421);
nor U20553 (N_20553,N_15640,N_18759);
nor U20554 (N_20554,N_18544,N_17129);
and U20555 (N_20555,N_17413,N_19968);
and U20556 (N_20556,N_15843,N_16905);
nand U20557 (N_20557,N_18067,N_15945);
xor U20558 (N_20558,N_16657,N_16590);
and U20559 (N_20559,N_17699,N_18529);
and U20560 (N_20560,N_16781,N_15280);
xnor U20561 (N_20561,N_17262,N_16877);
nand U20562 (N_20562,N_17138,N_19856);
or U20563 (N_20563,N_15648,N_15011);
and U20564 (N_20564,N_15254,N_15740);
or U20565 (N_20565,N_15621,N_16476);
nor U20566 (N_20566,N_16627,N_15555);
nor U20567 (N_20567,N_16043,N_19031);
and U20568 (N_20568,N_16995,N_16987);
nand U20569 (N_20569,N_19415,N_19341);
nand U20570 (N_20570,N_16568,N_17074);
and U20571 (N_20571,N_16514,N_15698);
nand U20572 (N_20572,N_16240,N_15995);
or U20573 (N_20573,N_15589,N_19956);
xnor U20574 (N_20574,N_19497,N_19231);
nor U20575 (N_20575,N_19742,N_16985);
nand U20576 (N_20576,N_19861,N_18684);
or U20577 (N_20577,N_16170,N_15459);
xnor U20578 (N_20578,N_19238,N_18714);
nand U20579 (N_20579,N_18154,N_19000);
nand U20580 (N_20580,N_18150,N_17401);
xnor U20581 (N_20581,N_17414,N_18151);
or U20582 (N_20582,N_15796,N_16036);
and U20583 (N_20583,N_18792,N_17780);
or U20584 (N_20584,N_17505,N_18856);
and U20585 (N_20585,N_15675,N_17787);
and U20586 (N_20586,N_19078,N_16926);
and U20587 (N_20587,N_18369,N_18475);
nor U20588 (N_20588,N_16232,N_15267);
and U20589 (N_20589,N_17601,N_16418);
xor U20590 (N_20590,N_16993,N_16029);
xor U20591 (N_20591,N_19092,N_16817);
nor U20592 (N_20592,N_19447,N_17442);
xnor U20593 (N_20593,N_17715,N_15003);
or U20594 (N_20594,N_18118,N_16196);
and U20595 (N_20595,N_18679,N_17192);
nor U20596 (N_20596,N_15420,N_16134);
nor U20597 (N_20597,N_16660,N_19129);
and U20598 (N_20598,N_16818,N_16346);
nand U20599 (N_20599,N_17557,N_15988);
xnor U20600 (N_20600,N_18305,N_16546);
nand U20601 (N_20601,N_16867,N_16061);
nor U20602 (N_20602,N_19029,N_16138);
nand U20603 (N_20603,N_19076,N_17334);
nor U20604 (N_20604,N_18833,N_18190);
and U20605 (N_20605,N_18873,N_18795);
nand U20606 (N_20606,N_17254,N_15294);
nand U20607 (N_20607,N_16774,N_17751);
and U20608 (N_20608,N_19181,N_17793);
or U20609 (N_20609,N_15830,N_16822);
and U20610 (N_20610,N_17647,N_19794);
nor U20611 (N_20611,N_17940,N_19362);
nand U20612 (N_20612,N_18260,N_15028);
xor U20613 (N_20613,N_16122,N_16374);
nor U20614 (N_20614,N_16358,N_17438);
nand U20615 (N_20615,N_16652,N_16777);
and U20616 (N_20616,N_19868,N_15539);
xor U20617 (N_20617,N_19884,N_17358);
nand U20618 (N_20618,N_17415,N_18435);
or U20619 (N_20619,N_15758,N_17432);
xnor U20620 (N_20620,N_16659,N_19148);
or U20621 (N_20621,N_18042,N_16868);
and U20622 (N_20622,N_19066,N_19837);
nand U20623 (N_20623,N_16010,N_15672);
nand U20624 (N_20624,N_19193,N_16364);
nor U20625 (N_20625,N_15415,N_16691);
or U20626 (N_20626,N_18726,N_19623);
or U20627 (N_20627,N_17482,N_19783);
or U20628 (N_20628,N_17892,N_19536);
and U20629 (N_20629,N_18793,N_15895);
or U20630 (N_20630,N_19699,N_19391);
and U20631 (N_20631,N_17541,N_16185);
nor U20632 (N_20632,N_19344,N_18006);
nand U20633 (N_20633,N_19304,N_16524);
or U20634 (N_20634,N_17143,N_16758);
nor U20635 (N_20635,N_17724,N_17812);
or U20636 (N_20636,N_16357,N_17345);
and U20637 (N_20637,N_17239,N_18509);
nor U20638 (N_20638,N_19401,N_19001);
and U20639 (N_20639,N_19818,N_18474);
and U20640 (N_20640,N_15455,N_16237);
and U20641 (N_20641,N_18052,N_16160);
nor U20642 (N_20642,N_17913,N_19210);
and U20643 (N_20643,N_16743,N_16903);
or U20644 (N_20644,N_18575,N_18806);
nand U20645 (N_20645,N_15004,N_18017);
nor U20646 (N_20646,N_19823,N_15434);
or U20647 (N_20647,N_17106,N_16205);
nand U20648 (N_20648,N_19540,N_15799);
nand U20649 (N_20649,N_16714,N_17324);
and U20650 (N_20650,N_19695,N_16625);
or U20651 (N_20651,N_15106,N_16727);
xor U20652 (N_20652,N_19408,N_19299);
or U20653 (N_20653,N_18329,N_15190);
nor U20654 (N_20654,N_16457,N_17680);
xor U20655 (N_20655,N_15363,N_15695);
or U20656 (N_20656,N_19677,N_19959);
or U20657 (N_20657,N_19526,N_18041);
nand U20658 (N_20658,N_19282,N_18662);
nand U20659 (N_20659,N_16274,N_19392);
or U20660 (N_20660,N_17115,N_16593);
xnor U20661 (N_20661,N_19199,N_19205);
or U20662 (N_20662,N_17854,N_19254);
and U20663 (N_20663,N_15427,N_18334);
nand U20664 (N_20664,N_15316,N_17103);
or U20665 (N_20665,N_15001,N_17418);
nand U20666 (N_20666,N_17385,N_16646);
xor U20667 (N_20667,N_19683,N_16137);
or U20668 (N_20668,N_16911,N_19022);
xor U20669 (N_20669,N_17089,N_15147);
nand U20670 (N_20670,N_19115,N_15436);
and U20671 (N_20671,N_19289,N_19705);
xor U20672 (N_20672,N_19501,N_18326);
xnor U20673 (N_20673,N_16793,N_16376);
xor U20674 (N_20674,N_17306,N_15252);
nand U20675 (N_20675,N_18616,N_16612);
and U20676 (N_20676,N_19744,N_16373);
or U20677 (N_20677,N_19649,N_19313);
nand U20678 (N_20678,N_15256,N_19527);
nor U20679 (N_20679,N_17720,N_19314);
or U20680 (N_20680,N_19503,N_16257);
xor U20681 (N_20681,N_19145,N_15703);
nand U20682 (N_20682,N_17079,N_15242);
and U20683 (N_20683,N_19578,N_17615);
xor U20684 (N_20684,N_18705,N_16991);
and U20685 (N_20685,N_17256,N_18741);
nand U20686 (N_20686,N_15319,N_17942);
xnor U20687 (N_20687,N_19019,N_15322);
nor U20688 (N_20688,N_16125,N_17011);
xnor U20689 (N_20689,N_17341,N_18164);
nor U20690 (N_20690,N_17668,N_18838);
xor U20691 (N_20691,N_16445,N_17219);
xor U20692 (N_20692,N_17497,N_17005);
nor U20693 (N_20693,N_19836,N_19662);
and U20694 (N_20694,N_16212,N_17097);
nor U20695 (N_20695,N_17923,N_17993);
or U20696 (N_20696,N_16680,N_19748);
and U20697 (N_20697,N_19023,N_15960);
and U20698 (N_20698,N_16684,N_17273);
and U20699 (N_20699,N_15887,N_15053);
xnor U20700 (N_20700,N_17360,N_19780);
and U20701 (N_20701,N_15431,N_16379);
and U20702 (N_20702,N_15272,N_15213);
nand U20703 (N_20703,N_15498,N_16767);
and U20704 (N_20704,N_19523,N_17042);
and U20705 (N_20705,N_17568,N_18950);
nand U20706 (N_20706,N_17384,N_19495);
xor U20707 (N_20707,N_18767,N_15215);
nor U20708 (N_20708,N_19734,N_18546);
or U20709 (N_20709,N_18907,N_18931);
nor U20710 (N_20710,N_18669,N_16190);
xnor U20711 (N_20711,N_15170,N_18841);
and U20712 (N_20712,N_16016,N_19652);
and U20713 (N_20713,N_18869,N_18724);
xnor U20714 (N_20714,N_18501,N_16348);
nand U20715 (N_20715,N_17021,N_18773);
and U20716 (N_20716,N_17572,N_19058);
or U20717 (N_20717,N_15523,N_19796);
and U20718 (N_20718,N_16858,N_15552);
and U20719 (N_20719,N_19643,N_17926);
nand U20720 (N_20720,N_19545,N_16006);
and U20721 (N_20721,N_19621,N_19083);
and U20722 (N_20722,N_17309,N_19656);
xor U20723 (N_20723,N_19208,N_17159);
or U20724 (N_20724,N_18327,N_18712);
nand U20725 (N_20725,N_16387,N_19218);
xnor U20726 (N_20726,N_19802,N_17738);
xor U20727 (N_20727,N_15567,N_15574);
nand U20728 (N_20728,N_17883,N_18973);
nor U20729 (N_20729,N_17285,N_15663);
and U20730 (N_20730,N_16496,N_15248);
or U20731 (N_20731,N_17534,N_18953);
nor U20732 (N_20732,N_17792,N_15611);
and U20733 (N_20733,N_19756,N_18930);
nor U20734 (N_20734,N_16436,N_18734);
and U20735 (N_20735,N_18865,N_15955);
nor U20736 (N_20736,N_19376,N_15676);
nor U20737 (N_20737,N_18755,N_15384);
or U20738 (N_20738,N_19351,N_17260);
nor U20739 (N_20739,N_17464,N_17339);
or U20740 (N_20740,N_17470,N_18682);
nand U20741 (N_20741,N_18991,N_19352);
nor U20742 (N_20742,N_16518,N_19419);
and U20743 (N_20743,N_15699,N_17997);
xnor U20744 (N_20744,N_15343,N_17865);
and U20745 (N_20745,N_16340,N_19196);
nand U20746 (N_20746,N_15317,N_19466);
nor U20747 (N_20747,N_16981,N_16226);
nor U20748 (N_20748,N_15578,N_15668);
xor U20749 (N_20749,N_15912,N_18285);
and U20750 (N_20750,N_15448,N_16854);
or U20751 (N_20751,N_18934,N_15969);
and U20752 (N_20752,N_16567,N_18729);
and U20753 (N_20753,N_15627,N_17169);
nand U20754 (N_20754,N_16615,N_17566);
nor U20755 (N_20755,N_19830,N_18183);
or U20756 (N_20756,N_19477,N_16566);
nor U20757 (N_20757,N_15601,N_19551);
xor U20758 (N_20758,N_16516,N_15480);
nor U20759 (N_20759,N_19017,N_17654);
xor U20760 (N_20760,N_16478,N_15379);
nand U20761 (N_20761,N_19831,N_19378);
xor U20762 (N_20762,N_15231,N_16056);
and U20763 (N_20763,N_19885,N_15968);
and U20764 (N_20764,N_15339,N_17469);
xor U20765 (N_20765,N_19319,N_19624);
nor U20766 (N_20766,N_18492,N_18766);
or U20767 (N_20767,N_16055,N_18012);
or U20768 (N_20768,N_19187,N_16077);
nand U20769 (N_20769,N_19758,N_16820);
xor U20770 (N_20770,N_16677,N_18590);
nor U20771 (N_20771,N_19672,N_16735);
or U20772 (N_20772,N_16944,N_18948);
and U20773 (N_20773,N_19939,N_19062);
nor U20774 (N_20774,N_19733,N_18446);
nor U20775 (N_20775,N_16350,N_18397);
nand U20776 (N_20776,N_17308,N_18702);
or U20777 (N_20777,N_19943,N_15572);
nor U20778 (N_20778,N_19316,N_19971);
xor U20779 (N_20779,N_16120,N_18473);
nand U20780 (N_20780,N_19242,N_16180);
nor U20781 (N_20781,N_19214,N_17825);
xor U20782 (N_20782,N_18959,N_18016);
and U20783 (N_20783,N_16108,N_16008);
and U20784 (N_20784,N_15458,N_19816);
or U20785 (N_20785,N_16025,N_19227);
or U20786 (N_20786,N_18360,N_16764);
nor U20787 (N_20787,N_16603,N_17211);
nand U20788 (N_20788,N_17003,N_16658);
nor U20789 (N_20789,N_18942,N_17910);
nand U20790 (N_20790,N_16616,N_16359);
and U20791 (N_20791,N_19037,N_17898);
or U20792 (N_20792,N_18106,N_18623);
nand U20793 (N_20793,N_17866,N_17644);
or U20794 (N_20794,N_16506,N_17475);
nand U20795 (N_20795,N_16795,N_19576);
nand U20796 (N_20796,N_16095,N_18330);
and U20797 (N_20797,N_16965,N_18302);
nand U20798 (N_20798,N_16509,N_17605);
or U20799 (N_20799,N_16464,N_15857);
or U20800 (N_20800,N_17370,N_16809);
xor U20801 (N_20801,N_18021,N_19149);
nor U20802 (N_20802,N_17575,N_16648);
nor U20803 (N_20803,N_15511,N_18728);
or U20804 (N_20804,N_15760,N_17173);
nand U20805 (N_20805,N_17125,N_18550);
nand U20806 (N_20806,N_17985,N_16427);
or U20807 (N_20807,N_18350,N_15471);
xnor U20808 (N_20808,N_16919,N_19848);
and U20809 (N_20809,N_15293,N_17964);
nand U20810 (N_20810,N_19615,N_18229);
nor U20811 (N_20811,N_16813,N_15929);
nand U20812 (N_20812,N_17477,N_15930);
nand U20813 (N_20813,N_18047,N_18760);
nand U20814 (N_20814,N_17767,N_17269);
nor U20815 (N_20815,N_15462,N_17035);
and U20816 (N_20816,N_19709,N_19226);
and U20817 (N_20817,N_16713,N_16688);
or U20818 (N_20818,N_15120,N_16083);
xor U20819 (N_20819,N_16182,N_17880);
xor U20820 (N_20820,N_16974,N_18640);
and U20821 (N_20821,N_15064,N_18919);
and U20822 (N_20822,N_16441,N_15831);
xor U20823 (N_20823,N_15399,N_18168);
nor U20824 (N_20824,N_18690,N_19967);
and U20825 (N_20825,N_19666,N_19552);
nor U20826 (N_20826,N_15808,N_17075);
and U20827 (N_20827,N_17361,N_18850);
nand U20828 (N_20828,N_19180,N_15176);
nand U20829 (N_20829,N_15557,N_17795);
or U20830 (N_20830,N_17310,N_15257);
nand U20831 (N_20831,N_18747,N_16037);
nand U20832 (N_20832,N_17503,N_18434);
nor U20833 (N_20833,N_15059,N_17156);
and U20834 (N_20834,N_19451,N_18637);
xor U20835 (N_20835,N_15300,N_19932);
or U20836 (N_20836,N_19692,N_15755);
nor U20837 (N_20837,N_16682,N_19887);
nor U20838 (N_20838,N_17733,N_19012);
or U20839 (N_20839,N_15367,N_18517);
or U20840 (N_20840,N_19456,N_18238);
and U20841 (N_20841,N_19194,N_17282);
nor U20842 (N_20842,N_15264,N_17278);
nand U20843 (N_20843,N_18113,N_15372);
nor U20844 (N_20844,N_18002,N_17045);
or U20845 (N_20845,N_17537,N_16859);
nand U20846 (N_20846,N_15060,N_18654);
nand U20847 (N_20847,N_16152,N_18868);
nand U20848 (N_20848,N_17808,N_15865);
nand U20849 (N_20849,N_15800,N_17419);
or U20850 (N_20850,N_19829,N_19107);
and U20851 (N_20851,N_19361,N_16007);
nor U20852 (N_20852,N_18341,N_15103);
xor U20853 (N_20853,N_16650,N_17824);
xnor U20854 (N_20854,N_19772,N_16087);
or U20855 (N_20855,N_18304,N_16872);
nand U20856 (N_20856,N_19679,N_17678);
or U20857 (N_20857,N_19957,N_18422);
xor U20858 (N_20858,N_15327,N_19161);
nand U20859 (N_20859,N_19718,N_15477);
and U20860 (N_20860,N_18809,N_17353);
nor U20861 (N_20861,N_16486,N_15587);
xnor U20862 (N_20862,N_15329,N_17111);
or U20863 (N_20863,N_19087,N_19388);
nor U20864 (N_20864,N_17048,N_19070);
or U20865 (N_20865,N_15043,N_15396);
or U20866 (N_20866,N_16806,N_15664);
xor U20867 (N_20867,N_17643,N_19871);
xor U20868 (N_20868,N_18964,N_16005);
nand U20869 (N_20869,N_19570,N_16198);
xnor U20870 (N_20870,N_19881,N_15287);
or U20871 (N_20871,N_19893,N_16178);
xor U20872 (N_20872,N_15094,N_17987);
and U20873 (N_20873,N_16722,N_18758);
nand U20874 (N_20874,N_18849,N_18762);
or U20875 (N_20875,N_15647,N_19749);
and U20876 (N_20876,N_16284,N_15151);
xnor U20877 (N_20877,N_17142,N_18979);
nor U20878 (N_20878,N_19886,N_19397);
or U20879 (N_20879,N_18612,N_17020);
nand U20880 (N_20880,N_19259,N_19068);
nor U20881 (N_20881,N_18512,N_19914);
or U20882 (N_20882,N_17137,N_18386);
nand U20883 (N_20883,N_15183,N_15013);
and U20884 (N_20884,N_19455,N_17164);
and U20885 (N_20885,N_15871,N_17220);
nor U20886 (N_20886,N_17933,N_15710);
xnor U20887 (N_20887,N_17914,N_19604);
and U20888 (N_20888,N_19358,N_16760);
nor U20889 (N_20889,N_15956,N_15468);
nor U20890 (N_20890,N_18472,N_19285);
nor U20891 (N_20891,N_15086,N_19735);
and U20892 (N_20892,N_17405,N_19165);
xnor U20893 (N_20893,N_15532,N_18697);
nand U20894 (N_20894,N_19395,N_17902);
nand U20895 (N_20895,N_17237,N_15376);
xor U20896 (N_20896,N_17487,N_15000);
or U20897 (N_20897,N_16236,N_15373);
xor U20898 (N_20898,N_15522,N_16845);
and U20899 (N_20899,N_18427,N_18576);
nor U20900 (N_20900,N_15097,N_15366);
nor U20901 (N_20901,N_17001,N_19755);
or U20902 (N_20902,N_16247,N_19232);
and U20903 (N_20903,N_18095,N_18483);
nand U20904 (N_20904,N_17437,N_17214);
nor U20905 (N_20905,N_19026,N_17489);
or U20906 (N_20906,N_18034,N_16153);
nor U20907 (N_20907,N_15944,N_16365);
xnor U20908 (N_20908,N_17510,N_17468);
nor U20909 (N_20909,N_18915,N_16179);
and U20910 (N_20910,N_15353,N_19111);
xnor U20911 (N_20911,N_19470,N_18107);
xor U20912 (N_20912,N_19310,N_18814);
nand U20913 (N_20913,N_17957,N_19926);
nor U20914 (N_20914,N_16312,N_18453);
or U20915 (N_20915,N_16044,N_19368);
or U20916 (N_20916,N_15612,N_18822);
and U20917 (N_20917,N_15642,N_17915);
nor U20918 (N_20918,N_17014,N_16208);
and U20919 (N_20919,N_18441,N_17459);
or U20920 (N_20920,N_17149,N_16269);
and U20921 (N_20921,N_18035,N_18402);
and U20922 (N_20922,N_19303,N_16491);
or U20923 (N_20923,N_15116,N_18859);
and U20924 (N_20924,N_17894,N_15402);
xor U20925 (N_20925,N_15303,N_16081);
xor U20926 (N_20926,N_17434,N_16811);
xor U20927 (N_20927,N_18228,N_18980);
and U20928 (N_20928,N_16847,N_19778);
and U20929 (N_20929,N_19459,N_17709);
or U20930 (N_20930,N_19543,N_19452);
and U20931 (N_20931,N_16664,N_16543);
nor U20932 (N_20932,N_15198,N_19240);
nand U20933 (N_20933,N_16611,N_15138);
and U20934 (N_20934,N_19424,N_17059);
nor U20935 (N_20935,N_16698,N_15302);
nor U20936 (N_20936,N_19880,N_18646);
xnor U20937 (N_20937,N_19905,N_18438);
xor U20938 (N_20938,N_19525,N_16280);
and U20939 (N_20939,N_17768,N_15206);
nor U20940 (N_20940,N_18686,N_15128);
xnor U20941 (N_20941,N_17344,N_18063);
nor U20942 (N_20942,N_17759,N_17595);
or U20943 (N_20943,N_17873,N_17066);
nor U20944 (N_20944,N_17186,N_18802);
nand U20945 (N_20945,N_15503,N_18431);
xnor U20946 (N_20946,N_16255,N_19020);
xnor U20947 (N_20947,N_19620,N_16929);
nand U20948 (N_20948,N_15337,N_19274);
nand U20949 (N_20949,N_15842,N_17072);
nand U20950 (N_20950,N_19614,N_17296);
and U20951 (N_20951,N_15902,N_19038);
nor U20952 (N_20952,N_17594,N_16204);
and U20953 (N_20953,N_16827,N_19216);
and U20954 (N_20954,N_16191,N_16881);
or U20955 (N_20955,N_17386,N_15289);
and U20956 (N_20956,N_15687,N_16270);
or U20957 (N_20957,N_19263,N_16203);
xor U20958 (N_20958,N_17655,N_15159);
xor U20959 (N_20959,N_19607,N_17971);
nand U20960 (N_20960,N_15125,N_19590);
nor U20961 (N_20961,N_19207,N_18967);
or U20962 (N_20962,N_19387,N_15037);
xor U20963 (N_20963,N_15785,N_17889);
xnor U20964 (N_20964,N_15966,N_17752);
xor U20965 (N_20965,N_16595,N_15278);
nor U20966 (N_20966,N_16670,N_16574);
or U20967 (N_20967,N_19219,N_19307);
nand U20968 (N_20968,N_17659,N_17410);
or U20969 (N_20969,N_16925,N_16206);
nor U20970 (N_20970,N_18060,N_15717);
xnor U20971 (N_20971,N_19267,N_15364);
nor U20972 (N_20972,N_18425,N_19659);
xnor U20973 (N_20973,N_16263,N_18132);
xnor U20974 (N_20974,N_17663,N_16986);
and U20975 (N_20975,N_16846,N_17180);
and U20976 (N_20976,N_15745,N_16111);
and U20977 (N_20977,N_18338,N_19800);
nand U20978 (N_20978,N_17857,N_19626);
and U20979 (N_20979,N_17666,N_15982);
nor U20980 (N_20980,N_18092,N_17744);
nor U20981 (N_20981,N_19918,N_17706);
and U20982 (N_20982,N_18296,N_16917);
and U20983 (N_20983,N_18834,N_17105);
xnor U20984 (N_20984,N_15819,N_17815);
or U20985 (N_20985,N_19188,N_15006);
nand U20986 (N_20986,N_16322,N_19349);
nand U20987 (N_20987,N_15365,N_19389);
and U20988 (N_20988,N_19565,N_19015);
nand U20989 (N_20989,N_18906,N_18756);
xnor U20990 (N_20990,N_16425,N_17935);
and U20991 (N_20991,N_18487,N_18225);
nand U20992 (N_20992,N_18267,N_15951);
or U20993 (N_20993,N_18605,N_15425);
nand U20994 (N_20994,N_19645,N_17778);
xor U20995 (N_20995,N_17387,N_16901);
or U20996 (N_20996,N_18031,N_16575);
nand U20997 (N_20997,N_18401,N_15320);
nor U20998 (N_20998,N_16482,N_19592);
nand U20999 (N_20999,N_16344,N_17363);
and U21000 (N_21000,N_15101,N_17184);
or U21001 (N_21001,N_15599,N_15451);
nand U21002 (N_21002,N_17697,N_16253);
xor U21003 (N_21003,N_16821,N_18204);
xor U21004 (N_21004,N_17258,N_16787);
or U21005 (N_21005,N_19407,N_17837);
nor U21006 (N_21006,N_18098,N_16465);
nand U21007 (N_21007,N_19190,N_16686);
xor U21008 (N_21008,N_15124,N_19597);
nor U21009 (N_21009,N_15014,N_15464);
nand U21010 (N_21010,N_17618,N_17104);
and U21011 (N_21011,N_15255,N_17514);
and U21012 (N_21012,N_19779,N_16002);
nor U21013 (N_21013,N_17597,N_17986);
and U21014 (N_21014,N_16381,N_19287);
xnor U21015 (N_21015,N_19917,N_18357);
or U21016 (N_21016,N_19764,N_17231);
or U21017 (N_21017,N_16661,N_19867);
and U21018 (N_21018,N_19869,N_16530);
xnor U21019 (N_21019,N_17078,N_18004);
nor U21020 (N_21020,N_17408,N_18406);
xor U21021 (N_21021,N_17612,N_19409);
nand U21022 (N_21022,N_16423,N_19532);
nand U21023 (N_21023,N_19061,N_18900);
or U21024 (N_21024,N_19991,N_18037);
and U21025 (N_21025,N_17732,N_18245);
nor U21026 (N_21026,N_19910,N_17646);
or U21027 (N_21027,N_16561,N_15034);
and U21028 (N_21028,N_17672,N_15314);
or U21029 (N_21029,N_18216,N_16946);
and U21030 (N_21030,N_16989,N_16635);
nand U21031 (N_21031,N_17261,N_17340);
nand U21032 (N_21032,N_17980,N_17215);
or U21033 (N_21033,N_15594,N_18497);
or U21034 (N_21034,N_19152,N_17495);
nand U21035 (N_21035,N_15265,N_18146);
and U21036 (N_21036,N_16862,N_19512);
and U21037 (N_21037,N_15251,N_17455);
nor U21038 (N_21038,N_17703,N_16258);
and U21039 (N_21039,N_19273,N_15562);
xnor U21040 (N_21040,N_19815,N_15375);
or U21041 (N_21041,N_19345,N_17210);
nor U21042 (N_21042,N_15432,N_15344);
xor U21043 (N_21043,N_19859,N_17945);
nor U21044 (N_21044,N_15168,N_15456);
nand U21045 (N_21045,N_17938,N_17454);
or U21046 (N_21046,N_19954,N_15681);
or U21047 (N_21047,N_18783,N_16221);
and U21048 (N_21048,N_19266,N_18315);
xor U21049 (N_21049,N_19762,N_15697);
xor U21050 (N_21050,N_15156,N_16961);
xnor U21051 (N_21051,N_19157,N_18584);
nand U21052 (N_21052,N_17007,N_17856);
xor U21053 (N_21053,N_17010,N_15953);
or U21054 (N_21054,N_16505,N_16529);
xor U21055 (N_21055,N_18252,N_18465);
nand U21056 (N_21056,N_17995,N_15258);
or U21057 (N_21057,N_17362,N_16631);
nand U21058 (N_21058,N_17818,N_15090);
and U21059 (N_21059,N_15350,N_17550);
nand U21060 (N_21060,N_19482,N_16938);
nand U21061 (N_21061,N_19256,N_17052);
nor U21062 (N_21062,N_19931,N_17124);
nand U21063 (N_21063,N_18195,N_16325);
nor U21064 (N_21064,N_16294,N_16394);
and U21065 (N_21065,N_19460,N_16702);
or U21066 (N_21066,N_17424,N_19651);
nor U21067 (N_21067,N_17540,N_17693);
or U21068 (N_21068,N_18440,N_16317);
or U21069 (N_21069,N_19144,N_18055);
and U21070 (N_21070,N_17429,N_16703);
and U21071 (N_21071,N_16329,N_15044);
nand U21072 (N_21072,N_16484,N_17189);
xor U21073 (N_21073,N_18261,N_15360);
nand U21074 (N_21074,N_15805,N_16708);
and U21075 (N_21075,N_19838,N_16109);
nand U21076 (N_21076,N_16469,N_16912);
and U21077 (N_21077,N_18393,N_15920);
and U21078 (N_21078,N_15727,N_19575);
and U21079 (N_21079,N_19731,N_18804);
or U21080 (N_21080,N_17748,N_15309);
nor U21081 (N_21081,N_18244,N_19228);
xor U21082 (N_21082,N_15092,N_19686);
nand U21083 (N_21083,N_18658,N_15246);
nand U21084 (N_21084,N_19787,N_16316);
or U21085 (N_21085,N_18490,N_19184);
nand U21086 (N_21086,N_18998,N_16177);
nor U21087 (N_21087,N_15993,N_17163);
or U21088 (N_21088,N_18194,N_17652);
xor U21089 (N_21089,N_15290,N_19164);
xnor U21090 (N_21090,N_16653,N_18496);
xnor U21091 (N_21091,N_15786,N_15224);
or U21092 (N_21092,N_18161,N_15551);
xor U21093 (N_21093,N_18001,N_19434);
xnor U21094 (N_21094,N_18881,N_18056);
nor U21095 (N_21095,N_15149,N_16149);
nor U21096 (N_21096,N_16802,N_15862);
nand U21097 (N_21097,N_16780,N_15163);
nor U21098 (N_21098,N_19502,N_18949);
or U21099 (N_21099,N_16906,N_19668);
nand U21100 (N_21100,N_19739,N_15947);
or U21101 (N_21101,N_16831,N_16967);
or U21102 (N_21102,N_16260,N_18087);
or U21103 (N_21103,N_15352,N_18482);
xnor U21104 (N_21104,N_16222,N_15918);
or U21105 (N_21105,N_16739,N_19398);
or U21106 (N_21106,N_16753,N_16129);
nor U21107 (N_21107,N_19961,N_15913);
nor U21108 (N_21108,N_15347,N_19907);
nand U21109 (N_21109,N_16966,N_15782);
nor U21110 (N_21110,N_16826,N_16146);
or U21111 (N_21111,N_18088,N_15541);
nor U21112 (N_21112,N_16220,N_19414);
or U21113 (N_21113,N_17616,N_19209);
or U21114 (N_21114,N_16528,N_17322);
nor U21115 (N_21115,N_16707,N_19357);
nor U21116 (N_21116,N_18955,N_19069);
or U21117 (N_21117,N_17937,N_18180);
nor U21118 (N_21118,N_16366,N_19644);
and U21119 (N_21119,N_16172,N_17907);
or U21120 (N_21120,N_17132,N_18254);
nor U21121 (N_21121,N_18944,N_17026);
nand U21122 (N_21122,N_17126,N_15171);
and U21123 (N_21123,N_19243,N_16352);
nor U21124 (N_21124,N_15450,N_15696);
nand U21125 (N_21125,N_15978,N_15547);
xor U21126 (N_21126,N_18707,N_18009);
or U21127 (N_21127,N_19191,N_17101);
xnor U21128 (N_21128,N_19582,N_17267);
or U21129 (N_21129,N_17891,N_16880);
nor U21130 (N_21130,N_18061,N_19151);
nor U21131 (N_21131,N_16649,N_17301);
nand U21132 (N_21132,N_17695,N_16199);
xnor U21133 (N_21133,N_16285,N_16145);
nand U21134 (N_21134,N_19089,N_18751);
and U21135 (N_21135,N_16458,N_17867);
nand U21136 (N_21136,N_16499,N_16923);
nor U21137 (N_21137,N_18404,N_16766);
nor U21138 (N_21138,N_19518,N_18935);
xor U21139 (N_21139,N_17496,N_16015);
xnor U21140 (N_21140,N_15946,N_15714);
xnor U21141 (N_21141,N_19811,N_15614);
xor U21142 (N_21142,N_18207,N_16580);
or U21143 (N_21143,N_19529,N_17564);
or U21144 (N_21144,N_19708,N_18489);
xor U21145 (N_21145,N_19091,N_17421);
nor U21146 (N_21146,N_17661,N_19250);
xor U21147 (N_21147,N_19169,N_16174);
nor U21148 (N_21148,N_17004,N_15305);
xnor U21149 (N_21149,N_19283,N_15494);
nor U21150 (N_21150,N_18905,N_19788);
or U21151 (N_21151,N_17968,N_15694);
nor U21152 (N_21152,N_15196,N_16385);
nand U21153 (N_21153,N_18174,N_15654);
nor U21154 (N_21154,N_17948,N_18952);
or U21155 (N_21155,N_17545,N_18191);
nor U21156 (N_21156,N_19754,N_15491);
or U21157 (N_21157,N_17625,N_18831);
nand U21158 (N_21158,N_16429,N_15882);
and U21159 (N_21159,N_15306,N_19975);
and U21160 (N_21160,N_17832,N_19172);
xor U21161 (N_21161,N_19810,N_17764);
xor U21162 (N_21162,N_18153,N_17209);
nor U21163 (N_21163,N_19390,N_19097);
and U21164 (N_21164,N_19539,N_16229);
nor U21165 (N_21165,N_15910,N_19281);
or U21166 (N_21166,N_19746,N_15204);
nor U21167 (N_21167,N_16209,N_15665);
and U21168 (N_21168,N_17535,N_16042);
nand U21169 (N_21169,N_19577,N_17015);
or U21170 (N_21170,N_16955,N_15704);
nor U21171 (N_21171,N_15931,N_18177);
nor U21172 (N_21172,N_17027,N_15741);
nand U21173 (N_21173,N_16759,N_18884);
or U21174 (N_21174,N_19635,N_17349);
nor U21175 (N_21175,N_19542,N_19839);
xor U21176 (N_21176,N_16400,N_16613);
nand U21177 (N_21177,N_15954,N_15115);
and U21178 (N_21178,N_18896,N_16706);
or U21179 (N_21179,N_17840,N_15571);
xor U21180 (N_21180,N_17774,N_16000);
or U21181 (N_21181,N_16931,N_16958);
nand U21182 (N_21182,N_17337,N_17578);
xnor U21183 (N_21183,N_16757,N_16596);
xnor U21184 (N_21184,N_15325,N_18947);
or U21185 (N_21185,N_16662,N_17133);
or U21186 (N_21186,N_18105,N_17417);
and U21187 (N_21187,N_16443,N_15405);
and U21188 (N_21188,N_19936,N_19701);
xor U21189 (N_21189,N_19100,N_19347);
or U21190 (N_21190,N_16503,N_15602);
and U21191 (N_21191,N_15997,N_17717);
nor U21192 (N_21192,N_16021,N_17221);
or U21193 (N_21193,N_15069,N_15722);
or U21194 (N_21194,N_15990,N_18008);
or U21195 (N_21195,N_16705,N_17485);
or U21196 (N_21196,N_16068,N_19322);
nand U21197 (N_21197,N_19435,N_15038);
nor U21198 (N_21198,N_16085,N_15548);
and U21199 (N_21199,N_15880,N_16184);
or U21200 (N_21200,N_19373,N_19958);
and U21201 (N_21201,N_17392,N_16328);
or U21202 (N_21202,N_15051,N_15813);
and U21203 (N_21203,N_16301,N_19028);
and U21204 (N_21204,N_15818,N_19302);
nor U21205 (N_21205,N_18265,N_16789);
or U21206 (N_21206,N_18978,N_18782);
nand U21207 (N_21207,N_19483,N_16143);
or U21208 (N_21208,N_18770,N_19589);
xnor U21209 (N_21209,N_16587,N_19396);
xnor U21210 (N_21210,N_16571,N_18813);
nor U21211 (N_21211,N_15513,N_15406);
xnor U21212 (N_21212,N_18495,N_15870);
nor U21213 (N_21213,N_19993,N_19853);
nand U21214 (N_21214,N_16866,N_17474);
nand U21215 (N_21215,N_16131,N_15903);
nand U21216 (N_21216,N_18982,N_18940);
and U21217 (N_21217,N_16803,N_16033);
or U21218 (N_21218,N_17202,N_19433);
and U21219 (N_21219,N_15414,N_19601);
nand U21220 (N_21220,N_15884,N_18801);
nand U21221 (N_21221,N_18555,N_15747);
xor U21222 (N_21222,N_18255,N_16563);
xor U21223 (N_21223,N_19364,N_17516);
nor U21224 (N_21224,N_19653,N_16327);
or U21225 (N_21225,N_15046,N_19916);
xor U21226 (N_21226,N_16335,N_15975);
or U21227 (N_21227,N_16642,N_16953);
xnor U21228 (N_21228,N_17225,N_17217);
nand U21229 (N_21229,N_19298,N_15223);
nand U21230 (N_21230,N_17053,N_17118);
or U21231 (N_21231,N_19080,N_18989);
or U21232 (N_21232,N_18580,N_16135);
nor U21233 (N_21233,N_17093,N_17976);
or U21234 (N_21234,N_19425,N_19826);
and U21235 (N_21235,N_19333,N_15023);
xor U21236 (N_21236,N_19416,N_17681);
or U21237 (N_21237,N_16565,N_18966);
or U21238 (N_21238,N_15162,N_16169);
nor U21239 (N_21239,N_18203,N_19244);
and U21240 (N_21240,N_19750,N_19382);
and U21241 (N_21241,N_17375,N_16126);
nor U21242 (N_21242,N_18144,N_17043);
nor U21243 (N_21243,N_15218,N_18971);
nand U21244 (N_21244,N_19457,N_15054);
nand U21245 (N_21245,N_18284,N_15273);
xnor U21246 (N_21246,N_19241,N_18030);
and U21247 (N_21247,N_16304,N_19966);
or U21248 (N_21248,N_17704,N_18007);
nand U21249 (N_21249,N_16101,N_17592);
or U21250 (N_21250,N_18757,N_18281);
nand U21251 (N_21251,N_18513,N_17293);
nor U21252 (N_21252,N_18527,N_18855);
and U21253 (N_21253,N_19265,N_18867);
xnor U21254 (N_21254,N_15629,N_17667);
and U21255 (N_21255,N_16098,N_18218);
nor U21256 (N_21256,N_17236,N_17051);
xnor U21257 (N_21257,N_16272,N_17554);
or U21258 (N_21258,N_19761,N_17763);
nor U21259 (N_21259,N_18419,N_18036);
and U21260 (N_21260,N_16936,N_16167);
xnor U21261 (N_21261,N_18011,N_19671);
nand U21262 (N_21262,N_18921,N_19309);
and U21263 (N_21263,N_18205,N_18241);
nand U21264 (N_21264,N_18974,N_16521);
nand U21265 (N_21265,N_18461,N_15568);
nand U21266 (N_21266,N_19379,N_15492);
nor U21267 (N_21267,N_16156,N_15315);
nor U21268 (N_21268,N_17200,N_16992);
nor U21269 (N_21269,N_18000,N_18644);
nor U21270 (N_21270,N_18167,N_15178);
or U21271 (N_21271,N_16823,N_18988);
nor U21272 (N_21272,N_18227,N_19096);
and U21273 (N_21273,N_17274,N_19612);
or U21274 (N_21274,N_16158,N_18389);
and U21275 (N_21275,N_16161,N_17929);
nand U21276 (N_21276,N_18632,N_16045);
or U21277 (N_21277,N_18114,N_16607);
nand U21278 (N_21278,N_17478,N_17990);
and U21279 (N_21279,N_16578,N_15585);
xnor U21280 (N_21280,N_15062,N_18264);
nor U21281 (N_21281,N_17809,N_15864);
nand U21282 (N_21282,N_15438,N_17242);
nand U21283 (N_21283,N_15119,N_19353);
or U21284 (N_21284,N_16402,N_16584);
xnor U21285 (N_21285,N_19473,N_17374);
or U21286 (N_21286,N_18511,N_18081);
nor U21287 (N_21287,N_16875,N_18540);
xor U21288 (N_21288,N_19860,N_19065);
nand U21289 (N_21289,N_19505,N_15299);
xnor U21290 (N_21290,N_16834,N_17348);
and U21291 (N_21291,N_16896,N_17552);
nor U21292 (N_21292,N_18965,N_16748);
nor U21293 (N_21293,N_16550,N_16927);
nand U21294 (N_21294,N_16681,N_19935);
xor U21295 (N_21295,N_18336,N_15888);
and U21296 (N_21296,N_18650,N_16752);
and U21297 (N_21297,N_17373,N_16276);
nand U21298 (N_21298,N_17598,N_17530);
nor U21299 (N_21299,N_15403,N_16020);
and U21300 (N_21300,N_15114,N_19567);
and U21301 (N_21301,N_19573,N_17922);
or U21302 (N_21302,N_16013,N_19318);
xnor U21303 (N_21303,N_17785,N_18574);
and U21304 (N_21304,N_17250,N_16127);
xnor U21305 (N_21305,N_17140,N_16730);
and U21306 (N_21306,N_18909,N_16583);
and U21307 (N_21307,N_18383,N_15774);
xor U21308 (N_21308,N_16784,N_17297);
xor U21309 (N_21309,N_16022,N_17800);
and U21310 (N_21310,N_18706,N_19405);
nand U21311 (N_21311,N_18651,N_15537);
nand U21312 (N_21312,N_16250,N_15342);
xnor U21313 (N_21313,N_15221,N_19014);
nand U21314 (N_21314,N_16363,N_19952);
or U21315 (N_21315,N_16408,N_17544);
or U21316 (N_21316,N_17897,N_19611);
or U21317 (N_21317,N_16075,N_16279);
nand U21318 (N_21318,N_16119,N_19702);
or U21319 (N_21319,N_19365,N_16026);
or U21320 (N_21320,N_16833,N_18547);
or U21321 (N_21321,N_16751,N_18075);
nand U21322 (N_21322,N_19646,N_19321);
nor U21323 (N_21323,N_15144,N_16522);
and U21324 (N_21324,N_16526,N_17783);
xor U21325 (N_21325,N_16474,N_17247);
or U21326 (N_21326,N_17187,N_15783);
and U21327 (N_21327,N_18201,N_15260);
nand U21328 (N_21328,N_19293,N_15655);
or U21329 (N_21329,N_18866,N_19198);
nand U21330 (N_21330,N_15768,N_18117);
and U21331 (N_21331,N_15388,N_18520);
nand U21332 (N_21332,N_16771,N_15232);
nor U21333 (N_21333,N_19682,N_19311);
and U21334 (N_21334,N_17617,N_19258);
nor U21335 (N_21335,N_17150,N_15700);
nor U21336 (N_21336,N_19402,N_16663);
or U21337 (N_21337,N_15096,N_15501);
and U21338 (N_21338,N_16654,N_15559);
nor U21339 (N_21339,N_18676,N_16467);
nand U21340 (N_21340,N_19042,N_19195);
or U21341 (N_21341,N_18337,N_16861);
nand U21342 (N_21342,N_16104,N_16538);
and U21343 (N_21343,N_18688,N_16779);
xnor U21344 (N_21344,N_17218,N_16569);
nor U21345 (N_21345,N_18874,N_19928);
or U21346 (N_21346,N_18663,N_17162);
xor U21347 (N_21347,N_17729,N_15820);
nand U21348 (N_21348,N_15973,N_17613);
nand U21349 (N_21349,N_18808,N_17488);
nor U21350 (N_21350,N_18961,N_15355);
nand U21351 (N_21351,N_17058,N_15195);
or U21352 (N_21352,N_15067,N_16701);
or U21353 (N_21353,N_18077,N_16556);
or U21354 (N_21354,N_19088,N_15295);
nor U21355 (N_21355,N_18805,N_19663);
or U21356 (N_21356,N_17057,N_19463);
xor U21357 (N_21357,N_15226,N_18920);
nand U21358 (N_21358,N_15334,N_17547);
and U21359 (N_21359,N_18541,N_15702);
nor U21360 (N_21360,N_15262,N_18450);
nor U21361 (N_21361,N_19337,N_16570);
nand U21362 (N_21362,N_16420,N_18449);
nor U21363 (N_21363,N_16333,N_17318);
and U21364 (N_21364,N_16532,N_19493);
xor U21365 (N_21365,N_16339,N_15772);
nor U21366 (N_21366,N_19237,N_18879);
or U21367 (N_21367,N_17999,N_18468);
nor U21368 (N_21368,N_17243,N_16372);
or U21369 (N_21369,N_18916,N_19173);
or U21370 (N_21370,N_16132,N_15605);
nand U21371 (N_21371,N_19478,N_17288);
nand U21372 (N_21372,N_19855,N_16788);
nor U21373 (N_21373,N_16066,N_15943);
and U21374 (N_21374,N_19833,N_19271);
and U21375 (N_21375,N_17718,N_19847);
and U21376 (N_21376,N_17877,N_16403);
and U21377 (N_21377,N_19678,N_17018);
nand U21378 (N_21378,N_16281,N_15478);
nand U21379 (N_21379,N_17381,N_16492);
nand U21380 (N_21380,N_15656,N_18485);
xor U21381 (N_21381,N_17095,N_15331);
nand U21382 (N_21382,N_16920,N_16401);
or U21383 (N_21383,N_16604,N_17369);
nor U21384 (N_21384,N_17640,N_19824);
or U21385 (N_21385,N_17395,N_18538);
and U21386 (N_21386,N_18003,N_19557);
xnor U21387 (N_21387,N_18689,N_17805);
nor U21388 (N_21388,N_15590,N_16594);
nand U21389 (N_21389,N_18589,N_15504);
nand U21390 (N_21390,N_16096,N_15174);
xor U21391 (N_21391,N_19685,N_15029);
or U21392 (N_21392,N_16268,N_15948);
nor U21393 (N_21393,N_18391,N_15519);
nor U21394 (N_21394,N_17665,N_17906);
xnor U21395 (N_21395,N_19099,N_15597);
or U21396 (N_21396,N_16378,N_17801);
and U21397 (N_21397,N_17323,N_17621);
and U21398 (N_21398,N_15078,N_18108);
nand U21399 (N_21399,N_18083,N_19737);
nor U21400 (N_21400,N_17589,N_18157);
nor U21401 (N_21401,N_19976,N_18857);
or U21402 (N_21402,N_15777,N_15934);
or U21403 (N_21403,N_18780,N_19689);
nor U21404 (N_21404,N_16940,N_17198);
nand U21405 (N_21405,N_16144,N_16216);
or U21406 (N_21406,N_19660,N_18778);
nor U21407 (N_21407,N_15310,N_18169);
xnor U21408 (N_21408,N_17694,N_17604);
or U21409 (N_21409,N_18648,N_18039);
xor U21410 (N_21410,N_17728,N_18142);
and U21411 (N_21411,N_17371,N_18358);
or U21412 (N_21412,N_15917,N_18395);
or U21413 (N_21413,N_18452,N_15238);
or U21414 (N_21414,N_18882,N_15609);
nor U21415 (N_21415,N_17131,N_18396);
and U21416 (N_21416,N_16591,N_18424);
nor U21417 (N_21417,N_18781,N_18481);
xnor U21418 (N_21418,N_17862,N_17245);
or U21419 (N_21419,N_16231,N_16349);
or U21420 (N_21420,N_15441,N_15240);
nor U21421 (N_21421,N_18206,N_16057);
and U21422 (N_21422,N_17264,N_18958);
xor U21423 (N_21423,N_18433,N_15349);
nor U21424 (N_21424,N_17569,N_18268);
xnor U21425 (N_21425,N_16256,N_19086);
xnor U21426 (N_21426,N_15457,N_16885);
nor U21427 (N_21427,N_17919,N_17091);
or U21428 (N_21428,N_15770,N_19825);
nor U21429 (N_21429,N_19305,N_19127);
and U21430 (N_21430,N_15192,N_15841);
and U21431 (N_21431,N_17603,N_19712);
nor U21432 (N_21432,N_16323,N_18249);
and U21433 (N_21433,N_17565,N_19938);
xor U21434 (N_21434,N_17740,N_15230);
or U21435 (N_21435,N_18346,N_17492);
nand U21436 (N_21436,N_18657,N_15730);
nor U21437 (N_21437,N_15209,N_18996);
xor U21438 (N_21438,N_15861,N_18595);
or U21439 (N_21439,N_17725,N_19275);
and U21440 (N_21440,N_18983,N_15045);
and U21441 (N_21441,N_19548,N_16063);
xor U21442 (N_21442,N_18639,N_19223);
nor U21443 (N_21443,N_15643,N_19960);
nor U21444 (N_21444,N_19011,N_17879);
or U21445 (N_21445,N_16749,N_19384);
nand U21446 (N_21446,N_15160,N_19619);
xor U21447 (N_21447,N_15393,N_16902);
xor U21448 (N_21448,N_15193,N_17203);
nand U21449 (N_21449,N_18382,N_18275);
or U21450 (N_21450,N_15641,N_18761);
nor U21451 (N_21451,N_18274,N_19053);
xnor U21452 (N_21452,N_18775,N_17518);
nor U21453 (N_21453,N_15214,N_19446);
xor U21454 (N_21454,N_18723,N_17871);
and U21455 (N_21455,N_17543,N_18076);
xnor U21456 (N_21456,N_16027,N_18656);
xor U21457 (N_21457,N_19360,N_15217);
nand U21458 (N_21458,N_15277,N_17828);
or U21459 (N_21459,N_15922,N_19694);
nand U21460 (N_21460,N_15613,N_19832);
nor U21461 (N_21461,N_18800,N_18885);
and U21462 (N_21462,N_17719,N_17602);
xnor U21463 (N_21463,N_18339,N_18786);
nor U21464 (N_21464,N_16259,N_15031);
nor U21465 (N_21465,N_18532,N_16554);
and U21466 (N_21466,N_18668,N_15839);
xor U21467 (N_21467,N_17549,N_19510);
xnor U21468 (N_21468,N_15199,N_16988);
nor U21469 (N_21469,N_16028,N_19410);
nor U21470 (N_21470,N_19752,N_18491);
xnor U21471 (N_21471,N_17462,N_17789);
or U21472 (N_21472,N_17398,N_15666);
nand U21473 (N_21473,N_17773,N_16878);
xor U21474 (N_21474,N_17954,N_16687);
xor U21475 (N_21475,N_19229,N_16356);
xor U21476 (N_21476,N_16797,N_17567);
nor U21477 (N_21477,N_19903,N_15598);
nand U21478 (N_21478,N_16982,N_16975);
or U21479 (N_21479,N_16715,N_19714);
xor U21480 (N_21480,N_18043,N_19736);
nor U21481 (N_21481,N_17542,N_17593);
nor U21482 (N_21482,N_17289,N_18262);
xor U21483 (N_21483,N_17300,N_17500);
or U21484 (N_21484,N_17491,N_18347);
and U21485 (N_21485,N_19367,N_18165);
xor U21486 (N_21486,N_19538,N_19403);
or U21487 (N_21487,N_18862,N_15497);
and U21488 (N_21488,N_17034,N_19331);
and U21489 (N_21489,N_18139,N_19834);
nand U21490 (N_21490,N_18870,N_17326);
nor U21491 (N_21491,N_15422,N_17833);
xnor U21492 (N_21492,N_15952,N_17268);
and U21493 (N_21493,N_15243,N_15624);
xor U21494 (N_21494,N_15906,N_18525);
and U21495 (N_21495,N_16369,N_17486);
and U21496 (N_21496,N_16856,N_19717);
xnor U21497 (N_21497,N_17433,N_16410);
xor U21498 (N_21498,N_17743,N_19044);
nand U21499 (N_21499,N_18430,N_17090);
nor U21500 (N_21500,N_16155,N_18199);
nor U21501 (N_21501,N_15661,N_15283);
nor U21502 (N_21502,N_15618,N_15356);
nor U21503 (N_21503,N_19399,N_16949);
nor U21504 (N_21504,N_19513,N_17523);
or U21505 (N_21505,N_17240,N_15019);
and U21506 (N_21506,N_17574,N_18649);
or U21507 (N_21507,N_19864,N_17481);
nor U21508 (N_21508,N_16389,N_18558);
and U21509 (N_21509,N_18090,N_17580);
nand U21510 (N_21510,N_17754,N_19440);
or U21511 (N_21511,N_17811,N_16078);
nand U21512 (N_21512,N_17166,N_17465);
nor U21513 (N_21513,N_16890,N_17102);
nand U21514 (N_21514,N_19437,N_15732);
nand U21515 (N_21515,N_16183,N_18776);
nand U21516 (N_21516,N_16726,N_16770);
or U21517 (N_21517,N_18565,N_15650);
and U21518 (N_21518,N_17702,N_18409);
or U21519 (N_21519,N_19420,N_17259);
nand U21520 (N_21520,N_19476,N_17887);
xor U21521 (N_21521,N_18464,N_15411);
and U21522 (N_21522,N_15039,N_16455);
xnor U21523 (N_21523,N_19338,N_17416);
and U21524 (N_21524,N_15476,N_18126);
or U21525 (N_21525,N_16589,N_19521);
nor U21526 (N_21526,N_19687,N_15657);
nand U21527 (N_21527,N_19795,N_17197);
xnor U21528 (N_21528,N_17941,N_15965);
xnor U21529 (N_21529,N_15625,N_17821);
nand U21530 (N_21530,N_19454,N_15490);
xor U21531 (N_21531,N_18200,N_17896);
nor U21532 (N_21532,N_18744,N_17190);
and U21533 (N_21533,N_16299,N_15068);
xor U21534 (N_21534,N_17852,N_16879);
and U21535 (N_21535,N_16825,N_16894);
xor U21536 (N_21536,N_17651,N_19638);
or U21537 (N_21537,N_19568,N_19925);
xor U21538 (N_21538,N_19131,N_16303);
and U21539 (N_21539,N_15104,N_19032);
xor U21540 (N_21540,N_17266,N_16900);
nor U21541 (N_21541,N_17939,N_17112);
xor U21542 (N_21542,N_18611,N_15845);
nand U21543 (N_21543,N_15113,N_17494);
nand U21544 (N_21544,N_16405,N_18112);
nand U21545 (N_21545,N_16622,N_18476);
nand U21546 (N_21546,N_19574,N_16588);
nor U21547 (N_21547,N_17788,N_16468);
nor U21548 (N_21548,N_16741,N_16808);
nor U21549 (N_21549,N_17483,N_17539);
and U21550 (N_21550,N_19247,N_16432);
and U21551 (N_21551,N_18020,N_15892);
or U21552 (N_21552,N_16058,N_18796);
or U21553 (N_21553,N_17532,N_15662);
and U21554 (N_21554,N_19278,N_17493);
and U21555 (N_21555,N_15974,N_16937);
nand U21556 (N_21556,N_16954,N_16717);
xor U21557 (N_21557,N_16041,N_17044);
nand U21558 (N_21558,N_16140,N_16630);
xnor U21559 (N_21559,N_16893,N_16054);
nand U21560 (N_21560,N_16935,N_18160);
and U21561 (N_21561,N_19300,N_17443);
and U21562 (N_21562,N_15925,N_15804);
and U21563 (N_21563,N_17444,N_15362);
or U21564 (N_21564,N_17025,N_17936);
and U21565 (N_21565,N_19201,N_16676);
nand U21566 (N_21566,N_17144,N_16639);
or U21567 (N_21567,N_16397,N_19876);
and U21568 (N_21568,N_18263,N_15024);
and U21569 (N_21569,N_16023,N_15671);
or U21570 (N_21570,N_19517,N_15047);
and U21571 (N_21571,N_18969,N_16228);
nand U21572 (N_21572,N_16052,N_16501);
xnor U21573 (N_21573,N_15989,N_16117);
and U21574 (N_21574,N_17755,N_15311);
and U21575 (N_21575,N_18442,N_17771);
nor U21576 (N_21576,N_19569,N_16579);
nor U21577 (N_21577,N_15771,N_18573);
or U21578 (N_21578,N_16414,N_15761);
nand U21579 (N_21579,N_15878,N_18631);
nand U21580 (N_21580,N_19919,N_16883);
or U21581 (N_21581,N_17875,N_19436);
nand U21582 (N_21582,N_18366,N_17782);
nand U21583 (N_21583,N_15651,N_18621);
or U21584 (N_21584,N_15834,N_15711);
and U21585 (N_21585,N_17739,N_16539);
xor U21586 (N_21586,N_18120,N_17983);
and U21587 (N_21587,N_18607,N_18709);
nor U21588 (N_21588,N_16320,N_16776);
nor U21589 (N_21589,N_17357,N_18572);
or U21590 (N_21590,N_17290,N_15081);
nand U21591 (N_21591,N_18910,N_19394);
nand U21592 (N_21592,N_19982,N_17445);
and U21593 (N_21593,N_18152,N_18889);
nand U21594 (N_21594,N_17838,N_16489);
nand U21595 (N_21595,N_16971,N_15575);
and U21596 (N_21596,N_18322,N_19781);
nand U21597 (N_21597,N_16778,N_16651);
nor U21598 (N_21598,N_18655,N_15102);
xnor U21599 (N_21599,N_18407,N_15767);
nand U21600 (N_21600,N_16577,N_15586);
nand U21601 (N_21601,N_16133,N_16884);
or U21602 (N_21602,N_17504,N_18447);
or U21603 (N_21603,N_17476,N_17529);
and U21604 (N_21604,N_19236,N_16592);
nand U21605 (N_21605,N_18539,N_15110);
or U21606 (N_21606,N_18799,N_18819);
xnor U21607 (N_21607,N_18997,N_17506);
nor U21608 (N_21608,N_17033,N_17303);
nor U21609 (N_21609,N_16626,N_17777);
or U21610 (N_21610,N_19370,N_16480);
nor U21611 (N_21611,N_16097,N_19054);
or U21612 (N_21612,N_18659,N_17819);
xor U21613 (N_21613,N_16624,N_17947);
or U21614 (N_21614,N_19033,N_19317);
and U21615 (N_21615,N_17671,N_19295);
xor U21616 (N_21616,N_16553,N_19784);
and U21617 (N_21617,N_18788,N_16306);
nand U21618 (N_21618,N_17365,N_19820);
nor U21619 (N_21619,N_16291,N_19004);
nor U21620 (N_21620,N_16599,N_19617);
or U21621 (N_21621,N_17581,N_19985);
or U21622 (N_21622,N_16562,N_17073);
nor U21623 (N_21623,N_15234,N_16475);
nor U21624 (N_21624,N_18359,N_17393);
xnor U21625 (N_21625,N_16899,N_19639);
and U21626 (N_21626,N_16791,N_18469);
and U21627 (N_21627,N_19048,N_17737);
xor U21628 (N_21628,N_18586,N_19082);
and U21629 (N_21629,N_19981,N_15440);
or U21630 (N_21630,N_19174,N_19426);
nor U21631 (N_21631,N_16210,N_17336);
nand U21632 (N_21632,N_15250,N_17136);
xnor U21633 (N_21633,N_16842,N_16371);
or U21634 (N_21634,N_19693,N_16915);
xnor U21635 (N_21635,N_16347,N_17076);
nor U21636 (N_21636,N_17979,N_19051);
nor U21637 (N_21637,N_17167,N_18115);
or U21638 (N_21638,N_19770,N_15359);
xnor U21639 (N_21639,N_16059,N_19950);
and U21640 (N_21640,N_19427,N_18908);
or U21641 (N_21641,N_17727,N_18548);
and U21642 (N_21642,N_18053,N_18384);
xnor U21643 (N_21643,N_15754,N_16815);
or U21644 (N_21644,N_16755,N_18960);
nor U21645 (N_21645,N_15475,N_17946);
xnor U21646 (N_21646,N_15923,N_18321);
and U21647 (N_21647,N_16608,N_18977);
and U21648 (N_21648,N_17314,N_15705);
and U21649 (N_21649,N_17686,N_18622);
or U21650 (N_21650,N_19990,N_16248);
and U21651 (N_21651,N_15449,N_15239);
nand U21652 (N_21652,N_19123,N_16621);
and U21653 (N_21653,N_17148,N_15576);
and U21654 (N_21654,N_19923,N_15637);
and U21655 (N_21655,N_18209,N_15225);
nand U21656 (N_21656,N_15916,N_15052);
and U21657 (N_21657,N_17965,N_17050);
nor U21658 (N_21658,N_18563,N_18508);
and U21659 (N_21659,N_17590,N_18828);
xor U21660 (N_21660,N_19320,N_17596);
xor U21661 (N_21661,N_19108,N_15400);
nand U21662 (N_21662,N_16215,N_19413);
and U21663 (N_21663,N_18283,N_19167);
xor U21664 (N_21664,N_17194,N_17963);
and U21665 (N_21665,N_15131,N_17151);
or U21666 (N_21666,N_16510,N_19292);
and U21667 (N_21667,N_19315,N_15603);
nor U21668 (N_21668,N_18236,N_19212);
or U21669 (N_21669,N_18602,N_15914);
or U21670 (N_21670,N_16737,N_17056);
or U21671 (N_21671,N_19817,N_16996);
nand U21672 (N_21672,N_16330,N_19480);
nand U21673 (N_21673,N_16738,N_19138);
xor U21674 (N_21674,N_16725,N_17607);
and U21675 (N_21675,N_15088,N_17925);
and U21676 (N_21676,N_18893,N_17587);
and U21677 (N_21677,N_19063,N_19110);
nand U21678 (N_21678,N_16110,N_19987);
or U21679 (N_21679,N_17031,N_19913);
xor U21680 (N_21680,N_17441,N_17662);
xnor U21681 (N_21681,N_16176,N_16375);
nor U21682 (N_21682,N_15798,N_19602);
and U21683 (N_21683,N_18562,N_19775);
or U21684 (N_21684,N_17252,N_17038);
xor U21685 (N_21685,N_17861,N_19908);
or U21686 (N_21686,N_19132,N_18187);
xor U21687 (N_21687,N_17352,N_18771);
nor U21688 (N_21688,N_15057,N_19897);
or U21689 (N_21689,N_19738,N_19633);
xor U21690 (N_21690,N_15298,N_16689);
or U21691 (N_21691,N_18111,N_17711);
nand U21692 (N_21692,N_18552,N_16406);
nor U21693 (N_21693,N_16162,N_15801);
or U21694 (N_21694,N_17846,N_16175);
or U21695 (N_21695,N_19675,N_18840);
nand U21696 (N_21696,N_18288,N_19490);
and U21697 (N_21697,N_17321,N_17641);
nor U21698 (N_21698,N_16038,N_15018);
nor U21699 (N_21699,N_19462,N_16039);
nor U21700 (N_21700,N_18749,N_19335);
nor U21701 (N_21701,N_19458,N_16786);
xor U21702 (N_21702,N_18189,N_15429);
xor U21703 (N_21703,N_16090,N_18066);
nor U21704 (N_21704,N_18903,N_17176);
nor U21705 (N_21705,N_18166,N_15619);
nand U21706 (N_21706,N_16396,N_18703);
xnor U21707 (N_21707,N_19423,N_19090);
nor U21708 (N_21708,N_16331,N_18519);
nand U21709 (N_21709,N_16207,N_18410);
and U21710 (N_21710,N_17383,N_18826);
or U21711 (N_21711,N_16511,N_16273);
and U21712 (N_21712,N_18951,N_16136);
and U21713 (N_21713,N_19721,N_19200);
nand U21714 (N_21714,N_16452,N_15744);
and U21715 (N_21715,N_19857,N_15166);
xnor U21716 (N_21716,N_15134,N_17473);
and U21717 (N_21717,N_15719,N_16605);
or U21718 (N_21718,N_18247,N_18933);
or U21719 (N_21719,N_17399,N_18058);
and U21720 (N_21720,N_15323,N_16572);
xor U21721 (N_21721,N_15623,N_15016);
or U21722 (N_21722,N_17577,N_15145);
xnor U21723 (N_21723,N_18170,N_19230);
nand U21724 (N_21724,N_17177,N_19354);
xnor U21725 (N_21725,N_17956,N_18954);
nand U21726 (N_21726,N_15797,N_19261);
nand U21727 (N_21727,N_16309,N_15538);
and U21728 (N_21728,N_18415,N_16719);
and U21729 (N_21729,N_16310,N_18990);
xnor U21730 (N_21730,N_16051,N_16336);
or U21731 (N_21731,N_19710,N_19767);
and U21732 (N_21732,N_15970,N_15634);
or U21733 (N_21733,N_17707,N_15180);
or U21734 (N_21734,N_17154,N_16241);
nor U21735 (N_21735,N_16342,N_16728);
or U21736 (N_21736,N_17253,N_17292);
and U21737 (N_21737,N_16549,N_15991);
nand U21738 (N_21738,N_17388,N_17984);
nand U21739 (N_21739,N_19312,N_15669);
or U21740 (N_21740,N_17172,N_19515);
or U21741 (N_21741,N_16951,N_16536);
nand U21742 (N_21742,N_18220,N_16669);
nand U21743 (N_21743,N_18470,N_19600);
or U21744 (N_21744,N_18681,N_19706);
nand U21745 (N_21745,N_16750,N_17347);
and U21746 (N_21746,N_17630,N_17786);
or U21747 (N_21747,N_16437,N_19791);
or U21748 (N_21748,N_19814,N_17775);
nand U21749 (N_21749,N_16873,N_15579);
and U21750 (N_21750,N_15435,N_16947);
xor U21751 (N_21751,N_19027,N_18911);
xor U21752 (N_21752,N_18992,N_18276);
xor U21753 (N_21753,N_19955,N_17390);
xor U21754 (N_21754,N_16573,N_19940);
nand U21755 (N_21755,N_18198,N_19142);
nand U21756 (N_21756,N_17682,N_19369);
and U21757 (N_21757,N_17320,N_17814);
or U21758 (N_21758,N_17899,N_18567);
and U21759 (N_21759,N_17046,N_18328);
nor U21760 (N_21760,N_15964,N_17981);
nor U21761 (N_21761,N_15593,N_16262);
and U21762 (N_21762,N_15829,N_16067);
and U21763 (N_21763,N_19075,N_19141);
and U21764 (N_21764,N_17796,N_19769);
nor U21765 (N_21765,N_19894,N_17526);
nor U21766 (N_21766,N_19989,N_15900);
or U21767 (N_21767,N_19895,N_18271);
or U21768 (N_21768,N_16064,N_15153);
nor U21769 (N_21769,N_19962,N_18531);
nand U21770 (N_21770,N_16460,N_18310);
or U21771 (N_21771,N_15890,N_15158);
nand U21772 (N_21772,N_19732,N_18403);
and U21773 (N_21773,N_18155,N_15789);
nor U21774 (N_21774,N_18692,N_19942);
xor U21775 (N_21775,N_19197,N_16392);
and U21776 (N_21776,N_16837,N_16442);
or U21777 (N_21777,N_16785,N_17456);
and U21778 (N_21778,N_16889,N_19630);
and U21779 (N_21779,N_19598,N_19381);
or U21780 (N_21780,N_15211,N_15549);
nor U21781 (N_21781,N_19658,N_18566);
nor U21782 (N_21782,N_17524,N_16942);
or U21783 (N_21783,N_17611,N_18510);
xor U21784 (N_21784,N_16909,N_16907);
xor U21785 (N_21785,N_16393,N_15130);
xnor U21786 (N_21786,N_19948,N_17157);
nand U21787 (N_21787,N_16433,N_18420);
or U21788 (N_21788,N_16860,N_19594);
and U21789 (N_21789,N_15980,N_16897);
xnor U21790 (N_21790,N_16017,N_15167);
or U21791 (N_21791,N_18257,N_18025);
and U21792 (N_21792,N_16481,N_19039);
or U21793 (N_21793,N_19797,N_19673);
and U21794 (N_21794,N_16252,N_18925);
or U21795 (N_21795,N_16693,N_18629);
nand U21796 (N_21796,N_16775,N_17991);
and U21797 (N_21797,N_18503,N_18588);
nor U21798 (N_21798,N_16586,N_18224);
and U21799 (N_21799,N_19192,N_18158);
and U21800 (N_21800,N_17803,N_18821);
or U21801 (N_21801,N_15307,N_16417);
xnor U21802 (N_21802,N_16601,N_17900);
or U21803 (N_21803,N_19146,N_15276);
or U21804 (N_21804,N_19655,N_17689);
nor U21805 (N_21805,N_15638,N_18918);
nand U21806 (N_21806,N_18443,N_17721);
or U21807 (N_21807,N_15141,N_16633);
and U21808 (N_21808,N_15370,N_16783);
xor U21809 (N_21809,N_18798,N_15129);
and U21810 (N_21810,N_18693,N_16718);
or U21811 (N_21811,N_17430,N_18591);
or U21812 (N_21812,N_16459,N_16638);
nor U21813 (N_21813,N_15827,N_15825);
nor U21814 (N_21814,N_17835,N_18022);
nor U21815 (N_21815,N_19269,N_17440);
or U21816 (N_21816,N_18240,N_16557);
nand U21817 (N_21817,N_18387,N_18104);
nand U21818 (N_21818,N_17257,N_16999);
and U21819 (N_21819,N_19158,N_17969);
nor U21820 (N_21820,N_15886,N_15550);
or U21821 (N_21821,N_15460,N_15566);
xnor U21822 (N_21822,N_15063,N_19204);
and U21823 (N_21823,N_15085,N_16640);
xor U21824 (N_21824,N_18968,N_15963);
and U21825 (N_21825,N_17766,N_15268);
nor U21826 (N_21826,N_17119,N_15726);
or U21827 (N_21827,N_18134,N_15470);
and U21828 (N_21828,N_16227,N_15150);
and U21829 (N_21829,N_16159,N_16904);
xnor U21830 (N_21830,N_15596,N_17878);
nand U21831 (N_21831,N_17872,N_16049);
or U21832 (N_21832,N_19553,N_18710);
nor U21833 (N_21833,N_16620,N_18486);
nor U21834 (N_21834,N_18215,N_17560);
and U21835 (N_21835,N_16502,N_15823);
and U21836 (N_21836,N_15584,N_16747);
nand U21837 (N_21837,N_15607,N_19642);
and U21838 (N_21838,N_17684,N_19951);
or U21839 (N_21839,N_17249,N_16892);
and U21840 (N_21840,N_15765,N_19429);
and U21841 (N_21841,N_16576,N_15926);
or U21842 (N_21842,N_17028,N_19464);
xor U21843 (N_21843,N_18295,N_16419);
xnor U21844 (N_21844,N_18311,N_15713);
or U21845 (N_21845,N_17583,N_16014);
and U21846 (N_21846,N_16112,N_17758);
or U21847 (N_21847,N_18014,N_17458);
and U21848 (N_21848,N_19603,N_16171);
xnor U21849 (N_21849,N_17637,N_19323);
or U21850 (N_21850,N_18530,N_15065);
or U21851 (N_21851,N_15397,N_18928);
and U21852 (N_21852,N_18349,N_18880);
xnor U21853 (N_21853,N_17633,N_18626);
and U21854 (N_21854,N_16498,N_16921);
nor U21855 (N_21855,N_16704,N_17750);
nor U21856 (N_21856,N_17307,N_19120);
nand U21857 (N_21857,N_16399,N_16508);
nor U21858 (N_21858,N_18674,N_18143);
nor U21859 (N_21859,N_15721,N_18742);
or U21860 (N_21860,N_16337,N_16047);
or U21861 (N_21861,N_16754,N_18484);
nor U21862 (N_21862,N_17714,N_17649);
nand U21863 (N_21863,N_16957,N_16962);
and U21864 (N_21864,N_18592,N_16792);
and U21865 (N_21865,N_15516,N_19060);
xnor U21866 (N_21866,N_17893,N_19257);
nor U21867 (N_21867,N_16800,N_15728);
nor U21868 (N_21868,N_19654,N_15866);
nor U21869 (N_21869,N_19580,N_19866);
and U21870 (N_21870,N_17734,N_15759);
nand U21871 (N_21871,N_18713,N_18769);
and U21872 (N_21872,N_16976,N_18292);
nor U21873 (N_21873,N_16515,N_15154);
nand U21874 (N_21874,N_15025,N_17563);
or U21875 (N_21875,N_15742,N_18212);
xor U21876 (N_21876,N_15493,N_19443);
xnor U21877 (N_21877,N_17562,N_18456);
nand U21878 (N_21878,N_18089,N_19049);
or U21879 (N_21879,N_16062,N_16675);
xnor U21880 (N_21880,N_19980,N_19997);
xnor U21881 (N_21881,N_18962,N_18883);
nand U21882 (N_21882,N_17970,N_18091);
and U21883 (N_21883,N_18124,N_15826);
or U21884 (N_21884,N_17712,N_16084);
or U21885 (N_21885,N_17988,N_18695);
nand U21886 (N_21886,N_15846,N_18343);
or U21887 (N_21887,N_17208,N_16380);
xor U21888 (N_21888,N_19840,N_15486);
nor U21889 (N_21889,N_19290,N_15253);
or U21890 (N_21890,N_17716,N_18914);
xor U21891 (N_21891,N_17299,N_16513);
xor U21892 (N_21892,N_19533,N_16485);
nor U21893 (N_21893,N_18897,N_17746);
and U21894 (N_21894,N_18272,N_18313);
nand U21895 (N_21895,N_17404,N_18768);
and U21896 (N_21896,N_17234,N_17627);
nor U21897 (N_21897,N_17512,N_18524);
nand U21898 (N_21898,N_17460,N_19674);
or U21899 (N_21899,N_19628,N_16163);
or U21900 (N_21900,N_15565,N_18253);
or U21901 (N_21901,N_17860,N_15279);
nor U21902 (N_21902,N_15898,N_18571);
nor U21903 (N_21903,N_17584,N_17850);
nor U21904 (N_21904,N_19355,N_18362);
nor U21905 (N_21905,N_17146,N_19450);
nand U21906 (N_21906,N_17519,N_18286);
or U21907 (N_21907,N_16150,N_16542);
nand U21908 (N_21908,N_19009,N_18641);
xnor U21909 (N_21909,N_18324,N_17480);
nor U21910 (N_21910,N_18136,N_19371);
xor U21911 (N_21911,N_17435,N_16411);
and U21912 (N_21912,N_15465,N_15608);
xor U21913 (N_21913,N_18100,N_19272);
and U21914 (N_21914,N_17246,N_15285);
nor U21915 (N_21915,N_15055,N_19873);
and U21916 (N_21916,N_15296,N_19634);
nand U21917 (N_21917,N_18045,N_15533);
xor U21918 (N_21918,N_17400,N_16692);
and U21919 (N_21919,N_16383,N_15332);
and U21920 (N_21920,N_18032,N_18135);
xnor U21921 (N_21921,N_16721,N_18300);
or U21922 (N_21922,N_17351,N_19326);
or U21923 (N_21923,N_19441,N_18145);
nand U21924 (N_21924,N_17201,N_19544);
or U21925 (N_21925,N_17520,N_16711);
or U21926 (N_21926,N_15850,N_17255);
xnor U21927 (N_21927,N_15854,N_19782);
xnor U21928 (N_21928,N_15247,N_17009);
nand U21929 (N_21929,N_17904,N_15108);
and U21930 (N_21930,N_16857,N_15734);
nand U21931 (N_21931,N_17008,N_16107);
xnor U21932 (N_21932,N_17736,N_19128);
or U21933 (N_21933,N_15219,N_18259);
and U21934 (N_21934,N_17931,N_19156);
and U21935 (N_21935,N_18140,N_18578);
xnor U21936 (N_21936,N_17847,N_18478);
nor U21937 (N_21937,N_19511,N_17722);
or U21938 (N_21938,N_16891,N_15216);
nor U21939 (N_21939,N_16968,N_18791);
nand U21940 (N_21940,N_16830,N_15689);
and U21941 (N_21941,N_19519,N_17270);
or U21942 (N_21942,N_18895,N_17412);
nand U21943 (N_21943,N_15111,N_17998);
xor U21944 (N_21944,N_19915,N_15794);
xor U21945 (N_21945,N_19559,N_16245);
nand U21946 (N_21946,N_19077,N_17319);
nand U21947 (N_21947,N_18127,N_15620);
nand U21948 (N_21948,N_16790,N_17141);
xor U21949 (N_21949,N_15308,N_18994);
nand U21950 (N_21950,N_19485,N_17676);
nor U21951 (N_21951,N_17713,N_17992);
nand U21952 (N_21952,N_19730,N_15649);
nor U21953 (N_21953,N_18186,N_19994);
nand U21954 (N_21954,N_15915,N_19587);
xnor U21955 (N_21955,N_18888,N_17765);
and U21956 (N_21956,N_18269,N_17016);
nand U21957 (N_21957,N_18131,N_15652);
and U21958 (N_21958,N_19725,N_16723);
and U21959 (N_21959,N_17022,N_19109);
and U21960 (N_21960,N_15452,N_19759);
nor U21961 (N_21961,N_18033,N_19785);
and U21962 (N_21962,N_17342,N_19850);
nor U21963 (N_21963,N_16234,N_17628);
xor U21964 (N_21964,N_17927,N_18846);
nand U21965 (N_21965,N_16040,N_19616);
xor U21966 (N_21966,N_16585,N_16810);
or U21967 (N_21967,N_15374,N_15639);
and U21968 (N_21968,N_15210,N_16404);
and U21969 (N_21969,N_19385,N_17784);
nand U21970 (N_21970,N_17109,N_18026);
nor U21971 (N_21971,N_18727,N_16128);
nand U21972 (N_21972,N_18096,N_16762);
nor U21973 (N_21973,N_15026,N_18149);
nor U21974 (N_21974,N_19902,N_18156);
and U21975 (N_21975,N_19618,N_15984);
xor U21976 (N_21976,N_17974,N_17924);
or U21977 (N_21977,N_15142,N_17749);
and U21978 (N_21978,N_16541,N_17579);
or U21979 (N_21979,N_15030,N_18445);
or U21980 (N_21980,N_17359,N_16960);
and U21981 (N_21981,N_19328,N_19016);
or U21982 (N_21982,N_17032,N_16950);
and U21983 (N_21983,N_18148,N_19160);
nand U21984 (N_21984,N_16523,N_15530);
nand U21985 (N_21985,N_19339,N_17610);
nand U21986 (N_21986,N_19438,N_19934);
or U21987 (N_21987,N_16265,N_18777);
or U21988 (N_21988,N_15089,N_15182);
nor U21989 (N_21989,N_19676,N_16123);
nor U21990 (N_21990,N_15536,N_18568);
or U21991 (N_21991,N_16151,N_16984);
or U21992 (N_21992,N_18642,N_15885);
xnor U21993 (N_21993,N_17263,N_18704);
xor U21994 (N_21994,N_15169,N_17425);
xor U21995 (N_21995,N_16978,N_17546);
or U21996 (N_21996,N_17521,N_16472);
or U21997 (N_21997,N_17881,N_17099);
or U21998 (N_21998,N_18732,N_19359);
nand U21999 (N_21999,N_18995,N_17450);
xor U22000 (N_22000,N_17411,N_16471);
nand U22001 (N_22001,N_17012,N_16426);
nor U22002 (N_22002,N_18516,N_15949);
or U22003 (N_22003,N_17692,N_17069);
or U22004 (N_22004,N_17055,N_15348);
nand U22005 (N_22005,N_15883,N_15288);
and U22006 (N_22006,N_15684,N_16283);
nand U22007 (N_22007,N_15233,N_16181);
nor U22008 (N_22008,N_19560,N_15208);
or U22009 (N_22009,N_19045,N_19878);
nor U22010 (N_22010,N_19324,N_18309);
and U22011 (N_22011,N_19963,N_17279);
nor U22012 (N_22012,N_15301,N_17265);
and U22013 (N_22013,N_18405,N_16672);
and U22014 (N_22014,N_19792,N_19500);
nand U22015 (N_22015,N_16094,N_19334);
and U22016 (N_22016,N_15133,N_17829);
or U22017 (N_22017,N_19276,N_15773);
xor U22018 (N_22018,N_19059,N_16048);
or U22019 (N_22019,N_16610,N_19119);
and U22020 (N_22020,N_15136,N_18972);
or U22021 (N_22021,N_18899,N_19849);
and U22022 (N_22022,N_17836,N_19094);
nor U22023 (N_22023,N_19147,N_19249);
nor U22024 (N_22024,N_15237,N_18373);
xor U22025 (N_22025,N_15385,N_17531);
or U22026 (N_22026,N_17114,N_15856);
nand U22027 (N_22027,N_19901,N_17077);
and U22028 (N_22028,N_17096,N_16710);
xnor U22029 (N_22029,N_17498,N_19356);
or U22030 (N_22030,N_17834,N_17298);
nand U22031 (N_22031,N_15437,N_15049);
and U22032 (N_22032,N_16012,N_18553);
and U22033 (N_22033,N_19586,N_18943);
nor U22034 (N_22034,N_19786,N_19900);
xor U22035 (N_22035,N_16969,N_18243);
nand U22036 (N_22036,N_15015,N_16614);
nor U22037 (N_22037,N_16493,N_16736);
and U22038 (N_22038,N_15957,N_16533);
nand U22039 (N_22039,N_18239,N_16623);
xor U22040 (N_22040,N_18986,N_17930);
nor U22041 (N_22041,N_17515,N_15172);
or U22042 (N_22042,N_15904,N_15573);
nand U22043 (N_22043,N_15495,N_17092);
or U22044 (N_22044,N_18810,N_18514);
and U22045 (N_22045,N_15795,N_19777);
nor U22046 (N_22046,N_17304,N_19471);
nand U22047 (N_22047,N_17436,N_15528);
xor U22048 (N_22048,N_18027,N_17409);
or U22049 (N_22049,N_15479,N_16898);
nor U22050 (N_22050,N_16093,N_19067);
xnor U22051 (N_22051,N_17638,N_18234);
nand U22052 (N_22052,N_17431,N_15849);
nor U22053 (N_22053,N_15275,N_15582);
and U22054 (N_22054,N_19465,N_17402);
or U22055 (N_22055,N_17826,N_16243);
or U22056 (N_22056,N_18976,N_19605);
xor U22057 (N_22057,N_16598,N_15828);
nand U22058 (N_22058,N_16600,N_19342);
xor U22059 (N_22059,N_19085,N_16239);
or U22060 (N_22060,N_18345,N_19404);
xor U22061 (N_22061,N_17585,N_15444);
nand U22062 (N_22062,N_18564,N_18772);
and U22063 (N_22063,N_19182,N_17620);
nand U22064 (N_22064,N_17178,N_17207);
or U22065 (N_22065,N_15766,N_17745);
or U22066 (N_22066,N_17368,N_16343);
or U22067 (N_22067,N_19751,N_19727);
nand U22068 (N_22068,N_15446,N_19892);
nor U22069 (N_22069,N_15855,N_16368);
xor U22070 (N_22070,N_18223,N_19813);
or U22071 (N_22071,N_17950,N_17972);
xnor U22072 (N_22072,N_15764,N_18412);
xnor U22073 (N_22073,N_18518,N_15410);
xnor U22074 (N_22074,N_19073,N_18214);
nor U22075 (N_22075,N_15860,N_19021);
xnor U22076 (N_22076,N_19724,N_18123);
or U22077 (N_22077,N_19789,N_16186);
nand U22078 (N_22078,N_15891,N_19383);
nand U22079 (N_22079,N_17139,N_18073);
and U22080 (N_22080,N_16983,N_16416);
nor U22081 (N_22081,N_18348,N_19217);
nor U22082 (N_22082,N_15184,N_16447);
and U22083 (N_22083,N_19105,N_15508);
and U22084 (N_22084,N_19308,N_16963);
or U22085 (N_22085,N_18463,N_17513);
xor U22086 (N_22086,N_15107,N_19805);
nand U22087 (N_22087,N_19697,N_17561);
and U22088 (N_22088,N_17275,N_18050);
nand U22089 (N_22089,N_16439,N_15919);
nor U22090 (N_22090,N_16756,N_19400);
xor U22091 (N_22091,N_18740,N_19842);
nor U22092 (N_22092,N_19168,N_17551);
nor U22093 (N_22093,N_17116,N_16214);
or U22094 (N_22094,N_17206,N_18365);
and U22095 (N_22095,N_16908,N_18624);
and U22096 (N_22096,N_19431,N_19098);
and U22097 (N_22097,N_16679,N_18745);
xor U22098 (N_22098,N_18502,N_15542);
or U22099 (N_22099,N_19079,N_15853);
and U22100 (N_22100,N_15986,N_19492);
nor U22101 (N_22101,N_15527,N_15506);
and U22102 (N_22102,N_19650,N_19534);
nor U22103 (N_22103,N_18924,N_17127);
and U22104 (N_22104,N_15041,N_18956);
nor U22105 (N_22105,N_18937,N_16080);
and U22106 (N_22106,N_16641,N_15036);
xor U22107 (N_22107,N_17928,N_18643);
xor U22108 (N_22108,N_19776,N_18333);
and U22109 (N_22109,N_19432,N_16113);
nor U22110 (N_22110,N_19558,N_19103);
nand U22111 (N_22111,N_15077,N_18379);
xnor U22112 (N_22112,N_15518,N_19696);
xor U22113 (N_22113,N_15692,N_18820);
and U22114 (N_22114,N_17670,N_17070);
nor U22115 (N_22115,N_15706,N_18421);
nor U22116 (N_22116,N_17648,N_16685);
or U22117 (N_22117,N_15534,N_15483);
xor U22118 (N_22118,N_16606,N_15369);
and U22119 (N_22119,N_18708,N_17452);
or U22120 (N_22120,N_15271,N_19213);
or U22121 (N_22121,N_15207,N_15500);
nor U22122 (N_22122,N_18671,N_15179);
or U22123 (N_22123,N_19489,N_18765);
nand U22124 (N_22124,N_15175,N_16980);
and U22125 (N_22125,N_15832,N_18318);
and U22126 (N_22126,N_16678,N_18159);
or U22127 (N_22127,N_15979,N_18411);
nand U22128 (N_22128,N_16189,N_16683);
and U22129 (N_22129,N_16278,N_18827);
nand U22130 (N_22130,N_17660,N_17507);
or U22131 (N_22131,N_16224,N_18556);
and U22132 (N_22132,N_15874,N_15994);
and U22133 (N_22133,N_16647,N_15673);
xnor U22134 (N_22134,N_15241,N_18372);
nand U22135 (N_22135,N_17735,N_15851);
nor U22136 (N_22136,N_15286,N_18594);
xnor U22137 (N_22137,N_17688,N_18581);
and U22138 (N_22138,N_19745,N_15409);
and U22139 (N_22139,N_17917,N_16100);
or U22140 (N_22140,N_17797,N_15723);
nor U22141 (N_22141,N_16841,N_17216);
xor U22142 (N_22142,N_18634,N_17996);
or U22143 (N_22143,N_17165,N_17158);
or U22144 (N_22144,N_16288,N_15658);
xor U22145 (N_22145,N_19268,N_15977);
nand U22146 (N_22146,N_18537,N_15784);
and U22147 (N_22147,N_15404,N_16733);
or U22148 (N_22148,N_17839,N_19579);
xor U22149 (N_22149,N_19921,N_18428);
and U22150 (N_22150,N_15600,N_15418);
or U22151 (N_22151,N_17858,N_15164);
xor U22152 (N_22152,N_18178,N_19972);
nand U22153 (N_22153,N_19720,N_18122);
or U22154 (N_22154,N_15646,N_17502);
nand U22155 (N_22155,N_19555,N_15012);
xor U22156 (N_22156,N_18752,N_17943);
nor U22157 (N_22157,N_18230,N_15936);
xor U22158 (N_22158,N_16655,N_17958);
or U22159 (N_22159,N_19771,N_15430);
xor U22160 (N_22160,N_17912,N_18432);
or U22161 (N_22161,N_18844,N_15595);
or U22162 (N_22162,N_18523,N_18886);
nand U22163 (N_22163,N_18685,N_19136);
xnor U22164 (N_22164,N_18023,N_16295);
and U22165 (N_22165,N_18342,N_15525);
and U22166 (N_22166,N_19946,N_15606);
and U22167 (N_22167,N_17885,N_17614);
nand U22168 (N_22168,N_17283,N_15244);
nor U22169 (N_22169,N_17642,N_19713);
nand U22170 (N_22170,N_18617,N_19163);
or U22171 (N_22171,N_15817,N_16242);
and U22172 (N_22172,N_19591,N_18970);
and U22173 (N_22173,N_19106,N_15340);
nand U22174 (N_22174,N_17403,N_16370);
and U22175 (N_22175,N_18221,N_15757);
xor U22176 (N_22176,N_17302,N_18945);
nand U22177 (N_22177,N_19488,N_19498);
nand U22178 (N_22178,N_19691,N_15005);
xor U22179 (N_22179,N_18133,N_17806);
or U22180 (N_22180,N_15197,N_17205);
nor U22181 (N_22181,N_17656,N_18815);
nor U22182 (N_22182,N_17327,N_16072);
and U22183 (N_22183,N_18299,N_19428);
and U22184 (N_22184,N_19286,N_19760);
and U22185 (N_22185,N_18176,N_15729);
nor U22186 (N_22186,N_15791,N_17088);
or U22187 (N_22187,N_18208,N_15781);
and U22188 (N_22188,N_15035,N_19595);
or U22189 (N_22189,N_16829,N_18444);
and U22190 (N_22190,N_15481,N_15008);
or U22191 (N_22191,N_17017,N_19877);
nand U22192 (N_22192,N_17000,N_16354);
or U22193 (N_22193,N_15869,N_18138);
or U22194 (N_22194,N_19670,N_18904);
and U22195 (N_22195,N_16201,N_15048);
nor U22196 (N_22196,N_19854,N_17376);
nor U22197 (N_22197,N_16768,N_15346);
nand U22198 (N_22198,N_15173,N_15333);
nor U22199 (N_22199,N_16520,N_17423);
or U22200 (N_22200,N_17908,N_16934);
nor U22201 (N_22201,N_17312,N_19346);
nand U22202 (N_22202,N_15070,N_17916);
nand U22203 (N_22203,N_16377,N_19514);
xnor U22204 (N_22204,N_19992,N_15408);
nor U22205 (N_22205,N_16290,N_17600);
nand U22206 (N_22206,N_18718,N_16463);
xor U22207 (N_22207,N_19430,N_18385);
or U22208 (N_22208,N_19723,N_17731);
nand U22209 (N_22209,N_16948,N_19179);
nor U22210 (N_22210,N_19220,N_18455);
xor U22211 (N_22211,N_15775,N_18071);
or U22212 (N_22212,N_19606,N_17586);
or U22213 (N_22213,N_16223,N_15080);
and U22214 (N_22214,N_17183,N_18340);
xnor U22215 (N_22215,N_18439,N_15091);
and U22216 (N_22216,N_18454,N_18354);
or U22217 (N_22217,N_17619,N_19566);
or U22218 (N_22218,N_17013,N_18522);
xor U22219 (N_22219,N_17623,N_19071);
nor U22220 (N_22220,N_18528,N_17499);
and U22221 (N_22221,N_19306,N_15837);
and U22222 (N_22222,N_19516,N_16438);
and U22223 (N_22223,N_16544,N_19715);
and U22224 (N_22224,N_17064,N_16254);
xnor U22225 (N_22225,N_19808,N_16069);
nor U22226 (N_22226,N_15137,N_17241);
nor U22227 (N_22227,N_17330,N_18735);
xor U22228 (N_22228,N_16313,N_16454);
nor U22229 (N_22229,N_17556,N_19375);
nor U22230 (N_22230,N_15270,N_17679);
or U22231 (N_22231,N_19363,N_18499);
xnor U22232 (N_22232,N_16448,N_16932);
xor U22233 (N_22233,N_15382,N_18864);
and U22234 (N_22234,N_17673,N_19896);
and U22235 (N_22235,N_17762,N_16293);
nor U22236 (N_22236,N_17490,N_17447);
and U22237 (N_22237,N_17196,N_15688);
nand U22238 (N_22238,N_16147,N_18816);
or U22239 (N_22239,N_17223,N_17966);
and U22240 (N_22240,N_15631,N_18763);
and U22241 (N_22241,N_17831,N_17204);
nor U22242 (N_22242,N_17471,N_19074);
nor U22243 (N_22243,N_18044,N_17870);
nand U22244 (N_22244,N_15093,N_15560);
and U22245 (N_22245,N_16292,N_15873);
and U22246 (N_22246,N_16053,N_15859);
nor U22247 (N_22247,N_16666,N_15229);
nand U22248 (N_22248,N_15324,N_17062);
and U22249 (N_22249,N_18029,N_17230);
nand U22250 (N_22250,N_16564,N_17317);
and U22251 (N_22251,N_19583,N_17023);
nor U22252 (N_22252,N_16407,N_15082);
nor U22253 (N_22253,N_15987,N_19294);
nand U22254 (N_22254,N_18596,N_18308);
or U22255 (N_22255,N_18175,N_17049);
or U22256 (N_22256,N_18390,N_18005);
nand U22257 (N_22257,N_16545,N_15445);
or U22258 (N_22258,N_17108,N_16009);
or U22259 (N_22259,N_19899,N_15635);
or U22260 (N_22260,N_18197,N_19883);
or U22261 (N_22261,N_17406,N_19506);
nand U22262 (N_22262,N_18162,N_17799);
nor U22263 (N_22263,N_16716,N_17650);
xnor U22264 (N_22264,N_18878,N_19665);
nor U22265 (N_22265,N_16314,N_19719);
or U22266 (N_22266,N_16275,N_18270);
and U22267 (N_22267,N_18790,N_17844);
nor U22268 (N_22268,N_19496,N_15788);
xnor U22269 (N_22269,N_15907,N_18219);
nor U22270 (N_22270,N_15838,N_18680);
nand U22271 (N_22271,N_19546,N_15423);
or U22272 (N_22272,N_17338,N_19596);
nand U22273 (N_22273,N_16763,N_16105);
nor U22274 (N_22274,N_18619,N_15146);
or U22275 (N_22275,N_15189,N_19171);
xnor U22276 (N_22276,N_17346,N_15391);
and U22277 (N_22277,N_18182,N_15061);
and U22278 (N_22278,N_18789,N_18137);
and U22279 (N_22279,N_19608,N_15235);
nand U22280 (N_22280,N_15967,N_19852);
nand U22281 (N_22281,N_19822,N_15909);
and U22282 (N_22282,N_15633,N_15386);
xnor U22283 (N_22283,N_18493,N_19222);
nor U22284 (N_22284,N_19057,N_16674);
xnor U22285 (N_22285,N_17380,N_17085);
nor U22286 (N_22286,N_17810,N_15152);
and U22287 (N_22287,N_17790,N_15269);
nor U22288 (N_22288,N_19135,N_15750);
xor U22289 (N_22289,N_16282,N_18368);
nand U22290 (N_22290,N_15616,N_16814);
nor U22291 (N_22291,N_18981,N_15670);
and U22292 (N_22292,N_15143,N_15546);
xor U22293 (N_22293,N_17723,N_17538);
nor U22294 (N_22294,N_16560,N_17823);
and U22295 (N_22295,N_15407,N_15181);
and U22296 (N_22296,N_19889,N_17629);
or U22297 (N_22297,N_16019,N_17509);
nand U22298 (N_22298,N_15588,N_19803);
or U22299 (N_22299,N_15563,N_17060);
nor U22300 (N_22300,N_18235,N_17094);
nor U22301 (N_22301,N_18277,N_16712);
nand U22302 (N_22302,N_19444,N_18722);
xor U22303 (N_22303,N_17525,N_15463);
and U22304 (N_22304,N_17466,N_15454);
and U22305 (N_22305,N_15261,N_16487);
nand U22306 (N_22306,N_16261,N_18608);
or U22307 (N_22307,N_15076,N_16534);
nor U22308 (N_22308,N_18028,N_15720);
and U22309 (N_22309,N_19233,N_17335);
xor U22310 (N_22310,N_19741,N_15958);
nand U22311 (N_22311,N_18233,N_19640);
nor U22312 (N_22312,N_18609,N_15718);
nand U22313 (N_22313,N_18730,N_18845);
nor U22314 (N_22314,N_18103,N_17372);
nand U22315 (N_22315,N_18193,N_18380);
and U22316 (N_22316,N_15017,N_19648);
and U22317 (N_22317,N_16731,N_16618);
and U22318 (N_22318,N_15099,N_18462);
or U22319 (N_22319,N_15467,N_18109);
nand U22320 (N_22320,N_15292,N_17559);
nor U22321 (N_22321,N_17905,N_18645);
xnor U22322 (N_22322,N_18818,N_15682);
and U22323 (N_22323,N_18667,N_17227);
or U22324 (N_22324,N_15326,N_16450);
xor U22325 (N_22325,N_19812,N_18015);
nand U22326 (N_22326,N_15079,N_19095);
xnor U22327 (N_22327,N_17853,N_17677);
xnor U22328 (N_22328,N_15312,N_15908);
xor U22329 (N_22329,N_18835,N_18633);
nor U22330 (N_22330,N_17121,N_18963);
or U22331 (N_22331,N_15746,N_17849);
nand U22332 (N_22332,N_15447,N_15881);
xor U22333 (N_22333,N_19716,N_18307);
and U22334 (N_22334,N_19941,N_19239);
or U22335 (N_22335,N_17635,N_17281);
nand U22336 (N_22336,N_19704,N_16828);
and U22337 (N_22337,N_15453,N_16772);
xnor U22338 (N_22338,N_15735,N_16218);
xnor U22339 (N_22339,N_15872,N_16488);
nor U22340 (N_22340,N_18832,N_17086);
and U22341 (N_22341,N_16141,N_19898);
nor U22342 (N_22342,N_17029,N_16517);
and U22343 (N_22343,N_18811,N_15780);
and U22344 (N_22344,N_18875,N_15157);
xnor U22345 (N_22345,N_15032,N_16864);
xor U22346 (N_22346,N_19251,N_16696);
nand U22347 (N_22347,N_16324,N_17911);
or U22348 (N_22348,N_19947,N_16166);
nand U22349 (N_22349,N_19929,N_18417);
or U22350 (N_22350,N_18851,N_15615);
nor U22351 (N_22351,N_18097,N_18559);
nor U22352 (N_22352,N_18388,N_18289);
nand U22353 (N_22353,N_16089,N_18172);
or U22354 (N_22354,N_16882,N_17634);
or U22355 (N_22355,N_16835,N_18890);
xor U22356 (N_22356,N_15709,N_15126);
or U22357 (N_22357,N_15526,N_17087);
nand U22358 (N_22358,N_19927,N_17280);
xnor U22359 (N_22359,N_19206,N_19969);
and U22360 (N_22360,N_17036,N_19537);
or U22361 (N_22361,N_18018,N_16796);
or U22362 (N_22362,N_15395,N_16888);
nor U22363 (N_22363,N_16507,N_15377);
nor U22364 (N_22364,N_15725,N_19904);
or U22365 (N_22365,N_17573,N_17396);
nor U22366 (N_22366,N_15938,N_15544);
xor U22367 (N_22367,N_16326,N_15281);
nand U22368 (N_22368,N_18306,N_18297);
xnor U22369 (N_22369,N_15894,N_19421);
nor U22370 (N_22370,N_16351,N_18314);
nand U22371 (N_22371,N_15105,N_18613);
nor U22372 (N_22372,N_17100,N_16046);
or U22373 (N_22373,N_16914,N_19801);
and U22374 (N_22374,N_18837,N_19118);
xor U22375 (N_22375,N_18927,N_18817);
and U22376 (N_22376,N_17700,N_19872);
xnor U22377 (N_22377,N_19002,N_19030);
xor U22378 (N_22378,N_17355,N_19729);
xor U22379 (N_22379,N_16495,N_16267);
xnor U22380 (N_22380,N_15263,N_15058);
and U22381 (N_22381,N_15824,N_17955);
xnor U22382 (N_22382,N_18460,N_18392);
and U22383 (N_22383,N_17407,N_15769);
or U22384 (N_22384,N_19155,N_15496);
nor U22385 (N_22385,N_19499,N_15489);
and U22386 (N_22386,N_16308,N_15132);
nand U22387 (N_22387,N_18664,N_17284);
or U22388 (N_22388,N_18507,N_18687);
and U22389 (N_22389,N_19909,N_18830);
nand U22390 (N_22390,N_17083,N_16116);
and U22391 (N_22391,N_15188,N_17511);
nand U22392 (N_22392,N_17329,N_18582);
xnor U22393 (N_22393,N_16233,N_16844);
xor U22394 (N_22394,N_19547,N_15412);
xnor U22395 (N_22395,N_19625,N_16540);
and U22396 (N_22396,N_18079,N_17328);
or U22397 (N_22397,N_19753,N_16118);
nand U22398 (N_22398,N_19117,N_15999);
xnor U22399 (N_22399,N_19162,N_17960);
and U22400 (N_22400,N_18561,N_17350);
nand U22401 (N_22401,N_19010,N_19632);
xnor U22402 (N_22402,N_15972,N_15521);
or U22403 (N_22403,N_15617,N_16918);
xnor U22404 (N_22404,N_19475,N_19486);
nor U22405 (N_22405,N_18625,N_19851);
or U22406 (N_22406,N_17683,N_19530);
xor U22407 (N_22407,N_15793,N_16099);
nand U22408 (N_22408,N_19116,N_18901);
and U22409 (N_22409,N_15122,N_18371);
nand U22410 (N_22410,N_16973,N_16032);
nor U22411 (N_22411,N_19202,N_15473);
or U22412 (N_22412,N_16848,N_15398);
and U22413 (N_22413,N_18458,N_16745);
nor U22414 (N_22414,N_17420,N_15186);
or U22415 (N_22415,N_15212,N_15580);
xor U22416 (N_22416,N_18068,N_19681);
nor U22417 (N_22417,N_16071,N_18698);
or U22418 (N_22418,N_17884,N_18660);
and U22419 (N_22419,N_16449,N_18860);
or U22420 (N_22420,N_16139,N_18593);
xnor U22421 (N_22421,N_18361,N_17030);
nand U22422 (N_22422,N_16535,N_16277);
and U22423 (N_22423,N_16409,N_15840);
nand U22424 (N_22424,N_17065,N_19863);
or U22425 (N_22425,N_19680,N_17842);
or U22426 (N_22426,N_17377,N_19974);
or U22427 (N_22427,N_18731,N_19979);
or U22428 (N_22428,N_19858,N_17978);
nand U22429 (N_22429,N_19102,N_18936);
xor U22430 (N_22430,N_18691,N_18672);
xor U22431 (N_22431,N_19301,N_17232);
xnor U22432 (N_22432,N_18610,N_19329);
and U22433 (N_22433,N_19728,N_15911);
nor U22434 (N_22434,N_17813,N_15417);
or U22435 (N_22435,N_16874,N_18332);
and U22436 (N_22436,N_18784,N_19535);
and U22437 (N_22437,N_16519,N_17463);
nor U22438 (N_22438,N_18494,N_19599);
xnor U22439 (N_22439,N_16034,N_16729);
or U22440 (N_22440,N_16832,N_15778);
nand U22441 (N_22441,N_17325,N_19047);
and U22442 (N_22442,N_15220,N_19978);
nand U22443 (N_22443,N_17769,N_15118);
or U22444 (N_22444,N_18975,N_19722);
or U22445 (N_22445,N_19740,N_18627);
nor U22446 (N_22446,N_19844,N_17741);
or U22447 (N_22447,N_15792,N_19467);
nor U22448 (N_22448,N_19774,N_16251);
nand U22449 (N_22449,N_19262,N_16913);
or U22450 (N_22450,N_19561,N_15752);
xor U22451 (N_22451,N_16746,N_19726);
nand U22452 (N_22452,N_16395,N_15998);
nand U22453 (N_22453,N_18785,N_18871);
nand U22454 (N_22454,N_18353,N_17110);
and U22455 (N_22455,N_19845,N_16311);
and U22456 (N_22456,N_18665,N_18320);
nor U22457 (N_22457,N_17536,N_19988);
and U22458 (N_22458,N_18599,N_19279);
and U22459 (N_22459,N_18298,N_15482);
or U22460 (N_22460,N_18738,N_19297);
nand U22461 (N_22461,N_19461,N_18536);
nand U22462 (N_22462,N_15095,N_18606);
nand U22463 (N_22463,N_16807,N_15806);
and U22464 (N_22464,N_18250,N_17657);
xnor U22465 (N_22465,N_18628,N_19700);
or U22466 (N_22466,N_16812,N_17658);
and U22467 (N_22467,N_15073,N_19970);
nand U22468 (N_22468,N_18377,N_19224);
nand U22469 (N_22469,N_16065,N_16106);
or U22470 (N_22470,N_17047,N_16024);
nor U22471 (N_22471,N_16744,N_18437);
nand U22472 (N_22472,N_16030,N_15581);
nand U22473 (N_22473,N_16548,N_15282);
nand U22474 (N_22474,N_19296,N_17962);
or U22475 (N_22475,N_15645,N_19911);
nor U22476 (N_22476,N_18957,N_17888);
nand U22477 (N_22477,N_15812,N_16440);
xnor U22478 (N_22478,N_17967,N_18378);
nand U22479 (N_22479,N_17622,N_17084);
xor U22480 (N_22480,N_18892,N_15636);
xnor U22481 (N_22481,N_17153,N_16998);
or U22482 (N_22482,N_15401,N_19133);
and U22483 (N_22483,N_19104,N_17439);
nand U22484 (N_22484,N_17170,N_16895);
or U22485 (N_22485,N_18477,N_16157);
and U22486 (N_22486,N_16720,N_18251);
and U22487 (N_22487,N_18093,N_18051);
nand U22488 (N_22488,N_16668,N_18119);
xnor U22489 (N_22489,N_16527,N_16244);
nor U22490 (N_22490,N_15381,N_16415);
and U22491 (N_22491,N_18010,N_18733);
nor U22492 (N_22492,N_19875,N_15707);
nand U22493 (N_22493,N_19790,N_16031);
xor U22494 (N_22494,N_19052,N_18696);
and U22495 (N_22495,N_18064,N_17332);
or U22496 (N_22496,N_17179,N_15738);
and U22497 (N_22497,N_17134,N_15739);
nand U22498 (N_22498,N_19277,N_15139);
xor U22499 (N_22499,N_15554,N_18736);
xor U22500 (N_22500,N_17416,N_19037);
and U22501 (N_22501,N_18585,N_18974);
and U22502 (N_22502,N_17910,N_18409);
nor U22503 (N_22503,N_15957,N_16441);
nor U22504 (N_22504,N_19055,N_19089);
and U22505 (N_22505,N_17280,N_18508);
xnor U22506 (N_22506,N_19556,N_16089);
nor U22507 (N_22507,N_18267,N_15302);
or U22508 (N_22508,N_17079,N_18927);
and U22509 (N_22509,N_17312,N_19264);
xor U22510 (N_22510,N_19669,N_15503);
and U22511 (N_22511,N_18362,N_18351);
nor U22512 (N_22512,N_16843,N_19478);
and U22513 (N_22513,N_16355,N_18233);
xor U22514 (N_22514,N_19094,N_18527);
and U22515 (N_22515,N_19317,N_15935);
nor U22516 (N_22516,N_18001,N_15039);
nand U22517 (N_22517,N_16402,N_19529);
xor U22518 (N_22518,N_19465,N_17353);
or U22519 (N_22519,N_15851,N_18797);
or U22520 (N_22520,N_18269,N_18552);
xnor U22521 (N_22521,N_18019,N_15371);
nand U22522 (N_22522,N_18321,N_18760);
and U22523 (N_22523,N_19082,N_16997);
or U22524 (N_22524,N_19228,N_15958);
or U22525 (N_22525,N_15804,N_19500);
nor U22526 (N_22526,N_18476,N_15112);
xnor U22527 (N_22527,N_15660,N_16072);
and U22528 (N_22528,N_16880,N_18674);
nor U22529 (N_22529,N_18850,N_15283);
or U22530 (N_22530,N_15204,N_16545);
nor U22531 (N_22531,N_18305,N_17785);
and U22532 (N_22532,N_18126,N_19302);
xnor U22533 (N_22533,N_17855,N_16934);
or U22534 (N_22534,N_16624,N_18478);
xor U22535 (N_22535,N_16836,N_17108);
nand U22536 (N_22536,N_16531,N_17758);
nor U22537 (N_22537,N_19281,N_16670);
or U22538 (N_22538,N_15065,N_15460);
xor U22539 (N_22539,N_16601,N_19734);
or U22540 (N_22540,N_19485,N_17556);
nor U22541 (N_22541,N_18855,N_17598);
xor U22542 (N_22542,N_18089,N_15911);
and U22543 (N_22543,N_18569,N_17620);
and U22544 (N_22544,N_19478,N_16123);
or U22545 (N_22545,N_15990,N_15511);
nor U22546 (N_22546,N_17631,N_16410);
nand U22547 (N_22547,N_16512,N_17128);
xor U22548 (N_22548,N_15864,N_18791);
or U22549 (N_22549,N_19492,N_15395);
and U22550 (N_22550,N_15147,N_19582);
xor U22551 (N_22551,N_16701,N_17310);
and U22552 (N_22552,N_17917,N_15690);
nand U22553 (N_22553,N_19883,N_16268);
and U22554 (N_22554,N_16909,N_15255);
xnor U22555 (N_22555,N_15360,N_15086);
nand U22556 (N_22556,N_15670,N_17343);
xor U22557 (N_22557,N_15181,N_16056);
and U22558 (N_22558,N_19881,N_15040);
xor U22559 (N_22559,N_19826,N_17740);
nor U22560 (N_22560,N_18766,N_19589);
or U22561 (N_22561,N_15486,N_17778);
or U22562 (N_22562,N_15434,N_18747);
nor U22563 (N_22563,N_15173,N_18473);
xor U22564 (N_22564,N_19018,N_17796);
xor U22565 (N_22565,N_16598,N_17414);
nor U22566 (N_22566,N_18553,N_17740);
and U22567 (N_22567,N_15361,N_15497);
nand U22568 (N_22568,N_16301,N_19009);
xnor U22569 (N_22569,N_19449,N_15687);
or U22570 (N_22570,N_16523,N_16949);
or U22571 (N_22571,N_19465,N_18823);
or U22572 (N_22572,N_17651,N_19716);
or U22573 (N_22573,N_17478,N_16420);
xnor U22574 (N_22574,N_19957,N_18903);
nand U22575 (N_22575,N_19730,N_17486);
xnor U22576 (N_22576,N_16766,N_16447);
or U22577 (N_22577,N_19325,N_18296);
xnor U22578 (N_22578,N_16172,N_19123);
or U22579 (N_22579,N_15009,N_19821);
and U22580 (N_22580,N_18369,N_15186);
and U22581 (N_22581,N_17662,N_15774);
or U22582 (N_22582,N_16111,N_16068);
and U22583 (N_22583,N_18596,N_19221);
or U22584 (N_22584,N_16518,N_19533);
or U22585 (N_22585,N_16333,N_18789);
xor U22586 (N_22586,N_17801,N_19233);
or U22587 (N_22587,N_17153,N_17978);
or U22588 (N_22588,N_17760,N_19348);
or U22589 (N_22589,N_19851,N_19773);
xor U22590 (N_22590,N_17658,N_17750);
xnor U22591 (N_22591,N_18980,N_19212);
or U22592 (N_22592,N_15113,N_18248);
nand U22593 (N_22593,N_19785,N_19896);
nor U22594 (N_22594,N_17842,N_15834);
and U22595 (N_22595,N_19283,N_18553);
xor U22596 (N_22596,N_15574,N_18404);
nor U22597 (N_22597,N_17629,N_18241);
nand U22598 (N_22598,N_19846,N_15671);
nand U22599 (N_22599,N_15139,N_17399);
nand U22600 (N_22600,N_18386,N_18080);
nand U22601 (N_22601,N_16805,N_18088);
and U22602 (N_22602,N_15991,N_19642);
and U22603 (N_22603,N_16950,N_19466);
xnor U22604 (N_22604,N_19657,N_19968);
xnor U22605 (N_22605,N_16415,N_18625);
xor U22606 (N_22606,N_16268,N_16928);
nand U22607 (N_22607,N_19206,N_19967);
and U22608 (N_22608,N_16369,N_16221);
and U22609 (N_22609,N_17254,N_16949);
nor U22610 (N_22610,N_16177,N_17603);
and U22611 (N_22611,N_18397,N_19270);
nor U22612 (N_22612,N_18860,N_19757);
nand U22613 (N_22613,N_17588,N_19326);
xnor U22614 (N_22614,N_18839,N_17259);
nor U22615 (N_22615,N_19122,N_15139);
xor U22616 (N_22616,N_18871,N_19013);
nor U22617 (N_22617,N_15009,N_16439);
nor U22618 (N_22618,N_16692,N_16257);
or U22619 (N_22619,N_16792,N_17018);
xor U22620 (N_22620,N_19555,N_17559);
xor U22621 (N_22621,N_19349,N_19319);
nand U22622 (N_22622,N_17713,N_16917);
nor U22623 (N_22623,N_18619,N_16126);
xnor U22624 (N_22624,N_18077,N_19705);
or U22625 (N_22625,N_19793,N_16646);
nor U22626 (N_22626,N_15334,N_17065);
nor U22627 (N_22627,N_18522,N_16360);
and U22628 (N_22628,N_18312,N_17293);
or U22629 (N_22629,N_19133,N_16760);
nor U22630 (N_22630,N_16964,N_17147);
or U22631 (N_22631,N_15480,N_15931);
xor U22632 (N_22632,N_18626,N_19678);
and U22633 (N_22633,N_19806,N_16240);
nand U22634 (N_22634,N_18516,N_18031);
xnor U22635 (N_22635,N_16409,N_19895);
and U22636 (N_22636,N_19118,N_15051);
nor U22637 (N_22637,N_17469,N_17110);
and U22638 (N_22638,N_19695,N_19541);
and U22639 (N_22639,N_18438,N_19060);
xor U22640 (N_22640,N_18225,N_17679);
and U22641 (N_22641,N_17072,N_15231);
nand U22642 (N_22642,N_17128,N_17811);
xnor U22643 (N_22643,N_15308,N_15739);
and U22644 (N_22644,N_19379,N_17418);
nand U22645 (N_22645,N_19059,N_16472);
nor U22646 (N_22646,N_15106,N_17189);
nand U22647 (N_22647,N_15590,N_17764);
or U22648 (N_22648,N_17905,N_16504);
or U22649 (N_22649,N_15582,N_15421);
and U22650 (N_22650,N_15787,N_17962);
nor U22651 (N_22651,N_19674,N_19224);
and U22652 (N_22652,N_18745,N_15406);
or U22653 (N_22653,N_19732,N_18660);
or U22654 (N_22654,N_19630,N_15636);
xnor U22655 (N_22655,N_16764,N_16659);
nand U22656 (N_22656,N_15401,N_17916);
xnor U22657 (N_22657,N_17256,N_17698);
and U22658 (N_22658,N_17346,N_18585);
or U22659 (N_22659,N_16072,N_17094);
xnor U22660 (N_22660,N_19928,N_16803);
or U22661 (N_22661,N_15669,N_17599);
nor U22662 (N_22662,N_17193,N_19849);
nor U22663 (N_22663,N_18102,N_16989);
or U22664 (N_22664,N_15433,N_17411);
xnor U22665 (N_22665,N_19965,N_18509);
or U22666 (N_22666,N_19250,N_18292);
or U22667 (N_22667,N_18326,N_18891);
and U22668 (N_22668,N_18803,N_17266);
and U22669 (N_22669,N_17445,N_16448);
and U22670 (N_22670,N_17362,N_19415);
or U22671 (N_22671,N_16453,N_19920);
or U22672 (N_22672,N_17402,N_16419);
xnor U22673 (N_22673,N_19516,N_19444);
nand U22674 (N_22674,N_16338,N_16175);
or U22675 (N_22675,N_16059,N_19843);
or U22676 (N_22676,N_17111,N_19011);
nor U22677 (N_22677,N_17950,N_15424);
xnor U22678 (N_22678,N_18006,N_18280);
or U22679 (N_22679,N_17385,N_17555);
nor U22680 (N_22680,N_17995,N_18335);
nor U22681 (N_22681,N_15148,N_15565);
or U22682 (N_22682,N_17600,N_16469);
and U22683 (N_22683,N_16845,N_15717);
or U22684 (N_22684,N_18982,N_18275);
and U22685 (N_22685,N_18284,N_16539);
nand U22686 (N_22686,N_15341,N_18513);
and U22687 (N_22687,N_17124,N_17184);
or U22688 (N_22688,N_19162,N_16775);
nand U22689 (N_22689,N_17745,N_15628);
and U22690 (N_22690,N_15491,N_17405);
nand U22691 (N_22691,N_16862,N_19222);
or U22692 (N_22692,N_15385,N_16803);
nor U22693 (N_22693,N_16885,N_15029);
and U22694 (N_22694,N_19925,N_18388);
nor U22695 (N_22695,N_18996,N_15224);
and U22696 (N_22696,N_17310,N_16474);
xor U22697 (N_22697,N_15418,N_16775);
or U22698 (N_22698,N_15589,N_18722);
xnor U22699 (N_22699,N_15529,N_16453);
xor U22700 (N_22700,N_16134,N_15146);
nand U22701 (N_22701,N_16990,N_19366);
or U22702 (N_22702,N_19828,N_15305);
or U22703 (N_22703,N_17894,N_18410);
or U22704 (N_22704,N_16846,N_18863);
xnor U22705 (N_22705,N_19452,N_18529);
xor U22706 (N_22706,N_17615,N_19195);
or U22707 (N_22707,N_19113,N_19956);
nand U22708 (N_22708,N_18570,N_16374);
nand U22709 (N_22709,N_18248,N_19627);
nand U22710 (N_22710,N_18584,N_15597);
and U22711 (N_22711,N_19534,N_17017);
nor U22712 (N_22712,N_15260,N_17467);
or U22713 (N_22713,N_19409,N_16141);
and U22714 (N_22714,N_16021,N_16854);
nand U22715 (N_22715,N_17331,N_19197);
and U22716 (N_22716,N_15753,N_19610);
nand U22717 (N_22717,N_16981,N_15740);
and U22718 (N_22718,N_16258,N_16830);
xnor U22719 (N_22719,N_16943,N_18902);
xnor U22720 (N_22720,N_15417,N_19452);
xnor U22721 (N_22721,N_16695,N_16830);
or U22722 (N_22722,N_18911,N_16670);
or U22723 (N_22723,N_19408,N_17970);
nor U22724 (N_22724,N_17957,N_18770);
nand U22725 (N_22725,N_19807,N_15539);
and U22726 (N_22726,N_15310,N_15831);
nor U22727 (N_22727,N_17983,N_18162);
xnor U22728 (N_22728,N_16769,N_15680);
nor U22729 (N_22729,N_16445,N_15003);
nand U22730 (N_22730,N_19736,N_18464);
and U22731 (N_22731,N_15717,N_19927);
nor U22732 (N_22732,N_17329,N_18957);
nand U22733 (N_22733,N_17163,N_19938);
nand U22734 (N_22734,N_19939,N_17865);
or U22735 (N_22735,N_18221,N_19766);
xnor U22736 (N_22736,N_18812,N_15689);
nand U22737 (N_22737,N_19446,N_17196);
nor U22738 (N_22738,N_17190,N_16547);
nor U22739 (N_22739,N_18312,N_15792);
or U22740 (N_22740,N_16972,N_16495);
xnor U22741 (N_22741,N_18428,N_16583);
nor U22742 (N_22742,N_17435,N_16316);
nand U22743 (N_22743,N_19495,N_16447);
xor U22744 (N_22744,N_17451,N_17000);
or U22745 (N_22745,N_17871,N_18597);
and U22746 (N_22746,N_15508,N_19494);
xor U22747 (N_22747,N_19167,N_18781);
xnor U22748 (N_22748,N_16470,N_17541);
nand U22749 (N_22749,N_17993,N_19975);
nand U22750 (N_22750,N_17285,N_16798);
xnor U22751 (N_22751,N_18209,N_17039);
xnor U22752 (N_22752,N_17194,N_18334);
nand U22753 (N_22753,N_18165,N_18643);
nor U22754 (N_22754,N_17978,N_18324);
xor U22755 (N_22755,N_18636,N_17618);
or U22756 (N_22756,N_16897,N_18223);
nor U22757 (N_22757,N_19785,N_17630);
and U22758 (N_22758,N_19461,N_16965);
or U22759 (N_22759,N_15180,N_18427);
nor U22760 (N_22760,N_19824,N_19203);
nand U22761 (N_22761,N_17667,N_15935);
nand U22762 (N_22762,N_19278,N_19014);
or U22763 (N_22763,N_16874,N_18479);
nor U22764 (N_22764,N_17961,N_18735);
nand U22765 (N_22765,N_15075,N_17841);
and U22766 (N_22766,N_18550,N_16067);
and U22767 (N_22767,N_17932,N_17759);
nand U22768 (N_22768,N_18904,N_16405);
xnor U22769 (N_22769,N_19920,N_15500);
nand U22770 (N_22770,N_16176,N_18113);
nor U22771 (N_22771,N_17295,N_17220);
and U22772 (N_22772,N_15678,N_17843);
nand U22773 (N_22773,N_18982,N_19676);
or U22774 (N_22774,N_18763,N_17883);
and U22775 (N_22775,N_18755,N_18279);
or U22776 (N_22776,N_19720,N_19372);
or U22777 (N_22777,N_16038,N_15574);
and U22778 (N_22778,N_16887,N_16913);
nor U22779 (N_22779,N_16057,N_15134);
or U22780 (N_22780,N_19075,N_19187);
or U22781 (N_22781,N_16132,N_15561);
xnor U22782 (N_22782,N_15736,N_15622);
xnor U22783 (N_22783,N_15762,N_19640);
or U22784 (N_22784,N_16334,N_17440);
nand U22785 (N_22785,N_17706,N_17674);
and U22786 (N_22786,N_16938,N_15041);
xor U22787 (N_22787,N_16091,N_17823);
or U22788 (N_22788,N_17171,N_19030);
nor U22789 (N_22789,N_19728,N_19537);
and U22790 (N_22790,N_15359,N_19619);
xor U22791 (N_22791,N_19878,N_17381);
nand U22792 (N_22792,N_16023,N_18759);
or U22793 (N_22793,N_19734,N_18281);
and U22794 (N_22794,N_19727,N_18285);
nor U22795 (N_22795,N_19556,N_15844);
nor U22796 (N_22796,N_19462,N_17030);
nor U22797 (N_22797,N_16412,N_16153);
or U22798 (N_22798,N_18763,N_17908);
and U22799 (N_22799,N_15856,N_18927);
and U22800 (N_22800,N_18852,N_19663);
and U22801 (N_22801,N_16798,N_17778);
and U22802 (N_22802,N_18815,N_18908);
xor U22803 (N_22803,N_16984,N_18735);
nor U22804 (N_22804,N_17907,N_16535);
and U22805 (N_22805,N_17315,N_18585);
nand U22806 (N_22806,N_16080,N_15593);
nand U22807 (N_22807,N_19271,N_18025);
nand U22808 (N_22808,N_15372,N_16330);
or U22809 (N_22809,N_19121,N_15070);
xor U22810 (N_22810,N_19227,N_18603);
and U22811 (N_22811,N_17820,N_18339);
or U22812 (N_22812,N_16742,N_16395);
xnor U22813 (N_22813,N_19350,N_16840);
or U22814 (N_22814,N_15885,N_18686);
xor U22815 (N_22815,N_16984,N_17284);
and U22816 (N_22816,N_15963,N_15354);
nor U22817 (N_22817,N_15206,N_15740);
nor U22818 (N_22818,N_15117,N_16552);
xnor U22819 (N_22819,N_19363,N_16715);
nor U22820 (N_22820,N_19976,N_19201);
and U22821 (N_22821,N_15331,N_16414);
xnor U22822 (N_22822,N_16877,N_16673);
or U22823 (N_22823,N_19230,N_18993);
nand U22824 (N_22824,N_17914,N_15114);
nor U22825 (N_22825,N_19573,N_17265);
nor U22826 (N_22826,N_18286,N_19053);
and U22827 (N_22827,N_18694,N_16711);
nor U22828 (N_22828,N_15317,N_18009);
nor U22829 (N_22829,N_18901,N_18381);
nor U22830 (N_22830,N_18915,N_16559);
nand U22831 (N_22831,N_16289,N_16816);
xor U22832 (N_22832,N_19122,N_18672);
xnor U22833 (N_22833,N_19703,N_18936);
nand U22834 (N_22834,N_17880,N_18579);
and U22835 (N_22835,N_16685,N_18439);
or U22836 (N_22836,N_18854,N_17889);
nor U22837 (N_22837,N_15537,N_19779);
or U22838 (N_22838,N_15049,N_17417);
nor U22839 (N_22839,N_16158,N_17433);
or U22840 (N_22840,N_16438,N_15191);
and U22841 (N_22841,N_19489,N_18875);
nand U22842 (N_22842,N_19244,N_16919);
and U22843 (N_22843,N_17259,N_15867);
nand U22844 (N_22844,N_18090,N_15223);
xnor U22845 (N_22845,N_19436,N_15332);
or U22846 (N_22846,N_19929,N_16745);
or U22847 (N_22847,N_15827,N_18837);
xor U22848 (N_22848,N_16010,N_19482);
or U22849 (N_22849,N_18398,N_19437);
nor U22850 (N_22850,N_15181,N_17551);
and U22851 (N_22851,N_15049,N_17757);
nand U22852 (N_22852,N_15264,N_17321);
or U22853 (N_22853,N_17347,N_18383);
nor U22854 (N_22854,N_16715,N_16877);
nand U22855 (N_22855,N_15425,N_16004);
nor U22856 (N_22856,N_15928,N_17338);
xor U22857 (N_22857,N_18825,N_16012);
and U22858 (N_22858,N_17740,N_15435);
xnor U22859 (N_22859,N_16324,N_17709);
nand U22860 (N_22860,N_17901,N_16804);
nand U22861 (N_22861,N_15367,N_18478);
or U22862 (N_22862,N_16080,N_17284);
nand U22863 (N_22863,N_19594,N_18383);
xnor U22864 (N_22864,N_16497,N_18453);
and U22865 (N_22865,N_15164,N_17846);
xnor U22866 (N_22866,N_18371,N_15389);
and U22867 (N_22867,N_15526,N_17932);
xnor U22868 (N_22868,N_15038,N_15292);
or U22869 (N_22869,N_17386,N_17049);
nand U22870 (N_22870,N_16756,N_16266);
xnor U22871 (N_22871,N_19364,N_17177);
nor U22872 (N_22872,N_15589,N_18617);
or U22873 (N_22873,N_18181,N_16680);
xor U22874 (N_22874,N_19688,N_18363);
nor U22875 (N_22875,N_15065,N_16157);
or U22876 (N_22876,N_16347,N_16067);
or U22877 (N_22877,N_15481,N_15562);
or U22878 (N_22878,N_17170,N_15269);
nor U22879 (N_22879,N_16052,N_15762);
and U22880 (N_22880,N_18408,N_19897);
xor U22881 (N_22881,N_17210,N_18176);
xor U22882 (N_22882,N_17940,N_16776);
or U22883 (N_22883,N_16043,N_18419);
or U22884 (N_22884,N_17583,N_16849);
xnor U22885 (N_22885,N_17344,N_18372);
nand U22886 (N_22886,N_19555,N_19182);
and U22887 (N_22887,N_19474,N_17248);
nand U22888 (N_22888,N_18114,N_17295);
xor U22889 (N_22889,N_19677,N_15146);
xor U22890 (N_22890,N_19142,N_15064);
nand U22891 (N_22891,N_15160,N_15321);
nand U22892 (N_22892,N_19154,N_15856);
or U22893 (N_22893,N_18078,N_16194);
nor U22894 (N_22894,N_19432,N_18942);
and U22895 (N_22895,N_18860,N_19573);
or U22896 (N_22896,N_18398,N_16897);
and U22897 (N_22897,N_17212,N_19861);
nor U22898 (N_22898,N_18363,N_15481);
and U22899 (N_22899,N_18613,N_17726);
or U22900 (N_22900,N_19699,N_17042);
and U22901 (N_22901,N_17782,N_16715);
xnor U22902 (N_22902,N_19674,N_17402);
nor U22903 (N_22903,N_16867,N_17842);
or U22904 (N_22904,N_15851,N_17457);
and U22905 (N_22905,N_16192,N_15625);
nand U22906 (N_22906,N_15063,N_17874);
or U22907 (N_22907,N_15280,N_19308);
nor U22908 (N_22908,N_16043,N_18963);
or U22909 (N_22909,N_16428,N_18661);
nand U22910 (N_22910,N_16766,N_18484);
and U22911 (N_22911,N_16165,N_18700);
or U22912 (N_22912,N_15083,N_18098);
or U22913 (N_22913,N_16072,N_18270);
nand U22914 (N_22914,N_17326,N_15469);
and U22915 (N_22915,N_18648,N_19296);
or U22916 (N_22916,N_16179,N_19252);
xnor U22917 (N_22917,N_19020,N_17663);
nand U22918 (N_22918,N_18767,N_15300);
nand U22919 (N_22919,N_17851,N_19937);
nand U22920 (N_22920,N_17665,N_15031);
xor U22921 (N_22921,N_18099,N_15757);
nand U22922 (N_22922,N_17164,N_17720);
xor U22923 (N_22923,N_15650,N_18987);
nand U22924 (N_22924,N_16438,N_18372);
nor U22925 (N_22925,N_18245,N_19884);
and U22926 (N_22926,N_16568,N_18895);
nand U22927 (N_22927,N_18870,N_17559);
and U22928 (N_22928,N_15148,N_18539);
nor U22929 (N_22929,N_19319,N_16470);
nor U22930 (N_22930,N_15509,N_19324);
nand U22931 (N_22931,N_16278,N_17146);
xnor U22932 (N_22932,N_19584,N_19664);
xnor U22933 (N_22933,N_16739,N_15734);
nor U22934 (N_22934,N_18319,N_15006);
xor U22935 (N_22935,N_17319,N_19404);
nor U22936 (N_22936,N_15006,N_19477);
nor U22937 (N_22937,N_16692,N_15178);
and U22938 (N_22938,N_15344,N_19674);
and U22939 (N_22939,N_19693,N_19179);
nor U22940 (N_22940,N_18610,N_17669);
or U22941 (N_22941,N_16638,N_15724);
nand U22942 (N_22942,N_18120,N_17739);
and U22943 (N_22943,N_17424,N_18883);
nor U22944 (N_22944,N_18444,N_15734);
xor U22945 (N_22945,N_15068,N_17120);
nor U22946 (N_22946,N_16224,N_17466);
nand U22947 (N_22947,N_19569,N_17354);
and U22948 (N_22948,N_17964,N_19577);
xnor U22949 (N_22949,N_18267,N_17812);
xor U22950 (N_22950,N_19935,N_15577);
or U22951 (N_22951,N_19854,N_18611);
and U22952 (N_22952,N_15035,N_19431);
or U22953 (N_22953,N_15839,N_16193);
nor U22954 (N_22954,N_17335,N_16119);
and U22955 (N_22955,N_18226,N_15991);
or U22956 (N_22956,N_16013,N_19559);
xnor U22957 (N_22957,N_19481,N_16513);
nor U22958 (N_22958,N_18935,N_16030);
or U22959 (N_22959,N_18469,N_18965);
and U22960 (N_22960,N_17301,N_15353);
nor U22961 (N_22961,N_19878,N_18671);
and U22962 (N_22962,N_19602,N_16056);
nand U22963 (N_22963,N_19379,N_15127);
or U22964 (N_22964,N_19121,N_17808);
nor U22965 (N_22965,N_15374,N_18598);
nor U22966 (N_22966,N_15092,N_17718);
and U22967 (N_22967,N_19817,N_15186);
nand U22968 (N_22968,N_17106,N_19661);
xor U22969 (N_22969,N_15670,N_16260);
nor U22970 (N_22970,N_19623,N_18754);
nor U22971 (N_22971,N_18287,N_16601);
xor U22972 (N_22972,N_15934,N_15204);
or U22973 (N_22973,N_18609,N_19012);
nand U22974 (N_22974,N_18182,N_16356);
xor U22975 (N_22975,N_18787,N_17979);
and U22976 (N_22976,N_15563,N_19078);
and U22977 (N_22977,N_18106,N_18874);
and U22978 (N_22978,N_18147,N_16488);
and U22979 (N_22979,N_15233,N_17620);
or U22980 (N_22980,N_18194,N_15442);
nand U22981 (N_22981,N_16281,N_19635);
nor U22982 (N_22982,N_17513,N_18501);
xnor U22983 (N_22983,N_17190,N_19708);
and U22984 (N_22984,N_18029,N_15397);
or U22985 (N_22985,N_16395,N_18432);
nand U22986 (N_22986,N_17318,N_15244);
nor U22987 (N_22987,N_16969,N_15094);
xor U22988 (N_22988,N_18920,N_18503);
and U22989 (N_22989,N_16852,N_18284);
or U22990 (N_22990,N_17230,N_16291);
xnor U22991 (N_22991,N_18150,N_19374);
or U22992 (N_22992,N_18649,N_18725);
nand U22993 (N_22993,N_18678,N_16186);
or U22994 (N_22994,N_15946,N_16109);
and U22995 (N_22995,N_15830,N_16486);
xnor U22996 (N_22996,N_17170,N_19468);
and U22997 (N_22997,N_18697,N_18819);
or U22998 (N_22998,N_19266,N_16690);
nand U22999 (N_22999,N_19167,N_18303);
and U23000 (N_23000,N_16033,N_18647);
and U23001 (N_23001,N_16936,N_18807);
nand U23002 (N_23002,N_19624,N_16780);
xor U23003 (N_23003,N_19782,N_15067);
and U23004 (N_23004,N_18767,N_15418);
and U23005 (N_23005,N_18673,N_16429);
nand U23006 (N_23006,N_15786,N_15370);
xor U23007 (N_23007,N_18922,N_16742);
nand U23008 (N_23008,N_19407,N_17615);
or U23009 (N_23009,N_19400,N_15239);
and U23010 (N_23010,N_17138,N_16810);
and U23011 (N_23011,N_19457,N_17628);
nand U23012 (N_23012,N_15140,N_17092);
nand U23013 (N_23013,N_16692,N_18128);
xnor U23014 (N_23014,N_19374,N_15296);
xor U23015 (N_23015,N_16218,N_16112);
nand U23016 (N_23016,N_15818,N_18432);
and U23017 (N_23017,N_18444,N_16365);
and U23018 (N_23018,N_17428,N_16417);
xor U23019 (N_23019,N_17318,N_18163);
and U23020 (N_23020,N_17777,N_16075);
xor U23021 (N_23021,N_18414,N_19782);
nand U23022 (N_23022,N_17019,N_19272);
and U23023 (N_23023,N_15615,N_17167);
xnor U23024 (N_23024,N_19565,N_17021);
xnor U23025 (N_23025,N_16571,N_19091);
xnor U23026 (N_23026,N_17790,N_15850);
nand U23027 (N_23027,N_16186,N_16637);
nand U23028 (N_23028,N_19352,N_17434);
nand U23029 (N_23029,N_19275,N_17521);
or U23030 (N_23030,N_19798,N_16450);
nor U23031 (N_23031,N_19584,N_17767);
xor U23032 (N_23032,N_15367,N_16122);
or U23033 (N_23033,N_19272,N_17651);
nor U23034 (N_23034,N_16645,N_16086);
or U23035 (N_23035,N_18189,N_17616);
or U23036 (N_23036,N_18691,N_16880);
or U23037 (N_23037,N_18209,N_19336);
or U23038 (N_23038,N_19848,N_18967);
or U23039 (N_23039,N_18741,N_16670);
nor U23040 (N_23040,N_18050,N_17342);
or U23041 (N_23041,N_17429,N_19982);
nor U23042 (N_23042,N_17997,N_15992);
nor U23043 (N_23043,N_15972,N_16807);
xnor U23044 (N_23044,N_16526,N_19601);
nor U23045 (N_23045,N_18208,N_17218);
or U23046 (N_23046,N_15057,N_19002);
and U23047 (N_23047,N_16057,N_19977);
nand U23048 (N_23048,N_17604,N_17161);
and U23049 (N_23049,N_16171,N_16282);
xor U23050 (N_23050,N_18087,N_18669);
or U23051 (N_23051,N_18910,N_17604);
or U23052 (N_23052,N_18307,N_19806);
nor U23053 (N_23053,N_16467,N_15620);
nor U23054 (N_23054,N_16778,N_15018);
or U23055 (N_23055,N_17919,N_15614);
nor U23056 (N_23056,N_17463,N_15474);
nand U23057 (N_23057,N_17275,N_18256);
nand U23058 (N_23058,N_17329,N_18819);
or U23059 (N_23059,N_16702,N_19018);
or U23060 (N_23060,N_15953,N_19271);
xnor U23061 (N_23061,N_15093,N_16101);
or U23062 (N_23062,N_19409,N_18194);
nor U23063 (N_23063,N_16032,N_17012);
nand U23064 (N_23064,N_16669,N_16823);
or U23065 (N_23065,N_18240,N_18890);
nor U23066 (N_23066,N_19017,N_19946);
xnor U23067 (N_23067,N_15575,N_15110);
nand U23068 (N_23068,N_15716,N_18477);
or U23069 (N_23069,N_16682,N_18045);
xor U23070 (N_23070,N_18352,N_15429);
nand U23071 (N_23071,N_17514,N_17595);
or U23072 (N_23072,N_17631,N_19180);
nor U23073 (N_23073,N_15304,N_15092);
nand U23074 (N_23074,N_19637,N_15057);
and U23075 (N_23075,N_18714,N_17736);
and U23076 (N_23076,N_17384,N_17049);
nand U23077 (N_23077,N_17980,N_18873);
nor U23078 (N_23078,N_16234,N_15679);
xnor U23079 (N_23079,N_15208,N_19612);
nand U23080 (N_23080,N_17174,N_18566);
nor U23081 (N_23081,N_18781,N_16184);
xor U23082 (N_23082,N_16424,N_17054);
nand U23083 (N_23083,N_17638,N_15012);
xor U23084 (N_23084,N_17777,N_18466);
or U23085 (N_23085,N_17018,N_16321);
or U23086 (N_23086,N_15335,N_15177);
and U23087 (N_23087,N_16252,N_19667);
or U23088 (N_23088,N_16509,N_16595);
xnor U23089 (N_23089,N_15626,N_15380);
nor U23090 (N_23090,N_17873,N_16380);
nand U23091 (N_23091,N_17060,N_17110);
xnor U23092 (N_23092,N_16362,N_16797);
and U23093 (N_23093,N_17200,N_18500);
nor U23094 (N_23094,N_15307,N_17255);
xor U23095 (N_23095,N_18861,N_18546);
nor U23096 (N_23096,N_19154,N_18752);
and U23097 (N_23097,N_16230,N_16412);
xor U23098 (N_23098,N_16788,N_19204);
nor U23099 (N_23099,N_15731,N_18388);
nor U23100 (N_23100,N_18403,N_18548);
nand U23101 (N_23101,N_16021,N_17934);
nand U23102 (N_23102,N_16361,N_17037);
xor U23103 (N_23103,N_16171,N_19182);
and U23104 (N_23104,N_15221,N_19724);
and U23105 (N_23105,N_18173,N_15760);
nor U23106 (N_23106,N_17102,N_18050);
nand U23107 (N_23107,N_19691,N_17755);
and U23108 (N_23108,N_18982,N_15276);
xnor U23109 (N_23109,N_17240,N_16066);
and U23110 (N_23110,N_16878,N_17558);
or U23111 (N_23111,N_15204,N_19299);
and U23112 (N_23112,N_15632,N_16569);
nand U23113 (N_23113,N_18171,N_19485);
nand U23114 (N_23114,N_17838,N_17628);
xor U23115 (N_23115,N_15874,N_16501);
and U23116 (N_23116,N_18483,N_16878);
and U23117 (N_23117,N_17663,N_19897);
and U23118 (N_23118,N_16671,N_17658);
nor U23119 (N_23119,N_19610,N_17958);
nand U23120 (N_23120,N_18556,N_18161);
and U23121 (N_23121,N_17130,N_19106);
and U23122 (N_23122,N_17225,N_19754);
nand U23123 (N_23123,N_19738,N_17214);
nand U23124 (N_23124,N_16287,N_18674);
and U23125 (N_23125,N_17810,N_16998);
or U23126 (N_23126,N_18863,N_19723);
or U23127 (N_23127,N_15749,N_17651);
nor U23128 (N_23128,N_15398,N_15472);
nor U23129 (N_23129,N_19735,N_16070);
nand U23130 (N_23130,N_15818,N_15080);
nor U23131 (N_23131,N_17425,N_17073);
nand U23132 (N_23132,N_17012,N_18844);
and U23133 (N_23133,N_18800,N_15768);
and U23134 (N_23134,N_16960,N_19350);
or U23135 (N_23135,N_17564,N_16797);
xnor U23136 (N_23136,N_19896,N_15076);
and U23137 (N_23137,N_16223,N_18884);
nor U23138 (N_23138,N_19163,N_15131);
nand U23139 (N_23139,N_15781,N_18997);
nand U23140 (N_23140,N_16042,N_17048);
xnor U23141 (N_23141,N_17103,N_15716);
and U23142 (N_23142,N_16903,N_15629);
nor U23143 (N_23143,N_18449,N_18990);
and U23144 (N_23144,N_17209,N_19460);
nor U23145 (N_23145,N_17491,N_16273);
and U23146 (N_23146,N_17766,N_16426);
xor U23147 (N_23147,N_17185,N_15099);
xnor U23148 (N_23148,N_16464,N_18371);
or U23149 (N_23149,N_17757,N_19759);
and U23150 (N_23150,N_15958,N_15917);
or U23151 (N_23151,N_17987,N_19820);
or U23152 (N_23152,N_18415,N_15817);
or U23153 (N_23153,N_16805,N_16079);
xnor U23154 (N_23154,N_15555,N_19002);
and U23155 (N_23155,N_17727,N_17618);
and U23156 (N_23156,N_19535,N_15999);
or U23157 (N_23157,N_18541,N_18033);
xnor U23158 (N_23158,N_17128,N_17887);
and U23159 (N_23159,N_18958,N_15565);
xnor U23160 (N_23160,N_17010,N_16108);
nand U23161 (N_23161,N_16487,N_19001);
xor U23162 (N_23162,N_17023,N_19941);
and U23163 (N_23163,N_15369,N_18525);
nor U23164 (N_23164,N_15984,N_15011);
xor U23165 (N_23165,N_19463,N_19304);
xor U23166 (N_23166,N_16579,N_16058);
or U23167 (N_23167,N_17029,N_19070);
nor U23168 (N_23168,N_16630,N_17178);
or U23169 (N_23169,N_19568,N_17694);
nor U23170 (N_23170,N_16848,N_15599);
nand U23171 (N_23171,N_18475,N_18772);
nor U23172 (N_23172,N_18334,N_18862);
nand U23173 (N_23173,N_15895,N_17407);
nand U23174 (N_23174,N_16051,N_16364);
xnor U23175 (N_23175,N_15642,N_15817);
nand U23176 (N_23176,N_17890,N_16390);
or U23177 (N_23177,N_15701,N_15764);
nand U23178 (N_23178,N_18639,N_19512);
or U23179 (N_23179,N_17240,N_19897);
or U23180 (N_23180,N_18798,N_16101);
or U23181 (N_23181,N_17223,N_17189);
xor U23182 (N_23182,N_19429,N_16188);
nor U23183 (N_23183,N_15219,N_17991);
xnor U23184 (N_23184,N_15040,N_17761);
nand U23185 (N_23185,N_19877,N_16715);
or U23186 (N_23186,N_19302,N_16835);
nand U23187 (N_23187,N_18206,N_18662);
or U23188 (N_23188,N_16399,N_16741);
and U23189 (N_23189,N_19907,N_18909);
or U23190 (N_23190,N_19447,N_15295);
xor U23191 (N_23191,N_16154,N_19086);
xor U23192 (N_23192,N_17869,N_16337);
or U23193 (N_23193,N_17331,N_17179);
and U23194 (N_23194,N_18127,N_18796);
nor U23195 (N_23195,N_17214,N_17163);
nor U23196 (N_23196,N_16786,N_16275);
or U23197 (N_23197,N_16170,N_19080);
and U23198 (N_23198,N_15575,N_17131);
xor U23199 (N_23199,N_17289,N_17951);
or U23200 (N_23200,N_15493,N_19677);
or U23201 (N_23201,N_15336,N_16745);
or U23202 (N_23202,N_17442,N_19875);
or U23203 (N_23203,N_18115,N_17746);
nand U23204 (N_23204,N_17833,N_19450);
nand U23205 (N_23205,N_18785,N_19651);
and U23206 (N_23206,N_19431,N_15017);
xor U23207 (N_23207,N_16425,N_18449);
and U23208 (N_23208,N_19498,N_19199);
nor U23209 (N_23209,N_16683,N_19414);
xnor U23210 (N_23210,N_17564,N_18227);
or U23211 (N_23211,N_15917,N_17872);
xnor U23212 (N_23212,N_19978,N_18785);
nor U23213 (N_23213,N_18283,N_18816);
and U23214 (N_23214,N_16242,N_15744);
or U23215 (N_23215,N_18415,N_18334);
xnor U23216 (N_23216,N_17717,N_19541);
and U23217 (N_23217,N_19193,N_18662);
or U23218 (N_23218,N_18203,N_19951);
xnor U23219 (N_23219,N_16586,N_17286);
or U23220 (N_23220,N_17727,N_16433);
nor U23221 (N_23221,N_15833,N_16650);
nor U23222 (N_23222,N_16909,N_18538);
nand U23223 (N_23223,N_16273,N_17135);
or U23224 (N_23224,N_17130,N_16385);
and U23225 (N_23225,N_19169,N_19500);
nor U23226 (N_23226,N_16480,N_17558);
nand U23227 (N_23227,N_19129,N_17811);
nand U23228 (N_23228,N_17553,N_19621);
xor U23229 (N_23229,N_19880,N_17277);
or U23230 (N_23230,N_16212,N_15610);
nor U23231 (N_23231,N_18181,N_19174);
and U23232 (N_23232,N_17700,N_16815);
or U23233 (N_23233,N_16947,N_17304);
nor U23234 (N_23234,N_17015,N_19098);
nor U23235 (N_23235,N_15445,N_18928);
nor U23236 (N_23236,N_15028,N_19302);
and U23237 (N_23237,N_15779,N_17607);
xor U23238 (N_23238,N_15176,N_16347);
and U23239 (N_23239,N_19911,N_18161);
nor U23240 (N_23240,N_15606,N_18672);
nand U23241 (N_23241,N_15478,N_16043);
xnor U23242 (N_23242,N_19389,N_16630);
xor U23243 (N_23243,N_18976,N_19822);
nand U23244 (N_23244,N_15297,N_19102);
nor U23245 (N_23245,N_15214,N_15552);
and U23246 (N_23246,N_15783,N_18317);
or U23247 (N_23247,N_17441,N_17626);
nor U23248 (N_23248,N_16481,N_19131);
nor U23249 (N_23249,N_16162,N_16500);
nand U23250 (N_23250,N_18909,N_17972);
nor U23251 (N_23251,N_17617,N_15512);
xnor U23252 (N_23252,N_15713,N_19968);
and U23253 (N_23253,N_16486,N_17651);
or U23254 (N_23254,N_19098,N_15538);
and U23255 (N_23255,N_19684,N_15357);
xnor U23256 (N_23256,N_16144,N_15367);
xor U23257 (N_23257,N_18396,N_19014);
nand U23258 (N_23258,N_18531,N_15203);
and U23259 (N_23259,N_15147,N_19318);
nand U23260 (N_23260,N_19195,N_17925);
or U23261 (N_23261,N_18916,N_19677);
nor U23262 (N_23262,N_17704,N_19861);
nor U23263 (N_23263,N_15583,N_18663);
xor U23264 (N_23264,N_15772,N_15085);
xor U23265 (N_23265,N_18922,N_18131);
or U23266 (N_23266,N_15136,N_16276);
or U23267 (N_23267,N_16451,N_15385);
and U23268 (N_23268,N_19524,N_17663);
nor U23269 (N_23269,N_19591,N_17331);
nand U23270 (N_23270,N_18741,N_19092);
nand U23271 (N_23271,N_18858,N_17786);
nand U23272 (N_23272,N_18233,N_18104);
and U23273 (N_23273,N_18694,N_16970);
or U23274 (N_23274,N_17043,N_18506);
xnor U23275 (N_23275,N_15326,N_15217);
nor U23276 (N_23276,N_17804,N_17670);
xor U23277 (N_23277,N_16929,N_18145);
nand U23278 (N_23278,N_18111,N_18930);
or U23279 (N_23279,N_16616,N_19147);
and U23280 (N_23280,N_17867,N_16074);
or U23281 (N_23281,N_18302,N_17220);
nor U23282 (N_23282,N_18478,N_18535);
and U23283 (N_23283,N_17620,N_19027);
or U23284 (N_23284,N_17467,N_18227);
or U23285 (N_23285,N_16747,N_19668);
nor U23286 (N_23286,N_19933,N_19190);
and U23287 (N_23287,N_16204,N_16212);
nand U23288 (N_23288,N_18248,N_19703);
nand U23289 (N_23289,N_17639,N_18168);
or U23290 (N_23290,N_15080,N_19375);
nand U23291 (N_23291,N_19677,N_17223);
xnor U23292 (N_23292,N_16653,N_19195);
and U23293 (N_23293,N_19451,N_16544);
or U23294 (N_23294,N_16612,N_17024);
nor U23295 (N_23295,N_18326,N_17367);
nand U23296 (N_23296,N_15683,N_17112);
nand U23297 (N_23297,N_19717,N_15897);
nand U23298 (N_23298,N_18474,N_16286);
xnor U23299 (N_23299,N_18895,N_17349);
and U23300 (N_23300,N_19282,N_18737);
or U23301 (N_23301,N_17246,N_17534);
or U23302 (N_23302,N_19139,N_15841);
xor U23303 (N_23303,N_15313,N_18646);
or U23304 (N_23304,N_19647,N_17879);
and U23305 (N_23305,N_16410,N_17632);
and U23306 (N_23306,N_16074,N_16726);
xor U23307 (N_23307,N_15637,N_15930);
xnor U23308 (N_23308,N_17001,N_18015);
or U23309 (N_23309,N_16827,N_19815);
or U23310 (N_23310,N_15258,N_18801);
and U23311 (N_23311,N_18614,N_18055);
nand U23312 (N_23312,N_17508,N_16390);
and U23313 (N_23313,N_19744,N_16602);
nor U23314 (N_23314,N_18880,N_15582);
and U23315 (N_23315,N_17424,N_15508);
nor U23316 (N_23316,N_17427,N_15834);
or U23317 (N_23317,N_16622,N_19765);
or U23318 (N_23318,N_16906,N_18443);
xnor U23319 (N_23319,N_16913,N_18763);
xor U23320 (N_23320,N_18670,N_18202);
nand U23321 (N_23321,N_19041,N_15532);
or U23322 (N_23322,N_18114,N_19191);
nor U23323 (N_23323,N_17399,N_15790);
or U23324 (N_23324,N_18175,N_15619);
nand U23325 (N_23325,N_17521,N_17538);
or U23326 (N_23326,N_17008,N_19362);
or U23327 (N_23327,N_17816,N_18559);
xor U23328 (N_23328,N_17075,N_16096);
xor U23329 (N_23329,N_19399,N_16836);
or U23330 (N_23330,N_16114,N_19187);
or U23331 (N_23331,N_18609,N_17682);
xnor U23332 (N_23332,N_19424,N_17942);
or U23333 (N_23333,N_19930,N_16146);
nor U23334 (N_23334,N_16455,N_18719);
nand U23335 (N_23335,N_19974,N_17490);
nor U23336 (N_23336,N_19563,N_16577);
nand U23337 (N_23337,N_15299,N_19057);
and U23338 (N_23338,N_16296,N_18998);
xnor U23339 (N_23339,N_19945,N_19221);
and U23340 (N_23340,N_15155,N_19967);
or U23341 (N_23341,N_19422,N_15914);
nand U23342 (N_23342,N_17030,N_15030);
xor U23343 (N_23343,N_17461,N_18814);
xor U23344 (N_23344,N_17509,N_15283);
nor U23345 (N_23345,N_19292,N_18508);
xnor U23346 (N_23346,N_16686,N_16261);
or U23347 (N_23347,N_18823,N_19232);
nor U23348 (N_23348,N_19526,N_15528);
nor U23349 (N_23349,N_16002,N_17931);
xor U23350 (N_23350,N_18940,N_17545);
xor U23351 (N_23351,N_19310,N_16281);
xnor U23352 (N_23352,N_15868,N_18626);
xnor U23353 (N_23353,N_15199,N_19757);
xnor U23354 (N_23354,N_15965,N_17251);
nor U23355 (N_23355,N_18572,N_17800);
nand U23356 (N_23356,N_17994,N_19026);
nand U23357 (N_23357,N_16663,N_15110);
xor U23358 (N_23358,N_19067,N_15620);
xnor U23359 (N_23359,N_15733,N_16867);
and U23360 (N_23360,N_18082,N_15006);
nand U23361 (N_23361,N_16944,N_16755);
xnor U23362 (N_23362,N_16585,N_15731);
nor U23363 (N_23363,N_15086,N_18631);
and U23364 (N_23364,N_19875,N_17234);
nand U23365 (N_23365,N_19531,N_18620);
nand U23366 (N_23366,N_18202,N_18192);
nand U23367 (N_23367,N_17879,N_17032);
xor U23368 (N_23368,N_17773,N_15151);
nand U23369 (N_23369,N_16765,N_16538);
nor U23370 (N_23370,N_16926,N_19142);
xor U23371 (N_23371,N_18924,N_16851);
or U23372 (N_23372,N_18950,N_18591);
nand U23373 (N_23373,N_15624,N_19563);
or U23374 (N_23374,N_15360,N_19763);
nor U23375 (N_23375,N_19019,N_18155);
nor U23376 (N_23376,N_17158,N_16529);
and U23377 (N_23377,N_19426,N_18236);
nor U23378 (N_23378,N_19252,N_17765);
nand U23379 (N_23379,N_19177,N_19094);
or U23380 (N_23380,N_18570,N_15330);
nor U23381 (N_23381,N_18102,N_16264);
nor U23382 (N_23382,N_19638,N_16154);
nor U23383 (N_23383,N_19507,N_15934);
nor U23384 (N_23384,N_19397,N_15950);
nor U23385 (N_23385,N_16201,N_15578);
nor U23386 (N_23386,N_17182,N_18809);
nand U23387 (N_23387,N_17682,N_19885);
xnor U23388 (N_23388,N_17420,N_18822);
nand U23389 (N_23389,N_15990,N_17417);
nor U23390 (N_23390,N_17430,N_18622);
or U23391 (N_23391,N_17640,N_19141);
or U23392 (N_23392,N_17672,N_16129);
nand U23393 (N_23393,N_16102,N_17139);
and U23394 (N_23394,N_15692,N_18720);
or U23395 (N_23395,N_17633,N_15726);
or U23396 (N_23396,N_15949,N_16827);
nand U23397 (N_23397,N_18450,N_18150);
or U23398 (N_23398,N_17135,N_15363);
nor U23399 (N_23399,N_15349,N_16833);
nand U23400 (N_23400,N_15221,N_16826);
nor U23401 (N_23401,N_18719,N_15861);
nand U23402 (N_23402,N_19955,N_17611);
nor U23403 (N_23403,N_17024,N_18633);
or U23404 (N_23404,N_16346,N_17717);
or U23405 (N_23405,N_16777,N_18569);
nand U23406 (N_23406,N_16919,N_17642);
xnor U23407 (N_23407,N_19519,N_19630);
or U23408 (N_23408,N_19269,N_19268);
or U23409 (N_23409,N_15014,N_19933);
nor U23410 (N_23410,N_17674,N_16472);
nand U23411 (N_23411,N_19517,N_17693);
nand U23412 (N_23412,N_17179,N_19707);
or U23413 (N_23413,N_19288,N_19172);
and U23414 (N_23414,N_19050,N_15969);
and U23415 (N_23415,N_15219,N_19183);
nand U23416 (N_23416,N_15453,N_19303);
nand U23417 (N_23417,N_19885,N_18793);
xor U23418 (N_23418,N_16533,N_17030);
and U23419 (N_23419,N_16336,N_17299);
xnor U23420 (N_23420,N_15756,N_18229);
nor U23421 (N_23421,N_19528,N_18368);
xnor U23422 (N_23422,N_19105,N_17323);
xnor U23423 (N_23423,N_17946,N_17712);
and U23424 (N_23424,N_15091,N_19303);
and U23425 (N_23425,N_16599,N_19941);
or U23426 (N_23426,N_16476,N_19865);
and U23427 (N_23427,N_19713,N_15641);
or U23428 (N_23428,N_16299,N_19366);
nor U23429 (N_23429,N_19618,N_17616);
or U23430 (N_23430,N_16135,N_17955);
or U23431 (N_23431,N_15440,N_18612);
or U23432 (N_23432,N_17985,N_16690);
xor U23433 (N_23433,N_16682,N_18871);
nor U23434 (N_23434,N_18152,N_18779);
and U23435 (N_23435,N_15344,N_18693);
and U23436 (N_23436,N_16227,N_15681);
nand U23437 (N_23437,N_19651,N_15828);
xnor U23438 (N_23438,N_18529,N_16369);
or U23439 (N_23439,N_18074,N_19804);
and U23440 (N_23440,N_17902,N_16840);
xnor U23441 (N_23441,N_19745,N_17065);
or U23442 (N_23442,N_15402,N_19445);
xor U23443 (N_23443,N_16466,N_19858);
and U23444 (N_23444,N_18791,N_16982);
xor U23445 (N_23445,N_19198,N_16937);
nor U23446 (N_23446,N_18559,N_15933);
and U23447 (N_23447,N_17603,N_17334);
or U23448 (N_23448,N_19508,N_19326);
xnor U23449 (N_23449,N_16652,N_16026);
nor U23450 (N_23450,N_15674,N_15339);
nor U23451 (N_23451,N_17802,N_15850);
nand U23452 (N_23452,N_19796,N_18526);
xor U23453 (N_23453,N_15958,N_18525);
xor U23454 (N_23454,N_17366,N_15869);
nand U23455 (N_23455,N_15703,N_16524);
and U23456 (N_23456,N_18118,N_18882);
and U23457 (N_23457,N_17668,N_16994);
and U23458 (N_23458,N_15929,N_19030);
or U23459 (N_23459,N_15266,N_19169);
nor U23460 (N_23460,N_19957,N_19965);
nor U23461 (N_23461,N_19583,N_15016);
xnor U23462 (N_23462,N_19554,N_17328);
nor U23463 (N_23463,N_15722,N_19230);
nor U23464 (N_23464,N_16527,N_15489);
nand U23465 (N_23465,N_15740,N_16420);
nor U23466 (N_23466,N_17795,N_18014);
nand U23467 (N_23467,N_16769,N_15944);
or U23468 (N_23468,N_18263,N_18193);
or U23469 (N_23469,N_19173,N_17265);
nor U23470 (N_23470,N_18588,N_18227);
nor U23471 (N_23471,N_19584,N_16504);
nand U23472 (N_23472,N_18436,N_16163);
nand U23473 (N_23473,N_18931,N_19308);
or U23474 (N_23474,N_16089,N_16236);
nand U23475 (N_23475,N_16998,N_15575);
and U23476 (N_23476,N_15768,N_16573);
nand U23477 (N_23477,N_16953,N_17245);
and U23478 (N_23478,N_19019,N_19111);
or U23479 (N_23479,N_16826,N_18076);
nand U23480 (N_23480,N_15815,N_19472);
nand U23481 (N_23481,N_15863,N_18665);
nand U23482 (N_23482,N_17262,N_17978);
and U23483 (N_23483,N_18512,N_16874);
and U23484 (N_23484,N_15052,N_16874);
and U23485 (N_23485,N_15108,N_19972);
or U23486 (N_23486,N_19271,N_18219);
nand U23487 (N_23487,N_15747,N_17343);
or U23488 (N_23488,N_16255,N_19495);
nor U23489 (N_23489,N_19012,N_17985);
and U23490 (N_23490,N_19385,N_17309);
or U23491 (N_23491,N_19976,N_19325);
nand U23492 (N_23492,N_15438,N_16389);
or U23493 (N_23493,N_15670,N_17890);
nor U23494 (N_23494,N_17364,N_15677);
and U23495 (N_23495,N_17066,N_16178);
nand U23496 (N_23496,N_15129,N_16109);
or U23497 (N_23497,N_19837,N_18348);
xor U23498 (N_23498,N_18138,N_15573);
xnor U23499 (N_23499,N_18730,N_17154);
nor U23500 (N_23500,N_18942,N_19961);
or U23501 (N_23501,N_17994,N_17842);
nand U23502 (N_23502,N_19846,N_17951);
nor U23503 (N_23503,N_16713,N_17356);
or U23504 (N_23504,N_17605,N_19087);
nand U23505 (N_23505,N_17125,N_16032);
xnor U23506 (N_23506,N_19002,N_19337);
or U23507 (N_23507,N_18629,N_17140);
nand U23508 (N_23508,N_18026,N_19562);
nand U23509 (N_23509,N_19534,N_15798);
nand U23510 (N_23510,N_15723,N_15286);
or U23511 (N_23511,N_19145,N_18782);
or U23512 (N_23512,N_17495,N_19623);
nand U23513 (N_23513,N_19259,N_17974);
xnor U23514 (N_23514,N_19182,N_15465);
xor U23515 (N_23515,N_18250,N_17959);
nand U23516 (N_23516,N_18584,N_15273);
xnor U23517 (N_23517,N_18717,N_18394);
or U23518 (N_23518,N_15219,N_15546);
nand U23519 (N_23519,N_19750,N_19536);
or U23520 (N_23520,N_16050,N_18375);
nor U23521 (N_23521,N_15128,N_16179);
nor U23522 (N_23522,N_18072,N_16177);
xor U23523 (N_23523,N_17692,N_16158);
or U23524 (N_23524,N_17199,N_16738);
nand U23525 (N_23525,N_16066,N_15992);
and U23526 (N_23526,N_19122,N_18949);
or U23527 (N_23527,N_19982,N_17081);
or U23528 (N_23528,N_15718,N_19011);
xnor U23529 (N_23529,N_16210,N_16655);
and U23530 (N_23530,N_16533,N_18156);
nor U23531 (N_23531,N_19131,N_15601);
nor U23532 (N_23532,N_17988,N_17774);
nand U23533 (N_23533,N_19163,N_18264);
nor U23534 (N_23534,N_19254,N_18618);
or U23535 (N_23535,N_19885,N_16286);
or U23536 (N_23536,N_16734,N_19495);
nor U23537 (N_23537,N_18880,N_19845);
or U23538 (N_23538,N_19377,N_16697);
xor U23539 (N_23539,N_17916,N_16889);
and U23540 (N_23540,N_18936,N_19658);
nor U23541 (N_23541,N_15262,N_19208);
xor U23542 (N_23542,N_15103,N_17117);
nor U23543 (N_23543,N_15849,N_16325);
nor U23544 (N_23544,N_15171,N_19058);
or U23545 (N_23545,N_17504,N_17286);
nor U23546 (N_23546,N_18939,N_17210);
xor U23547 (N_23547,N_18015,N_19555);
and U23548 (N_23548,N_16495,N_15281);
or U23549 (N_23549,N_15046,N_17827);
nand U23550 (N_23550,N_19145,N_18378);
xor U23551 (N_23551,N_17801,N_18805);
nor U23552 (N_23552,N_16499,N_15886);
nor U23553 (N_23553,N_17431,N_17734);
nor U23554 (N_23554,N_15632,N_18636);
nand U23555 (N_23555,N_17884,N_18131);
xor U23556 (N_23556,N_17582,N_17539);
and U23557 (N_23557,N_16435,N_19265);
xor U23558 (N_23558,N_16173,N_18031);
and U23559 (N_23559,N_16937,N_18220);
nand U23560 (N_23560,N_18330,N_19314);
xnor U23561 (N_23561,N_15027,N_16037);
nand U23562 (N_23562,N_16726,N_19809);
nand U23563 (N_23563,N_15995,N_15413);
or U23564 (N_23564,N_17200,N_18540);
nor U23565 (N_23565,N_16977,N_18343);
nand U23566 (N_23566,N_17467,N_15308);
xor U23567 (N_23567,N_17106,N_18841);
nand U23568 (N_23568,N_15239,N_15317);
and U23569 (N_23569,N_18644,N_19018);
and U23570 (N_23570,N_15039,N_15720);
and U23571 (N_23571,N_18106,N_18164);
xnor U23572 (N_23572,N_17750,N_16884);
nor U23573 (N_23573,N_15327,N_16014);
nand U23574 (N_23574,N_19306,N_17344);
or U23575 (N_23575,N_16272,N_17286);
nand U23576 (N_23576,N_18040,N_16486);
nand U23577 (N_23577,N_18888,N_15263);
and U23578 (N_23578,N_19366,N_17779);
and U23579 (N_23579,N_19574,N_16820);
or U23580 (N_23580,N_18589,N_16743);
xor U23581 (N_23581,N_19443,N_16636);
and U23582 (N_23582,N_18065,N_15208);
and U23583 (N_23583,N_15178,N_18769);
or U23584 (N_23584,N_17414,N_17311);
or U23585 (N_23585,N_18106,N_16240);
and U23586 (N_23586,N_15145,N_19513);
nor U23587 (N_23587,N_19458,N_18019);
xor U23588 (N_23588,N_19389,N_15034);
or U23589 (N_23589,N_17328,N_17819);
nand U23590 (N_23590,N_15613,N_19870);
nand U23591 (N_23591,N_16405,N_17143);
or U23592 (N_23592,N_17314,N_16315);
nor U23593 (N_23593,N_15582,N_15991);
and U23594 (N_23594,N_19450,N_18070);
nand U23595 (N_23595,N_15020,N_19412);
or U23596 (N_23596,N_15736,N_17693);
nand U23597 (N_23597,N_15862,N_15354);
nand U23598 (N_23598,N_16688,N_17596);
xnor U23599 (N_23599,N_17656,N_18195);
nor U23600 (N_23600,N_17840,N_16856);
nor U23601 (N_23601,N_15257,N_19994);
xnor U23602 (N_23602,N_18645,N_18204);
nand U23603 (N_23603,N_18028,N_18437);
nand U23604 (N_23604,N_18736,N_18108);
xor U23605 (N_23605,N_19742,N_16726);
nand U23606 (N_23606,N_15936,N_17995);
xnor U23607 (N_23607,N_17646,N_15424);
and U23608 (N_23608,N_16713,N_18346);
nand U23609 (N_23609,N_16733,N_15293);
xor U23610 (N_23610,N_18357,N_15533);
nand U23611 (N_23611,N_17316,N_15224);
and U23612 (N_23612,N_16526,N_18550);
xor U23613 (N_23613,N_16734,N_18169);
nor U23614 (N_23614,N_17501,N_16806);
xnor U23615 (N_23615,N_19002,N_19633);
xor U23616 (N_23616,N_16141,N_15864);
and U23617 (N_23617,N_18537,N_15279);
nand U23618 (N_23618,N_18026,N_18715);
xor U23619 (N_23619,N_15058,N_19789);
or U23620 (N_23620,N_17613,N_15726);
and U23621 (N_23621,N_17060,N_15810);
nand U23622 (N_23622,N_16590,N_17929);
or U23623 (N_23623,N_18888,N_18937);
xnor U23624 (N_23624,N_17509,N_19954);
and U23625 (N_23625,N_15972,N_17297);
xor U23626 (N_23626,N_16535,N_19892);
nand U23627 (N_23627,N_16424,N_17093);
nor U23628 (N_23628,N_19002,N_18950);
xor U23629 (N_23629,N_19650,N_15456);
nor U23630 (N_23630,N_16337,N_19518);
nor U23631 (N_23631,N_18453,N_15340);
or U23632 (N_23632,N_15486,N_17730);
nor U23633 (N_23633,N_15855,N_15652);
xor U23634 (N_23634,N_15897,N_15111);
nand U23635 (N_23635,N_16114,N_19917);
nor U23636 (N_23636,N_17425,N_15243);
and U23637 (N_23637,N_16722,N_16958);
and U23638 (N_23638,N_19448,N_15135);
xnor U23639 (N_23639,N_18194,N_16513);
nand U23640 (N_23640,N_15093,N_16019);
nor U23641 (N_23641,N_19223,N_18078);
xnor U23642 (N_23642,N_19445,N_16293);
nor U23643 (N_23643,N_18085,N_18159);
nor U23644 (N_23644,N_18106,N_17909);
or U23645 (N_23645,N_16834,N_17747);
nand U23646 (N_23646,N_17475,N_18742);
nand U23647 (N_23647,N_18370,N_15207);
and U23648 (N_23648,N_18288,N_15787);
nand U23649 (N_23649,N_19030,N_17136);
nor U23650 (N_23650,N_19761,N_15923);
nor U23651 (N_23651,N_18870,N_15725);
and U23652 (N_23652,N_17318,N_15785);
xor U23653 (N_23653,N_15030,N_16608);
and U23654 (N_23654,N_18156,N_17303);
nand U23655 (N_23655,N_15835,N_16441);
nand U23656 (N_23656,N_15319,N_15016);
or U23657 (N_23657,N_16560,N_18115);
xor U23658 (N_23658,N_17606,N_15593);
nor U23659 (N_23659,N_17785,N_17577);
or U23660 (N_23660,N_19083,N_15118);
xor U23661 (N_23661,N_15420,N_17581);
or U23662 (N_23662,N_18480,N_18412);
or U23663 (N_23663,N_18260,N_17895);
nand U23664 (N_23664,N_17134,N_15270);
and U23665 (N_23665,N_16041,N_18299);
and U23666 (N_23666,N_17707,N_19105);
xnor U23667 (N_23667,N_18252,N_19364);
or U23668 (N_23668,N_18578,N_15455);
and U23669 (N_23669,N_19161,N_19432);
nor U23670 (N_23670,N_16105,N_16218);
nand U23671 (N_23671,N_17988,N_18169);
nor U23672 (N_23672,N_17357,N_16592);
and U23673 (N_23673,N_19114,N_18260);
xnor U23674 (N_23674,N_15296,N_17084);
xnor U23675 (N_23675,N_18145,N_17322);
nand U23676 (N_23676,N_17596,N_17457);
and U23677 (N_23677,N_16102,N_17643);
nand U23678 (N_23678,N_15133,N_15564);
or U23679 (N_23679,N_16428,N_18711);
nand U23680 (N_23680,N_18606,N_16701);
or U23681 (N_23681,N_18464,N_18653);
xor U23682 (N_23682,N_16577,N_18947);
nor U23683 (N_23683,N_17722,N_19500);
and U23684 (N_23684,N_16917,N_17621);
xor U23685 (N_23685,N_19263,N_15199);
or U23686 (N_23686,N_15936,N_16688);
nor U23687 (N_23687,N_17283,N_19352);
xnor U23688 (N_23688,N_16246,N_16052);
xnor U23689 (N_23689,N_16412,N_17674);
and U23690 (N_23690,N_19870,N_16058);
and U23691 (N_23691,N_19311,N_18084);
and U23692 (N_23692,N_16318,N_19015);
nor U23693 (N_23693,N_17564,N_15768);
and U23694 (N_23694,N_19620,N_16834);
or U23695 (N_23695,N_18609,N_18097);
nor U23696 (N_23696,N_15632,N_17413);
xor U23697 (N_23697,N_16396,N_18004);
xnor U23698 (N_23698,N_16589,N_16198);
or U23699 (N_23699,N_17881,N_19126);
and U23700 (N_23700,N_16666,N_15671);
and U23701 (N_23701,N_18023,N_15150);
nand U23702 (N_23702,N_17223,N_19403);
nor U23703 (N_23703,N_15689,N_15559);
xnor U23704 (N_23704,N_15278,N_19185);
nand U23705 (N_23705,N_18656,N_17709);
xnor U23706 (N_23706,N_15952,N_17177);
and U23707 (N_23707,N_18879,N_19463);
nand U23708 (N_23708,N_18228,N_19156);
and U23709 (N_23709,N_16052,N_15553);
and U23710 (N_23710,N_15586,N_16339);
nor U23711 (N_23711,N_16087,N_17435);
or U23712 (N_23712,N_16763,N_17686);
and U23713 (N_23713,N_15509,N_18476);
nor U23714 (N_23714,N_17564,N_18974);
and U23715 (N_23715,N_17507,N_19675);
nand U23716 (N_23716,N_19894,N_16120);
xor U23717 (N_23717,N_17867,N_19275);
nand U23718 (N_23718,N_15672,N_19162);
xor U23719 (N_23719,N_15871,N_16083);
or U23720 (N_23720,N_17138,N_18557);
xor U23721 (N_23721,N_17651,N_19784);
nand U23722 (N_23722,N_16936,N_15327);
xor U23723 (N_23723,N_17170,N_15950);
and U23724 (N_23724,N_18115,N_15092);
xnor U23725 (N_23725,N_18995,N_17001);
or U23726 (N_23726,N_16495,N_19615);
and U23727 (N_23727,N_16203,N_15359);
nor U23728 (N_23728,N_17880,N_15742);
xnor U23729 (N_23729,N_16720,N_19131);
nor U23730 (N_23730,N_17214,N_18367);
xnor U23731 (N_23731,N_19409,N_19993);
xnor U23732 (N_23732,N_19898,N_17340);
nor U23733 (N_23733,N_15929,N_18490);
nor U23734 (N_23734,N_15045,N_19677);
or U23735 (N_23735,N_17372,N_15774);
nor U23736 (N_23736,N_15779,N_19191);
and U23737 (N_23737,N_18642,N_19016);
xor U23738 (N_23738,N_17556,N_17904);
nand U23739 (N_23739,N_16227,N_16425);
and U23740 (N_23740,N_17139,N_18169);
and U23741 (N_23741,N_17587,N_17853);
and U23742 (N_23742,N_16162,N_19501);
and U23743 (N_23743,N_18765,N_15866);
or U23744 (N_23744,N_15668,N_18128);
nand U23745 (N_23745,N_16350,N_18366);
nor U23746 (N_23746,N_16652,N_15036);
or U23747 (N_23747,N_16608,N_19900);
or U23748 (N_23748,N_18216,N_19965);
or U23749 (N_23749,N_15790,N_15730);
xnor U23750 (N_23750,N_19550,N_16768);
or U23751 (N_23751,N_18266,N_19189);
nand U23752 (N_23752,N_18769,N_16722);
nand U23753 (N_23753,N_18736,N_15003);
xnor U23754 (N_23754,N_18392,N_18133);
or U23755 (N_23755,N_15420,N_16159);
or U23756 (N_23756,N_19746,N_17765);
and U23757 (N_23757,N_15033,N_15497);
xnor U23758 (N_23758,N_17729,N_18800);
and U23759 (N_23759,N_17226,N_19898);
and U23760 (N_23760,N_17708,N_17996);
and U23761 (N_23761,N_17012,N_19260);
and U23762 (N_23762,N_15995,N_18459);
xor U23763 (N_23763,N_17117,N_16590);
and U23764 (N_23764,N_18560,N_16937);
and U23765 (N_23765,N_17638,N_15494);
nand U23766 (N_23766,N_15808,N_16314);
nand U23767 (N_23767,N_16271,N_17301);
nor U23768 (N_23768,N_19642,N_15710);
nand U23769 (N_23769,N_19511,N_17974);
xnor U23770 (N_23770,N_16772,N_19506);
nand U23771 (N_23771,N_18185,N_17515);
or U23772 (N_23772,N_17974,N_15154);
nor U23773 (N_23773,N_18608,N_19747);
or U23774 (N_23774,N_19360,N_15363);
nand U23775 (N_23775,N_17480,N_17158);
or U23776 (N_23776,N_19618,N_15557);
or U23777 (N_23777,N_16196,N_17648);
and U23778 (N_23778,N_19310,N_19046);
nor U23779 (N_23779,N_17186,N_15074);
xor U23780 (N_23780,N_15312,N_15984);
or U23781 (N_23781,N_17916,N_15309);
and U23782 (N_23782,N_16958,N_18664);
nand U23783 (N_23783,N_16099,N_17703);
nand U23784 (N_23784,N_18615,N_16651);
and U23785 (N_23785,N_16583,N_19253);
nor U23786 (N_23786,N_19280,N_16278);
and U23787 (N_23787,N_15500,N_16185);
nor U23788 (N_23788,N_16864,N_18061);
and U23789 (N_23789,N_15392,N_16062);
or U23790 (N_23790,N_17450,N_18277);
and U23791 (N_23791,N_18601,N_16975);
nand U23792 (N_23792,N_17733,N_18662);
nand U23793 (N_23793,N_19133,N_19765);
or U23794 (N_23794,N_17154,N_19724);
nor U23795 (N_23795,N_15720,N_15748);
nor U23796 (N_23796,N_16478,N_19766);
xnor U23797 (N_23797,N_17853,N_19852);
nor U23798 (N_23798,N_16915,N_18005);
or U23799 (N_23799,N_15661,N_18794);
nor U23800 (N_23800,N_16964,N_17226);
nor U23801 (N_23801,N_16799,N_19207);
nor U23802 (N_23802,N_19345,N_15348);
or U23803 (N_23803,N_17223,N_17927);
and U23804 (N_23804,N_17545,N_19748);
or U23805 (N_23805,N_16550,N_18094);
or U23806 (N_23806,N_17611,N_16179);
xnor U23807 (N_23807,N_17640,N_16074);
or U23808 (N_23808,N_18683,N_15977);
nor U23809 (N_23809,N_15881,N_17064);
and U23810 (N_23810,N_16776,N_17843);
and U23811 (N_23811,N_16157,N_16937);
xor U23812 (N_23812,N_17577,N_19102);
nor U23813 (N_23813,N_15667,N_15044);
nor U23814 (N_23814,N_15390,N_16029);
nor U23815 (N_23815,N_18645,N_16259);
xnor U23816 (N_23816,N_16118,N_16772);
xor U23817 (N_23817,N_18090,N_16027);
xor U23818 (N_23818,N_17932,N_17004);
nor U23819 (N_23819,N_17924,N_19717);
nand U23820 (N_23820,N_17526,N_15504);
nor U23821 (N_23821,N_15889,N_15605);
and U23822 (N_23822,N_18145,N_17553);
or U23823 (N_23823,N_16379,N_19997);
nand U23824 (N_23824,N_16883,N_16882);
nand U23825 (N_23825,N_15640,N_16630);
or U23826 (N_23826,N_18673,N_19571);
or U23827 (N_23827,N_16509,N_15343);
xor U23828 (N_23828,N_16925,N_19999);
xor U23829 (N_23829,N_16885,N_16065);
or U23830 (N_23830,N_17548,N_19684);
and U23831 (N_23831,N_15619,N_19099);
or U23832 (N_23832,N_19284,N_15991);
nand U23833 (N_23833,N_18947,N_17736);
or U23834 (N_23834,N_17398,N_18383);
nor U23835 (N_23835,N_19707,N_17764);
xor U23836 (N_23836,N_18963,N_18065);
xor U23837 (N_23837,N_18444,N_17066);
or U23838 (N_23838,N_16061,N_16823);
or U23839 (N_23839,N_18467,N_15674);
and U23840 (N_23840,N_16008,N_15608);
xor U23841 (N_23841,N_19968,N_16319);
nand U23842 (N_23842,N_17461,N_17269);
or U23843 (N_23843,N_19557,N_15619);
xnor U23844 (N_23844,N_17262,N_19205);
or U23845 (N_23845,N_18584,N_16020);
nor U23846 (N_23846,N_16725,N_19609);
nand U23847 (N_23847,N_15352,N_18825);
nand U23848 (N_23848,N_17527,N_18383);
xor U23849 (N_23849,N_18819,N_19654);
nand U23850 (N_23850,N_18470,N_19681);
nand U23851 (N_23851,N_16358,N_16156);
xnor U23852 (N_23852,N_16556,N_15051);
nand U23853 (N_23853,N_15335,N_18000);
or U23854 (N_23854,N_15498,N_19758);
nor U23855 (N_23855,N_16361,N_18991);
and U23856 (N_23856,N_17054,N_17788);
nor U23857 (N_23857,N_18697,N_15709);
or U23858 (N_23858,N_16849,N_17822);
xor U23859 (N_23859,N_18076,N_18541);
xor U23860 (N_23860,N_18328,N_15397);
and U23861 (N_23861,N_15189,N_17823);
xnor U23862 (N_23862,N_15706,N_15289);
nand U23863 (N_23863,N_17278,N_15482);
nand U23864 (N_23864,N_15980,N_17172);
or U23865 (N_23865,N_16096,N_17864);
nand U23866 (N_23866,N_18370,N_18076);
xnor U23867 (N_23867,N_15398,N_16338);
xnor U23868 (N_23868,N_18340,N_18055);
and U23869 (N_23869,N_18911,N_17378);
xnor U23870 (N_23870,N_17279,N_19744);
xnor U23871 (N_23871,N_16780,N_19560);
or U23872 (N_23872,N_19552,N_17494);
nand U23873 (N_23873,N_19082,N_19609);
and U23874 (N_23874,N_16067,N_17990);
or U23875 (N_23875,N_18255,N_16795);
nor U23876 (N_23876,N_16177,N_15860);
xor U23877 (N_23877,N_17423,N_17958);
and U23878 (N_23878,N_15818,N_17830);
xor U23879 (N_23879,N_18304,N_19212);
or U23880 (N_23880,N_17950,N_15913);
nand U23881 (N_23881,N_18616,N_19430);
nand U23882 (N_23882,N_15726,N_15617);
nor U23883 (N_23883,N_18568,N_15736);
nor U23884 (N_23884,N_18873,N_15465);
nor U23885 (N_23885,N_17732,N_16011);
nor U23886 (N_23886,N_19522,N_15999);
xor U23887 (N_23887,N_18125,N_16366);
and U23888 (N_23888,N_16548,N_16761);
nor U23889 (N_23889,N_16991,N_16535);
or U23890 (N_23890,N_19624,N_16706);
and U23891 (N_23891,N_15367,N_17338);
nor U23892 (N_23892,N_16343,N_15986);
xnor U23893 (N_23893,N_18079,N_19579);
nor U23894 (N_23894,N_19880,N_19499);
nand U23895 (N_23895,N_16714,N_19890);
nor U23896 (N_23896,N_19416,N_15123);
nor U23897 (N_23897,N_17448,N_18137);
nor U23898 (N_23898,N_19028,N_17781);
and U23899 (N_23899,N_19871,N_17537);
nor U23900 (N_23900,N_17641,N_17176);
xnor U23901 (N_23901,N_17521,N_15470);
nand U23902 (N_23902,N_18506,N_17626);
or U23903 (N_23903,N_19870,N_16378);
or U23904 (N_23904,N_16062,N_15326);
nand U23905 (N_23905,N_17363,N_17136);
or U23906 (N_23906,N_16385,N_19848);
nand U23907 (N_23907,N_15569,N_17230);
and U23908 (N_23908,N_16967,N_17611);
xnor U23909 (N_23909,N_19496,N_15168);
or U23910 (N_23910,N_16554,N_17403);
nor U23911 (N_23911,N_15540,N_15911);
xor U23912 (N_23912,N_19904,N_18999);
or U23913 (N_23913,N_15190,N_15544);
nand U23914 (N_23914,N_18427,N_15476);
nor U23915 (N_23915,N_17309,N_17939);
or U23916 (N_23916,N_16657,N_15154);
xor U23917 (N_23917,N_19020,N_17893);
nor U23918 (N_23918,N_19447,N_17976);
nand U23919 (N_23919,N_17709,N_18505);
and U23920 (N_23920,N_16498,N_17067);
nand U23921 (N_23921,N_17920,N_16206);
and U23922 (N_23922,N_18061,N_19450);
and U23923 (N_23923,N_16923,N_18349);
nand U23924 (N_23924,N_16442,N_16718);
nand U23925 (N_23925,N_17091,N_18008);
xnor U23926 (N_23926,N_16392,N_15470);
xor U23927 (N_23927,N_16297,N_16525);
and U23928 (N_23928,N_18825,N_15069);
nor U23929 (N_23929,N_17293,N_18836);
nor U23930 (N_23930,N_19816,N_17050);
and U23931 (N_23931,N_16855,N_19210);
nand U23932 (N_23932,N_16197,N_15893);
nor U23933 (N_23933,N_17934,N_19501);
xor U23934 (N_23934,N_16854,N_16446);
nand U23935 (N_23935,N_16969,N_15970);
or U23936 (N_23936,N_15145,N_17722);
nand U23937 (N_23937,N_16078,N_17696);
or U23938 (N_23938,N_19685,N_17606);
nand U23939 (N_23939,N_18625,N_15856);
and U23940 (N_23940,N_18526,N_17935);
xnor U23941 (N_23941,N_15451,N_15141);
and U23942 (N_23942,N_15121,N_19733);
nand U23943 (N_23943,N_15532,N_16283);
and U23944 (N_23944,N_15238,N_16704);
nor U23945 (N_23945,N_17546,N_19333);
and U23946 (N_23946,N_15251,N_18520);
xnor U23947 (N_23947,N_18790,N_17089);
or U23948 (N_23948,N_15112,N_16299);
and U23949 (N_23949,N_16922,N_19735);
or U23950 (N_23950,N_17658,N_16864);
and U23951 (N_23951,N_17724,N_19081);
and U23952 (N_23952,N_17908,N_16855);
or U23953 (N_23953,N_18065,N_16802);
or U23954 (N_23954,N_15079,N_16779);
nor U23955 (N_23955,N_18380,N_18895);
or U23956 (N_23956,N_16704,N_18228);
xor U23957 (N_23957,N_19485,N_17714);
nor U23958 (N_23958,N_16863,N_18655);
xor U23959 (N_23959,N_19366,N_16135);
and U23960 (N_23960,N_16444,N_17670);
nor U23961 (N_23961,N_16483,N_16738);
nor U23962 (N_23962,N_16649,N_18716);
and U23963 (N_23963,N_19254,N_17453);
nand U23964 (N_23964,N_15972,N_16203);
and U23965 (N_23965,N_19875,N_15530);
nor U23966 (N_23966,N_17483,N_17808);
nor U23967 (N_23967,N_18003,N_18475);
nor U23968 (N_23968,N_16207,N_16741);
nor U23969 (N_23969,N_19980,N_16819);
xor U23970 (N_23970,N_18828,N_17876);
nor U23971 (N_23971,N_15188,N_18954);
and U23972 (N_23972,N_19902,N_18146);
nor U23973 (N_23973,N_15038,N_18605);
and U23974 (N_23974,N_19225,N_19133);
nand U23975 (N_23975,N_17771,N_18560);
or U23976 (N_23976,N_16122,N_19858);
or U23977 (N_23977,N_19966,N_19322);
nor U23978 (N_23978,N_16162,N_18831);
nor U23979 (N_23979,N_19334,N_18105);
or U23980 (N_23980,N_15194,N_16447);
nand U23981 (N_23981,N_17904,N_15452);
and U23982 (N_23982,N_19050,N_16365);
xnor U23983 (N_23983,N_18521,N_17471);
nand U23984 (N_23984,N_19567,N_16438);
and U23985 (N_23985,N_15221,N_15733);
xor U23986 (N_23986,N_18459,N_15658);
xnor U23987 (N_23987,N_19655,N_17494);
xor U23988 (N_23988,N_19759,N_15099);
and U23989 (N_23989,N_15740,N_15465);
xor U23990 (N_23990,N_15321,N_17214);
xor U23991 (N_23991,N_16781,N_19606);
xnor U23992 (N_23992,N_16119,N_17293);
and U23993 (N_23993,N_19239,N_15621);
nor U23994 (N_23994,N_17888,N_15271);
or U23995 (N_23995,N_17837,N_18713);
nand U23996 (N_23996,N_18774,N_19898);
nand U23997 (N_23997,N_15974,N_18743);
nand U23998 (N_23998,N_16268,N_17188);
and U23999 (N_23999,N_19810,N_19874);
or U24000 (N_24000,N_18062,N_15322);
nand U24001 (N_24001,N_19622,N_18676);
nand U24002 (N_24002,N_16106,N_17333);
nand U24003 (N_24003,N_17137,N_17737);
nor U24004 (N_24004,N_17741,N_16785);
nor U24005 (N_24005,N_15711,N_18344);
and U24006 (N_24006,N_18993,N_19343);
or U24007 (N_24007,N_16988,N_18189);
nand U24008 (N_24008,N_16368,N_17637);
or U24009 (N_24009,N_19174,N_17821);
xor U24010 (N_24010,N_19998,N_16774);
nor U24011 (N_24011,N_15364,N_18405);
or U24012 (N_24012,N_15595,N_15501);
xnor U24013 (N_24013,N_16318,N_19810);
nor U24014 (N_24014,N_16753,N_19121);
and U24015 (N_24015,N_18564,N_17857);
or U24016 (N_24016,N_15276,N_17937);
or U24017 (N_24017,N_18433,N_19934);
and U24018 (N_24018,N_16532,N_18580);
nand U24019 (N_24019,N_16882,N_15408);
and U24020 (N_24020,N_19695,N_16771);
nor U24021 (N_24021,N_15569,N_19167);
or U24022 (N_24022,N_15171,N_16287);
xnor U24023 (N_24023,N_16753,N_17391);
nor U24024 (N_24024,N_17519,N_17743);
xnor U24025 (N_24025,N_19007,N_18932);
or U24026 (N_24026,N_17641,N_16768);
xnor U24027 (N_24027,N_16760,N_18881);
xor U24028 (N_24028,N_16071,N_16863);
or U24029 (N_24029,N_18141,N_18843);
nor U24030 (N_24030,N_15216,N_19457);
nand U24031 (N_24031,N_18039,N_17780);
xor U24032 (N_24032,N_19548,N_16381);
and U24033 (N_24033,N_19822,N_17651);
xnor U24034 (N_24034,N_19023,N_19282);
nor U24035 (N_24035,N_19290,N_16963);
nor U24036 (N_24036,N_15294,N_19525);
and U24037 (N_24037,N_17555,N_19027);
and U24038 (N_24038,N_18232,N_19011);
or U24039 (N_24039,N_16571,N_15023);
xor U24040 (N_24040,N_19902,N_17111);
xor U24041 (N_24041,N_16931,N_18873);
and U24042 (N_24042,N_17368,N_16169);
xor U24043 (N_24043,N_18254,N_19638);
or U24044 (N_24044,N_15956,N_18982);
nand U24045 (N_24045,N_18018,N_18767);
nand U24046 (N_24046,N_19738,N_19050);
xor U24047 (N_24047,N_15212,N_16310);
or U24048 (N_24048,N_19233,N_16894);
xor U24049 (N_24049,N_17995,N_17925);
and U24050 (N_24050,N_19211,N_19207);
and U24051 (N_24051,N_15216,N_16076);
nor U24052 (N_24052,N_17867,N_18744);
or U24053 (N_24053,N_16734,N_18432);
nor U24054 (N_24054,N_15608,N_17267);
xor U24055 (N_24055,N_19754,N_17590);
nand U24056 (N_24056,N_15555,N_17807);
xnor U24057 (N_24057,N_15950,N_19984);
or U24058 (N_24058,N_17979,N_17025);
nor U24059 (N_24059,N_19454,N_19622);
and U24060 (N_24060,N_16297,N_18408);
nand U24061 (N_24061,N_15291,N_16228);
xor U24062 (N_24062,N_17531,N_16005);
nand U24063 (N_24063,N_16814,N_15098);
and U24064 (N_24064,N_18216,N_15536);
nand U24065 (N_24065,N_15571,N_17607);
and U24066 (N_24066,N_15057,N_16158);
nand U24067 (N_24067,N_19436,N_19732);
nand U24068 (N_24068,N_18690,N_16513);
or U24069 (N_24069,N_18263,N_15560);
nor U24070 (N_24070,N_18735,N_16228);
nor U24071 (N_24071,N_19912,N_17214);
nor U24072 (N_24072,N_19147,N_15459);
nand U24073 (N_24073,N_19556,N_17924);
nor U24074 (N_24074,N_17325,N_15844);
and U24075 (N_24075,N_15543,N_17445);
nand U24076 (N_24076,N_17261,N_17935);
nand U24077 (N_24077,N_19785,N_16771);
or U24078 (N_24078,N_18094,N_19402);
and U24079 (N_24079,N_17721,N_16505);
and U24080 (N_24080,N_15311,N_15497);
nor U24081 (N_24081,N_18497,N_18472);
nor U24082 (N_24082,N_19436,N_15765);
or U24083 (N_24083,N_16081,N_18934);
nor U24084 (N_24084,N_16159,N_19561);
nor U24085 (N_24085,N_16416,N_19139);
nand U24086 (N_24086,N_17218,N_18513);
nor U24087 (N_24087,N_16581,N_16637);
or U24088 (N_24088,N_18676,N_16849);
nor U24089 (N_24089,N_17864,N_16936);
or U24090 (N_24090,N_19094,N_16518);
or U24091 (N_24091,N_17737,N_16535);
and U24092 (N_24092,N_18167,N_15187);
xnor U24093 (N_24093,N_16708,N_19756);
nand U24094 (N_24094,N_18250,N_17929);
or U24095 (N_24095,N_19499,N_17598);
nand U24096 (N_24096,N_18720,N_17702);
xor U24097 (N_24097,N_17884,N_15959);
or U24098 (N_24098,N_18827,N_18493);
and U24099 (N_24099,N_18723,N_17017);
and U24100 (N_24100,N_19064,N_16813);
nor U24101 (N_24101,N_17011,N_18832);
nor U24102 (N_24102,N_15731,N_16799);
or U24103 (N_24103,N_18816,N_17081);
xor U24104 (N_24104,N_15562,N_19940);
nand U24105 (N_24105,N_16068,N_18754);
nand U24106 (N_24106,N_18465,N_16059);
or U24107 (N_24107,N_15990,N_17505);
or U24108 (N_24108,N_16728,N_19894);
nor U24109 (N_24109,N_18825,N_19513);
nor U24110 (N_24110,N_17018,N_17903);
xnor U24111 (N_24111,N_16686,N_18134);
xor U24112 (N_24112,N_17475,N_15701);
nand U24113 (N_24113,N_17036,N_18203);
nor U24114 (N_24114,N_18092,N_17898);
and U24115 (N_24115,N_16132,N_16721);
or U24116 (N_24116,N_17351,N_19499);
and U24117 (N_24117,N_19518,N_16904);
nand U24118 (N_24118,N_18570,N_18014);
xnor U24119 (N_24119,N_17684,N_19320);
xor U24120 (N_24120,N_19803,N_16681);
nand U24121 (N_24121,N_15927,N_17999);
nand U24122 (N_24122,N_19965,N_18494);
or U24123 (N_24123,N_18757,N_18432);
nand U24124 (N_24124,N_17871,N_16344);
nor U24125 (N_24125,N_15083,N_16811);
and U24126 (N_24126,N_15349,N_17325);
xnor U24127 (N_24127,N_16200,N_18487);
nor U24128 (N_24128,N_18283,N_15967);
or U24129 (N_24129,N_17420,N_18504);
and U24130 (N_24130,N_18035,N_17127);
or U24131 (N_24131,N_15824,N_16589);
nor U24132 (N_24132,N_19835,N_17597);
or U24133 (N_24133,N_19087,N_18668);
nor U24134 (N_24134,N_19327,N_17575);
nand U24135 (N_24135,N_18147,N_18794);
nand U24136 (N_24136,N_18318,N_19940);
nand U24137 (N_24137,N_17827,N_19303);
xor U24138 (N_24138,N_15329,N_19660);
nand U24139 (N_24139,N_18307,N_17881);
xor U24140 (N_24140,N_18276,N_19776);
nand U24141 (N_24141,N_15022,N_19038);
and U24142 (N_24142,N_19805,N_18672);
and U24143 (N_24143,N_15524,N_19623);
nor U24144 (N_24144,N_15180,N_16526);
and U24145 (N_24145,N_19517,N_18394);
and U24146 (N_24146,N_16330,N_18601);
nand U24147 (N_24147,N_16264,N_15130);
nor U24148 (N_24148,N_18049,N_18918);
or U24149 (N_24149,N_15680,N_15500);
xnor U24150 (N_24150,N_16409,N_17815);
nor U24151 (N_24151,N_18709,N_18849);
xor U24152 (N_24152,N_19348,N_19652);
nor U24153 (N_24153,N_15325,N_18661);
and U24154 (N_24154,N_17812,N_15023);
xor U24155 (N_24155,N_15052,N_15192);
or U24156 (N_24156,N_15434,N_17931);
nand U24157 (N_24157,N_15956,N_16506);
xor U24158 (N_24158,N_17672,N_16125);
xnor U24159 (N_24159,N_18569,N_16304);
nor U24160 (N_24160,N_17233,N_16909);
and U24161 (N_24161,N_15352,N_17682);
xnor U24162 (N_24162,N_16354,N_18843);
xnor U24163 (N_24163,N_16231,N_17407);
or U24164 (N_24164,N_18154,N_16213);
nand U24165 (N_24165,N_17519,N_15584);
nor U24166 (N_24166,N_18471,N_17489);
or U24167 (N_24167,N_15219,N_17187);
xnor U24168 (N_24168,N_15087,N_17793);
nor U24169 (N_24169,N_15350,N_16023);
or U24170 (N_24170,N_16727,N_19434);
nor U24171 (N_24171,N_19078,N_19251);
xor U24172 (N_24172,N_18829,N_16303);
xor U24173 (N_24173,N_15474,N_18289);
or U24174 (N_24174,N_18625,N_16067);
and U24175 (N_24175,N_18379,N_18012);
xor U24176 (N_24176,N_15708,N_15207);
and U24177 (N_24177,N_18838,N_16868);
nand U24178 (N_24178,N_17026,N_19791);
nand U24179 (N_24179,N_15789,N_18137);
xor U24180 (N_24180,N_15083,N_15984);
nor U24181 (N_24181,N_15932,N_18176);
xor U24182 (N_24182,N_16630,N_18470);
and U24183 (N_24183,N_19017,N_19401);
or U24184 (N_24184,N_18902,N_15020);
nor U24185 (N_24185,N_18544,N_18376);
and U24186 (N_24186,N_17007,N_17103);
nor U24187 (N_24187,N_17063,N_17070);
xor U24188 (N_24188,N_18511,N_18364);
xor U24189 (N_24189,N_15568,N_19250);
nand U24190 (N_24190,N_17357,N_16007);
nand U24191 (N_24191,N_15416,N_16432);
nand U24192 (N_24192,N_18349,N_19060);
nor U24193 (N_24193,N_19243,N_15714);
xnor U24194 (N_24194,N_17292,N_16732);
nand U24195 (N_24195,N_18207,N_19529);
xnor U24196 (N_24196,N_16321,N_17917);
xnor U24197 (N_24197,N_15893,N_16905);
xnor U24198 (N_24198,N_16048,N_17731);
xnor U24199 (N_24199,N_15029,N_19854);
nor U24200 (N_24200,N_18078,N_17159);
xnor U24201 (N_24201,N_16666,N_15916);
xor U24202 (N_24202,N_15932,N_17249);
nand U24203 (N_24203,N_17272,N_15033);
nor U24204 (N_24204,N_16811,N_19253);
nand U24205 (N_24205,N_16123,N_18617);
xor U24206 (N_24206,N_17946,N_19539);
nor U24207 (N_24207,N_19067,N_18395);
nor U24208 (N_24208,N_19990,N_16247);
nor U24209 (N_24209,N_17304,N_15608);
and U24210 (N_24210,N_17687,N_18842);
or U24211 (N_24211,N_15213,N_17764);
and U24212 (N_24212,N_18566,N_19391);
xnor U24213 (N_24213,N_19284,N_19097);
and U24214 (N_24214,N_18887,N_19793);
xor U24215 (N_24215,N_18965,N_19641);
xor U24216 (N_24216,N_16519,N_15521);
xor U24217 (N_24217,N_16082,N_19844);
and U24218 (N_24218,N_19634,N_15176);
nand U24219 (N_24219,N_19920,N_15562);
and U24220 (N_24220,N_18202,N_15361);
and U24221 (N_24221,N_17535,N_19764);
xnor U24222 (N_24222,N_19932,N_19059);
nand U24223 (N_24223,N_15504,N_17818);
nor U24224 (N_24224,N_15000,N_19825);
or U24225 (N_24225,N_17249,N_17796);
nand U24226 (N_24226,N_18537,N_16261);
or U24227 (N_24227,N_17384,N_15549);
xnor U24228 (N_24228,N_15238,N_15267);
and U24229 (N_24229,N_18643,N_17117);
and U24230 (N_24230,N_18863,N_18043);
and U24231 (N_24231,N_16712,N_16488);
nor U24232 (N_24232,N_18357,N_18324);
nor U24233 (N_24233,N_15776,N_18645);
nand U24234 (N_24234,N_16945,N_16788);
nand U24235 (N_24235,N_19314,N_19060);
xnor U24236 (N_24236,N_17252,N_19961);
nand U24237 (N_24237,N_17702,N_15132);
nor U24238 (N_24238,N_16336,N_18373);
and U24239 (N_24239,N_17320,N_19584);
nand U24240 (N_24240,N_17481,N_17180);
or U24241 (N_24241,N_18764,N_19866);
nand U24242 (N_24242,N_18822,N_17949);
nor U24243 (N_24243,N_17896,N_18114);
nand U24244 (N_24244,N_18447,N_18076);
and U24245 (N_24245,N_17786,N_15763);
and U24246 (N_24246,N_18037,N_17272);
or U24247 (N_24247,N_18985,N_16187);
nand U24248 (N_24248,N_16390,N_17453);
or U24249 (N_24249,N_17256,N_15827);
nor U24250 (N_24250,N_18767,N_15882);
xnor U24251 (N_24251,N_17844,N_18777);
nand U24252 (N_24252,N_17800,N_19151);
nand U24253 (N_24253,N_18818,N_19611);
and U24254 (N_24254,N_19423,N_15723);
or U24255 (N_24255,N_18534,N_18041);
and U24256 (N_24256,N_19641,N_18417);
and U24257 (N_24257,N_19102,N_15371);
nor U24258 (N_24258,N_15057,N_15432);
or U24259 (N_24259,N_19693,N_18117);
or U24260 (N_24260,N_15261,N_19638);
and U24261 (N_24261,N_16706,N_15453);
nor U24262 (N_24262,N_15649,N_19888);
xnor U24263 (N_24263,N_18536,N_17740);
and U24264 (N_24264,N_16580,N_17206);
nor U24265 (N_24265,N_17043,N_17127);
or U24266 (N_24266,N_17905,N_17705);
or U24267 (N_24267,N_15654,N_19106);
or U24268 (N_24268,N_15437,N_18252);
nand U24269 (N_24269,N_17813,N_18897);
or U24270 (N_24270,N_15316,N_18153);
or U24271 (N_24271,N_19908,N_19848);
xnor U24272 (N_24272,N_19186,N_17997);
nand U24273 (N_24273,N_17514,N_18819);
nor U24274 (N_24274,N_18488,N_17091);
xor U24275 (N_24275,N_15793,N_19084);
or U24276 (N_24276,N_16398,N_15234);
and U24277 (N_24277,N_16342,N_17607);
and U24278 (N_24278,N_16459,N_19943);
xor U24279 (N_24279,N_16591,N_17125);
and U24280 (N_24280,N_18744,N_19885);
nor U24281 (N_24281,N_15996,N_18459);
xor U24282 (N_24282,N_16102,N_17857);
xnor U24283 (N_24283,N_15885,N_18185);
or U24284 (N_24284,N_15574,N_16550);
nand U24285 (N_24285,N_16039,N_15893);
nor U24286 (N_24286,N_19187,N_16969);
or U24287 (N_24287,N_15592,N_16188);
or U24288 (N_24288,N_15402,N_17564);
or U24289 (N_24289,N_18313,N_19735);
or U24290 (N_24290,N_18994,N_17029);
nand U24291 (N_24291,N_19056,N_15656);
nor U24292 (N_24292,N_19396,N_17146);
or U24293 (N_24293,N_19756,N_17014);
nor U24294 (N_24294,N_17162,N_19449);
xor U24295 (N_24295,N_15487,N_18603);
and U24296 (N_24296,N_18943,N_17156);
nand U24297 (N_24297,N_15654,N_19770);
nand U24298 (N_24298,N_18770,N_18059);
xnor U24299 (N_24299,N_17944,N_18869);
nor U24300 (N_24300,N_15981,N_15273);
xnor U24301 (N_24301,N_19393,N_15512);
nand U24302 (N_24302,N_15721,N_16723);
and U24303 (N_24303,N_17248,N_19992);
and U24304 (N_24304,N_19308,N_18859);
or U24305 (N_24305,N_16035,N_15412);
nor U24306 (N_24306,N_15133,N_19334);
and U24307 (N_24307,N_19875,N_18489);
and U24308 (N_24308,N_19727,N_16938);
xnor U24309 (N_24309,N_18204,N_19264);
nor U24310 (N_24310,N_16522,N_18929);
xor U24311 (N_24311,N_15338,N_19536);
xor U24312 (N_24312,N_19596,N_17973);
xnor U24313 (N_24313,N_16359,N_16130);
nand U24314 (N_24314,N_16044,N_16577);
nand U24315 (N_24315,N_17943,N_18509);
xor U24316 (N_24316,N_19627,N_15880);
nand U24317 (N_24317,N_16714,N_15796);
and U24318 (N_24318,N_17006,N_15938);
xnor U24319 (N_24319,N_18210,N_18959);
or U24320 (N_24320,N_19770,N_19993);
and U24321 (N_24321,N_18460,N_18306);
and U24322 (N_24322,N_16143,N_15250);
or U24323 (N_24323,N_15625,N_16992);
nor U24324 (N_24324,N_16425,N_16303);
nor U24325 (N_24325,N_15487,N_15606);
and U24326 (N_24326,N_16977,N_15190);
and U24327 (N_24327,N_19793,N_19262);
xnor U24328 (N_24328,N_16154,N_17165);
xor U24329 (N_24329,N_19825,N_15021);
and U24330 (N_24330,N_18324,N_18018);
nand U24331 (N_24331,N_16233,N_17721);
nor U24332 (N_24332,N_17633,N_15757);
and U24333 (N_24333,N_16640,N_17988);
xor U24334 (N_24334,N_17268,N_17322);
and U24335 (N_24335,N_16489,N_16957);
nor U24336 (N_24336,N_17966,N_15533);
and U24337 (N_24337,N_18084,N_19659);
xor U24338 (N_24338,N_17014,N_16562);
or U24339 (N_24339,N_15831,N_18730);
or U24340 (N_24340,N_15525,N_16037);
xnor U24341 (N_24341,N_16459,N_16958);
xnor U24342 (N_24342,N_17175,N_15618);
nand U24343 (N_24343,N_15138,N_18541);
xor U24344 (N_24344,N_18083,N_15989);
nor U24345 (N_24345,N_17987,N_19865);
and U24346 (N_24346,N_17679,N_16522);
xor U24347 (N_24347,N_15377,N_18454);
xor U24348 (N_24348,N_19732,N_17868);
or U24349 (N_24349,N_19707,N_15215);
nand U24350 (N_24350,N_17255,N_17911);
xor U24351 (N_24351,N_15354,N_18390);
xor U24352 (N_24352,N_18366,N_18682);
xor U24353 (N_24353,N_15712,N_16592);
or U24354 (N_24354,N_19601,N_18123);
or U24355 (N_24355,N_18651,N_19323);
or U24356 (N_24356,N_19293,N_15322);
nor U24357 (N_24357,N_18021,N_17680);
nand U24358 (N_24358,N_19695,N_16039);
xnor U24359 (N_24359,N_19531,N_16719);
and U24360 (N_24360,N_16185,N_16059);
and U24361 (N_24361,N_19052,N_15784);
xor U24362 (N_24362,N_19486,N_17118);
xor U24363 (N_24363,N_16403,N_17054);
nor U24364 (N_24364,N_18608,N_17226);
xor U24365 (N_24365,N_18555,N_19595);
xnor U24366 (N_24366,N_15148,N_16517);
nand U24367 (N_24367,N_18530,N_15181);
or U24368 (N_24368,N_19187,N_15952);
nand U24369 (N_24369,N_17082,N_17880);
and U24370 (N_24370,N_18463,N_17742);
and U24371 (N_24371,N_18234,N_18445);
or U24372 (N_24372,N_16910,N_15388);
or U24373 (N_24373,N_15181,N_16024);
nand U24374 (N_24374,N_18798,N_17078);
nand U24375 (N_24375,N_16017,N_17052);
nand U24376 (N_24376,N_17026,N_19561);
nand U24377 (N_24377,N_19726,N_15521);
xor U24378 (N_24378,N_15189,N_16092);
xor U24379 (N_24379,N_18629,N_19716);
nand U24380 (N_24380,N_15523,N_18248);
nor U24381 (N_24381,N_15822,N_17979);
xor U24382 (N_24382,N_15715,N_15077);
nor U24383 (N_24383,N_19844,N_18222);
nor U24384 (N_24384,N_16014,N_17914);
nor U24385 (N_24385,N_19709,N_18026);
and U24386 (N_24386,N_16603,N_19075);
nand U24387 (N_24387,N_15270,N_19497);
and U24388 (N_24388,N_18690,N_15026);
nor U24389 (N_24389,N_19196,N_18374);
xor U24390 (N_24390,N_15963,N_17568);
nand U24391 (N_24391,N_16030,N_16660);
and U24392 (N_24392,N_15106,N_19405);
xor U24393 (N_24393,N_15102,N_18516);
xor U24394 (N_24394,N_16440,N_17534);
xor U24395 (N_24395,N_19024,N_18137);
nor U24396 (N_24396,N_18000,N_16112);
xnor U24397 (N_24397,N_17671,N_19986);
nor U24398 (N_24398,N_16907,N_19489);
and U24399 (N_24399,N_17504,N_19568);
and U24400 (N_24400,N_19905,N_18499);
xnor U24401 (N_24401,N_16747,N_19459);
nand U24402 (N_24402,N_16316,N_17631);
nand U24403 (N_24403,N_17535,N_17613);
and U24404 (N_24404,N_19052,N_18785);
or U24405 (N_24405,N_17342,N_16097);
xnor U24406 (N_24406,N_18662,N_17289);
nand U24407 (N_24407,N_15843,N_18473);
or U24408 (N_24408,N_19318,N_19586);
xor U24409 (N_24409,N_18458,N_16586);
nand U24410 (N_24410,N_16057,N_19639);
and U24411 (N_24411,N_15767,N_16941);
xnor U24412 (N_24412,N_17742,N_19514);
nor U24413 (N_24413,N_15409,N_16046);
xnor U24414 (N_24414,N_16114,N_18529);
nand U24415 (N_24415,N_19181,N_16409);
xor U24416 (N_24416,N_16337,N_15498);
nand U24417 (N_24417,N_15672,N_16899);
and U24418 (N_24418,N_15403,N_17034);
or U24419 (N_24419,N_17194,N_19798);
nand U24420 (N_24420,N_15119,N_16331);
xnor U24421 (N_24421,N_19752,N_15385);
and U24422 (N_24422,N_16472,N_16661);
nor U24423 (N_24423,N_15465,N_15702);
or U24424 (N_24424,N_19091,N_17168);
xor U24425 (N_24425,N_18892,N_16131);
xor U24426 (N_24426,N_18931,N_18435);
or U24427 (N_24427,N_16918,N_17172);
xnor U24428 (N_24428,N_18735,N_16707);
nor U24429 (N_24429,N_19919,N_18263);
or U24430 (N_24430,N_17795,N_15759);
and U24431 (N_24431,N_16056,N_16570);
and U24432 (N_24432,N_17804,N_15325);
and U24433 (N_24433,N_15215,N_16334);
xnor U24434 (N_24434,N_18392,N_18200);
nor U24435 (N_24435,N_19559,N_19167);
and U24436 (N_24436,N_18322,N_19547);
xor U24437 (N_24437,N_16429,N_16924);
and U24438 (N_24438,N_19215,N_18239);
or U24439 (N_24439,N_16134,N_18238);
and U24440 (N_24440,N_18198,N_15875);
xnor U24441 (N_24441,N_18100,N_15616);
nand U24442 (N_24442,N_16247,N_15562);
nor U24443 (N_24443,N_17769,N_15387);
and U24444 (N_24444,N_17051,N_16927);
xnor U24445 (N_24445,N_19952,N_17565);
nand U24446 (N_24446,N_19502,N_16946);
nor U24447 (N_24447,N_16702,N_16551);
and U24448 (N_24448,N_17094,N_15995);
nor U24449 (N_24449,N_17668,N_19948);
or U24450 (N_24450,N_18446,N_19108);
nor U24451 (N_24451,N_18720,N_15977);
and U24452 (N_24452,N_17548,N_17970);
xor U24453 (N_24453,N_19629,N_16614);
xor U24454 (N_24454,N_19822,N_17895);
and U24455 (N_24455,N_19673,N_16228);
and U24456 (N_24456,N_15517,N_19547);
nand U24457 (N_24457,N_19765,N_17021);
nand U24458 (N_24458,N_16792,N_19342);
or U24459 (N_24459,N_16686,N_15128);
nor U24460 (N_24460,N_15238,N_15724);
nand U24461 (N_24461,N_18927,N_15892);
nand U24462 (N_24462,N_15296,N_19951);
and U24463 (N_24463,N_17269,N_17076);
and U24464 (N_24464,N_19888,N_16488);
or U24465 (N_24465,N_18745,N_17838);
xnor U24466 (N_24466,N_15135,N_19294);
or U24467 (N_24467,N_19618,N_17728);
nor U24468 (N_24468,N_18868,N_15835);
and U24469 (N_24469,N_16673,N_15809);
nor U24470 (N_24470,N_17682,N_15579);
nor U24471 (N_24471,N_16741,N_15808);
xnor U24472 (N_24472,N_19729,N_19142);
nor U24473 (N_24473,N_16490,N_17081);
nor U24474 (N_24474,N_18902,N_16431);
and U24475 (N_24475,N_18104,N_18109);
nor U24476 (N_24476,N_17407,N_19554);
or U24477 (N_24477,N_16043,N_16495);
xor U24478 (N_24478,N_15770,N_18466);
and U24479 (N_24479,N_15584,N_19395);
and U24480 (N_24480,N_17545,N_16139);
and U24481 (N_24481,N_16658,N_16398);
or U24482 (N_24482,N_17038,N_15513);
xor U24483 (N_24483,N_15923,N_19927);
xor U24484 (N_24484,N_16172,N_17550);
and U24485 (N_24485,N_16773,N_19982);
nand U24486 (N_24486,N_15053,N_19485);
and U24487 (N_24487,N_16514,N_17401);
xnor U24488 (N_24488,N_17873,N_15715);
nor U24489 (N_24489,N_18161,N_17345);
nand U24490 (N_24490,N_16885,N_16871);
nor U24491 (N_24491,N_18876,N_17675);
and U24492 (N_24492,N_15443,N_18704);
nand U24493 (N_24493,N_17712,N_17623);
nand U24494 (N_24494,N_18395,N_17959);
nand U24495 (N_24495,N_16316,N_15808);
or U24496 (N_24496,N_16458,N_15536);
xnor U24497 (N_24497,N_16777,N_17630);
and U24498 (N_24498,N_16272,N_19389);
nand U24499 (N_24499,N_19006,N_16972);
or U24500 (N_24500,N_17402,N_16665);
xnor U24501 (N_24501,N_19537,N_19692);
nand U24502 (N_24502,N_15303,N_16380);
and U24503 (N_24503,N_19253,N_19094);
and U24504 (N_24504,N_15033,N_16812);
nor U24505 (N_24505,N_17242,N_15960);
xor U24506 (N_24506,N_19312,N_17583);
or U24507 (N_24507,N_19577,N_18496);
nor U24508 (N_24508,N_15765,N_15546);
nand U24509 (N_24509,N_16108,N_15581);
xor U24510 (N_24510,N_18048,N_19806);
nand U24511 (N_24511,N_18657,N_15585);
nand U24512 (N_24512,N_16129,N_15343);
nand U24513 (N_24513,N_18137,N_16616);
and U24514 (N_24514,N_16484,N_19905);
or U24515 (N_24515,N_19083,N_15999);
xor U24516 (N_24516,N_19415,N_17654);
nand U24517 (N_24517,N_16384,N_17539);
and U24518 (N_24518,N_18215,N_19813);
or U24519 (N_24519,N_15314,N_18162);
and U24520 (N_24520,N_18804,N_18447);
or U24521 (N_24521,N_18871,N_17990);
or U24522 (N_24522,N_17622,N_18694);
or U24523 (N_24523,N_17594,N_17657);
nor U24524 (N_24524,N_19695,N_19175);
xnor U24525 (N_24525,N_18327,N_18670);
nor U24526 (N_24526,N_17625,N_17027);
xor U24527 (N_24527,N_17321,N_17588);
nand U24528 (N_24528,N_17974,N_15962);
nand U24529 (N_24529,N_18910,N_17339);
nor U24530 (N_24530,N_15701,N_17332);
xnor U24531 (N_24531,N_15378,N_17490);
and U24532 (N_24532,N_19908,N_18936);
nor U24533 (N_24533,N_19760,N_15072);
nor U24534 (N_24534,N_18787,N_19730);
and U24535 (N_24535,N_18604,N_18569);
nor U24536 (N_24536,N_18778,N_15566);
xnor U24537 (N_24537,N_18713,N_18346);
nand U24538 (N_24538,N_19692,N_17321);
xnor U24539 (N_24539,N_17002,N_17359);
and U24540 (N_24540,N_18129,N_16385);
nor U24541 (N_24541,N_18992,N_19614);
nand U24542 (N_24542,N_16089,N_15411);
nand U24543 (N_24543,N_16220,N_17001);
nand U24544 (N_24544,N_18098,N_19415);
or U24545 (N_24545,N_17979,N_17277);
nand U24546 (N_24546,N_18986,N_17296);
nand U24547 (N_24547,N_16759,N_15343);
xor U24548 (N_24548,N_18813,N_17930);
xnor U24549 (N_24549,N_18594,N_17013);
nand U24550 (N_24550,N_18996,N_19838);
nor U24551 (N_24551,N_17732,N_15025);
nor U24552 (N_24552,N_19345,N_19141);
nor U24553 (N_24553,N_16724,N_18667);
nor U24554 (N_24554,N_15702,N_15530);
and U24555 (N_24555,N_18312,N_18624);
nor U24556 (N_24556,N_16137,N_16879);
nor U24557 (N_24557,N_15912,N_16452);
xnor U24558 (N_24558,N_16890,N_19413);
nor U24559 (N_24559,N_15125,N_18339);
nor U24560 (N_24560,N_17152,N_16333);
or U24561 (N_24561,N_17424,N_19122);
and U24562 (N_24562,N_16777,N_19983);
and U24563 (N_24563,N_16803,N_15080);
nand U24564 (N_24564,N_19503,N_19581);
or U24565 (N_24565,N_19329,N_16631);
nand U24566 (N_24566,N_15947,N_17975);
or U24567 (N_24567,N_17576,N_19993);
nand U24568 (N_24568,N_19078,N_19730);
xnor U24569 (N_24569,N_15611,N_19210);
and U24570 (N_24570,N_18860,N_19665);
and U24571 (N_24571,N_19873,N_15421);
or U24572 (N_24572,N_15281,N_18038);
xor U24573 (N_24573,N_16887,N_19655);
or U24574 (N_24574,N_17983,N_17318);
or U24575 (N_24575,N_15371,N_19784);
nand U24576 (N_24576,N_19647,N_17975);
xor U24577 (N_24577,N_15889,N_16000);
nand U24578 (N_24578,N_19112,N_15785);
and U24579 (N_24579,N_15336,N_19036);
xnor U24580 (N_24580,N_19143,N_19268);
or U24581 (N_24581,N_16902,N_16506);
nor U24582 (N_24582,N_17576,N_15043);
and U24583 (N_24583,N_17258,N_18986);
and U24584 (N_24584,N_19041,N_15329);
nand U24585 (N_24585,N_17452,N_15682);
nor U24586 (N_24586,N_18367,N_18997);
nand U24587 (N_24587,N_16351,N_18414);
xnor U24588 (N_24588,N_16984,N_18531);
nand U24589 (N_24589,N_16650,N_19432);
and U24590 (N_24590,N_18486,N_15750);
or U24591 (N_24591,N_17099,N_16802);
xnor U24592 (N_24592,N_15851,N_15668);
nand U24593 (N_24593,N_17939,N_17675);
or U24594 (N_24594,N_19184,N_17233);
nor U24595 (N_24595,N_16826,N_17284);
xnor U24596 (N_24596,N_17984,N_17438);
xnor U24597 (N_24597,N_17586,N_17897);
nand U24598 (N_24598,N_17867,N_18464);
nand U24599 (N_24599,N_18776,N_17572);
nor U24600 (N_24600,N_15555,N_15216);
nor U24601 (N_24601,N_18923,N_19755);
nand U24602 (N_24602,N_19975,N_19089);
xor U24603 (N_24603,N_19976,N_19233);
xor U24604 (N_24604,N_17318,N_15691);
or U24605 (N_24605,N_19457,N_18006);
nand U24606 (N_24606,N_19332,N_19899);
nor U24607 (N_24607,N_19157,N_17775);
nand U24608 (N_24608,N_19353,N_16993);
nor U24609 (N_24609,N_18925,N_15970);
nor U24610 (N_24610,N_19240,N_16083);
nand U24611 (N_24611,N_18629,N_18382);
nand U24612 (N_24612,N_19038,N_16432);
or U24613 (N_24613,N_16144,N_15587);
or U24614 (N_24614,N_19865,N_15559);
and U24615 (N_24615,N_19908,N_16465);
nor U24616 (N_24616,N_18260,N_16749);
xnor U24617 (N_24617,N_17339,N_16629);
nor U24618 (N_24618,N_16308,N_17012);
xor U24619 (N_24619,N_15622,N_19982);
and U24620 (N_24620,N_16930,N_18275);
nand U24621 (N_24621,N_19085,N_19205);
nand U24622 (N_24622,N_17042,N_15847);
xnor U24623 (N_24623,N_19660,N_16521);
nand U24624 (N_24624,N_18146,N_16766);
nand U24625 (N_24625,N_19442,N_19986);
nor U24626 (N_24626,N_18067,N_18215);
and U24627 (N_24627,N_19271,N_19199);
and U24628 (N_24628,N_16493,N_17715);
nand U24629 (N_24629,N_19089,N_17888);
and U24630 (N_24630,N_16015,N_16751);
xnor U24631 (N_24631,N_15224,N_19770);
and U24632 (N_24632,N_17118,N_19645);
nand U24633 (N_24633,N_16715,N_16881);
and U24634 (N_24634,N_18738,N_17348);
nand U24635 (N_24635,N_17343,N_19793);
or U24636 (N_24636,N_15341,N_17789);
or U24637 (N_24637,N_15133,N_16612);
nand U24638 (N_24638,N_17183,N_15213);
nor U24639 (N_24639,N_18977,N_18753);
nand U24640 (N_24640,N_16050,N_17410);
nand U24641 (N_24641,N_19524,N_15345);
and U24642 (N_24642,N_15490,N_16666);
nand U24643 (N_24643,N_17130,N_17397);
and U24644 (N_24644,N_17963,N_17236);
or U24645 (N_24645,N_16995,N_19635);
or U24646 (N_24646,N_18038,N_15678);
nor U24647 (N_24647,N_19107,N_16554);
or U24648 (N_24648,N_15973,N_18029);
nand U24649 (N_24649,N_16364,N_18165);
nor U24650 (N_24650,N_15457,N_16769);
xor U24651 (N_24651,N_18051,N_15476);
nor U24652 (N_24652,N_18124,N_18772);
xor U24653 (N_24653,N_19534,N_18175);
xor U24654 (N_24654,N_16131,N_16840);
and U24655 (N_24655,N_18130,N_15790);
xor U24656 (N_24656,N_19057,N_18170);
xor U24657 (N_24657,N_15158,N_15990);
or U24658 (N_24658,N_16956,N_17425);
or U24659 (N_24659,N_19032,N_16511);
or U24660 (N_24660,N_15314,N_18074);
nand U24661 (N_24661,N_15173,N_16997);
and U24662 (N_24662,N_18106,N_16910);
or U24663 (N_24663,N_15519,N_17539);
nand U24664 (N_24664,N_16292,N_16087);
or U24665 (N_24665,N_15609,N_19186);
nor U24666 (N_24666,N_15071,N_18954);
nand U24667 (N_24667,N_18793,N_18945);
and U24668 (N_24668,N_15341,N_18026);
nor U24669 (N_24669,N_18298,N_15573);
xnor U24670 (N_24670,N_18038,N_19060);
and U24671 (N_24671,N_18466,N_15973);
xnor U24672 (N_24672,N_17587,N_17406);
nand U24673 (N_24673,N_19631,N_17822);
nand U24674 (N_24674,N_15716,N_18553);
nand U24675 (N_24675,N_16562,N_15792);
xnor U24676 (N_24676,N_15699,N_18751);
nor U24677 (N_24677,N_18700,N_15484);
and U24678 (N_24678,N_17854,N_17336);
nand U24679 (N_24679,N_19687,N_18679);
nor U24680 (N_24680,N_15544,N_19661);
nand U24681 (N_24681,N_16010,N_15032);
and U24682 (N_24682,N_16374,N_17731);
nor U24683 (N_24683,N_15427,N_19171);
or U24684 (N_24684,N_19150,N_16514);
xor U24685 (N_24685,N_16629,N_18696);
nand U24686 (N_24686,N_18637,N_15065);
nand U24687 (N_24687,N_18215,N_16690);
nor U24688 (N_24688,N_16892,N_19329);
or U24689 (N_24689,N_18081,N_17019);
or U24690 (N_24690,N_16135,N_17818);
nor U24691 (N_24691,N_15988,N_17123);
nor U24692 (N_24692,N_17117,N_18538);
xor U24693 (N_24693,N_18517,N_19544);
nor U24694 (N_24694,N_18586,N_19038);
or U24695 (N_24695,N_17484,N_16283);
nor U24696 (N_24696,N_17432,N_15658);
or U24697 (N_24697,N_17057,N_19891);
nand U24698 (N_24698,N_17463,N_19706);
or U24699 (N_24699,N_16589,N_19668);
xor U24700 (N_24700,N_15992,N_15373);
xnor U24701 (N_24701,N_17779,N_17934);
nand U24702 (N_24702,N_18434,N_17422);
or U24703 (N_24703,N_16959,N_18236);
nand U24704 (N_24704,N_17655,N_15948);
or U24705 (N_24705,N_18038,N_17503);
or U24706 (N_24706,N_16331,N_16089);
nand U24707 (N_24707,N_17298,N_17157);
nand U24708 (N_24708,N_19327,N_19767);
or U24709 (N_24709,N_16257,N_16839);
or U24710 (N_24710,N_17641,N_15495);
or U24711 (N_24711,N_17152,N_16669);
xor U24712 (N_24712,N_16822,N_19137);
and U24713 (N_24713,N_19850,N_17364);
or U24714 (N_24714,N_17005,N_16029);
or U24715 (N_24715,N_15094,N_19116);
nand U24716 (N_24716,N_15147,N_15744);
or U24717 (N_24717,N_16648,N_19658);
xnor U24718 (N_24718,N_16258,N_18930);
nor U24719 (N_24719,N_16782,N_15039);
nand U24720 (N_24720,N_19061,N_19959);
nand U24721 (N_24721,N_19001,N_18831);
nor U24722 (N_24722,N_16956,N_17330);
nand U24723 (N_24723,N_16601,N_16447);
nor U24724 (N_24724,N_15842,N_18292);
nor U24725 (N_24725,N_19310,N_19475);
xor U24726 (N_24726,N_17755,N_19950);
xnor U24727 (N_24727,N_16090,N_18584);
or U24728 (N_24728,N_19561,N_16717);
nor U24729 (N_24729,N_17709,N_19717);
or U24730 (N_24730,N_16794,N_16056);
or U24731 (N_24731,N_17729,N_17373);
and U24732 (N_24732,N_16640,N_19671);
nand U24733 (N_24733,N_15711,N_15542);
xnor U24734 (N_24734,N_15741,N_19543);
or U24735 (N_24735,N_18818,N_15075);
and U24736 (N_24736,N_18537,N_18952);
and U24737 (N_24737,N_15334,N_15832);
nand U24738 (N_24738,N_17108,N_19741);
or U24739 (N_24739,N_17036,N_19882);
nor U24740 (N_24740,N_15501,N_17773);
xnor U24741 (N_24741,N_15498,N_15425);
nor U24742 (N_24742,N_15571,N_18833);
and U24743 (N_24743,N_15764,N_18514);
or U24744 (N_24744,N_17868,N_17125);
and U24745 (N_24745,N_18752,N_17080);
xnor U24746 (N_24746,N_18740,N_15042);
and U24747 (N_24747,N_16886,N_19065);
nor U24748 (N_24748,N_18246,N_18520);
xor U24749 (N_24749,N_18418,N_17582);
and U24750 (N_24750,N_18161,N_17385);
nor U24751 (N_24751,N_15994,N_19789);
nor U24752 (N_24752,N_16242,N_15283);
and U24753 (N_24753,N_18094,N_15357);
and U24754 (N_24754,N_15155,N_18710);
nand U24755 (N_24755,N_15119,N_15658);
xor U24756 (N_24756,N_19712,N_19747);
nor U24757 (N_24757,N_18389,N_16087);
nand U24758 (N_24758,N_17500,N_18236);
xnor U24759 (N_24759,N_18341,N_18408);
or U24760 (N_24760,N_18466,N_16515);
and U24761 (N_24761,N_18478,N_16144);
or U24762 (N_24762,N_17610,N_15088);
or U24763 (N_24763,N_19887,N_16559);
xor U24764 (N_24764,N_19853,N_18937);
nor U24765 (N_24765,N_15267,N_18583);
nor U24766 (N_24766,N_16544,N_17884);
xor U24767 (N_24767,N_16070,N_17477);
nor U24768 (N_24768,N_15875,N_17545);
nor U24769 (N_24769,N_17402,N_17094);
nand U24770 (N_24770,N_16172,N_16554);
nand U24771 (N_24771,N_17933,N_16542);
xor U24772 (N_24772,N_18127,N_17464);
xor U24773 (N_24773,N_16933,N_18714);
xnor U24774 (N_24774,N_16934,N_18823);
nand U24775 (N_24775,N_17928,N_18049);
xor U24776 (N_24776,N_19541,N_19992);
nand U24777 (N_24777,N_19901,N_17150);
and U24778 (N_24778,N_18024,N_18005);
or U24779 (N_24779,N_16613,N_15400);
xor U24780 (N_24780,N_19842,N_16080);
or U24781 (N_24781,N_18837,N_17806);
or U24782 (N_24782,N_16186,N_16948);
xor U24783 (N_24783,N_18723,N_16002);
and U24784 (N_24784,N_19670,N_17761);
or U24785 (N_24785,N_17719,N_18274);
and U24786 (N_24786,N_18910,N_19377);
xnor U24787 (N_24787,N_17081,N_15903);
or U24788 (N_24788,N_18463,N_19093);
nor U24789 (N_24789,N_18435,N_19976);
nand U24790 (N_24790,N_17094,N_15112);
xor U24791 (N_24791,N_17123,N_16348);
and U24792 (N_24792,N_19534,N_15134);
nand U24793 (N_24793,N_15775,N_18416);
or U24794 (N_24794,N_15045,N_15464);
nor U24795 (N_24795,N_19208,N_17768);
xor U24796 (N_24796,N_16595,N_16204);
or U24797 (N_24797,N_17064,N_17789);
and U24798 (N_24798,N_15827,N_17700);
nor U24799 (N_24799,N_18068,N_18376);
or U24800 (N_24800,N_17367,N_17853);
and U24801 (N_24801,N_19822,N_17671);
or U24802 (N_24802,N_15734,N_17786);
xnor U24803 (N_24803,N_18915,N_18311);
and U24804 (N_24804,N_17651,N_15689);
or U24805 (N_24805,N_16636,N_16092);
or U24806 (N_24806,N_19510,N_16543);
nand U24807 (N_24807,N_16012,N_16163);
nand U24808 (N_24808,N_18592,N_16512);
xnor U24809 (N_24809,N_18117,N_18771);
nor U24810 (N_24810,N_17215,N_16147);
or U24811 (N_24811,N_17205,N_17154);
nor U24812 (N_24812,N_17866,N_15918);
and U24813 (N_24813,N_15084,N_19001);
nor U24814 (N_24814,N_16148,N_19014);
or U24815 (N_24815,N_16301,N_19783);
xnor U24816 (N_24816,N_16777,N_16311);
or U24817 (N_24817,N_17941,N_17601);
and U24818 (N_24818,N_19554,N_15622);
nor U24819 (N_24819,N_16672,N_19890);
and U24820 (N_24820,N_16845,N_16975);
xnor U24821 (N_24821,N_15263,N_19535);
nand U24822 (N_24822,N_15354,N_16445);
and U24823 (N_24823,N_18181,N_17462);
or U24824 (N_24824,N_18858,N_17117);
nor U24825 (N_24825,N_19696,N_17327);
and U24826 (N_24826,N_18515,N_19460);
nand U24827 (N_24827,N_15223,N_17965);
nor U24828 (N_24828,N_15961,N_19358);
nor U24829 (N_24829,N_17190,N_18005);
or U24830 (N_24830,N_18088,N_15554);
or U24831 (N_24831,N_19381,N_18318);
and U24832 (N_24832,N_17662,N_17131);
and U24833 (N_24833,N_16137,N_18006);
or U24834 (N_24834,N_15865,N_15204);
or U24835 (N_24835,N_17475,N_15468);
nand U24836 (N_24836,N_16876,N_19387);
xnor U24837 (N_24837,N_19408,N_17258);
xor U24838 (N_24838,N_15348,N_18495);
nor U24839 (N_24839,N_15110,N_15138);
or U24840 (N_24840,N_19866,N_15109);
and U24841 (N_24841,N_19295,N_15831);
or U24842 (N_24842,N_19114,N_19926);
and U24843 (N_24843,N_18909,N_19660);
nor U24844 (N_24844,N_19078,N_15053);
and U24845 (N_24845,N_19496,N_18653);
xnor U24846 (N_24846,N_17917,N_16708);
nor U24847 (N_24847,N_17915,N_15643);
nand U24848 (N_24848,N_16328,N_18151);
nand U24849 (N_24849,N_19698,N_18096);
and U24850 (N_24850,N_17366,N_19890);
or U24851 (N_24851,N_18899,N_15896);
xor U24852 (N_24852,N_15495,N_17167);
nand U24853 (N_24853,N_15990,N_16945);
and U24854 (N_24854,N_19473,N_15386);
xnor U24855 (N_24855,N_18663,N_15417);
nand U24856 (N_24856,N_15682,N_18101);
nand U24857 (N_24857,N_16944,N_19905);
nand U24858 (N_24858,N_19422,N_15978);
nand U24859 (N_24859,N_19353,N_16923);
and U24860 (N_24860,N_19473,N_18169);
nor U24861 (N_24861,N_16748,N_19713);
nand U24862 (N_24862,N_19463,N_15448);
nand U24863 (N_24863,N_19351,N_18629);
and U24864 (N_24864,N_17662,N_17949);
nand U24865 (N_24865,N_17982,N_15198);
nor U24866 (N_24866,N_17454,N_15910);
or U24867 (N_24867,N_18302,N_16559);
or U24868 (N_24868,N_15411,N_16984);
and U24869 (N_24869,N_15462,N_15387);
nand U24870 (N_24870,N_15726,N_18593);
nand U24871 (N_24871,N_18841,N_18335);
and U24872 (N_24872,N_15738,N_19381);
nand U24873 (N_24873,N_19649,N_16465);
nand U24874 (N_24874,N_16061,N_16977);
nand U24875 (N_24875,N_19094,N_16903);
nand U24876 (N_24876,N_16661,N_19458);
nand U24877 (N_24877,N_19262,N_19861);
and U24878 (N_24878,N_19472,N_16679);
xnor U24879 (N_24879,N_18845,N_15827);
xor U24880 (N_24880,N_16722,N_16608);
or U24881 (N_24881,N_17137,N_18857);
xor U24882 (N_24882,N_15307,N_18698);
or U24883 (N_24883,N_15164,N_15236);
and U24884 (N_24884,N_17479,N_16286);
nand U24885 (N_24885,N_15278,N_17721);
xor U24886 (N_24886,N_16010,N_16807);
or U24887 (N_24887,N_15694,N_18938);
and U24888 (N_24888,N_15805,N_16619);
nand U24889 (N_24889,N_18598,N_16015);
and U24890 (N_24890,N_16019,N_15772);
nor U24891 (N_24891,N_19884,N_18833);
or U24892 (N_24892,N_19758,N_16146);
and U24893 (N_24893,N_15716,N_15533);
nand U24894 (N_24894,N_19331,N_15611);
nand U24895 (N_24895,N_18643,N_17921);
xnor U24896 (N_24896,N_19950,N_16926);
xor U24897 (N_24897,N_15304,N_18166);
nand U24898 (N_24898,N_18458,N_17339);
or U24899 (N_24899,N_19907,N_18340);
or U24900 (N_24900,N_16225,N_15667);
and U24901 (N_24901,N_17722,N_19061);
nand U24902 (N_24902,N_18884,N_15987);
and U24903 (N_24903,N_17417,N_18866);
and U24904 (N_24904,N_18035,N_18553);
nor U24905 (N_24905,N_16309,N_17520);
nor U24906 (N_24906,N_17390,N_19875);
nand U24907 (N_24907,N_16010,N_18073);
nand U24908 (N_24908,N_16787,N_15843);
nor U24909 (N_24909,N_18200,N_19577);
or U24910 (N_24910,N_18172,N_19436);
nor U24911 (N_24911,N_16068,N_17477);
or U24912 (N_24912,N_15764,N_17663);
xnor U24913 (N_24913,N_19193,N_18110);
nand U24914 (N_24914,N_16854,N_18721);
nand U24915 (N_24915,N_15687,N_15129);
and U24916 (N_24916,N_18177,N_18246);
nor U24917 (N_24917,N_16569,N_15628);
xor U24918 (N_24918,N_16685,N_18842);
and U24919 (N_24919,N_19853,N_18137);
and U24920 (N_24920,N_16950,N_19506);
xnor U24921 (N_24921,N_18106,N_18314);
or U24922 (N_24922,N_18670,N_19033);
xnor U24923 (N_24923,N_15367,N_16001);
and U24924 (N_24924,N_16892,N_19479);
or U24925 (N_24925,N_15122,N_18868);
nand U24926 (N_24926,N_15293,N_15615);
nor U24927 (N_24927,N_17608,N_18797);
xnor U24928 (N_24928,N_16655,N_15946);
or U24929 (N_24929,N_16528,N_15549);
and U24930 (N_24930,N_15935,N_19607);
and U24931 (N_24931,N_18112,N_19253);
nor U24932 (N_24932,N_18511,N_19241);
and U24933 (N_24933,N_17167,N_18189);
xnor U24934 (N_24934,N_17121,N_18134);
nor U24935 (N_24935,N_18705,N_19580);
nor U24936 (N_24936,N_16014,N_16381);
and U24937 (N_24937,N_17250,N_19454);
nor U24938 (N_24938,N_19751,N_18957);
or U24939 (N_24939,N_17605,N_19090);
nor U24940 (N_24940,N_15341,N_19591);
nand U24941 (N_24941,N_15242,N_19387);
xor U24942 (N_24942,N_18756,N_18577);
xor U24943 (N_24943,N_16515,N_18002);
and U24944 (N_24944,N_18916,N_18896);
and U24945 (N_24945,N_17219,N_16122);
and U24946 (N_24946,N_19543,N_15975);
xnor U24947 (N_24947,N_17169,N_16195);
xnor U24948 (N_24948,N_16190,N_17152);
and U24949 (N_24949,N_16090,N_15783);
nor U24950 (N_24950,N_18153,N_15264);
or U24951 (N_24951,N_17224,N_17500);
xnor U24952 (N_24952,N_15250,N_16546);
and U24953 (N_24953,N_17702,N_15179);
and U24954 (N_24954,N_16003,N_17654);
xor U24955 (N_24955,N_19801,N_15291);
or U24956 (N_24956,N_17678,N_19741);
xor U24957 (N_24957,N_15603,N_18677);
or U24958 (N_24958,N_15411,N_18025);
xnor U24959 (N_24959,N_18453,N_19698);
xnor U24960 (N_24960,N_19089,N_19569);
xor U24961 (N_24961,N_18675,N_19911);
and U24962 (N_24962,N_18280,N_19266);
nor U24963 (N_24963,N_17080,N_19523);
and U24964 (N_24964,N_17744,N_17063);
nor U24965 (N_24965,N_18105,N_18015);
nor U24966 (N_24966,N_19444,N_19371);
xnor U24967 (N_24967,N_15273,N_16939);
and U24968 (N_24968,N_16738,N_15579);
xnor U24969 (N_24969,N_15605,N_16835);
nor U24970 (N_24970,N_18974,N_18683);
and U24971 (N_24971,N_16090,N_19861);
or U24972 (N_24972,N_19842,N_16497);
nor U24973 (N_24973,N_15940,N_17748);
nand U24974 (N_24974,N_18822,N_16482);
nand U24975 (N_24975,N_16785,N_19572);
and U24976 (N_24976,N_15728,N_18138);
xor U24977 (N_24977,N_18235,N_18683);
and U24978 (N_24978,N_16401,N_15945);
or U24979 (N_24979,N_15850,N_15407);
and U24980 (N_24980,N_19632,N_15717);
nand U24981 (N_24981,N_19584,N_19435);
xor U24982 (N_24982,N_17609,N_15106);
nor U24983 (N_24983,N_19836,N_16437);
nor U24984 (N_24984,N_16929,N_15051);
and U24985 (N_24985,N_16296,N_17076);
or U24986 (N_24986,N_17590,N_16138);
nor U24987 (N_24987,N_16168,N_15311);
or U24988 (N_24988,N_19472,N_15879);
nand U24989 (N_24989,N_15946,N_17196);
xor U24990 (N_24990,N_18563,N_19439);
xor U24991 (N_24991,N_18656,N_19227);
and U24992 (N_24992,N_19427,N_17783);
or U24993 (N_24993,N_15817,N_15035);
or U24994 (N_24994,N_16305,N_18835);
or U24995 (N_24995,N_16897,N_15182);
nor U24996 (N_24996,N_17888,N_15568);
nor U24997 (N_24997,N_15287,N_18176);
nor U24998 (N_24998,N_15509,N_17247);
nor U24999 (N_24999,N_16926,N_19899);
and UO_0 (O_0,N_24481,N_24064);
or UO_1 (O_1,N_20882,N_21817);
or UO_2 (O_2,N_24025,N_20087);
xnor UO_3 (O_3,N_24988,N_22924);
nor UO_4 (O_4,N_21418,N_21573);
nand UO_5 (O_5,N_20509,N_23052);
and UO_6 (O_6,N_23714,N_21597);
nand UO_7 (O_7,N_21047,N_23545);
nor UO_8 (O_8,N_23834,N_22124);
xor UO_9 (O_9,N_21333,N_22860);
nand UO_10 (O_10,N_22346,N_24100);
xor UO_11 (O_11,N_23594,N_24029);
nor UO_12 (O_12,N_22699,N_23198);
xor UO_13 (O_13,N_21759,N_20492);
nor UO_14 (O_14,N_20999,N_22022);
or UO_15 (O_15,N_22423,N_22900);
nand UO_16 (O_16,N_20285,N_22286);
nand UO_17 (O_17,N_21571,N_22232);
and UO_18 (O_18,N_22329,N_23266);
xnor UO_19 (O_19,N_21528,N_20456);
nand UO_20 (O_20,N_23434,N_21001);
and UO_21 (O_21,N_21598,N_21673);
nor UO_22 (O_22,N_23194,N_20115);
nand UO_23 (O_23,N_24812,N_24341);
nand UO_24 (O_24,N_20817,N_21715);
or UO_25 (O_25,N_21002,N_21622);
or UO_26 (O_26,N_24084,N_23452);
nand UO_27 (O_27,N_20311,N_21379);
nand UO_28 (O_28,N_20338,N_22103);
or UO_29 (O_29,N_21820,N_22717);
nor UO_30 (O_30,N_21752,N_21319);
and UO_31 (O_31,N_24779,N_21375);
and UO_32 (O_32,N_20761,N_21708);
xor UO_33 (O_33,N_21810,N_22130);
and UO_34 (O_34,N_21056,N_23917);
nor UO_35 (O_35,N_22869,N_22009);
nand UO_36 (O_36,N_23382,N_21701);
or UO_37 (O_37,N_20126,N_20365);
nand UO_38 (O_38,N_24081,N_22040);
nand UO_39 (O_39,N_24174,N_21758);
and UO_40 (O_40,N_24499,N_24076);
or UO_41 (O_41,N_21142,N_23497);
xnor UO_42 (O_42,N_22219,N_21407);
nor UO_43 (O_43,N_23312,N_22207);
and UO_44 (O_44,N_20652,N_21464);
or UO_45 (O_45,N_20467,N_21412);
or UO_46 (O_46,N_20432,N_24284);
xor UO_47 (O_47,N_22969,N_24620);
and UO_48 (O_48,N_20972,N_24317);
or UO_49 (O_49,N_20867,N_24408);
and UO_50 (O_50,N_20757,N_22691);
nand UO_51 (O_51,N_23618,N_23164);
nor UO_52 (O_52,N_22623,N_23478);
or UO_53 (O_53,N_22029,N_22045);
or UO_54 (O_54,N_24947,N_24855);
nor UO_55 (O_55,N_21267,N_21702);
xnor UO_56 (O_56,N_24963,N_21683);
xor UO_57 (O_57,N_22920,N_20546);
or UO_58 (O_58,N_23852,N_22039);
and UO_59 (O_59,N_20109,N_23946);
xnor UO_60 (O_60,N_23649,N_20657);
nand UO_61 (O_61,N_24336,N_23664);
xor UO_62 (O_62,N_24601,N_24639);
xnor UO_63 (O_63,N_20805,N_21886);
nor UO_64 (O_64,N_23627,N_23785);
nand UO_65 (O_65,N_20500,N_24810);
nand UO_66 (O_66,N_22562,N_22706);
nand UO_67 (O_67,N_20890,N_22633);
and UO_68 (O_68,N_20874,N_21014);
nand UO_69 (O_69,N_22988,N_23445);
nand UO_70 (O_70,N_22795,N_21525);
or UO_71 (O_71,N_23994,N_21939);
or UO_72 (O_72,N_23125,N_24889);
xor UO_73 (O_73,N_24367,N_21157);
nand UO_74 (O_74,N_24490,N_23463);
xor UO_75 (O_75,N_24980,N_23626);
nand UO_76 (O_76,N_20489,N_24063);
xnor UO_77 (O_77,N_23555,N_24722);
or UO_78 (O_78,N_22689,N_21740);
and UO_79 (O_79,N_21247,N_20577);
and UO_80 (O_80,N_23993,N_23591);
nand UO_81 (O_81,N_20935,N_22125);
or UO_82 (O_82,N_20856,N_20097);
or UO_83 (O_83,N_21467,N_24672);
nand UO_84 (O_84,N_20244,N_21544);
nor UO_85 (O_85,N_21484,N_24933);
nand UO_86 (O_86,N_22823,N_22761);
nand UO_87 (O_87,N_22858,N_20584);
xor UO_88 (O_88,N_23022,N_22181);
xor UO_89 (O_89,N_23127,N_20322);
xor UO_90 (O_90,N_23830,N_21881);
and UO_91 (O_91,N_21489,N_22553);
and UO_92 (O_92,N_23997,N_24679);
and UO_93 (O_93,N_24124,N_24348);
and UO_94 (O_94,N_20634,N_23751);
xnor UO_95 (O_95,N_20715,N_20305);
nor UO_96 (O_96,N_21951,N_22282);
or UO_97 (O_97,N_23256,N_23531);
nand UO_98 (O_98,N_23988,N_24079);
and UO_99 (O_99,N_23914,N_23066);
and UO_100 (O_100,N_22978,N_24460);
or UO_101 (O_101,N_22873,N_21200);
or UO_102 (O_102,N_21018,N_24383);
nor UO_103 (O_103,N_21588,N_23747);
nand UO_104 (O_104,N_20737,N_24182);
and UO_105 (O_105,N_22440,N_21317);
nor UO_106 (O_106,N_22109,N_22825);
or UO_107 (O_107,N_20818,N_21383);
nor UO_108 (O_108,N_22250,N_22437);
nand UO_109 (O_109,N_21378,N_24016);
and UO_110 (O_110,N_23344,N_24128);
and UO_111 (O_111,N_21746,N_22494);
nand UO_112 (O_112,N_22670,N_21616);
xnor UO_113 (O_113,N_22913,N_20175);
xor UO_114 (O_114,N_24010,N_21648);
and UO_115 (O_115,N_24188,N_23244);
and UO_116 (O_116,N_22237,N_21025);
xnor UO_117 (O_117,N_24323,N_21459);
or UO_118 (O_118,N_22031,N_23701);
nor UO_119 (O_119,N_23204,N_21520);
and UO_120 (O_120,N_21431,N_24739);
xnor UO_121 (O_121,N_20402,N_24822);
xnor UO_122 (O_122,N_20098,N_21635);
or UO_123 (O_123,N_20736,N_24516);
nand UO_124 (O_124,N_21633,N_21727);
xor UO_125 (O_125,N_22407,N_23778);
or UO_126 (O_126,N_24417,N_24036);
nand UO_127 (O_127,N_24600,N_21154);
xor UO_128 (O_128,N_23425,N_20060);
xnor UO_129 (O_129,N_22887,N_20021);
or UO_130 (O_130,N_23119,N_21837);
and UO_131 (O_131,N_20096,N_22327);
and UO_132 (O_132,N_24451,N_20672);
nor UO_133 (O_133,N_22656,N_24576);
or UO_134 (O_134,N_20202,N_23813);
nand UO_135 (O_135,N_23854,N_24609);
nand UO_136 (O_136,N_23697,N_21706);
nor UO_137 (O_137,N_23279,N_20531);
nand UO_138 (O_138,N_23487,N_24015);
nand UO_139 (O_139,N_20862,N_24617);
or UO_140 (O_140,N_22069,N_23527);
and UO_141 (O_141,N_23176,N_20441);
xnor UO_142 (O_142,N_24682,N_23982);
xnor UO_143 (O_143,N_21032,N_22740);
and UO_144 (O_144,N_20340,N_23901);
nand UO_145 (O_145,N_23058,N_23687);
and UO_146 (O_146,N_20300,N_24935);
nor UO_147 (O_147,N_24753,N_23357);
nor UO_148 (O_148,N_22291,N_20947);
xor UO_149 (O_149,N_23375,N_21092);
xnor UO_150 (O_150,N_22230,N_22246);
and UO_151 (O_151,N_22905,N_21191);
or UO_152 (O_152,N_21285,N_22963);
nand UO_153 (O_153,N_21495,N_22324);
nor UO_154 (O_154,N_23289,N_20783);
and UO_155 (O_155,N_21127,N_23328);
and UO_156 (O_156,N_20752,N_20259);
xnor UO_157 (O_157,N_20496,N_23325);
or UO_158 (O_158,N_20477,N_20434);
xnor UO_159 (O_159,N_20996,N_24102);
and UO_160 (O_160,N_23908,N_22629);
or UO_161 (O_161,N_22196,N_24241);
xnor UO_162 (O_162,N_21907,N_22059);
and UO_163 (O_163,N_24998,N_23689);
nand UO_164 (O_164,N_20258,N_23799);
or UO_165 (O_165,N_24320,N_20237);
or UO_166 (O_166,N_21862,N_20483);
and UO_167 (O_167,N_21090,N_23568);
or UO_168 (O_168,N_23932,N_20049);
and UO_169 (O_169,N_20325,N_24519);
and UO_170 (O_170,N_22742,N_21481);
xor UO_171 (O_171,N_20036,N_24007);
or UO_172 (O_172,N_20457,N_24254);
nor UO_173 (O_173,N_23306,N_24240);
xor UO_174 (O_174,N_21334,N_23303);
and UO_175 (O_175,N_21404,N_20583);
or UO_176 (O_176,N_20621,N_23313);
and UO_177 (O_177,N_20829,N_24875);
and UO_178 (O_178,N_24528,N_21754);
and UO_179 (O_179,N_20560,N_21680);
nand UO_180 (O_180,N_21340,N_24194);
nand UO_181 (O_181,N_22087,N_24986);
nor UO_182 (O_182,N_20134,N_21714);
and UO_183 (O_183,N_22228,N_22705);
nand UO_184 (O_184,N_21162,N_20253);
xnor UO_185 (O_185,N_20607,N_24273);
nor UO_186 (O_186,N_20662,N_20385);
nand UO_187 (O_187,N_21362,N_24234);
nor UO_188 (O_188,N_23742,N_24390);
xnor UO_189 (O_189,N_24313,N_22410);
nor UO_190 (O_190,N_22068,N_21436);
or UO_191 (O_191,N_22077,N_23953);
nand UO_192 (O_192,N_24665,N_24982);
and UO_193 (O_193,N_24835,N_20241);
nand UO_194 (O_194,N_24981,N_24031);
and UO_195 (O_195,N_21729,N_21562);
and UO_196 (O_196,N_21400,N_22431);
or UO_197 (O_197,N_21087,N_24400);
or UO_198 (O_198,N_24940,N_20376);
and UO_199 (O_199,N_21380,N_24869);
nor UO_200 (O_200,N_24013,N_24728);
or UO_201 (O_201,N_23524,N_23784);
nor UO_202 (O_202,N_24326,N_23581);
nand UO_203 (O_203,N_21813,N_21197);
and UO_204 (O_204,N_24120,N_24233);
or UO_205 (O_205,N_20886,N_24337);
xnor UO_206 (O_206,N_24813,N_23061);
or UO_207 (O_207,N_20991,N_20388);
and UO_208 (O_208,N_23758,N_20027);
and UO_209 (O_209,N_21647,N_24589);
or UO_210 (O_210,N_21377,N_22436);
xor UO_211 (O_211,N_22121,N_22006);
and UO_212 (O_212,N_21411,N_20112);
nor UO_213 (O_213,N_20361,N_22719);
nor UO_214 (O_214,N_21438,N_24177);
or UO_215 (O_215,N_24842,N_22676);
nand UO_216 (O_216,N_23647,N_21839);
xnor UO_217 (O_217,N_20077,N_22734);
nor UO_218 (O_218,N_21114,N_24072);
xnor UO_219 (O_219,N_22395,N_21156);
nand UO_220 (O_220,N_24692,N_23596);
or UO_221 (O_221,N_20278,N_21630);
or UO_222 (O_222,N_24069,N_20415);
and UO_223 (O_223,N_21892,N_23317);
and UO_224 (O_224,N_22642,N_20083);
nor UO_225 (O_225,N_21560,N_23835);
or UO_226 (O_226,N_24185,N_20032);
or UO_227 (O_227,N_23533,N_23214);
and UO_228 (O_228,N_22224,N_24238);
xnor UO_229 (O_229,N_21576,N_24474);
nand UO_230 (O_230,N_24643,N_21624);
or UO_231 (O_231,N_24555,N_20649);
xor UO_232 (O_232,N_21502,N_21969);
xor UO_233 (O_233,N_20460,N_23693);
xnor UO_234 (O_234,N_20919,N_22620);
or UO_235 (O_235,N_23959,N_20254);
nor UO_236 (O_236,N_20616,N_22217);
or UO_237 (O_237,N_22752,N_23020);
or UO_238 (O_238,N_24514,N_21337);
xor UO_239 (O_239,N_24138,N_24738);
or UO_240 (O_240,N_24274,N_23404);
and UO_241 (O_241,N_20262,N_24552);
or UO_242 (O_242,N_20288,N_20085);
nor UO_243 (O_243,N_20143,N_23105);
nor UO_244 (O_244,N_20110,N_21711);
xor UO_245 (O_245,N_21444,N_20487);
and UO_246 (O_246,N_20863,N_22094);
or UO_247 (O_247,N_21475,N_21718);
xor UO_248 (O_248,N_20786,N_22764);
and UO_249 (O_249,N_23838,N_21026);
or UO_250 (O_250,N_21970,N_21590);
xnor UO_251 (O_251,N_24494,N_20068);
nor UO_252 (O_252,N_21141,N_21028);
xnor UO_253 (O_253,N_23674,N_24463);
and UO_254 (O_254,N_20824,N_22892);
or UO_255 (O_255,N_23707,N_21572);
and UO_256 (O_256,N_23358,N_23002);
xor UO_257 (O_257,N_21486,N_20756);
nor UO_258 (O_258,N_24428,N_20907);
nand UO_259 (O_259,N_21506,N_20104);
or UO_260 (O_260,N_20810,N_23226);
nand UO_261 (O_261,N_21239,N_22152);
nor UO_262 (O_262,N_21356,N_22527);
nor UO_263 (O_263,N_23826,N_23655);
or UO_264 (O_264,N_23297,N_21720);
xnor UO_265 (O_265,N_22162,N_23413);
or UO_266 (O_266,N_20592,N_20732);
or UO_267 (O_267,N_22991,N_23130);
nor UO_268 (O_268,N_24533,N_21973);
nor UO_269 (O_269,N_22272,N_22730);
nand UO_270 (O_270,N_21555,N_24252);
nor UO_271 (O_271,N_20050,N_21504);
and UO_272 (O_272,N_21921,N_20651);
nor UO_273 (O_273,N_22400,N_20895);
nor UO_274 (O_274,N_20357,N_23380);
or UO_275 (O_275,N_22409,N_24741);
nor UO_276 (O_276,N_21498,N_23639);
and UO_277 (O_277,N_21449,N_20681);
and UO_278 (O_278,N_21113,N_24944);
or UO_279 (O_279,N_24155,N_21744);
xnor UO_280 (O_280,N_21645,N_23819);
or UO_281 (O_281,N_23072,N_21363);
or UO_282 (O_282,N_24698,N_24640);
and UO_283 (O_283,N_20427,N_24894);
or UO_284 (O_284,N_21046,N_24635);
nand UO_285 (O_285,N_24838,N_23873);
and UO_286 (O_286,N_20881,N_23666);
and UO_287 (O_287,N_24293,N_23498);
nand UO_288 (O_288,N_21210,N_22159);
or UO_289 (O_289,N_22360,N_24342);
and UO_290 (O_290,N_23461,N_22770);
and UO_291 (O_291,N_21726,N_20696);
nand UO_292 (O_292,N_20464,N_22451);
nand UO_293 (O_293,N_20225,N_20885);
or UO_294 (O_294,N_22231,N_22502);
xor UO_295 (O_295,N_23050,N_20426);
xnor UO_296 (O_296,N_20216,N_20312);
and UO_297 (O_297,N_21294,N_21250);
or UO_298 (O_298,N_24937,N_23171);
and UO_299 (O_299,N_21768,N_21173);
or UO_300 (O_300,N_21721,N_24677);
and UO_301 (O_301,N_22321,N_24794);
or UO_302 (O_302,N_23848,N_24189);
nand UO_303 (O_303,N_24118,N_21261);
xor UO_304 (O_304,N_21343,N_24203);
nor UO_305 (O_305,N_20428,N_22611);
or UO_306 (O_306,N_22809,N_22533);
and UO_307 (O_307,N_23321,N_21183);
xnor UO_308 (O_308,N_24903,N_22627);
or UO_309 (O_309,N_21834,N_23169);
or UO_310 (O_310,N_21688,N_23146);
nor UO_311 (O_311,N_22118,N_21619);
and UO_312 (O_312,N_22772,N_23391);
xor UO_313 (O_313,N_24051,N_21426);
xor UO_314 (O_314,N_20948,N_21086);
or UO_315 (O_315,N_22080,N_20327);
nor UO_316 (O_316,N_21697,N_23717);
nor UO_317 (O_317,N_20835,N_23045);
nor UO_318 (O_318,N_23109,N_24167);
nor UO_319 (O_319,N_20822,N_22540);
xnor UO_320 (O_320,N_23642,N_21083);
and UO_321 (O_321,N_23347,N_23235);
xnor UO_322 (O_322,N_23730,N_20580);
and UO_323 (O_323,N_22514,N_22669);
and UO_324 (O_324,N_21566,N_22235);
and UO_325 (O_325,N_24422,N_22391);
and UO_326 (O_326,N_24222,N_20292);
or UO_327 (O_327,N_22163,N_20277);
xor UO_328 (O_328,N_22551,N_23978);
xnor UO_329 (O_329,N_24922,N_22542);
nand UO_330 (O_330,N_20058,N_20722);
or UO_331 (O_331,N_21344,N_23557);
xor UO_332 (O_332,N_22380,N_22608);
xor UO_333 (O_333,N_22267,N_23032);
and UO_334 (O_334,N_24615,N_24042);
nand UO_335 (O_335,N_20753,N_22979);
and UO_336 (O_336,N_21620,N_22322);
and UO_337 (O_337,N_24163,N_21845);
or UO_338 (O_338,N_20392,N_24153);
nand UO_339 (O_339,N_24668,N_23910);
and UO_340 (O_340,N_24066,N_24476);
nand UO_341 (O_341,N_23180,N_22161);
nor UO_342 (O_342,N_23775,N_24994);
nor UO_343 (O_343,N_23054,N_24987);
or UO_344 (O_344,N_23904,N_21736);
nand UO_345 (O_345,N_24696,N_20780);
nor UO_346 (O_346,N_21403,N_21109);
xor UO_347 (O_347,N_22845,N_23995);
and UO_348 (O_348,N_24578,N_21098);
xnor UO_349 (O_349,N_21865,N_24159);
and UO_350 (O_350,N_22573,N_22702);
nor UO_351 (O_351,N_20564,N_22644);
nor UO_352 (O_352,N_21454,N_22754);
or UO_353 (O_353,N_20576,N_24502);
nand UO_354 (O_354,N_23603,N_20941);
nand UO_355 (O_355,N_20670,N_24393);
xnor UO_356 (O_356,N_24046,N_23671);
or UO_357 (O_357,N_22496,N_20196);
and UO_358 (O_358,N_22142,N_22106);
or UO_359 (O_359,N_24955,N_20799);
and UO_360 (O_360,N_24095,N_24478);
and UO_361 (O_361,N_21996,N_24127);
nor UO_362 (O_362,N_20301,N_22057);
xor UO_363 (O_363,N_21552,N_22976);
or UO_364 (O_364,N_23165,N_23966);
xnor UO_365 (O_365,N_24917,N_20107);
nor UO_366 (O_366,N_20313,N_23365);
xor UO_367 (O_367,N_24763,N_21871);
nor UO_368 (O_368,N_21473,N_24641);
and UO_369 (O_369,N_20724,N_20820);
and UO_370 (O_370,N_24769,N_24629);
xnor UO_371 (O_371,N_22585,N_21565);
and UO_372 (O_372,N_20199,N_20589);
xor UO_373 (O_373,N_20610,N_22332);
and UO_374 (O_374,N_22749,N_23532);
and UO_375 (O_375,N_20035,N_22659);
nor UO_376 (O_376,N_23475,N_20429);
or UO_377 (O_377,N_23691,N_22671);
nor UO_378 (O_378,N_23299,N_22790);
xor UO_379 (O_379,N_21185,N_24397);
or UO_380 (O_380,N_20678,N_23203);
nand UO_381 (O_381,N_20559,N_20029);
and UO_382 (O_382,N_20934,N_20072);
and UO_383 (O_383,N_20166,N_20513);
xnor UO_384 (O_384,N_23415,N_24693);
nand UO_385 (O_385,N_20446,N_20228);
xor UO_386 (O_386,N_23196,N_22424);
xor UO_387 (O_387,N_23473,N_24656);
nor UO_388 (O_388,N_20011,N_23315);
nor UO_389 (O_389,N_23629,N_23309);
and UO_390 (O_390,N_23055,N_21206);
xor UO_391 (O_391,N_24958,N_23341);
or UO_392 (O_392,N_24403,N_24827);
or UO_393 (O_393,N_20578,N_24398);
or UO_394 (O_394,N_21848,N_22794);
xor UO_395 (O_395,N_20495,N_22884);
nor UO_396 (O_396,N_20575,N_22516);
or UO_397 (O_397,N_21887,N_23120);
nor UO_398 (O_398,N_20679,N_22647);
or UO_399 (O_399,N_22276,N_20154);
or UO_400 (O_400,N_24910,N_22355);
and UO_401 (O_401,N_24003,N_22971);
xnor UO_402 (O_402,N_22397,N_24250);
and UO_403 (O_403,N_24627,N_21190);
xor UO_404 (O_404,N_20062,N_20791);
or UO_405 (O_405,N_22549,N_21822);
or UO_406 (O_406,N_22003,N_23928);
xor UO_407 (O_407,N_24520,N_22984);
nand UO_408 (O_408,N_20986,N_24811);
nand UO_409 (O_409,N_24564,N_24420);
and UO_410 (O_410,N_21600,N_20527);
or UO_411 (O_411,N_21789,N_20958);
nor UO_412 (O_412,N_20116,N_23593);
xnor UO_413 (O_413,N_21452,N_23571);
and UO_414 (O_414,N_22122,N_23046);
xnor UO_415 (O_415,N_22615,N_22927);
nand UO_416 (O_416,N_23484,N_21609);
nand UO_417 (O_417,N_24591,N_24198);
nor UO_418 (O_418,N_20615,N_24957);
or UO_419 (O_419,N_23148,N_23121);
or UO_420 (O_420,N_23939,N_21877);
and UO_421 (O_421,N_22413,N_24898);
or UO_422 (O_422,N_24268,N_22505);
or UO_423 (O_423,N_20565,N_21612);
xnor UO_424 (O_424,N_24626,N_24733);
xnor UO_425 (O_425,N_24357,N_22762);
and UO_426 (O_426,N_21500,N_20984);
xor UO_427 (O_427,N_23869,N_21347);
and UO_428 (O_428,N_21443,N_22193);
xnor UO_429 (O_429,N_21488,N_20105);
xor UO_430 (O_430,N_23016,N_22715);
or UO_431 (O_431,N_21260,N_20498);
and UO_432 (O_432,N_23175,N_24884);
or UO_433 (O_433,N_24784,N_23678);
or UO_434 (O_434,N_23034,N_20544);
or UO_435 (O_435,N_23736,N_21584);
or UO_436 (O_436,N_20725,N_21802);
nand UO_437 (O_437,N_23703,N_20102);
and UO_438 (O_438,N_21149,N_21796);
nand UO_439 (O_439,N_21636,N_22567);
and UO_440 (O_440,N_22070,N_20369);
and UO_441 (O_441,N_21825,N_23223);
nor UO_442 (O_442,N_23417,N_21487);
nor UO_443 (O_443,N_24888,N_23464);
xor UO_444 (O_444,N_22359,N_24447);
nand UO_445 (O_445,N_21263,N_23424);
or UO_446 (O_446,N_22830,N_22782);
nand UO_447 (O_447,N_23560,N_20066);
or UO_448 (O_448,N_20450,N_23709);
xor UO_449 (O_449,N_21331,N_20612);
xnor UO_450 (O_450,N_23349,N_24325);
nor UO_451 (O_451,N_21017,N_24833);
nand UO_452 (O_452,N_21880,N_21942);
nand UO_453 (O_453,N_22390,N_20730);
or UO_454 (O_454,N_20337,N_24686);
xnor UO_455 (O_455,N_21042,N_24122);
nand UO_456 (O_456,N_20316,N_24251);
nor UO_457 (O_457,N_23123,N_23828);
xor UO_458 (O_458,N_20447,N_22067);
and UO_459 (O_459,N_20229,N_22019);
and UO_460 (O_460,N_22385,N_23757);
nand UO_461 (O_461,N_24773,N_21523);
nand UO_462 (O_462,N_23047,N_20242);
xnor UO_463 (O_463,N_20088,N_22089);
and UO_464 (O_464,N_22895,N_24288);
or UO_465 (O_465,N_23433,N_20604);
and UO_466 (O_466,N_21237,N_21777);
and UO_467 (O_467,N_22428,N_23019);
xnor UO_468 (O_468,N_21513,N_24700);
xnor UO_469 (O_469,N_23961,N_23488);
xor UO_470 (O_470,N_20410,N_23902);
or UO_471 (O_471,N_21976,N_21195);
nor UO_472 (O_472,N_20482,N_24923);
nand UO_473 (O_473,N_23956,N_21815);
nor UO_474 (O_474,N_23481,N_24642);
and UO_475 (O_475,N_21073,N_20960);
xor UO_476 (O_476,N_24558,N_21009);
nor UO_477 (O_477,N_22743,N_23777);
nor UO_478 (O_478,N_21447,N_21159);
or UO_479 (O_479,N_22723,N_20664);
nor UO_480 (O_480,N_21072,N_23036);
and UO_481 (O_481,N_20860,N_20600);
xor UO_482 (O_482,N_20371,N_23364);
nand UO_483 (O_483,N_22662,N_21468);
nand UO_484 (O_484,N_23716,N_21230);
nor UO_485 (O_485,N_22587,N_24532);
or UO_486 (O_486,N_24916,N_21258);
nor UO_487 (O_487,N_24862,N_23547);
nor UO_488 (O_488,N_23168,N_22677);
nor UO_489 (O_489,N_22954,N_20086);
nor UO_490 (O_490,N_20218,N_24680);
nor UO_491 (O_491,N_22960,N_21988);
xor UO_492 (O_492,N_20833,N_21607);
and UO_493 (O_493,N_20748,N_23506);
nand UO_494 (O_494,N_20334,N_24941);
and UO_495 (O_495,N_22568,N_24966);
xnor UO_496 (O_496,N_22599,N_22041);
and UO_497 (O_497,N_24756,N_22883);
and UO_498 (O_498,N_20406,N_24395);
nand UO_499 (O_499,N_20391,N_23494);
xnor UO_500 (O_500,N_24782,N_23903);
nand UO_501 (O_501,N_20048,N_21783);
or UO_502 (O_502,N_21686,N_22733);
and UO_503 (O_503,N_24765,N_20843);
or UO_504 (O_504,N_21643,N_23082);
or UO_505 (O_505,N_22249,N_21549);
xnor UO_506 (O_506,N_20004,N_22510);
xnor UO_507 (O_507,N_21164,N_22526);
xnor UO_508 (O_508,N_24071,N_24147);
nand UO_509 (O_509,N_21656,N_21662);
or UO_510 (O_510,N_24820,N_24551);
xor UO_511 (O_511,N_22784,N_21563);
and UO_512 (O_512,N_24676,N_20466);
nor UO_513 (O_513,N_22443,N_21466);
xor UO_514 (O_514,N_21559,N_22074);
xor UO_515 (O_515,N_24452,N_22961);
nor UO_516 (O_516,N_24535,N_20992);
and UO_517 (O_517,N_21359,N_22925);
xor UO_518 (O_518,N_20682,N_23035);
nand UO_519 (O_519,N_23285,N_20266);
nor UO_520 (O_520,N_24942,N_22777);
or UO_521 (O_521,N_22233,N_22801);
nand UO_522 (O_522,N_21291,N_24370);
xor UO_523 (O_523,N_23888,N_21695);
nand UO_524 (O_524,N_22641,N_22799);
or UO_525 (O_525,N_21310,N_24705);
xnor UO_526 (O_526,N_22223,N_20981);
xnor UO_527 (O_527,N_23437,N_22366);
nand UO_528 (O_528,N_23291,N_24992);
or UO_529 (O_529,N_23040,N_24570);
and UO_530 (O_530,N_21629,N_20632);
and UO_531 (O_531,N_23849,N_20894);
or UO_532 (O_532,N_22315,N_21307);
nand UO_533 (O_533,N_22192,N_24825);
nand UO_534 (O_534,N_20403,N_23030);
nor UO_535 (O_535,N_21071,N_21006);
or UO_536 (O_536,N_20452,N_23114);
nand UO_537 (O_537,N_24116,N_20117);
nor UO_538 (O_538,N_21535,N_24237);
or UO_539 (O_539,N_24045,N_20906);
or UO_540 (O_540,N_22508,N_21255);
xnor UO_541 (O_541,N_24526,N_20430);
nand UO_542 (O_542,N_20461,N_21215);
nor UO_543 (O_543,N_23393,N_24841);
or UO_544 (O_544,N_20603,N_24734);
nand UO_545 (O_545,N_22236,N_24895);
or UO_546 (O_546,N_24160,N_24664);
or UO_547 (O_547,N_20852,N_24780);
nor UO_548 (O_548,N_21642,N_20869);
nor UO_549 (O_549,N_22968,N_21091);
xnor UO_550 (O_550,N_24653,N_24377);
and UO_551 (O_551,N_22054,N_22406);
nor UO_552 (O_552,N_21278,N_23384);
xnor UO_553 (O_553,N_21855,N_20212);
nand UO_554 (O_554,N_24651,N_22268);
or UO_555 (O_555,N_21445,N_21501);
and UO_556 (O_556,N_23001,N_23833);
or UO_557 (O_557,N_23962,N_24628);
nand UO_558 (O_558,N_22763,N_20596);
and UO_559 (O_559,N_20462,N_24356);
or UO_560 (O_560,N_21193,N_20930);
nand UO_561 (O_561,N_21076,N_20059);
nand UO_562 (O_562,N_20622,N_21891);
nor UO_563 (O_563,N_22907,N_23343);
or UO_564 (O_564,N_22273,N_21345);
nand UO_565 (O_565,N_21064,N_24823);
nor UO_566 (O_566,N_23859,N_23278);
xnor UO_567 (O_567,N_20157,N_24201);
and UO_568 (O_568,N_22725,N_22950);
or UO_569 (O_569,N_23702,N_22622);
nand UO_570 (O_570,N_23954,N_21872);
xor UO_571 (O_571,N_24097,N_22745);
xnor UO_572 (O_572,N_22822,N_23658);
and UO_573 (O_573,N_23097,N_20716);
xor UO_574 (O_574,N_24857,N_22708);
nand UO_575 (O_575,N_20911,N_24266);
or UO_576 (O_576,N_21264,N_20647);
nor UO_577 (O_577,N_20271,N_24960);
nor UO_578 (O_578,N_22281,N_23483);
or UO_579 (O_579,N_20453,N_22561);
nand UO_580 (O_580,N_21423,N_20840);
or UO_581 (O_581,N_21846,N_24021);
and UO_582 (O_582,N_22471,N_24145);
nor UO_583 (O_583,N_23081,N_20142);
nor UO_584 (O_584,N_21806,N_23261);
or UO_585 (O_585,N_23871,N_20508);
xnor UO_586 (O_586,N_23276,N_24285);
nand UO_587 (O_587,N_21306,N_24757);
nor UO_588 (O_588,N_21987,N_20702);
nor UO_589 (O_589,N_24971,N_23955);
or UO_590 (O_590,N_24086,N_21569);
xor UO_591 (O_591,N_22726,N_22747);
and UO_592 (O_592,N_22867,N_24432);
nand UO_593 (O_593,N_20892,N_22264);
xor UO_594 (O_594,N_22361,N_23916);
and UO_595 (O_595,N_23632,N_23606);
nand UO_596 (O_596,N_20005,N_23720);
xor UO_597 (O_597,N_24671,N_22490);
xnor UO_598 (O_598,N_21733,N_24711);
nand UO_599 (O_599,N_23782,N_23354);
nand UO_600 (O_600,N_20187,N_23013);
xnor UO_601 (O_601,N_22750,N_22517);
and UO_602 (O_602,N_21671,N_24737);
nor UO_603 (O_603,N_20942,N_20859);
and UO_604 (O_604,N_23469,N_23446);
nand UO_605 (O_605,N_24495,N_20363);
and UO_606 (O_606,N_23983,N_24294);
nor UO_607 (O_607,N_21554,N_24389);
or UO_608 (O_608,N_22596,N_22803);
nor UO_609 (O_609,N_20248,N_22613);
nor UO_610 (O_610,N_22776,N_21069);
xor UO_611 (O_611,N_22016,N_23808);
xnor UO_612 (O_612,N_22441,N_24953);
or UO_613 (O_613,N_20971,N_23288);
or UO_614 (O_614,N_22491,N_23769);
nor UO_615 (O_615,N_22129,N_24993);
and UO_616 (O_616,N_23124,N_23143);
nor UO_617 (O_617,N_23044,N_22082);
or UO_618 (O_618,N_24496,N_23153);
or UO_619 (O_619,N_23794,N_24312);
xnor UO_620 (O_620,N_23554,N_23352);
xnor UO_621 (O_621,N_24421,N_24062);
nand UO_622 (O_622,N_20937,N_21130);
nor UO_623 (O_623,N_22805,N_20965);
or UO_624 (O_624,N_22580,N_22903);
nand UO_625 (O_625,N_24573,N_21879);
xor UO_626 (O_626,N_23844,N_23300);
or UO_627 (O_627,N_24448,N_24675);
and UO_628 (O_628,N_24028,N_20101);
nand UO_629 (O_629,N_22243,N_20397);
nand UO_630 (O_630,N_21248,N_23329);
xor UO_631 (O_631,N_24379,N_20586);
nor UO_632 (O_632,N_21672,N_24979);
nor UO_633 (O_633,N_20220,N_23511);
and UO_634 (O_634,N_22197,N_22185);
and UO_635 (O_635,N_22373,N_21676);
nand UO_636 (O_636,N_21348,N_23608);
and UO_637 (O_637,N_21265,N_21112);
or UO_638 (O_638,N_22866,N_23057);
or UO_639 (O_639,N_24101,N_24852);
nor UO_640 (O_640,N_20067,N_22085);
or UO_641 (O_641,N_24702,N_20121);
and UO_642 (O_642,N_24039,N_23841);
or UO_643 (O_643,N_21856,N_24774);
and UO_644 (O_644,N_22310,N_21593);
xnor UO_645 (O_645,N_23907,N_23396);
nand UO_646 (O_646,N_24430,N_23420);
xor UO_647 (O_647,N_21958,N_21152);
nor UO_648 (O_648,N_21795,N_20328);
nor UO_649 (O_649,N_21661,N_23867);
and UO_650 (O_650,N_22157,N_20557);
nand UO_651 (O_651,N_22601,N_21510);
or UO_652 (O_652,N_22545,N_21794);
and UO_653 (O_653,N_22078,N_24295);
or UO_654 (O_654,N_23346,N_22429);
and UO_655 (O_655,N_20697,N_23652);
or UO_656 (O_656,N_22712,N_22415);
nor UO_657 (O_657,N_22947,N_22831);
nor UO_658 (O_658,N_23177,N_20714);
and UO_659 (O_659,N_24638,N_20037);
nor UO_660 (O_660,N_23984,N_24866);
nor UO_661 (O_661,N_20421,N_24724);
nor UO_662 (O_662,N_21209,N_24392);
xnor UO_663 (O_663,N_24244,N_20138);
xor UO_664 (O_664,N_20997,N_23017);
or UO_665 (O_665,N_21297,N_22941);
or UO_666 (O_666,N_23783,N_23379);
xor UO_667 (O_667,N_20000,N_20518);
or UO_668 (O_668,N_24681,N_20054);
nor UO_669 (O_669,N_22881,N_24175);
xor UO_670 (O_670,N_23422,N_23875);
and UO_671 (O_671,N_20235,N_20710);
nor UO_672 (O_672,N_21088,N_24310);
and UO_673 (O_673,N_23144,N_20370);
and UO_674 (O_674,N_21705,N_21719);
nor UO_675 (O_675,N_22820,N_23265);
nor UO_676 (O_676,N_20548,N_21304);
nand UO_677 (O_677,N_22792,N_20039);
or UO_678 (O_678,N_22002,N_23683);
nor UO_679 (O_679,N_24845,N_21791);
and UO_680 (O_680,N_21919,N_22987);
xnor UO_681 (O_681,N_20667,N_24501);
or UO_682 (O_682,N_22843,N_24470);
or UO_683 (O_683,N_24119,N_22303);
nand UO_684 (O_684,N_24709,N_20661);
and UO_685 (O_685,N_22476,N_23926);
or UO_686 (O_686,N_23861,N_22638);
nand UO_687 (O_687,N_23412,N_21787);
xor UO_688 (O_688,N_22886,N_20320);
nor UO_689 (O_689,N_20413,N_24776);
xor UO_690 (O_690,N_20283,N_23729);
xnor UO_691 (O_691,N_20517,N_21997);
nand UO_692 (O_692,N_23301,N_22957);
or UO_693 (O_693,N_23170,N_23041);
nor UO_694 (O_694,N_23509,N_23377);
and UO_695 (O_695,N_21460,N_23722);
or UO_696 (O_696,N_22084,N_24414);
or UO_697 (O_697,N_20599,N_22500);
and UO_698 (O_698,N_20849,N_22316);
nor UO_699 (O_699,N_23653,N_24488);
xnor UO_700 (O_700,N_23520,N_22506);
and UO_701 (O_701,N_23373,N_24246);
xor UO_702 (O_702,N_22401,N_21370);
or UO_703 (O_703,N_22675,N_24190);
nor UO_704 (O_704,N_21451,N_22445);
xnor UO_705 (O_705,N_21021,N_23431);
xnor UO_706 (O_706,N_20782,N_24110);
or UO_707 (O_707,N_20550,N_20465);
and UO_708 (O_708,N_23847,N_22394);
and UO_709 (O_709,N_21772,N_20974);
nand UO_710 (O_710,N_21780,N_23476);
xnor UO_711 (O_711,N_23980,N_23460);
xnor UO_712 (O_712,N_20257,N_23711);
and UO_713 (O_713,N_21875,N_24506);
nor UO_714 (O_714,N_20916,N_24208);
nand UO_715 (O_715,N_24058,N_24793);
or UO_716 (O_716,N_21059,N_21830);
nor UO_717 (O_717,N_20323,N_22875);
or UO_718 (O_718,N_23942,N_20893);
or UO_719 (O_719,N_22910,N_23385);
nand UO_720 (O_720,N_24446,N_22470);
nand UO_721 (O_721,N_21015,N_21315);
and UO_722 (O_722,N_23311,N_20870);
nand UO_723 (O_723,N_22478,N_23376);
or UO_724 (O_724,N_20291,N_23245);
or UO_725 (O_725,N_24646,N_20198);
nand UO_726 (O_726,N_22855,N_23274);
or UO_727 (O_727,N_22010,N_21128);
xor UO_728 (O_728,N_21446,N_23135);
xor UO_729 (O_729,N_24851,N_23340);
xor UO_730 (O_730,N_21392,N_23911);
or UO_731 (O_731,N_23187,N_24450);
and UO_732 (O_732,N_23977,N_21024);
nor UO_733 (O_733,N_20648,N_23803);
nor UO_734 (O_734,N_23374,N_24111);
nor UO_735 (O_735,N_20940,N_22826);
xnor UO_736 (O_736,N_24350,N_21354);
or UO_737 (O_737,N_22046,N_20319);
and UO_738 (O_738,N_24547,N_21888);
xor UO_739 (O_739,N_24130,N_22135);
or UO_740 (O_740,N_23269,N_23832);
and UO_741 (O_741,N_24537,N_23156);
and UO_742 (O_742,N_22475,N_24315);
xnor UO_743 (O_743,N_24832,N_22835);
xor UO_744 (O_744,N_22270,N_23793);
nand UO_745 (O_745,N_23512,N_21805);
nor UO_746 (O_746,N_20633,N_24632);
or UO_747 (O_747,N_21147,N_22174);
or UO_748 (O_748,N_20899,N_22612);
nand UO_749 (O_749,N_20970,N_23905);
nand UO_750 (O_750,N_21691,N_21959);
nor UO_751 (O_751,N_21353,N_22848);
or UO_752 (O_752,N_24267,N_22917);
and UO_753 (O_753,N_21937,N_20132);
xnor UO_754 (O_754,N_23132,N_23704);
and UO_755 (O_755,N_24605,N_23686);
xnor UO_756 (O_756,N_22972,N_21203);
nor UO_757 (O_757,N_21229,N_21840);
or UO_758 (O_758,N_22036,N_23870);
nor UO_759 (O_759,N_22464,N_22838);
nor UO_760 (O_760,N_21453,N_24275);
or UO_761 (O_761,N_20902,N_24919);
and UO_762 (O_762,N_22985,N_23216);
nand UO_763 (O_763,N_21932,N_20135);
or UO_764 (O_764,N_20865,N_22351);
or UO_765 (O_765,N_22062,N_20289);
and UO_766 (O_766,N_21730,N_20219);
and UO_767 (O_767,N_23444,N_24707);
and UO_768 (O_768,N_24731,N_21242);
nor UO_769 (O_769,N_20435,N_24215);
xor UO_770 (O_770,N_20476,N_23508);
nand UO_771 (O_771,N_23877,N_22076);
nand UO_772 (O_772,N_23615,N_21222);
or UO_773 (O_773,N_24806,N_24004);
nor UO_774 (O_774,N_20014,N_20922);
or UO_775 (O_775,N_21398,N_20781);
nand UO_776 (O_776,N_23286,N_21043);
nor UO_777 (O_777,N_24074,N_24673);
or UO_778 (O_778,N_21929,N_24819);
nor UO_779 (O_779,N_20139,N_21761);
and UO_780 (O_780,N_20873,N_24808);
or UO_781 (O_781,N_24314,N_24235);
or UO_782 (O_782,N_22635,N_20264);
xnor UO_783 (O_783,N_21005,N_23083);
nor UO_784 (O_784,N_22785,N_23699);
xnor UO_785 (O_785,N_22487,N_22259);
xor UO_786 (O_786,N_24689,N_24459);
nor UO_787 (O_787,N_21476,N_24000);
xor UO_788 (O_788,N_22956,N_23558);
nand UO_789 (O_789,N_23957,N_22603);
and UO_790 (O_790,N_23580,N_23335);
xor UO_791 (O_791,N_21631,N_23898);
and UO_792 (O_792,N_22757,N_20073);
nor UO_793 (O_793,N_20438,N_22744);
nor UO_794 (O_794,N_21166,N_22834);
and UO_795 (O_795,N_22829,N_21225);
or UO_796 (O_796,N_20846,N_22643);
xnor UO_797 (O_797,N_23804,N_22600);
nand UO_798 (O_798,N_22104,N_20170);
nor UO_799 (O_799,N_20272,N_21409);
or UO_800 (O_800,N_20484,N_21666);
xnor UO_801 (O_801,N_24150,N_21421);
xor UO_802 (O_802,N_21725,N_22014);
nand UO_803 (O_803,N_22468,N_21551);
and UO_804 (O_804,N_24892,N_20252);
or UO_805 (O_805,N_21603,N_21982);
nand UO_806 (O_806,N_20020,N_23116);
or UO_807 (O_807,N_22586,N_22543);
and UO_808 (O_808,N_22850,N_23567);
nand UO_809 (O_809,N_24732,N_22579);
or UO_810 (O_810,N_24885,N_20162);
nor UO_811 (O_811,N_23451,N_23967);
xor UO_812 (O_812,N_21270,N_24223);
nand UO_813 (O_813,N_22389,N_22444);
or UO_814 (O_814,N_20912,N_23272);
xor UO_815 (O_815,N_24410,N_23268);
xnor UO_816 (O_816,N_24358,N_22929);
nor UO_817 (O_817,N_21391,N_24157);
xor UO_818 (O_818,N_23403,N_23964);
and UO_819 (O_819,N_23688,N_23392);
xnor UO_820 (O_820,N_24754,N_21859);
nand UO_821 (O_821,N_23800,N_21008);
or UO_822 (O_822,N_20887,N_24109);
and UO_823 (O_823,N_20405,N_24736);
nand UO_824 (O_824,N_23113,N_22165);
nor UO_825 (O_825,N_24248,N_22458);
xnor UO_826 (O_826,N_24141,N_24001);
and UO_827 (O_827,N_24962,N_24382);
nor UO_828 (O_828,N_21681,N_22811);
xor UO_829 (O_829,N_23913,N_20074);
nand UO_830 (O_830,N_24005,N_24492);
nand UO_831 (O_831,N_22371,N_22636);
nor UO_832 (O_832,N_20743,N_24726);
and UO_833 (O_833,N_23564,N_24435);
xor UO_834 (O_834,N_23450,N_20480);
nor UO_835 (O_835,N_24824,N_24844);
and UO_836 (O_836,N_24684,N_21771);
nand UO_837 (O_837,N_22571,N_23470);
and UO_838 (O_838,N_22184,N_22108);
nor UO_839 (O_839,N_20223,N_24997);
and UO_840 (O_840,N_24049,N_21081);
xnor UO_841 (O_841,N_23038,N_21786);
and UO_842 (O_842,N_24316,N_22617);
or UO_843 (O_843,N_20944,N_20929);
and UO_844 (O_844,N_21479,N_24817);
xor UO_845 (O_845,N_20789,N_20030);
xnor UO_846 (O_846,N_24493,N_20536);
or UO_847 (O_847,N_20267,N_24645);
xor UO_848 (O_848,N_23548,N_21575);
or UO_849 (O_849,N_23536,N_20931);
and UO_850 (O_850,N_21196,N_24137);
or UO_851 (O_851,N_21275,N_23383);
or UO_852 (O_852,N_21328,N_22759);
nand UO_853 (O_853,N_24974,N_21991);
or UO_854 (O_854,N_21923,N_21956);
or UO_855 (O_855,N_22846,N_24670);
nor UO_856 (O_856,N_23234,N_24710);
xnor UO_857 (O_857,N_24374,N_24455);
and UO_858 (O_858,N_21868,N_23263);
or UO_859 (O_859,N_21538,N_22336);
nor UO_860 (O_860,N_22583,N_21968);
xnor UO_861 (O_861,N_24572,N_22800);
nand UO_862 (O_862,N_23607,N_24669);
and UO_863 (O_863,N_20635,N_20031);
xnor UO_864 (O_864,N_24727,N_21568);
xnor UO_865 (O_865,N_23233,N_23489);
nor UO_866 (O_866,N_22402,N_24995);
nor UO_867 (O_867,N_22344,N_23786);
nand UO_868 (O_868,N_20918,N_24789);
xnor UO_869 (O_869,N_21927,N_21536);
nand UO_870 (O_870,N_24108,N_24790);
nor UO_871 (O_871,N_22296,N_22050);
nand UO_872 (O_872,N_22285,N_24587);
nand UO_873 (O_873,N_22387,N_21763);
and UO_874 (O_874,N_21346,N_22173);
and UO_875 (O_875,N_21954,N_22710);
or UO_876 (O_876,N_24816,N_22651);
or UO_877 (O_877,N_20923,N_22837);
or UO_878 (O_878,N_21402,N_20091);
nor UO_879 (O_879,N_23694,N_22806);
nor UO_880 (O_880,N_23796,N_21163);
nor UO_881 (O_881,N_22450,N_22483);
or UO_882 (O_882,N_24018,N_23212);
xnor UO_883 (O_883,N_24596,N_21717);
and UO_884 (O_884,N_23122,N_20964);
and UO_885 (O_885,N_21060,N_21150);
nor UO_886 (O_886,N_24804,N_20668);
xnor UO_887 (O_887,N_24242,N_21639);
and UO_888 (O_888,N_23337,N_23356);
nor UO_889 (O_889,N_22731,N_24399);
nand UO_890 (O_890,N_22964,N_22265);
nor UO_891 (O_891,N_21177,N_21300);
nand UO_892 (O_892,N_20018,N_23136);
xor UO_893 (O_893,N_21318,N_21769);
xnor UO_894 (O_894,N_23851,N_23405);
xnor UO_895 (O_895,N_24206,N_23535);
nor UO_896 (O_896,N_20364,N_22575);
xnor UO_897 (O_897,N_21483,N_20206);
nand UO_898 (O_898,N_22928,N_22460);
nor UO_899 (O_899,N_22755,N_20876);
xnor UO_900 (O_900,N_24444,N_24978);
and UO_901 (O_901,N_24930,N_20542);
nand UO_902 (O_902,N_20394,N_21605);
xor UO_903 (O_903,N_22091,N_21170);
xor UO_904 (O_904,N_20879,N_24660);
and UO_905 (O_905,N_23853,N_24454);
or UO_906 (O_906,N_23739,N_20680);
nand UO_907 (O_907,N_20345,N_24351);
xnor UO_908 (O_908,N_20349,N_22597);
or UO_909 (O_909,N_24772,N_20197);
nor UO_910 (O_910,N_22926,N_23999);
xnor UO_911 (O_911,N_21148,N_23881);
and UO_912 (O_912,N_23398,N_23918);
nand UO_913 (O_913,N_21401,N_23202);
nor UO_914 (O_914,N_22756,N_22448);
xnor UO_915 (O_915,N_20767,N_23387);
or UO_916 (O_916,N_21063,N_22630);
and UO_917 (O_917,N_22172,N_24324);
nand UO_918 (O_918,N_24619,N_22427);
or UO_919 (O_919,N_24956,N_22973);
xnor UO_920 (O_920,N_21417,N_24290);
xnor UO_921 (O_921,N_22962,N_20977);
and UO_922 (O_922,N_22292,N_24767);
nor UO_923 (O_923,N_20131,N_23840);
or UO_924 (O_924,N_24796,N_22728);
nor UO_925 (O_925,N_22334,N_22482);
xor UO_926 (O_926,N_23951,N_21180);
xnor UO_927 (O_927,N_21186,N_23302);
and UO_928 (O_928,N_23355,N_22347);
and UO_929 (O_929,N_21007,N_24327);
or UO_930 (O_930,N_21490,N_24777);
xnor UO_931 (O_931,N_21037,N_22877);
and UO_932 (O_932,N_23906,N_22247);
nor UO_933 (O_933,N_21670,N_24803);
and UO_934 (O_934,N_21223,N_21548);
nor UO_935 (O_935,N_23681,N_22556);
xnor UO_936 (O_936,N_24152,N_23490);
xnor UO_937 (O_937,N_21169,N_22673);
or UO_938 (O_938,N_21462,N_23866);
nand UO_939 (O_939,N_24716,N_22631);
nor UO_940 (O_940,N_23496,N_20145);
nor UO_941 (O_941,N_21517,N_21341);
xnor UO_942 (O_942,N_22188,N_21816);
xor UO_943 (O_943,N_21687,N_22095);
nand UO_944 (O_944,N_24440,N_20249);
or UO_945 (O_945,N_22519,N_24087);
nor UO_946 (O_946,N_22375,N_21732);
and UO_947 (O_947,N_20847,N_22363);
and UO_948 (O_948,N_23528,N_23719);
xnor UO_949 (O_949,N_22945,N_24859);
or UO_950 (O_950,N_21082,N_22052);
and UO_951 (O_951,N_22923,N_21033);
or UO_952 (O_952,N_20100,N_21030);
nor UO_953 (O_953,N_20700,N_20915);
and UO_954 (O_954,N_24913,N_21075);
and UO_955 (O_955,N_20007,N_20352);
xnor UO_956 (O_956,N_23160,N_20342);
nor UO_957 (O_957,N_21273,N_22736);
and UO_958 (O_958,N_24394,N_22682);
nor UO_959 (O_959,N_21302,N_21540);
or UO_960 (O_960,N_20260,N_24229);
and UO_961 (O_961,N_21271,N_21917);
nor UO_962 (O_962,N_22199,N_23351);
xnor UO_963 (O_963,N_23790,N_20286);
xor UO_964 (O_964,N_22119,N_21692);
and UO_965 (O_965,N_24561,N_20034);
or UO_966 (O_966,N_22381,N_23798);
or UO_967 (O_967,N_24900,N_20555);
nand UO_968 (O_968,N_22664,N_20404);
nor UO_969 (O_969,N_21004,N_22143);
xnor UO_970 (O_970,N_23432,N_21945);
nor UO_971 (O_971,N_24603,N_20269);
nand UO_972 (O_972,N_20374,N_21448);
nand UO_973 (O_973,N_20384,N_22727);
nor UO_974 (O_974,N_20674,N_20701);
xnor UO_975 (O_975,N_20501,N_20141);
nor UO_976 (O_976,N_23051,N_24523);
nand UO_977 (O_977,N_21863,N_20185);
xnor UO_978 (O_978,N_23936,N_24745);
nor UO_979 (O_979,N_24818,N_24829);
nor UO_980 (O_980,N_20823,N_20848);
and UO_981 (O_981,N_21122,N_21308);
nor UO_982 (O_982,N_21934,N_22333);
or UO_983 (O_983,N_20172,N_23173);
xnor UO_984 (O_984,N_21950,N_23353);
nand UO_985 (O_985,N_20547,N_22075);
and UO_986 (O_986,N_23048,N_23237);
nor UO_987 (O_987,N_21099,N_22819);
or UO_988 (O_988,N_20174,N_21541);
or UO_989 (O_989,N_23619,N_20279);
nand UO_990 (O_990,N_20038,N_20226);
xnor UO_991 (O_991,N_23110,N_22220);
and UO_992 (O_992,N_20980,N_22341);
and UO_993 (O_993,N_24936,N_22027);
nand UO_994 (O_994,N_23421,N_23106);
and UO_995 (O_995,N_21778,N_22299);
nand UO_996 (O_996,N_20900,N_22026);
or UO_997 (O_997,N_23656,N_22195);
nand UO_998 (O_998,N_24183,N_21061);
or UO_999 (O_999,N_22107,N_22694);
or UO_1000 (O_1000,N_24286,N_23884);
or UO_1001 (O_1001,N_22098,N_22015);
nor UO_1002 (O_1002,N_21724,N_20831);
nand UO_1003 (O_1003,N_23779,N_23088);
nand UO_1004 (O_1004,N_22861,N_22072);
and UO_1005 (O_1005,N_24814,N_22320);
nor UO_1006 (O_1006,N_22628,N_24618);
nor UO_1007 (O_1007,N_20772,N_23846);
or UO_1008 (O_1008,N_22241,N_24964);
or UO_1009 (O_1009,N_20768,N_23651);
and UO_1010 (O_1010,N_23574,N_22729);
and UO_1011 (O_1011,N_22840,N_24052);
or UO_1012 (O_1012,N_20002,N_23154);
or UO_1013 (O_1013,N_23005,N_22012);
xnor UO_1014 (O_1014,N_24180,N_21118);
or UO_1015 (O_1015,N_23076,N_23222);
nor UO_1016 (O_1016,N_24217,N_22936);
nand UO_1017 (O_1017,N_24105,N_24322);
xor UO_1018 (O_1018,N_24037,N_24429);
or UO_1019 (O_1019,N_23660,N_22665);
or UO_1020 (O_1020,N_24658,N_23712);
nor UO_1021 (O_1021,N_24475,N_20524);
nand UO_1022 (O_1022,N_24291,N_21482);
and UO_1023 (O_1023,N_22714,N_24270);
xor UO_1024 (O_1024,N_21136,N_21930);
nand UO_1025 (O_1025,N_23084,N_23150);
and UO_1026 (O_1026,N_22064,N_21522);
xnor UO_1027 (O_1027,N_20173,N_22513);
nor UO_1028 (O_1028,N_20080,N_24197);
and UO_1029 (O_1029,N_22548,N_22531);
nand UO_1030 (O_1030,N_23454,N_22824);
nor UO_1031 (O_1031,N_21640,N_23631);
or UO_1032 (O_1032,N_21889,N_22854);
xor UO_1033 (O_1033,N_22206,N_21884);
xnor UO_1034 (O_1034,N_20914,N_23295);
xnor UO_1035 (O_1035,N_20106,N_22088);
xor UO_1036 (O_1036,N_24017,N_23028);
or UO_1037 (O_1037,N_21187,N_24623);
or UO_1038 (O_1038,N_20505,N_21985);
nor UO_1039 (O_1039,N_20735,N_23314);
or UO_1040 (O_1040,N_20396,N_22774);
nor UO_1041 (O_1041,N_22150,N_22225);
or UO_1042 (O_1042,N_22943,N_21947);
nand UO_1043 (O_1043,N_22547,N_20309);
nor UO_1044 (O_1044,N_22481,N_20321);
nor UO_1045 (O_1045,N_20164,N_20795);
xnor UO_1046 (O_1046,N_20263,N_22261);
nor UO_1047 (O_1047,N_23529,N_23795);
nor UO_1048 (O_1048,N_24630,N_23305);
nor UO_1049 (O_1049,N_21394,N_21110);
or UO_1050 (O_1050,N_22377,N_22975);
nand UO_1051 (O_1051,N_20246,N_20936);
or UO_1052 (O_1052,N_22780,N_20570);
or UO_1053 (O_1053,N_22263,N_22833);
xnor UO_1054 (O_1054,N_24542,N_21325);
nand UO_1055 (O_1055,N_21798,N_23900);
nand UO_1056 (O_1056,N_21442,N_20033);
nand UO_1057 (O_1057,N_24424,N_22123);
nand UO_1058 (O_1058,N_22179,N_24697);
nor UO_1059 (O_1059,N_20961,N_23708);
or UO_1060 (O_1060,N_21125,N_21981);
or UO_1061 (O_1061,N_22859,N_21351);
nor UO_1062 (O_1062,N_23492,N_21589);
and UO_1063 (O_1063,N_22836,N_23937);
nand UO_1064 (O_1064,N_20793,N_24549);
and UO_1065 (O_1065,N_22452,N_21003);
xor UO_1066 (O_1066,N_20713,N_23665);
or UO_1067 (O_1067,N_24277,N_22732);
nor UO_1068 (O_1068,N_21703,N_20089);
or UO_1069 (O_1069,N_23940,N_20160);
or UO_1070 (O_1070,N_21895,N_21167);
or UO_1071 (O_1071,N_22528,N_24477);
xor UO_1072 (O_1072,N_23505,N_24985);
or UO_1073 (O_1073,N_23053,N_24531);
or UO_1074 (O_1074,N_20836,N_23159);
xor UO_1075 (O_1075,N_22751,N_21870);
xnor UO_1076 (O_1076,N_22529,N_21457);
xnor UO_1077 (O_1077,N_20122,N_22696);
or UO_1078 (O_1078,N_21545,N_23247);
nor UO_1079 (O_1079,N_23070,N_22949);
nor UO_1080 (O_1080,N_22594,N_23876);
or UO_1081 (O_1081,N_21361,N_20491);
or UO_1082 (O_1082,N_23864,N_20842);
nor UO_1083 (O_1083,N_20618,N_23510);
xnor UO_1084 (O_1084,N_24685,N_24033);
nor UO_1085 (O_1085,N_21883,N_24498);
or UO_1086 (O_1086,N_22403,N_22626);
nor UO_1087 (O_1087,N_21801,N_21980);
nor UO_1088 (O_1088,N_24178,N_23746);
nand UO_1089 (O_1089,N_21365,N_23827);
nand UO_1090 (O_1090,N_20152,N_20744);
and UO_1091 (O_1091,N_21084,N_20515);
or UO_1092 (O_1092,N_20333,N_23590);
nor UO_1093 (O_1093,N_24746,N_21685);
nor UO_1094 (O_1094,N_20400,N_20623);
and UO_1095 (O_1095,N_22934,N_20766);
xnor UO_1096 (O_1096,N_20282,N_23947);
nand UO_1097 (O_1097,N_24881,N_23640);
nor UO_1098 (O_1098,N_21277,N_20693);
or UO_1099 (O_1099,N_22555,N_21139);
and UO_1100 (O_1100,N_20056,N_21623);
xnor UO_1101 (O_1101,N_22619,N_24800);
xor UO_1102 (O_1102,N_20332,N_24289);
nor UO_1103 (O_1103,N_20075,N_21519);
xnor UO_1104 (O_1104,N_21595,N_23836);
and UO_1105 (O_1105,N_20927,N_22748);
and UO_1106 (O_1106,N_23477,N_20758);
and UO_1107 (O_1107,N_24434,N_22417);
or UO_1108 (O_1108,N_21626,N_20706);
or UO_1109 (O_1109,N_24186,N_24038);
nor UO_1110 (O_1110,N_22769,N_22300);
and UO_1111 (O_1111,N_24385,N_24195);
or UO_1112 (O_1112,N_23991,N_22958);
xnor UO_1113 (O_1113,N_23416,N_23990);
and UO_1114 (O_1114,N_20493,N_24593);
nor UO_1115 (O_1115,N_24309,N_22828);
nand UO_1116 (O_1116,N_22983,N_23267);
and UO_1117 (O_1117,N_20012,N_20597);
xnor UO_1118 (O_1118,N_24723,N_21478);
nor UO_1119 (O_1119,N_23397,N_23760);
xnor UO_1120 (O_1120,N_20978,N_24085);
or UO_1121 (O_1121,N_22666,N_24973);
and UO_1122 (O_1122,N_21779,N_22539);
xnor UO_1123 (O_1123,N_20192,N_23003);
nand UO_1124 (O_1124,N_24518,N_20051);
and UO_1125 (O_1125,N_24179,N_23102);
xnor UO_1126 (O_1126,N_21581,N_21531);
xor UO_1127 (O_1127,N_20979,N_24461);
nor UO_1128 (O_1128,N_22812,N_24990);
nand UO_1129 (O_1129,N_23868,N_23588);
and UO_1130 (O_1130,N_20184,N_22564);
or UO_1131 (O_1131,N_22986,N_23208);
nor UO_1132 (O_1132,N_20468,N_23394);
and UO_1133 (O_1133,N_23662,N_23973);
or UO_1134 (O_1134,N_23850,N_21922);
or UO_1135 (O_1135,N_21625,N_22065);
and UO_1136 (O_1136,N_22721,N_21627);
and UO_1137 (O_1137,N_24581,N_24582);
nor UO_1138 (O_1138,N_22590,N_20023);
nand UO_1139 (O_1139,N_21674,N_23569);
and UO_1140 (O_1140,N_21596,N_20314);
and UO_1141 (O_1141,N_22099,N_23033);
nand UO_1142 (O_1142,N_22253,N_22352);
or UO_1143 (O_1143,N_21807,N_21244);
xor UO_1144 (O_1144,N_23131,N_21456);
nand UO_1145 (O_1145,N_24504,N_21679);
nand UO_1146 (O_1146,N_23254,N_23455);
nand UO_1147 (O_1147,N_20568,N_23099);
nor UO_1148 (O_1148,N_24667,N_24830);
nor UO_1149 (O_1149,N_20136,N_21342);
nand UO_1150 (O_1150,N_21129,N_20362);
or UO_1151 (O_1151,N_20828,N_22993);
or UO_1152 (O_1152,N_23667,N_22667);
nand UO_1153 (O_1153,N_21819,N_24034);
xnor UO_1154 (O_1154,N_22852,N_21322);
or UO_1155 (O_1155,N_24172,N_20144);
nor UO_1156 (O_1156,N_23491,N_21918);
nand UO_1157 (O_1157,N_22646,N_21429);
and UO_1158 (O_1158,N_24965,N_24093);
and UO_1159 (O_1159,N_20562,N_22138);
xor UO_1160 (O_1160,N_21866,N_20798);
nand UO_1161 (O_1161,N_23324,N_23814);
xnor UO_1162 (O_1162,N_22128,N_20092);
or UO_1163 (O_1163,N_24517,N_22678);
or UO_1164 (O_1164,N_24113,N_22211);
and UO_1165 (O_1165,N_20433,N_20627);
and UO_1166 (O_1166,N_20663,N_20151);
or UO_1167 (O_1167,N_23893,N_24946);
or UO_1168 (O_1168,N_21664,N_23613);
or UO_1169 (O_1169,N_23400,N_24778);
and UO_1170 (O_1170,N_20356,N_22115);
or UO_1171 (O_1171,N_23262,N_23780);
xor UO_1172 (O_1172,N_20825,N_23430);
and UO_1173 (O_1173,N_21066,N_22537);
nor UO_1174 (O_1174,N_22841,N_21103);
nor UO_1175 (O_1175,N_21389,N_21330);
xor UO_1176 (O_1176,N_22338,N_22416);
xnor UO_1177 (O_1177,N_20455,N_20078);
nor UO_1178 (O_1178,N_21077,N_24012);
or UO_1179 (O_1179,N_21080,N_22037);
xnor UO_1180 (O_1180,N_23008,N_22141);
nor UO_1181 (O_1181,N_24674,N_24546);
or UO_1182 (O_1182,N_21770,N_24088);
nand UO_1183 (O_1183,N_23190,N_23323);
xor UO_1184 (O_1184,N_24343,N_23974);
or UO_1185 (O_1185,N_22025,N_20819);
nand UO_1186 (O_1186,N_21804,N_23698);
nor UO_1187 (O_1187,N_22557,N_22952);
and UO_1188 (O_1188,N_21966,N_20691);
and UO_1189 (O_1189,N_22698,N_24704);
and UO_1190 (O_1190,N_23251,N_22538);
nor UO_1191 (O_1191,N_24353,N_23583);
or UO_1192 (O_1192,N_20205,N_23103);
nand UO_1193 (O_1193,N_20864,N_20777);
xnor UO_1194 (O_1194,N_22872,N_22868);
nand UO_1195 (O_1195,N_21885,N_22996);
nand UO_1196 (O_1196,N_20111,N_24748);
and UO_1197 (O_1197,N_24166,N_20390);
nor UO_1198 (O_1198,N_24560,N_23895);
nor UO_1199 (O_1199,N_23100,N_24148);
and UO_1200 (O_1200,N_20796,N_24788);
nand UO_1201 (O_1201,N_20270,N_22432);
nand UO_1202 (O_1202,N_22396,N_22245);
and UO_1203 (O_1203,N_21108,N_22328);
and UO_1204 (O_1204,N_24969,N_21408);
and UO_1205 (O_1205,N_23338,N_20734);
nor UO_1206 (O_1206,N_20255,N_23727);
and UO_1207 (O_1207,N_24156,N_21858);
or UO_1208 (O_1208,N_22032,N_23467);
xor UO_1209 (O_1209,N_22899,N_21010);
or UO_1210 (O_1210,N_21313,N_22703);
or UO_1211 (O_1211,N_22817,N_24729);
nor UO_1212 (O_1212,N_24725,N_23646);
nand UO_1213 (O_1213,N_22942,N_23378);
or UO_1214 (O_1214,N_23753,N_20913);
nor UO_1215 (O_1215,N_22974,N_20989);
and UO_1216 (O_1216,N_23563,N_24861);
nor UO_1217 (O_1217,N_24339,N_23273);
xnor UO_1218 (O_1218,N_22319,N_24809);
and UO_1219 (O_1219,N_24181,N_20956);
or UO_1220 (O_1220,N_23534,N_23806);
nand UO_1221 (O_1221,N_21874,N_23968);
and UO_1222 (O_1222,N_22499,N_21216);
nor UO_1223 (O_1223,N_22305,N_20497);
nor UO_1224 (O_1224,N_20265,N_21857);
nor UO_1225 (O_1225,N_22145,N_23635);
nor UO_1226 (O_1226,N_20133,N_21054);
nand UO_1227 (O_1227,N_20538,N_22796);
nor UO_1228 (O_1228,N_20488,N_21902);
nor UO_1229 (O_1229,N_21512,N_24075);
and UO_1230 (O_1230,N_22781,N_22204);
nand UO_1231 (O_1231,N_22182,N_21774);
nor UO_1232 (O_1232,N_23112,N_22215);
nor UO_1233 (O_1233,N_23059,N_23682);
nor UO_1234 (O_1234,N_20448,N_23448);
or UO_1235 (O_1235,N_24214,N_24467);
or UO_1236 (O_1236,N_20069,N_22455);
nor UO_1237 (O_1237,N_22312,N_24530);
nor UO_1238 (O_1238,N_21766,N_22607);
nor UO_1239 (O_1239,N_20726,N_23332);
xnor UO_1240 (O_1240,N_20094,N_23086);
nand UO_1241 (O_1241,N_24799,N_24065);
nand UO_1242 (O_1242,N_22255,N_22294);
xnor UO_1243 (O_1243,N_22536,N_22541);
and UO_1244 (O_1244,N_24925,N_23342);
and UO_1245 (O_1245,N_23231,N_23151);
xnor UO_1246 (O_1246,N_20955,N_24426);
nand UO_1247 (O_1247,N_23367,N_21621);
or UO_1248 (O_1248,N_20826,N_20420);
or UO_1249 (O_1249,N_20641,N_23650);
xor UO_1250 (O_1250,N_20998,N_23362);
nand UO_1251 (O_1251,N_23992,N_21124);
nor UO_1252 (O_1252,N_20626,N_23577);
xor UO_1253 (O_1253,N_23501,N_20123);
xnor UO_1254 (O_1254,N_21728,N_22133);
nand UO_1255 (O_1255,N_20380,N_22532);
xor UO_1256 (O_1256,N_23931,N_23654);
or UO_1257 (O_1257,N_24621,N_21594);
and UO_1258 (O_1258,N_23781,N_22383);
xnor UO_1259 (O_1259,N_20821,N_21433);
nor UO_1260 (O_1260,N_20827,N_21924);
nand UO_1261 (O_1261,N_24360,N_23429);
nor UO_1262 (O_1262,N_24607,N_20631);
or UO_1263 (O_1263,N_22660,N_21192);
and UO_1264 (O_1264,N_20326,N_24764);
and UO_1265 (O_1265,N_22331,N_23705);
and UO_1266 (O_1266,N_20177,N_20602);
and UO_1267 (O_1267,N_21963,N_21580);
nor UO_1268 (O_1268,N_24114,N_20169);
and UO_1269 (O_1269,N_22313,N_23715);
nor UO_1270 (O_1270,N_23012,N_24335);
and UO_1271 (O_1271,N_20537,N_23440);
and UO_1272 (O_1272,N_24586,N_20525);
and UO_1273 (O_1273,N_22339,N_23690);
xnor UO_1274 (O_1274,N_22158,N_21386);
nor UO_1275 (O_1275,N_22935,N_20802);
and UO_1276 (O_1276,N_24239,N_21240);
or UO_1277 (O_1277,N_23766,N_20230);
or UO_1278 (O_1278,N_24169,N_22509);
xnor UO_1279 (O_1279,N_24760,N_20108);
or UO_1280 (O_1280,N_23179,N_21537);
xnor UO_1281 (O_1281,N_23334,N_20490);
nor UO_1282 (O_1282,N_22915,N_23225);
and UO_1283 (O_1283,N_22367,N_21957);
and UO_1284 (O_1284,N_22842,N_23889);
nand UO_1285 (O_1285,N_20814,N_22966);
xor UO_1286 (O_1286,N_22808,N_23723);
nor UO_1287 (O_1287,N_21707,N_23009);
xor UO_1288 (O_1288,N_22876,N_23695);
xnor UO_1289 (O_1289,N_21105,N_24624);
xor UO_1290 (O_1290,N_24743,N_20308);
or UO_1291 (O_1291,N_21078,N_22126);
and UO_1292 (O_1292,N_24292,N_22497);
nor UO_1293 (O_1293,N_20797,N_21920);
nand UO_1294 (O_1294,N_24453,N_22190);
and UO_1295 (O_1295,N_22144,N_24436);
nand UO_1296 (O_1296,N_21734,N_21036);
nor UO_1297 (O_1297,N_23541,N_22880);
and UO_1298 (O_1298,N_20140,N_21606);
nor UO_1299 (O_1299,N_20861,N_21381);
nor UO_1300 (O_1300,N_24216,N_23155);
or UO_1301 (O_1301,N_20256,N_24483);
or UO_1302 (O_1302,N_24703,N_23242);
nor UO_1303 (O_1303,N_21539,N_20227);
and UO_1304 (O_1304,N_21750,N_21441);
or UO_1305 (O_1305,N_24303,N_23220);
or UO_1306 (O_1306,N_24199,N_23614);
nand UO_1307 (O_1307,N_24056,N_20719);
nor UO_1308 (O_1308,N_21217,N_21843);
nor UO_1309 (O_1309,N_22577,N_20617);
xnor UO_1310 (O_1310,N_24505,N_22530);
nor UO_1311 (O_1311,N_21765,N_23486);
and UO_1312 (O_1312,N_23419,N_23068);
nand UO_1313 (O_1313,N_23934,N_20611);
nor UO_1314 (O_1314,N_21644,N_23761);
nor UO_1315 (O_1315,N_22569,N_21428);
nor UO_1316 (O_1316,N_20156,N_22918);
and UO_1317 (O_1317,N_21093,N_21660);
and UO_1318 (O_1318,N_20572,N_22507);
nand UO_1319 (O_1319,N_20355,N_21419);
nand UO_1320 (O_1320,N_24129,N_23857);
and UO_1321 (O_1321,N_24032,N_23389);
nand UO_1322 (O_1322,N_20951,N_24610);
nor UO_1323 (O_1323,N_20877,N_22768);
or UO_1324 (O_1324,N_22980,N_21089);
and UO_1325 (O_1325,N_20790,N_24482);
or UO_1326 (O_1326,N_24598,N_24691);
nand UO_1327 (O_1327,N_22127,N_24545);
and UO_1328 (O_1328,N_23229,N_23821);
nand UO_1329 (O_1329,N_24847,N_22120);
or UO_1330 (O_1330,N_22463,N_22024);
xnor UO_1331 (O_1331,N_20966,N_22882);
or UO_1332 (O_1332,N_24387,N_24272);
and UO_1333 (O_1333,N_20574,N_21085);
or UO_1334 (O_1334,N_23933,N_22634);
and UO_1335 (O_1335,N_20511,N_24334);
xnor UO_1336 (O_1336,N_23465,N_21511);
nor UO_1337 (O_1337,N_20377,N_23890);
or UO_1338 (O_1338,N_21878,N_20485);
xnor UO_1339 (O_1339,N_23628,N_23987);
xor UO_1340 (O_1340,N_20924,N_23157);
or UO_1341 (O_1341,N_20921,N_21543);
or UO_1342 (O_1342,N_20437,N_24164);
or UO_1343 (O_1343,N_21743,N_23246);
and UO_1344 (O_1344,N_21904,N_24281);
and UO_1345 (O_1345,N_23685,N_20582);
and UO_1346 (O_1346,N_23661,N_24359);
and UO_1347 (O_1347,N_20839,N_20359);
and UO_1348 (O_1348,N_23572,N_23787);
and UO_1349 (O_1349,N_21586,N_23517);
nor UO_1350 (O_1350,N_24507,N_22147);
nor UO_1351 (O_1351,N_23283,N_23919);
nor UO_1352 (O_1352,N_21809,N_21901);
nor UO_1353 (O_1353,N_24173,N_20884);
or UO_1354 (O_1354,N_23537,N_22480);
xnor UO_1355 (O_1355,N_23927,N_21373);
xnor UO_1356 (O_1356,N_23912,N_23310);
nor UO_1357 (O_1357,N_21546,N_23408);
nand UO_1358 (O_1358,N_23252,N_22709);
or UO_1359 (O_1359,N_21272,N_22202);
nand UO_1360 (O_1360,N_23676,N_21738);
xor UO_1361 (O_1361,N_23217,N_20529);
nor UO_1362 (O_1362,N_24009,N_23294);
and UO_1363 (O_1363,N_24500,N_22939);
xnor UO_1364 (O_1364,N_21591,N_22071);
nand UO_1365 (O_1365,N_22849,N_20245);
nand UO_1366 (O_1366,N_23858,N_23042);
nor UO_1367 (O_1367,N_23238,N_23915);
or UO_1368 (O_1368,N_22595,N_24055);
or UO_1369 (O_1369,N_24721,N_21913);
or UO_1370 (O_1370,N_23345,N_24104);
nand UO_1371 (O_1371,N_24228,N_22183);
nand UO_1372 (O_1372,N_20815,N_22093);
nand UO_1373 (O_1373,N_23950,N_21788);
and UO_1374 (O_1374,N_24151,N_20530);
nor UO_1375 (O_1375,N_21058,N_22092);
and UO_1376 (O_1376,N_23172,N_20521);
nand UO_1377 (O_1377,N_21145,N_20556);
xnor UO_1378 (O_1378,N_20167,N_22198);
or UO_1379 (O_1379,N_20302,N_21556);
xor UO_1380 (O_1380,N_22815,N_22283);
and UO_1381 (O_1381,N_22008,N_21742);
nand UO_1382 (O_1382,N_23623,N_21931);
and UO_1383 (O_1383,N_22214,N_24302);
and UO_1384 (O_1384,N_22898,N_23561);
nand UO_1385 (O_1385,N_24384,N_23474);
and UO_1386 (O_1386,N_22906,N_22827);
xnor UO_1387 (O_1387,N_22574,N_20047);
nor UO_1388 (O_1388,N_23007,N_22293);
and UO_1389 (O_1389,N_24245,N_23449);
and UO_1390 (O_1390,N_22683,N_20408);
nand UO_1391 (O_1391,N_20171,N_21599);
nor UO_1392 (O_1392,N_21420,N_20898);
nor UO_1393 (O_1393,N_21201,N_20458);
or UO_1394 (O_1394,N_22151,N_23200);
nand UO_1395 (O_1395,N_21465,N_21301);
xor UO_1396 (O_1396,N_23207,N_23117);
xor UO_1397 (O_1397,N_24134,N_20608);
nor UO_1398 (O_1398,N_22937,N_22798);
or UO_1399 (O_1399,N_23952,N_23773);
nand UO_1400 (O_1400,N_24868,N_23768);
nand UO_1401 (O_1401,N_22180,N_22314);
or UO_1402 (O_1402,N_24924,N_23181);
or UO_1403 (O_1403,N_20813,N_23330);
nand UO_1404 (O_1404,N_22581,N_20699);
or UO_1405 (O_1405,N_21851,N_23791);
or UO_1406 (O_1406,N_21792,N_20129);
and UO_1407 (O_1407,N_24230,N_20358);
xor UO_1408 (O_1408,N_22090,N_21847);
nor UO_1409 (O_1409,N_24301,N_22372);
nor UO_1410 (O_1410,N_23885,N_20975);
and UO_1411 (O_1411,N_21906,N_21867);
nand UO_1412 (O_1412,N_21214,N_24943);
or UO_1413 (O_1413,N_20686,N_22287);
or UO_1414 (O_1414,N_20963,N_22086);
xnor UO_1415 (O_1415,N_20595,N_21663);
nor UO_1416 (O_1416,N_21507,N_23069);
nor UO_1417 (O_1417,N_21698,N_24932);
nand UO_1418 (O_1418,N_22269,N_23407);
nand UO_1419 (O_1419,N_23731,N_23570);
xor UO_1420 (O_1420,N_21137,N_21279);
nand UO_1421 (O_1421,N_20844,N_23210);
xnor UO_1422 (O_1422,N_22365,N_23549);
or UO_1423 (O_1423,N_23257,N_22649);
nor UO_1424 (O_1424,N_21735,N_21757);
and UO_1425 (O_1425,N_21281,N_22693);
or UO_1426 (O_1426,N_23270,N_24752);
and UO_1427 (O_1427,N_24040,N_22166);
nand UO_1428 (O_1428,N_21094,N_20019);
xnor UO_1429 (O_1429,N_21289,N_24311);
nor UO_1430 (O_1430,N_21570,N_22278);
and UO_1431 (O_1431,N_24836,N_23369);
xor UO_1432 (O_1432,N_20261,N_20317);
nor UO_1433 (O_1433,N_21387,N_20168);
xor UO_1434 (O_1434,N_22252,N_20816);
or UO_1435 (O_1435,N_23192,N_21040);
and UO_1436 (O_1436,N_21477,N_22222);
nor UO_1437 (O_1437,N_24657,N_24368);
or UO_1438 (O_1438,N_20475,N_20209);
nor UO_1439 (O_1439,N_24257,N_21284);
or UO_1440 (O_1440,N_21184,N_21582);
or UO_1441 (O_1441,N_20306,N_20784);
xor UO_1442 (O_1442,N_20741,N_20967);
nand UO_1443 (O_1443,N_22254,N_24123);
xnor UO_1444 (O_1444,N_22672,N_23184);
nand UO_1445 (O_1445,N_24014,N_20910);
or UO_1446 (O_1446,N_22177,N_23145);
nand UO_1447 (O_1447,N_22602,N_21762);
nor UO_1448 (O_1448,N_20901,N_24579);
nor UO_1449 (O_1449,N_20375,N_21493);
nand UO_1450 (O_1450,N_20330,N_23586);
or UO_1451 (O_1451,N_22862,N_22559);
xnor UO_1452 (O_1452,N_23079,N_23372);
and UO_1453 (O_1453,N_24536,N_20275);
nor UO_1454 (O_1454,N_23899,N_24655);
xnor UO_1455 (O_1455,N_21175,N_20211);
xnor UO_1456 (O_1456,N_24613,N_22655);
and UO_1457 (O_1457,N_22081,N_24340);
xnor UO_1458 (O_1458,N_21470,N_24758);
or UO_1459 (O_1459,N_23186,N_21316);
nand UO_1460 (O_1460,N_21893,N_24849);
or UO_1461 (O_1461,N_21909,N_24439);
xnor UO_1462 (O_1462,N_23767,N_23350);
nand UO_1463 (O_1463,N_24365,N_24487);
xnor UO_1464 (O_1464,N_20746,N_24149);
nand UO_1465 (O_1465,N_24945,N_24699);
and UO_1466 (O_1466,N_24486,N_23971);
xor UO_1467 (O_1467,N_22716,N_23860);
and UO_1468 (O_1468,N_21020,N_21153);
xor UO_1469 (O_1469,N_22357,N_22111);
xor UO_1470 (O_1470,N_21231,N_20001);
or UO_1471 (O_1471,N_20727,N_22226);
xnor UO_1472 (O_1472,N_20566,N_24372);
nand UO_1473 (O_1473,N_21057,N_21041);
nor UO_1474 (O_1474,N_24271,N_24649);
nor UO_1475 (O_1475,N_20373,N_20551);
nor UO_1476 (O_1476,N_21526,N_21693);
nor UO_1477 (O_1477,N_24443,N_24795);
nor UO_1478 (O_1478,N_23896,N_23095);
nor UO_1479 (O_1479,N_23706,N_21677);
nor UO_1480 (O_1480,N_20176,N_20329);
or UO_1481 (O_1481,N_22512,N_20659);
nor UO_1482 (O_1482,N_20065,N_24759);
xnor UO_1483 (O_1483,N_21873,N_24427);
nor UO_1484 (O_1484,N_21745,N_20628);
nand UO_1485 (O_1485,N_20987,N_24950);
nand UO_1486 (O_1486,N_21235,N_24094);
or UO_1487 (O_1487,N_22904,N_24751);
and UO_1488 (O_1488,N_20469,N_24874);
nand UO_1489 (O_1489,N_20988,N_23049);
or UO_1490 (O_1490,N_24209,N_23713);
or UO_1491 (O_1491,N_21749,N_20411);
and UO_1492 (O_1492,N_24090,N_23975);
nand UO_1493 (O_1493,N_20017,N_22870);
xor UO_1494 (O_1494,N_24469,N_22456);
nor UO_1495 (O_1495,N_22688,N_21650);
nor UO_1496 (O_1496,N_20803,N_20295);
nand UO_1497 (O_1497,N_23240,N_22606);
or UO_1498 (O_1498,N_23025,N_23576);
nor UO_1499 (O_1499,N_22399,N_21276);
nand UO_1500 (O_1500,N_20801,N_20210);
and UO_1501 (O_1501,N_22653,N_20381);
and UO_1502 (O_1502,N_22582,N_24355);
nand UO_1503 (O_1503,N_21369,N_22982);
and UO_1504 (O_1504,N_23163,N_21355);
nor UO_1505 (O_1505,N_23457,N_21494);
nor UO_1506 (O_1506,N_24606,N_22061);
nand UO_1507 (O_1507,N_24952,N_20854);
nand UO_1508 (O_1508,N_20983,N_21413);
nand UO_1509 (O_1509,N_24636,N_23663);
nand UO_1510 (O_1510,N_21529,N_21828);
xnor UO_1511 (O_1511,N_23770,N_24253);
and UO_1512 (O_1512,N_23174,N_23809);
and UO_1513 (O_1513,N_21135,N_20287);
nand UO_1514 (O_1514,N_21577,N_20897);
xor UO_1515 (O_1515,N_20858,N_20351);
nor UO_1516 (O_1516,N_21269,N_23255);
and UO_1517 (O_1517,N_20516,N_23322);
and UO_1518 (O_1518,N_24837,N_23948);
nand UO_1519 (O_1519,N_20418,N_21349);
and UO_1520 (O_1520,N_23162,N_21505);
or UO_1521 (O_1521,N_23630,N_22946);
xor UO_1522 (O_1522,N_24577,N_24712);
nor UO_1523 (O_1523,N_21305,N_21329);
or UO_1524 (O_1524,N_21869,N_23645);
xor UO_1525 (O_1525,N_21323,N_24863);
nand UO_1526 (O_1526,N_23260,N_21256);
and UO_1527 (O_1527,N_23230,N_21374);
xnor UO_1528 (O_1528,N_21023,N_21925);
nor UO_1529 (O_1529,N_24747,N_20208);
nor UO_1530 (O_1530,N_23579,N_22368);
xnor UO_1531 (O_1531,N_20990,N_20830);
xnor UO_1532 (O_1532,N_21132,N_21835);
nand UO_1533 (O_1533,N_21027,N_20189);
nand UO_1534 (O_1534,N_24264,N_20591);
xnor UO_1535 (O_1535,N_22645,N_21611);
or UO_1536 (O_1536,N_24931,N_21303);
nor UO_1537 (O_1537,N_21106,N_24328);
or UO_1538 (O_1538,N_22189,N_20889);
xor UO_1539 (O_1539,N_23929,N_23585);
nor UO_1540 (O_1540,N_23891,N_22614);
and UO_1541 (O_1541,N_22056,N_20439);
nor UO_1542 (O_1542,N_22216,N_21534);
nand UO_1543 (O_1543,N_24976,N_20721);
xor UO_1544 (O_1544,N_23513,N_24364);
nor UO_1545 (O_1545,N_21808,N_24583);
or UO_1546 (O_1546,N_20424,N_21882);
xor UO_1547 (O_1547,N_20868,N_20543);
nand UO_1548 (O_1548,N_22467,N_24260);
nand UO_1549 (O_1549,N_20445,N_21045);
and UO_1550 (O_1550,N_24708,N_20650);
nor UO_1551 (O_1551,N_20347,N_20360);
or UO_1552 (O_1552,N_22105,N_20006);
or UO_1553 (O_1553,N_21508,N_22408);
and UO_1554 (O_1554,N_20250,N_23239);
and UO_1555 (O_1555,N_24485,N_20239);
and UO_1556 (O_1556,N_21034,N_22797);
nor UO_1557 (O_1557,N_22418,N_20190);
or UO_1558 (O_1558,N_20620,N_23601);
nor UO_1559 (O_1559,N_22650,N_21327);
or UO_1560 (O_1560,N_24801,N_23924);
nand UO_1561 (O_1561,N_22035,N_20658);
nand UO_1562 (O_1562,N_20280,N_23725);
and UO_1563 (O_1563,N_23183,N_23788);
xnor UO_1564 (O_1564,N_24574,N_23519);
nand UO_1565 (O_1565,N_24694,N_23178);
xnor UO_1566 (O_1566,N_20506,N_22386);
nor UO_1567 (O_1567,N_20052,N_24840);
nor UO_1568 (O_1568,N_23456,N_21321);
or UO_1569 (O_1569,N_23339,N_20103);
or UO_1570 (O_1570,N_20773,N_20425);
xor UO_1571 (O_1571,N_22722,N_20837);
nand UO_1572 (O_1572,N_20731,N_22325);
nand UO_1573 (O_1573,N_20348,N_24225);
or UO_1574 (O_1574,N_22023,N_24786);
and UO_1575 (O_1575,N_24720,N_21911);
xnor UO_1576 (O_1576,N_21912,N_23638);
or UO_1577 (O_1577,N_24276,N_24652);
nand UO_1578 (O_1578,N_23282,N_20717);
xor UO_1579 (O_1579,N_20523,N_23604);
nand UO_1580 (O_1580,N_22724,N_23060);
xnor UO_1581 (O_1581,N_21992,N_24456);
nand UO_1582 (O_1582,N_21022,N_21773);
nand UO_1583 (O_1583,N_23718,N_24247);
xor UO_1584 (O_1584,N_23985,N_20315);
or UO_1585 (O_1585,N_24298,N_24807);
nor UO_1586 (O_1586,N_21019,N_22302);
nand UO_1587 (O_1587,N_22083,N_23318);
xor UO_1588 (O_1588,N_24438,N_23466);
xor UO_1589 (O_1589,N_21812,N_22663);
or UO_1590 (O_1590,N_20382,N_23197);
nand UO_1591 (O_1591,N_21516,N_22767);
and UO_1592 (O_1592,N_23644,N_20593);
nand UO_1593 (O_1593,N_22187,N_23074);
nor UO_1594 (O_1594,N_22425,N_24465);
or UO_1595 (O_1595,N_24867,N_20507);
xor UO_1596 (O_1596,N_23829,N_22260);
nor UO_1597 (O_1597,N_21434,N_24078);
nand UO_1598 (O_1598,N_20994,N_24184);
nor UO_1599 (O_1599,N_24715,N_23308);
nor UO_1600 (O_1600,N_23087,N_20297);
xor UO_1601 (O_1601,N_22349,N_24831);
xnor UO_1602 (O_1602,N_22169,N_21262);
xor UO_1603 (O_1603,N_24255,N_20733);
nand UO_1604 (O_1604,N_22878,N_23887);
nand UO_1605 (O_1605,N_21366,N_20957);
or UO_1606 (O_1606,N_22485,N_23161);
and UO_1607 (O_1607,N_23280,N_21463);
xnor UO_1608 (O_1608,N_22323,N_22753);
nor UO_1609 (O_1609,N_21251,N_24458);
nor UO_1610 (O_1610,N_23410,N_24462);
and UO_1611 (O_1611,N_22625,N_21296);
xnor UO_1612 (O_1612,N_24879,N_23368);
nor UO_1613 (O_1613,N_20646,N_24489);
and UO_1614 (O_1614,N_22864,N_20904);
nand UO_1615 (O_1615,N_24419,N_23227);
xnor UO_1616 (O_1616,N_21011,N_20240);
and UO_1617 (O_1617,N_20563,N_21637);
nand UO_1618 (O_1618,N_24468,N_22488);
nor UO_1619 (O_1619,N_21415,N_24346);
nor UO_1620 (O_1620,N_23004,N_21741);
nand UO_1621 (O_1621,N_23831,N_23426);
nor UO_1622 (O_1622,N_24595,N_22778);
and UO_1623 (O_1623,N_22690,N_22258);
nor UO_1624 (O_1624,N_20150,N_24647);
or UO_1625 (O_1625,N_20120,N_22970);
and UO_1626 (O_1626,N_22297,N_22570);
nor UO_1627 (O_1627,N_24366,N_24269);
nand UO_1628 (O_1628,N_20463,N_21140);
nor UO_1629 (O_1629,N_24265,N_24024);
nand UO_1630 (O_1630,N_24219,N_22149);
and UO_1631 (O_1631,N_23759,N_23599);
and UO_1632 (O_1632,N_24928,N_21266);
and UO_1633 (O_1633,N_23611,N_23096);
xor UO_1634 (O_1634,N_23118,N_20028);
nand UO_1635 (O_1635,N_21211,N_21899);
and UO_1636 (O_1636,N_24566,N_21960);
and UO_1637 (O_1637,N_24631,N_20878);
nor UO_1638 (O_1638,N_22592,N_21101);
xnor UO_1639 (O_1639,N_24409,N_22894);
nand UO_1640 (O_1640,N_21632,N_20124);
nand UO_1641 (O_1641,N_23842,N_22922);
or UO_1642 (O_1642,N_20331,N_21338);
xnor UO_1643 (O_1643,N_22909,N_20222);
or UO_1644 (O_1644,N_24521,N_24300);
xor UO_1645 (O_1645,N_23923,N_24132);
xor UO_1646 (O_1646,N_20389,N_24584);
or UO_1647 (O_1647,N_20273,N_24761);
and UO_1648 (O_1648,N_20754,N_24106);
and UO_1649 (O_1649,N_21416,N_23221);
xnor UO_1650 (O_1650,N_22051,N_21811);
xor UO_1651 (O_1651,N_20440,N_21998);
xor UO_1652 (O_1652,N_21120,N_24442);
nand UO_1653 (O_1653,N_24344,N_23411);
xor UO_1654 (O_1654,N_20594,N_20040);
and UO_1655 (O_1655,N_23427,N_21716);
nand UO_1656 (O_1656,N_21824,N_22398);
and UO_1657 (O_1657,N_24053,N_20514);
nand UO_1658 (O_1658,N_24590,N_24967);
xnor UO_1659 (O_1659,N_24687,N_21979);
nor UO_1660 (O_1660,N_24915,N_21731);
xnor UO_1661 (O_1661,N_21309,N_24534);
nand UO_1662 (O_1662,N_21751,N_21908);
or UO_1663 (O_1663,N_20585,N_21435);
or UO_1664 (O_1664,N_23726,N_20939);
nor UO_1665 (O_1665,N_24232,N_23189);
nor UO_1666 (O_1666,N_20695,N_23166);
and UO_1667 (O_1667,N_21995,N_21243);
xnor UO_1668 (O_1668,N_24977,N_20472);
xor UO_1669 (O_1669,N_24479,N_20690);
and UO_1670 (O_1670,N_21048,N_24020);
nand UO_1671 (O_1671,N_23922,N_22994);
nand UO_1672 (O_1672,N_24690,N_21713);
or UO_1673 (O_1673,N_24352,N_24329);
and UO_1674 (O_1674,N_24103,N_20422);
or UO_1675 (O_1675,N_22897,N_20788);
nand UO_1676 (O_1676,N_24893,N_22550);
or UO_1677 (O_1677,N_20749,N_22889);
xor UO_1678 (O_1678,N_21583,N_24914);
or UO_1679 (O_1679,N_21614,N_24783);
or UO_1680 (O_1680,N_23137,N_24614);
or UO_1681 (O_1681,N_22999,N_23441);
xor UO_1682 (O_1682,N_23472,N_21111);
nand UO_1683 (O_1683,N_23670,N_22309);
nand UO_1684 (O_1684,N_22004,N_24117);
and UO_1685 (O_1685,N_21393,N_23503);
xor UO_1686 (O_1686,N_20624,N_24508);
xnor UO_1687 (O_1687,N_23843,N_21049);
xnor UO_1688 (O_1688,N_20750,N_21364);
or UO_1689 (O_1689,N_20399,N_24401);
xnor UO_1690 (O_1690,N_24280,N_22786);
and UO_1691 (O_1691,N_22358,N_22454);
nand UO_1692 (O_1692,N_20407,N_22821);
nand UO_1693 (O_1693,N_23801,N_23023);
or UO_1694 (O_1694,N_21961,N_22171);
xor UO_1695 (O_1695,N_24473,N_21439);
nand UO_1696 (O_1696,N_24961,N_21896);
nand UO_1697 (O_1697,N_23543,N_23522);
nand UO_1698 (O_1698,N_22738,N_24441);
nand UO_1699 (O_1699,N_24161,N_21684);
xor UO_1700 (O_1700,N_22388,N_22735);
and UO_1701 (O_1701,N_21827,N_22758);
or UO_1702 (O_1702,N_23776,N_21399);
xnor UO_1703 (O_1703,N_20684,N_22043);
nand UO_1704 (O_1704,N_21965,N_22350);
nand UO_1705 (O_1705,N_20552,N_24597);
or UO_1706 (O_1706,N_22364,N_22501);
nor UO_1707 (O_1707,N_21550,N_21553);
nor UO_1708 (O_1708,N_20606,N_21029);
xnor UO_1709 (O_1709,N_24211,N_20412);
or UO_1710 (O_1710,N_24375,N_23284);
or UO_1711 (O_1711,N_23972,N_23482);
nor UO_1712 (O_1712,N_22661,N_24562);
nor UO_1713 (O_1713,N_20494,N_24853);
nor UO_1714 (O_1714,N_22680,N_21823);
nor UO_1715 (O_1715,N_24585,N_22140);
nor UO_1716 (O_1716,N_23856,N_22891);
nand UO_1717 (O_1717,N_22136,N_22609);
nand UO_1718 (O_1718,N_21204,N_22965);
or UO_1719 (O_1719,N_24870,N_22298);
or UO_1720 (O_1720,N_24791,N_23874);
xnor UO_1721 (O_1721,N_23965,N_24527);
xnor UO_1722 (O_1722,N_21864,N_23566);
or UO_1723 (O_1723,N_22021,N_21422);
xnor UO_1724 (O_1724,N_23182,N_23209);
or UO_1725 (O_1725,N_21694,N_21944);
and UO_1726 (O_1726,N_21188,N_24787);
and UO_1727 (O_1727,N_22279,N_20855);
and UO_1728 (O_1728,N_20003,N_23721);
and UO_1729 (O_1729,N_20776,N_24484);
xor UO_1730 (O_1730,N_22047,N_20063);
nand UO_1731 (O_1731,N_24213,N_23595);
and UO_1732 (O_1732,N_22566,N_23232);
nor UO_1733 (O_1733,N_22813,N_20569);
nand UO_1734 (O_1734,N_21051,N_22354);
or UO_1735 (O_1735,N_21117,N_20609);
nand UO_1736 (O_1736,N_23480,N_24999);
nor UO_1737 (O_1737,N_22167,N_20811);
nand UO_1738 (O_1738,N_24839,N_20567);
nor UO_1739 (O_1739,N_24951,N_21935);
xor UO_1740 (O_1740,N_20473,N_23188);
nor UO_1741 (O_1741,N_20759,N_21781);
xnor UO_1742 (O_1742,N_21013,N_20774);
nor UO_1743 (O_1743,N_22955,N_22457);
nor UO_1744 (O_1744,N_24538,N_24404);
nand UO_1745 (O_1745,N_21861,N_20195);
nor UO_1746 (O_1746,N_20294,N_20368);
and UO_1747 (O_1747,N_21972,N_20459);
xnor UO_1748 (O_1748,N_21450,N_20689);
xor UO_1749 (O_1749,N_23733,N_21613);
nor UO_1750 (O_1750,N_20694,N_21168);
xnor UO_1751 (O_1751,N_24073,N_24856);
xnor UO_1752 (O_1752,N_23789,N_20976);
xor UO_1753 (O_1753,N_22244,N_22704);
xor UO_1754 (O_1754,N_24730,N_23093);
or UO_1755 (O_1755,N_20008,N_22218);
or UO_1756 (O_1756,N_24540,N_23741);
xnor UO_1757 (O_1757,N_22791,N_23243);
xnor UO_1758 (O_1758,N_24091,N_21314);
nand UO_1759 (O_1759,N_21371,N_24006);
or UO_1760 (O_1760,N_22598,N_20723);
xnor UO_1761 (O_1761,N_23807,N_24529);
xnor UO_1762 (O_1762,N_21915,N_22832);
or UO_1763 (O_1763,N_23659,N_20945);
nand UO_1764 (O_1764,N_23094,N_21295);
and UO_1765 (O_1765,N_21739,N_22030);
nand UO_1766 (O_1766,N_21096,N_23307);
and UO_1767 (O_1767,N_24491,N_20675);
and UO_1768 (O_1768,N_20845,N_22271);
and UO_1769 (O_1769,N_21668,N_23360);
and UO_1770 (O_1770,N_22902,N_24929);
or UO_1771 (O_1771,N_20296,N_22116);
xor UO_1772 (O_1772,N_20808,N_24047);
xor UO_1773 (O_1773,N_24934,N_23399);
xor UO_1774 (O_1774,N_24411,N_24512);
xor UO_1775 (O_1775,N_22096,N_24077);
and UO_1776 (O_1776,N_22604,N_22430);
and UO_1777 (O_1777,N_22066,N_24154);
xnor UO_1778 (O_1778,N_21990,N_20708);
and UO_1779 (O_1779,N_24361,N_20807);
xor UO_1780 (O_1780,N_22701,N_21767);
nor UO_1781 (O_1781,N_24921,N_24871);
and UO_1782 (O_1782,N_23546,N_23462);
and UO_1783 (O_1783,N_23771,N_23802);
and UO_1784 (O_1784,N_21799,N_24880);
xor UO_1785 (O_1785,N_22814,N_21176);
or UO_1786 (O_1786,N_23471,N_23039);
xnor UO_1787 (O_1787,N_23043,N_20071);
nand UO_1788 (O_1788,N_20969,N_24030);
xor UO_1789 (O_1789,N_24926,N_23752);
nor UO_1790 (O_1790,N_22718,N_24858);
or UO_1791 (O_1791,N_21116,N_22931);
nor UO_1792 (O_1792,N_23882,N_20395);
nand UO_1793 (O_1793,N_20740,N_21234);
xnor UO_1794 (O_1794,N_21833,N_21425);
nor UO_1795 (O_1795,N_24338,N_21286);
xor UO_1796 (O_1796,N_22787,N_24050);
xnor UO_1797 (O_1797,N_23215,N_20926);
and UO_1798 (O_1798,N_24554,N_22393);
nor UO_1799 (O_1799,N_21776,N_24098);
nor UO_1800 (O_1800,N_23562,N_23824);
nor UO_1801 (O_1801,N_23219,N_21634);
nor UO_1802 (O_1802,N_22248,N_20119);
xor UO_1803 (O_1803,N_21897,N_22544);
or UO_1804 (O_1804,N_20386,N_21172);
and UO_1805 (O_1805,N_23140,N_24550);
and UO_1806 (O_1806,N_23091,N_20676);
nand UO_1807 (O_1807,N_24661,N_20718);
nor UO_1808 (O_1808,N_22446,N_23921);
or UO_1809 (O_1809,N_23556,N_23744);
and UO_1810 (O_1810,N_21160,N_22989);
nand UO_1811 (O_1811,N_24717,N_21360);
and UO_1812 (O_1812,N_24539,N_24306);
or UO_1813 (O_1813,N_21890,N_23837);
or UO_1814 (O_1814,N_21119,N_21199);
xor UO_1815 (O_1815,N_22113,N_24509);
and UO_1816 (O_1816,N_24625,N_22584);
xor UO_1817 (O_1817,N_21382,N_21228);
nand UO_1818 (O_1818,N_24332,N_21161);
nor UO_1819 (O_1819,N_20729,N_24541);
nor UO_1820 (O_1820,N_24515,N_20765);
xor UO_1821 (O_1821,N_23015,N_23669);
and UO_1822 (O_1822,N_24821,N_21527);
and UO_1823 (O_1823,N_23575,N_20481);
nand UO_1824 (O_1824,N_22284,N_21760);
and UO_1825 (O_1825,N_24158,N_24896);
xor UO_1826 (O_1826,N_20180,N_22370);
nand UO_1827 (O_1827,N_24802,N_23822);
nand UO_1828 (O_1828,N_21194,N_20298);
nor UO_1829 (O_1829,N_20238,N_24362);
xor UO_1830 (O_1830,N_21213,N_23544);
nor UO_1831 (O_1831,N_22477,N_21268);
and UO_1832 (O_1832,N_20871,N_22462);
or UO_1833 (O_1833,N_23925,N_21320);
or UO_1834 (O_1834,N_22100,N_21949);
nor UO_1835 (O_1835,N_23823,N_24663);
nor UO_1836 (O_1836,N_20993,N_22422);
or UO_1837 (O_1837,N_21638,N_20644);
nor UO_1838 (O_1838,N_20346,N_22439);
xor UO_1839 (O_1839,N_23443,N_21358);
or UO_1840 (O_1840,N_22739,N_22658);
nand UO_1841 (O_1841,N_23609,N_21311);
xnor UO_1842 (O_1842,N_22914,N_21293);
nand UO_1843 (O_1843,N_20224,N_24226);
nand UO_1844 (O_1844,N_24457,N_24433);
xnor UO_1845 (O_1845,N_20113,N_23748);
xnor UO_1846 (O_1846,N_23762,N_23941);
or UO_1847 (O_1847,N_24902,N_22844);
and UO_1848 (O_1848,N_23754,N_22442);
xor UO_1849 (O_1849,N_21989,N_24405);
and UO_1850 (O_1850,N_20276,N_20638);
or UO_1851 (O_1851,N_23089,N_22684);
and UO_1852 (O_1852,N_24654,N_21126);
xnor UO_1853 (O_1853,N_20950,N_24171);
xor UO_1854 (O_1854,N_21601,N_22896);
xor UO_1855 (O_1855,N_21933,N_20738);
xor UO_1856 (O_1856,N_21704,N_23348);
and UO_1857 (O_1857,N_20419,N_23897);
xnor UO_1858 (O_1858,N_24354,N_21179);
or UO_1859 (O_1859,N_24634,N_20571);
or UO_1860 (O_1860,N_23129,N_20581);
or UO_1861 (O_1861,N_21121,N_24373);
nor UO_1862 (O_1862,N_21700,N_22885);
or UO_1863 (O_1863,N_22378,N_22229);
or UO_1864 (O_1864,N_23518,N_20076);
and UO_1865 (O_1865,N_24082,N_20379);
and UO_1866 (O_1866,N_20470,N_21916);
xor UO_1867 (O_1867,N_22242,N_22472);
nand UO_1868 (O_1868,N_24860,N_20891);
and UO_1869 (O_1869,N_24380,N_21458);
and UO_1870 (O_1870,N_22469,N_22560);
or UO_1871 (O_1871,N_20949,N_21753);
nand UO_1872 (O_1872,N_24873,N_21397);
and UO_1873 (O_1873,N_24771,N_23550);
xnor UO_1874 (O_1874,N_22879,N_20203);
nor UO_1875 (O_1875,N_21953,N_24650);
and UO_1876 (O_1876,N_24588,N_21496);
and UO_1877 (O_1877,N_23981,N_23085);
or UO_1878 (O_1878,N_20478,N_24565);
nor UO_1879 (O_1879,N_20535,N_23316);
nor UO_1880 (O_1880,N_23963,N_20764);
nand UO_1881 (O_1881,N_24890,N_22317);
or UO_1882 (O_1882,N_22239,N_24828);
xor UO_1883 (O_1883,N_21850,N_23878);
nor UO_1884 (O_1884,N_20372,N_21189);
nand UO_1885 (O_1885,N_24781,N_24391);
nand UO_1886 (O_1886,N_24221,N_24865);
and UO_1887 (O_1887,N_22376,N_21775);
and UO_1888 (O_1888,N_23684,N_20155);
or UO_1889 (O_1889,N_22565,N_20745);
or UO_1890 (O_1890,N_20812,N_21938);
or UO_1891 (O_1891,N_23986,N_23195);
and UO_1892 (O_1892,N_23815,N_24243);
and UO_1893 (O_1893,N_20775,N_23539);
xor UO_1894 (O_1894,N_21678,N_20499);
nand UO_1895 (O_1895,N_23018,N_21384);
nor UO_1896 (O_1896,N_23818,N_21831);
or UO_1897 (O_1897,N_22175,N_22554);
xnor UO_1898 (O_1898,N_20044,N_23402);
or UO_1899 (O_1899,N_24369,N_20933);
nand UO_1900 (O_1900,N_21782,N_23111);
and UO_1901 (O_1901,N_20968,N_24556);
nor UO_1902 (O_1902,N_20401,N_22318);
nor UO_1903 (O_1903,N_21038,N_20640);
xnor UO_1904 (O_1904,N_22330,N_21324);
xnor UO_1905 (O_1905,N_23743,N_22856);
nor UO_1906 (O_1906,N_21232,N_20200);
xor UO_1907 (O_1907,N_23637,N_22102);
or UO_1908 (O_1908,N_20214,N_23078);
or UO_1909 (O_1909,N_22525,N_20779);
xor UO_1910 (O_1910,N_22055,N_23211);
nand UO_1911 (O_1911,N_24797,N_22326);
or UO_1912 (O_1912,N_23880,N_23657);
xor UO_1913 (O_1913,N_20335,N_24418);
nor UO_1914 (O_1914,N_21039,N_20479);
xor UO_1915 (O_1915,N_21350,N_22576);
nor UO_1916 (O_1916,N_21221,N_23616);
nor UO_1917 (O_1917,N_23142,N_23149);
or UO_1918 (O_1918,N_22044,N_20704);
or UO_1919 (O_1919,N_21578,N_20041);
and UO_1920 (O_1920,N_23573,N_24297);
nor UO_1921 (O_1921,N_20573,N_24210);
xnor UO_1922 (O_1922,N_24719,N_23879);
xor UO_1923 (O_1923,N_21784,N_23582);
xnor UO_1924 (O_1924,N_23945,N_21335);
and UO_1925 (O_1925,N_23740,N_22804);
nor UO_1926 (O_1926,N_23361,N_23507);
and UO_1927 (O_1927,N_22110,N_21288);
and UO_1928 (O_1928,N_20204,N_22308);
nand UO_1929 (O_1929,N_23735,N_20629);
nor UO_1930 (O_1930,N_23732,N_20872);
nand UO_1931 (O_1931,N_24878,N_21657);
and UO_1932 (O_1932,N_21155,N_22932);
nand UO_1933 (O_1933,N_23281,N_20598);
nor UO_1934 (O_1934,N_20015,N_23014);
xor UO_1935 (O_1935,N_21564,N_21689);
nand UO_1936 (O_1936,N_24876,N_21651);
or UO_1937 (O_1937,N_20147,N_21471);
or UO_1938 (O_1938,N_21390,N_20217);
nor UO_1939 (O_1939,N_20274,N_22807);
xnor UO_1940 (O_1940,N_24200,N_21144);
nor UO_1941 (O_1941,N_22194,N_24511);
or UO_1942 (O_1942,N_24026,N_24041);
and UO_1943 (O_1943,N_22465,N_20742);
or UO_1944 (O_1944,N_22563,N_20251);
and UO_1945 (O_1945,N_23553,N_23134);
and UO_1946 (O_1946,N_23371,N_20917);
and UO_1947 (O_1947,N_24279,N_23763);
nand UO_1948 (O_1948,N_21245,N_20095);
and UO_1949 (O_1949,N_22521,N_20778);
and UO_1950 (O_1950,N_20553,N_24524);
or UO_1951 (O_1951,N_24848,N_24815);
nand UO_1952 (O_1952,N_22414,N_21368);
nand UO_1953 (O_1953,N_24258,N_23331);
or UO_1954 (O_1954,N_20705,N_21259);
nand UO_1955 (O_1955,N_24569,N_21238);
xor UO_1956 (O_1956,N_24054,N_22266);
xor UO_1957 (O_1957,N_20436,N_23597);
nand UO_1958 (O_1958,N_22773,N_22492);
xnor UO_1959 (O_1959,N_21178,N_23010);
nand UO_1960 (O_1960,N_21252,N_21853);
or UO_1961 (O_1961,N_21532,N_22374);
or UO_1962 (O_1962,N_20449,N_21290);
nor UO_1963 (O_1963,N_21712,N_20601);
and UO_1964 (O_1964,N_24212,N_22771);
nor UO_1965 (O_1965,N_23500,N_23077);
xnor UO_1966 (O_1966,N_20163,N_20213);
or UO_1967 (O_1967,N_20043,N_21737);
or UO_1968 (O_1968,N_24231,N_20688);
or UO_1969 (O_1969,N_24843,N_23820);
nand UO_1970 (O_1970,N_21405,N_21618);
nor UO_1971 (O_1971,N_20545,N_24349);
or UO_1972 (O_1972,N_22523,N_22038);
xnor UO_1973 (O_1973,N_24144,N_23249);
nor UO_1974 (O_1974,N_23459,N_22301);
nand UO_1975 (O_1975,N_21832,N_23065);
nor UO_1976 (O_1976,N_23810,N_24864);
and UO_1977 (O_1977,N_21226,N_24023);
nor UO_1978 (O_1978,N_24775,N_22221);
xnor UO_1979 (O_1979,N_20673,N_23075);
or UO_1980 (O_1980,N_23128,N_24224);
xor UO_1981 (O_1981,N_21437,N_23598);
nor UO_1982 (O_1982,N_21962,N_23515);
or UO_1983 (O_1983,N_20146,N_21579);
nor UO_1984 (O_1984,N_23648,N_24192);
nand UO_1985 (O_1985,N_20042,N_23333);
nor UO_1986 (O_1986,N_21469,N_24371);
or UO_1987 (O_1987,N_20653,N_22369);
xor UO_1988 (O_1988,N_21860,N_24133);
nand UO_1989 (O_1989,N_23453,N_22534);
nor UO_1990 (O_1990,N_20148,N_22001);
nand UO_1991 (O_1991,N_21793,N_24425);
and UO_1992 (O_1992,N_20642,N_20013);
and UO_1993 (O_1993,N_24503,N_22697);
xor UO_1994 (O_1994,N_24920,N_23565);
or UO_1995 (O_1995,N_20760,N_20613);
xor UO_1996 (O_1996,N_22356,N_22155);
and UO_1997 (O_1997,N_22137,N_20118);
nor UO_1998 (O_1998,N_20561,N_22435);
or UO_1999 (O_1999,N_22411,N_24193);
and UO_2000 (O_2000,N_20442,N_24019);
nand UO_2001 (O_2001,N_22493,N_20070);
nor UO_2002 (O_2002,N_24989,N_22449);
xor UO_2003 (O_2003,N_21747,N_22713);
or UO_2004 (O_2004,N_22209,N_22793);
nor UO_2005 (O_2005,N_21646,N_24396);
nand UO_2006 (O_2006,N_20630,N_23592);
xnor UO_2007 (O_2007,N_24022,N_20792);
nand UO_2008 (O_2008,N_21044,N_22101);
and UO_2009 (O_2009,N_20905,N_21065);
xnor UO_2010 (O_2010,N_20025,N_23193);
or UO_2011 (O_2011,N_24544,N_23998);
xnor UO_2012 (O_2012,N_20946,N_23516);
nand UO_2013 (O_2013,N_23935,N_21709);
nand UO_2014 (O_2014,N_21424,N_21659);
or UO_2015 (O_2015,N_22919,N_21682);
or UO_2016 (O_2016,N_22518,N_22343);
nor UO_2017 (O_2017,N_20055,N_20064);
nor UO_2018 (O_2018,N_21067,N_22668);
nand UO_2019 (O_2019,N_22720,N_21654);
and UO_2020 (O_2020,N_21274,N_24407);
xor UO_2021 (O_2021,N_24472,N_24445);
nand UO_2022 (O_2022,N_21710,N_20755);
nand UO_2023 (O_2023,N_20534,N_21800);
or UO_2024 (O_2024,N_20711,N_23728);
nand UO_2025 (O_2025,N_24259,N_21838);
or UO_2026 (O_2026,N_20698,N_20938);
and UO_2027 (O_2027,N_23080,N_24906);
xor UO_2028 (O_2028,N_23938,N_21372);
and UO_2029 (O_2029,N_22998,N_20114);
xnor UO_2030 (O_2030,N_22073,N_24449);
nand UO_2031 (O_2031,N_23248,N_21842);
nand UO_2032 (O_2032,N_21410,N_24386);
nand UO_2033 (O_2033,N_23098,N_20353);
nor UO_2034 (O_2034,N_21357,N_24204);
nor UO_2035 (O_2035,N_23750,N_21978);
and UO_2036 (O_2036,N_22433,N_22079);
nand UO_2037 (O_2037,N_21031,N_20804);
xor UO_2038 (O_2038,N_22707,N_24911);
or UO_2039 (O_2039,N_23439,N_21836);
xnor UO_2040 (O_2040,N_21514,N_20215);
xnor UO_2041 (O_2041,N_22007,N_22992);
and UO_2042 (O_2042,N_24568,N_21764);
nor UO_2043 (O_2043,N_20324,N_23493);
nand UO_2044 (O_2044,N_22160,N_20304);
or UO_2045 (O_2045,N_24287,N_23892);
nor UO_2046 (O_2046,N_23540,N_24218);
or UO_2047 (O_2047,N_21928,N_21894);
and UO_2048 (O_2048,N_22434,N_24406);
and UO_2049 (O_2049,N_21946,N_23817);
and UO_2050 (O_2050,N_22654,N_21955);
xor UO_2051 (O_2051,N_22981,N_21246);
and UO_2052 (O_2052,N_24901,N_24755);
xnor UO_2053 (O_2053,N_22474,N_22186);
or UO_2054 (O_2054,N_21655,N_22711);
nor UO_2055 (O_2055,N_21756,N_22382);
nand UO_2056 (O_2056,N_24908,N_20709);
or UO_2057 (O_2057,N_20880,N_23692);
or UO_2058 (O_2058,N_20303,N_23108);
or UO_2059 (O_2059,N_21557,N_24008);
xnor UO_2060 (O_2060,N_22921,N_20953);
nor UO_2061 (O_2061,N_24522,N_20233);
nand UO_2062 (O_2062,N_21254,N_21984);
nand UO_2063 (O_2063,N_20165,N_21948);
xor UO_2064 (O_2064,N_20343,N_22637);
xnor UO_2065 (O_2065,N_21138,N_22146);
or UO_2066 (O_2066,N_23617,N_21900);
nor UO_2067 (O_2067,N_21699,N_22234);
nor UO_2068 (O_2068,N_21012,N_23228);
xor UO_2069 (O_2069,N_20182,N_20443);
xnor UO_2070 (O_2070,N_21975,N_22156);
or UO_2071 (O_2071,N_23673,N_20683);
nand UO_2072 (O_2072,N_23250,N_22020);
nand UO_2073 (O_2073,N_22495,N_20236);
or UO_2074 (O_2074,N_23259,N_23442);
nor UO_2075 (O_2075,N_20851,N_23605);
and UO_2076 (O_2076,N_23067,N_22621);
or UO_2077 (O_2077,N_22857,N_22940);
xor UO_2078 (O_2078,N_21283,N_23612);
nor UO_2079 (O_2079,N_20655,N_20875);
or UO_2080 (O_2080,N_23479,N_20636);
or UO_2081 (O_2081,N_24968,N_20985);
or UO_2082 (O_2082,N_24883,N_21208);
nor UO_2083 (O_2083,N_20336,N_20838);
nor UO_2084 (O_2084,N_21171,N_23386);
nor UO_2085 (O_2085,N_21326,N_21406);
xnor UO_2086 (O_2086,N_24991,N_20179);
or UO_2087 (O_2087,N_21803,N_23602);
and UO_2088 (O_2088,N_20354,N_23026);
nand UO_2089 (O_2089,N_22097,N_24877);
xnor UO_2090 (O_2090,N_23213,N_23679);
and UO_2091 (O_2091,N_20502,N_21207);
xor UO_2092 (O_2092,N_22132,N_22033);
nor UO_2093 (O_2093,N_21967,N_20973);
or UO_2094 (O_2094,N_23236,N_24431);
and UO_2095 (O_2095,N_21050,N_20834);
nor UO_2096 (O_2096,N_23191,N_24899);
nor UO_2097 (O_2097,N_24886,N_22018);
nand UO_2098 (O_2098,N_23359,N_20995);
nor UO_2099 (O_2099,N_23126,N_24061);
nor UO_2100 (O_2100,N_24826,N_24648);
xor UO_2101 (O_2101,N_20344,N_23700);
xnor UO_2102 (O_2102,N_24602,N_22139);
and UO_2103 (O_2103,N_21615,N_24319);
and UO_2104 (O_2104,N_23370,N_21533);
xnor UO_2105 (O_2105,N_22953,N_23863);
or UO_2106 (O_2106,N_20614,N_21299);
nand UO_2107 (O_2107,N_21158,N_21146);
or UO_2108 (O_2108,N_22134,N_22420);
xnor UO_2109 (O_2109,N_24168,N_22154);
and UO_2110 (O_2110,N_20398,N_23989);
nand UO_2111 (O_2111,N_22810,N_22053);
nand UO_2112 (O_2112,N_23258,N_21610);
or UO_2113 (O_2113,N_21000,N_20299);
and UO_2114 (O_2114,N_22624,N_24416);
nand UO_2115 (O_2115,N_20954,N_24939);
nor UO_2116 (O_2116,N_23816,N_21993);
xor UO_2117 (O_2117,N_21952,N_20769);
nor UO_2118 (O_2118,N_23167,N_24770);
and UO_2119 (O_2119,N_22737,N_20232);
or UO_2120 (O_2120,N_23293,N_20474);
or UO_2121 (O_2121,N_24205,N_23578);
nor UO_2122 (O_2122,N_23064,N_21218);
nand UO_2123 (O_2123,N_22681,N_21649);
nand UO_2124 (O_2124,N_24713,N_20896);
or UO_2125 (O_2125,N_21062,N_21224);
and UO_2126 (O_2126,N_22783,N_23063);
xor UO_2127 (O_2127,N_24805,N_23745);
or UO_2128 (O_2128,N_21983,N_21826);
and UO_2129 (O_2129,N_23418,N_21070);
or UO_2130 (O_2130,N_24283,N_24706);
nor UO_2131 (O_2131,N_24202,N_20318);
nor UO_2132 (O_2132,N_24412,N_23839);
nor UO_2133 (O_2133,N_22498,N_23037);
xor UO_2134 (O_2134,N_24165,N_23756);
nor UO_2135 (O_2135,N_22503,N_24092);
or UO_2136 (O_2136,N_24471,N_23523);
xnor UO_2137 (O_2137,N_20787,N_20181);
xnor UO_2138 (O_2138,N_22908,N_23388);
xor UO_2139 (O_2139,N_24236,N_22203);
and UO_2140 (O_2140,N_23734,N_20888);
nor UO_2141 (O_2141,N_21143,N_21414);
xor UO_2142 (O_2142,N_21257,N_22307);
nand UO_2143 (O_2143,N_20183,N_22990);
and UO_2144 (O_2144,N_22353,N_20866);
or UO_2145 (O_2145,N_24112,N_24882);
or UO_2146 (O_2146,N_20687,N_23825);
xor UO_2147 (O_2147,N_23680,N_21914);
xor UO_2148 (O_2148,N_20128,N_24662);
nor UO_2149 (O_2149,N_22995,N_23406);
xnor UO_2150 (O_2150,N_23969,N_23327);
xnor UO_2151 (O_2151,N_24548,N_23090);
xor UO_2152 (O_2152,N_21814,N_24261);
xor UO_2153 (O_2153,N_24002,N_20857);
nand UO_2154 (O_2154,N_20024,N_23224);
xor UO_2155 (O_2155,N_24011,N_20785);
xnor UO_2156 (O_2156,N_23883,N_21016);
or UO_2157 (O_2157,N_22674,N_24575);
or UO_2158 (O_2158,N_24330,N_24140);
nor UO_2159 (O_2159,N_24749,N_20558);
nand UO_2160 (O_2160,N_21219,N_21100);
nand UO_2161 (O_2161,N_21797,N_23755);
or UO_2162 (O_2162,N_23620,N_22117);
nand UO_2163 (O_2163,N_22257,N_22640);
nand UO_2164 (O_2164,N_22486,N_22405);
and UO_2165 (O_2165,N_22605,N_24701);
nor UO_2166 (O_2166,N_23158,N_23438);
or UO_2167 (O_2167,N_23624,N_24905);
xor UO_2168 (O_2168,N_20712,N_24904);
xor UO_2169 (O_2169,N_24115,N_20605);
nor UO_2170 (O_2170,N_24249,N_20503);
and UO_2171 (O_2171,N_23107,N_23622);
nor UO_2172 (O_2172,N_20770,N_23943);
or UO_2173 (O_2173,N_20130,N_23092);
xor UO_2174 (O_2174,N_23320,N_20656);
nand UO_2175 (O_2175,N_20669,N_21499);
nor UO_2176 (O_2176,N_21236,N_24543);
nand UO_2177 (O_2177,N_21844,N_24121);
xnor UO_2178 (O_2178,N_23436,N_21905);
nand UO_2179 (O_2179,N_23326,N_22912);
nor UO_2180 (O_2180,N_23336,N_20366);
or UO_2181 (O_2181,N_20850,N_21220);
nand UO_2182 (O_2182,N_24318,N_23409);
nor UO_2183 (O_2183,N_21994,N_22789);
xor UO_2184 (O_2184,N_24321,N_22060);
and UO_2185 (O_2185,N_24666,N_21604);
xnor UO_2186 (O_2186,N_22522,N_24378);
nor UO_2187 (O_2187,N_23401,N_24035);
nor UO_2188 (O_2188,N_23737,N_20625);
and UO_2189 (O_2189,N_24345,N_21282);
nand UO_2190 (O_2190,N_24304,N_21376);
and UO_2191 (O_2191,N_24718,N_23764);
nor UO_2192 (O_2192,N_21472,N_22426);
or UO_2193 (O_2193,N_23610,N_24622);
nor UO_2194 (O_2194,N_23774,N_22412);
nor UO_2195 (O_2195,N_22766,N_23587);
and UO_2196 (O_2196,N_23435,N_24608);
and UO_2197 (O_2197,N_24207,N_23696);
or UO_2198 (O_2198,N_20188,N_22632);
xnor UO_2199 (O_2199,N_24347,N_22049);
nor UO_2200 (O_2200,N_21561,N_20841);
nand UO_2201 (O_2201,N_20883,N_22657);
xor UO_2202 (O_2202,N_24563,N_24510);
xor UO_2203 (O_2203,N_22013,N_22005);
xnor UO_2204 (O_2204,N_20082,N_20193);
nor UO_2205 (O_2205,N_22944,N_22788);
nor UO_2206 (O_2206,N_21943,N_22888);
and UO_2207 (O_2207,N_22572,N_21940);
nor UO_2208 (O_2208,N_22977,N_20952);
or UO_2209 (O_2209,N_22616,N_21617);
nand UO_2210 (O_2210,N_20677,N_21440);
or UO_2211 (O_2211,N_23298,N_20643);
nand UO_2212 (O_2212,N_23872,N_21849);
xnor UO_2213 (O_2213,N_20540,N_23139);
or UO_2214 (O_2214,N_23514,N_22240);
xor UO_2215 (O_2215,N_20522,N_22967);
xnor UO_2216 (O_2216,N_23677,N_22679);
xnor UO_2217 (O_2217,N_24262,N_23970);
xnor UO_2218 (O_2218,N_24126,N_22901);
nand UO_2219 (O_2219,N_20671,N_20090);
and UO_2220 (O_2220,N_20137,N_22213);
xnor UO_2221 (O_2221,N_21396,N_24891);
xor UO_2222 (O_2222,N_21585,N_21653);
nor UO_2223 (O_2223,N_23979,N_23589);
xnor UO_2224 (O_2224,N_23643,N_20414);
nand UO_2225 (O_2225,N_23152,N_20045);
nand UO_2226 (O_2226,N_21986,N_22459);
nor UO_2227 (O_2227,N_23797,N_21748);
and UO_2228 (O_2228,N_21292,N_24938);
or UO_2229 (O_2229,N_24559,N_21497);
nor UO_2230 (O_2230,N_21910,N_21755);
nor UO_2231 (O_2231,N_20590,N_21971);
or UO_2232 (O_2232,N_23292,N_24107);
nor UO_2233 (O_2233,N_22362,N_24187);
xnor UO_2234 (O_2234,N_22345,N_21336);
xor UO_2235 (O_2235,N_22337,N_22170);
xor UO_2236 (O_2236,N_20666,N_20451);
nand UO_2237 (O_2237,N_22348,N_23006);
and UO_2238 (O_2238,N_24080,N_20541);
or UO_2239 (O_2239,N_21102,N_22447);
nor UO_2240 (O_2240,N_22153,N_24196);
and UO_2241 (O_2241,N_23909,N_24135);
nor UO_2242 (O_2242,N_20125,N_24068);
xor UO_2243 (O_2243,N_24376,N_20920);
and UO_2244 (O_2244,N_22874,N_22392);
xor UO_2245 (O_2245,N_24282,N_21964);
xor UO_2246 (O_2246,N_20692,N_23559);
nand UO_2247 (O_2247,N_23206,N_21926);
xnor UO_2248 (O_2248,N_20528,N_21280);
nand UO_2249 (O_2249,N_23185,N_24854);
nand UO_2250 (O_2250,N_20579,N_22853);
nor UO_2251 (O_2251,N_20191,N_22588);
and UO_2252 (O_2252,N_22178,N_23812);
and UO_2253 (O_2253,N_24136,N_23521);
nor UO_2254 (O_2254,N_21898,N_21385);
and UO_2255 (O_2255,N_24972,N_21052);
nand UO_2256 (O_2256,N_24599,N_22779);
or UO_2257 (O_2257,N_24220,N_22685);
and UO_2258 (O_2258,N_23920,N_23062);
nand UO_2259 (O_2259,N_23894,N_22274);
xnor UO_2260 (O_2260,N_22131,N_21903);
xor UO_2261 (O_2261,N_24983,N_22205);
xnor UO_2262 (O_2262,N_20751,N_20794);
nand UO_2263 (O_2263,N_21182,N_20293);
nor UO_2264 (O_2264,N_22610,N_24191);
xor UO_2265 (O_2265,N_20186,N_21430);
or UO_2266 (O_2266,N_20207,N_24927);
nor UO_2267 (O_2267,N_23672,N_21455);
nor UO_2268 (O_2268,N_22558,N_21587);
xnor UO_2269 (O_2269,N_20739,N_23542);
and UO_2270 (O_2270,N_20925,N_20016);
or UO_2271 (O_2271,N_23101,N_23366);
or UO_2272 (O_2272,N_22639,N_22916);
and UO_2273 (O_2273,N_22277,N_21492);
nand UO_2274 (O_2274,N_23525,N_22017);
nor UO_2275 (O_2275,N_20639,N_20554);
nand UO_2276 (O_2276,N_23458,N_24984);
nand UO_2277 (O_2277,N_20665,N_22191);
nand UO_2278 (O_2278,N_20928,N_22593);
nor UO_2279 (O_2279,N_20161,N_22453);
xnor UO_2280 (O_2280,N_20526,N_22280);
nor UO_2281 (O_2281,N_24146,N_20908);
or UO_2282 (O_2282,N_24996,N_23290);
and UO_2283 (O_2283,N_23621,N_22148);
nand UO_2284 (O_2284,N_24415,N_24131);
or UO_2285 (O_2285,N_24678,N_24278);
and UO_2286 (O_2286,N_24048,N_24766);
nand UO_2287 (O_2287,N_20158,N_23710);
nor UO_2288 (O_2288,N_23502,N_22042);
nand UO_2289 (O_2289,N_23390,N_20932);
xnor UO_2290 (O_2290,N_23275,N_21312);
xor UO_2291 (O_2291,N_23584,N_20486);
and UO_2292 (O_2292,N_20341,N_24162);
or UO_2293 (O_2293,N_20247,N_22839);
and UO_2294 (O_2294,N_21852,N_20423);
nand UO_2295 (O_2295,N_20809,N_22687);
and UO_2296 (O_2296,N_20093,N_20201);
nand UO_2297 (O_2297,N_24308,N_24897);
nor UO_2298 (O_2298,N_22000,N_22058);
nand UO_2299 (O_2299,N_24959,N_24307);
nor UO_2300 (O_2300,N_21608,N_24027);
or UO_2301 (O_2301,N_22201,N_23414);
nand UO_2302 (O_2302,N_21491,N_24043);
or UO_2303 (O_2303,N_21547,N_23277);
xor UO_2304 (O_2304,N_22535,N_21133);
and UO_2305 (O_2305,N_24057,N_21115);
nand UO_2306 (O_2306,N_21722,N_22063);
nor UO_2307 (O_2307,N_20046,N_20685);
or UO_2308 (O_2308,N_23495,N_21249);
xor UO_2309 (O_2309,N_20378,N_20471);
nor UO_2310 (O_2310,N_21095,N_22306);
or UO_2311 (O_2311,N_23071,N_22295);
nor UO_2312 (O_2312,N_20009,N_21690);
nor UO_2313 (O_2313,N_23526,N_21165);
xnor UO_2314 (O_2314,N_22484,N_24714);
nand UO_2315 (O_2315,N_24571,N_20243);
xnor UO_2316 (O_2316,N_20619,N_21999);
nand UO_2317 (O_2317,N_22404,N_22227);
nor UO_2318 (O_2318,N_21974,N_23724);
nor UO_2319 (O_2319,N_24616,N_23538);
xor UO_2320 (O_2320,N_22340,N_24970);
nand UO_2321 (O_2321,N_23363,N_23772);
xnor UO_2322 (O_2322,N_20084,N_22311);
nor UO_2323 (O_2323,N_20409,N_21198);
xnor UO_2324 (O_2324,N_21352,N_22591);
nor UO_2325 (O_2325,N_22948,N_21941);
or UO_2326 (O_2326,N_22951,N_20383);
xor UO_2327 (O_2327,N_22473,N_21667);
xor UO_2328 (O_2328,N_22700,N_22112);
nor UO_2329 (O_2329,N_23949,N_21518);
nor UO_2330 (O_2330,N_20853,N_22933);
nor UO_2331 (O_2331,N_23141,N_22652);
nor UO_2332 (O_2332,N_22816,N_20057);
nand UO_2333 (O_2333,N_22997,N_20707);
nand UO_2334 (O_2334,N_23675,N_20387);
or UO_2335 (O_2335,N_22775,N_24413);
or UO_2336 (O_2336,N_22930,N_22176);
and UO_2337 (O_2337,N_20153,N_20159);
xnor UO_2338 (O_2338,N_20587,N_24949);
or UO_2339 (O_2339,N_24388,N_21104);
nand UO_2340 (O_2340,N_23485,N_24683);
xnor UO_2341 (O_2341,N_23996,N_21669);
nand UO_2342 (O_2342,N_22419,N_24688);
or UO_2343 (O_2343,N_22200,N_21174);
nor UO_2344 (O_2344,N_23031,N_24296);
nor UO_2345 (O_2345,N_21068,N_23886);
xor UO_2346 (O_2346,N_20943,N_24735);
nand UO_2347 (O_2347,N_23765,N_20367);
or UO_2348 (O_2348,N_21298,N_22865);
or UO_2349 (O_2349,N_22048,N_24740);
and UO_2350 (O_2350,N_20416,N_21503);
nor UO_2351 (O_2351,N_21395,N_20800);
xnor UO_2352 (O_2352,N_20061,N_21339);
nor UO_2353 (O_2353,N_22290,N_23958);
nand UO_2354 (O_2354,N_24256,N_21641);
and UO_2355 (O_2355,N_23738,N_24792);
or UO_2356 (O_2356,N_20290,N_21785);
nand UO_2357 (O_2357,N_23201,N_23633);
xor UO_2358 (O_2358,N_23024,N_23199);
and UO_2359 (O_2359,N_23104,N_21524);
or UO_2360 (O_2360,N_24227,N_21592);
nor UO_2361 (O_2361,N_20053,N_22618);
xnor UO_2362 (O_2362,N_20149,N_23792);
or UO_2363 (O_2363,N_20081,N_22578);
nand UO_2364 (O_2364,N_23147,N_22034);
nor UO_2365 (O_2365,N_21977,N_24513);
nand UO_2366 (O_2366,N_22479,N_21521);
nor UO_2367 (O_2367,N_22511,N_22208);
xor UO_2368 (O_2368,N_21790,N_22515);
xnor UO_2369 (O_2369,N_24912,N_21936);
nor UO_2370 (O_2370,N_21509,N_24975);
nand UO_2371 (O_2371,N_20178,N_24067);
nor UO_2372 (O_2372,N_24768,N_24125);
nor UO_2373 (O_2373,N_21602,N_24909);
nor UO_2374 (O_2374,N_22818,N_22524);
nand UO_2375 (O_2375,N_22520,N_20431);
and UO_2376 (O_2376,N_20417,N_22384);
or UO_2377 (O_2377,N_24363,N_20099);
or UO_2378 (O_2378,N_23395,N_20194);
nor UO_2379 (O_2379,N_20310,N_21202);
nor UO_2380 (O_2380,N_23749,N_24592);
xnor UO_2381 (O_2381,N_24633,N_24099);
or UO_2382 (O_2382,N_22256,N_20959);
nor UO_2383 (O_2383,N_20806,N_24497);
or UO_2384 (O_2384,N_21821,N_21841);
and UO_2385 (O_2385,N_20520,N_24423);
and UO_2386 (O_2386,N_23552,N_22304);
and UO_2387 (O_2387,N_23625,N_21542);
nor UO_2388 (O_2388,N_22342,N_21558);
nor UO_2389 (O_2389,N_20504,N_20909);
nand UO_2390 (O_2390,N_22765,N_24567);
nor UO_2391 (O_2391,N_20393,N_22164);
or UO_2392 (O_2392,N_24785,N_23115);
xor UO_2393 (O_2393,N_22421,N_22741);
nand UO_2394 (O_2394,N_23027,N_23504);
and UO_2395 (O_2395,N_24176,N_21876);
xor UO_2396 (O_2396,N_21055,N_20026);
and UO_2397 (O_2397,N_24742,N_23428);
and UO_2398 (O_2398,N_23056,N_23381);
nor UO_2399 (O_2399,N_21675,N_22011);
and UO_2400 (O_2400,N_23668,N_20903);
nor UO_2401 (O_2401,N_22546,N_22911);
nor UO_2402 (O_2402,N_24480,N_22760);
nand UO_2403 (O_2403,N_22871,N_22288);
xnor UO_2404 (O_2404,N_21485,N_24464);
xor UO_2405 (O_2405,N_24872,N_23319);
and UO_2406 (O_2406,N_21131,N_22275);
and UO_2407 (O_2407,N_24798,N_22802);
xnor UO_2408 (O_2408,N_22648,N_20982);
nand UO_2409 (O_2409,N_20454,N_20307);
or UO_2410 (O_2410,N_20747,N_23930);
and UO_2411 (O_2411,N_24850,N_24887);
nor UO_2412 (O_2412,N_24580,N_21097);
xnor UO_2413 (O_2413,N_23253,N_21474);
or UO_2414 (O_2414,N_20645,N_23138);
and UO_2415 (O_2415,N_21628,N_23287);
nand UO_2416 (O_2416,N_21205,N_24525);
nand UO_2417 (O_2417,N_22289,N_21461);
nand UO_2418 (O_2418,N_24402,N_22466);
and UO_2419 (O_2419,N_21665,N_20284);
nand UO_2420 (O_2420,N_24612,N_24834);
xor UO_2421 (O_2421,N_23960,N_24381);
nand UO_2422 (O_2422,N_24637,N_20549);
xor UO_2423 (O_2423,N_23634,N_24096);
xor UO_2424 (O_2424,N_24263,N_22262);
nor UO_2425 (O_2425,N_23205,N_24918);
xnor UO_2426 (O_2426,N_22851,N_21480);
or UO_2427 (O_2427,N_22212,N_20231);
nor UO_2428 (O_2428,N_21723,N_20962);
or UO_2429 (O_2429,N_24846,N_24948);
nor UO_2430 (O_2430,N_22589,N_21079);
nor UO_2431 (O_2431,N_23600,N_22695);
xor UO_2432 (O_2432,N_22438,N_21332);
nor UO_2433 (O_2433,N_20720,N_23218);
nand UO_2434 (O_2434,N_21530,N_23805);
nand UO_2435 (O_2435,N_24170,N_20010);
or UO_2436 (O_2436,N_23855,N_24142);
nand UO_2437 (O_2437,N_23862,N_20588);
and UO_2438 (O_2438,N_22028,N_24594);
xnor UO_2439 (O_2439,N_20539,N_21818);
and UO_2440 (O_2440,N_22210,N_24557);
xnor UO_2441 (O_2441,N_21151,N_23499);
xnor UO_2442 (O_2442,N_21212,N_21253);
nor UO_2443 (O_2443,N_23423,N_20763);
or UO_2444 (O_2444,N_23447,N_22168);
and UO_2445 (O_2445,N_20234,N_24044);
and UO_2446 (O_2446,N_23271,N_21854);
xnor UO_2447 (O_2447,N_23021,N_21233);
xnor UO_2448 (O_2448,N_21053,N_21367);
or UO_2449 (O_2449,N_20127,N_24907);
xor UO_2450 (O_2450,N_24604,N_23551);
nand UO_2451 (O_2451,N_22379,N_21287);
nand UO_2452 (O_2452,N_20654,N_21829);
or UO_2453 (O_2453,N_22863,N_23241);
nor UO_2454 (O_2454,N_23073,N_21241);
nor UO_2455 (O_2455,N_21696,N_22504);
and UO_2456 (O_2456,N_21652,N_24954);
and UO_2457 (O_2457,N_21123,N_21574);
xor UO_2458 (O_2458,N_21388,N_20268);
nor UO_2459 (O_2459,N_24644,N_20221);
and UO_2460 (O_2460,N_20079,N_21427);
or UO_2461 (O_2461,N_21074,N_21658);
nor UO_2462 (O_2462,N_20512,N_22847);
or UO_2463 (O_2463,N_22335,N_23530);
xor UO_2464 (O_2464,N_22959,N_22114);
and UO_2465 (O_2465,N_24083,N_23029);
nand UO_2466 (O_2466,N_23468,N_22890);
and UO_2467 (O_2467,N_24070,N_22686);
nor UO_2468 (O_2468,N_21107,N_24611);
and UO_2469 (O_2469,N_23865,N_24553);
nor UO_2470 (O_2470,N_20510,N_22552);
or UO_2471 (O_2471,N_20637,N_23304);
xor UO_2472 (O_2472,N_20444,N_24744);
and UO_2473 (O_2473,N_23641,N_24060);
nand UO_2474 (O_2474,N_20832,N_20728);
nand UO_2475 (O_2475,N_24659,N_20281);
nor UO_2476 (O_2476,N_24762,N_24059);
and UO_2477 (O_2477,N_21227,N_24466);
or UO_2478 (O_2478,N_24089,N_20022);
nand UO_2479 (O_2479,N_22692,N_24333);
and UO_2480 (O_2480,N_22489,N_24143);
xor UO_2481 (O_2481,N_22893,N_23811);
and UO_2482 (O_2482,N_21035,N_22251);
nor UO_2483 (O_2483,N_23296,N_23944);
and UO_2484 (O_2484,N_20532,N_24331);
nor UO_2485 (O_2485,N_24750,N_20660);
or UO_2486 (O_2486,N_20519,N_20350);
xnor UO_2487 (O_2487,N_20762,N_23845);
and UO_2488 (O_2488,N_23011,N_23976);
or UO_2489 (O_2489,N_22461,N_21567);
xor UO_2490 (O_2490,N_21515,N_24305);
xnor UO_2491 (O_2491,N_24437,N_20533);
xor UO_2492 (O_2492,N_21432,N_21134);
xnor UO_2493 (O_2493,N_23264,N_20339);
xor UO_2494 (O_2494,N_24695,N_22938);
xor UO_2495 (O_2495,N_23636,N_24299);
nand UO_2496 (O_2496,N_23000,N_20771);
xnor UO_2497 (O_2497,N_24139,N_22238);
nand UO_2498 (O_2498,N_23133,N_20703);
or UO_2499 (O_2499,N_22746,N_21181);
and UO_2500 (O_2500,N_23320,N_24235);
nor UO_2501 (O_2501,N_23486,N_20021);
nor UO_2502 (O_2502,N_20805,N_23736);
xor UO_2503 (O_2503,N_24971,N_20683);
nor UO_2504 (O_2504,N_21486,N_23768);
nor UO_2505 (O_2505,N_23714,N_23178);
and UO_2506 (O_2506,N_20872,N_24073);
or UO_2507 (O_2507,N_21665,N_22243);
xor UO_2508 (O_2508,N_23050,N_22392);
xnor UO_2509 (O_2509,N_22003,N_23589);
nand UO_2510 (O_2510,N_24727,N_23332);
nor UO_2511 (O_2511,N_22577,N_24311);
xor UO_2512 (O_2512,N_23461,N_20223);
nand UO_2513 (O_2513,N_22248,N_22949);
nor UO_2514 (O_2514,N_24639,N_24508);
xor UO_2515 (O_2515,N_23635,N_20609);
nand UO_2516 (O_2516,N_24181,N_20401);
xnor UO_2517 (O_2517,N_21486,N_24433);
nand UO_2518 (O_2518,N_24813,N_22928);
xnor UO_2519 (O_2519,N_23104,N_22993);
and UO_2520 (O_2520,N_24295,N_21943);
or UO_2521 (O_2521,N_22340,N_24545);
or UO_2522 (O_2522,N_22488,N_21105);
xnor UO_2523 (O_2523,N_23474,N_20207);
xor UO_2524 (O_2524,N_20632,N_22203);
and UO_2525 (O_2525,N_22401,N_21315);
nor UO_2526 (O_2526,N_24050,N_23814);
xnor UO_2527 (O_2527,N_22740,N_20753);
nor UO_2528 (O_2528,N_21719,N_20477);
nand UO_2529 (O_2529,N_24219,N_20949);
xor UO_2530 (O_2530,N_23850,N_22638);
or UO_2531 (O_2531,N_20154,N_21573);
nor UO_2532 (O_2532,N_23869,N_24060);
xor UO_2533 (O_2533,N_20503,N_24351);
and UO_2534 (O_2534,N_22316,N_24798);
or UO_2535 (O_2535,N_21312,N_21062);
xnor UO_2536 (O_2536,N_20262,N_21116);
xor UO_2537 (O_2537,N_21816,N_24283);
and UO_2538 (O_2538,N_23960,N_22755);
nand UO_2539 (O_2539,N_24966,N_22920);
and UO_2540 (O_2540,N_23498,N_21567);
and UO_2541 (O_2541,N_24836,N_23835);
nand UO_2542 (O_2542,N_20999,N_23120);
nand UO_2543 (O_2543,N_21315,N_23771);
nand UO_2544 (O_2544,N_22912,N_22951);
or UO_2545 (O_2545,N_21120,N_21917);
nor UO_2546 (O_2546,N_22768,N_24800);
and UO_2547 (O_2547,N_21854,N_22163);
and UO_2548 (O_2548,N_24910,N_20975);
nor UO_2549 (O_2549,N_22506,N_23852);
nand UO_2550 (O_2550,N_23440,N_20765);
or UO_2551 (O_2551,N_20277,N_21926);
xor UO_2552 (O_2552,N_21920,N_21350);
or UO_2553 (O_2553,N_21836,N_22889);
nor UO_2554 (O_2554,N_20170,N_23060);
nor UO_2555 (O_2555,N_20551,N_22382);
and UO_2556 (O_2556,N_20384,N_23815);
xnor UO_2557 (O_2557,N_21874,N_23136);
xor UO_2558 (O_2558,N_22871,N_20089);
xor UO_2559 (O_2559,N_22731,N_23117);
or UO_2560 (O_2560,N_21662,N_21916);
nor UO_2561 (O_2561,N_22084,N_24369);
nand UO_2562 (O_2562,N_23846,N_24427);
nand UO_2563 (O_2563,N_22015,N_24446);
xor UO_2564 (O_2564,N_24200,N_24406);
or UO_2565 (O_2565,N_24161,N_20198);
nor UO_2566 (O_2566,N_21365,N_24941);
nor UO_2567 (O_2567,N_22993,N_20679);
or UO_2568 (O_2568,N_22958,N_24524);
and UO_2569 (O_2569,N_22493,N_20204);
xnor UO_2570 (O_2570,N_24172,N_20910);
and UO_2571 (O_2571,N_23473,N_23110);
nand UO_2572 (O_2572,N_23476,N_20656);
nor UO_2573 (O_2573,N_22834,N_21723);
nor UO_2574 (O_2574,N_20746,N_20539);
xnor UO_2575 (O_2575,N_22680,N_22595);
nand UO_2576 (O_2576,N_23651,N_21147);
nand UO_2577 (O_2577,N_23193,N_20631);
and UO_2578 (O_2578,N_21554,N_23235);
nor UO_2579 (O_2579,N_21037,N_23310);
or UO_2580 (O_2580,N_24407,N_24649);
nand UO_2581 (O_2581,N_20373,N_21736);
or UO_2582 (O_2582,N_21232,N_23440);
xor UO_2583 (O_2583,N_22844,N_21806);
or UO_2584 (O_2584,N_24376,N_21058);
and UO_2585 (O_2585,N_20067,N_20603);
xor UO_2586 (O_2586,N_20759,N_23295);
or UO_2587 (O_2587,N_20194,N_21118);
nand UO_2588 (O_2588,N_22289,N_20584);
and UO_2589 (O_2589,N_23346,N_20213);
and UO_2590 (O_2590,N_22109,N_20769);
or UO_2591 (O_2591,N_20930,N_23423);
or UO_2592 (O_2592,N_21523,N_20887);
nand UO_2593 (O_2593,N_22409,N_24540);
nand UO_2594 (O_2594,N_20763,N_22083);
nor UO_2595 (O_2595,N_23980,N_20400);
nor UO_2596 (O_2596,N_20898,N_23126);
nor UO_2597 (O_2597,N_24391,N_22550);
nor UO_2598 (O_2598,N_22740,N_23331);
or UO_2599 (O_2599,N_23020,N_20286);
or UO_2600 (O_2600,N_23547,N_22876);
nand UO_2601 (O_2601,N_20141,N_24560);
or UO_2602 (O_2602,N_23917,N_22476);
or UO_2603 (O_2603,N_22629,N_22541);
nand UO_2604 (O_2604,N_20710,N_21273);
or UO_2605 (O_2605,N_23266,N_21799);
or UO_2606 (O_2606,N_24236,N_23645);
xor UO_2607 (O_2607,N_20845,N_23334);
nor UO_2608 (O_2608,N_23364,N_20363);
nand UO_2609 (O_2609,N_24656,N_22941);
and UO_2610 (O_2610,N_24191,N_22160);
nand UO_2611 (O_2611,N_21925,N_24846);
nand UO_2612 (O_2612,N_20582,N_22673);
nor UO_2613 (O_2613,N_20821,N_21100);
or UO_2614 (O_2614,N_20773,N_23870);
nor UO_2615 (O_2615,N_22101,N_24961);
xnor UO_2616 (O_2616,N_21668,N_23940);
xnor UO_2617 (O_2617,N_21274,N_22421);
or UO_2618 (O_2618,N_20384,N_22757);
or UO_2619 (O_2619,N_23046,N_21888);
xor UO_2620 (O_2620,N_22028,N_21188);
xnor UO_2621 (O_2621,N_23498,N_22013);
nor UO_2622 (O_2622,N_22640,N_20790);
nor UO_2623 (O_2623,N_24858,N_24087);
and UO_2624 (O_2624,N_22269,N_20719);
nand UO_2625 (O_2625,N_22637,N_22630);
nand UO_2626 (O_2626,N_21042,N_22291);
nor UO_2627 (O_2627,N_20354,N_20001);
nor UO_2628 (O_2628,N_20731,N_21294);
xor UO_2629 (O_2629,N_20351,N_22324);
xor UO_2630 (O_2630,N_21242,N_23060);
xor UO_2631 (O_2631,N_22011,N_21847);
nor UO_2632 (O_2632,N_22135,N_23773);
and UO_2633 (O_2633,N_20968,N_21940);
xnor UO_2634 (O_2634,N_24930,N_20992);
and UO_2635 (O_2635,N_20100,N_24037);
and UO_2636 (O_2636,N_21148,N_20883);
nand UO_2637 (O_2637,N_20056,N_20263);
xnor UO_2638 (O_2638,N_21835,N_21539);
or UO_2639 (O_2639,N_23963,N_23065);
nor UO_2640 (O_2640,N_24621,N_24206);
nor UO_2641 (O_2641,N_23736,N_21017);
or UO_2642 (O_2642,N_20825,N_21967);
or UO_2643 (O_2643,N_24284,N_21986);
and UO_2644 (O_2644,N_23599,N_20658);
xor UO_2645 (O_2645,N_21033,N_20247);
and UO_2646 (O_2646,N_23765,N_22639);
nand UO_2647 (O_2647,N_22870,N_24317);
xor UO_2648 (O_2648,N_22836,N_21692);
xnor UO_2649 (O_2649,N_20669,N_24019);
nor UO_2650 (O_2650,N_23926,N_22507);
or UO_2651 (O_2651,N_24458,N_20361);
nand UO_2652 (O_2652,N_22177,N_24296);
and UO_2653 (O_2653,N_24356,N_23160);
nand UO_2654 (O_2654,N_23892,N_22765);
nand UO_2655 (O_2655,N_24884,N_23959);
or UO_2656 (O_2656,N_20287,N_23591);
and UO_2657 (O_2657,N_20604,N_22988);
nor UO_2658 (O_2658,N_24451,N_24391);
xnor UO_2659 (O_2659,N_20316,N_20705);
or UO_2660 (O_2660,N_24485,N_20771);
nand UO_2661 (O_2661,N_21978,N_24962);
xor UO_2662 (O_2662,N_24301,N_24728);
xnor UO_2663 (O_2663,N_22663,N_22857);
xor UO_2664 (O_2664,N_21029,N_22371);
and UO_2665 (O_2665,N_22762,N_23727);
nor UO_2666 (O_2666,N_22987,N_23238);
nor UO_2667 (O_2667,N_21491,N_21284);
and UO_2668 (O_2668,N_22700,N_21198);
xnor UO_2669 (O_2669,N_20223,N_22962);
xor UO_2670 (O_2670,N_20584,N_20881);
and UO_2671 (O_2671,N_23411,N_21421);
nand UO_2672 (O_2672,N_23213,N_20805);
and UO_2673 (O_2673,N_24483,N_21379);
xnor UO_2674 (O_2674,N_24192,N_21526);
xor UO_2675 (O_2675,N_23490,N_21946);
nand UO_2676 (O_2676,N_23113,N_24959);
or UO_2677 (O_2677,N_20884,N_23853);
nor UO_2678 (O_2678,N_21144,N_23420);
nand UO_2679 (O_2679,N_23156,N_23712);
nor UO_2680 (O_2680,N_22426,N_22024);
nand UO_2681 (O_2681,N_24516,N_22436);
nor UO_2682 (O_2682,N_23891,N_24843);
nor UO_2683 (O_2683,N_24473,N_24290);
and UO_2684 (O_2684,N_20405,N_23987);
nand UO_2685 (O_2685,N_24605,N_21540);
nand UO_2686 (O_2686,N_20439,N_22328);
or UO_2687 (O_2687,N_21711,N_20464);
and UO_2688 (O_2688,N_20456,N_22238);
nor UO_2689 (O_2689,N_24185,N_23178);
and UO_2690 (O_2690,N_24584,N_21044);
nor UO_2691 (O_2691,N_21348,N_22876);
nor UO_2692 (O_2692,N_24478,N_22665);
or UO_2693 (O_2693,N_21370,N_24227);
and UO_2694 (O_2694,N_24158,N_21044);
nor UO_2695 (O_2695,N_23059,N_24685);
or UO_2696 (O_2696,N_24416,N_23219);
or UO_2697 (O_2697,N_24055,N_20807);
xor UO_2698 (O_2698,N_24792,N_24981);
nand UO_2699 (O_2699,N_20842,N_20382);
nor UO_2700 (O_2700,N_23619,N_24157);
nand UO_2701 (O_2701,N_20425,N_23759);
or UO_2702 (O_2702,N_20164,N_21593);
xor UO_2703 (O_2703,N_20875,N_21000);
and UO_2704 (O_2704,N_24575,N_21474);
and UO_2705 (O_2705,N_23189,N_21353);
nand UO_2706 (O_2706,N_21378,N_22830);
xor UO_2707 (O_2707,N_20402,N_23929);
or UO_2708 (O_2708,N_22453,N_20368);
nand UO_2709 (O_2709,N_23339,N_21386);
or UO_2710 (O_2710,N_22189,N_23654);
nand UO_2711 (O_2711,N_24020,N_20660);
and UO_2712 (O_2712,N_21804,N_21764);
nor UO_2713 (O_2713,N_22900,N_24952);
xor UO_2714 (O_2714,N_21862,N_20065);
xor UO_2715 (O_2715,N_20597,N_24229);
nor UO_2716 (O_2716,N_22815,N_22144);
nor UO_2717 (O_2717,N_22090,N_21322);
or UO_2718 (O_2718,N_20255,N_24471);
nand UO_2719 (O_2719,N_22018,N_21487);
or UO_2720 (O_2720,N_22995,N_22068);
or UO_2721 (O_2721,N_22463,N_21926);
nor UO_2722 (O_2722,N_24983,N_23655);
xnor UO_2723 (O_2723,N_20892,N_23308);
xor UO_2724 (O_2724,N_22458,N_21002);
and UO_2725 (O_2725,N_23458,N_22673);
or UO_2726 (O_2726,N_21440,N_22113);
or UO_2727 (O_2727,N_23085,N_23865);
xnor UO_2728 (O_2728,N_21394,N_23893);
or UO_2729 (O_2729,N_20806,N_24062);
or UO_2730 (O_2730,N_21365,N_23442);
nor UO_2731 (O_2731,N_20357,N_24464);
xnor UO_2732 (O_2732,N_24252,N_22510);
and UO_2733 (O_2733,N_20288,N_24979);
nand UO_2734 (O_2734,N_21175,N_24928);
or UO_2735 (O_2735,N_21192,N_20033);
and UO_2736 (O_2736,N_21506,N_21985);
or UO_2737 (O_2737,N_23151,N_24517);
xnor UO_2738 (O_2738,N_21153,N_23940);
xnor UO_2739 (O_2739,N_22755,N_23656);
nor UO_2740 (O_2740,N_23388,N_20265);
and UO_2741 (O_2741,N_20653,N_22883);
and UO_2742 (O_2742,N_24959,N_24769);
nor UO_2743 (O_2743,N_22949,N_21098);
xor UO_2744 (O_2744,N_22162,N_22449);
or UO_2745 (O_2745,N_24153,N_22535);
xnor UO_2746 (O_2746,N_23989,N_21507);
nor UO_2747 (O_2747,N_23163,N_21142);
nor UO_2748 (O_2748,N_20639,N_20851);
nor UO_2749 (O_2749,N_21376,N_24848);
nand UO_2750 (O_2750,N_20015,N_23283);
or UO_2751 (O_2751,N_21321,N_21221);
and UO_2752 (O_2752,N_21426,N_20507);
nor UO_2753 (O_2753,N_20534,N_24561);
nand UO_2754 (O_2754,N_23438,N_20242);
nor UO_2755 (O_2755,N_24825,N_23208);
or UO_2756 (O_2756,N_20359,N_21055);
or UO_2757 (O_2757,N_22360,N_21960);
nor UO_2758 (O_2758,N_23030,N_23386);
nand UO_2759 (O_2759,N_23696,N_20667);
nor UO_2760 (O_2760,N_21329,N_24754);
and UO_2761 (O_2761,N_24501,N_20717);
and UO_2762 (O_2762,N_20352,N_24642);
xor UO_2763 (O_2763,N_24474,N_23524);
nand UO_2764 (O_2764,N_23338,N_21256);
xnor UO_2765 (O_2765,N_20748,N_21326);
or UO_2766 (O_2766,N_21220,N_20936);
or UO_2767 (O_2767,N_23072,N_22695);
nand UO_2768 (O_2768,N_20115,N_24193);
xnor UO_2769 (O_2769,N_23767,N_20194);
nand UO_2770 (O_2770,N_22289,N_21779);
nand UO_2771 (O_2771,N_20850,N_23296);
xor UO_2772 (O_2772,N_24512,N_24847);
nand UO_2773 (O_2773,N_22906,N_20657);
nor UO_2774 (O_2774,N_20444,N_22274);
nand UO_2775 (O_2775,N_23993,N_22395);
nor UO_2776 (O_2776,N_22725,N_22754);
nor UO_2777 (O_2777,N_20006,N_20662);
nor UO_2778 (O_2778,N_21945,N_23497);
nor UO_2779 (O_2779,N_24035,N_24640);
nand UO_2780 (O_2780,N_21950,N_21415);
nor UO_2781 (O_2781,N_22312,N_21346);
and UO_2782 (O_2782,N_21054,N_20382);
or UO_2783 (O_2783,N_24300,N_21929);
xor UO_2784 (O_2784,N_20697,N_23919);
or UO_2785 (O_2785,N_21934,N_23588);
nor UO_2786 (O_2786,N_24107,N_24667);
nand UO_2787 (O_2787,N_21788,N_22772);
xor UO_2788 (O_2788,N_24934,N_21752);
xnor UO_2789 (O_2789,N_22134,N_20347);
or UO_2790 (O_2790,N_20558,N_24022);
nor UO_2791 (O_2791,N_22463,N_24777);
or UO_2792 (O_2792,N_23067,N_23083);
xnor UO_2793 (O_2793,N_20779,N_24160);
xnor UO_2794 (O_2794,N_24435,N_22975);
or UO_2795 (O_2795,N_20150,N_21426);
xor UO_2796 (O_2796,N_22883,N_21039);
nand UO_2797 (O_2797,N_23562,N_20988);
nand UO_2798 (O_2798,N_21501,N_20862);
nor UO_2799 (O_2799,N_21782,N_21090);
or UO_2800 (O_2800,N_22629,N_22527);
nand UO_2801 (O_2801,N_20024,N_21337);
xnor UO_2802 (O_2802,N_24633,N_23838);
and UO_2803 (O_2803,N_24613,N_23400);
nor UO_2804 (O_2804,N_20861,N_20592);
nand UO_2805 (O_2805,N_23173,N_23227);
xor UO_2806 (O_2806,N_21690,N_24218);
or UO_2807 (O_2807,N_23638,N_22408);
nor UO_2808 (O_2808,N_21033,N_22855);
or UO_2809 (O_2809,N_24316,N_20566);
nor UO_2810 (O_2810,N_21126,N_24189);
nand UO_2811 (O_2811,N_20639,N_21291);
and UO_2812 (O_2812,N_21320,N_22170);
and UO_2813 (O_2813,N_24682,N_22862);
or UO_2814 (O_2814,N_20423,N_24164);
nor UO_2815 (O_2815,N_20658,N_24935);
nor UO_2816 (O_2816,N_23680,N_20246);
nor UO_2817 (O_2817,N_24444,N_22008);
or UO_2818 (O_2818,N_23189,N_22314);
nand UO_2819 (O_2819,N_20423,N_20579);
and UO_2820 (O_2820,N_22275,N_21781);
nor UO_2821 (O_2821,N_20664,N_21727);
and UO_2822 (O_2822,N_22722,N_24385);
or UO_2823 (O_2823,N_22983,N_22190);
and UO_2824 (O_2824,N_24997,N_20511);
and UO_2825 (O_2825,N_21187,N_21613);
and UO_2826 (O_2826,N_23800,N_22563);
or UO_2827 (O_2827,N_24942,N_22664);
and UO_2828 (O_2828,N_21519,N_20799);
xor UO_2829 (O_2829,N_20883,N_21877);
nor UO_2830 (O_2830,N_20603,N_20973);
nor UO_2831 (O_2831,N_21944,N_24451);
or UO_2832 (O_2832,N_23145,N_20485);
and UO_2833 (O_2833,N_21525,N_22245);
or UO_2834 (O_2834,N_21641,N_23479);
nor UO_2835 (O_2835,N_20472,N_24630);
and UO_2836 (O_2836,N_20294,N_23364);
nor UO_2837 (O_2837,N_24740,N_20671);
nand UO_2838 (O_2838,N_21016,N_23377);
or UO_2839 (O_2839,N_23288,N_23132);
or UO_2840 (O_2840,N_21529,N_24377);
nor UO_2841 (O_2841,N_22965,N_21830);
or UO_2842 (O_2842,N_23725,N_24366);
or UO_2843 (O_2843,N_23923,N_21739);
or UO_2844 (O_2844,N_24011,N_23991);
and UO_2845 (O_2845,N_23040,N_24355);
nand UO_2846 (O_2846,N_23645,N_22783);
xnor UO_2847 (O_2847,N_22693,N_23358);
nor UO_2848 (O_2848,N_20781,N_23010);
nor UO_2849 (O_2849,N_24993,N_23425);
and UO_2850 (O_2850,N_23670,N_23978);
or UO_2851 (O_2851,N_23176,N_21767);
xor UO_2852 (O_2852,N_24828,N_24122);
nand UO_2853 (O_2853,N_23767,N_22565);
and UO_2854 (O_2854,N_20676,N_20026);
xnor UO_2855 (O_2855,N_23548,N_22703);
or UO_2856 (O_2856,N_22134,N_21405);
xor UO_2857 (O_2857,N_24295,N_23457);
xnor UO_2858 (O_2858,N_24855,N_21609);
nor UO_2859 (O_2859,N_21703,N_21205);
and UO_2860 (O_2860,N_24508,N_20552);
and UO_2861 (O_2861,N_23550,N_22421);
nand UO_2862 (O_2862,N_22984,N_22528);
xnor UO_2863 (O_2863,N_24000,N_24182);
xnor UO_2864 (O_2864,N_22876,N_23904);
nand UO_2865 (O_2865,N_21458,N_22535);
nand UO_2866 (O_2866,N_20683,N_24849);
and UO_2867 (O_2867,N_21292,N_20653);
xor UO_2868 (O_2868,N_20690,N_20984);
and UO_2869 (O_2869,N_21622,N_24722);
nor UO_2870 (O_2870,N_21968,N_22485);
and UO_2871 (O_2871,N_23123,N_23342);
xor UO_2872 (O_2872,N_23985,N_21951);
nand UO_2873 (O_2873,N_24382,N_21888);
or UO_2874 (O_2874,N_22329,N_20354);
nor UO_2875 (O_2875,N_24099,N_24796);
xnor UO_2876 (O_2876,N_21677,N_22621);
nand UO_2877 (O_2877,N_22618,N_20836);
xnor UO_2878 (O_2878,N_24538,N_22698);
or UO_2879 (O_2879,N_22526,N_21836);
nor UO_2880 (O_2880,N_24229,N_23261);
nand UO_2881 (O_2881,N_23250,N_24288);
xnor UO_2882 (O_2882,N_24907,N_21688);
and UO_2883 (O_2883,N_21023,N_23540);
or UO_2884 (O_2884,N_24442,N_21271);
nor UO_2885 (O_2885,N_23464,N_23156);
xnor UO_2886 (O_2886,N_24079,N_23171);
and UO_2887 (O_2887,N_24480,N_22013);
nor UO_2888 (O_2888,N_24369,N_21194);
or UO_2889 (O_2889,N_22571,N_22557);
nor UO_2890 (O_2890,N_22447,N_20320);
nor UO_2891 (O_2891,N_23108,N_22959);
or UO_2892 (O_2892,N_24529,N_22583);
nand UO_2893 (O_2893,N_22629,N_24084);
xnor UO_2894 (O_2894,N_23458,N_24250);
xnor UO_2895 (O_2895,N_21012,N_23243);
nand UO_2896 (O_2896,N_24931,N_23583);
nor UO_2897 (O_2897,N_24830,N_24579);
or UO_2898 (O_2898,N_21244,N_24384);
nand UO_2899 (O_2899,N_22633,N_24091);
xor UO_2900 (O_2900,N_24887,N_24773);
or UO_2901 (O_2901,N_22360,N_21547);
nand UO_2902 (O_2902,N_24737,N_23736);
xor UO_2903 (O_2903,N_23025,N_22750);
xnor UO_2904 (O_2904,N_22978,N_21374);
nor UO_2905 (O_2905,N_22766,N_24162);
nand UO_2906 (O_2906,N_20115,N_23821);
or UO_2907 (O_2907,N_23824,N_21033);
nor UO_2908 (O_2908,N_22442,N_23462);
nor UO_2909 (O_2909,N_21358,N_20061);
nand UO_2910 (O_2910,N_21709,N_20592);
and UO_2911 (O_2911,N_20862,N_20418);
nor UO_2912 (O_2912,N_22967,N_21196);
nor UO_2913 (O_2913,N_21478,N_21459);
nand UO_2914 (O_2914,N_21695,N_22449);
or UO_2915 (O_2915,N_24356,N_23652);
and UO_2916 (O_2916,N_20890,N_20220);
nand UO_2917 (O_2917,N_23077,N_23683);
nand UO_2918 (O_2918,N_23943,N_21218);
nand UO_2919 (O_2919,N_24328,N_24690);
or UO_2920 (O_2920,N_22139,N_21169);
xnor UO_2921 (O_2921,N_22508,N_21771);
nand UO_2922 (O_2922,N_20553,N_21035);
xor UO_2923 (O_2923,N_20635,N_20584);
nand UO_2924 (O_2924,N_21033,N_21645);
nor UO_2925 (O_2925,N_22025,N_23703);
nor UO_2926 (O_2926,N_21585,N_21592);
and UO_2927 (O_2927,N_21141,N_24645);
and UO_2928 (O_2928,N_22543,N_23311);
xor UO_2929 (O_2929,N_24081,N_24457);
or UO_2930 (O_2930,N_20234,N_22784);
and UO_2931 (O_2931,N_22203,N_21785);
xor UO_2932 (O_2932,N_21380,N_22334);
nor UO_2933 (O_2933,N_21539,N_21809);
nand UO_2934 (O_2934,N_20171,N_21586);
nor UO_2935 (O_2935,N_21346,N_20627);
or UO_2936 (O_2936,N_21583,N_24450);
xor UO_2937 (O_2937,N_20162,N_20787);
nor UO_2938 (O_2938,N_21301,N_21807);
nand UO_2939 (O_2939,N_20125,N_21463);
nand UO_2940 (O_2940,N_24513,N_24012);
nor UO_2941 (O_2941,N_23513,N_20214);
xnor UO_2942 (O_2942,N_23422,N_22946);
nand UO_2943 (O_2943,N_20935,N_21970);
nand UO_2944 (O_2944,N_24995,N_21461);
xor UO_2945 (O_2945,N_21423,N_22869);
and UO_2946 (O_2946,N_24796,N_20470);
xor UO_2947 (O_2947,N_23534,N_21618);
nand UO_2948 (O_2948,N_23369,N_24421);
nor UO_2949 (O_2949,N_24276,N_20322);
or UO_2950 (O_2950,N_23414,N_22528);
and UO_2951 (O_2951,N_20875,N_20387);
or UO_2952 (O_2952,N_24518,N_21996);
nor UO_2953 (O_2953,N_22315,N_23808);
nor UO_2954 (O_2954,N_21266,N_23623);
nor UO_2955 (O_2955,N_21504,N_21774);
nand UO_2956 (O_2956,N_23016,N_21290);
xor UO_2957 (O_2957,N_23935,N_21046);
nand UO_2958 (O_2958,N_21982,N_24730);
or UO_2959 (O_2959,N_22611,N_21923);
and UO_2960 (O_2960,N_21393,N_24826);
and UO_2961 (O_2961,N_21401,N_21846);
xor UO_2962 (O_2962,N_24584,N_22322);
xnor UO_2963 (O_2963,N_23028,N_24142);
or UO_2964 (O_2964,N_20472,N_22632);
xnor UO_2965 (O_2965,N_23924,N_20670);
and UO_2966 (O_2966,N_23927,N_23082);
or UO_2967 (O_2967,N_23065,N_20420);
xnor UO_2968 (O_2968,N_24524,N_24552);
and UO_2969 (O_2969,N_23653,N_22315);
nand UO_2970 (O_2970,N_24935,N_24561);
or UO_2971 (O_2971,N_23148,N_22986);
and UO_2972 (O_2972,N_22981,N_20277);
nor UO_2973 (O_2973,N_24052,N_20697);
and UO_2974 (O_2974,N_23944,N_24246);
or UO_2975 (O_2975,N_21461,N_22926);
or UO_2976 (O_2976,N_20182,N_22608);
xor UO_2977 (O_2977,N_23945,N_20022);
nand UO_2978 (O_2978,N_24031,N_24026);
xor UO_2979 (O_2979,N_20746,N_22436);
nand UO_2980 (O_2980,N_20841,N_24693);
nor UO_2981 (O_2981,N_24740,N_20850);
or UO_2982 (O_2982,N_23836,N_20206);
nor UO_2983 (O_2983,N_21665,N_23180);
and UO_2984 (O_2984,N_20686,N_24097);
nor UO_2985 (O_2985,N_21716,N_23111);
or UO_2986 (O_2986,N_23171,N_21836);
nor UO_2987 (O_2987,N_22374,N_24512);
or UO_2988 (O_2988,N_22586,N_22959);
xor UO_2989 (O_2989,N_22591,N_20477);
nor UO_2990 (O_2990,N_22886,N_22804);
nor UO_2991 (O_2991,N_23122,N_23680);
nand UO_2992 (O_2992,N_23121,N_21624);
nor UO_2993 (O_2993,N_21600,N_23490);
nor UO_2994 (O_2994,N_20020,N_21345);
or UO_2995 (O_2995,N_20941,N_24875);
nand UO_2996 (O_2996,N_24873,N_23841);
and UO_2997 (O_2997,N_23110,N_24161);
nand UO_2998 (O_2998,N_20553,N_22466);
or UO_2999 (O_2999,N_22664,N_22869);
endmodule