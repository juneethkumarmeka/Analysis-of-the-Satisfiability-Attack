module basic_500_3000_500_15_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_344,In_298);
or U1 (N_1,In_198,In_309);
nand U2 (N_2,In_53,In_85);
nand U3 (N_3,In_318,In_362);
and U4 (N_4,In_444,In_72);
nand U5 (N_5,In_329,In_285);
nand U6 (N_6,In_189,In_268);
or U7 (N_7,In_414,In_252);
nand U8 (N_8,In_98,In_185);
or U9 (N_9,In_417,In_325);
nand U10 (N_10,In_293,In_308);
or U11 (N_11,In_391,In_431);
xor U12 (N_12,In_256,In_33);
and U13 (N_13,In_240,In_234);
nand U14 (N_14,In_123,In_388);
and U15 (N_15,In_21,In_369);
nor U16 (N_16,In_255,In_379);
nand U17 (N_17,In_287,In_399);
nor U18 (N_18,In_222,In_387);
or U19 (N_19,In_310,In_106);
nand U20 (N_20,In_415,In_396);
nand U21 (N_21,In_109,In_15);
or U22 (N_22,In_233,In_457);
nand U23 (N_23,In_436,In_407);
nand U24 (N_24,In_342,In_131);
nand U25 (N_25,In_251,In_94);
nand U26 (N_26,In_420,In_341);
and U27 (N_27,In_257,In_367);
nand U28 (N_28,In_317,In_182);
and U29 (N_29,In_156,In_348);
and U30 (N_30,In_52,In_110);
and U31 (N_31,In_203,In_32);
nor U32 (N_32,In_258,In_118);
or U33 (N_33,In_90,In_193);
and U34 (N_34,In_459,In_354);
nor U35 (N_35,In_449,In_35);
and U36 (N_36,In_475,In_116);
or U37 (N_37,In_401,In_84);
and U38 (N_38,In_199,In_357);
or U39 (N_39,In_191,In_400);
and U40 (N_40,In_147,In_439);
nor U41 (N_41,In_454,In_280);
or U42 (N_42,In_478,In_76);
nand U43 (N_43,In_276,In_340);
and U44 (N_44,In_266,In_167);
and U45 (N_45,In_321,In_187);
nand U46 (N_46,In_212,In_411);
or U47 (N_47,In_283,In_181);
or U48 (N_48,In_350,In_159);
and U49 (N_49,In_278,In_225);
nand U50 (N_50,In_305,In_81);
or U51 (N_51,In_75,In_382);
and U52 (N_52,In_179,In_103);
nand U53 (N_53,In_370,In_485);
and U54 (N_54,In_9,In_323);
and U55 (N_55,In_270,In_300);
nor U56 (N_56,In_465,In_163);
and U57 (N_57,In_200,In_107);
and U58 (N_58,In_336,In_339);
or U59 (N_59,In_334,In_490);
nand U60 (N_60,In_219,In_92);
nor U61 (N_61,In_237,In_441);
nand U62 (N_62,In_78,In_172);
nand U63 (N_63,In_289,In_104);
nand U64 (N_64,In_260,In_2);
nor U65 (N_65,In_429,In_442);
and U66 (N_66,In_322,In_26);
nor U67 (N_67,In_450,In_236);
nor U68 (N_68,In_499,In_176);
nor U69 (N_69,In_5,In_223);
nor U70 (N_70,In_67,In_360);
xnor U71 (N_71,In_139,In_273);
and U72 (N_72,In_148,In_169);
nand U73 (N_73,In_271,In_132);
nand U74 (N_74,In_101,In_385);
or U75 (N_75,In_13,In_453);
or U76 (N_76,In_166,In_384);
nand U77 (N_77,In_41,In_218);
and U78 (N_78,In_142,In_297);
and U79 (N_79,In_491,In_445);
nand U80 (N_80,In_313,In_238);
nand U81 (N_81,In_291,In_57);
and U82 (N_82,In_31,In_144);
nor U83 (N_83,In_58,In_428);
nand U84 (N_84,In_375,In_358);
nand U85 (N_85,In_54,In_229);
nor U86 (N_86,In_351,In_468);
or U87 (N_87,In_173,In_122);
xor U88 (N_88,In_8,In_365);
nor U89 (N_89,In_483,In_488);
nor U90 (N_90,In_83,In_346);
or U91 (N_91,In_279,In_331);
and U92 (N_92,In_37,In_267);
nor U93 (N_93,In_112,In_239);
and U94 (N_94,In_27,In_0);
nand U95 (N_95,In_18,In_337);
or U96 (N_96,In_17,In_363);
nand U97 (N_97,In_183,In_143);
nand U98 (N_98,In_497,In_250);
nor U99 (N_99,In_335,In_42);
and U100 (N_100,In_154,In_220);
nor U101 (N_101,In_460,In_25);
and U102 (N_102,In_63,In_302);
and U103 (N_103,In_77,In_467);
and U104 (N_104,In_338,In_494);
nand U105 (N_105,In_412,In_416);
nand U106 (N_106,In_146,In_286);
and U107 (N_107,In_440,In_97);
or U108 (N_108,In_165,In_205);
or U109 (N_109,In_424,In_192);
nor U110 (N_110,In_277,In_319);
nor U111 (N_111,In_421,In_214);
or U112 (N_112,In_153,In_418);
nand U113 (N_113,In_7,In_190);
or U114 (N_114,In_152,In_23);
or U115 (N_115,In_11,In_175);
nor U116 (N_116,In_96,In_221);
or U117 (N_117,In_364,In_60);
or U118 (N_118,In_217,In_327);
and U119 (N_119,In_133,In_356);
nand U120 (N_120,In_324,In_315);
nor U121 (N_121,In_117,In_484);
and U122 (N_122,In_487,In_68);
nor U123 (N_123,In_311,In_208);
and U124 (N_124,In_119,In_177);
nor U125 (N_125,In_432,In_125);
nand U126 (N_126,In_4,In_393);
or U127 (N_127,In_374,In_377);
or U128 (N_128,In_381,In_126);
or U129 (N_129,In_124,In_366);
nor U130 (N_130,In_188,In_12);
nand U131 (N_131,In_137,In_292);
nor U132 (N_132,In_328,In_409);
xnor U133 (N_133,In_332,In_207);
or U134 (N_134,In_56,In_368);
or U135 (N_135,In_426,In_66);
nand U136 (N_136,In_88,In_473);
nor U137 (N_137,In_171,In_64);
nor U138 (N_138,In_51,In_19);
xor U139 (N_139,In_435,In_194);
and U140 (N_140,In_86,In_326);
nand U141 (N_141,In_113,In_46);
nor U142 (N_142,In_69,In_406);
nand U143 (N_143,In_299,In_20);
or U144 (N_144,In_437,In_231);
nand U145 (N_145,In_296,In_145);
or U146 (N_146,In_355,In_290);
and U147 (N_147,In_164,In_30);
nand U148 (N_148,In_455,In_71);
nand U149 (N_149,In_288,In_130);
nand U150 (N_150,In_247,In_269);
or U151 (N_151,In_433,In_245);
or U152 (N_152,In_38,In_28);
and U153 (N_153,In_249,In_330);
nor U154 (N_154,In_272,In_446);
and U155 (N_155,In_474,In_486);
or U156 (N_156,In_448,In_158);
or U157 (N_157,In_394,In_472);
nor U158 (N_158,In_482,In_34);
nand U159 (N_159,In_496,In_295);
nand U160 (N_160,In_99,In_253);
nor U161 (N_161,In_134,In_39);
or U162 (N_162,In_135,In_498);
or U163 (N_163,In_95,In_157);
or U164 (N_164,In_371,In_456);
or U165 (N_165,In_306,In_349);
nand U166 (N_166,In_423,In_49);
nor U167 (N_167,In_359,In_178);
and U168 (N_168,In_162,In_211);
nor U169 (N_169,In_136,In_138);
and U170 (N_170,In_241,In_43);
nor U171 (N_171,In_216,In_452);
or U172 (N_172,In_438,In_224);
nor U173 (N_173,In_151,In_372);
or U174 (N_174,In_481,In_392);
or U175 (N_175,In_89,In_170);
and U176 (N_176,In_470,In_378);
or U177 (N_177,In_150,In_24);
nor U178 (N_178,In_74,In_413);
or U179 (N_179,In_422,In_471);
or U180 (N_180,In_65,In_186);
or U181 (N_181,In_195,In_48);
or U182 (N_182,In_235,In_202);
and U183 (N_183,In_140,In_206);
or U184 (N_184,In_248,In_73);
and U185 (N_185,In_59,In_149);
and U186 (N_186,In_463,In_93);
nand U187 (N_187,In_303,In_213);
nor U188 (N_188,In_476,In_102);
and U189 (N_189,In_204,In_201);
and U190 (N_190,In_114,In_232);
and U191 (N_191,In_210,In_160);
and U192 (N_192,In_398,In_121);
nand U193 (N_193,In_3,In_307);
nor U194 (N_194,In_373,In_469);
or U195 (N_195,In_264,In_492);
or U196 (N_196,In_87,In_294);
and U197 (N_197,In_120,In_108);
and U198 (N_198,In_79,In_129);
or U199 (N_199,In_480,In_495);
and U200 (N_200,N_22,In_447);
nand U201 (N_201,N_101,N_145);
nand U202 (N_202,In_29,N_191);
or U203 (N_203,N_59,N_100);
nor U204 (N_204,In_380,N_12);
nand U205 (N_205,In_489,In_389);
nor U206 (N_206,In_40,N_155);
nor U207 (N_207,N_54,N_109);
and U208 (N_208,N_30,N_131);
or U209 (N_209,N_68,N_80);
or U210 (N_210,N_7,In_314);
nor U211 (N_211,In_47,N_2);
nor U212 (N_212,N_50,In_62);
and U213 (N_213,N_94,N_38);
or U214 (N_214,In_312,N_64);
and U215 (N_215,In_259,In_242);
and U216 (N_216,N_127,In_353);
and U217 (N_217,N_24,N_110);
or U218 (N_218,N_129,In_262);
and U219 (N_219,In_451,N_157);
nand U220 (N_220,N_0,N_105);
nand U221 (N_221,In_184,N_161);
or U222 (N_222,N_188,In_383);
nand U223 (N_223,In_50,In_347);
and U224 (N_224,N_90,In_461);
and U225 (N_225,N_190,N_153);
nor U226 (N_226,N_160,N_196);
or U227 (N_227,N_11,N_88);
nor U228 (N_228,In_410,N_20);
nand U229 (N_229,In_282,N_171);
or U230 (N_230,N_185,N_163);
and U231 (N_231,N_8,N_198);
nor U232 (N_232,N_3,N_169);
and U233 (N_233,In_361,N_35);
or U234 (N_234,In_434,In_91);
nand U235 (N_235,N_76,N_149);
or U236 (N_236,In_284,N_26);
or U237 (N_237,N_167,N_132);
nor U238 (N_238,In_301,In_403);
and U239 (N_239,N_115,In_390);
nor U240 (N_240,N_58,N_92);
nand U241 (N_241,N_125,N_21);
nor U242 (N_242,N_174,N_87);
and U243 (N_243,N_77,In_493);
or U244 (N_244,N_23,In_226);
nor U245 (N_245,N_83,In_45);
or U246 (N_246,In_376,N_166);
or U247 (N_247,In_333,N_95);
nand U248 (N_248,N_122,In_386);
and U249 (N_249,In_477,In_100);
and U250 (N_250,In_479,N_195);
or U251 (N_251,In_196,N_52);
nor U252 (N_252,N_78,In_243);
nor U253 (N_253,N_170,N_85);
or U254 (N_254,N_107,In_111);
nor U255 (N_255,In_16,N_61);
nor U256 (N_256,N_67,N_71);
nand U257 (N_257,N_1,N_173);
and U258 (N_258,N_74,N_151);
nor U259 (N_259,N_47,In_61);
nor U260 (N_260,N_194,In_80);
or U261 (N_261,In_70,In_209);
and U262 (N_262,In_404,In_425);
nor U263 (N_263,N_126,N_108);
and U264 (N_264,In_316,N_27);
nor U265 (N_265,In_105,N_103);
nand U266 (N_266,In_464,N_82);
and U267 (N_267,N_102,N_84);
and U268 (N_268,N_178,N_45);
nor U269 (N_269,N_13,N_25);
and U270 (N_270,N_33,N_57);
and U271 (N_271,N_4,N_159);
nand U272 (N_272,N_139,N_98);
or U273 (N_273,N_53,N_97);
nor U274 (N_274,In_395,N_133);
nor U275 (N_275,In_14,N_147);
nand U276 (N_276,N_42,In_419);
and U277 (N_277,N_96,In_82);
or U278 (N_278,N_31,N_89);
or U279 (N_279,In_244,N_136);
and U280 (N_280,In_155,In_180);
and U281 (N_281,N_135,N_120);
nor U282 (N_282,N_179,In_128);
nand U283 (N_283,N_168,N_37);
or U284 (N_284,N_43,N_62);
nor U285 (N_285,N_73,N_143);
and U286 (N_286,N_142,In_430);
or U287 (N_287,N_17,N_162);
nand U288 (N_288,N_65,N_10);
nand U289 (N_289,In_1,N_49);
nand U290 (N_290,N_141,N_18);
or U291 (N_291,In_345,N_181);
nand U292 (N_292,N_29,N_177);
nand U293 (N_293,N_158,N_119);
or U294 (N_294,In_405,In_343);
or U295 (N_295,N_199,N_14);
and U296 (N_296,N_28,In_462);
nor U297 (N_297,N_140,In_228);
nor U298 (N_298,N_113,In_227);
nor U299 (N_299,N_69,N_79);
nor U300 (N_300,N_99,In_397);
or U301 (N_301,N_187,N_180);
nand U302 (N_302,N_154,N_152);
nand U303 (N_303,N_128,In_320);
nor U304 (N_304,N_172,N_111);
or U305 (N_305,N_114,In_261);
nor U306 (N_306,N_144,N_32);
nor U307 (N_307,N_91,In_168);
nor U308 (N_308,N_189,N_106);
or U309 (N_309,N_86,N_75);
and U310 (N_310,In_275,N_72);
nand U311 (N_311,In_127,N_60);
and U312 (N_312,In_22,N_176);
nor U313 (N_313,N_104,In_10);
and U314 (N_314,In_36,N_15);
and U315 (N_315,In_6,N_70);
and U316 (N_316,N_164,In_352);
nand U317 (N_317,In_281,In_55);
nor U318 (N_318,N_156,N_112);
nand U319 (N_319,N_36,N_5);
and U320 (N_320,N_44,N_137);
and U321 (N_321,N_186,In_458);
nand U322 (N_322,In_230,N_6);
nor U323 (N_323,In_246,N_93);
and U324 (N_324,N_146,N_39);
or U325 (N_325,N_183,In_254);
nor U326 (N_326,N_150,N_56);
nand U327 (N_327,N_16,In_263);
nor U328 (N_328,N_197,N_81);
or U329 (N_329,N_41,N_40);
nand U330 (N_330,N_121,N_124);
nor U331 (N_331,In_466,N_9);
nand U332 (N_332,N_51,In_265);
or U333 (N_333,N_116,N_123);
nor U334 (N_334,In_44,In_115);
xor U335 (N_335,In_141,In_304);
and U336 (N_336,N_117,N_184);
and U337 (N_337,N_55,N_175);
or U338 (N_338,N_46,N_63);
or U339 (N_339,In_443,In_408);
and U340 (N_340,N_134,N_192);
nand U341 (N_341,In_402,N_19);
or U342 (N_342,In_427,N_182);
or U343 (N_343,N_138,N_148);
nand U344 (N_344,In_215,In_197);
nand U345 (N_345,In_274,N_165);
nand U346 (N_346,N_118,N_193);
nor U347 (N_347,N_66,In_174);
or U348 (N_348,In_161,N_130);
or U349 (N_349,N_34,N_48);
and U350 (N_350,N_15,N_112);
and U351 (N_351,N_157,N_149);
nor U352 (N_352,N_90,N_22);
nor U353 (N_353,N_12,In_168);
or U354 (N_354,N_51,In_47);
xor U355 (N_355,In_464,N_167);
or U356 (N_356,In_262,N_50);
xor U357 (N_357,In_100,In_425);
xnor U358 (N_358,N_127,N_193);
and U359 (N_359,N_52,In_397);
nand U360 (N_360,N_49,In_259);
and U361 (N_361,In_493,N_106);
nor U362 (N_362,N_0,In_345);
nand U363 (N_363,N_119,N_22);
nor U364 (N_364,N_58,In_61);
nand U365 (N_365,N_115,In_284);
and U366 (N_366,N_83,N_85);
and U367 (N_367,N_32,N_17);
nand U368 (N_368,N_113,N_16);
and U369 (N_369,In_230,N_111);
nor U370 (N_370,In_127,N_74);
or U371 (N_371,In_36,N_104);
nor U372 (N_372,In_301,N_176);
and U373 (N_373,N_93,N_148);
nor U374 (N_374,In_115,N_61);
or U375 (N_375,In_376,N_153);
and U376 (N_376,N_2,N_166);
and U377 (N_377,N_3,In_244);
nand U378 (N_378,N_198,N_33);
nor U379 (N_379,N_104,N_29);
or U380 (N_380,N_109,N_17);
nor U381 (N_381,N_120,N_21);
nor U382 (N_382,N_63,N_38);
and U383 (N_383,In_320,N_139);
nand U384 (N_384,N_87,In_168);
nor U385 (N_385,In_397,N_178);
nand U386 (N_386,N_63,In_376);
or U387 (N_387,In_128,N_97);
and U388 (N_388,N_144,N_149);
nand U389 (N_389,In_61,In_443);
and U390 (N_390,In_47,N_126);
or U391 (N_391,In_312,N_176);
xor U392 (N_392,N_46,N_2);
and U393 (N_393,N_54,N_147);
and U394 (N_394,N_53,N_135);
or U395 (N_395,In_115,N_193);
nor U396 (N_396,N_93,N_36);
or U397 (N_397,N_166,In_443);
nor U398 (N_398,N_175,In_361);
nand U399 (N_399,In_55,In_259);
nor U400 (N_400,N_397,N_233);
nand U401 (N_401,N_213,N_364);
or U402 (N_402,N_373,N_349);
nor U403 (N_403,N_235,N_234);
or U404 (N_404,N_289,N_273);
or U405 (N_405,N_225,N_293);
and U406 (N_406,N_308,N_219);
nor U407 (N_407,N_292,N_276);
nand U408 (N_408,N_228,N_386);
or U409 (N_409,N_328,N_361);
nand U410 (N_410,N_326,N_329);
and U411 (N_411,N_313,N_348);
or U412 (N_412,N_223,N_330);
or U413 (N_413,N_218,N_227);
nor U414 (N_414,N_217,N_238);
and U415 (N_415,N_256,N_381);
nor U416 (N_416,N_239,N_297);
nor U417 (N_417,N_271,N_207);
nor U418 (N_418,N_291,N_378);
nor U419 (N_419,N_316,N_254);
nor U420 (N_420,N_312,N_251);
and U421 (N_421,N_353,N_355);
or U422 (N_422,N_249,N_319);
nor U423 (N_423,N_206,N_241);
nand U424 (N_424,N_321,N_237);
and U425 (N_425,N_243,N_315);
nand U426 (N_426,N_242,N_262);
and U427 (N_427,N_352,N_248);
or U428 (N_428,N_377,N_382);
and U429 (N_429,N_310,N_332);
nor U430 (N_430,N_286,N_287);
or U431 (N_431,N_222,N_296);
or U432 (N_432,N_362,N_246);
nor U433 (N_433,N_343,N_285);
and U434 (N_434,N_359,N_277);
or U435 (N_435,N_281,N_224);
nand U436 (N_436,N_300,N_302);
and U437 (N_437,N_269,N_270);
nor U438 (N_438,N_365,N_320);
nor U439 (N_439,N_267,N_324);
and U440 (N_440,N_356,N_395);
and U441 (N_441,N_205,N_384);
and U442 (N_442,N_389,N_396);
or U443 (N_443,N_290,N_317);
nor U444 (N_444,N_393,N_230);
or U445 (N_445,N_259,N_226);
nor U446 (N_446,N_379,N_390);
and U447 (N_447,N_357,N_231);
and U448 (N_448,N_311,N_360);
nor U449 (N_449,N_376,N_268);
nor U450 (N_450,N_342,N_331);
or U451 (N_451,N_266,N_301);
nand U452 (N_452,N_265,N_275);
nand U453 (N_453,N_383,N_354);
nand U454 (N_454,N_298,N_372);
and U455 (N_455,N_264,N_366);
and U456 (N_456,N_305,N_398);
nor U457 (N_457,N_337,N_303);
nor U458 (N_458,N_318,N_334);
nor U459 (N_459,N_229,N_261);
or U460 (N_460,N_388,N_347);
or U461 (N_461,N_274,N_351);
and U462 (N_462,N_333,N_279);
nand U463 (N_463,N_304,N_341);
or U464 (N_464,N_363,N_255);
nand U465 (N_465,N_250,N_215);
nand U466 (N_466,N_232,N_212);
or U467 (N_467,N_247,N_323);
nor U468 (N_468,N_209,N_336);
or U469 (N_469,N_385,N_252);
nor U470 (N_470,N_208,N_201);
and U471 (N_471,N_371,N_263);
nor U472 (N_472,N_392,N_210);
nor U473 (N_473,N_220,N_387);
nor U474 (N_474,N_200,N_374);
and U475 (N_475,N_367,N_283);
nand U476 (N_476,N_391,N_309);
or U477 (N_477,N_399,N_204);
or U478 (N_478,N_245,N_370);
and U479 (N_479,N_272,N_294);
and U480 (N_480,N_350,N_258);
nand U481 (N_481,N_394,N_335);
or U482 (N_482,N_380,N_221);
and U483 (N_483,N_280,N_244);
and U484 (N_484,N_202,N_375);
nor U485 (N_485,N_346,N_327);
nand U486 (N_486,N_295,N_284);
or U487 (N_487,N_358,N_211);
nor U488 (N_488,N_203,N_369);
and U489 (N_489,N_278,N_288);
or U490 (N_490,N_306,N_339);
nor U491 (N_491,N_257,N_325);
nand U492 (N_492,N_344,N_282);
nor U493 (N_493,N_340,N_236);
and U494 (N_494,N_253,N_307);
nor U495 (N_495,N_299,N_240);
nor U496 (N_496,N_214,N_322);
nor U497 (N_497,N_345,N_260);
nand U498 (N_498,N_368,N_314);
or U499 (N_499,N_338,N_216);
nor U500 (N_500,N_340,N_247);
and U501 (N_501,N_376,N_299);
and U502 (N_502,N_306,N_290);
nor U503 (N_503,N_243,N_384);
or U504 (N_504,N_250,N_334);
nand U505 (N_505,N_329,N_300);
nand U506 (N_506,N_367,N_291);
or U507 (N_507,N_298,N_267);
and U508 (N_508,N_349,N_383);
nand U509 (N_509,N_331,N_370);
and U510 (N_510,N_222,N_324);
nand U511 (N_511,N_257,N_383);
nor U512 (N_512,N_392,N_310);
or U513 (N_513,N_380,N_286);
nor U514 (N_514,N_267,N_333);
nand U515 (N_515,N_330,N_352);
or U516 (N_516,N_219,N_227);
or U517 (N_517,N_361,N_284);
nor U518 (N_518,N_346,N_320);
and U519 (N_519,N_297,N_252);
nor U520 (N_520,N_206,N_229);
nor U521 (N_521,N_338,N_373);
and U522 (N_522,N_289,N_261);
nand U523 (N_523,N_239,N_242);
or U524 (N_524,N_204,N_235);
nand U525 (N_525,N_321,N_269);
or U526 (N_526,N_309,N_332);
nand U527 (N_527,N_233,N_246);
nor U528 (N_528,N_389,N_305);
or U529 (N_529,N_309,N_263);
or U530 (N_530,N_366,N_319);
nor U531 (N_531,N_377,N_317);
or U532 (N_532,N_279,N_254);
nand U533 (N_533,N_273,N_396);
nor U534 (N_534,N_200,N_242);
nand U535 (N_535,N_273,N_357);
nor U536 (N_536,N_307,N_361);
nand U537 (N_537,N_350,N_307);
and U538 (N_538,N_212,N_391);
nand U539 (N_539,N_390,N_284);
and U540 (N_540,N_239,N_322);
nand U541 (N_541,N_251,N_358);
nor U542 (N_542,N_222,N_287);
or U543 (N_543,N_239,N_259);
or U544 (N_544,N_317,N_368);
and U545 (N_545,N_336,N_348);
or U546 (N_546,N_339,N_238);
nand U547 (N_547,N_368,N_204);
nand U548 (N_548,N_396,N_301);
and U549 (N_549,N_320,N_349);
nand U550 (N_550,N_214,N_268);
and U551 (N_551,N_313,N_377);
or U552 (N_552,N_389,N_283);
nor U553 (N_553,N_287,N_326);
or U554 (N_554,N_217,N_373);
and U555 (N_555,N_267,N_349);
or U556 (N_556,N_250,N_253);
nor U557 (N_557,N_341,N_319);
or U558 (N_558,N_344,N_361);
and U559 (N_559,N_393,N_311);
or U560 (N_560,N_264,N_208);
or U561 (N_561,N_279,N_365);
xor U562 (N_562,N_257,N_232);
and U563 (N_563,N_248,N_385);
and U564 (N_564,N_268,N_339);
nand U565 (N_565,N_259,N_298);
nand U566 (N_566,N_340,N_208);
or U567 (N_567,N_207,N_247);
nand U568 (N_568,N_385,N_378);
or U569 (N_569,N_315,N_296);
nor U570 (N_570,N_365,N_358);
nand U571 (N_571,N_200,N_376);
nor U572 (N_572,N_344,N_218);
or U573 (N_573,N_262,N_312);
or U574 (N_574,N_333,N_260);
nor U575 (N_575,N_323,N_217);
nand U576 (N_576,N_261,N_226);
nor U577 (N_577,N_351,N_328);
nand U578 (N_578,N_289,N_387);
nor U579 (N_579,N_256,N_278);
nor U580 (N_580,N_386,N_271);
nand U581 (N_581,N_215,N_369);
nor U582 (N_582,N_395,N_368);
nand U583 (N_583,N_341,N_376);
nor U584 (N_584,N_331,N_349);
nor U585 (N_585,N_375,N_254);
and U586 (N_586,N_355,N_200);
nor U587 (N_587,N_305,N_207);
nand U588 (N_588,N_217,N_308);
nand U589 (N_589,N_206,N_310);
and U590 (N_590,N_266,N_233);
nand U591 (N_591,N_214,N_376);
or U592 (N_592,N_263,N_380);
nor U593 (N_593,N_379,N_344);
nor U594 (N_594,N_359,N_343);
and U595 (N_595,N_397,N_230);
or U596 (N_596,N_248,N_204);
and U597 (N_597,N_356,N_248);
and U598 (N_598,N_345,N_378);
nor U599 (N_599,N_211,N_249);
nand U600 (N_600,N_416,N_468);
or U601 (N_601,N_433,N_592);
or U602 (N_602,N_409,N_429);
nand U603 (N_603,N_589,N_505);
nor U604 (N_604,N_400,N_462);
nor U605 (N_605,N_483,N_456);
nor U606 (N_606,N_594,N_586);
and U607 (N_607,N_434,N_516);
and U608 (N_608,N_534,N_509);
nand U609 (N_609,N_583,N_442);
nand U610 (N_610,N_437,N_538);
nand U611 (N_611,N_481,N_487);
nor U612 (N_612,N_427,N_501);
or U613 (N_613,N_529,N_474);
and U614 (N_614,N_473,N_493);
and U615 (N_615,N_507,N_447);
and U616 (N_616,N_420,N_565);
or U617 (N_617,N_457,N_441);
or U618 (N_618,N_458,N_494);
and U619 (N_619,N_547,N_557);
nand U620 (N_620,N_504,N_422);
or U621 (N_621,N_552,N_492);
and U622 (N_622,N_524,N_506);
nand U623 (N_623,N_431,N_446);
and U624 (N_624,N_580,N_412);
and U625 (N_625,N_566,N_471);
nand U626 (N_626,N_523,N_593);
or U627 (N_627,N_403,N_485);
nor U628 (N_628,N_528,N_502);
nand U629 (N_629,N_495,N_527);
nand U630 (N_630,N_454,N_448);
or U631 (N_631,N_572,N_450);
and U632 (N_632,N_568,N_533);
or U633 (N_633,N_445,N_575);
nor U634 (N_634,N_556,N_587);
or U635 (N_635,N_436,N_554);
or U636 (N_636,N_408,N_535);
or U637 (N_637,N_512,N_551);
nand U638 (N_638,N_511,N_479);
nor U639 (N_639,N_596,N_496);
and U640 (N_640,N_526,N_497);
and U641 (N_641,N_463,N_590);
or U642 (N_642,N_424,N_548);
nor U643 (N_643,N_561,N_550);
or U644 (N_644,N_537,N_599);
or U645 (N_645,N_449,N_573);
or U646 (N_646,N_542,N_582);
or U647 (N_647,N_521,N_418);
nor U648 (N_648,N_508,N_543);
and U649 (N_649,N_432,N_452);
nor U650 (N_650,N_544,N_540);
nand U651 (N_651,N_419,N_559);
nor U652 (N_652,N_401,N_482);
and U653 (N_653,N_518,N_579);
nand U654 (N_654,N_578,N_480);
nor U655 (N_655,N_574,N_541);
nand U656 (N_656,N_440,N_478);
nor U657 (N_657,N_499,N_539);
nor U658 (N_658,N_571,N_563);
and U659 (N_659,N_466,N_530);
and U660 (N_660,N_555,N_510);
or U661 (N_661,N_549,N_461);
nand U662 (N_662,N_564,N_598);
and U663 (N_663,N_428,N_536);
nor U664 (N_664,N_477,N_414);
nand U665 (N_665,N_489,N_464);
and U666 (N_666,N_570,N_584);
or U667 (N_667,N_460,N_597);
nor U668 (N_668,N_588,N_514);
xnor U669 (N_669,N_577,N_558);
nor U670 (N_670,N_522,N_546);
or U671 (N_671,N_443,N_488);
or U672 (N_672,N_402,N_467);
nor U673 (N_673,N_498,N_595);
and U674 (N_674,N_519,N_435);
nand U675 (N_675,N_425,N_476);
nor U676 (N_676,N_532,N_413);
nand U677 (N_677,N_404,N_439);
or U678 (N_678,N_417,N_455);
and U679 (N_679,N_569,N_517);
or U680 (N_680,N_591,N_438);
nand U681 (N_681,N_513,N_581);
nor U682 (N_682,N_451,N_562);
nor U683 (N_683,N_585,N_531);
and U684 (N_684,N_490,N_426);
nand U685 (N_685,N_444,N_430);
and U686 (N_686,N_453,N_503);
nand U687 (N_687,N_472,N_405);
and U688 (N_688,N_500,N_470);
and U689 (N_689,N_520,N_553);
xor U690 (N_690,N_411,N_576);
or U691 (N_691,N_484,N_525);
nor U692 (N_692,N_491,N_515);
nor U693 (N_693,N_406,N_560);
and U694 (N_694,N_465,N_421);
nand U695 (N_695,N_415,N_475);
nor U696 (N_696,N_423,N_545);
nand U697 (N_697,N_567,N_407);
or U698 (N_698,N_486,N_410);
nand U699 (N_699,N_469,N_459);
nand U700 (N_700,N_414,N_541);
or U701 (N_701,N_430,N_588);
or U702 (N_702,N_558,N_539);
nor U703 (N_703,N_405,N_439);
and U704 (N_704,N_583,N_453);
nor U705 (N_705,N_502,N_533);
or U706 (N_706,N_530,N_562);
nand U707 (N_707,N_580,N_483);
nor U708 (N_708,N_566,N_469);
or U709 (N_709,N_474,N_458);
nand U710 (N_710,N_491,N_462);
or U711 (N_711,N_527,N_419);
or U712 (N_712,N_410,N_560);
or U713 (N_713,N_581,N_457);
nor U714 (N_714,N_534,N_459);
and U715 (N_715,N_463,N_517);
nor U716 (N_716,N_426,N_495);
and U717 (N_717,N_541,N_461);
or U718 (N_718,N_586,N_574);
and U719 (N_719,N_487,N_567);
or U720 (N_720,N_565,N_401);
nand U721 (N_721,N_566,N_420);
nor U722 (N_722,N_473,N_517);
nand U723 (N_723,N_442,N_553);
and U724 (N_724,N_487,N_563);
nand U725 (N_725,N_459,N_415);
nor U726 (N_726,N_423,N_517);
and U727 (N_727,N_538,N_548);
nand U728 (N_728,N_412,N_490);
nor U729 (N_729,N_438,N_512);
or U730 (N_730,N_445,N_473);
or U731 (N_731,N_462,N_466);
nand U732 (N_732,N_473,N_407);
nand U733 (N_733,N_561,N_479);
and U734 (N_734,N_569,N_456);
xor U735 (N_735,N_428,N_449);
nor U736 (N_736,N_533,N_432);
nand U737 (N_737,N_555,N_535);
nand U738 (N_738,N_481,N_550);
and U739 (N_739,N_581,N_485);
nor U740 (N_740,N_460,N_451);
nand U741 (N_741,N_522,N_511);
or U742 (N_742,N_424,N_545);
or U743 (N_743,N_462,N_457);
and U744 (N_744,N_468,N_558);
nand U745 (N_745,N_579,N_516);
nor U746 (N_746,N_461,N_422);
and U747 (N_747,N_550,N_526);
and U748 (N_748,N_482,N_475);
and U749 (N_749,N_450,N_500);
nand U750 (N_750,N_431,N_413);
nand U751 (N_751,N_403,N_597);
nor U752 (N_752,N_586,N_570);
or U753 (N_753,N_505,N_499);
or U754 (N_754,N_427,N_426);
nand U755 (N_755,N_406,N_536);
and U756 (N_756,N_496,N_431);
and U757 (N_757,N_570,N_560);
nand U758 (N_758,N_432,N_502);
and U759 (N_759,N_497,N_588);
nor U760 (N_760,N_445,N_517);
nand U761 (N_761,N_565,N_526);
and U762 (N_762,N_571,N_434);
nand U763 (N_763,N_559,N_565);
nand U764 (N_764,N_580,N_548);
or U765 (N_765,N_429,N_512);
or U766 (N_766,N_472,N_505);
or U767 (N_767,N_556,N_555);
or U768 (N_768,N_541,N_550);
xnor U769 (N_769,N_446,N_551);
nand U770 (N_770,N_550,N_571);
and U771 (N_771,N_598,N_591);
xnor U772 (N_772,N_522,N_540);
nand U773 (N_773,N_595,N_478);
nor U774 (N_774,N_522,N_480);
or U775 (N_775,N_579,N_483);
nor U776 (N_776,N_511,N_493);
or U777 (N_777,N_543,N_563);
nor U778 (N_778,N_517,N_503);
and U779 (N_779,N_561,N_588);
and U780 (N_780,N_435,N_565);
and U781 (N_781,N_465,N_425);
and U782 (N_782,N_518,N_493);
nand U783 (N_783,N_581,N_570);
or U784 (N_784,N_541,N_532);
and U785 (N_785,N_500,N_400);
nand U786 (N_786,N_539,N_442);
xnor U787 (N_787,N_440,N_532);
nor U788 (N_788,N_556,N_508);
or U789 (N_789,N_463,N_469);
nor U790 (N_790,N_488,N_420);
xor U791 (N_791,N_509,N_486);
xor U792 (N_792,N_475,N_435);
or U793 (N_793,N_574,N_476);
nor U794 (N_794,N_557,N_551);
nand U795 (N_795,N_403,N_566);
or U796 (N_796,N_431,N_445);
nor U797 (N_797,N_463,N_567);
nand U798 (N_798,N_494,N_591);
or U799 (N_799,N_402,N_499);
nor U800 (N_800,N_727,N_784);
nor U801 (N_801,N_648,N_733);
nor U802 (N_802,N_712,N_684);
nor U803 (N_803,N_782,N_666);
and U804 (N_804,N_748,N_639);
nor U805 (N_805,N_798,N_640);
and U806 (N_806,N_627,N_645);
or U807 (N_807,N_797,N_749);
and U808 (N_808,N_769,N_722);
nand U809 (N_809,N_672,N_658);
and U810 (N_810,N_623,N_786);
nand U811 (N_811,N_759,N_783);
nor U812 (N_812,N_760,N_656);
nand U813 (N_813,N_650,N_767);
and U814 (N_814,N_775,N_789);
nor U815 (N_815,N_703,N_696);
and U816 (N_816,N_710,N_788);
and U817 (N_817,N_719,N_664);
or U818 (N_818,N_742,N_678);
and U819 (N_819,N_621,N_763);
and U820 (N_820,N_635,N_793);
or U821 (N_821,N_725,N_606);
or U822 (N_822,N_706,N_750);
nand U823 (N_823,N_714,N_785);
nor U824 (N_824,N_607,N_734);
and U825 (N_825,N_701,N_673);
or U826 (N_826,N_751,N_735);
nor U827 (N_827,N_756,N_729);
or U828 (N_828,N_713,N_632);
or U829 (N_829,N_795,N_711);
nor U830 (N_830,N_705,N_616);
nor U831 (N_831,N_700,N_668);
or U832 (N_832,N_772,N_693);
or U833 (N_833,N_610,N_644);
nor U834 (N_834,N_625,N_726);
nor U835 (N_835,N_665,N_694);
or U836 (N_836,N_773,N_758);
nor U837 (N_837,N_702,N_651);
nor U838 (N_838,N_614,N_660);
nand U839 (N_839,N_646,N_667);
nor U840 (N_840,N_780,N_659);
nand U841 (N_841,N_600,N_681);
or U842 (N_842,N_690,N_718);
nand U843 (N_843,N_686,N_695);
nor U844 (N_844,N_732,N_604);
nor U845 (N_845,N_754,N_674);
or U846 (N_846,N_708,N_762);
or U847 (N_847,N_791,N_716);
or U848 (N_848,N_634,N_728);
nor U849 (N_849,N_671,N_765);
and U850 (N_850,N_641,N_670);
or U851 (N_851,N_720,N_643);
or U852 (N_852,N_796,N_636);
nor U853 (N_853,N_685,N_655);
and U854 (N_854,N_740,N_611);
and U855 (N_855,N_717,N_633);
or U856 (N_856,N_778,N_608);
nor U857 (N_857,N_662,N_692);
nand U858 (N_858,N_624,N_637);
nor U859 (N_859,N_629,N_777);
or U860 (N_860,N_743,N_683);
and U861 (N_861,N_738,N_675);
and U862 (N_862,N_715,N_709);
and U863 (N_863,N_792,N_642);
nor U864 (N_864,N_746,N_697);
nand U865 (N_865,N_663,N_661);
nor U866 (N_866,N_790,N_618);
or U867 (N_867,N_745,N_669);
or U868 (N_868,N_619,N_761);
nand U869 (N_869,N_652,N_609);
or U870 (N_870,N_622,N_724);
nor U871 (N_871,N_603,N_620);
nand U872 (N_872,N_730,N_736);
nor U873 (N_873,N_677,N_723);
nor U874 (N_874,N_601,N_771);
or U875 (N_875,N_766,N_779);
nor U876 (N_876,N_764,N_794);
and U877 (N_877,N_747,N_770);
nand U878 (N_878,N_698,N_657);
nor U879 (N_879,N_688,N_752);
and U880 (N_880,N_768,N_757);
or U881 (N_881,N_731,N_741);
nor U882 (N_882,N_676,N_744);
nand U883 (N_883,N_753,N_707);
xor U884 (N_884,N_626,N_699);
or U885 (N_885,N_617,N_631);
nor U886 (N_886,N_653,N_613);
nand U887 (N_887,N_649,N_781);
and U888 (N_888,N_704,N_689);
nor U889 (N_889,N_630,N_799);
and U890 (N_890,N_612,N_739);
nand U891 (N_891,N_682,N_787);
or U892 (N_892,N_755,N_654);
xor U893 (N_893,N_605,N_774);
and U894 (N_894,N_680,N_776);
nand U895 (N_895,N_687,N_615);
or U896 (N_896,N_602,N_628);
xor U897 (N_897,N_737,N_679);
nand U898 (N_898,N_647,N_691);
nand U899 (N_899,N_721,N_638);
nand U900 (N_900,N_639,N_739);
nand U901 (N_901,N_752,N_613);
nand U902 (N_902,N_683,N_771);
nor U903 (N_903,N_677,N_786);
nor U904 (N_904,N_747,N_705);
nand U905 (N_905,N_632,N_658);
or U906 (N_906,N_651,N_733);
nand U907 (N_907,N_607,N_633);
or U908 (N_908,N_785,N_710);
and U909 (N_909,N_755,N_700);
nand U910 (N_910,N_776,N_643);
and U911 (N_911,N_675,N_671);
or U912 (N_912,N_749,N_603);
nor U913 (N_913,N_611,N_638);
nor U914 (N_914,N_747,N_777);
and U915 (N_915,N_692,N_618);
nor U916 (N_916,N_697,N_715);
nand U917 (N_917,N_766,N_791);
nor U918 (N_918,N_680,N_613);
nor U919 (N_919,N_781,N_684);
nand U920 (N_920,N_774,N_713);
and U921 (N_921,N_671,N_677);
xor U922 (N_922,N_682,N_742);
and U923 (N_923,N_605,N_733);
nand U924 (N_924,N_692,N_654);
nor U925 (N_925,N_717,N_789);
and U926 (N_926,N_798,N_644);
or U927 (N_927,N_653,N_636);
or U928 (N_928,N_776,N_701);
nand U929 (N_929,N_666,N_718);
nand U930 (N_930,N_698,N_682);
nor U931 (N_931,N_786,N_761);
and U932 (N_932,N_781,N_692);
nor U933 (N_933,N_655,N_720);
nor U934 (N_934,N_728,N_646);
and U935 (N_935,N_711,N_720);
nand U936 (N_936,N_711,N_745);
nand U937 (N_937,N_775,N_691);
and U938 (N_938,N_680,N_634);
and U939 (N_939,N_613,N_608);
and U940 (N_940,N_602,N_754);
or U941 (N_941,N_685,N_728);
nor U942 (N_942,N_688,N_679);
nand U943 (N_943,N_677,N_736);
and U944 (N_944,N_726,N_712);
or U945 (N_945,N_729,N_671);
nand U946 (N_946,N_701,N_683);
and U947 (N_947,N_775,N_694);
nand U948 (N_948,N_723,N_630);
and U949 (N_949,N_650,N_636);
and U950 (N_950,N_642,N_679);
nand U951 (N_951,N_750,N_683);
and U952 (N_952,N_651,N_620);
nand U953 (N_953,N_782,N_667);
or U954 (N_954,N_645,N_605);
nand U955 (N_955,N_731,N_761);
nand U956 (N_956,N_660,N_691);
nand U957 (N_957,N_778,N_626);
nor U958 (N_958,N_792,N_761);
nor U959 (N_959,N_768,N_637);
nand U960 (N_960,N_692,N_748);
nor U961 (N_961,N_683,N_657);
nor U962 (N_962,N_684,N_707);
nor U963 (N_963,N_761,N_610);
or U964 (N_964,N_758,N_717);
nand U965 (N_965,N_772,N_776);
and U966 (N_966,N_713,N_660);
nor U967 (N_967,N_676,N_731);
or U968 (N_968,N_745,N_761);
or U969 (N_969,N_652,N_773);
or U970 (N_970,N_767,N_759);
or U971 (N_971,N_660,N_647);
nand U972 (N_972,N_668,N_673);
or U973 (N_973,N_745,N_616);
and U974 (N_974,N_658,N_693);
nand U975 (N_975,N_705,N_666);
and U976 (N_976,N_719,N_661);
nand U977 (N_977,N_782,N_784);
nand U978 (N_978,N_736,N_789);
nand U979 (N_979,N_660,N_612);
nor U980 (N_980,N_607,N_646);
or U981 (N_981,N_674,N_755);
and U982 (N_982,N_602,N_601);
or U983 (N_983,N_720,N_736);
nor U984 (N_984,N_722,N_714);
and U985 (N_985,N_765,N_709);
and U986 (N_986,N_651,N_716);
nor U987 (N_987,N_659,N_608);
nor U988 (N_988,N_639,N_624);
and U989 (N_989,N_782,N_696);
nor U990 (N_990,N_671,N_790);
nand U991 (N_991,N_774,N_775);
nor U992 (N_992,N_659,N_698);
and U993 (N_993,N_653,N_614);
or U994 (N_994,N_711,N_794);
nor U995 (N_995,N_741,N_693);
and U996 (N_996,N_778,N_611);
or U997 (N_997,N_653,N_718);
nand U998 (N_998,N_731,N_627);
nand U999 (N_999,N_626,N_743);
or U1000 (N_1000,N_857,N_855);
or U1001 (N_1001,N_968,N_838);
nor U1002 (N_1002,N_813,N_890);
and U1003 (N_1003,N_920,N_905);
or U1004 (N_1004,N_891,N_930);
nor U1005 (N_1005,N_990,N_875);
or U1006 (N_1006,N_965,N_814);
and U1007 (N_1007,N_841,N_966);
nor U1008 (N_1008,N_877,N_852);
nor U1009 (N_1009,N_975,N_961);
or U1010 (N_1010,N_911,N_839);
nand U1011 (N_1011,N_835,N_806);
or U1012 (N_1012,N_886,N_873);
nand U1013 (N_1013,N_866,N_989);
and U1014 (N_1014,N_820,N_952);
nor U1015 (N_1015,N_812,N_900);
nor U1016 (N_1016,N_956,N_963);
nor U1017 (N_1017,N_982,N_861);
xor U1018 (N_1018,N_889,N_985);
and U1019 (N_1019,N_954,N_816);
or U1020 (N_1020,N_818,N_808);
nand U1021 (N_1021,N_996,N_910);
or U1022 (N_1022,N_896,N_976);
or U1023 (N_1023,N_827,N_869);
and U1024 (N_1024,N_822,N_942);
nor U1025 (N_1025,N_874,N_870);
xor U1026 (N_1026,N_811,N_955);
nor U1027 (N_1027,N_845,N_935);
nand U1028 (N_1028,N_937,N_871);
nand U1029 (N_1029,N_946,N_971);
and U1030 (N_1030,N_885,N_936);
nand U1031 (N_1031,N_926,N_803);
nand U1032 (N_1032,N_899,N_940);
nor U1033 (N_1033,N_846,N_938);
or U1034 (N_1034,N_804,N_919);
and U1035 (N_1035,N_817,N_878);
nand U1036 (N_1036,N_842,N_922);
nand U1037 (N_1037,N_957,N_932);
nand U1038 (N_1038,N_950,N_978);
nor U1039 (N_1039,N_906,N_964);
or U1040 (N_1040,N_892,N_948);
nand U1041 (N_1041,N_974,N_831);
or U1042 (N_1042,N_988,N_981);
and U1043 (N_1043,N_918,N_863);
nand U1044 (N_1044,N_879,N_883);
or U1045 (N_1045,N_925,N_972);
nor U1046 (N_1046,N_980,N_898);
or U1047 (N_1047,N_909,N_805);
or U1048 (N_1048,N_800,N_984);
and U1049 (N_1049,N_833,N_903);
or U1050 (N_1050,N_843,N_872);
nand U1051 (N_1051,N_902,N_832);
or U1052 (N_1052,N_801,N_823);
nor U1053 (N_1053,N_858,N_962);
or U1054 (N_1054,N_904,N_921);
nand U1055 (N_1055,N_880,N_848);
or U1056 (N_1056,N_850,N_840);
and U1057 (N_1057,N_959,N_928);
nand U1058 (N_1058,N_970,N_829);
nor U1059 (N_1059,N_893,N_998);
and U1060 (N_1060,N_924,N_836);
or U1061 (N_1061,N_809,N_815);
nor U1062 (N_1062,N_994,N_826);
and U1063 (N_1063,N_897,N_923);
and U1064 (N_1064,N_868,N_951);
or U1065 (N_1065,N_933,N_912);
nor U1066 (N_1066,N_810,N_882);
and U1067 (N_1067,N_825,N_943);
nor U1068 (N_1068,N_819,N_802);
or U1069 (N_1069,N_945,N_979);
or U1070 (N_1070,N_837,N_851);
and U1071 (N_1071,N_939,N_987);
nand U1072 (N_1072,N_949,N_941);
and U1073 (N_1073,N_999,N_867);
nor U1074 (N_1074,N_960,N_847);
and U1075 (N_1075,N_824,N_934);
xor U1076 (N_1076,N_888,N_807);
or U1077 (N_1077,N_864,N_953);
nand U1078 (N_1078,N_929,N_876);
or U1079 (N_1079,N_916,N_881);
nand U1080 (N_1080,N_862,N_995);
nor U1081 (N_1081,N_856,N_853);
or U1082 (N_1082,N_967,N_973);
nor U1083 (N_1083,N_977,N_887);
or U1084 (N_1084,N_849,N_884);
or U1085 (N_1085,N_997,N_907);
nor U1086 (N_1086,N_913,N_860);
nand U1087 (N_1087,N_914,N_944);
and U1088 (N_1088,N_901,N_992);
or U1089 (N_1089,N_983,N_927);
nor U1090 (N_1090,N_986,N_894);
or U1091 (N_1091,N_908,N_895);
and U1092 (N_1092,N_834,N_947);
nor U1093 (N_1093,N_859,N_917);
or U1094 (N_1094,N_821,N_991);
nor U1095 (N_1095,N_830,N_828);
or U1096 (N_1096,N_844,N_854);
and U1097 (N_1097,N_993,N_958);
nand U1098 (N_1098,N_915,N_969);
or U1099 (N_1099,N_865,N_931);
nand U1100 (N_1100,N_892,N_888);
nand U1101 (N_1101,N_856,N_994);
and U1102 (N_1102,N_892,N_990);
nor U1103 (N_1103,N_967,N_858);
nor U1104 (N_1104,N_810,N_946);
and U1105 (N_1105,N_866,N_962);
nor U1106 (N_1106,N_963,N_925);
nor U1107 (N_1107,N_972,N_850);
nor U1108 (N_1108,N_806,N_931);
and U1109 (N_1109,N_976,N_964);
nand U1110 (N_1110,N_870,N_926);
nor U1111 (N_1111,N_848,N_855);
or U1112 (N_1112,N_983,N_899);
and U1113 (N_1113,N_976,N_907);
or U1114 (N_1114,N_820,N_832);
nand U1115 (N_1115,N_920,N_917);
and U1116 (N_1116,N_914,N_993);
or U1117 (N_1117,N_838,N_820);
or U1118 (N_1118,N_863,N_844);
or U1119 (N_1119,N_889,N_960);
xnor U1120 (N_1120,N_992,N_991);
nand U1121 (N_1121,N_905,N_907);
and U1122 (N_1122,N_889,N_880);
nand U1123 (N_1123,N_845,N_873);
nor U1124 (N_1124,N_993,N_935);
and U1125 (N_1125,N_823,N_811);
nand U1126 (N_1126,N_955,N_999);
nand U1127 (N_1127,N_967,N_952);
nor U1128 (N_1128,N_878,N_994);
and U1129 (N_1129,N_963,N_993);
nand U1130 (N_1130,N_833,N_870);
xnor U1131 (N_1131,N_966,N_864);
nand U1132 (N_1132,N_872,N_927);
nor U1133 (N_1133,N_809,N_960);
and U1134 (N_1134,N_876,N_990);
nand U1135 (N_1135,N_800,N_856);
nand U1136 (N_1136,N_803,N_904);
and U1137 (N_1137,N_907,N_849);
or U1138 (N_1138,N_942,N_981);
or U1139 (N_1139,N_804,N_883);
nor U1140 (N_1140,N_837,N_938);
nand U1141 (N_1141,N_953,N_926);
or U1142 (N_1142,N_904,N_909);
and U1143 (N_1143,N_901,N_812);
and U1144 (N_1144,N_827,N_985);
nand U1145 (N_1145,N_866,N_862);
and U1146 (N_1146,N_808,N_932);
nor U1147 (N_1147,N_853,N_999);
or U1148 (N_1148,N_894,N_989);
xnor U1149 (N_1149,N_875,N_833);
or U1150 (N_1150,N_886,N_961);
and U1151 (N_1151,N_941,N_972);
and U1152 (N_1152,N_999,N_872);
nand U1153 (N_1153,N_827,N_978);
nor U1154 (N_1154,N_923,N_943);
nand U1155 (N_1155,N_932,N_948);
nand U1156 (N_1156,N_929,N_955);
and U1157 (N_1157,N_952,N_992);
or U1158 (N_1158,N_904,N_940);
nor U1159 (N_1159,N_917,N_882);
or U1160 (N_1160,N_801,N_861);
and U1161 (N_1161,N_903,N_955);
and U1162 (N_1162,N_934,N_914);
nor U1163 (N_1163,N_923,N_947);
and U1164 (N_1164,N_947,N_901);
and U1165 (N_1165,N_952,N_996);
nor U1166 (N_1166,N_811,N_849);
nand U1167 (N_1167,N_880,N_827);
nor U1168 (N_1168,N_972,N_960);
and U1169 (N_1169,N_813,N_878);
and U1170 (N_1170,N_958,N_876);
nor U1171 (N_1171,N_914,N_857);
or U1172 (N_1172,N_958,N_957);
nand U1173 (N_1173,N_888,N_917);
nand U1174 (N_1174,N_887,N_916);
nand U1175 (N_1175,N_983,N_905);
nand U1176 (N_1176,N_960,N_859);
and U1177 (N_1177,N_857,N_991);
or U1178 (N_1178,N_926,N_971);
nand U1179 (N_1179,N_813,N_833);
nand U1180 (N_1180,N_975,N_901);
nand U1181 (N_1181,N_803,N_884);
or U1182 (N_1182,N_836,N_961);
or U1183 (N_1183,N_937,N_900);
or U1184 (N_1184,N_875,N_870);
nand U1185 (N_1185,N_811,N_885);
or U1186 (N_1186,N_923,N_967);
nand U1187 (N_1187,N_911,N_915);
and U1188 (N_1188,N_857,N_910);
or U1189 (N_1189,N_864,N_929);
and U1190 (N_1190,N_924,N_865);
nand U1191 (N_1191,N_807,N_829);
and U1192 (N_1192,N_977,N_910);
or U1193 (N_1193,N_837,N_985);
and U1194 (N_1194,N_895,N_998);
nor U1195 (N_1195,N_896,N_993);
and U1196 (N_1196,N_852,N_873);
nor U1197 (N_1197,N_904,N_925);
nor U1198 (N_1198,N_871,N_917);
nand U1199 (N_1199,N_898,N_955);
or U1200 (N_1200,N_1185,N_1182);
nor U1201 (N_1201,N_1179,N_1136);
or U1202 (N_1202,N_1156,N_1036);
and U1203 (N_1203,N_1132,N_1034);
nand U1204 (N_1204,N_1039,N_1121);
and U1205 (N_1205,N_1157,N_1052);
and U1206 (N_1206,N_1014,N_1099);
or U1207 (N_1207,N_1002,N_1012);
or U1208 (N_1208,N_1146,N_1147);
nand U1209 (N_1209,N_1126,N_1024);
or U1210 (N_1210,N_1118,N_1045);
or U1211 (N_1211,N_1074,N_1088);
nand U1212 (N_1212,N_1163,N_1107);
nor U1213 (N_1213,N_1153,N_1116);
nand U1214 (N_1214,N_1187,N_1075);
and U1215 (N_1215,N_1098,N_1047);
or U1216 (N_1216,N_1007,N_1000);
nand U1217 (N_1217,N_1040,N_1051);
and U1218 (N_1218,N_1095,N_1104);
nand U1219 (N_1219,N_1139,N_1180);
nand U1220 (N_1220,N_1111,N_1066);
or U1221 (N_1221,N_1031,N_1169);
nor U1222 (N_1222,N_1117,N_1113);
and U1223 (N_1223,N_1044,N_1164);
nand U1224 (N_1224,N_1033,N_1019);
xnor U1225 (N_1225,N_1127,N_1166);
and U1226 (N_1226,N_1178,N_1076);
or U1227 (N_1227,N_1027,N_1142);
and U1228 (N_1228,N_1056,N_1125);
nand U1229 (N_1229,N_1080,N_1188);
or U1230 (N_1230,N_1137,N_1120);
or U1231 (N_1231,N_1108,N_1124);
and U1232 (N_1232,N_1050,N_1170);
nor U1233 (N_1233,N_1054,N_1195);
or U1234 (N_1234,N_1059,N_1109);
or U1235 (N_1235,N_1097,N_1068);
nor U1236 (N_1236,N_1023,N_1143);
or U1237 (N_1237,N_1029,N_1155);
xnor U1238 (N_1238,N_1003,N_1189);
or U1239 (N_1239,N_1140,N_1094);
or U1240 (N_1240,N_1082,N_1055);
and U1241 (N_1241,N_1165,N_1061);
or U1242 (N_1242,N_1130,N_1010);
and U1243 (N_1243,N_1148,N_1158);
or U1244 (N_1244,N_1176,N_1053);
or U1245 (N_1245,N_1115,N_1042);
nand U1246 (N_1246,N_1102,N_1199);
nand U1247 (N_1247,N_1114,N_1135);
and U1248 (N_1248,N_1167,N_1192);
nor U1249 (N_1249,N_1020,N_1028);
nand U1250 (N_1250,N_1183,N_1089);
nand U1251 (N_1251,N_1069,N_1101);
nor U1252 (N_1252,N_1058,N_1175);
nor U1253 (N_1253,N_1022,N_1048);
and U1254 (N_1254,N_1090,N_1122);
nor U1255 (N_1255,N_1057,N_1083);
nor U1256 (N_1256,N_1173,N_1103);
or U1257 (N_1257,N_1065,N_1017);
or U1258 (N_1258,N_1062,N_1144);
and U1259 (N_1259,N_1123,N_1145);
or U1260 (N_1260,N_1138,N_1006);
and U1261 (N_1261,N_1073,N_1043);
nand U1262 (N_1262,N_1193,N_1079);
nand U1263 (N_1263,N_1149,N_1141);
nor U1264 (N_1264,N_1096,N_1021);
or U1265 (N_1265,N_1004,N_1035);
or U1266 (N_1266,N_1106,N_1060);
or U1267 (N_1267,N_1197,N_1009);
nor U1268 (N_1268,N_1011,N_1131);
and U1269 (N_1269,N_1190,N_1133);
nand U1270 (N_1270,N_1150,N_1085);
and U1271 (N_1271,N_1008,N_1161);
and U1272 (N_1272,N_1037,N_1159);
nor U1273 (N_1273,N_1026,N_1078);
or U1274 (N_1274,N_1100,N_1071);
or U1275 (N_1275,N_1032,N_1086);
and U1276 (N_1276,N_1198,N_1105);
or U1277 (N_1277,N_1018,N_1063);
and U1278 (N_1278,N_1194,N_1001);
nor U1279 (N_1279,N_1191,N_1110);
nand U1280 (N_1280,N_1046,N_1013);
and U1281 (N_1281,N_1072,N_1015);
nor U1282 (N_1282,N_1152,N_1041);
nand U1283 (N_1283,N_1174,N_1092);
nor U1284 (N_1284,N_1064,N_1160);
and U1285 (N_1285,N_1162,N_1067);
nand U1286 (N_1286,N_1172,N_1168);
or U1287 (N_1287,N_1091,N_1049);
or U1288 (N_1288,N_1077,N_1016);
nand U1289 (N_1289,N_1184,N_1171);
or U1290 (N_1290,N_1087,N_1030);
nand U1291 (N_1291,N_1070,N_1093);
or U1292 (N_1292,N_1081,N_1154);
nor U1293 (N_1293,N_1038,N_1177);
nand U1294 (N_1294,N_1181,N_1196);
and U1295 (N_1295,N_1025,N_1112);
or U1296 (N_1296,N_1084,N_1128);
or U1297 (N_1297,N_1129,N_1119);
nor U1298 (N_1298,N_1151,N_1005);
nor U1299 (N_1299,N_1134,N_1186);
and U1300 (N_1300,N_1089,N_1060);
nor U1301 (N_1301,N_1176,N_1119);
and U1302 (N_1302,N_1000,N_1187);
nor U1303 (N_1303,N_1118,N_1016);
and U1304 (N_1304,N_1109,N_1100);
nor U1305 (N_1305,N_1081,N_1086);
or U1306 (N_1306,N_1046,N_1091);
or U1307 (N_1307,N_1148,N_1081);
nand U1308 (N_1308,N_1043,N_1048);
nor U1309 (N_1309,N_1022,N_1113);
and U1310 (N_1310,N_1119,N_1158);
or U1311 (N_1311,N_1022,N_1149);
and U1312 (N_1312,N_1012,N_1004);
or U1313 (N_1313,N_1192,N_1067);
nand U1314 (N_1314,N_1071,N_1137);
or U1315 (N_1315,N_1135,N_1019);
and U1316 (N_1316,N_1039,N_1161);
or U1317 (N_1317,N_1048,N_1109);
nor U1318 (N_1318,N_1166,N_1002);
or U1319 (N_1319,N_1072,N_1029);
nor U1320 (N_1320,N_1024,N_1150);
nor U1321 (N_1321,N_1009,N_1097);
and U1322 (N_1322,N_1061,N_1103);
and U1323 (N_1323,N_1020,N_1149);
nand U1324 (N_1324,N_1158,N_1187);
nor U1325 (N_1325,N_1098,N_1054);
or U1326 (N_1326,N_1016,N_1161);
nand U1327 (N_1327,N_1113,N_1126);
and U1328 (N_1328,N_1104,N_1050);
and U1329 (N_1329,N_1002,N_1058);
or U1330 (N_1330,N_1026,N_1140);
nand U1331 (N_1331,N_1114,N_1195);
and U1332 (N_1332,N_1122,N_1169);
or U1333 (N_1333,N_1167,N_1139);
and U1334 (N_1334,N_1133,N_1131);
and U1335 (N_1335,N_1082,N_1018);
or U1336 (N_1336,N_1132,N_1108);
xor U1337 (N_1337,N_1086,N_1056);
or U1338 (N_1338,N_1019,N_1175);
or U1339 (N_1339,N_1051,N_1042);
nand U1340 (N_1340,N_1106,N_1085);
and U1341 (N_1341,N_1106,N_1022);
nor U1342 (N_1342,N_1126,N_1135);
and U1343 (N_1343,N_1075,N_1101);
nor U1344 (N_1344,N_1042,N_1009);
nand U1345 (N_1345,N_1033,N_1083);
and U1346 (N_1346,N_1004,N_1107);
or U1347 (N_1347,N_1056,N_1023);
and U1348 (N_1348,N_1125,N_1075);
nor U1349 (N_1349,N_1004,N_1124);
or U1350 (N_1350,N_1039,N_1177);
and U1351 (N_1351,N_1000,N_1164);
nor U1352 (N_1352,N_1176,N_1166);
nand U1353 (N_1353,N_1011,N_1054);
nand U1354 (N_1354,N_1124,N_1128);
nand U1355 (N_1355,N_1101,N_1134);
and U1356 (N_1356,N_1000,N_1190);
xnor U1357 (N_1357,N_1165,N_1059);
and U1358 (N_1358,N_1154,N_1100);
or U1359 (N_1359,N_1173,N_1049);
and U1360 (N_1360,N_1112,N_1178);
or U1361 (N_1361,N_1182,N_1003);
or U1362 (N_1362,N_1079,N_1113);
nor U1363 (N_1363,N_1033,N_1097);
nand U1364 (N_1364,N_1031,N_1188);
or U1365 (N_1365,N_1150,N_1140);
or U1366 (N_1366,N_1103,N_1123);
or U1367 (N_1367,N_1154,N_1017);
nor U1368 (N_1368,N_1102,N_1067);
and U1369 (N_1369,N_1009,N_1117);
nor U1370 (N_1370,N_1198,N_1172);
nand U1371 (N_1371,N_1014,N_1138);
nor U1372 (N_1372,N_1184,N_1168);
or U1373 (N_1373,N_1166,N_1015);
nand U1374 (N_1374,N_1019,N_1049);
nand U1375 (N_1375,N_1081,N_1080);
and U1376 (N_1376,N_1057,N_1104);
nor U1377 (N_1377,N_1016,N_1050);
and U1378 (N_1378,N_1055,N_1100);
and U1379 (N_1379,N_1091,N_1084);
nor U1380 (N_1380,N_1009,N_1189);
nor U1381 (N_1381,N_1173,N_1071);
or U1382 (N_1382,N_1123,N_1187);
xor U1383 (N_1383,N_1035,N_1006);
and U1384 (N_1384,N_1020,N_1108);
nand U1385 (N_1385,N_1034,N_1140);
or U1386 (N_1386,N_1008,N_1170);
nor U1387 (N_1387,N_1013,N_1145);
nand U1388 (N_1388,N_1071,N_1183);
nand U1389 (N_1389,N_1167,N_1187);
and U1390 (N_1390,N_1091,N_1035);
nor U1391 (N_1391,N_1063,N_1131);
or U1392 (N_1392,N_1176,N_1175);
nand U1393 (N_1393,N_1031,N_1039);
or U1394 (N_1394,N_1179,N_1072);
and U1395 (N_1395,N_1111,N_1083);
nor U1396 (N_1396,N_1108,N_1025);
nor U1397 (N_1397,N_1023,N_1197);
or U1398 (N_1398,N_1131,N_1042);
or U1399 (N_1399,N_1135,N_1171);
or U1400 (N_1400,N_1361,N_1328);
nor U1401 (N_1401,N_1261,N_1365);
or U1402 (N_1402,N_1335,N_1256);
nand U1403 (N_1403,N_1314,N_1205);
or U1404 (N_1404,N_1350,N_1315);
nand U1405 (N_1405,N_1376,N_1390);
nand U1406 (N_1406,N_1282,N_1285);
xnor U1407 (N_1407,N_1312,N_1207);
nor U1408 (N_1408,N_1373,N_1331);
nand U1409 (N_1409,N_1351,N_1334);
nand U1410 (N_1410,N_1341,N_1380);
nand U1411 (N_1411,N_1228,N_1306);
or U1412 (N_1412,N_1379,N_1319);
nor U1413 (N_1413,N_1269,N_1291);
nor U1414 (N_1414,N_1245,N_1253);
nand U1415 (N_1415,N_1243,N_1333);
nor U1416 (N_1416,N_1302,N_1398);
nor U1417 (N_1417,N_1215,N_1294);
and U1418 (N_1418,N_1235,N_1286);
and U1419 (N_1419,N_1381,N_1384);
nor U1420 (N_1420,N_1227,N_1304);
or U1421 (N_1421,N_1206,N_1281);
nor U1422 (N_1422,N_1236,N_1326);
or U1423 (N_1423,N_1283,N_1208);
nor U1424 (N_1424,N_1318,N_1367);
and U1425 (N_1425,N_1284,N_1349);
nor U1426 (N_1426,N_1303,N_1378);
nand U1427 (N_1427,N_1389,N_1250);
nor U1428 (N_1428,N_1226,N_1219);
nand U1429 (N_1429,N_1336,N_1241);
xnor U1430 (N_1430,N_1358,N_1316);
or U1431 (N_1431,N_1385,N_1259);
or U1432 (N_1432,N_1289,N_1295);
nor U1433 (N_1433,N_1340,N_1338);
nand U1434 (N_1434,N_1260,N_1290);
or U1435 (N_1435,N_1267,N_1355);
and U1436 (N_1436,N_1305,N_1268);
and U1437 (N_1437,N_1357,N_1313);
nand U1438 (N_1438,N_1265,N_1272);
nand U1439 (N_1439,N_1214,N_1363);
or U1440 (N_1440,N_1242,N_1320);
or U1441 (N_1441,N_1274,N_1388);
nor U1442 (N_1442,N_1292,N_1310);
nor U1443 (N_1443,N_1202,N_1298);
nand U1444 (N_1444,N_1270,N_1240);
nor U1445 (N_1445,N_1217,N_1383);
nand U1446 (N_1446,N_1393,N_1354);
and U1447 (N_1447,N_1273,N_1308);
nand U1448 (N_1448,N_1264,N_1399);
nand U1449 (N_1449,N_1266,N_1279);
and U1450 (N_1450,N_1211,N_1307);
nand U1451 (N_1451,N_1251,N_1257);
or U1452 (N_1452,N_1329,N_1311);
or U1453 (N_1453,N_1330,N_1271);
nor U1454 (N_1454,N_1247,N_1222);
nor U1455 (N_1455,N_1321,N_1233);
or U1456 (N_1456,N_1299,N_1345);
nand U1457 (N_1457,N_1263,N_1386);
or U1458 (N_1458,N_1201,N_1394);
and U1459 (N_1459,N_1344,N_1374);
or U1460 (N_1460,N_1397,N_1325);
and U1461 (N_1461,N_1348,N_1218);
nor U1462 (N_1462,N_1209,N_1237);
nor U1463 (N_1463,N_1287,N_1342);
nor U1464 (N_1464,N_1293,N_1301);
nor U1465 (N_1465,N_1232,N_1352);
nor U1466 (N_1466,N_1370,N_1221);
or U1467 (N_1467,N_1223,N_1346);
and U1468 (N_1468,N_1368,N_1216);
and U1469 (N_1469,N_1224,N_1396);
nand U1470 (N_1470,N_1220,N_1258);
nand U1471 (N_1471,N_1255,N_1392);
and U1472 (N_1472,N_1332,N_1353);
nor U1473 (N_1473,N_1364,N_1337);
and U1474 (N_1474,N_1244,N_1248);
nand U1475 (N_1475,N_1296,N_1347);
or U1476 (N_1476,N_1317,N_1377);
or U1477 (N_1477,N_1297,N_1323);
nand U1478 (N_1478,N_1200,N_1339);
and U1479 (N_1479,N_1366,N_1210);
nand U1480 (N_1480,N_1262,N_1371);
or U1481 (N_1481,N_1372,N_1234);
or U1482 (N_1482,N_1212,N_1277);
and U1483 (N_1483,N_1288,N_1322);
nor U1484 (N_1484,N_1275,N_1387);
and U1485 (N_1485,N_1375,N_1382);
nand U1486 (N_1486,N_1249,N_1391);
nand U1487 (N_1487,N_1276,N_1225);
nor U1488 (N_1488,N_1213,N_1300);
nand U1489 (N_1489,N_1369,N_1343);
nor U1490 (N_1490,N_1327,N_1362);
and U1491 (N_1491,N_1324,N_1229);
and U1492 (N_1492,N_1395,N_1238);
nor U1493 (N_1493,N_1252,N_1359);
and U1494 (N_1494,N_1239,N_1230);
nand U1495 (N_1495,N_1278,N_1246);
nor U1496 (N_1496,N_1360,N_1309);
nand U1497 (N_1497,N_1204,N_1280);
or U1498 (N_1498,N_1231,N_1356);
and U1499 (N_1499,N_1254,N_1203);
nor U1500 (N_1500,N_1335,N_1277);
nor U1501 (N_1501,N_1310,N_1315);
and U1502 (N_1502,N_1373,N_1369);
or U1503 (N_1503,N_1208,N_1380);
and U1504 (N_1504,N_1294,N_1254);
and U1505 (N_1505,N_1391,N_1216);
and U1506 (N_1506,N_1224,N_1377);
nor U1507 (N_1507,N_1353,N_1330);
nor U1508 (N_1508,N_1345,N_1312);
or U1509 (N_1509,N_1313,N_1237);
or U1510 (N_1510,N_1383,N_1338);
nor U1511 (N_1511,N_1332,N_1290);
and U1512 (N_1512,N_1291,N_1315);
nand U1513 (N_1513,N_1205,N_1231);
nand U1514 (N_1514,N_1307,N_1279);
nand U1515 (N_1515,N_1200,N_1353);
and U1516 (N_1516,N_1242,N_1300);
and U1517 (N_1517,N_1226,N_1383);
nor U1518 (N_1518,N_1256,N_1207);
or U1519 (N_1519,N_1241,N_1240);
nor U1520 (N_1520,N_1311,N_1327);
nor U1521 (N_1521,N_1262,N_1370);
nor U1522 (N_1522,N_1325,N_1385);
nor U1523 (N_1523,N_1282,N_1204);
nand U1524 (N_1524,N_1341,N_1212);
or U1525 (N_1525,N_1271,N_1254);
nand U1526 (N_1526,N_1240,N_1389);
and U1527 (N_1527,N_1277,N_1223);
nand U1528 (N_1528,N_1263,N_1380);
and U1529 (N_1529,N_1294,N_1289);
nand U1530 (N_1530,N_1303,N_1308);
nand U1531 (N_1531,N_1289,N_1263);
nor U1532 (N_1532,N_1207,N_1224);
nor U1533 (N_1533,N_1372,N_1256);
or U1534 (N_1534,N_1241,N_1320);
nand U1535 (N_1535,N_1377,N_1311);
nand U1536 (N_1536,N_1200,N_1304);
nor U1537 (N_1537,N_1344,N_1339);
nand U1538 (N_1538,N_1382,N_1215);
nor U1539 (N_1539,N_1240,N_1352);
nand U1540 (N_1540,N_1355,N_1259);
or U1541 (N_1541,N_1254,N_1323);
nor U1542 (N_1542,N_1272,N_1211);
or U1543 (N_1543,N_1312,N_1318);
nor U1544 (N_1544,N_1304,N_1273);
nand U1545 (N_1545,N_1270,N_1313);
xor U1546 (N_1546,N_1351,N_1332);
or U1547 (N_1547,N_1249,N_1248);
nor U1548 (N_1548,N_1369,N_1376);
nand U1549 (N_1549,N_1354,N_1377);
nor U1550 (N_1550,N_1246,N_1301);
and U1551 (N_1551,N_1398,N_1211);
and U1552 (N_1552,N_1360,N_1253);
or U1553 (N_1553,N_1238,N_1320);
nand U1554 (N_1554,N_1243,N_1336);
or U1555 (N_1555,N_1285,N_1243);
and U1556 (N_1556,N_1249,N_1244);
or U1557 (N_1557,N_1306,N_1394);
and U1558 (N_1558,N_1203,N_1265);
nand U1559 (N_1559,N_1390,N_1207);
nand U1560 (N_1560,N_1350,N_1320);
nor U1561 (N_1561,N_1355,N_1247);
nor U1562 (N_1562,N_1271,N_1284);
xor U1563 (N_1563,N_1361,N_1334);
nand U1564 (N_1564,N_1362,N_1257);
nor U1565 (N_1565,N_1205,N_1375);
nand U1566 (N_1566,N_1341,N_1247);
nand U1567 (N_1567,N_1308,N_1267);
and U1568 (N_1568,N_1250,N_1302);
nand U1569 (N_1569,N_1395,N_1279);
and U1570 (N_1570,N_1292,N_1346);
or U1571 (N_1571,N_1278,N_1300);
and U1572 (N_1572,N_1275,N_1356);
and U1573 (N_1573,N_1339,N_1274);
and U1574 (N_1574,N_1227,N_1231);
and U1575 (N_1575,N_1244,N_1231);
or U1576 (N_1576,N_1293,N_1299);
and U1577 (N_1577,N_1241,N_1281);
nor U1578 (N_1578,N_1279,N_1289);
nor U1579 (N_1579,N_1218,N_1294);
and U1580 (N_1580,N_1381,N_1240);
or U1581 (N_1581,N_1260,N_1215);
or U1582 (N_1582,N_1224,N_1286);
and U1583 (N_1583,N_1346,N_1270);
nor U1584 (N_1584,N_1335,N_1239);
nor U1585 (N_1585,N_1326,N_1208);
nand U1586 (N_1586,N_1380,N_1201);
nor U1587 (N_1587,N_1268,N_1201);
and U1588 (N_1588,N_1364,N_1247);
xnor U1589 (N_1589,N_1248,N_1345);
nand U1590 (N_1590,N_1399,N_1267);
nor U1591 (N_1591,N_1258,N_1237);
nand U1592 (N_1592,N_1235,N_1274);
nand U1593 (N_1593,N_1232,N_1392);
nand U1594 (N_1594,N_1209,N_1254);
or U1595 (N_1595,N_1322,N_1353);
nand U1596 (N_1596,N_1213,N_1254);
nand U1597 (N_1597,N_1399,N_1352);
and U1598 (N_1598,N_1252,N_1321);
nor U1599 (N_1599,N_1257,N_1363);
and U1600 (N_1600,N_1418,N_1462);
and U1601 (N_1601,N_1599,N_1555);
nand U1602 (N_1602,N_1492,N_1544);
nand U1603 (N_1603,N_1499,N_1406);
nor U1604 (N_1604,N_1509,N_1573);
or U1605 (N_1605,N_1505,N_1478);
nand U1606 (N_1606,N_1534,N_1421);
xnor U1607 (N_1607,N_1459,N_1480);
or U1608 (N_1608,N_1494,N_1550);
nand U1609 (N_1609,N_1542,N_1496);
nor U1610 (N_1610,N_1488,N_1476);
or U1611 (N_1611,N_1562,N_1556);
and U1612 (N_1612,N_1463,N_1551);
nor U1613 (N_1613,N_1595,N_1433);
nand U1614 (N_1614,N_1596,N_1412);
nor U1615 (N_1615,N_1422,N_1501);
or U1616 (N_1616,N_1519,N_1587);
nand U1617 (N_1617,N_1526,N_1580);
nand U1618 (N_1618,N_1558,N_1465);
nand U1619 (N_1619,N_1432,N_1436);
and U1620 (N_1620,N_1513,N_1517);
nor U1621 (N_1621,N_1424,N_1477);
nor U1622 (N_1622,N_1438,N_1518);
and U1623 (N_1623,N_1411,N_1549);
or U1624 (N_1624,N_1548,N_1557);
nand U1625 (N_1625,N_1510,N_1597);
and U1626 (N_1626,N_1554,N_1588);
or U1627 (N_1627,N_1401,N_1404);
or U1628 (N_1628,N_1407,N_1443);
and U1629 (N_1629,N_1442,N_1541);
nand U1630 (N_1630,N_1449,N_1524);
and U1631 (N_1631,N_1435,N_1583);
nor U1632 (N_1632,N_1520,N_1452);
nor U1633 (N_1633,N_1483,N_1482);
and U1634 (N_1634,N_1409,N_1437);
nand U1635 (N_1635,N_1473,N_1455);
or U1636 (N_1636,N_1460,N_1419);
nor U1637 (N_1637,N_1414,N_1582);
nand U1638 (N_1638,N_1594,N_1445);
nand U1639 (N_1639,N_1585,N_1527);
nor U1640 (N_1640,N_1589,N_1584);
and U1641 (N_1641,N_1467,N_1408);
or U1642 (N_1642,N_1538,N_1507);
nor U1643 (N_1643,N_1565,N_1486);
and U1644 (N_1644,N_1495,N_1561);
and U1645 (N_1645,N_1434,N_1586);
nand U1646 (N_1646,N_1572,N_1559);
nand U1647 (N_1647,N_1575,N_1456);
nand U1648 (N_1648,N_1498,N_1454);
or U1649 (N_1649,N_1515,N_1576);
nor U1650 (N_1650,N_1566,N_1571);
nand U1651 (N_1651,N_1487,N_1415);
nor U1652 (N_1652,N_1431,N_1423);
and U1653 (N_1653,N_1593,N_1536);
nor U1654 (N_1654,N_1491,N_1440);
or U1655 (N_1655,N_1451,N_1564);
or U1656 (N_1656,N_1441,N_1410);
and U1657 (N_1657,N_1540,N_1420);
nor U1658 (N_1658,N_1446,N_1522);
nand U1659 (N_1659,N_1416,N_1457);
nor U1660 (N_1660,N_1428,N_1592);
and U1661 (N_1661,N_1591,N_1444);
and U1662 (N_1662,N_1503,N_1511);
nor U1663 (N_1663,N_1490,N_1405);
nor U1664 (N_1664,N_1447,N_1532);
or U1665 (N_1665,N_1426,N_1523);
and U1666 (N_1666,N_1552,N_1506);
or U1667 (N_1667,N_1429,N_1461);
or U1668 (N_1668,N_1413,N_1474);
nand U1669 (N_1669,N_1504,N_1458);
nor U1670 (N_1670,N_1533,N_1514);
nand U1671 (N_1671,N_1535,N_1516);
or U1672 (N_1672,N_1563,N_1508);
and U1673 (N_1673,N_1469,N_1471);
nor U1674 (N_1674,N_1425,N_1590);
nand U1675 (N_1675,N_1485,N_1493);
and U1676 (N_1676,N_1484,N_1568);
nand U1677 (N_1677,N_1531,N_1574);
and U1678 (N_1678,N_1453,N_1430);
or U1679 (N_1679,N_1464,N_1466);
or U1680 (N_1680,N_1569,N_1577);
or U1681 (N_1681,N_1475,N_1545);
nor U1682 (N_1682,N_1479,N_1489);
nand U1683 (N_1683,N_1546,N_1560);
or U1684 (N_1684,N_1427,N_1439);
or U1685 (N_1685,N_1528,N_1525);
nand U1686 (N_1686,N_1500,N_1570);
and U1687 (N_1687,N_1529,N_1403);
nor U1688 (N_1688,N_1530,N_1481);
nand U1689 (N_1689,N_1581,N_1448);
and U1690 (N_1690,N_1567,N_1547);
or U1691 (N_1691,N_1579,N_1468);
and U1692 (N_1692,N_1539,N_1450);
or U1693 (N_1693,N_1417,N_1472);
nand U1694 (N_1694,N_1598,N_1400);
or U1695 (N_1695,N_1537,N_1497);
nor U1696 (N_1696,N_1470,N_1502);
or U1697 (N_1697,N_1543,N_1553);
nand U1698 (N_1698,N_1578,N_1521);
nor U1699 (N_1699,N_1402,N_1512);
or U1700 (N_1700,N_1433,N_1501);
or U1701 (N_1701,N_1481,N_1563);
or U1702 (N_1702,N_1507,N_1569);
nand U1703 (N_1703,N_1457,N_1536);
or U1704 (N_1704,N_1527,N_1430);
and U1705 (N_1705,N_1587,N_1575);
xnor U1706 (N_1706,N_1454,N_1543);
and U1707 (N_1707,N_1410,N_1547);
nor U1708 (N_1708,N_1436,N_1491);
and U1709 (N_1709,N_1496,N_1423);
and U1710 (N_1710,N_1511,N_1561);
nor U1711 (N_1711,N_1421,N_1545);
nand U1712 (N_1712,N_1567,N_1415);
and U1713 (N_1713,N_1501,N_1428);
or U1714 (N_1714,N_1483,N_1470);
nor U1715 (N_1715,N_1554,N_1549);
nand U1716 (N_1716,N_1498,N_1470);
or U1717 (N_1717,N_1415,N_1510);
and U1718 (N_1718,N_1583,N_1589);
nor U1719 (N_1719,N_1551,N_1584);
or U1720 (N_1720,N_1482,N_1466);
nand U1721 (N_1721,N_1484,N_1424);
nand U1722 (N_1722,N_1549,N_1562);
and U1723 (N_1723,N_1407,N_1427);
nand U1724 (N_1724,N_1478,N_1570);
nor U1725 (N_1725,N_1422,N_1406);
and U1726 (N_1726,N_1560,N_1538);
xor U1727 (N_1727,N_1558,N_1594);
and U1728 (N_1728,N_1486,N_1523);
or U1729 (N_1729,N_1550,N_1434);
nand U1730 (N_1730,N_1589,N_1597);
or U1731 (N_1731,N_1496,N_1526);
nor U1732 (N_1732,N_1555,N_1525);
nor U1733 (N_1733,N_1537,N_1534);
and U1734 (N_1734,N_1525,N_1548);
or U1735 (N_1735,N_1418,N_1425);
nor U1736 (N_1736,N_1406,N_1551);
nand U1737 (N_1737,N_1510,N_1520);
nor U1738 (N_1738,N_1479,N_1529);
nor U1739 (N_1739,N_1467,N_1435);
and U1740 (N_1740,N_1482,N_1420);
or U1741 (N_1741,N_1509,N_1448);
and U1742 (N_1742,N_1576,N_1591);
or U1743 (N_1743,N_1590,N_1539);
and U1744 (N_1744,N_1470,N_1422);
nor U1745 (N_1745,N_1427,N_1419);
nand U1746 (N_1746,N_1430,N_1461);
nand U1747 (N_1747,N_1433,N_1428);
nand U1748 (N_1748,N_1426,N_1535);
and U1749 (N_1749,N_1483,N_1403);
or U1750 (N_1750,N_1465,N_1431);
nor U1751 (N_1751,N_1423,N_1438);
and U1752 (N_1752,N_1402,N_1508);
xnor U1753 (N_1753,N_1449,N_1582);
or U1754 (N_1754,N_1544,N_1566);
nand U1755 (N_1755,N_1583,N_1514);
nor U1756 (N_1756,N_1460,N_1527);
nor U1757 (N_1757,N_1534,N_1550);
or U1758 (N_1758,N_1466,N_1545);
nor U1759 (N_1759,N_1561,N_1428);
or U1760 (N_1760,N_1447,N_1552);
and U1761 (N_1761,N_1526,N_1560);
nand U1762 (N_1762,N_1539,N_1477);
or U1763 (N_1763,N_1527,N_1537);
nor U1764 (N_1764,N_1411,N_1503);
and U1765 (N_1765,N_1576,N_1528);
or U1766 (N_1766,N_1597,N_1457);
or U1767 (N_1767,N_1532,N_1445);
nand U1768 (N_1768,N_1509,N_1535);
nor U1769 (N_1769,N_1472,N_1593);
and U1770 (N_1770,N_1423,N_1454);
or U1771 (N_1771,N_1530,N_1443);
and U1772 (N_1772,N_1503,N_1586);
nor U1773 (N_1773,N_1463,N_1421);
and U1774 (N_1774,N_1581,N_1589);
nor U1775 (N_1775,N_1424,N_1527);
and U1776 (N_1776,N_1438,N_1455);
and U1777 (N_1777,N_1466,N_1517);
or U1778 (N_1778,N_1561,N_1579);
and U1779 (N_1779,N_1422,N_1589);
or U1780 (N_1780,N_1557,N_1595);
and U1781 (N_1781,N_1520,N_1506);
and U1782 (N_1782,N_1525,N_1560);
and U1783 (N_1783,N_1591,N_1501);
nand U1784 (N_1784,N_1535,N_1504);
xnor U1785 (N_1785,N_1482,N_1578);
nand U1786 (N_1786,N_1542,N_1469);
nand U1787 (N_1787,N_1524,N_1530);
and U1788 (N_1788,N_1590,N_1586);
and U1789 (N_1789,N_1421,N_1589);
and U1790 (N_1790,N_1486,N_1481);
nand U1791 (N_1791,N_1542,N_1455);
and U1792 (N_1792,N_1533,N_1491);
and U1793 (N_1793,N_1458,N_1534);
nor U1794 (N_1794,N_1557,N_1512);
or U1795 (N_1795,N_1486,N_1436);
or U1796 (N_1796,N_1423,N_1537);
or U1797 (N_1797,N_1454,N_1438);
nor U1798 (N_1798,N_1435,N_1588);
nand U1799 (N_1799,N_1485,N_1541);
and U1800 (N_1800,N_1694,N_1740);
and U1801 (N_1801,N_1671,N_1749);
nor U1802 (N_1802,N_1797,N_1675);
and U1803 (N_1803,N_1759,N_1697);
and U1804 (N_1804,N_1779,N_1665);
nand U1805 (N_1805,N_1658,N_1656);
or U1806 (N_1806,N_1687,N_1704);
nand U1807 (N_1807,N_1647,N_1638);
nor U1808 (N_1808,N_1734,N_1708);
and U1809 (N_1809,N_1725,N_1622);
xor U1810 (N_1810,N_1631,N_1706);
and U1811 (N_1811,N_1718,N_1775);
or U1812 (N_1812,N_1777,N_1745);
nand U1813 (N_1813,N_1651,N_1765);
nor U1814 (N_1814,N_1771,N_1657);
or U1815 (N_1815,N_1690,N_1660);
nand U1816 (N_1816,N_1785,N_1732);
and U1817 (N_1817,N_1667,N_1663);
nor U1818 (N_1818,N_1637,N_1644);
and U1819 (N_1819,N_1630,N_1608);
nor U1820 (N_1820,N_1791,N_1632);
nor U1821 (N_1821,N_1696,N_1648);
nor U1822 (N_1822,N_1618,N_1727);
and U1823 (N_1823,N_1733,N_1628);
nor U1824 (N_1824,N_1787,N_1707);
and U1825 (N_1825,N_1621,N_1680);
nor U1826 (N_1826,N_1738,N_1655);
nand U1827 (N_1827,N_1686,N_1620);
or U1828 (N_1828,N_1601,N_1755);
nor U1829 (N_1829,N_1705,N_1769);
nor U1830 (N_1830,N_1753,N_1763);
and U1831 (N_1831,N_1711,N_1607);
nor U1832 (N_1832,N_1788,N_1715);
nand U1833 (N_1833,N_1744,N_1737);
or U1834 (N_1834,N_1699,N_1683);
and U1835 (N_1835,N_1614,N_1645);
nor U1836 (N_1836,N_1764,N_1684);
and U1837 (N_1837,N_1702,N_1716);
nor U1838 (N_1838,N_1735,N_1703);
xor U1839 (N_1839,N_1762,N_1624);
and U1840 (N_1840,N_1606,N_1767);
nor U1841 (N_1841,N_1784,N_1709);
and U1842 (N_1842,N_1695,N_1676);
and U1843 (N_1843,N_1757,N_1770);
or U1844 (N_1844,N_1776,N_1633);
nand U1845 (N_1845,N_1758,N_1612);
and U1846 (N_1846,N_1692,N_1635);
and U1847 (N_1847,N_1602,N_1662);
or U1848 (N_1848,N_1605,N_1617);
xnor U1849 (N_1849,N_1778,N_1799);
nand U1850 (N_1850,N_1719,N_1780);
nand U1851 (N_1851,N_1688,N_1729);
and U1852 (N_1852,N_1677,N_1731);
nor U1853 (N_1853,N_1659,N_1634);
or U1854 (N_1854,N_1673,N_1782);
nor U1855 (N_1855,N_1795,N_1613);
and U1856 (N_1856,N_1600,N_1752);
nand U1857 (N_1857,N_1643,N_1790);
nor U1858 (N_1858,N_1750,N_1714);
nor U1859 (N_1859,N_1724,N_1685);
or U1860 (N_1860,N_1793,N_1641);
nand U1861 (N_1861,N_1781,N_1720);
and U1862 (N_1862,N_1654,N_1722);
nand U1863 (N_1863,N_1666,N_1728);
and U1864 (N_1864,N_1751,N_1736);
or U1865 (N_1865,N_1748,N_1682);
nor U1866 (N_1866,N_1639,N_1609);
nand U1867 (N_1867,N_1604,N_1642);
nor U1868 (N_1868,N_1610,N_1742);
nand U1869 (N_1869,N_1689,N_1783);
nor U1870 (N_1870,N_1698,N_1615);
or U1871 (N_1871,N_1723,N_1760);
nor U1872 (N_1872,N_1693,N_1739);
nor U1873 (N_1873,N_1743,N_1681);
and U1874 (N_1874,N_1741,N_1652);
nand U1875 (N_1875,N_1768,N_1772);
and U1876 (N_1876,N_1713,N_1653);
and U1877 (N_1877,N_1616,N_1646);
or U1878 (N_1878,N_1611,N_1773);
nor U1879 (N_1879,N_1712,N_1754);
or U1880 (N_1880,N_1747,N_1636);
or U1881 (N_1881,N_1668,N_1792);
and U1882 (N_1882,N_1700,N_1625);
nand U1883 (N_1883,N_1710,N_1730);
nor U1884 (N_1884,N_1717,N_1674);
and U1885 (N_1885,N_1701,N_1619);
or U1886 (N_1886,N_1629,N_1726);
nor U1887 (N_1887,N_1786,N_1796);
and U1888 (N_1888,N_1626,N_1789);
nor U1889 (N_1889,N_1678,N_1669);
and U1890 (N_1890,N_1798,N_1640);
nand U1891 (N_1891,N_1691,N_1623);
and U1892 (N_1892,N_1761,N_1664);
nand U1893 (N_1893,N_1661,N_1670);
nor U1894 (N_1894,N_1721,N_1794);
nor U1895 (N_1895,N_1679,N_1756);
or U1896 (N_1896,N_1766,N_1774);
nand U1897 (N_1897,N_1650,N_1627);
nand U1898 (N_1898,N_1672,N_1603);
nand U1899 (N_1899,N_1746,N_1649);
or U1900 (N_1900,N_1603,N_1656);
and U1901 (N_1901,N_1708,N_1735);
or U1902 (N_1902,N_1680,N_1786);
nand U1903 (N_1903,N_1706,N_1774);
nand U1904 (N_1904,N_1697,N_1601);
nand U1905 (N_1905,N_1658,N_1765);
nand U1906 (N_1906,N_1689,N_1653);
xnor U1907 (N_1907,N_1678,N_1623);
nor U1908 (N_1908,N_1616,N_1645);
and U1909 (N_1909,N_1775,N_1696);
nor U1910 (N_1910,N_1646,N_1674);
nor U1911 (N_1911,N_1729,N_1768);
or U1912 (N_1912,N_1700,N_1772);
xor U1913 (N_1913,N_1627,N_1724);
or U1914 (N_1914,N_1750,N_1768);
nand U1915 (N_1915,N_1756,N_1623);
nand U1916 (N_1916,N_1648,N_1758);
or U1917 (N_1917,N_1783,N_1709);
and U1918 (N_1918,N_1630,N_1676);
or U1919 (N_1919,N_1715,N_1686);
and U1920 (N_1920,N_1641,N_1660);
nand U1921 (N_1921,N_1660,N_1630);
and U1922 (N_1922,N_1604,N_1744);
nand U1923 (N_1923,N_1660,N_1757);
nand U1924 (N_1924,N_1680,N_1705);
nand U1925 (N_1925,N_1678,N_1706);
nor U1926 (N_1926,N_1687,N_1722);
or U1927 (N_1927,N_1662,N_1778);
nor U1928 (N_1928,N_1612,N_1653);
or U1929 (N_1929,N_1760,N_1638);
and U1930 (N_1930,N_1656,N_1773);
nand U1931 (N_1931,N_1754,N_1624);
and U1932 (N_1932,N_1605,N_1706);
xor U1933 (N_1933,N_1617,N_1771);
nor U1934 (N_1934,N_1638,N_1723);
or U1935 (N_1935,N_1629,N_1649);
nand U1936 (N_1936,N_1650,N_1653);
nand U1937 (N_1937,N_1673,N_1700);
and U1938 (N_1938,N_1619,N_1618);
and U1939 (N_1939,N_1684,N_1631);
nand U1940 (N_1940,N_1664,N_1605);
nor U1941 (N_1941,N_1729,N_1780);
and U1942 (N_1942,N_1764,N_1748);
or U1943 (N_1943,N_1651,N_1602);
or U1944 (N_1944,N_1693,N_1665);
and U1945 (N_1945,N_1772,N_1767);
and U1946 (N_1946,N_1657,N_1743);
nand U1947 (N_1947,N_1717,N_1766);
nor U1948 (N_1948,N_1688,N_1611);
and U1949 (N_1949,N_1611,N_1741);
and U1950 (N_1950,N_1614,N_1768);
nor U1951 (N_1951,N_1601,N_1645);
and U1952 (N_1952,N_1601,N_1674);
nand U1953 (N_1953,N_1664,N_1775);
or U1954 (N_1954,N_1655,N_1722);
and U1955 (N_1955,N_1780,N_1700);
or U1956 (N_1956,N_1775,N_1741);
nand U1957 (N_1957,N_1718,N_1676);
nand U1958 (N_1958,N_1702,N_1685);
xor U1959 (N_1959,N_1670,N_1648);
nand U1960 (N_1960,N_1690,N_1645);
nand U1961 (N_1961,N_1726,N_1702);
nand U1962 (N_1962,N_1709,N_1673);
or U1963 (N_1963,N_1757,N_1627);
and U1964 (N_1964,N_1765,N_1744);
or U1965 (N_1965,N_1608,N_1600);
nor U1966 (N_1966,N_1717,N_1788);
nand U1967 (N_1967,N_1744,N_1769);
nand U1968 (N_1968,N_1717,N_1646);
nand U1969 (N_1969,N_1772,N_1656);
nand U1970 (N_1970,N_1669,N_1796);
nand U1971 (N_1971,N_1680,N_1731);
nor U1972 (N_1972,N_1766,N_1665);
and U1973 (N_1973,N_1643,N_1663);
and U1974 (N_1974,N_1600,N_1739);
nor U1975 (N_1975,N_1662,N_1680);
and U1976 (N_1976,N_1739,N_1659);
nor U1977 (N_1977,N_1734,N_1600);
nand U1978 (N_1978,N_1605,N_1600);
nand U1979 (N_1979,N_1652,N_1734);
nor U1980 (N_1980,N_1716,N_1735);
and U1981 (N_1981,N_1617,N_1703);
or U1982 (N_1982,N_1774,N_1665);
or U1983 (N_1983,N_1781,N_1649);
or U1984 (N_1984,N_1782,N_1609);
and U1985 (N_1985,N_1660,N_1679);
and U1986 (N_1986,N_1622,N_1705);
and U1987 (N_1987,N_1608,N_1732);
or U1988 (N_1988,N_1604,N_1657);
and U1989 (N_1989,N_1758,N_1630);
and U1990 (N_1990,N_1760,N_1730);
and U1991 (N_1991,N_1704,N_1733);
or U1992 (N_1992,N_1710,N_1793);
nand U1993 (N_1993,N_1772,N_1780);
nand U1994 (N_1994,N_1635,N_1724);
nor U1995 (N_1995,N_1675,N_1641);
or U1996 (N_1996,N_1681,N_1700);
or U1997 (N_1997,N_1684,N_1622);
or U1998 (N_1998,N_1723,N_1769);
and U1999 (N_1999,N_1614,N_1620);
or U2000 (N_2000,N_1911,N_1927);
nor U2001 (N_2001,N_1808,N_1974);
nor U2002 (N_2002,N_1830,N_1868);
nand U2003 (N_2003,N_1972,N_1824);
or U2004 (N_2004,N_1811,N_1806);
or U2005 (N_2005,N_1930,N_1926);
xnor U2006 (N_2006,N_1891,N_1858);
or U2007 (N_2007,N_1860,N_1944);
nor U2008 (N_2008,N_1905,N_1897);
nor U2009 (N_2009,N_1872,N_1938);
nor U2010 (N_2010,N_1867,N_1948);
nor U2011 (N_2011,N_1870,N_1816);
and U2012 (N_2012,N_1864,N_1960);
or U2013 (N_2013,N_1940,N_1908);
and U2014 (N_2014,N_1980,N_1900);
nor U2015 (N_2015,N_1925,N_1801);
and U2016 (N_2016,N_1886,N_1871);
or U2017 (N_2017,N_1840,N_1943);
and U2018 (N_2018,N_1854,N_1996);
or U2019 (N_2019,N_1805,N_1861);
or U2020 (N_2020,N_1982,N_1896);
nor U2021 (N_2021,N_1903,N_1910);
nor U2022 (N_2022,N_1991,N_1950);
and U2023 (N_2023,N_1914,N_1822);
nor U2024 (N_2024,N_1906,N_1947);
nor U2025 (N_2025,N_1928,N_1856);
or U2026 (N_2026,N_1804,N_1841);
nor U2027 (N_2027,N_1931,N_1919);
or U2028 (N_2028,N_1848,N_1847);
nand U2029 (N_2029,N_1802,N_1971);
nor U2030 (N_2030,N_1998,N_1933);
and U2031 (N_2031,N_1877,N_1952);
nor U2032 (N_2032,N_1878,N_1865);
and U2033 (N_2033,N_1829,N_1941);
or U2034 (N_2034,N_1898,N_1812);
nor U2035 (N_2035,N_1885,N_1881);
nand U2036 (N_2036,N_1888,N_1907);
and U2037 (N_2037,N_1849,N_1855);
and U2038 (N_2038,N_1909,N_1922);
and U2039 (N_2039,N_1815,N_1875);
or U2040 (N_2040,N_1934,N_1969);
or U2041 (N_2041,N_1955,N_1874);
or U2042 (N_2042,N_1817,N_1992);
nor U2043 (N_2043,N_1857,N_1884);
nand U2044 (N_2044,N_1846,N_1820);
or U2045 (N_2045,N_1985,N_1995);
xnor U2046 (N_2046,N_1899,N_1832);
nand U2047 (N_2047,N_1945,N_1842);
or U2048 (N_2048,N_1895,N_1921);
and U2049 (N_2049,N_1970,N_1957);
or U2050 (N_2050,N_1976,N_1924);
or U2051 (N_2051,N_1892,N_1913);
nor U2052 (N_2052,N_1827,N_1862);
nor U2053 (N_2053,N_1978,N_1839);
and U2054 (N_2054,N_1965,N_1997);
or U2055 (N_2055,N_1828,N_1918);
or U2056 (N_2056,N_1807,N_1963);
and U2057 (N_2057,N_1959,N_1831);
or U2058 (N_2058,N_1939,N_1979);
nor U2059 (N_2059,N_1893,N_1879);
nor U2060 (N_2060,N_1835,N_1813);
nor U2061 (N_2061,N_1966,N_1958);
or U2062 (N_2062,N_1850,N_1912);
nand U2063 (N_2063,N_1826,N_1935);
or U2064 (N_2064,N_1803,N_1964);
or U2065 (N_2065,N_1956,N_1977);
and U2066 (N_2066,N_1929,N_1843);
nor U2067 (N_2067,N_1984,N_1880);
or U2068 (N_2068,N_1836,N_1818);
nand U2069 (N_2069,N_1988,N_1876);
or U2070 (N_2070,N_1953,N_1810);
nand U2071 (N_2071,N_1962,N_1869);
nor U2072 (N_2072,N_1983,N_1989);
nor U2073 (N_2073,N_1967,N_1890);
nand U2074 (N_2074,N_1916,N_1994);
nand U2075 (N_2075,N_1859,N_1981);
nor U2076 (N_2076,N_1999,N_1968);
nand U2077 (N_2077,N_1814,N_1961);
or U2078 (N_2078,N_1993,N_1904);
or U2079 (N_2079,N_1866,N_1894);
and U2080 (N_2080,N_1973,N_1821);
and U2081 (N_2081,N_1833,N_1863);
and U2082 (N_2082,N_1932,N_1987);
nand U2083 (N_2083,N_1873,N_1951);
nand U2084 (N_2084,N_1901,N_1853);
and U2085 (N_2085,N_1986,N_1949);
nand U2086 (N_2086,N_1837,N_1838);
nand U2087 (N_2087,N_1923,N_1845);
or U2088 (N_2088,N_1954,N_1946);
or U2089 (N_2089,N_1937,N_1825);
and U2090 (N_2090,N_1917,N_1851);
nor U2091 (N_2091,N_1809,N_1936);
nor U2092 (N_2092,N_1883,N_1902);
and U2093 (N_2093,N_1819,N_1882);
or U2094 (N_2094,N_1942,N_1975);
or U2095 (N_2095,N_1800,N_1852);
or U2096 (N_2096,N_1920,N_1887);
or U2097 (N_2097,N_1915,N_1823);
or U2098 (N_2098,N_1990,N_1844);
nor U2099 (N_2099,N_1834,N_1889);
nor U2100 (N_2100,N_1966,N_1909);
or U2101 (N_2101,N_1970,N_1864);
or U2102 (N_2102,N_1845,N_1905);
nor U2103 (N_2103,N_1846,N_1906);
nor U2104 (N_2104,N_1821,N_1978);
and U2105 (N_2105,N_1921,N_1966);
nor U2106 (N_2106,N_1816,N_1837);
nand U2107 (N_2107,N_1850,N_1806);
nor U2108 (N_2108,N_1821,N_1908);
nand U2109 (N_2109,N_1832,N_1895);
or U2110 (N_2110,N_1997,N_1868);
nand U2111 (N_2111,N_1890,N_1965);
nand U2112 (N_2112,N_1939,N_1880);
nand U2113 (N_2113,N_1973,N_1854);
or U2114 (N_2114,N_1991,N_1957);
and U2115 (N_2115,N_1868,N_1984);
and U2116 (N_2116,N_1907,N_1831);
nor U2117 (N_2117,N_1862,N_1876);
or U2118 (N_2118,N_1933,N_1815);
and U2119 (N_2119,N_1969,N_1833);
and U2120 (N_2120,N_1926,N_1993);
and U2121 (N_2121,N_1945,N_1952);
or U2122 (N_2122,N_1962,N_1971);
and U2123 (N_2123,N_1977,N_1803);
and U2124 (N_2124,N_1998,N_1818);
nor U2125 (N_2125,N_1819,N_1803);
or U2126 (N_2126,N_1885,N_1812);
nand U2127 (N_2127,N_1994,N_1816);
and U2128 (N_2128,N_1845,N_1812);
xnor U2129 (N_2129,N_1918,N_1945);
and U2130 (N_2130,N_1803,N_1847);
or U2131 (N_2131,N_1836,N_1976);
or U2132 (N_2132,N_1883,N_1848);
and U2133 (N_2133,N_1898,N_1827);
nand U2134 (N_2134,N_1997,N_1847);
nand U2135 (N_2135,N_1941,N_1802);
nand U2136 (N_2136,N_1831,N_1874);
nor U2137 (N_2137,N_1997,N_1848);
nand U2138 (N_2138,N_1848,N_1868);
nand U2139 (N_2139,N_1987,N_1880);
and U2140 (N_2140,N_1966,N_1854);
and U2141 (N_2141,N_1829,N_1811);
nand U2142 (N_2142,N_1938,N_1936);
nand U2143 (N_2143,N_1807,N_1904);
or U2144 (N_2144,N_1945,N_1869);
or U2145 (N_2145,N_1824,N_1880);
or U2146 (N_2146,N_1813,N_1802);
nand U2147 (N_2147,N_1896,N_1978);
or U2148 (N_2148,N_1820,N_1983);
nor U2149 (N_2149,N_1998,N_1803);
or U2150 (N_2150,N_1999,N_1854);
and U2151 (N_2151,N_1937,N_1885);
nand U2152 (N_2152,N_1866,N_1808);
nor U2153 (N_2153,N_1851,N_1801);
nand U2154 (N_2154,N_1947,N_1827);
nor U2155 (N_2155,N_1843,N_1893);
and U2156 (N_2156,N_1977,N_1887);
nand U2157 (N_2157,N_1998,N_1987);
and U2158 (N_2158,N_1939,N_1802);
and U2159 (N_2159,N_1952,N_1983);
and U2160 (N_2160,N_1855,N_1885);
or U2161 (N_2161,N_1856,N_1984);
nand U2162 (N_2162,N_1982,N_1865);
or U2163 (N_2163,N_1884,N_1947);
and U2164 (N_2164,N_1912,N_1863);
nor U2165 (N_2165,N_1836,N_1966);
nor U2166 (N_2166,N_1961,N_1970);
nand U2167 (N_2167,N_1839,N_1863);
and U2168 (N_2168,N_1816,N_1917);
or U2169 (N_2169,N_1878,N_1956);
nor U2170 (N_2170,N_1958,N_1933);
or U2171 (N_2171,N_1962,N_1826);
nand U2172 (N_2172,N_1997,N_1805);
nand U2173 (N_2173,N_1952,N_1950);
or U2174 (N_2174,N_1924,N_1811);
nor U2175 (N_2175,N_1897,N_1904);
and U2176 (N_2176,N_1968,N_1947);
nor U2177 (N_2177,N_1999,N_1865);
or U2178 (N_2178,N_1824,N_1976);
nor U2179 (N_2179,N_1933,N_1979);
or U2180 (N_2180,N_1854,N_1935);
or U2181 (N_2181,N_1992,N_1874);
or U2182 (N_2182,N_1810,N_1961);
and U2183 (N_2183,N_1970,N_1956);
and U2184 (N_2184,N_1823,N_1965);
and U2185 (N_2185,N_1894,N_1902);
nand U2186 (N_2186,N_1878,N_1967);
and U2187 (N_2187,N_1814,N_1937);
nor U2188 (N_2188,N_1964,N_1910);
or U2189 (N_2189,N_1948,N_1872);
nor U2190 (N_2190,N_1866,N_1820);
nor U2191 (N_2191,N_1911,N_1866);
and U2192 (N_2192,N_1992,N_1908);
or U2193 (N_2193,N_1834,N_1913);
or U2194 (N_2194,N_1884,N_1904);
and U2195 (N_2195,N_1912,N_1890);
nand U2196 (N_2196,N_1990,N_1981);
and U2197 (N_2197,N_1810,N_1903);
and U2198 (N_2198,N_1810,N_1937);
nand U2199 (N_2199,N_1805,N_1918);
and U2200 (N_2200,N_2153,N_2187);
or U2201 (N_2201,N_2087,N_2168);
nand U2202 (N_2202,N_2192,N_2091);
or U2203 (N_2203,N_2020,N_2054);
nor U2204 (N_2204,N_2171,N_2195);
or U2205 (N_2205,N_2036,N_2141);
or U2206 (N_2206,N_2169,N_2142);
and U2207 (N_2207,N_2010,N_2130);
nand U2208 (N_2208,N_2112,N_2197);
nand U2209 (N_2209,N_2066,N_2006);
and U2210 (N_2210,N_2179,N_2182);
nand U2211 (N_2211,N_2023,N_2085);
or U2212 (N_2212,N_2069,N_2031);
or U2213 (N_2213,N_2021,N_2003);
nor U2214 (N_2214,N_2181,N_2042);
and U2215 (N_2215,N_2198,N_2047);
or U2216 (N_2216,N_2022,N_2073);
or U2217 (N_2217,N_2136,N_2117);
and U2218 (N_2218,N_2034,N_2148);
and U2219 (N_2219,N_2164,N_2176);
nor U2220 (N_2220,N_2051,N_2184);
or U2221 (N_2221,N_2027,N_2009);
and U2222 (N_2222,N_2144,N_2055);
nor U2223 (N_2223,N_2107,N_2033);
nor U2224 (N_2224,N_2172,N_2167);
or U2225 (N_2225,N_2156,N_2145);
nor U2226 (N_2226,N_2143,N_2185);
and U2227 (N_2227,N_2123,N_2188);
and U2228 (N_2228,N_2108,N_2175);
xnor U2229 (N_2229,N_2100,N_2030);
or U2230 (N_2230,N_2097,N_2140);
and U2231 (N_2231,N_2056,N_2163);
nand U2232 (N_2232,N_2190,N_2057);
or U2233 (N_2233,N_2150,N_2102);
or U2234 (N_2234,N_2118,N_2154);
and U2235 (N_2235,N_2071,N_2060);
nand U2236 (N_2236,N_2106,N_2158);
and U2237 (N_2237,N_2129,N_2093);
or U2238 (N_2238,N_2196,N_2099);
and U2239 (N_2239,N_2132,N_2098);
nand U2240 (N_2240,N_2183,N_2008);
and U2241 (N_2241,N_2089,N_2079);
nand U2242 (N_2242,N_2090,N_2065);
nand U2243 (N_2243,N_2165,N_2180);
and U2244 (N_2244,N_2159,N_2084);
nor U2245 (N_2245,N_2124,N_2007);
nand U2246 (N_2246,N_2170,N_2199);
or U2247 (N_2247,N_2160,N_2113);
and U2248 (N_2248,N_2151,N_2037);
and U2249 (N_2249,N_2013,N_2149);
or U2250 (N_2250,N_2080,N_2041);
and U2251 (N_2251,N_2011,N_2146);
or U2252 (N_2252,N_2039,N_2038);
nand U2253 (N_2253,N_2194,N_2128);
or U2254 (N_2254,N_2035,N_2045);
and U2255 (N_2255,N_2127,N_2070);
and U2256 (N_2256,N_2024,N_2119);
nand U2257 (N_2257,N_2189,N_2115);
or U2258 (N_2258,N_2092,N_2072);
nand U2259 (N_2259,N_2001,N_2044);
nand U2260 (N_2260,N_2101,N_2178);
or U2261 (N_2261,N_2120,N_2116);
nor U2262 (N_2262,N_2134,N_2052);
nand U2263 (N_2263,N_2025,N_2053);
and U2264 (N_2264,N_2177,N_2138);
nor U2265 (N_2265,N_2157,N_2068);
nor U2266 (N_2266,N_2193,N_2147);
and U2267 (N_2267,N_2135,N_2046);
nor U2268 (N_2268,N_2064,N_2109);
nor U2269 (N_2269,N_2000,N_2152);
nor U2270 (N_2270,N_2078,N_2174);
or U2271 (N_2271,N_2014,N_2081);
or U2272 (N_2272,N_2186,N_2166);
and U2273 (N_2273,N_2032,N_2018);
nand U2274 (N_2274,N_2026,N_2058);
nand U2275 (N_2275,N_2004,N_2083);
nand U2276 (N_2276,N_2061,N_2076);
nor U2277 (N_2277,N_2050,N_2040);
or U2278 (N_2278,N_2049,N_2110);
nor U2279 (N_2279,N_2173,N_2028);
nand U2280 (N_2280,N_2122,N_2137);
and U2281 (N_2281,N_2017,N_2077);
or U2282 (N_2282,N_2074,N_2133);
and U2283 (N_2283,N_2059,N_2048);
and U2284 (N_2284,N_2094,N_2002);
or U2285 (N_2285,N_2121,N_2088);
xor U2286 (N_2286,N_2005,N_2114);
and U2287 (N_2287,N_2067,N_2191);
or U2288 (N_2288,N_2162,N_2096);
or U2289 (N_2289,N_2095,N_2155);
or U2290 (N_2290,N_2082,N_2015);
nand U2291 (N_2291,N_2043,N_2131);
or U2292 (N_2292,N_2016,N_2126);
nor U2293 (N_2293,N_2139,N_2029);
nand U2294 (N_2294,N_2103,N_2105);
or U2295 (N_2295,N_2062,N_2125);
and U2296 (N_2296,N_2075,N_2063);
or U2297 (N_2297,N_2012,N_2019);
and U2298 (N_2298,N_2086,N_2104);
nor U2299 (N_2299,N_2111,N_2161);
nor U2300 (N_2300,N_2031,N_2099);
nand U2301 (N_2301,N_2179,N_2011);
and U2302 (N_2302,N_2084,N_2073);
or U2303 (N_2303,N_2078,N_2125);
nor U2304 (N_2304,N_2048,N_2193);
nor U2305 (N_2305,N_2157,N_2072);
xor U2306 (N_2306,N_2109,N_2184);
nand U2307 (N_2307,N_2058,N_2117);
nor U2308 (N_2308,N_2044,N_2199);
nor U2309 (N_2309,N_2104,N_2028);
nor U2310 (N_2310,N_2166,N_2117);
nand U2311 (N_2311,N_2092,N_2040);
and U2312 (N_2312,N_2055,N_2016);
and U2313 (N_2313,N_2074,N_2159);
nand U2314 (N_2314,N_2199,N_2102);
nor U2315 (N_2315,N_2173,N_2185);
or U2316 (N_2316,N_2178,N_2009);
nand U2317 (N_2317,N_2038,N_2140);
or U2318 (N_2318,N_2100,N_2173);
nor U2319 (N_2319,N_2078,N_2013);
nor U2320 (N_2320,N_2079,N_2030);
or U2321 (N_2321,N_2100,N_2022);
nand U2322 (N_2322,N_2066,N_2018);
and U2323 (N_2323,N_2053,N_2136);
nand U2324 (N_2324,N_2022,N_2130);
nor U2325 (N_2325,N_2185,N_2011);
nand U2326 (N_2326,N_2075,N_2021);
nand U2327 (N_2327,N_2095,N_2093);
nand U2328 (N_2328,N_2146,N_2111);
or U2329 (N_2329,N_2048,N_2191);
nand U2330 (N_2330,N_2122,N_2108);
or U2331 (N_2331,N_2141,N_2030);
nand U2332 (N_2332,N_2114,N_2046);
nand U2333 (N_2333,N_2037,N_2076);
and U2334 (N_2334,N_2175,N_2042);
nand U2335 (N_2335,N_2076,N_2048);
or U2336 (N_2336,N_2139,N_2121);
and U2337 (N_2337,N_2113,N_2165);
nor U2338 (N_2338,N_2031,N_2109);
xor U2339 (N_2339,N_2066,N_2013);
nand U2340 (N_2340,N_2135,N_2113);
nand U2341 (N_2341,N_2169,N_2181);
nor U2342 (N_2342,N_2046,N_2071);
and U2343 (N_2343,N_2094,N_2129);
nor U2344 (N_2344,N_2130,N_2129);
nand U2345 (N_2345,N_2143,N_2186);
nor U2346 (N_2346,N_2053,N_2012);
nand U2347 (N_2347,N_2057,N_2051);
or U2348 (N_2348,N_2099,N_2067);
nand U2349 (N_2349,N_2008,N_2139);
xnor U2350 (N_2350,N_2079,N_2082);
and U2351 (N_2351,N_2167,N_2099);
nor U2352 (N_2352,N_2062,N_2185);
nand U2353 (N_2353,N_2108,N_2001);
and U2354 (N_2354,N_2128,N_2134);
nor U2355 (N_2355,N_2158,N_2099);
xor U2356 (N_2356,N_2011,N_2012);
or U2357 (N_2357,N_2185,N_2068);
and U2358 (N_2358,N_2140,N_2183);
or U2359 (N_2359,N_2059,N_2134);
nor U2360 (N_2360,N_2165,N_2135);
and U2361 (N_2361,N_2058,N_2012);
nand U2362 (N_2362,N_2031,N_2016);
and U2363 (N_2363,N_2084,N_2070);
nand U2364 (N_2364,N_2130,N_2072);
nor U2365 (N_2365,N_2094,N_2030);
and U2366 (N_2366,N_2199,N_2050);
or U2367 (N_2367,N_2057,N_2152);
and U2368 (N_2368,N_2083,N_2164);
or U2369 (N_2369,N_2058,N_2021);
nor U2370 (N_2370,N_2198,N_2089);
nand U2371 (N_2371,N_2141,N_2039);
or U2372 (N_2372,N_2073,N_2035);
or U2373 (N_2373,N_2058,N_2050);
or U2374 (N_2374,N_2096,N_2095);
and U2375 (N_2375,N_2046,N_2163);
and U2376 (N_2376,N_2088,N_2077);
nand U2377 (N_2377,N_2136,N_2145);
nand U2378 (N_2378,N_2164,N_2111);
nand U2379 (N_2379,N_2095,N_2048);
nor U2380 (N_2380,N_2105,N_2118);
nor U2381 (N_2381,N_2188,N_2103);
or U2382 (N_2382,N_2107,N_2061);
nor U2383 (N_2383,N_2150,N_2082);
nor U2384 (N_2384,N_2191,N_2152);
and U2385 (N_2385,N_2105,N_2042);
nand U2386 (N_2386,N_2046,N_2167);
nor U2387 (N_2387,N_2096,N_2063);
nand U2388 (N_2388,N_2027,N_2001);
or U2389 (N_2389,N_2196,N_2027);
and U2390 (N_2390,N_2153,N_2173);
nand U2391 (N_2391,N_2117,N_2193);
and U2392 (N_2392,N_2002,N_2140);
and U2393 (N_2393,N_2173,N_2122);
nor U2394 (N_2394,N_2096,N_2115);
or U2395 (N_2395,N_2020,N_2088);
and U2396 (N_2396,N_2073,N_2116);
nand U2397 (N_2397,N_2116,N_2093);
and U2398 (N_2398,N_2075,N_2053);
nand U2399 (N_2399,N_2009,N_2189);
nand U2400 (N_2400,N_2394,N_2359);
and U2401 (N_2401,N_2296,N_2294);
nand U2402 (N_2402,N_2271,N_2253);
or U2403 (N_2403,N_2309,N_2389);
nor U2404 (N_2404,N_2258,N_2300);
and U2405 (N_2405,N_2265,N_2344);
nand U2406 (N_2406,N_2384,N_2313);
nand U2407 (N_2407,N_2332,N_2319);
or U2408 (N_2408,N_2361,N_2301);
nor U2409 (N_2409,N_2208,N_2213);
or U2410 (N_2410,N_2312,N_2298);
nand U2411 (N_2411,N_2318,N_2293);
or U2412 (N_2412,N_2235,N_2368);
and U2413 (N_2413,N_2287,N_2207);
and U2414 (N_2414,N_2348,N_2383);
nor U2415 (N_2415,N_2279,N_2311);
nor U2416 (N_2416,N_2275,N_2218);
and U2417 (N_2417,N_2374,N_2393);
nand U2418 (N_2418,N_2222,N_2203);
and U2419 (N_2419,N_2372,N_2257);
and U2420 (N_2420,N_2283,N_2321);
nand U2421 (N_2421,N_2280,N_2270);
or U2422 (N_2422,N_2200,N_2328);
and U2423 (N_2423,N_2367,N_2205);
nor U2424 (N_2424,N_2269,N_2391);
nand U2425 (N_2425,N_2333,N_2288);
and U2426 (N_2426,N_2251,N_2291);
and U2427 (N_2427,N_2286,N_2252);
nor U2428 (N_2428,N_2254,N_2365);
and U2429 (N_2429,N_2375,N_2201);
nand U2430 (N_2430,N_2336,N_2340);
nor U2431 (N_2431,N_2234,N_2307);
nand U2432 (N_2432,N_2337,N_2245);
and U2433 (N_2433,N_2237,N_2354);
nand U2434 (N_2434,N_2268,N_2266);
and U2435 (N_2435,N_2238,N_2241);
nand U2436 (N_2436,N_2386,N_2398);
or U2437 (N_2437,N_2284,N_2343);
and U2438 (N_2438,N_2210,N_2352);
nor U2439 (N_2439,N_2338,N_2216);
nand U2440 (N_2440,N_2285,N_2320);
or U2441 (N_2441,N_2292,N_2364);
nor U2442 (N_2442,N_2395,N_2360);
or U2443 (N_2443,N_2295,N_2347);
or U2444 (N_2444,N_2370,N_2228);
and U2445 (N_2445,N_2224,N_2388);
and U2446 (N_2446,N_2304,N_2274);
and U2447 (N_2447,N_2392,N_2261);
nor U2448 (N_2448,N_2363,N_2249);
nor U2449 (N_2449,N_2366,N_2378);
or U2450 (N_2450,N_2263,N_2240);
or U2451 (N_2451,N_2396,N_2273);
and U2452 (N_2452,N_2331,N_2310);
or U2453 (N_2453,N_2248,N_2277);
or U2454 (N_2454,N_2397,N_2369);
nor U2455 (N_2455,N_2305,N_2390);
or U2456 (N_2456,N_2330,N_2355);
nand U2457 (N_2457,N_2329,N_2223);
nor U2458 (N_2458,N_2317,N_2204);
and U2459 (N_2459,N_2242,N_2399);
and U2460 (N_2460,N_2356,N_2231);
nor U2461 (N_2461,N_2385,N_2221);
or U2462 (N_2462,N_2316,N_2247);
and U2463 (N_2463,N_2230,N_2236);
or U2464 (N_2464,N_2358,N_2233);
nor U2465 (N_2465,N_2350,N_2353);
nand U2466 (N_2466,N_2219,N_2243);
and U2467 (N_2467,N_2299,N_2209);
nand U2468 (N_2468,N_2346,N_2227);
and U2469 (N_2469,N_2256,N_2267);
nand U2470 (N_2470,N_2325,N_2302);
or U2471 (N_2471,N_2308,N_2327);
nand U2472 (N_2472,N_2373,N_2381);
nor U2473 (N_2473,N_2206,N_2255);
or U2474 (N_2474,N_2239,N_2351);
nor U2475 (N_2475,N_2259,N_2377);
nand U2476 (N_2476,N_2212,N_2281);
nor U2477 (N_2477,N_2297,N_2289);
nand U2478 (N_2478,N_2315,N_2244);
and U2479 (N_2479,N_2246,N_2272);
nand U2480 (N_2480,N_2326,N_2362);
or U2481 (N_2481,N_2260,N_2282);
and U2482 (N_2482,N_2220,N_2323);
nand U2483 (N_2483,N_2229,N_2349);
and U2484 (N_2484,N_2339,N_2226);
nand U2485 (N_2485,N_2290,N_2376);
and U2486 (N_2486,N_2303,N_2306);
or U2487 (N_2487,N_2341,N_2314);
or U2488 (N_2488,N_2322,N_2382);
or U2489 (N_2489,N_2379,N_2214);
and U2490 (N_2490,N_2225,N_2357);
nand U2491 (N_2491,N_2371,N_2380);
nor U2492 (N_2492,N_2264,N_2342);
and U2493 (N_2493,N_2335,N_2232);
and U2494 (N_2494,N_2215,N_2345);
nand U2495 (N_2495,N_2250,N_2278);
nor U2496 (N_2496,N_2211,N_2334);
and U2497 (N_2497,N_2202,N_2217);
and U2498 (N_2498,N_2276,N_2262);
or U2499 (N_2499,N_2387,N_2324);
and U2500 (N_2500,N_2273,N_2203);
nand U2501 (N_2501,N_2219,N_2358);
nand U2502 (N_2502,N_2280,N_2328);
nor U2503 (N_2503,N_2235,N_2228);
nor U2504 (N_2504,N_2378,N_2208);
and U2505 (N_2505,N_2332,N_2352);
nand U2506 (N_2506,N_2214,N_2383);
and U2507 (N_2507,N_2231,N_2375);
and U2508 (N_2508,N_2245,N_2211);
nand U2509 (N_2509,N_2302,N_2393);
nor U2510 (N_2510,N_2254,N_2212);
nand U2511 (N_2511,N_2273,N_2307);
nor U2512 (N_2512,N_2245,N_2222);
and U2513 (N_2513,N_2341,N_2317);
and U2514 (N_2514,N_2245,N_2355);
nor U2515 (N_2515,N_2228,N_2304);
nor U2516 (N_2516,N_2356,N_2335);
or U2517 (N_2517,N_2252,N_2287);
nor U2518 (N_2518,N_2317,N_2216);
or U2519 (N_2519,N_2384,N_2303);
or U2520 (N_2520,N_2217,N_2335);
nor U2521 (N_2521,N_2307,N_2257);
or U2522 (N_2522,N_2313,N_2348);
and U2523 (N_2523,N_2256,N_2217);
nor U2524 (N_2524,N_2290,N_2357);
nor U2525 (N_2525,N_2266,N_2289);
nor U2526 (N_2526,N_2298,N_2319);
nand U2527 (N_2527,N_2201,N_2240);
nand U2528 (N_2528,N_2247,N_2293);
nor U2529 (N_2529,N_2383,N_2200);
or U2530 (N_2530,N_2254,N_2287);
or U2531 (N_2531,N_2247,N_2323);
nand U2532 (N_2532,N_2213,N_2254);
or U2533 (N_2533,N_2325,N_2376);
or U2534 (N_2534,N_2290,N_2258);
and U2535 (N_2535,N_2337,N_2305);
nand U2536 (N_2536,N_2385,N_2280);
nand U2537 (N_2537,N_2358,N_2250);
or U2538 (N_2538,N_2310,N_2275);
or U2539 (N_2539,N_2291,N_2286);
nor U2540 (N_2540,N_2203,N_2218);
nor U2541 (N_2541,N_2259,N_2303);
nor U2542 (N_2542,N_2272,N_2291);
nor U2543 (N_2543,N_2375,N_2385);
or U2544 (N_2544,N_2258,N_2251);
and U2545 (N_2545,N_2203,N_2391);
and U2546 (N_2546,N_2333,N_2369);
nor U2547 (N_2547,N_2395,N_2376);
nor U2548 (N_2548,N_2257,N_2240);
and U2549 (N_2549,N_2222,N_2286);
or U2550 (N_2550,N_2202,N_2259);
nor U2551 (N_2551,N_2200,N_2385);
nor U2552 (N_2552,N_2322,N_2294);
nor U2553 (N_2553,N_2248,N_2229);
and U2554 (N_2554,N_2262,N_2313);
nand U2555 (N_2555,N_2360,N_2289);
or U2556 (N_2556,N_2219,N_2259);
nor U2557 (N_2557,N_2308,N_2305);
and U2558 (N_2558,N_2317,N_2316);
nand U2559 (N_2559,N_2311,N_2356);
and U2560 (N_2560,N_2387,N_2269);
and U2561 (N_2561,N_2314,N_2324);
nand U2562 (N_2562,N_2343,N_2214);
nor U2563 (N_2563,N_2323,N_2222);
and U2564 (N_2564,N_2313,N_2381);
and U2565 (N_2565,N_2253,N_2385);
nor U2566 (N_2566,N_2217,N_2369);
and U2567 (N_2567,N_2298,N_2330);
nand U2568 (N_2568,N_2214,N_2273);
or U2569 (N_2569,N_2234,N_2245);
or U2570 (N_2570,N_2254,N_2307);
nand U2571 (N_2571,N_2285,N_2222);
and U2572 (N_2572,N_2361,N_2331);
nand U2573 (N_2573,N_2270,N_2351);
or U2574 (N_2574,N_2368,N_2261);
nand U2575 (N_2575,N_2218,N_2265);
nor U2576 (N_2576,N_2349,N_2212);
or U2577 (N_2577,N_2220,N_2354);
or U2578 (N_2578,N_2389,N_2265);
nand U2579 (N_2579,N_2395,N_2319);
and U2580 (N_2580,N_2204,N_2205);
or U2581 (N_2581,N_2316,N_2371);
nor U2582 (N_2582,N_2339,N_2233);
nand U2583 (N_2583,N_2249,N_2240);
nand U2584 (N_2584,N_2214,N_2317);
nand U2585 (N_2585,N_2332,N_2320);
nand U2586 (N_2586,N_2220,N_2246);
nand U2587 (N_2587,N_2320,N_2358);
nand U2588 (N_2588,N_2255,N_2389);
nor U2589 (N_2589,N_2334,N_2357);
or U2590 (N_2590,N_2313,N_2234);
nand U2591 (N_2591,N_2332,N_2219);
and U2592 (N_2592,N_2225,N_2288);
xnor U2593 (N_2593,N_2364,N_2387);
nor U2594 (N_2594,N_2373,N_2337);
or U2595 (N_2595,N_2306,N_2299);
nand U2596 (N_2596,N_2311,N_2260);
nand U2597 (N_2597,N_2352,N_2295);
and U2598 (N_2598,N_2324,N_2261);
and U2599 (N_2599,N_2273,N_2376);
and U2600 (N_2600,N_2497,N_2402);
or U2601 (N_2601,N_2512,N_2415);
or U2602 (N_2602,N_2541,N_2517);
or U2603 (N_2603,N_2563,N_2555);
and U2604 (N_2604,N_2448,N_2592);
nor U2605 (N_2605,N_2521,N_2476);
nand U2606 (N_2606,N_2425,N_2525);
or U2607 (N_2607,N_2407,N_2438);
or U2608 (N_2608,N_2470,N_2573);
or U2609 (N_2609,N_2428,N_2460);
nor U2610 (N_2610,N_2458,N_2534);
nand U2611 (N_2611,N_2400,N_2499);
nor U2612 (N_2612,N_2440,N_2526);
xor U2613 (N_2613,N_2543,N_2432);
or U2614 (N_2614,N_2447,N_2467);
or U2615 (N_2615,N_2597,N_2430);
nand U2616 (N_2616,N_2527,N_2477);
or U2617 (N_2617,N_2533,N_2551);
nor U2618 (N_2618,N_2565,N_2537);
and U2619 (N_2619,N_2519,N_2417);
nor U2620 (N_2620,N_2464,N_2511);
nand U2621 (N_2621,N_2596,N_2548);
xor U2622 (N_2622,N_2446,N_2578);
and U2623 (N_2623,N_2462,N_2404);
or U2624 (N_2624,N_2522,N_2545);
and U2625 (N_2625,N_2479,N_2556);
nand U2626 (N_2626,N_2427,N_2410);
or U2627 (N_2627,N_2546,N_2564);
nand U2628 (N_2628,N_2593,N_2409);
nor U2629 (N_2629,N_2496,N_2408);
nor U2630 (N_2630,N_2406,N_2574);
nand U2631 (N_2631,N_2450,N_2444);
or U2632 (N_2632,N_2507,N_2423);
or U2633 (N_2633,N_2435,N_2481);
and U2634 (N_2634,N_2572,N_2535);
or U2635 (N_2635,N_2513,N_2530);
nand U2636 (N_2636,N_2516,N_2552);
nand U2637 (N_2637,N_2451,N_2480);
nor U2638 (N_2638,N_2472,N_2567);
nand U2639 (N_2639,N_2580,N_2598);
or U2640 (N_2640,N_2483,N_2413);
nor U2641 (N_2641,N_2579,N_2532);
nor U2642 (N_2642,N_2515,N_2494);
nor U2643 (N_2643,N_2431,N_2503);
or U2644 (N_2644,N_2436,N_2416);
and U2645 (N_2645,N_2456,N_2487);
nand U2646 (N_2646,N_2424,N_2520);
and U2647 (N_2647,N_2581,N_2455);
or U2648 (N_2648,N_2486,N_2412);
nor U2649 (N_2649,N_2506,N_2557);
and U2650 (N_2650,N_2585,N_2569);
nand U2651 (N_2651,N_2442,N_2586);
nand U2652 (N_2652,N_2414,N_2489);
nand U2653 (N_2653,N_2491,N_2492);
nand U2654 (N_2654,N_2550,N_2590);
nand U2655 (N_2655,N_2478,N_2401);
and U2656 (N_2656,N_2473,N_2419);
and U2657 (N_2657,N_2547,N_2453);
nand U2658 (N_2658,N_2509,N_2465);
nand U2659 (N_2659,N_2544,N_2421);
nor U2660 (N_2660,N_2463,N_2576);
nor U2661 (N_2661,N_2488,N_2538);
nor U2662 (N_2662,N_2536,N_2542);
nand U2663 (N_2663,N_2434,N_2518);
or U2664 (N_2664,N_2452,N_2571);
nand U2665 (N_2665,N_2474,N_2403);
or U2666 (N_2666,N_2498,N_2549);
nor U2667 (N_2667,N_2469,N_2554);
or U2668 (N_2668,N_2568,N_2422);
or U2669 (N_2669,N_2495,N_2587);
or U2670 (N_2670,N_2457,N_2594);
or U2671 (N_2671,N_2529,N_2466);
or U2672 (N_2672,N_2405,N_2454);
or U2673 (N_2673,N_2539,N_2429);
nand U2674 (N_2674,N_2584,N_2540);
or U2675 (N_2675,N_2411,N_2500);
and U2676 (N_2676,N_2468,N_2426);
or U2677 (N_2677,N_2583,N_2553);
or U2678 (N_2678,N_2504,N_2591);
nor U2679 (N_2679,N_2441,N_2418);
nor U2680 (N_2680,N_2501,N_2439);
or U2681 (N_2681,N_2433,N_2570);
nor U2682 (N_2682,N_2475,N_2459);
nand U2683 (N_2683,N_2582,N_2490);
and U2684 (N_2684,N_2562,N_2485);
nor U2685 (N_2685,N_2589,N_2599);
or U2686 (N_2686,N_2505,N_2445);
xor U2687 (N_2687,N_2566,N_2528);
nor U2688 (N_2688,N_2493,N_2523);
nor U2689 (N_2689,N_2449,N_2461);
and U2690 (N_2690,N_2577,N_2482);
xnor U2691 (N_2691,N_2531,N_2595);
nand U2692 (N_2692,N_2560,N_2559);
and U2693 (N_2693,N_2524,N_2420);
or U2694 (N_2694,N_2471,N_2502);
or U2695 (N_2695,N_2510,N_2484);
or U2696 (N_2696,N_2575,N_2588);
nand U2697 (N_2697,N_2561,N_2514);
nor U2698 (N_2698,N_2437,N_2443);
nor U2699 (N_2699,N_2558,N_2508);
and U2700 (N_2700,N_2455,N_2406);
nand U2701 (N_2701,N_2538,N_2418);
nor U2702 (N_2702,N_2597,N_2486);
or U2703 (N_2703,N_2483,N_2404);
nand U2704 (N_2704,N_2571,N_2537);
or U2705 (N_2705,N_2421,N_2433);
nand U2706 (N_2706,N_2404,N_2484);
nand U2707 (N_2707,N_2530,N_2407);
and U2708 (N_2708,N_2470,N_2574);
or U2709 (N_2709,N_2598,N_2495);
nor U2710 (N_2710,N_2492,N_2549);
nand U2711 (N_2711,N_2518,N_2535);
nor U2712 (N_2712,N_2475,N_2466);
nor U2713 (N_2713,N_2424,N_2584);
or U2714 (N_2714,N_2511,N_2595);
nand U2715 (N_2715,N_2558,N_2493);
nor U2716 (N_2716,N_2566,N_2543);
and U2717 (N_2717,N_2408,N_2555);
or U2718 (N_2718,N_2506,N_2438);
nor U2719 (N_2719,N_2431,N_2417);
nor U2720 (N_2720,N_2453,N_2483);
and U2721 (N_2721,N_2412,N_2562);
or U2722 (N_2722,N_2588,N_2568);
nand U2723 (N_2723,N_2478,N_2519);
and U2724 (N_2724,N_2565,N_2463);
and U2725 (N_2725,N_2488,N_2442);
and U2726 (N_2726,N_2483,N_2531);
nor U2727 (N_2727,N_2580,N_2444);
or U2728 (N_2728,N_2503,N_2591);
nor U2729 (N_2729,N_2565,N_2417);
or U2730 (N_2730,N_2472,N_2465);
and U2731 (N_2731,N_2510,N_2458);
and U2732 (N_2732,N_2432,N_2570);
xor U2733 (N_2733,N_2532,N_2530);
or U2734 (N_2734,N_2482,N_2400);
or U2735 (N_2735,N_2536,N_2482);
and U2736 (N_2736,N_2562,N_2453);
and U2737 (N_2737,N_2446,N_2416);
nand U2738 (N_2738,N_2458,N_2408);
nand U2739 (N_2739,N_2467,N_2582);
nor U2740 (N_2740,N_2424,N_2540);
and U2741 (N_2741,N_2475,N_2574);
nand U2742 (N_2742,N_2576,N_2418);
nand U2743 (N_2743,N_2400,N_2414);
or U2744 (N_2744,N_2575,N_2495);
or U2745 (N_2745,N_2554,N_2462);
or U2746 (N_2746,N_2532,N_2425);
nor U2747 (N_2747,N_2488,N_2536);
nor U2748 (N_2748,N_2599,N_2419);
nor U2749 (N_2749,N_2415,N_2471);
nor U2750 (N_2750,N_2436,N_2441);
or U2751 (N_2751,N_2438,N_2443);
or U2752 (N_2752,N_2411,N_2529);
nor U2753 (N_2753,N_2486,N_2449);
or U2754 (N_2754,N_2469,N_2400);
nand U2755 (N_2755,N_2569,N_2541);
or U2756 (N_2756,N_2437,N_2526);
nor U2757 (N_2757,N_2564,N_2513);
nor U2758 (N_2758,N_2567,N_2436);
and U2759 (N_2759,N_2557,N_2498);
and U2760 (N_2760,N_2591,N_2564);
nor U2761 (N_2761,N_2486,N_2533);
nor U2762 (N_2762,N_2514,N_2549);
or U2763 (N_2763,N_2466,N_2408);
and U2764 (N_2764,N_2512,N_2441);
nor U2765 (N_2765,N_2546,N_2512);
nand U2766 (N_2766,N_2508,N_2503);
or U2767 (N_2767,N_2456,N_2569);
or U2768 (N_2768,N_2525,N_2570);
and U2769 (N_2769,N_2574,N_2459);
nand U2770 (N_2770,N_2573,N_2505);
or U2771 (N_2771,N_2524,N_2488);
and U2772 (N_2772,N_2527,N_2495);
and U2773 (N_2773,N_2573,N_2551);
nand U2774 (N_2774,N_2460,N_2432);
nand U2775 (N_2775,N_2473,N_2465);
nand U2776 (N_2776,N_2483,N_2578);
nor U2777 (N_2777,N_2442,N_2445);
or U2778 (N_2778,N_2486,N_2538);
or U2779 (N_2779,N_2495,N_2546);
or U2780 (N_2780,N_2500,N_2563);
and U2781 (N_2781,N_2515,N_2521);
or U2782 (N_2782,N_2432,N_2540);
nor U2783 (N_2783,N_2599,N_2453);
or U2784 (N_2784,N_2578,N_2563);
nor U2785 (N_2785,N_2430,N_2557);
xnor U2786 (N_2786,N_2508,N_2585);
nor U2787 (N_2787,N_2434,N_2499);
nand U2788 (N_2788,N_2561,N_2509);
nand U2789 (N_2789,N_2593,N_2580);
nand U2790 (N_2790,N_2552,N_2446);
or U2791 (N_2791,N_2578,N_2564);
and U2792 (N_2792,N_2469,N_2527);
nand U2793 (N_2793,N_2489,N_2438);
xor U2794 (N_2794,N_2564,N_2511);
and U2795 (N_2795,N_2407,N_2527);
or U2796 (N_2796,N_2478,N_2485);
and U2797 (N_2797,N_2423,N_2417);
and U2798 (N_2798,N_2510,N_2404);
and U2799 (N_2799,N_2512,N_2463);
or U2800 (N_2800,N_2613,N_2633);
and U2801 (N_2801,N_2722,N_2745);
or U2802 (N_2802,N_2796,N_2636);
or U2803 (N_2803,N_2632,N_2711);
nand U2804 (N_2804,N_2799,N_2716);
nand U2805 (N_2805,N_2659,N_2752);
and U2806 (N_2806,N_2753,N_2707);
and U2807 (N_2807,N_2750,N_2611);
and U2808 (N_2808,N_2790,N_2676);
nand U2809 (N_2809,N_2762,N_2712);
and U2810 (N_2810,N_2781,N_2774);
and U2811 (N_2811,N_2673,N_2657);
nor U2812 (N_2812,N_2728,N_2714);
nor U2813 (N_2813,N_2688,N_2606);
and U2814 (N_2814,N_2637,N_2685);
nand U2815 (N_2815,N_2620,N_2610);
and U2816 (N_2816,N_2731,N_2699);
and U2817 (N_2817,N_2694,N_2737);
xor U2818 (N_2818,N_2776,N_2644);
nand U2819 (N_2819,N_2618,N_2643);
and U2820 (N_2820,N_2623,N_2721);
and U2821 (N_2821,N_2603,N_2748);
and U2822 (N_2822,N_2706,N_2769);
nor U2823 (N_2823,N_2746,N_2786);
nand U2824 (N_2824,N_2635,N_2780);
and U2825 (N_2825,N_2718,N_2724);
nand U2826 (N_2826,N_2624,N_2761);
nor U2827 (N_2827,N_2678,N_2634);
and U2828 (N_2828,N_2649,N_2726);
or U2829 (N_2829,N_2640,N_2729);
or U2830 (N_2830,N_2691,N_2646);
nand U2831 (N_2831,N_2742,N_2789);
nand U2832 (N_2832,N_2720,N_2677);
nor U2833 (N_2833,N_2642,N_2681);
nor U2834 (N_2834,N_2604,N_2704);
or U2835 (N_2835,N_2671,N_2727);
nor U2836 (N_2836,N_2669,N_2747);
or U2837 (N_2837,N_2626,N_2741);
nand U2838 (N_2838,N_2692,N_2791);
or U2839 (N_2839,N_2768,N_2738);
xnor U2840 (N_2840,N_2730,N_2775);
and U2841 (N_2841,N_2600,N_2725);
nand U2842 (N_2842,N_2693,N_2614);
nor U2843 (N_2843,N_2653,N_2700);
nand U2844 (N_2844,N_2703,N_2670);
nor U2845 (N_2845,N_2719,N_2663);
and U2846 (N_2846,N_2629,N_2661);
nor U2847 (N_2847,N_2602,N_2755);
and U2848 (N_2848,N_2638,N_2621);
and U2849 (N_2849,N_2680,N_2749);
and U2850 (N_2850,N_2788,N_2630);
nor U2851 (N_2851,N_2765,N_2645);
nand U2852 (N_2852,N_2708,N_2601);
nand U2853 (N_2853,N_2715,N_2784);
or U2854 (N_2854,N_2683,N_2734);
or U2855 (N_2855,N_2655,N_2713);
nand U2856 (N_2856,N_2664,N_2660);
and U2857 (N_2857,N_2736,N_2666);
nand U2858 (N_2858,N_2798,N_2619);
nand U2859 (N_2859,N_2639,N_2656);
nand U2860 (N_2860,N_2609,N_2735);
xor U2861 (N_2861,N_2760,N_2710);
or U2862 (N_2862,N_2701,N_2605);
and U2863 (N_2863,N_2665,N_2744);
and U2864 (N_2864,N_2687,N_2675);
or U2865 (N_2865,N_2773,N_2641);
nand U2866 (N_2866,N_2785,N_2672);
or U2867 (N_2867,N_2662,N_2758);
and U2868 (N_2868,N_2767,N_2771);
or U2869 (N_2869,N_2794,N_2782);
and U2870 (N_2870,N_2766,N_2770);
or U2871 (N_2871,N_2732,N_2757);
nor U2872 (N_2872,N_2612,N_2616);
nor U2873 (N_2873,N_2777,N_2608);
nor U2874 (N_2874,N_2651,N_2650);
or U2875 (N_2875,N_2743,N_2698);
and U2876 (N_2876,N_2695,N_2679);
and U2877 (N_2877,N_2607,N_2702);
nand U2878 (N_2878,N_2756,N_2690);
nor U2879 (N_2879,N_2686,N_2717);
or U2880 (N_2880,N_2668,N_2797);
and U2881 (N_2881,N_2625,N_2733);
and U2882 (N_2882,N_2648,N_2764);
nand U2883 (N_2883,N_2795,N_2763);
nor U2884 (N_2884,N_2652,N_2617);
nand U2885 (N_2885,N_2631,N_2772);
nor U2886 (N_2886,N_2759,N_2622);
nand U2887 (N_2887,N_2684,N_2723);
and U2888 (N_2888,N_2787,N_2783);
nand U2889 (N_2889,N_2647,N_2682);
and U2890 (N_2890,N_2696,N_2740);
or U2891 (N_2891,N_2658,N_2739);
and U2892 (N_2892,N_2792,N_2778);
or U2893 (N_2893,N_2628,N_2689);
nor U2894 (N_2894,N_2627,N_2754);
and U2895 (N_2895,N_2793,N_2674);
or U2896 (N_2896,N_2697,N_2779);
xor U2897 (N_2897,N_2667,N_2654);
nor U2898 (N_2898,N_2615,N_2705);
nand U2899 (N_2899,N_2751,N_2709);
nor U2900 (N_2900,N_2775,N_2702);
and U2901 (N_2901,N_2703,N_2786);
nand U2902 (N_2902,N_2631,N_2723);
nand U2903 (N_2903,N_2728,N_2691);
nand U2904 (N_2904,N_2726,N_2608);
or U2905 (N_2905,N_2728,N_2782);
and U2906 (N_2906,N_2724,N_2642);
nand U2907 (N_2907,N_2710,N_2742);
and U2908 (N_2908,N_2793,N_2656);
nor U2909 (N_2909,N_2723,N_2727);
and U2910 (N_2910,N_2637,N_2782);
nand U2911 (N_2911,N_2751,N_2670);
and U2912 (N_2912,N_2775,N_2688);
and U2913 (N_2913,N_2649,N_2702);
and U2914 (N_2914,N_2632,N_2623);
or U2915 (N_2915,N_2695,N_2622);
and U2916 (N_2916,N_2670,N_2665);
or U2917 (N_2917,N_2775,N_2665);
nand U2918 (N_2918,N_2685,N_2760);
and U2919 (N_2919,N_2719,N_2608);
nand U2920 (N_2920,N_2679,N_2657);
or U2921 (N_2921,N_2779,N_2767);
nor U2922 (N_2922,N_2624,N_2771);
or U2923 (N_2923,N_2718,N_2629);
nor U2924 (N_2924,N_2676,N_2785);
nor U2925 (N_2925,N_2623,N_2700);
nor U2926 (N_2926,N_2698,N_2769);
and U2927 (N_2927,N_2748,N_2636);
and U2928 (N_2928,N_2718,N_2635);
or U2929 (N_2929,N_2620,N_2629);
nor U2930 (N_2930,N_2748,N_2708);
and U2931 (N_2931,N_2623,N_2649);
and U2932 (N_2932,N_2743,N_2670);
or U2933 (N_2933,N_2627,N_2752);
and U2934 (N_2934,N_2727,N_2735);
or U2935 (N_2935,N_2763,N_2657);
or U2936 (N_2936,N_2753,N_2665);
nor U2937 (N_2937,N_2766,N_2630);
nor U2938 (N_2938,N_2789,N_2641);
nand U2939 (N_2939,N_2659,N_2701);
and U2940 (N_2940,N_2651,N_2680);
or U2941 (N_2941,N_2779,N_2686);
and U2942 (N_2942,N_2635,N_2646);
nor U2943 (N_2943,N_2689,N_2630);
nor U2944 (N_2944,N_2701,N_2620);
nor U2945 (N_2945,N_2777,N_2653);
and U2946 (N_2946,N_2725,N_2643);
nor U2947 (N_2947,N_2634,N_2740);
nand U2948 (N_2948,N_2617,N_2729);
xnor U2949 (N_2949,N_2743,N_2652);
nand U2950 (N_2950,N_2663,N_2642);
and U2951 (N_2951,N_2673,N_2675);
nor U2952 (N_2952,N_2750,N_2663);
and U2953 (N_2953,N_2605,N_2775);
nand U2954 (N_2954,N_2770,N_2719);
or U2955 (N_2955,N_2616,N_2785);
and U2956 (N_2956,N_2757,N_2600);
nand U2957 (N_2957,N_2730,N_2761);
and U2958 (N_2958,N_2700,N_2794);
or U2959 (N_2959,N_2714,N_2640);
or U2960 (N_2960,N_2649,N_2639);
nor U2961 (N_2961,N_2609,N_2698);
and U2962 (N_2962,N_2659,N_2755);
or U2963 (N_2963,N_2752,N_2735);
and U2964 (N_2964,N_2778,N_2690);
nor U2965 (N_2965,N_2632,N_2663);
nor U2966 (N_2966,N_2619,N_2639);
or U2967 (N_2967,N_2610,N_2687);
nor U2968 (N_2968,N_2753,N_2648);
nand U2969 (N_2969,N_2666,N_2641);
nor U2970 (N_2970,N_2715,N_2687);
nand U2971 (N_2971,N_2777,N_2722);
or U2972 (N_2972,N_2710,N_2650);
nand U2973 (N_2973,N_2725,N_2676);
or U2974 (N_2974,N_2678,N_2704);
nor U2975 (N_2975,N_2700,N_2662);
nand U2976 (N_2976,N_2783,N_2641);
nor U2977 (N_2977,N_2713,N_2605);
and U2978 (N_2978,N_2705,N_2675);
nor U2979 (N_2979,N_2737,N_2643);
or U2980 (N_2980,N_2686,N_2607);
and U2981 (N_2981,N_2652,N_2673);
or U2982 (N_2982,N_2703,N_2659);
nor U2983 (N_2983,N_2617,N_2772);
nand U2984 (N_2984,N_2674,N_2747);
nor U2985 (N_2985,N_2757,N_2692);
or U2986 (N_2986,N_2766,N_2731);
or U2987 (N_2987,N_2770,N_2708);
or U2988 (N_2988,N_2672,N_2794);
nor U2989 (N_2989,N_2629,N_2697);
nor U2990 (N_2990,N_2616,N_2776);
or U2991 (N_2991,N_2716,N_2680);
or U2992 (N_2992,N_2605,N_2771);
and U2993 (N_2993,N_2638,N_2663);
and U2994 (N_2994,N_2738,N_2611);
or U2995 (N_2995,N_2750,N_2691);
and U2996 (N_2996,N_2768,N_2709);
nand U2997 (N_2997,N_2670,N_2676);
and U2998 (N_2998,N_2637,N_2640);
and U2999 (N_2999,N_2630,N_2783);
nor UO_0 (O_0,N_2968,N_2813);
and UO_1 (O_1,N_2880,N_2920);
nor UO_2 (O_2,N_2898,N_2985);
nor UO_3 (O_3,N_2927,N_2815);
or UO_4 (O_4,N_2853,N_2888);
nand UO_5 (O_5,N_2944,N_2861);
nor UO_6 (O_6,N_2928,N_2940);
nor UO_7 (O_7,N_2834,N_2895);
or UO_8 (O_8,N_2903,N_2860);
nand UO_9 (O_9,N_2962,N_2823);
and UO_10 (O_10,N_2977,N_2907);
nor UO_11 (O_11,N_2837,N_2824);
nand UO_12 (O_12,N_2970,N_2878);
nor UO_13 (O_13,N_2805,N_2839);
and UO_14 (O_14,N_2992,N_2842);
or UO_15 (O_15,N_2800,N_2828);
or UO_16 (O_16,N_2885,N_2804);
or UO_17 (O_17,N_2955,N_2922);
nor UO_18 (O_18,N_2835,N_2929);
nand UO_19 (O_19,N_2990,N_2961);
nor UO_20 (O_20,N_2825,N_2986);
and UO_21 (O_21,N_2900,N_2877);
nand UO_22 (O_22,N_2971,N_2956);
and UO_23 (O_23,N_2984,N_2943);
and UO_24 (O_24,N_2879,N_2822);
and UO_25 (O_25,N_2848,N_2849);
and UO_26 (O_26,N_2965,N_2854);
nand UO_27 (O_27,N_2869,N_2840);
nor UO_28 (O_28,N_2978,N_2957);
nor UO_29 (O_29,N_2906,N_2942);
or UO_30 (O_30,N_2874,N_2843);
or UO_31 (O_31,N_2999,N_2806);
nor UO_32 (O_32,N_2864,N_2989);
nor UO_33 (O_33,N_2908,N_2807);
nor UO_34 (O_34,N_2951,N_2924);
or UO_35 (O_35,N_2882,N_2847);
or UO_36 (O_36,N_2933,N_2896);
or UO_37 (O_37,N_2850,N_2892);
nand UO_38 (O_38,N_2960,N_2974);
or UO_39 (O_39,N_2803,N_2831);
nand UO_40 (O_40,N_2949,N_2959);
and UO_41 (O_41,N_2901,N_2904);
nor UO_42 (O_42,N_2991,N_2988);
and UO_43 (O_43,N_2858,N_2919);
or UO_44 (O_44,N_2964,N_2866);
or UO_45 (O_45,N_2863,N_2975);
and UO_46 (O_46,N_2923,N_2870);
nor UO_47 (O_47,N_2820,N_2830);
or UO_48 (O_48,N_2954,N_2812);
nand UO_49 (O_49,N_2899,N_2859);
and UO_50 (O_50,N_2818,N_2994);
nand UO_51 (O_51,N_2941,N_2969);
nand UO_52 (O_52,N_2987,N_2829);
and UO_53 (O_53,N_2816,N_2979);
nand UO_54 (O_54,N_2801,N_2889);
nor UO_55 (O_55,N_2881,N_2814);
and UO_56 (O_56,N_2873,N_2894);
nand UO_57 (O_57,N_2857,N_2841);
nor UO_58 (O_58,N_2911,N_2921);
nand UO_59 (O_59,N_2909,N_2890);
nor UO_60 (O_60,N_2967,N_2905);
nand UO_61 (O_61,N_2862,N_2947);
and UO_62 (O_62,N_2811,N_2997);
nand UO_63 (O_63,N_2817,N_2983);
nor UO_64 (O_64,N_2832,N_2876);
nor UO_65 (O_65,N_2809,N_2925);
or UO_66 (O_66,N_2852,N_2915);
nor UO_67 (O_67,N_2917,N_2993);
nand UO_68 (O_68,N_2948,N_2998);
and UO_69 (O_69,N_2946,N_2980);
nand UO_70 (O_70,N_2945,N_2950);
and UO_71 (O_71,N_2939,N_2884);
nand UO_72 (O_72,N_2958,N_2902);
or UO_73 (O_73,N_2918,N_2953);
and UO_74 (O_74,N_2838,N_2936);
or UO_75 (O_75,N_2808,N_2897);
nand UO_76 (O_76,N_2886,N_2976);
and UO_77 (O_77,N_2934,N_2931);
nand UO_78 (O_78,N_2910,N_2937);
nor UO_79 (O_79,N_2845,N_2810);
and UO_80 (O_80,N_2887,N_2827);
nor UO_81 (O_81,N_2868,N_2883);
nand UO_82 (O_82,N_2821,N_2875);
or UO_83 (O_83,N_2836,N_2935);
nand UO_84 (O_84,N_2973,N_2851);
nand UO_85 (O_85,N_2926,N_2981);
nor UO_86 (O_86,N_2916,N_2972);
or UO_87 (O_87,N_2856,N_2930);
nand UO_88 (O_88,N_2826,N_2914);
nand UO_89 (O_89,N_2802,N_2867);
or UO_90 (O_90,N_2912,N_2952);
nor UO_91 (O_91,N_2932,N_2872);
or UO_92 (O_92,N_2891,N_2855);
nand UO_93 (O_93,N_2893,N_2963);
or UO_94 (O_94,N_2938,N_2833);
nand UO_95 (O_95,N_2913,N_2966);
nand UO_96 (O_96,N_2982,N_2846);
and UO_97 (O_97,N_2995,N_2996);
nor UO_98 (O_98,N_2819,N_2844);
or UO_99 (O_99,N_2865,N_2871);
nand UO_100 (O_100,N_2949,N_2901);
or UO_101 (O_101,N_2958,N_2988);
or UO_102 (O_102,N_2986,N_2859);
nor UO_103 (O_103,N_2990,N_2812);
nor UO_104 (O_104,N_2835,N_2980);
nor UO_105 (O_105,N_2835,N_2964);
or UO_106 (O_106,N_2918,N_2846);
nand UO_107 (O_107,N_2913,N_2861);
nor UO_108 (O_108,N_2802,N_2889);
or UO_109 (O_109,N_2913,N_2953);
nor UO_110 (O_110,N_2988,N_2850);
or UO_111 (O_111,N_2879,N_2951);
and UO_112 (O_112,N_2821,N_2944);
nor UO_113 (O_113,N_2820,N_2989);
nor UO_114 (O_114,N_2883,N_2948);
nor UO_115 (O_115,N_2823,N_2871);
or UO_116 (O_116,N_2872,N_2861);
nor UO_117 (O_117,N_2928,N_2855);
nand UO_118 (O_118,N_2948,N_2854);
and UO_119 (O_119,N_2852,N_2802);
nor UO_120 (O_120,N_2862,N_2965);
nor UO_121 (O_121,N_2952,N_2908);
nor UO_122 (O_122,N_2909,N_2963);
nand UO_123 (O_123,N_2978,N_2808);
nand UO_124 (O_124,N_2826,N_2992);
nor UO_125 (O_125,N_2929,N_2863);
nand UO_126 (O_126,N_2833,N_2881);
and UO_127 (O_127,N_2856,N_2903);
and UO_128 (O_128,N_2887,N_2957);
nor UO_129 (O_129,N_2913,N_2898);
or UO_130 (O_130,N_2860,N_2973);
nor UO_131 (O_131,N_2890,N_2936);
and UO_132 (O_132,N_2947,N_2943);
nor UO_133 (O_133,N_2812,N_2814);
or UO_134 (O_134,N_2962,N_2991);
nand UO_135 (O_135,N_2908,N_2884);
and UO_136 (O_136,N_2862,N_2865);
or UO_137 (O_137,N_2843,N_2924);
and UO_138 (O_138,N_2976,N_2957);
nor UO_139 (O_139,N_2935,N_2972);
or UO_140 (O_140,N_2804,N_2883);
nand UO_141 (O_141,N_2957,N_2970);
nor UO_142 (O_142,N_2947,N_2852);
nor UO_143 (O_143,N_2910,N_2807);
and UO_144 (O_144,N_2840,N_2913);
xor UO_145 (O_145,N_2993,N_2954);
nand UO_146 (O_146,N_2922,N_2836);
nand UO_147 (O_147,N_2897,N_2852);
nand UO_148 (O_148,N_2831,N_2945);
and UO_149 (O_149,N_2824,N_2957);
nor UO_150 (O_150,N_2862,N_2974);
and UO_151 (O_151,N_2997,N_2809);
nor UO_152 (O_152,N_2898,N_2944);
and UO_153 (O_153,N_2918,N_2982);
and UO_154 (O_154,N_2947,N_2865);
nor UO_155 (O_155,N_2812,N_2931);
and UO_156 (O_156,N_2865,N_2967);
nor UO_157 (O_157,N_2994,N_2893);
nand UO_158 (O_158,N_2966,N_2801);
nor UO_159 (O_159,N_2952,N_2991);
nand UO_160 (O_160,N_2990,N_2970);
nor UO_161 (O_161,N_2961,N_2951);
or UO_162 (O_162,N_2941,N_2816);
nand UO_163 (O_163,N_2959,N_2859);
and UO_164 (O_164,N_2880,N_2948);
or UO_165 (O_165,N_2924,N_2955);
nor UO_166 (O_166,N_2932,N_2841);
nand UO_167 (O_167,N_2961,N_2914);
nand UO_168 (O_168,N_2925,N_2894);
or UO_169 (O_169,N_2855,N_2888);
or UO_170 (O_170,N_2978,N_2977);
nand UO_171 (O_171,N_2842,N_2803);
or UO_172 (O_172,N_2871,N_2904);
nand UO_173 (O_173,N_2961,N_2944);
nand UO_174 (O_174,N_2931,N_2964);
or UO_175 (O_175,N_2935,N_2881);
nand UO_176 (O_176,N_2868,N_2944);
or UO_177 (O_177,N_2913,N_2979);
nor UO_178 (O_178,N_2919,N_2853);
nor UO_179 (O_179,N_2968,N_2990);
or UO_180 (O_180,N_2830,N_2951);
and UO_181 (O_181,N_2918,N_2905);
and UO_182 (O_182,N_2832,N_2936);
nand UO_183 (O_183,N_2842,N_2967);
nor UO_184 (O_184,N_2980,N_2936);
and UO_185 (O_185,N_2823,N_2866);
or UO_186 (O_186,N_2833,N_2914);
nand UO_187 (O_187,N_2805,N_2932);
or UO_188 (O_188,N_2908,N_2955);
nand UO_189 (O_189,N_2813,N_2924);
and UO_190 (O_190,N_2914,N_2861);
nor UO_191 (O_191,N_2945,N_2867);
nor UO_192 (O_192,N_2818,N_2803);
and UO_193 (O_193,N_2995,N_2974);
or UO_194 (O_194,N_2989,N_2999);
or UO_195 (O_195,N_2851,N_2932);
nor UO_196 (O_196,N_2924,N_2916);
nand UO_197 (O_197,N_2993,N_2956);
nand UO_198 (O_198,N_2930,N_2825);
nand UO_199 (O_199,N_2830,N_2801);
nor UO_200 (O_200,N_2984,N_2828);
and UO_201 (O_201,N_2943,N_2998);
or UO_202 (O_202,N_2874,N_2983);
nor UO_203 (O_203,N_2819,N_2973);
or UO_204 (O_204,N_2881,N_2992);
nor UO_205 (O_205,N_2911,N_2886);
or UO_206 (O_206,N_2889,N_2983);
nor UO_207 (O_207,N_2917,N_2988);
nand UO_208 (O_208,N_2984,N_2883);
nand UO_209 (O_209,N_2815,N_2925);
and UO_210 (O_210,N_2907,N_2915);
nand UO_211 (O_211,N_2859,N_2833);
and UO_212 (O_212,N_2804,N_2999);
or UO_213 (O_213,N_2836,N_2862);
and UO_214 (O_214,N_2884,N_2810);
and UO_215 (O_215,N_2885,N_2899);
and UO_216 (O_216,N_2866,N_2919);
or UO_217 (O_217,N_2982,N_2849);
and UO_218 (O_218,N_2970,N_2853);
nor UO_219 (O_219,N_2908,N_2924);
or UO_220 (O_220,N_2950,N_2997);
or UO_221 (O_221,N_2926,N_2918);
nand UO_222 (O_222,N_2893,N_2938);
or UO_223 (O_223,N_2800,N_2928);
and UO_224 (O_224,N_2907,N_2885);
and UO_225 (O_225,N_2891,N_2961);
or UO_226 (O_226,N_2867,N_2808);
nand UO_227 (O_227,N_2920,N_2909);
nand UO_228 (O_228,N_2891,N_2818);
or UO_229 (O_229,N_2906,N_2976);
or UO_230 (O_230,N_2951,N_2859);
or UO_231 (O_231,N_2918,N_2959);
and UO_232 (O_232,N_2997,N_2957);
and UO_233 (O_233,N_2912,N_2989);
and UO_234 (O_234,N_2982,N_2977);
and UO_235 (O_235,N_2902,N_2894);
and UO_236 (O_236,N_2831,N_2921);
or UO_237 (O_237,N_2923,N_2986);
and UO_238 (O_238,N_2822,N_2831);
nor UO_239 (O_239,N_2953,N_2990);
or UO_240 (O_240,N_2927,N_2909);
xor UO_241 (O_241,N_2907,N_2891);
nand UO_242 (O_242,N_2822,N_2829);
and UO_243 (O_243,N_2923,N_2984);
nand UO_244 (O_244,N_2843,N_2871);
nor UO_245 (O_245,N_2869,N_2946);
nor UO_246 (O_246,N_2941,N_2815);
nor UO_247 (O_247,N_2892,N_2899);
nand UO_248 (O_248,N_2904,N_2837);
nor UO_249 (O_249,N_2986,N_2807);
and UO_250 (O_250,N_2806,N_2816);
nor UO_251 (O_251,N_2915,N_2871);
and UO_252 (O_252,N_2866,N_2977);
nand UO_253 (O_253,N_2848,N_2975);
nor UO_254 (O_254,N_2961,N_2962);
and UO_255 (O_255,N_2872,N_2835);
and UO_256 (O_256,N_2829,N_2811);
nand UO_257 (O_257,N_2949,N_2850);
or UO_258 (O_258,N_2877,N_2828);
nor UO_259 (O_259,N_2925,N_2828);
or UO_260 (O_260,N_2995,N_2837);
nand UO_261 (O_261,N_2988,N_2965);
xor UO_262 (O_262,N_2923,N_2842);
nand UO_263 (O_263,N_2832,N_2867);
and UO_264 (O_264,N_2989,N_2971);
nor UO_265 (O_265,N_2990,N_2823);
and UO_266 (O_266,N_2905,N_2855);
and UO_267 (O_267,N_2913,N_2946);
or UO_268 (O_268,N_2871,N_2807);
or UO_269 (O_269,N_2975,N_2969);
nand UO_270 (O_270,N_2900,N_2966);
nand UO_271 (O_271,N_2996,N_2856);
xnor UO_272 (O_272,N_2954,N_2834);
nand UO_273 (O_273,N_2800,N_2924);
or UO_274 (O_274,N_2800,N_2955);
xor UO_275 (O_275,N_2890,N_2868);
nor UO_276 (O_276,N_2836,N_2882);
and UO_277 (O_277,N_2972,N_2966);
or UO_278 (O_278,N_2915,N_2936);
and UO_279 (O_279,N_2879,N_2892);
nand UO_280 (O_280,N_2923,N_2908);
or UO_281 (O_281,N_2980,N_2996);
and UO_282 (O_282,N_2879,N_2812);
nor UO_283 (O_283,N_2811,N_2801);
nand UO_284 (O_284,N_2876,N_2989);
nand UO_285 (O_285,N_2980,N_2869);
or UO_286 (O_286,N_2846,N_2855);
and UO_287 (O_287,N_2892,N_2818);
or UO_288 (O_288,N_2924,N_2921);
and UO_289 (O_289,N_2838,N_2835);
and UO_290 (O_290,N_2811,N_2940);
and UO_291 (O_291,N_2869,N_2894);
and UO_292 (O_292,N_2899,N_2984);
nor UO_293 (O_293,N_2926,N_2942);
and UO_294 (O_294,N_2823,N_2880);
or UO_295 (O_295,N_2923,N_2901);
and UO_296 (O_296,N_2987,N_2854);
or UO_297 (O_297,N_2884,N_2988);
or UO_298 (O_298,N_2807,N_2947);
nor UO_299 (O_299,N_2967,N_2867);
nor UO_300 (O_300,N_2951,N_2904);
nor UO_301 (O_301,N_2994,N_2811);
nand UO_302 (O_302,N_2891,N_2987);
and UO_303 (O_303,N_2872,N_2976);
or UO_304 (O_304,N_2849,N_2934);
nand UO_305 (O_305,N_2981,N_2999);
and UO_306 (O_306,N_2924,N_2887);
or UO_307 (O_307,N_2862,N_2961);
or UO_308 (O_308,N_2860,N_2834);
and UO_309 (O_309,N_2868,N_2844);
or UO_310 (O_310,N_2931,N_2952);
nor UO_311 (O_311,N_2909,N_2839);
and UO_312 (O_312,N_2842,N_2909);
nor UO_313 (O_313,N_2962,N_2881);
xnor UO_314 (O_314,N_2953,N_2985);
nand UO_315 (O_315,N_2927,N_2843);
nand UO_316 (O_316,N_2834,N_2852);
nor UO_317 (O_317,N_2807,N_2893);
nor UO_318 (O_318,N_2892,N_2888);
and UO_319 (O_319,N_2913,N_2832);
nor UO_320 (O_320,N_2995,N_2981);
nand UO_321 (O_321,N_2926,N_2989);
nor UO_322 (O_322,N_2827,N_2853);
nand UO_323 (O_323,N_2997,N_2912);
nand UO_324 (O_324,N_2801,N_2847);
or UO_325 (O_325,N_2984,N_2909);
xnor UO_326 (O_326,N_2802,N_2925);
and UO_327 (O_327,N_2925,N_2941);
nor UO_328 (O_328,N_2952,N_2980);
nand UO_329 (O_329,N_2897,N_2857);
nand UO_330 (O_330,N_2990,N_2914);
nor UO_331 (O_331,N_2915,N_2934);
nor UO_332 (O_332,N_2860,N_2924);
or UO_333 (O_333,N_2937,N_2960);
and UO_334 (O_334,N_2969,N_2865);
or UO_335 (O_335,N_2839,N_2821);
nor UO_336 (O_336,N_2893,N_2915);
and UO_337 (O_337,N_2915,N_2802);
nand UO_338 (O_338,N_2805,N_2920);
nand UO_339 (O_339,N_2905,N_2994);
nor UO_340 (O_340,N_2932,N_2960);
nand UO_341 (O_341,N_2841,N_2970);
nor UO_342 (O_342,N_2928,N_2811);
nand UO_343 (O_343,N_2918,N_2969);
and UO_344 (O_344,N_2813,N_2800);
nand UO_345 (O_345,N_2913,N_2921);
nand UO_346 (O_346,N_2830,N_2931);
nor UO_347 (O_347,N_2995,N_2972);
nor UO_348 (O_348,N_2880,N_2885);
nor UO_349 (O_349,N_2980,N_2983);
or UO_350 (O_350,N_2993,N_2818);
or UO_351 (O_351,N_2817,N_2886);
nor UO_352 (O_352,N_2829,N_2856);
nand UO_353 (O_353,N_2967,N_2916);
nor UO_354 (O_354,N_2884,N_2900);
and UO_355 (O_355,N_2985,N_2814);
and UO_356 (O_356,N_2935,N_2888);
and UO_357 (O_357,N_2829,N_2974);
and UO_358 (O_358,N_2973,N_2919);
and UO_359 (O_359,N_2951,N_2988);
nand UO_360 (O_360,N_2891,N_2965);
and UO_361 (O_361,N_2898,N_2836);
or UO_362 (O_362,N_2874,N_2896);
nand UO_363 (O_363,N_2840,N_2996);
nor UO_364 (O_364,N_2947,N_2988);
or UO_365 (O_365,N_2838,N_2923);
or UO_366 (O_366,N_2935,N_2856);
and UO_367 (O_367,N_2928,N_2979);
and UO_368 (O_368,N_2983,N_2804);
nand UO_369 (O_369,N_2875,N_2866);
nand UO_370 (O_370,N_2968,N_2983);
and UO_371 (O_371,N_2901,N_2889);
or UO_372 (O_372,N_2929,N_2886);
nand UO_373 (O_373,N_2860,N_2918);
or UO_374 (O_374,N_2914,N_2857);
or UO_375 (O_375,N_2869,N_2809);
xor UO_376 (O_376,N_2967,N_2832);
nand UO_377 (O_377,N_2979,N_2867);
nand UO_378 (O_378,N_2937,N_2906);
nand UO_379 (O_379,N_2853,N_2938);
or UO_380 (O_380,N_2995,N_2889);
and UO_381 (O_381,N_2989,N_2958);
nor UO_382 (O_382,N_2842,N_2802);
nor UO_383 (O_383,N_2933,N_2975);
or UO_384 (O_384,N_2929,N_2874);
nor UO_385 (O_385,N_2858,N_2950);
nand UO_386 (O_386,N_2934,N_2988);
and UO_387 (O_387,N_2973,N_2839);
nand UO_388 (O_388,N_2956,N_2897);
nand UO_389 (O_389,N_2848,N_2958);
and UO_390 (O_390,N_2949,N_2964);
nand UO_391 (O_391,N_2968,N_2882);
and UO_392 (O_392,N_2958,N_2851);
or UO_393 (O_393,N_2987,N_2911);
nand UO_394 (O_394,N_2866,N_2931);
and UO_395 (O_395,N_2850,N_2955);
nand UO_396 (O_396,N_2870,N_2856);
xor UO_397 (O_397,N_2995,N_2973);
nand UO_398 (O_398,N_2868,N_2931);
nor UO_399 (O_399,N_2887,N_2938);
and UO_400 (O_400,N_2954,N_2959);
nand UO_401 (O_401,N_2952,N_2929);
nor UO_402 (O_402,N_2859,N_2974);
nand UO_403 (O_403,N_2996,N_2849);
or UO_404 (O_404,N_2865,N_2852);
nor UO_405 (O_405,N_2840,N_2832);
nor UO_406 (O_406,N_2989,N_2963);
and UO_407 (O_407,N_2905,N_2947);
or UO_408 (O_408,N_2879,N_2883);
nor UO_409 (O_409,N_2818,N_2922);
or UO_410 (O_410,N_2993,N_2907);
and UO_411 (O_411,N_2910,N_2800);
and UO_412 (O_412,N_2902,N_2977);
or UO_413 (O_413,N_2971,N_2980);
and UO_414 (O_414,N_2980,N_2864);
nor UO_415 (O_415,N_2963,N_2855);
and UO_416 (O_416,N_2807,N_2946);
nor UO_417 (O_417,N_2846,N_2896);
nor UO_418 (O_418,N_2951,N_2851);
or UO_419 (O_419,N_2833,N_2977);
nand UO_420 (O_420,N_2874,N_2883);
nor UO_421 (O_421,N_2950,N_2899);
or UO_422 (O_422,N_2817,N_2831);
and UO_423 (O_423,N_2981,N_2858);
nand UO_424 (O_424,N_2872,N_2842);
or UO_425 (O_425,N_2948,N_2946);
nor UO_426 (O_426,N_2845,N_2899);
and UO_427 (O_427,N_2896,N_2908);
nor UO_428 (O_428,N_2807,N_2972);
nor UO_429 (O_429,N_2849,N_2882);
nor UO_430 (O_430,N_2966,N_2948);
nor UO_431 (O_431,N_2931,N_2995);
or UO_432 (O_432,N_2985,N_2878);
nand UO_433 (O_433,N_2848,N_2917);
nand UO_434 (O_434,N_2929,N_2855);
nor UO_435 (O_435,N_2955,N_2813);
nand UO_436 (O_436,N_2881,N_2974);
or UO_437 (O_437,N_2819,N_2825);
nand UO_438 (O_438,N_2940,N_2819);
and UO_439 (O_439,N_2868,N_2871);
and UO_440 (O_440,N_2977,N_2868);
and UO_441 (O_441,N_2957,N_2854);
nor UO_442 (O_442,N_2835,N_2857);
nand UO_443 (O_443,N_2878,N_2830);
nor UO_444 (O_444,N_2948,N_2974);
and UO_445 (O_445,N_2947,N_2870);
and UO_446 (O_446,N_2980,N_2949);
or UO_447 (O_447,N_2954,N_2836);
xnor UO_448 (O_448,N_2824,N_2872);
nand UO_449 (O_449,N_2885,N_2812);
or UO_450 (O_450,N_2969,N_2843);
or UO_451 (O_451,N_2913,N_2887);
and UO_452 (O_452,N_2944,N_2900);
nor UO_453 (O_453,N_2983,N_2956);
nand UO_454 (O_454,N_2829,N_2996);
nor UO_455 (O_455,N_2976,N_2855);
or UO_456 (O_456,N_2850,N_2802);
and UO_457 (O_457,N_2845,N_2806);
and UO_458 (O_458,N_2916,N_2813);
and UO_459 (O_459,N_2817,N_2844);
xor UO_460 (O_460,N_2962,N_2966);
nand UO_461 (O_461,N_2904,N_2984);
nand UO_462 (O_462,N_2922,N_2961);
or UO_463 (O_463,N_2959,N_2938);
nand UO_464 (O_464,N_2941,N_2866);
nor UO_465 (O_465,N_2826,N_2996);
or UO_466 (O_466,N_2829,N_2834);
and UO_467 (O_467,N_2823,N_2842);
and UO_468 (O_468,N_2889,N_2942);
nand UO_469 (O_469,N_2970,N_2892);
or UO_470 (O_470,N_2870,N_2932);
nor UO_471 (O_471,N_2892,N_2827);
or UO_472 (O_472,N_2925,N_2997);
nor UO_473 (O_473,N_2954,N_2869);
nand UO_474 (O_474,N_2956,N_2886);
nand UO_475 (O_475,N_2949,N_2968);
and UO_476 (O_476,N_2863,N_2887);
nand UO_477 (O_477,N_2895,N_2983);
nor UO_478 (O_478,N_2866,N_2967);
nor UO_479 (O_479,N_2965,N_2858);
nor UO_480 (O_480,N_2809,N_2867);
nand UO_481 (O_481,N_2811,N_2969);
nand UO_482 (O_482,N_2812,N_2960);
nor UO_483 (O_483,N_2848,N_2810);
nand UO_484 (O_484,N_2828,N_2953);
nand UO_485 (O_485,N_2894,N_2937);
nand UO_486 (O_486,N_2803,N_2921);
nand UO_487 (O_487,N_2963,N_2980);
and UO_488 (O_488,N_2970,N_2924);
nor UO_489 (O_489,N_2869,N_2961);
or UO_490 (O_490,N_2923,N_2803);
nand UO_491 (O_491,N_2999,N_2859);
and UO_492 (O_492,N_2873,N_2891);
nor UO_493 (O_493,N_2969,N_2999);
or UO_494 (O_494,N_2850,N_2911);
nor UO_495 (O_495,N_2851,N_2916);
nor UO_496 (O_496,N_2961,N_2968);
and UO_497 (O_497,N_2906,N_2815);
or UO_498 (O_498,N_2812,N_2847);
nor UO_499 (O_499,N_2934,N_2838);
endmodule