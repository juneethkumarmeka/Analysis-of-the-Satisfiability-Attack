module basic_500_3000_500_3_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_130,In_235);
and U1 (N_1,In_73,In_282);
or U2 (N_2,In_102,In_90);
or U3 (N_3,In_295,In_214);
nand U4 (N_4,In_459,In_298);
and U5 (N_5,In_338,In_225);
nand U6 (N_6,In_45,In_211);
nand U7 (N_7,In_131,In_482);
xnor U8 (N_8,In_244,In_422);
nand U9 (N_9,In_291,In_96);
or U10 (N_10,In_387,In_92);
nor U11 (N_11,In_265,In_187);
xnor U12 (N_12,In_401,In_234);
nor U13 (N_13,In_439,In_485);
xor U14 (N_14,In_409,In_432);
or U15 (N_15,In_243,In_88);
xnor U16 (N_16,In_224,In_495);
nor U17 (N_17,In_192,In_287);
and U18 (N_18,In_109,In_332);
xnor U19 (N_19,In_402,In_184);
nand U20 (N_20,In_271,In_430);
and U21 (N_21,In_273,In_348);
or U22 (N_22,In_388,In_356);
or U23 (N_23,In_286,In_391);
nand U24 (N_24,In_174,In_336);
nor U25 (N_25,In_108,In_204);
or U26 (N_26,In_160,In_418);
nor U27 (N_27,In_322,In_479);
nand U28 (N_28,In_170,In_355);
or U29 (N_29,In_285,In_70);
xor U30 (N_30,In_110,In_35);
and U31 (N_31,In_360,In_315);
or U32 (N_32,In_444,In_30);
nor U33 (N_33,In_80,In_167);
nand U34 (N_34,In_379,In_331);
or U35 (N_35,In_257,In_199);
xnor U36 (N_36,In_325,In_384);
or U37 (N_37,In_458,In_239);
nor U38 (N_38,In_343,In_254);
and U39 (N_39,In_324,In_292);
xnor U40 (N_40,In_116,In_38);
or U41 (N_41,In_437,In_252);
xor U42 (N_42,In_84,In_213);
and U43 (N_43,In_326,In_156);
and U44 (N_44,In_133,In_173);
or U45 (N_45,In_269,In_64);
nand U46 (N_46,In_469,In_375);
or U47 (N_47,In_405,In_0);
nand U48 (N_48,In_127,In_321);
nand U49 (N_49,In_306,In_3);
nand U50 (N_50,In_44,In_395);
and U51 (N_51,In_498,In_447);
nor U52 (N_52,In_303,In_163);
nand U53 (N_53,In_320,In_307);
nor U54 (N_54,In_374,In_144);
xor U55 (N_55,In_312,In_202);
nor U56 (N_56,In_435,In_261);
or U57 (N_57,In_29,In_123);
or U58 (N_58,In_350,In_208);
or U59 (N_59,In_408,In_4);
nand U60 (N_60,In_323,In_82);
or U61 (N_61,In_12,In_54);
and U62 (N_62,In_440,In_475);
or U63 (N_63,In_129,In_275);
nor U64 (N_64,In_474,In_63);
and U65 (N_65,In_397,In_329);
and U66 (N_66,In_7,In_240);
nor U67 (N_67,In_251,In_223);
and U68 (N_68,In_14,In_450);
xnor U69 (N_69,In_87,In_67);
or U70 (N_70,In_487,In_490);
nand U71 (N_71,In_13,In_162);
nand U72 (N_72,In_26,In_317);
xnor U73 (N_73,In_491,In_246);
nor U74 (N_74,In_148,In_158);
and U75 (N_75,In_238,In_346);
xor U76 (N_76,In_42,In_341);
nand U77 (N_77,In_171,In_277);
or U78 (N_78,In_86,In_168);
or U79 (N_79,In_369,In_107);
nor U80 (N_80,In_334,In_480);
and U81 (N_81,In_441,In_476);
or U82 (N_82,In_159,In_194);
nand U83 (N_83,In_274,In_125);
nor U84 (N_84,In_191,In_182);
xnor U85 (N_85,In_433,In_231);
nor U86 (N_86,In_169,In_18);
and U87 (N_87,In_53,In_386);
and U88 (N_88,In_382,In_345);
nor U89 (N_89,In_373,In_161);
nand U90 (N_90,In_114,In_446);
nand U91 (N_91,In_151,In_406);
or U92 (N_92,In_327,In_41);
and U93 (N_93,In_81,In_197);
or U94 (N_94,In_481,In_358);
nor U95 (N_95,In_85,In_328);
and U96 (N_96,In_380,In_172);
or U97 (N_97,In_147,In_46);
and U98 (N_98,In_478,In_203);
or U99 (N_99,In_443,In_362);
nand U100 (N_100,In_270,In_392);
nor U101 (N_101,In_75,In_242);
or U102 (N_102,In_453,In_178);
nand U103 (N_103,In_492,In_118);
nand U104 (N_104,In_353,In_72);
or U105 (N_105,In_417,In_48);
and U106 (N_106,In_473,In_318);
xor U107 (N_107,In_483,In_296);
or U108 (N_108,In_219,In_359);
and U109 (N_109,In_175,In_177);
or U110 (N_110,In_421,In_372);
xnor U111 (N_111,In_149,In_209);
nand U112 (N_112,In_23,In_137);
xnor U113 (N_113,In_484,In_337);
xnor U114 (N_114,In_28,In_61);
xor U115 (N_115,In_55,In_122);
nand U116 (N_116,In_233,In_313);
nand U117 (N_117,In_364,In_342);
nand U118 (N_118,In_25,In_494);
nand U119 (N_119,In_39,In_393);
and U120 (N_120,In_419,In_196);
or U121 (N_121,In_370,In_180);
nand U122 (N_122,In_247,In_352);
and U123 (N_123,In_100,In_221);
or U124 (N_124,In_267,In_457);
nor U125 (N_125,In_136,In_50);
nor U126 (N_126,In_205,In_215);
xnor U127 (N_127,In_24,In_377);
and U128 (N_128,In_354,In_52);
xor U129 (N_129,In_10,In_499);
nand U130 (N_130,In_367,In_216);
nor U131 (N_131,In_207,In_34);
and U132 (N_132,In_264,In_58);
nor U133 (N_133,In_294,In_27);
and U134 (N_134,In_124,In_276);
xor U135 (N_135,In_427,In_464);
and U136 (N_136,In_389,In_165);
or U137 (N_137,In_310,In_99);
and U138 (N_138,In_293,In_466);
xor U139 (N_139,In_414,In_228);
and U140 (N_140,In_220,In_89);
xor U141 (N_141,In_206,In_143);
nor U142 (N_142,In_410,In_248);
nand U143 (N_143,In_95,In_141);
and U144 (N_144,In_227,In_438);
and U145 (N_145,In_40,In_376);
nor U146 (N_146,In_451,In_188);
nand U147 (N_147,In_49,In_19);
and U148 (N_148,In_31,In_65);
nand U149 (N_149,In_339,In_425);
nor U150 (N_150,In_43,In_150);
or U151 (N_151,In_268,In_305);
or U152 (N_152,In_493,In_288);
and U153 (N_153,In_456,In_302);
xor U154 (N_154,In_212,In_497);
xnor U155 (N_155,In_138,In_93);
nand U156 (N_156,In_454,In_426);
nor U157 (N_157,In_195,In_279);
and U158 (N_158,In_299,In_83);
and U159 (N_159,In_62,In_128);
xor U160 (N_160,In_185,In_423);
xor U161 (N_161,In_20,In_200);
and U162 (N_162,In_60,In_78);
and U163 (N_163,In_399,In_452);
nor U164 (N_164,In_403,In_304);
xnor U165 (N_165,In_218,In_390);
xnor U166 (N_166,In_361,In_1);
or U167 (N_167,In_420,In_5);
xnor U168 (N_168,In_462,In_460);
or U169 (N_169,In_153,In_449);
nor U170 (N_170,In_98,In_436);
and U171 (N_171,In_398,In_121);
nand U172 (N_172,In_236,In_489);
nand U173 (N_173,In_237,In_349);
xnor U174 (N_174,In_37,In_146);
and U175 (N_175,In_434,In_135);
and U176 (N_176,In_465,In_112);
and U177 (N_177,In_266,In_139);
nand U178 (N_178,In_66,In_263);
xnor U179 (N_179,In_278,In_32);
nor U180 (N_180,In_229,In_486);
nor U181 (N_181,In_6,In_431);
xnor U182 (N_182,In_258,In_404);
or U183 (N_183,In_76,In_2);
nand U184 (N_184,In_415,In_210);
or U185 (N_185,In_250,In_120);
xor U186 (N_186,In_142,In_488);
nand U187 (N_187,In_428,In_259);
or U188 (N_188,In_11,In_22);
nand U189 (N_189,In_94,In_16);
and U190 (N_190,In_407,In_115);
xor U191 (N_191,In_308,In_105);
nor U192 (N_192,In_314,In_157);
and U193 (N_193,In_181,In_59);
nor U194 (N_194,In_412,In_117);
nand U195 (N_195,In_145,In_383);
nand U196 (N_196,In_301,In_289);
and U197 (N_197,In_179,In_132);
nor U198 (N_198,In_189,In_249);
nor U199 (N_199,In_47,In_253);
nand U200 (N_200,In_79,In_186);
or U201 (N_201,In_56,In_477);
or U202 (N_202,In_15,In_330);
and U203 (N_203,In_119,In_344);
nand U204 (N_204,In_222,In_103);
xor U205 (N_205,In_385,In_413);
nor U206 (N_206,In_400,In_69);
and U207 (N_207,In_33,In_232);
nand U208 (N_208,In_429,In_68);
nor U209 (N_209,In_316,In_378);
and U210 (N_210,In_176,In_290);
and U211 (N_211,In_363,In_17);
or U212 (N_212,In_351,In_198);
xor U213 (N_213,In_262,In_340);
nand U214 (N_214,In_455,In_461);
xor U215 (N_215,In_272,In_51);
or U216 (N_216,In_471,In_333);
and U217 (N_217,In_77,In_366);
xnor U218 (N_218,In_97,In_335);
or U219 (N_219,In_371,In_166);
nor U220 (N_220,In_468,In_113);
nor U221 (N_221,In_463,In_496);
and U222 (N_222,In_297,In_183);
and U223 (N_223,In_36,In_190);
xnor U224 (N_224,In_365,In_245);
or U225 (N_225,In_284,In_106);
nand U226 (N_226,In_319,In_300);
or U227 (N_227,In_260,In_256);
nor U228 (N_228,In_57,In_126);
or U229 (N_229,In_8,In_416);
and U230 (N_230,In_74,In_201);
nor U231 (N_231,In_396,In_217);
nand U232 (N_232,In_155,In_472);
nand U233 (N_233,In_309,In_281);
nor U234 (N_234,In_467,In_470);
nand U235 (N_235,In_283,In_134);
and U236 (N_236,In_140,In_91);
xor U237 (N_237,In_104,In_164);
nor U238 (N_238,In_71,In_381);
nor U239 (N_239,In_230,In_154);
nor U240 (N_240,In_357,In_255);
nand U241 (N_241,In_442,In_101);
and U242 (N_242,In_21,In_241);
nor U243 (N_243,In_152,In_448);
nand U244 (N_244,In_111,In_347);
nor U245 (N_245,In_280,In_193);
and U246 (N_246,In_445,In_368);
nor U247 (N_247,In_226,In_424);
and U248 (N_248,In_9,In_311);
xnor U249 (N_249,In_394,In_411);
nand U250 (N_250,In_101,In_238);
nor U251 (N_251,In_74,In_132);
and U252 (N_252,In_405,In_486);
and U253 (N_253,In_441,In_239);
and U254 (N_254,In_402,In_93);
and U255 (N_255,In_399,In_477);
or U256 (N_256,In_49,In_484);
nor U257 (N_257,In_159,In_7);
xor U258 (N_258,In_60,In_345);
nor U259 (N_259,In_151,In_100);
nand U260 (N_260,In_416,In_488);
nor U261 (N_261,In_96,In_238);
and U262 (N_262,In_490,In_302);
nand U263 (N_263,In_32,In_151);
and U264 (N_264,In_262,In_469);
nand U265 (N_265,In_166,In_375);
and U266 (N_266,In_279,In_125);
nand U267 (N_267,In_367,In_407);
or U268 (N_268,In_449,In_300);
nor U269 (N_269,In_214,In_291);
or U270 (N_270,In_174,In_366);
nand U271 (N_271,In_466,In_165);
xnor U272 (N_272,In_32,In_210);
nand U273 (N_273,In_53,In_364);
nor U274 (N_274,In_184,In_98);
nand U275 (N_275,In_448,In_262);
and U276 (N_276,In_297,In_282);
and U277 (N_277,In_409,In_147);
nand U278 (N_278,In_317,In_158);
and U279 (N_279,In_159,In_203);
or U280 (N_280,In_286,In_204);
nand U281 (N_281,In_380,In_325);
nand U282 (N_282,In_62,In_104);
nor U283 (N_283,In_117,In_253);
xor U284 (N_284,In_95,In_330);
nor U285 (N_285,In_189,In_15);
nand U286 (N_286,In_149,In_82);
nor U287 (N_287,In_172,In_418);
and U288 (N_288,In_382,In_434);
and U289 (N_289,In_455,In_442);
nor U290 (N_290,In_124,In_190);
nand U291 (N_291,In_69,In_50);
or U292 (N_292,In_455,In_127);
xnor U293 (N_293,In_168,In_403);
xor U294 (N_294,In_394,In_36);
or U295 (N_295,In_312,In_384);
xnor U296 (N_296,In_498,In_257);
and U297 (N_297,In_259,In_3);
nand U298 (N_298,In_163,In_266);
and U299 (N_299,In_491,In_284);
or U300 (N_300,In_327,In_61);
or U301 (N_301,In_449,In_18);
xor U302 (N_302,In_407,In_209);
or U303 (N_303,In_339,In_199);
xor U304 (N_304,In_497,In_286);
nand U305 (N_305,In_203,In_443);
nor U306 (N_306,In_406,In_18);
and U307 (N_307,In_428,In_218);
nand U308 (N_308,In_95,In_231);
or U309 (N_309,In_184,In_486);
xnor U310 (N_310,In_204,In_303);
and U311 (N_311,In_35,In_77);
xnor U312 (N_312,In_133,In_415);
nand U313 (N_313,In_319,In_117);
nand U314 (N_314,In_113,In_449);
nand U315 (N_315,In_497,In_477);
and U316 (N_316,In_85,In_468);
or U317 (N_317,In_40,In_11);
nor U318 (N_318,In_252,In_269);
nand U319 (N_319,In_342,In_207);
and U320 (N_320,In_216,In_412);
or U321 (N_321,In_457,In_20);
nand U322 (N_322,In_192,In_69);
and U323 (N_323,In_361,In_73);
and U324 (N_324,In_92,In_398);
xnor U325 (N_325,In_87,In_84);
and U326 (N_326,In_197,In_123);
and U327 (N_327,In_386,In_37);
and U328 (N_328,In_72,In_435);
nor U329 (N_329,In_374,In_222);
or U330 (N_330,In_132,In_249);
and U331 (N_331,In_299,In_351);
xnor U332 (N_332,In_1,In_244);
nor U333 (N_333,In_343,In_33);
xnor U334 (N_334,In_46,In_366);
and U335 (N_335,In_298,In_151);
and U336 (N_336,In_338,In_494);
and U337 (N_337,In_189,In_113);
nor U338 (N_338,In_332,In_414);
or U339 (N_339,In_195,In_369);
nor U340 (N_340,In_218,In_379);
nor U341 (N_341,In_153,In_51);
nand U342 (N_342,In_63,In_75);
nand U343 (N_343,In_295,In_3);
nand U344 (N_344,In_86,In_354);
nand U345 (N_345,In_177,In_429);
nand U346 (N_346,In_81,In_168);
and U347 (N_347,In_73,In_304);
or U348 (N_348,In_28,In_225);
nand U349 (N_349,In_440,In_106);
nor U350 (N_350,In_82,In_255);
or U351 (N_351,In_398,In_195);
or U352 (N_352,In_413,In_199);
nand U353 (N_353,In_450,In_306);
and U354 (N_354,In_30,In_298);
and U355 (N_355,In_219,In_142);
nor U356 (N_356,In_463,In_14);
nand U357 (N_357,In_155,In_56);
or U358 (N_358,In_293,In_156);
and U359 (N_359,In_385,In_495);
nand U360 (N_360,In_367,In_217);
nand U361 (N_361,In_357,In_150);
nor U362 (N_362,In_408,In_261);
and U363 (N_363,In_117,In_234);
or U364 (N_364,In_168,In_315);
or U365 (N_365,In_108,In_177);
and U366 (N_366,In_181,In_326);
and U367 (N_367,In_183,In_431);
and U368 (N_368,In_264,In_237);
or U369 (N_369,In_188,In_132);
and U370 (N_370,In_31,In_121);
nor U371 (N_371,In_310,In_153);
or U372 (N_372,In_341,In_356);
xnor U373 (N_373,In_106,In_444);
nor U374 (N_374,In_321,In_302);
or U375 (N_375,In_48,In_253);
or U376 (N_376,In_302,In_217);
xnor U377 (N_377,In_313,In_484);
and U378 (N_378,In_68,In_260);
or U379 (N_379,In_24,In_264);
nor U380 (N_380,In_298,In_446);
nand U381 (N_381,In_353,In_110);
and U382 (N_382,In_131,In_484);
and U383 (N_383,In_31,In_423);
xnor U384 (N_384,In_176,In_213);
nor U385 (N_385,In_417,In_391);
nand U386 (N_386,In_409,In_350);
or U387 (N_387,In_330,In_460);
xnor U388 (N_388,In_345,In_222);
or U389 (N_389,In_495,In_98);
nor U390 (N_390,In_166,In_20);
nand U391 (N_391,In_260,In_405);
or U392 (N_392,In_126,In_80);
nand U393 (N_393,In_136,In_445);
xor U394 (N_394,In_213,In_140);
and U395 (N_395,In_368,In_161);
xor U396 (N_396,In_464,In_127);
nand U397 (N_397,In_163,In_213);
xnor U398 (N_398,In_118,In_25);
and U399 (N_399,In_467,In_211);
and U400 (N_400,In_360,In_185);
nand U401 (N_401,In_204,In_222);
or U402 (N_402,In_453,In_368);
or U403 (N_403,In_112,In_199);
nand U404 (N_404,In_75,In_398);
or U405 (N_405,In_310,In_98);
nand U406 (N_406,In_223,In_399);
nand U407 (N_407,In_57,In_449);
and U408 (N_408,In_184,In_298);
nand U409 (N_409,In_288,In_279);
nor U410 (N_410,In_304,In_18);
or U411 (N_411,In_334,In_287);
xor U412 (N_412,In_382,In_432);
nand U413 (N_413,In_326,In_216);
xnor U414 (N_414,In_226,In_314);
xnor U415 (N_415,In_490,In_337);
xnor U416 (N_416,In_368,In_472);
nand U417 (N_417,In_41,In_246);
xor U418 (N_418,In_8,In_92);
nand U419 (N_419,In_264,In_280);
xnor U420 (N_420,In_3,In_224);
and U421 (N_421,In_370,In_157);
and U422 (N_422,In_91,In_46);
or U423 (N_423,In_211,In_76);
or U424 (N_424,In_101,In_262);
nor U425 (N_425,In_104,In_141);
nor U426 (N_426,In_275,In_416);
nand U427 (N_427,In_30,In_100);
nand U428 (N_428,In_314,In_204);
or U429 (N_429,In_373,In_360);
and U430 (N_430,In_138,In_19);
or U431 (N_431,In_422,In_25);
or U432 (N_432,In_8,In_37);
and U433 (N_433,In_393,In_132);
and U434 (N_434,In_68,In_170);
and U435 (N_435,In_210,In_405);
xnor U436 (N_436,In_297,In_352);
nand U437 (N_437,In_392,In_195);
xnor U438 (N_438,In_55,In_481);
nor U439 (N_439,In_362,In_95);
and U440 (N_440,In_412,In_30);
or U441 (N_441,In_296,In_412);
nand U442 (N_442,In_37,In_15);
nor U443 (N_443,In_499,In_274);
or U444 (N_444,In_276,In_280);
nor U445 (N_445,In_35,In_157);
nor U446 (N_446,In_80,In_14);
and U447 (N_447,In_28,In_489);
nand U448 (N_448,In_170,In_384);
nor U449 (N_449,In_144,In_355);
nor U450 (N_450,In_323,In_55);
nand U451 (N_451,In_305,In_455);
xor U452 (N_452,In_242,In_450);
or U453 (N_453,In_118,In_137);
and U454 (N_454,In_22,In_307);
nor U455 (N_455,In_473,In_222);
and U456 (N_456,In_92,In_215);
and U457 (N_457,In_207,In_172);
xnor U458 (N_458,In_44,In_271);
and U459 (N_459,In_338,In_196);
nor U460 (N_460,In_300,In_480);
nor U461 (N_461,In_249,In_459);
nor U462 (N_462,In_326,In_360);
or U463 (N_463,In_276,In_495);
nor U464 (N_464,In_373,In_419);
nor U465 (N_465,In_29,In_409);
nor U466 (N_466,In_430,In_268);
nor U467 (N_467,In_120,In_399);
xnor U468 (N_468,In_486,In_493);
or U469 (N_469,In_36,In_38);
xnor U470 (N_470,In_343,In_22);
and U471 (N_471,In_155,In_43);
and U472 (N_472,In_137,In_452);
nand U473 (N_473,In_453,In_20);
or U474 (N_474,In_317,In_56);
and U475 (N_475,In_236,In_188);
or U476 (N_476,In_54,In_361);
and U477 (N_477,In_305,In_483);
and U478 (N_478,In_319,In_246);
or U479 (N_479,In_425,In_46);
xnor U480 (N_480,In_494,In_325);
xnor U481 (N_481,In_246,In_181);
xor U482 (N_482,In_198,In_82);
xor U483 (N_483,In_336,In_398);
nor U484 (N_484,In_105,In_60);
xnor U485 (N_485,In_404,In_440);
and U486 (N_486,In_395,In_376);
nor U487 (N_487,In_271,In_157);
or U488 (N_488,In_144,In_470);
or U489 (N_489,In_46,In_159);
and U490 (N_490,In_487,In_297);
and U491 (N_491,In_306,In_369);
and U492 (N_492,In_401,In_450);
nand U493 (N_493,In_436,In_388);
and U494 (N_494,In_37,In_84);
nand U495 (N_495,In_132,In_190);
or U496 (N_496,In_275,In_282);
or U497 (N_497,In_405,In_271);
nor U498 (N_498,In_199,In_337);
and U499 (N_499,In_157,In_158);
xor U500 (N_500,In_470,In_185);
xor U501 (N_501,In_36,In_423);
or U502 (N_502,In_254,In_92);
and U503 (N_503,In_337,In_405);
and U504 (N_504,In_29,In_249);
nor U505 (N_505,In_373,In_6);
xnor U506 (N_506,In_72,In_398);
or U507 (N_507,In_100,In_38);
nand U508 (N_508,In_176,In_308);
and U509 (N_509,In_101,In_53);
xor U510 (N_510,In_297,In_467);
and U511 (N_511,In_459,In_433);
nor U512 (N_512,In_184,In_137);
or U513 (N_513,In_439,In_31);
xor U514 (N_514,In_262,In_418);
and U515 (N_515,In_444,In_19);
nand U516 (N_516,In_490,In_232);
nor U517 (N_517,In_406,In_263);
or U518 (N_518,In_418,In_289);
nand U519 (N_519,In_62,In_472);
or U520 (N_520,In_266,In_246);
or U521 (N_521,In_179,In_456);
xor U522 (N_522,In_351,In_35);
nand U523 (N_523,In_461,In_18);
or U524 (N_524,In_246,In_29);
nor U525 (N_525,In_102,In_230);
and U526 (N_526,In_348,In_319);
or U527 (N_527,In_12,In_268);
and U528 (N_528,In_78,In_244);
or U529 (N_529,In_435,In_339);
or U530 (N_530,In_162,In_448);
and U531 (N_531,In_15,In_461);
nand U532 (N_532,In_304,In_433);
and U533 (N_533,In_209,In_368);
and U534 (N_534,In_331,In_396);
nor U535 (N_535,In_425,In_460);
and U536 (N_536,In_265,In_353);
xor U537 (N_537,In_303,In_175);
xor U538 (N_538,In_13,In_452);
nand U539 (N_539,In_300,In_409);
nor U540 (N_540,In_281,In_326);
or U541 (N_541,In_441,In_112);
or U542 (N_542,In_25,In_165);
nand U543 (N_543,In_391,In_366);
nor U544 (N_544,In_380,In_476);
xor U545 (N_545,In_122,In_77);
nand U546 (N_546,In_302,In_98);
or U547 (N_547,In_447,In_469);
xor U548 (N_548,In_348,In_340);
nand U549 (N_549,In_154,In_255);
xnor U550 (N_550,In_157,In_221);
and U551 (N_551,In_357,In_395);
xnor U552 (N_552,In_98,In_63);
xnor U553 (N_553,In_9,In_102);
and U554 (N_554,In_492,In_419);
xnor U555 (N_555,In_217,In_160);
and U556 (N_556,In_316,In_55);
xnor U557 (N_557,In_103,In_96);
nand U558 (N_558,In_382,In_151);
nor U559 (N_559,In_152,In_73);
and U560 (N_560,In_412,In_385);
xor U561 (N_561,In_428,In_416);
nand U562 (N_562,In_447,In_9);
nor U563 (N_563,In_232,In_492);
nand U564 (N_564,In_133,In_66);
nand U565 (N_565,In_105,In_276);
nor U566 (N_566,In_64,In_480);
and U567 (N_567,In_305,In_157);
nand U568 (N_568,In_65,In_258);
nand U569 (N_569,In_78,In_292);
and U570 (N_570,In_465,In_210);
xnor U571 (N_571,In_61,In_94);
and U572 (N_572,In_5,In_111);
or U573 (N_573,In_11,In_19);
nor U574 (N_574,In_286,In_386);
xor U575 (N_575,In_413,In_113);
and U576 (N_576,In_489,In_135);
nor U577 (N_577,In_258,In_199);
nand U578 (N_578,In_16,In_71);
xor U579 (N_579,In_383,In_306);
nor U580 (N_580,In_291,In_11);
xnor U581 (N_581,In_79,In_34);
nor U582 (N_582,In_337,In_25);
nor U583 (N_583,In_472,In_239);
and U584 (N_584,In_164,In_335);
and U585 (N_585,In_332,In_301);
xnor U586 (N_586,In_181,In_438);
nor U587 (N_587,In_51,In_439);
xnor U588 (N_588,In_179,In_200);
nand U589 (N_589,In_5,In_235);
or U590 (N_590,In_18,In_215);
and U591 (N_591,In_120,In_148);
or U592 (N_592,In_345,In_24);
or U593 (N_593,In_387,In_214);
and U594 (N_594,In_145,In_316);
or U595 (N_595,In_441,In_256);
nand U596 (N_596,In_291,In_429);
xor U597 (N_597,In_434,In_431);
xnor U598 (N_598,In_38,In_91);
or U599 (N_599,In_291,In_285);
xnor U600 (N_600,In_492,In_356);
and U601 (N_601,In_9,In_306);
xnor U602 (N_602,In_101,In_20);
nand U603 (N_603,In_386,In_5);
or U604 (N_604,In_28,In_247);
nand U605 (N_605,In_213,In_272);
xnor U606 (N_606,In_425,In_458);
nor U607 (N_607,In_163,In_496);
or U608 (N_608,In_135,In_44);
and U609 (N_609,In_257,In_302);
nand U610 (N_610,In_403,In_115);
or U611 (N_611,In_328,In_337);
or U612 (N_612,In_161,In_359);
and U613 (N_613,In_206,In_207);
nand U614 (N_614,In_3,In_314);
and U615 (N_615,In_290,In_18);
nand U616 (N_616,In_103,In_139);
xor U617 (N_617,In_125,In_183);
xor U618 (N_618,In_122,In_85);
nor U619 (N_619,In_306,In_314);
xor U620 (N_620,In_269,In_47);
nand U621 (N_621,In_463,In_447);
nor U622 (N_622,In_395,In_210);
xnor U623 (N_623,In_378,In_356);
nand U624 (N_624,In_149,In_74);
and U625 (N_625,In_42,In_296);
and U626 (N_626,In_267,In_50);
nor U627 (N_627,In_390,In_266);
xor U628 (N_628,In_383,In_411);
xor U629 (N_629,In_212,In_31);
nor U630 (N_630,In_349,In_307);
and U631 (N_631,In_349,In_203);
nor U632 (N_632,In_358,In_400);
nand U633 (N_633,In_154,In_165);
xnor U634 (N_634,In_85,In_457);
nand U635 (N_635,In_264,In_36);
and U636 (N_636,In_107,In_332);
nand U637 (N_637,In_105,In_176);
or U638 (N_638,In_253,In_231);
and U639 (N_639,In_244,In_345);
nand U640 (N_640,In_81,In_175);
or U641 (N_641,In_211,In_27);
nor U642 (N_642,In_160,In_108);
or U643 (N_643,In_313,In_83);
and U644 (N_644,In_308,In_292);
or U645 (N_645,In_429,In_288);
xnor U646 (N_646,In_155,In_478);
nand U647 (N_647,In_365,In_165);
xnor U648 (N_648,In_466,In_71);
and U649 (N_649,In_181,In_274);
and U650 (N_650,In_196,In_269);
xnor U651 (N_651,In_260,In_358);
nor U652 (N_652,In_222,In_144);
and U653 (N_653,In_95,In_440);
xor U654 (N_654,In_145,In_188);
or U655 (N_655,In_442,In_469);
nor U656 (N_656,In_292,In_282);
or U657 (N_657,In_465,In_495);
and U658 (N_658,In_251,In_285);
nand U659 (N_659,In_19,In_345);
or U660 (N_660,In_18,In_1);
nand U661 (N_661,In_253,In_409);
and U662 (N_662,In_470,In_314);
xor U663 (N_663,In_10,In_86);
xnor U664 (N_664,In_190,In_63);
nor U665 (N_665,In_74,In_94);
and U666 (N_666,In_39,In_202);
nand U667 (N_667,In_499,In_17);
xnor U668 (N_668,In_140,In_222);
nand U669 (N_669,In_441,In_35);
nor U670 (N_670,In_77,In_152);
and U671 (N_671,In_260,In_344);
nand U672 (N_672,In_353,In_37);
nand U673 (N_673,In_25,In_268);
nor U674 (N_674,In_224,In_7);
or U675 (N_675,In_288,In_130);
nand U676 (N_676,In_263,In_79);
nor U677 (N_677,In_395,In_103);
nor U678 (N_678,In_30,In_452);
xor U679 (N_679,In_278,In_61);
or U680 (N_680,In_111,In_286);
xor U681 (N_681,In_183,In_256);
xor U682 (N_682,In_150,In_272);
nor U683 (N_683,In_399,In_345);
nand U684 (N_684,In_368,In_350);
and U685 (N_685,In_14,In_37);
nand U686 (N_686,In_381,In_20);
nand U687 (N_687,In_394,In_341);
nand U688 (N_688,In_203,In_466);
or U689 (N_689,In_108,In_315);
xor U690 (N_690,In_497,In_316);
nand U691 (N_691,In_98,In_213);
or U692 (N_692,In_218,In_241);
nor U693 (N_693,In_448,In_54);
nor U694 (N_694,In_324,In_367);
or U695 (N_695,In_427,In_180);
nand U696 (N_696,In_277,In_41);
or U697 (N_697,In_272,In_227);
nor U698 (N_698,In_483,In_473);
and U699 (N_699,In_383,In_369);
and U700 (N_700,In_440,In_223);
and U701 (N_701,In_376,In_316);
or U702 (N_702,In_162,In_26);
nand U703 (N_703,In_464,In_461);
or U704 (N_704,In_362,In_232);
or U705 (N_705,In_209,In_8);
or U706 (N_706,In_48,In_184);
nor U707 (N_707,In_60,In_19);
xnor U708 (N_708,In_208,In_445);
and U709 (N_709,In_208,In_287);
nand U710 (N_710,In_167,In_1);
and U711 (N_711,In_92,In_298);
xnor U712 (N_712,In_480,In_287);
and U713 (N_713,In_29,In_245);
nor U714 (N_714,In_251,In_310);
and U715 (N_715,In_110,In_298);
and U716 (N_716,In_335,In_291);
and U717 (N_717,In_336,In_266);
xor U718 (N_718,In_149,In_79);
xnor U719 (N_719,In_192,In_3);
or U720 (N_720,In_25,In_229);
and U721 (N_721,In_386,In_217);
nand U722 (N_722,In_447,In_5);
xor U723 (N_723,In_428,In_144);
nor U724 (N_724,In_69,In_38);
nor U725 (N_725,In_273,In_149);
and U726 (N_726,In_185,In_414);
nand U727 (N_727,In_314,In_430);
and U728 (N_728,In_332,In_305);
nor U729 (N_729,In_85,In_420);
xor U730 (N_730,In_335,In_490);
or U731 (N_731,In_387,In_38);
xor U732 (N_732,In_333,In_418);
nor U733 (N_733,In_113,In_38);
and U734 (N_734,In_334,In_237);
or U735 (N_735,In_378,In_312);
xor U736 (N_736,In_456,In_102);
nor U737 (N_737,In_428,In_304);
nor U738 (N_738,In_398,In_333);
or U739 (N_739,In_218,In_459);
nor U740 (N_740,In_160,In_163);
nor U741 (N_741,In_99,In_317);
and U742 (N_742,In_176,In_273);
xor U743 (N_743,In_76,In_411);
or U744 (N_744,In_25,In_451);
nand U745 (N_745,In_157,In_337);
and U746 (N_746,In_228,In_46);
or U747 (N_747,In_219,In_25);
nor U748 (N_748,In_124,In_138);
nand U749 (N_749,In_466,In_38);
nor U750 (N_750,In_488,In_296);
or U751 (N_751,In_33,In_245);
nand U752 (N_752,In_431,In_309);
and U753 (N_753,In_459,In_17);
nand U754 (N_754,In_108,In_156);
or U755 (N_755,In_442,In_490);
nor U756 (N_756,In_407,In_81);
nor U757 (N_757,In_192,In_245);
nor U758 (N_758,In_406,In_197);
nand U759 (N_759,In_482,In_166);
xnor U760 (N_760,In_313,In_134);
nor U761 (N_761,In_493,In_324);
or U762 (N_762,In_11,In_354);
nor U763 (N_763,In_286,In_475);
or U764 (N_764,In_359,In_313);
and U765 (N_765,In_408,In_152);
nor U766 (N_766,In_178,In_154);
nor U767 (N_767,In_207,In_165);
nor U768 (N_768,In_449,In_456);
nor U769 (N_769,In_316,In_460);
xnor U770 (N_770,In_17,In_423);
xnor U771 (N_771,In_424,In_22);
nor U772 (N_772,In_320,In_257);
nand U773 (N_773,In_169,In_446);
nand U774 (N_774,In_248,In_50);
nor U775 (N_775,In_311,In_331);
nand U776 (N_776,In_66,In_403);
nand U777 (N_777,In_322,In_476);
nor U778 (N_778,In_476,In_340);
xor U779 (N_779,In_482,In_353);
xnor U780 (N_780,In_46,In_389);
xor U781 (N_781,In_113,In_417);
xnor U782 (N_782,In_296,In_438);
nor U783 (N_783,In_342,In_175);
nand U784 (N_784,In_113,In_190);
or U785 (N_785,In_101,In_411);
nor U786 (N_786,In_452,In_170);
or U787 (N_787,In_224,In_324);
nand U788 (N_788,In_15,In_439);
xnor U789 (N_789,In_47,In_440);
nor U790 (N_790,In_212,In_282);
xnor U791 (N_791,In_152,In_488);
nor U792 (N_792,In_207,In_381);
nor U793 (N_793,In_375,In_283);
nand U794 (N_794,In_23,In_292);
or U795 (N_795,In_252,In_488);
or U796 (N_796,In_59,In_78);
or U797 (N_797,In_33,In_349);
and U798 (N_798,In_324,In_116);
nor U799 (N_799,In_267,In_120);
nor U800 (N_800,In_191,In_388);
nor U801 (N_801,In_456,In_283);
xor U802 (N_802,In_445,In_435);
xor U803 (N_803,In_296,In_459);
nand U804 (N_804,In_77,In_92);
xnor U805 (N_805,In_63,In_102);
and U806 (N_806,In_347,In_177);
and U807 (N_807,In_267,In_285);
or U808 (N_808,In_282,In_439);
nand U809 (N_809,In_274,In_153);
xnor U810 (N_810,In_20,In_253);
and U811 (N_811,In_468,In_45);
nand U812 (N_812,In_427,In_333);
or U813 (N_813,In_199,In_295);
nor U814 (N_814,In_438,In_86);
and U815 (N_815,In_192,In_210);
nand U816 (N_816,In_253,In_162);
or U817 (N_817,In_448,In_274);
or U818 (N_818,In_342,In_237);
nand U819 (N_819,In_0,In_235);
xnor U820 (N_820,In_292,In_168);
nand U821 (N_821,In_231,In_418);
nand U822 (N_822,In_322,In_318);
or U823 (N_823,In_283,In_471);
and U824 (N_824,In_117,In_492);
nand U825 (N_825,In_343,In_42);
nor U826 (N_826,In_167,In_51);
and U827 (N_827,In_341,In_270);
xnor U828 (N_828,In_198,In_390);
nand U829 (N_829,In_239,In_42);
nor U830 (N_830,In_460,In_435);
or U831 (N_831,In_73,In_31);
and U832 (N_832,In_282,In_258);
nand U833 (N_833,In_330,In_474);
nor U834 (N_834,In_152,In_441);
nand U835 (N_835,In_139,In_390);
xnor U836 (N_836,In_415,In_107);
and U837 (N_837,In_213,In_322);
nor U838 (N_838,In_405,In_385);
xor U839 (N_839,In_213,In_248);
or U840 (N_840,In_371,In_271);
nor U841 (N_841,In_362,In_470);
and U842 (N_842,In_405,In_63);
xnor U843 (N_843,In_6,In_168);
nor U844 (N_844,In_292,In_331);
nor U845 (N_845,In_378,In_227);
or U846 (N_846,In_333,In_215);
xnor U847 (N_847,In_17,In_41);
nand U848 (N_848,In_391,In_192);
xor U849 (N_849,In_429,In_245);
nor U850 (N_850,In_464,In_342);
nand U851 (N_851,In_489,In_230);
xnor U852 (N_852,In_353,In_57);
and U853 (N_853,In_32,In_363);
xnor U854 (N_854,In_381,In_158);
nor U855 (N_855,In_300,In_331);
or U856 (N_856,In_168,In_80);
or U857 (N_857,In_67,In_31);
xor U858 (N_858,In_490,In_39);
nor U859 (N_859,In_310,In_497);
and U860 (N_860,In_94,In_355);
and U861 (N_861,In_374,In_185);
nor U862 (N_862,In_334,In_194);
nand U863 (N_863,In_469,In_103);
and U864 (N_864,In_0,In_27);
and U865 (N_865,In_166,In_249);
nand U866 (N_866,In_50,In_371);
and U867 (N_867,In_180,In_184);
or U868 (N_868,In_167,In_499);
and U869 (N_869,In_68,In_207);
or U870 (N_870,In_84,In_50);
xnor U871 (N_871,In_140,In_71);
and U872 (N_872,In_222,In_82);
and U873 (N_873,In_358,In_196);
nand U874 (N_874,In_385,In_143);
and U875 (N_875,In_448,In_389);
and U876 (N_876,In_256,In_384);
and U877 (N_877,In_221,In_181);
and U878 (N_878,In_354,In_317);
nand U879 (N_879,In_58,In_348);
nand U880 (N_880,In_214,In_379);
nor U881 (N_881,In_0,In_416);
or U882 (N_882,In_175,In_438);
nand U883 (N_883,In_383,In_241);
nor U884 (N_884,In_272,In_329);
or U885 (N_885,In_61,In_349);
nor U886 (N_886,In_497,In_108);
nand U887 (N_887,In_468,In_80);
and U888 (N_888,In_391,In_291);
or U889 (N_889,In_28,In_277);
nor U890 (N_890,In_468,In_360);
xor U891 (N_891,In_379,In_198);
and U892 (N_892,In_27,In_451);
nor U893 (N_893,In_8,In_134);
nor U894 (N_894,In_463,In_297);
nand U895 (N_895,In_378,In_354);
nor U896 (N_896,In_171,In_348);
nor U897 (N_897,In_341,In_399);
nor U898 (N_898,In_290,In_193);
and U899 (N_899,In_312,In_149);
nor U900 (N_900,In_269,In_22);
and U901 (N_901,In_490,In_100);
or U902 (N_902,In_181,In_186);
nor U903 (N_903,In_196,In_13);
and U904 (N_904,In_35,In_135);
xnor U905 (N_905,In_359,In_71);
nor U906 (N_906,In_128,In_406);
nor U907 (N_907,In_311,In_349);
nor U908 (N_908,In_163,In_370);
nand U909 (N_909,In_393,In_48);
or U910 (N_910,In_262,In_397);
and U911 (N_911,In_425,In_186);
or U912 (N_912,In_250,In_262);
nand U913 (N_913,In_421,In_285);
or U914 (N_914,In_45,In_37);
xnor U915 (N_915,In_351,In_420);
nor U916 (N_916,In_325,In_141);
nand U917 (N_917,In_401,In_58);
and U918 (N_918,In_428,In_253);
nand U919 (N_919,In_22,In_334);
or U920 (N_920,In_35,In_390);
xnor U921 (N_921,In_79,In_192);
nand U922 (N_922,In_291,In_184);
or U923 (N_923,In_379,In_253);
and U924 (N_924,In_33,In_214);
nand U925 (N_925,In_110,In_57);
xnor U926 (N_926,In_120,In_147);
and U927 (N_927,In_25,In_103);
nand U928 (N_928,In_104,In_431);
and U929 (N_929,In_107,In_356);
xnor U930 (N_930,In_252,In_497);
xnor U931 (N_931,In_301,In_336);
nor U932 (N_932,In_25,In_76);
nand U933 (N_933,In_371,In_195);
and U934 (N_934,In_114,In_139);
nand U935 (N_935,In_87,In_231);
nand U936 (N_936,In_326,In_105);
nand U937 (N_937,In_329,In_177);
or U938 (N_938,In_413,In_435);
and U939 (N_939,In_496,In_9);
xor U940 (N_940,In_113,In_77);
nand U941 (N_941,In_376,In_193);
or U942 (N_942,In_245,In_375);
and U943 (N_943,In_21,In_119);
and U944 (N_944,In_264,In_18);
or U945 (N_945,In_176,In_19);
nand U946 (N_946,In_265,In_67);
nand U947 (N_947,In_8,In_330);
nand U948 (N_948,In_201,In_6);
nor U949 (N_949,In_364,In_368);
xor U950 (N_950,In_477,In_6);
and U951 (N_951,In_390,In_96);
and U952 (N_952,In_92,In_415);
and U953 (N_953,In_24,In_175);
nor U954 (N_954,In_400,In_305);
and U955 (N_955,In_282,In_342);
xor U956 (N_956,In_4,In_236);
nand U957 (N_957,In_45,In_277);
or U958 (N_958,In_227,In_382);
xnor U959 (N_959,In_433,In_83);
xor U960 (N_960,In_211,In_221);
and U961 (N_961,In_218,In_94);
and U962 (N_962,In_403,In_402);
or U963 (N_963,In_256,In_327);
and U964 (N_964,In_154,In_23);
or U965 (N_965,In_291,In_8);
nor U966 (N_966,In_7,In_168);
xor U967 (N_967,In_33,In_239);
xor U968 (N_968,In_345,In_101);
nor U969 (N_969,In_148,In_123);
nand U970 (N_970,In_2,In_6);
nor U971 (N_971,In_387,In_368);
and U972 (N_972,In_75,In_8);
or U973 (N_973,In_348,In_68);
nand U974 (N_974,In_277,In_481);
nand U975 (N_975,In_474,In_26);
nand U976 (N_976,In_468,In_223);
or U977 (N_977,In_151,In_25);
nand U978 (N_978,In_154,In_47);
nor U979 (N_979,In_490,In_179);
nand U980 (N_980,In_91,In_259);
nand U981 (N_981,In_174,In_470);
nand U982 (N_982,In_341,In_301);
nor U983 (N_983,In_441,In_87);
or U984 (N_984,In_476,In_201);
xnor U985 (N_985,In_55,In_242);
xor U986 (N_986,In_131,In_421);
nand U987 (N_987,In_142,In_37);
and U988 (N_988,In_481,In_205);
xor U989 (N_989,In_303,In_14);
and U990 (N_990,In_368,In_146);
xor U991 (N_991,In_51,In_364);
xnor U992 (N_992,In_88,In_393);
nor U993 (N_993,In_78,In_87);
nand U994 (N_994,In_316,In_427);
xor U995 (N_995,In_200,In_49);
nor U996 (N_996,In_231,In_406);
nor U997 (N_997,In_424,In_281);
and U998 (N_998,In_152,In_103);
xor U999 (N_999,In_379,In_222);
or U1000 (N_1000,N_979,N_804);
or U1001 (N_1001,N_7,N_430);
nand U1002 (N_1002,N_665,N_428);
nor U1003 (N_1003,N_135,N_862);
or U1004 (N_1004,N_825,N_578);
or U1005 (N_1005,N_499,N_86);
and U1006 (N_1006,N_95,N_706);
and U1007 (N_1007,N_128,N_652);
and U1008 (N_1008,N_259,N_580);
nor U1009 (N_1009,N_912,N_200);
or U1010 (N_1010,N_212,N_105);
xor U1011 (N_1011,N_208,N_348);
or U1012 (N_1012,N_799,N_643);
xor U1013 (N_1013,N_545,N_579);
nand U1014 (N_1014,N_368,N_424);
nor U1015 (N_1015,N_645,N_795);
or U1016 (N_1016,N_509,N_239);
nor U1017 (N_1017,N_951,N_561);
or U1018 (N_1018,N_699,N_146);
nand U1019 (N_1019,N_818,N_187);
nand U1020 (N_1020,N_589,N_680);
and U1021 (N_1021,N_185,N_925);
nor U1022 (N_1022,N_178,N_961);
and U1023 (N_1023,N_916,N_887);
xor U1024 (N_1024,N_759,N_232);
and U1025 (N_1025,N_634,N_924);
nand U1026 (N_1026,N_974,N_851);
and U1027 (N_1027,N_882,N_411);
nand U1028 (N_1028,N_560,N_385);
xnor U1029 (N_1029,N_553,N_326);
nand U1030 (N_1030,N_481,N_529);
nand U1031 (N_1031,N_418,N_335);
and U1032 (N_1032,N_915,N_911);
nand U1033 (N_1033,N_606,N_164);
or U1034 (N_1034,N_814,N_594);
nor U1035 (N_1035,N_447,N_848);
and U1036 (N_1036,N_253,N_454);
and U1037 (N_1037,N_453,N_0);
nand U1038 (N_1038,N_728,N_83);
nor U1039 (N_1039,N_38,N_391);
xnor U1040 (N_1040,N_715,N_46);
nor U1041 (N_1041,N_797,N_275);
xor U1042 (N_1042,N_931,N_539);
or U1043 (N_1043,N_605,N_96);
and U1044 (N_1044,N_803,N_279);
and U1045 (N_1045,N_273,N_521);
xor U1046 (N_1046,N_115,N_708);
xnor U1047 (N_1047,N_775,N_792);
xor U1048 (N_1048,N_733,N_767);
or U1049 (N_1049,N_150,N_888);
nor U1050 (N_1050,N_513,N_49);
or U1051 (N_1051,N_532,N_820);
and U1052 (N_1052,N_55,N_462);
or U1053 (N_1053,N_635,N_399);
nand U1054 (N_1054,N_928,N_197);
nor U1055 (N_1055,N_317,N_741);
or U1056 (N_1056,N_941,N_672);
or U1057 (N_1057,N_698,N_163);
nand U1058 (N_1058,N_495,N_396);
xnor U1059 (N_1059,N_661,N_547);
nand U1060 (N_1060,N_933,N_750);
and U1061 (N_1061,N_946,N_692);
xor U1062 (N_1062,N_423,N_686);
xor U1063 (N_1063,N_235,N_32);
nand U1064 (N_1064,N_303,N_439);
or U1065 (N_1065,N_821,N_768);
nor U1066 (N_1066,N_422,N_548);
xor U1067 (N_1067,N_190,N_774);
nor U1068 (N_1068,N_894,N_726);
and U1069 (N_1069,N_593,N_446);
or U1070 (N_1070,N_585,N_564);
or U1071 (N_1071,N_160,N_581);
and U1072 (N_1072,N_247,N_771);
nand U1073 (N_1073,N_963,N_909);
and U1074 (N_1074,N_568,N_230);
and U1075 (N_1075,N_754,N_215);
xor U1076 (N_1076,N_875,N_778);
or U1077 (N_1077,N_865,N_47);
xor U1078 (N_1078,N_267,N_196);
nand U1079 (N_1079,N_989,N_758);
xor U1080 (N_1080,N_709,N_808);
nor U1081 (N_1081,N_92,N_807);
or U1082 (N_1082,N_796,N_458);
nor U1083 (N_1083,N_588,N_631);
and U1084 (N_1084,N_638,N_50);
xnor U1085 (N_1085,N_477,N_650);
xor U1086 (N_1086,N_857,N_505);
nor U1087 (N_1087,N_188,N_78);
nor U1088 (N_1088,N_599,N_355);
and U1089 (N_1089,N_993,N_132);
and U1090 (N_1090,N_11,N_166);
xnor U1091 (N_1091,N_249,N_44);
nor U1092 (N_1092,N_297,N_877);
nor U1093 (N_1093,N_624,N_711);
or U1094 (N_1094,N_263,N_536);
and U1095 (N_1095,N_41,N_476);
xnor U1096 (N_1096,N_173,N_784);
xnor U1097 (N_1097,N_122,N_15);
or U1098 (N_1098,N_782,N_535);
nand U1099 (N_1099,N_710,N_25);
nand U1100 (N_1100,N_681,N_21);
nand U1101 (N_1101,N_633,N_881);
nor U1102 (N_1102,N_113,N_964);
nand U1103 (N_1103,N_359,N_981);
nor U1104 (N_1104,N_613,N_219);
nand U1105 (N_1105,N_492,N_443);
and U1106 (N_1106,N_859,N_378);
xor U1107 (N_1107,N_183,N_341);
nand U1108 (N_1108,N_660,N_864);
and U1109 (N_1109,N_811,N_838);
xor U1110 (N_1110,N_584,N_283);
and U1111 (N_1111,N_976,N_119);
and U1112 (N_1112,N_855,N_39);
xor U1113 (N_1113,N_969,N_436);
or U1114 (N_1114,N_468,N_318);
or U1115 (N_1115,N_842,N_9);
nand U1116 (N_1116,N_787,N_365);
or U1117 (N_1117,N_252,N_59);
and U1118 (N_1118,N_860,N_56);
or U1119 (N_1119,N_413,N_639);
xnor U1120 (N_1120,N_280,N_8);
nor U1121 (N_1121,N_270,N_383);
and U1122 (N_1122,N_824,N_421);
and U1123 (N_1123,N_432,N_702);
or U1124 (N_1124,N_497,N_556);
nand U1125 (N_1125,N_379,N_12);
or U1126 (N_1126,N_995,N_871);
and U1127 (N_1127,N_694,N_245);
or U1128 (N_1128,N_143,N_216);
or U1129 (N_1129,N_813,N_748);
nand U1130 (N_1130,N_389,N_986);
and U1131 (N_1131,N_337,N_696);
nand U1132 (N_1132,N_314,N_61);
nand U1133 (N_1133,N_193,N_919);
xor U1134 (N_1134,N_129,N_101);
nor U1135 (N_1135,N_316,N_576);
nand U1136 (N_1136,N_971,N_89);
nand U1137 (N_1137,N_721,N_308);
xor U1138 (N_1138,N_97,N_147);
nand U1139 (N_1139,N_315,N_831);
nor U1140 (N_1140,N_144,N_984);
xor U1141 (N_1141,N_414,N_222);
or U1142 (N_1142,N_701,N_401);
or U1143 (N_1143,N_338,N_358);
xnor U1144 (N_1144,N_177,N_372);
or U1145 (N_1145,N_408,N_920);
nand U1146 (N_1146,N_610,N_679);
xor U1147 (N_1147,N_623,N_134);
or U1148 (N_1148,N_714,N_171);
xnor U1149 (N_1149,N_738,N_781);
xor U1150 (N_1150,N_440,N_457);
and U1151 (N_1151,N_868,N_107);
or U1152 (N_1152,N_240,N_324);
or U1153 (N_1153,N_730,N_713);
nor U1154 (N_1154,N_640,N_843);
nand U1155 (N_1155,N_206,N_374);
and U1156 (N_1156,N_498,N_716);
xor U1157 (N_1157,N_571,N_675);
and U1158 (N_1158,N_935,N_646);
or U1159 (N_1159,N_35,N_116);
nand U1160 (N_1160,N_282,N_24);
and U1161 (N_1161,N_292,N_511);
xnor U1162 (N_1162,N_71,N_937);
or U1163 (N_1163,N_350,N_745);
nor U1164 (N_1164,N_298,N_910);
and U1165 (N_1165,N_583,N_494);
nand U1166 (N_1166,N_345,N_667);
nand U1167 (N_1167,N_75,N_563);
nand U1168 (N_1168,N_33,N_531);
and U1169 (N_1169,N_866,N_527);
xor U1170 (N_1170,N_697,N_203);
nor U1171 (N_1171,N_405,N_67);
or U1172 (N_1172,N_943,N_743);
nor U1173 (N_1173,N_471,N_63);
and U1174 (N_1174,N_788,N_344);
nand U1175 (N_1175,N_815,N_802);
nand U1176 (N_1176,N_102,N_123);
or U1177 (N_1177,N_22,N_671);
nor U1178 (N_1178,N_502,N_988);
or U1179 (N_1179,N_31,N_523);
nand U1180 (N_1180,N_977,N_844);
xor U1181 (N_1181,N_900,N_192);
nand U1182 (N_1182,N_210,N_966);
or U1183 (N_1183,N_947,N_729);
xnor U1184 (N_1184,N_172,N_668);
nor U1185 (N_1185,N_762,N_293);
nand U1186 (N_1186,N_903,N_742);
nand U1187 (N_1187,N_524,N_121);
and U1188 (N_1188,N_822,N_769);
xor U1189 (N_1189,N_908,N_373);
xnor U1190 (N_1190,N_306,N_510);
or U1191 (N_1191,N_978,N_948);
xnor U1192 (N_1192,N_334,N_836);
xnor U1193 (N_1193,N_357,N_112);
and U1194 (N_1194,N_403,N_323);
and U1195 (N_1195,N_707,N_299);
or U1196 (N_1196,N_154,N_155);
nor U1197 (N_1197,N_397,N_766);
nor U1198 (N_1198,N_213,N_609);
xnor U1199 (N_1199,N_780,N_256);
nand U1200 (N_1200,N_302,N_456);
and U1201 (N_1201,N_789,N_705);
or U1202 (N_1202,N_437,N_596);
and U1203 (N_1203,N_20,N_982);
xnor U1204 (N_1204,N_734,N_999);
or U1205 (N_1205,N_770,N_330);
and U1206 (N_1206,N_290,N_835);
nand U1207 (N_1207,N_79,N_930);
nand U1208 (N_1208,N_834,N_327);
xor U1209 (N_1209,N_281,N_258);
nor U1210 (N_1210,N_902,N_351);
xor U1211 (N_1211,N_179,N_597);
nor U1212 (N_1212,N_879,N_950);
xor U1213 (N_1213,N_313,N_74);
nand U1214 (N_1214,N_243,N_478);
or U1215 (N_1215,N_674,N_801);
xor U1216 (N_1216,N_572,N_817);
and U1217 (N_1217,N_174,N_914);
nor U1218 (N_1218,N_501,N_62);
or U1219 (N_1219,N_221,N_603);
nand U1220 (N_1220,N_242,N_990);
nand U1221 (N_1221,N_893,N_904);
nand U1222 (N_1222,N_136,N_783);
and U1223 (N_1223,N_225,N_170);
nand U1224 (N_1224,N_390,N_812);
and U1225 (N_1225,N_967,N_142);
xnor U1226 (N_1226,N_139,N_923);
and U1227 (N_1227,N_764,N_80);
and U1228 (N_1228,N_181,N_936);
nand U1229 (N_1229,N_255,N_410);
xor U1230 (N_1230,N_451,N_272);
nor U1231 (N_1231,N_231,N_870);
nand U1232 (N_1232,N_892,N_393);
or U1233 (N_1233,N_637,N_426);
nor U1234 (N_1234,N_991,N_354);
and U1235 (N_1235,N_490,N_541);
or U1236 (N_1236,N_333,N_574);
nor U1237 (N_1237,N_546,N_566);
nand U1238 (N_1238,N_994,N_305);
nor U1239 (N_1239,N_737,N_727);
nand U1240 (N_1240,N_100,N_890);
nor U1241 (N_1241,N_582,N_854);
or U1242 (N_1242,N_211,N_472);
and U1243 (N_1243,N_621,N_703);
and U1244 (N_1244,N_141,N_400);
nor U1245 (N_1245,N_678,N_538);
nand U1246 (N_1246,N_284,N_474);
and U1247 (N_1247,N_360,N_29);
nor U1248 (N_1248,N_406,N_427);
nand U1249 (N_1249,N_356,N_725);
or U1250 (N_1250,N_620,N_85);
nand U1251 (N_1251,N_772,N_244);
or U1252 (N_1252,N_328,N_684);
nor U1253 (N_1253,N_653,N_73);
nor U1254 (N_1254,N_312,N_677);
or U1255 (N_1255,N_590,N_885);
xnor U1256 (N_1256,N_189,N_852);
nand U1257 (N_1257,N_347,N_528);
and U1258 (N_1258,N_228,N_370);
xor U1259 (N_1259,N_214,N_809);
nor U1260 (N_1260,N_636,N_664);
nor U1261 (N_1261,N_644,N_901);
or U1262 (N_1262,N_839,N_630);
or U1263 (N_1263,N_987,N_223);
nand U1264 (N_1264,N_929,N_167);
and U1265 (N_1265,N_884,N_227);
or U1266 (N_1266,N_899,N_558);
nor U1267 (N_1267,N_309,N_632);
or U1268 (N_1268,N_688,N_786);
or U1269 (N_1269,N_118,N_199);
xnor U1270 (N_1270,N_626,N_550);
nor U1271 (N_1271,N_349,N_412);
xor U1272 (N_1272,N_957,N_570);
or U1273 (N_1273,N_878,N_233);
and U1274 (N_1274,N_180,N_450);
or U1275 (N_1275,N_549,N_869);
nand U1276 (N_1276,N_70,N_627);
and U1277 (N_1277,N_651,N_739);
xor U1278 (N_1278,N_717,N_751);
xor U1279 (N_1279,N_500,N_156);
or U1280 (N_1280,N_420,N_271);
nor U1281 (N_1281,N_525,N_286);
nand U1282 (N_1282,N_496,N_612);
or U1283 (N_1283,N_954,N_506);
nor U1284 (N_1284,N_704,N_891);
nor U1285 (N_1285,N_201,N_16);
or U1286 (N_1286,N_417,N_876);
nor U1287 (N_1287,N_598,N_322);
and U1288 (N_1288,N_998,N_441);
xnor U1289 (N_1289,N_830,N_922);
nor U1290 (N_1290,N_184,N_254);
nor U1291 (N_1291,N_310,N_514);
and U1292 (N_1292,N_618,N_301);
nand U1293 (N_1293,N_5,N_133);
xnor U1294 (N_1294,N_224,N_896);
xnor U1295 (N_1295,N_562,N_757);
nor U1296 (N_1296,N_387,N_36);
nor U1297 (N_1297,N_66,N_586);
nand U1298 (N_1298,N_266,N_269);
and U1299 (N_1299,N_724,N_104);
nand U1300 (N_1300,N_926,N_84);
nand U1301 (N_1301,N_37,N_274);
nand U1302 (N_1302,N_760,N_949);
and U1303 (N_1303,N_205,N_241);
nor U1304 (N_1304,N_491,N_176);
xor U1305 (N_1305,N_542,N_445);
nand U1306 (N_1306,N_264,N_980);
and U1307 (N_1307,N_13,N_518);
and U1308 (N_1308,N_194,N_601);
and U1309 (N_1309,N_87,N_395);
xor U1310 (N_1310,N_363,N_493);
and U1311 (N_1311,N_898,N_23);
nand U1312 (N_1312,N_939,N_676);
or U1313 (N_1313,N_960,N_431);
or U1314 (N_1314,N_559,N_459);
or U1315 (N_1315,N_364,N_693);
or U1316 (N_1316,N_861,N_889);
and U1317 (N_1317,N_433,N_968);
nor U1318 (N_1318,N_625,N_469);
and U1319 (N_1319,N_773,N_973);
nor U1320 (N_1320,N_319,N_700);
xor U1321 (N_1321,N_617,N_791);
and U1322 (N_1322,N_287,N_508);
or U1323 (N_1323,N_27,N_744);
nor U1324 (N_1324,N_465,N_735);
nor U1325 (N_1325,N_260,N_777);
nand U1326 (N_1326,N_366,N_666);
or U1327 (N_1327,N_731,N_261);
nand U1328 (N_1328,N_4,N_209);
nor U1329 (N_1329,N_392,N_806);
and U1330 (N_1330,N_753,N_856);
or U1331 (N_1331,N_161,N_845);
xnor U1332 (N_1332,N_198,N_793);
nor U1333 (N_1333,N_863,N_463);
and U1334 (N_1334,N_850,N_145);
xor U1335 (N_1335,N_402,N_448);
or U1336 (N_1336,N_934,N_763);
nor U1337 (N_1337,N_985,N_304);
nor U1338 (N_1338,N_19,N_43);
xnor U1339 (N_1339,N_880,N_220);
or U1340 (N_1340,N_654,N_40);
xnor U1341 (N_1341,N_26,N_776);
or U1342 (N_1342,N_77,N_289);
and U1343 (N_1343,N_157,N_690);
and U1344 (N_1344,N_996,N_386);
nor U1345 (N_1345,N_434,N_959);
nand U1346 (N_1346,N_460,N_992);
nor U1347 (N_1347,N_14,N_798);
or U1348 (N_1348,N_407,N_103);
or U1349 (N_1349,N_614,N_111);
nand U1350 (N_1350,N_276,N_153);
nand U1351 (N_1351,N_732,N_217);
nand U1352 (N_1352,N_554,N_873);
nor U1353 (N_1353,N_484,N_28);
or U1354 (N_1354,N_442,N_819);
or U1355 (N_1355,N_906,N_895);
or U1356 (N_1356,N_207,N_140);
nand U1357 (N_1357,N_51,N_6);
nor U1358 (N_1358,N_361,N_805);
nand U1359 (N_1359,N_695,N_965);
and U1360 (N_1360,N_332,N_1);
nand U1361 (N_1361,N_526,N_68);
and U1362 (N_1362,N_752,N_975);
and U1363 (N_1363,N_375,N_816);
and U1364 (N_1364,N_482,N_600);
xnor U1365 (N_1365,N_311,N_555);
xor U1366 (N_1366,N_246,N_486);
or U1367 (N_1367,N_503,N_747);
nand U1368 (N_1368,N_718,N_520);
or U1369 (N_1369,N_331,N_615);
nand U1370 (N_1370,N_336,N_91);
nand U1371 (N_1371,N_522,N_69);
nand U1372 (N_1372,N_883,N_234);
or U1373 (N_1373,N_565,N_321);
nand U1374 (N_1374,N_577,N_828);
nor U1375 (N_1375,N_685,N_250);
nor U1376 (N_1376,N_785,N_740);
nor U1377 (N_1377,N_339,N_353);
xnor U1378 (N_1378,N_972,N_874);
nand U1379 (N_1379,N_669,N_106);
and U1380 (N_1380,N_404,N_204);
or U1381 (N_1381,N_288,N_673);
xnor U1382 (N_1382,N_940,N_749);
and U1383 (N_1383,N_853,N_438);
nor U1384 (N_1384,N_48,N_682);
xnor U1385 (N_1385,N_186,N_569);
xor U1386 (N_1386,N_648,N_466);
nor U1387 (N_1387,N_997,N_125);
xor U1388 (N_1388,N_962,N_905);
and U1389 (N_1389,N_512,N_575);
xnor U1390 (N_1390,N_126,N_833);
and U1391 (N_1391,N_840,N_587);
nor U1392 (N_1392,N_64,N_544);
and U1393 (N_1393,N_218,N_592);
nand U1394 (N_1394,N_953,N_285);
nand U1395 (N_1395,N_983,N_921);
and U1396 (N_1396,N_380,N_124);
or U1397 (N_1397,N_779,N_109);
xnor U1398 (N_1398,N_352,N_425);
xnor U1399 (N_1399,N_226,N_191);
nand U1400 (N_1400,N_537,N_622);
xor U1401 (N_1401,N_483,N_300);
nand U1402 (N_1402,N_540,N_137);
or U1403 (N_1403,N_98,N_398);
and U1404 (N_1404,N_236,N_938);
nor U1405 (N_1405,N_159,N_543);
and U1406 (N_1406,N_719,N_641);
nand U1407 (N_1407,N_662,N_52);
xor U1408 (N_1408,N_473,N_670);
nand U1409 (N_1409,N_117,N_376);
xnor U1410 (N_1410,N_958,N_736);
nor U1411 (N_1411,N_794,N_165);
nor U1412 (N_1412,N_127,N_268);
and U1413 (N_1413,N_927,N_616);
and U1414 (N_1414,N_461,N_346);
xor U1415 (N_1415,N_872,N_608);
or U1416 (N_1416,N_534,N_573);
and U1417 (N_1417,N_278,N_151);
xor U1418 (N_1418,N_515,N_658);
nand U1419 (N_1419,N_800,N_384);
nand U1420 (N_1420,N_649,N_607);
xnor U1421 (N_1421,N_467,N_591);
nand U1422 (N_1422,N_294,N_53);
or U1423 (N_1423,N_970,N_381);
nor U1424 (N_1424,N_120,N_444);
or U1425 (N_1425,N_917,N_611);
nand U1426 (N_1426,N_507,N_683);
nor U1427 (N_1427,N_932,N_489);
xnor U1428 (N_1428,N_371,N_108);
nand U1429 (N_1429,N_504,N_94);
xor U1430 (N_1430,N_533,N_687);
nand U1431 (N_1431,N_82,N_913);
and U1432 (N_1432,N_148,N_790);
nand U1433 (N_1433,N_952,N_149);
nor U1434 (N_1434,N_761,N_195);
or U1435 (N_1435,N_659,N_846);
and U1436 (N_1436,N_168,N_60);
nand U1437 (N_1437,N_409,N_169);
or U1438 (N_1438,N_567,N_689);
xor U1439 (N_1439,N_452,N_756);
nand U1440 (N_1440,N_712,N_158);
nor U1441 (N_1441,N_76,N_867);
and U1442 (N_1442,N_897,N_602);
xor U1443 (N_1443,N_90,N_93);
or U1444 (N_1444,N_320,N_604);
and U1445 (N_1445,N_182,N_832);
nor U1446 (N_1446,N_394,N_340);
or U1447 (N_1447,N_628,N_595);
nand U1448 (N_1448,N_377,N_619);
nor U1449 (N_1449,N_918,N_829);
xor U1450 (N_1450,N_723,N_265);
xnor U1451 (N_1451,N_54,N_691);
nand U1452 (N_1452,N_647,N_480);
xor U1453 (N_1453,N_131,N_10);
nand U1454 (N_1454,N_858,N_519);
xnor U1455 (N_1455,N_202,N_362);
nor U1456 (N_1456,N_114,N_65);
or U1457 (N_1457,N_656,N_277);
and U1458 (N_1458,N_295,N_18);
nand U1459 (N_1459,N_942,N_517);
xnor U1460 (N_1460,N_837,N_30);
nor U1461 (N_1461,N_516,N_17);
nor U1462 (N_1462,N_435,N_765);
and U1463 (N_1463,N_956,N_629);
xnor U1464 (N_1464,N_826,N_475);
nor U1465 (N_1465,N_827,N_722);
and U1466 (N_1466,N_307,N_479);
and U1467 (N_1467,N_720,N_419);
or U1468 (N_1468,N_485,N_847);
nor U1469 (N_1469,N_57,N_944);
nor U1470 (N_1470,N_657,N_746);
nor U1471 (N_1471,N_382,N_557);
or U1472 (N_1472,N_130,N_110);
or U1473 (N_1473,N_449,N_470);
xor U1474 (N_1474,N_72,N_81);
nor U1475 (N_1475,N_369,N_88);
nor U1476 (N_1476,N_823,N_488);
and U1477 (N_1477,N_138,N_655);
xnor U1478 (N_1478,N_849,N_58);
nor U1479 (N_1479,N_251,N_464);
and U1480 (N_1480,N_175,N_329);
nor U1481 (N_1481,N_416,N_42);
or U1482 (N_1482,N_238,N_530);
or U1483 (N_1483,N_237,N_2);
or U1484 (N_1484,N_551,N_429);
and U1485 (N_1485,N_945,N_487);
and U1486 (N_1486,N_367,N_34);
nand U1487 (N_1487,N_886,N_907);
xnor U1488 (N_1488,N_415,N_343);
and U1489 (N_1489,N_755,N_841);
and U1490 (N_1490,N_257,N_642);
nor U1491 (N_1491,N_388,N_325);
nor U1492 (N_1492,N_248,N_663);
and U1493 (N_1493,N_45,N_342);
and U1494 (N_1494,N_99,N_810);
xnor U1495 (N_1495,N_3,N_955);
nor U1496 (N_1496,N_262,N_229);
nand U1497 (N_1497,N_455,N_296);
and U1498 (N_1498,N_552,N_152);
or U1499 (N_1499,N_162,N_291);
and U1500 (N_1500,N_387,N_741);
xor U1501 (N_1501,N_898,N_797);
nor U1502 (N_1502,N_47,N_155);
xnor U1503 (N_1503,N_514,N_778);
xor U1504 (N_1504,N_245,N_217);
nand U1505 (N_1505,N_746,N_119);
or U1506 (N_1506,N_880,N_289);
xnor U1507 (N_1507,N_450,N_26);
xnor U1508 (N_1508,N_436,N_384);
or U1509 (N_1509,N_352,N_25);
and U1510 (N_1510,N_378,N_13);
xnor U1511 (N_1511,N_159,N_667);
or U1512 (N_1512,N_540,N_584);
and U1513 (N_1513,N_174,N_249);
nand U1514 (N_1514,N_143,N_657);
or U1515 (N_1515,N_103,N_712);
or U1516 (N_1516,N_876,N_736);
nor U1517 (N_1517,N_865,N_522);
nand U1518 (N_1518,N_525,N_224);
nor U1519 (N_1519,N_808,N_578);
nand U1520 (N_1520,N_514,N_862);
xor U1521 (N_1521,N_495,N_723);
nor U1522 (N_1522,N_228,N_895);
nor U1523 (N_1523,N_256,N_259);
nor U1524 (N_1524,N_177,N_307);
xnor U1525 (N_1525,N_968,N_36);
or U1526 (N_1526,N_232,N_963);
or U1527 (N_1527,N_418,N_347);
nand U1528 (N_1528,N_470,N_745);
xnor U1529 (N_1529,N_776,N_19);
or U1530 (N_1530,N_3,N_893);
nor U1531 (N_1531,N_820,N_704);
or U1532 (N_1532,N_540,N_517);
nor U1533 (N_1533,N_922,N_288);
or U1534 (N_1534,N_231,N_477);
and U1535 (N_1535,N_195,N_806);
nand U1536 (N_1536,N_956,N_320);
nand U1537 (N_1537,N_876,N_998);
or U1538 (N_1538,N_166,N_488);
nand U1539 (N_1539,N_392,N_981);
or U1540 (N_1540,N_840,N_948);
nand U1541 (N_1541,N_308,N_560);
xnor U1542 (N_1542,N_453,N_902);
xor U1543 (N_1543,N_628,N_749);
or U1544 (N_1544,N_877,N_844);
xor U1545 (N_1545,N_115,N_849);
and U1546 (N_1546,N_615,N_699);
xnor U1547 (N_1547,N_616,N_98);
xor U1548 (N_1548,N_140,N_31);
and U1549 (N_1549,N_708,N_33);
nor U1550 (N_1550,N_621,N_214);
nand U1551 (N_1551,N_502,N_517);
and U1552 (N_1552,N_287,N_74);
nand U1553 (N_1553,N_496,N_471);
nor U1554 (N_1554,N_903,N_721);
nor U1555 (N_1555,N_918,N_759);
nand U1556 (N_1556,N_97,N_257);
nor U1557 (N_1557,N_634,N_855);
nor U1558 (N_1558,N_668,N_440);
and U1559 (N_1559,N_32,N_375);
or U1560 (N_1560,N_734,N_540);
and U1561 (N_1561,N_407,N_699);
xor U1562 (N_1562,N_689,N_933);
nor U1563 (N_1563,N_106,N_500);
nor U1564 (N_1564,N_113,N_934);
nand U1565 (N_1565,N_154,N_298);
xnor U1566 (N_1566,N_817,N_476);
or U1567 (N_1567,N_74,N_877);
xnor U1568 (N_1568,N_962,N_777);
xor U1569 (N_1569,N_24,N_524);
nor U1570 (N_1570,N_997,N_846);
nor U1571 (N_1571,N_883,N_792);
or U1572 (N_1572,N_654,N_269);
and U1573 (N_1573,N_604,N_178);
or U1574 (N_1574,N_977,N_736);
nor U1575 (N_1575,N_235,N_543);
xor U1576 (N_1576,N_498,N_515);
xnor U1577 (N_1577,N_788,N_506);
or U1578 (N_1578,N_933,N_952);
or U1579 (N_1579,N_35,N_115);
xor U1580 (N_1580,N_520,N_662);
xor U1581 (N_1581,N_698,N_324);
xnor U1582 (N_1582,N_937,N_910);
nor U1583 (N_1583,N_673,N_108);
or U1584 (N_1584,N_420,N_855);
xor U1585 (N_1585,N_256,N_288);
or U1586 (N_1586,N_771,N_876);
nand U1587 (N_1587,N_596,N_749);
nor U1588 (N_1588,N_251,N_687);
xnor U1589 (N_1589,N_255,N_388);
nand U1590 (N_1590,N_941,N_971);
or U1591 (N_1591,N_125,N_915);
nand U1592 (N_1592,N_87,N_373);
nand U1593 (N_1593,N_670,N_543);
xnor U1594 (N_1594,N_562,N_218);
nand U1595 (N_1595,N_603,N_878);
nand U1596 (N_1596,N_159,N_469);
or U1597 (N_1597,N_106,N_925);
xor U1598 (N_1598,N_927,N_890);
and U1599 (N_1599,N_14,N_337);
xnor U1600 (N_1600,N_665,N_180);
or U1601 (N_1601,N_394,N_828);
nor U1602 (N_1602,N_411,N_839);
xor U1603 (N_1603,N_25,N_650);
nor U1604 (N_1604,N_407,N_175);
or U1605 (N_1605,N_134,N_603);
and U1606 (N_1606,N_778,N_930);
xnor U1607 (N_1607,N_38,N_156);
nor U1608 (N_1608,N_34,N_634);
and U1609 (N_1609,N_337,N_594);
or U1610 (N_1610,N_246,N_720);
and U1611 (N_1611,N_455,N_755);
nor U1612 (N_1612,N_556,N_237);
nor U1613 (N_1613,N_79,N_332);
or U1614 (N_1614,N_291,N_46);
or U1615 (N_1615,N_389,N_802);
xnor U1616 (N_1616,N_728,N_463);
and U1617 (N_1617,N_741,N_673);
xnor U1618 (N_1618,N_62,N_410);
or U1619 (N_1619,N_736,N_441);
or U1620 (N_1620,N_767,N_941);
or U1621 (N_1621,N_823,N_518);
nor U1622 (N_1622,N_665,N_304);
and U1623 (N_1623,N_9,N_223);
xor U1624 (N_1624,N_129,N_845);
and U1625 (N_1625,N_962,N_985);
or U1626 (N_1626,N_885,N_360);
and U1627 (N_1627,N_123,N_581);
or U1628 (N_1628,N_329,N_591);
or U1629 (N_1629,N_285,N_916);
or U1630 (N_1630,N_914,N_241);
or U1631 (N_1631,N_888,N_249);
and U1632 (N_1632,N_412,N_875);
and U1633 (N_1633,N_176,N_321);
nor U1634 (N_1634,N_76,N_871);
nand U1635 (N_1635,N_624,N_655);
and U1636 (N_1636,N_455,N_774);
nand U1637 (N_1637,N_895,N_176);
nor U1638 (N_1638,N_986,N_348);
or U1639 (N_1639,N_936,N_352);
and U1640 (N_1640,N_539,N_585);
or U1641 (N_1641,N_120,N_221);
xnor U1642 (N_1642,N_762,N_930);
xor U1643 (N_1643,N_669,N_549);
or U1644 (N_1644,N_324,N_396);
nand U1645 (N_1645,N_454,N_191);
or U1646 (N_1646,N_347,N_661);
nor U1647 (N_1647,N_299,N_861);
nand U1648 (N_1648,N_677,N_16);
nand U1649 (N_1649,N_170,N_517);
nand U1650 (N_1650,N_433,N_428);
nand U1651 (N_1651,N_214,N_692);
or U1652 (N_1652,N_430,N_991);
xor U1653 (N_1653,N_574,N_565);
and U1654 (N_1654,N_345,N_8);
nor U1655 (N_1655,N_469,N_717);
and U1656 (N_1656,N_353,N_109);
or U1657 (N_1657,N_354,N_642);
xor U1658 (N_1658,N_747,N_219);
nand U1659 (N_1659,N_629,N_928);
nand U1660 (N_1660,N_239,N_295);
nand U1661 (N_1661,N_906,N_310);
or U1662 (N_1662,N_539,N_359);
or U1663 (N_1663,N_90,N_437);
or U1664 (N_1664,N_552,N_524);
xnor U1665 (N_1665,N_987,N_475);
or U1666 (N_1666,N_873,N_116);
nor U1667 (N_1667,N_43,N_103);
nand U1668 (N_1668,N_264,N_665);
or U1669 (N_1669,N_433,N_593);
xnor U1670 (N_1670,N_192,N_733);
nor U1671 (N_1671,N_209,N_176);
nand U1672 (N_1672,N_344,N_88);
and U1673 (N_1673,N_730,N_737);
and U1674 (N_1674,N_338,N_986);
or U1675 (N_1675,N_449,N_391);
nand U1676 (N_1676,N_720,N_173);
xor U1677 (N_1677,N_391,N_627);
xor U1678 (N_1678,N_916,N_713);
xnor U1679 (N_1679,N_640,N_515);
xor U1680 (N_1680,N_249,N_283);
nor U1681 (N_1681,N_877,N_453);
nor U1682 (N_1682,N_658,N_278);
xnor U1683 (N_1683,N_617,N_812);
and U1684 (N_1684,N_991,N_27);
nor U1685 (N_1685,N_77,N_541);
or U1686 (N_1686,N_372,N_874);
nor U1687 (N_1687,N_639,N_331);
nand U1688 (N_1688,N_822,N_973);
and U1689 (N_1689,N_375,N_416);
nand U1690 (N_1690,N_302,N_186);
and U1691 (N_1691,N_135,N_61);
nand U1692 (N_1692,N_498,N_113);
nor U1693 (N_1693,N_561,N_162);
xnor U1694 (N_1694,N_737,N_175);
nand U1695 (N_1695,N_162,N_710);
xnor U1696 (N_1696,N_55,N_47);
nand U1697 (N_1697,N_226,N_69);
xor U1698 (N_1698,N_616,N_146);
nand U1699 (N_1699,N_681,N_321);
or U1700 (N_1700,N_801,N_880);
nand U1701 (N_1701,N_483,N_841);
xnor U1702 (N_1702,N_66,N_619);
xor U1703 (N_1703,N_717,N_890);
xnor U1704 (N_1704,N_265,N_964);
xor U1705 (N_1705,N_265,N_536);
or U1706 (N_1706,N_906,N_924);
xor U1707 (N_1707,N_680,N_235);
nand U1708 (N_1708,N_607,N_172);
or U1709 (N_1709,N_395,N_657);
xnor U1710 (N_1710,N_41,N_699);
xnor U1711 (N_1711,N_881,N_566);
and U1712 (N_1712,N_580,N_689);
nor U1713 (N_1713,N_948,N_536);
nand U1714 (N_1714,N_481,N_592);
or U1715 (N_1715,N_106,N_708);
xor U1716 (N_1716,N_731,N_61);
and U1717 (N_1717,N_491,N_931);
nand U1718 (N_1718,N_334,N_969);
nor U1719 (N_1719,N_507,N_202);
nand U1720 (N_1720,N_847,N_255);
nor U1721 (N_1721,N_700,N_28);
and U1722 (N_1722,N_522,N_256);
xnor U1723 (N_1723,N_998,N_198);
xnor U1724 (N_1724,N_384,N_179);
or U1725 (N_1725,N_904,N_950);
nand U1726 (N_1726,N_803,N_655);
nand U1727 (N_1727,N_898,N_551);
and U1728 (N_1728,N_282,N_354);
nand U1729 (N_1729,N_477,N_434);
and U1730 (N_1730,N_763,N_579);
and U1731 (N_1731,N_416,N_437);
and U1732 (N_1732,N_266,N_260);
nand U1733 (N_1733,N_26,N_223);
or U1734 (N_1734,N_987,N_68);
and U1735 (N_1735,N_952,N_931);
xnor U1736 (N_1736,N_514,N_228);
nand U1737 (N_1737,N_896,N_209);
nor U1738 (N_1738,N_520,N_704);
nor U1739 (N_1739,N_206,N_97);
and U1740 (N_1740,N_774,N_8);
xor U1741 (N_1741,N_396,N_890);
or U1742 (N_1742,N_621,N_654);
nand U1743 (N_1743,N_101,N_952);
xnor U1744 (N_1744,N_926,N_987);
nand U1745 (N_1745,N_472,N_586);
xor U1746 (N_1746,N_170,N_34);
and U1747 (N_1747,N_740,N_153);
or U1748 (N_1748,N_257,N_315);
and U1749 (N_1749,N_577,N_590);
or U1750 (N_1750,N_281,N_919);
and U1751 (N_1751,N_790,N_223);
or U1752 (N_1752,N_880,N_267);
nor U1753 (N_1753,N_964,N_177);
nor U1754 (N_1754,N_445,N_165);
and U1755 (N_1755,N_499,N_516);
or U1756 (N_1756,N_347,N_990);
and U1757 (N_1757,N_452,N_627);
xor U1758 (N_1758,N_651,N_834);
or U1759 (N_1759,N_174,N_776);
nor U1760 (N_1760,N_123,N_976);
nor U1761 (N_1761,N_320,N_693);
nor U1762 (N_1762,N_486,N_146);
and U1763 (N_1763,N_40,N_199);
nand U1764 (N_1764,N_992,N_475);
and U1765 (N_1765,N_41,N_647);
nor U1766 (N_1766,N_169,N_644);
or U1767 (N_1767,N_845,N_558);
or U1768 (N_1768,N_703,N_518);
xnor U1769 (N_1769,N_271,N_201);
xor U1770 (N_1770,N_927,N_735);
xnor U1771 (N_1771,N_636,N_114);
and U1772 (N_1772,N_576,N_330);
xor U1773 (N_1773,N_991,N_9);
xnor U1774 (N_1774,N_763,N_165);
or U1775 (N_1775,N_573,N_446);
nor U1776 (N_1776,N_154,N_997);
and U1777 (N_1777,N_831,N_917);
and U1778 (N_1778,N_849,N_433);
nor U1779 (N_1779,N_606,N_363);
and U1780 (N_1780,N_499,N_142);
or U1781 (N_1781,N_673,N_727);
and U1782 (N_1782,N_143,N_547);
nor U1783 (N_1783,N_350,N_230);
or U1784 (N_1784,N_154,N_132);
xor U1785 (N_1785,N_278,N_324);
or U1786 (N_1786,N_346,N_699);
nand U1787 (N_1787,N_888,N_39);
or U1788 (N_1788,N_515,N_348);
xor U1789 (N_1789,N_289,N_850);
xor U1790 (N_1790,N_250,N_646);
or U1791 (N_1791,N_907,N_480);
and U1792 (N_1792,N_675,N_854);
and U1793 (N_1793,N_828,N_955);
and U1794 (N_1794,N_247,N_384);
xor U1795 (N_1795,N_643,N_34);
and U1796 (N_1796,N_762,N_562);
and U1797 (N_1797,N_7,N_233);
nor U1798 (N_1798,N_1,N_464);
xor U1799 (N_1799,N_232,N_791);
xor U1800 (N_1800,N_786,N_586);
nand U1801 (N_1801,N_965,N_694);
or U1802 (N_1802,N_741,N_687);
xnor U1803 (N_1803,N_900,N_271);
nand U1804 (N_1804,N_888,N_265);
and U1805 (N_1805,N_792,N_471);
or U1806 (N_1806,N_122,N_629);
or U1807 (N_1807,N_369,N_546);
or U1808 (N_1808,N_989,N_148);
or U1809 (N_1809,N_57,N_874);
xnor U1810 (N_1810,N_961,N_410);
nand U1811 (N_1811,N_253,N_350);
xnor U1812 (N_1812,N_954,N_535);
nor U1813 (N_1813,N_971,N_269);
and U1814 (N_1814,N_692,N_649);
or U1815 (N_1815,N_868,N_92);
and U1816 (N_1816,N_44,N_441);
and U1817 (N_1817,N_121,N_432);
and U1818 (N_1818,N_161,N_749);
or U1819 (N_1819,N_998,N_883);
nor U1820 (N_1820,N_400,N_919);
xnor U1821 (N_1821,N_274,N_684);
and U1822 (N_1822,N_592,N_23);
nand U1823 (N_1823,N_660,N_493);
nor U1824 (N_1824,N_663,N_21);
xor U1825 (N_1825,N_293,N_738);
nand U1826 (N_1826,N_353,N_218);
xor U1827 (N_1827,N_624,N_341);
nor U1828 (N_1828,N_896,N_539);
xnor U1829 (N_1829,N_782,N_400);
xnor U1830 (N_1830,N_790,N_338);
xnor U1831 (N_1831,N_765,N_916);
nor U1832 (N_1832,N_233,N_994);
nand U1833 (N_1833,N_818,N_742);
or U1834 (N_1834,N_759,N_783);
and U1835 (N_1835,N_972,N_363);
nor U1836 (N_1836,N_845,N_760);
nand U1837 (N_1837,N_971,N_323);
nor U1838 (N_1838,N_386,N_758);
and U1839 (N_1839,N_336,N_500);
nand U1840 (N_1840,N_274,N_146);
nand U1841 (N_1841,N_67,N_89);
or U1842 (N_1842,N_477,N_632);
nor U1843 (N_1843,N_53,N_494);
or U1844 (N_1844,N_815,N_582);
or U1845 (N_1845,N_573,N_433);
xor U1846 (N_1846,N_310,N_99);
and U1847 (N_1847,N_977,N_491);
nand U1848 (N_1848,N_63,N_75);
xor U1849 (N_1849,N_2,N_415);
xnor U1850 (N_1850,N_391,N_992);
or U1851 (N_1851,N_104,N_160);
nor U1852 (N_1852,N_54,N_804);
nand U1853 (N_1853,N_181,N_568);
nand U1854 (N_1854,N_974,N_606);
xor U1855 (N_1855,N_726,N_227);
or U1856 (N_1856,N_104,N_783);
or U1857 (N_1857,N_502,N_535);
xnor U1858 (N_1858,N_800,N_42);
and U1859 (N_1859,N_380,N_487);
or U1860 (N_1860,N_697,N_869);
xnor U1861 (N_1861,N_919,N_139);
xor U1862 (N_1862,N_741,N_968);
nand U1863 (N_1863,N_423,N_145);
and U1864 (N_1864,N_502,N_236);
nand U1865 (N_1865,N_894,N_396);
and U1866 (N_1866,N_405,N_170);
nor U1867 (N_1867,N_362,N_243);
and U1868 (N_1868,N_50,N_694);
or U1869 (N_1869,N_358,N_554);
nor U1870 (N_1870,N_327,N_541);
xor U1871 (N_1871,N_695,N_650);
or U1872 (N_1872,N_530,N_929);
xnor U1873 (N_1873,N_978,N_266);
xor U1874 (N_1874,N_607,N_231);
nor U1875 (N_1875,N_447,N_175);
nor U1876 (N_1876,N_646,N_633);
and U1877 (N_1877,N_784,N_886);
nand U1878 (N_1878,N_614,N_411);
and U1879 (N_1879,N_363,N_752);
or U1880 (N_1880,N_7,N_76);
nor U1881 (N_1881,N_704,N_667);
nand U1882 (N_1882,N_127,N_391);
or U1883 (N_1883,N_680,N_44);
nand U1884 (N_1884,N_712,N_107);
or U1885 (N_1885,N_654,N_736);
nand U1886 (N_1886,N_182,N_996);
xnor U1887 (N_1887,N_290,N_832);
nand U1888 (N_1888,N_685,N_774);
nor U1889 (N_1889,N_303,N_520);
and U1890 (N_1890,N_516,N_175);
and U1891 (N_1891,N_832,N_260);
and U1892 (N_1892,N_926,N_478);
xor U1893 (N_1893,N_900,N_579);
or U1894 (N_1894,N_138,N_571);
nor U1895 (N_1895,N_523,N_253);
xor U1896 (N_1896,N_396,N_197);
or U1897 (N_1897,N_577,N_903);
or U1898 (N_1898,N_655,N_951);
nand U1899 (N_1899,N_960,N_833);
nand U1900 (N_1900,N_466,N_254);
nor U1901 (N_1901,N_897,N_638);
and U1902 (N_1902,N_149,N_291);
nor U1903 (N_1903,N_581,N_733);
nand U1904 (N_1904,N_651,N_211);
nand U1905 (N_1905,N_194,N_216);
or U1906 (N_1906,N_855,N_805);
or U1907 (N_1907,N_669,N_198);
or U1908 (N_1908,N_115,N_216);
nor U1909 (N_1909,N_33,N_915);
nand U1910 (N_1910,N_239,N_821);
nor U1911 (N_1911,N_611,N_684);
xnor U1912 (N_1912,N_53,N_766);
and U1913 (N_1913,N_190,N_906);
nand U1914 (N_1914,N_760,N_685);
nand U1915 (N_1915,N_626,N_866);
xnor U1916 (N_1916,N_32,N_276);
nand U1917 (N_1917,N_914,N_862);
and U1918 (N_1918,N_202,N_49);
nand U1919 (N_1919,N_413,N_522);
nor U1920 (N_1920,N_91,N_724);
and U1921 (N_1921,N_371,N_131);
or U1922 (N_1922,N_97,N_342);
xnor U1923 (N_1923,N_352,N_552);
or U1924 (N_1924,N_417,N_415);
xor U1925 (N_1925,N_580,N_885);
nand U1926 (N_1926,N_837,N_369);
nand U1927 (N_1927,N_761,N_438);
or U1928 (N_1928,N_975,N_285);
nor U1929 (N_1929,N_583,N_375);
nor U1930 (N_1930,N_140,N_209);
or U1931 (N_1931,N_430,N_946);
and U1932 (N_1932,N_351,N_694);
xor U1933 (N_1933,N_994,N_421);
or U1934 (N_1934,N_582,N_69);
and U1935 (N_1935,N_110,N_452);
xnor U1936 (N_1936,N_842,N_930);
nand U1937 (N_1937,N_98,N_392);
and U1938 (N_1938,N_917,N_204);
nand U1939 (N_1939,N_39,N_720);
or U1940 (N_1940,N_202,N_240);
and U1941 (N_1941,N_866,N_138);
and U1942 (N_1942,N_354,N_849);
xnor U1943 (N_1943,N_456,N_309);
and U1944 (N_1944,N_151,N_58);
or U1945 (N_1945,N_744,N_290);
xor U1946 (N_1946,N_208,N_530);
and U1947 (N_1947,N_373,N_445);
and U1948 (N_1948,N_8,N_97);
nor U1949 (N_1949,N_997,N_202);
nor U1950 (N_1950,N_400,N_107);
or U1951 (N_1951,N_857,N_24);
and U1952 (N_1952,N_102,N_16);
nor U1953 (N_1953,N_750,N_402);
nand U1954 (N_1954,N_451,N_505);
nor U1955 (N_1955,N_54,N_68);
nor U1956 (N_1956,N_182,N_128);
xor U1957 (N_1957,N_670,N_287);
and U1958 (N_1958,N_163,N_483);
xor U1959 (N_1959,N_149,N_220);
or U1960 (N_1960,N_523,N_117);
xnor U1961 (N_1961,N_808,N_399);
xnor U1962 (N_1962,N_931,N_256);
xor U1963 (N_1963,N_888,N_765);
or U1964 (N_1964,N_617,N_435);
nor U1965 (N_1965,N_960,N_417);
or U1966 (N_1966,N_306,N_947);
nand U1967 (N_1967,N_711,N_82);
and U1968 (N_1968,N_727,N_970);
and U1969 (N_1969,N_312,N_667);
xor U1970 (N_1970,N_799,N_540);
nor U1971 (N_1971,N_194,N_91);
nand U1972 (N_1972,N_507,N_893);
or U1973 (N_1973,N_38,N_962);
or U1974 (N_1974,N_980,N_257);
or U1975 (N_1975,N_934,N_277);
and U1976 (N_1976,N_178,N_38);
nor U1977 (N_1977,N_589,N_672);
and U1978 (N_1978,N_235,N_355);
nand U1979 (N_1979,N_961,N_625);
nand U1980 (N_1980,N_780,N_703);
and U1981 (N_1981,N_541,N_878);
xor U1982 (N_1982,N_347,N_162);
nor U1983 (N_1983,N_958,N_469);
nor U1984 (N_1984,N_608,N_277);
nand U1985 (N_1985,N_330,N_152);
xnor U1986 (N_1986,N_184,N_25);
and U1987 (N_1987,N_613,N_532);
or U1988 (N_1988,N_123,N_898);
xor U1989 (N_1989,N_95,N_919);
or U1990 (N_1990,N_715,N_55);
nand U1991 (N_1991,N_909,N_524);
and U1992 (N_1992,N_743,N_90);
xnor U1993 (N_1993,N_690,N_132);
nor U1994 (N_1994,N_834,N_787);
and U1995 (N_1995,N_684,N_430);
xor U1996 (N_1996,N_644,N_597);
or U1997 (N_1997,N_728,N_196);
or U1998 (N_1998,N_15,N_647);
and U1999 (N_1999,N_5,N_599);
xor U2000 (N_2000,N_1656,N_1406);
and U2001 (N_2001,N_1454,N_1827);
nor U2002 (N_2002,N_1115,N_1931);
xnor U2003 (N_2003,N_1811,N_1308);
nand U2004 (N_2004,N_1780,N_1680);
and U2005 (N_2005,N_1280,N_1133);
nand U2006 (N_2006,N_1979,N_1694);
nor U2007 (N_2007,N_1587,N_1606);
nor U2008 (N_2008,N_1746,N_1019);
xnor U2009 (N_2009,N_1403,N_1121);
xnor U2010 (N_2010,N_1247,N_1614);
nor U2011 (N_2011,N_1268,N_1769);
nor U2012 (N_2012,N_1665,N_1547);
nor U2013 (N_2013,N_1253,N_1918);
xor U2014 (N_2014,N_1520,N_1230);
nor U2015 (N_2015,N_1279,N_1921);
or U2016 (N_2016,N_1251,N_1552);
nor U2017 (N_2017,N_1288,N_1119);
nand U2018 (N_2018,N_1296,N_1674);
nor U2019 (N_2019,N_1654,N_1319);
xor U2020 (N_2020,N_1053,N_1857);
nand U2021 (N_2021,N_1554,N_1408);
and U2022 (N_2022,N_1549,N_1417);
nand U2023 (N_2023,N_1726,N_1574);
xnor U2024 (N_2024,N_1820,N_1814);
nor U2025 (N_2025,N_1993,N_1592);
xor U2026 (N_2026,N_1607,N_1511);
nor U2027 (N_2027,N_1292,N_1977);
xnor U2028 (N_2028,N_1240,N_1492);
or U2029 (N_2029,N_1877,N_1739);
nand U2030 (N_2030,N_1781,N_1285);
nand U2031 (N_2031,N_1962,N_1476);
nor U2032 (N_2032,N_1161,N_1994);
and U2033 (N_2033,N_1947,N_1856);
nor U2034 (N_2034,N_1551,N_1736);
xnor U2035 (N_2035,N_1847,N_1721);
nor U2036 (N_2036,N_1001,N_1538);
xnor U2037 (N_2037,N_1718,N_1099);
nand U2038 (N_2038,N_1905,N_1682);
nand U2039 (N_2039,N_1495,N_1527);
nor U2040 (N_2040,N_1752,N_1205);
and U2041 (N_2041,N_1452,N_1843);
and U2042 (N_2042,N_1493,N_1088);
nand U2043 (N_2043,N_1257,N_1341);
xnor U2044 (N_2044,N_1346,N_1500);
nor U2045 (N_2045,N_1899,N_1621);
xnor U2046 (N_2046,N_1283,N_1953);
xor U2047 (N_2047,N_1920,N_1835);
or U2048 (N_2048,N_1715,N_1276);
and U2049 (N_2049,N_1955,N_1397);
nand U2050 (N_2050,N_1356,N_1686);
nand U2051 (N_2051,N_1690,N_1556);
nor U2052 (N_2052,N_1523,N_1434);
nand U2053 (N_2053,N_1627,N_1365);
nor U2054 (N_2054,N_1071,N_1139);
or U2055 (N_2055,N_1224,N_1046);
xor U2056 (N_2056,N_1405,N_1327);
or U2057 (N_2057,N_1353,N_1702);
nand U2058 (N_2058,N_1031,N_1803);
xnor U2059 (N_2059,N_1347,N_1234);
or U2060 (N_2060,N_1098,N_1060);
and U2061 (N_2061,N_1944,N_1613);
nor U2062 (N_2062,N_1532,N_1915);
or U2063 (N_2063,N_1582,N_1516);
nor U2064 (N_2064,N_1440,N_1713);
and U2065 (N_2065,N_1132,N_1318);
nor U2066 (N_2066,N_1841,N_1398);
nor U2067 (N_2067,N_1553,N_1072);
or U2068 (N_2068,N_1591,N_1764);
nor U2069 (N_2069,N_1120,N_1522);
nand U2070 (N_2070,N_1583,N_1174);
nand U2071 (N_2071,N_1533,N_1354);
xnor U2072 (N_2072,N_1943,N_1964);
xnor U2073 (N_2073,N_1800,N_1449);
nand U2074 (N_2074,N_1488,N_1238);
or U2075 (N_2075,N_1608,N_1486);
nor U2076 (N_2076,N_1630,N_1033);
xnor U2077 (N_2077,N_1442,N_1489);
nand U2078 (N_2078,N_1887,N_1952);
or U2079 (N_2079,N_1422,N_1469);
xor U2080 (N_2080,N_1380,N_1287);
or U2081 (N_2081,N_1661,N_1647);
and U2082 (N_2082,N_1300,N_1501);
or U2083 (N_2083,N_1368,N_1535);
nor U2084 (N_2084,N_1753,N_1640);
or U2085 (N_2085,N_1124,N_1762);
or U2086 (N_2086,N_1242,N_1867);
xor U2087 (N_2087,N_1540,N_1266);
nand U2088 (N_2088,N_1672,N_1770);
nand U2089 (N_2089,N_1151,N_1685);
and U2090 (N_2090,N_1515,N_1704);
and U2091 (N_2091,N_1941,N_1536);
nor U2092 (N_2092,N_1696,N_1277);
and U2093 (N_2093,N_1055,N_1080);
and U2094 (N_2094,N_1435,N_1975);
or U2095 (N_2095,N_1106,N_1874);
or U2096 (N_2096,N_1044,N_1963);
and U2097 (N_2097,N_1334,N_1862);
xnor U2098 (N_2098,N_1426,N_1503);
or U2099 (N_2099,N_1840,N_1385);
nor U2100 (N_2100,N_1624,N_1725);
and U2101 (N_2101,N_1004,N_1262);
or U2102 (N_2102,N_1249,N_1643);
nor U2103 (N_2103,N_1982,N_1082);
nor U2104 (N_2104,N_1997,N_1719);
xnor U2105 (N_2105,N_1797,N_1872);
nand U2106 (N_2106,N_1037,N_1147);
xor U2107 (N_2107,N_1271,N_1017);
nor U2108 (N_2108,N_1616,N_1988);
nand U2109 (N_2109,N_1441,N_1322);
xor U2110 (N_2110,N_1411,N_1415);
nor U2111 (N_2111,N_1848,N_1779);
xnor U2112 (N_2112,N_1926,N_1504);
and U2113 (N_2113,N_1444,N_1573);
xor U2114 (N_2114,N_1377,N_1076);
and U2115 (N_2115,N_1039,N_1577);
nor U2116 (N_2116,N_1569,N_1785);
and U2117 (N_2117,N_1360,N_1371);
or U2118 (N_2118,N_1073,N_1178);
and U2119 (N_2119,N_1973,N_1819);
and U2120 (N_2120,N_1677,N_1628);
nor U2121 (N_2121,N_1555,N_1974);
nor U2122 (N_2122,N_1667,N_1480);
or U2123 (N_2123,N_1231,N_1138);
xor U2124 (N_2124,N_1127,N_1061);
or U2125 (N_2125,N_1909,N_1730);
xnor U2126 (N_2126,N_1565,N_1419);
xnor U2127 (N_2127,N_1064,N_1557);
nor U2128 (N_2128,N_1485,N_1859);
xor U2129 (N_2129,N_1002,N_1875);
and U2130 (N_2130,N_1381,N_1866);
and U2131 (N_2131,N_1722,N_1293);
nor U2132 (N_2132,N_1016,N_1650);
xnor U2133 (N_2133,N_1747,N_1250);
xnor U2134 (N_2134,N_1939,N_1237);
and U2135 (N_2135,N_1390,N_1423);
nor U2136 (N_2136,N_1641,N_1833);
or U2137 (N_2137,N_1842,N_1898);
xnor U2138 (N_2138,N_1144,N_1471);
or U2139 (N_2139,N_1030,N_1883);
xor U2140 (N_2140,N_1946,N_1938);
nor U2141 (N_2141,N_1707,N_1258);
xor U2142 (N_2142,N_1684,N_1585);
xor U2143 (N_2143,N_1675,N_1945);
and U2144 (N_2144,N_1891,N_1387);
nor U2145 (N_2145,N_1999,N_1396);
nor U2146 (N_2146,N_1078,N_1756);
or U2147 (N_2147,N_1427,N_1281);
nor U2148 (N_2148,N_1546,N_1529);
and U2149 (N_2149,N_1373,N_1933);
xnor U2150 (N_2150,N_1812,N_1671);
nor U2151 (N_2151,N_1084,N_1468);
nor U2152 (N_2152,N_1225,N_1462);
nor U2153 (N_2153,N_1185,N_1751);
nand U2154 (N_2154,N_1761,N_1418);
or U2155 (N_2155,N_1776,N_1210);
and U2156 (N_2156,N_1709,N_1626);
and U2157 (N_2157,N_1652,N_1095);
nand U2158 (N_2158,N_1111,N_1141);
or U2159 (N_2159,N_1777,N_1359);
or U2160 (N_2160,N_1186,N_1985);
or U2161 (N_2161,N_1143,N_1213);
or U2162 (N_2162,N_1267,N_1497);
nor U2163 (N_2163,N_1733,N_1109);
xnor U2164 (N_2164,N_1050,N_1731);
xnor U2165 (N_2165,N_1393,N_1865);
xor U2166 (N_2166,N_1517,N_1090);
nor U2167 (N_2167,N_1871,N_1011);
or U2168 (N_2168,N_1303,N_1639);
and U2169 (N_2169,N_1789,N_1101);
xor U2170 (N_2170,N_1611,N_1742);
nand U2171 (N_2171,N_1294,N_1734);
and U2172 (N_2172,N_1135,N_1560);
or U2173 (N_2173,N_1760,N_1670);
and U2174 (N_2174,N_1934,N_1623);
and U2175 (N_2175,N_1765,N_1226);
or U2176 (N_2176,N_1459,N_1888);
and U2177 (N_2177,N_1420,N_1792);
and U2178 (N_2178,N_1983,N_1333);
or U2179 (N_2179,N_1919,N_1207);
xnor U2180 (N_2180,N_1625,N_1136);
nand U2181 (N_2181,N_1683,N_1311);
nor U2182 (N_2182,N_1309,N_1648);
xnor U2183 (N_2183,N_1023,N_1732);
and U2184 (N_2184,N_1506,N_1846);
or U2185 (N_2185,N_1027,N_1711);
nand U2186 (N_2186,N_1007,N_1069);
nor U2187 (N_2187,N_1180,N_1911);
nor U2188 (N_2188,N_1150,N_1477);
nor U2189 (N_2189,N_1163,N_1507);
nand U2190 (N_2190,N_1622,N_1048);
and U2191 (N_2191,N_1313,N_1113);
and U2192 (N_2192,N_1458,N_1110);
xnor U2193 (N_2193,N_1474,N_1935);
nor U2194 (N_2194,N_1208,N_1096);
xnor U2195 (N_2195,N_1496,N_1345);
and U2196 (N_2196,N_1603,N_1357);
xnor U2197 (N_2197,N_1633,N_1996);
and U2198 (N_2198,N_1595,N_1687);
or U2199 (N_2199,N_1085,N_1173);
xor U2200 (N_2200,N_1914,N_1352);
nor U2201 (N_2201,N_1699,N_1028);
xnor U2202 (N_2202,N_1724,N_1448);
xor U2203 (N_2203,N_1404,N_1457);
nand U2204 (N_2204,N_1837,N_1508);
nor U2205 (N_2205,N_1058,N_1669);
and U2206 (N_2206,N_1394,N_1787);
nor U2207 (N_2207,N_1430,N_1968);
nor U2208 (N_2208,N_1818,N_1370);
and U2209 (N_2209,N_1245,N_1763);
and U2210 (N_2210,N_1395,N_1826);
nor U2211 (N_2211,N_1563,N_1233);
and U2212 (N_2212,N_1428,N_1530);
nor U2213 (N_2213,N_1059,N_1297);
nand U2214 (N_2214,N_1122,N_1832);
nor U2215 (N_2215,N_1668,N_1291);
xnor U2216 (N_2216,N_1216,N_1793);
nor U2217 (N_2217,N_1795,N_1666);
xor U2218 (N_2218,N_1321,N_1984);
nor U2219 (N_2219,N_1617,N_1158);
or U2220 (N_2220,N_1681,N_1343);
and U2221 (N_2221,N_1850,N_1260);
nand U2222 (N_2222,N_1204,N_1490);
or U2223 (N_2223,N_1367,N_1118);
and U2224 (N_2224,N_1328,N_1013);
or U2225 (N_2225,N_1052,N_1706);
xor U2226 (N_2226,N_1550,N_1065);
and U2227 (N_2227,N_1881,N_1882);
and U2228 (N_2228,N_1439,N_1264);
or U2229 (N_2229,N_1599,N_1727);
or U2230 (N_2230,N_1068,N_1600);
nor U2231 (N_2231,N_1384,N_1810);
or U2232 (N_2232,N_1586,N_1214);
and U2233 (N_2233,N_1917,N_1539);
nand U2234 (N_2234,N_1924,N_1310);
or U2235 (N_2235,N_1544,N_1342);
nor U2236 (N_2236,N_1339,N_1852);
xnor U2237 (N_2237,N_1584,N_1610);
nor U2238 (N_2238,N_1154,N_1851);
nor U2239 (N_2239,N_1482,N_1438);
or U2240 (N_2240,N_1298,N_1189);
xor U2241 (N_2241,N_1137,N_1460);
or U2242 (N_2242,N_1379,N_1534);
or U2243 (N_2243,N_1894,N_1079);
or U2244 (N_2244,N_1971,N_1992);
nand U2245 (N_2245,N_1104,N_1995);
xor U2246 (N_2246,N_1041,N_1366);
nand U2247 (N_2247,N_1491,N_1807);
or U2248 (N_2248,N_1908,N_1304);
nor U2249 (N_2249,N_1796,N_1700);
nand U2250 (N_2250,N_1558,N_1604);
nor U2251 (N_2251,N_1155,N_1749);
nand U2252 (N_2252,N_1126,N_1056);
xor U2253 (N_2253,N_1658,N_1937);
nor U2254 (N_2254,N_1043,N_1103);
and U2255 (N_2255,N_1597,N_1657);
nor U2256 (N_2256,N_1940,N_1618);
nand U2257 (N_2257,N_1854,N_1767);
and U2258 (N_2258,N_1102,N_1615);
or U2259 (N_2259,N_1897,N_1369);
nor U2260 (N_2260,N_1223,N_1593);
nor U2261 (N_2261,N_1801,N_1688);
and U2262 (N_2262,N_1701,N_1198);
nand U2263 (N_2263,N_1128,N_1412);
nor U2264 (N_2264,N_1086,N_1958);
and U2265 (N_2265,N_1105,N_1246);
nor U2266 (N_2266,N_1083,N_1487);
xor U2267 (N_2267,N_1235,N_1049);
and U2268 (N_2268,N_1703,N_1956);
xnor U2269 (N_2269,N_1416,N_1159);
and U2270 (N_2270,N_1192,N_1187);
nand U2271 (N_2271,N_1097,N_1024);
xor U2272 (N_2272,N_1239,N_1986);
nor U2273 (N_2273,N_1087,N_1164);
nand U2274 (N_2274,N_1320,N_1382);
xor U2275 (N_2275,N_1123,N_1890);
nand U2276 (N_2276,N_1817,N_1008);
nor U2277 (N_2277,N_1316,N_1717);
nor U2278 (N_2278,N_1631,N_1160);
and U2279 (N_2279,N_1930,N_1182);
nand U2280 (N_2280,N_1860,N_1579);
or U2281 (N_2281,N_1012,N_1870);
nand U2282 (N_2282,N_1275,N_1619);
nor U2283 (N_2283,N_1548,N_1748);
nor U2284 (N_2284,N_1289,N_1849);
nand U2285 (N_2285,N_1823,N_1601);
nand U2286 (N_2286,N_1564,N_1567);
xor U2287 (N_2287,N_1910,N_1340);
nand U2288 (N_2288,N_1399,N_1094);
xnor U2289 (N_2289,N_1673,N_1199);
nor U2290 (N_2290,N_1323,N_1358);
or U2291 (N_2291,N_1450,N_1838);
and U2292 (N_2292,N_1000,N_1301);
nand U2293 (N_2293,N_1831,N_1034);
or U2294 (N_2294,N_1171,N_1759);
and U2295 (N_2295,N_1157,N_1219);
and U2296 (N_2296,N_1580,N_1659);
nand U2297 (N_2297,N_1217,N_1954);
xor U2298 (N_2298,N_1433,N_1662);
or U2299 (N_2299,N_1282,N_1168);
nand U2300 (N_2300,N_1645,N_1806);
nor U2301 (N_2301,N_1772,N_1927);
nand U2302 (N_2302,N_1032,N_1998);
xnor U2303 (N_2303,N_1775,N_1453);
xnor U2304 (N_2304,N_1502,N_1828);
nand U2305 (N_2305,N_1542,N_1197);
xor U2306 (N_2306,N_1483,N_1864);
or U2307 (N_2307,N_1757,N_1651);
or U2308 (N_2308,N_1844,N_1895);
and U2309 (N_2309,N_1075,N_1465);
or U2310 (N_2310,N_1009,N_1255);
and U2311 (N_2311,N_1689,N_1218);
nand U2312 (N_2312,N_1922,N_1456);
nand U2313 (N_2313,N_1788,N_1350);
and U2314 (N_2314,N_1620,N_1655);
or U2315 (N_2315,N_1773,N_1609);
nor U2316 (N_2316,N_1388,N_1286);
and U2317 (N_2317,N_1712,N_1195);
and U2318 (N_2318,N_1912,N_1472);
xor U2319 (N_2319,N_1066,N_1829);
and U2320 (N_2320,N_1274,N_1499);
nor U2321 (N_2321,N_1798,N_1879);
xnor U2322 (N_2322,N_1146,N_1220);
and U2323 (N_2323,N_1206,N_1928);
nor U2324 (N_2324,N_1265,N_1913);
nand U2325 (N_2325,N_1808,N_1885);
and U2326 (N_2326,N_1355,N_1990);
nor U2327 (N_2327,N_1351,N_1421);
or U2328 (N_2328,N_1960,N_1077);
xor U2329 (N_2329,N_1446,N_1424);
nand U2330 (N_2330,N_1447,N_1642);
or U2331 (N_2331,N_1152,N_1167);
nor U2332 (N_2332,N_1413,N_1475);
or U2333 (N_2333,N_1570,N_1302);
or U2334 (N_2334,N_1392,N_1589);
nand U2335 (N_2335,N_1822,N_1410);
or U2336 (N_2336,N_1705,N_1295);
and U2337 (N_2337,N_1526,N_1525);
nand U2338 (N_2338,N_1716,N_1362);
xnor U2339 (N_2339,N_1203,N_1378);
xor U2340 (N_2340,N_1566,N_1400);
and U2341 (N_2341,N_1873,N_1966);
nor U2342 (N_2342,N_1816,N_1653);
nand U2343 (N_2343,N_1695,N_1825);
nand U2344 (N_2344,N_1431,N_1855);
or U2345 (N_2345,N_1660,N_1256);
and U2346 (N_2346,N_1054,N_1679);
xor U2347 (N_2347,N_1375,N_1980);
nor U2348 (N_2348,N_1270,N_1212);
and U2349 (N_2349,N_1878,N_1361);
xnor U2350 (N_2350,N_1402,N_1884);
nand U2351 (N_2351,N_1042,N_1594);
nand U2352 (N_2352,N_1228,N_1272);
nand U2353 (N_2353,N_1035,N_1510);
xnor U2354 (N_2354,N_1783,N_1741);
and U2355 (N_2355,N_1602,N_1259);
nand U2356 (N_2356,N_1047,N_1081);
nand U2357 (N_2357,N_1886,N_1758);
xor U2358 (N_2358,N_1177,N_1575);
xor U2359 (N_2359,N_1129,N_1802);
nand U2360 (N_2360,N_1443,N_1211);
nand U2361 (N_2361,N_1693,N_1581);
or U2362 (N_2362,N_1559,N_1463);
or U2363 (N_2363,N_1200,N_1142);
and U2364 (N_2364,N_1750,N_1903);
xor U2365 (N_2365,N_1170,N_1074);
nand U2366 (N_2366,N_1172,N_1194);
nor U2367 (N_2367,N_1755,N_1509);
nor U2368 (N_2368,N_1470,N_1970);
or U2369 (N_2369,N_1543,N_1524);
xnor U2370 (N_2370,N_1790,N_1331);
and U2371 (N_2371,N_1202,N_1692);
or U2372 (N_2372,N_1436,N_1227);
xnor U2373 (N_2373,N_1005,N_1455);
or U2374 (N_2374,N_1479,N_1232);
and U2375 (N_2375,N_1188,N_1710);
and U2376 (N_2376,N_1728,N_1307);
nand U2377 (N_2377,N_1432,N_1698);
and U2378 (N_2378,N_1830,N_1338);
nand U2379 (N_2379,N_1987,N_1166);
nand U2380 (N_2380,N_1794,N_1858);
xnor U2381 (N_2381,N_1335,N_1176);
nor U2382 (N_2382,N_1637,N_1744);
and U2383 (N_2383,N_1799,N_1605);
or U2384 (N_2384,N_1782,N_1902);
nor U2385 (N_2385,N_1743,N_1805);
or U2386 (N_2386,N_1116,N_1429);
nand U2387 (N_2387,N_1386,N_1063);
nor U2388 (N_2388,N_1383,N_1089);
nand U2389 (N_2389,N_1766,N_1596);
nand U2390 (N_2390,N_1804,N_1942);
nand U2391 (N_2391,N_1969,N_1821);
xnor U2392 (N_2392,N_1664,N_1261);
nor U2393 (N_2393,N_1678,N_1332);
and U2394 (N_2394,N_1248,N_1029);
nand U2395 (N_2395,N_1519,N_1401);
and U2396 (N_2396,N_1907,N_1572);
nand U2397 (N_2397,N_1140,N_1349);
or U2398 (N_2398,N_1815,N_1134);
or U2399 (N_2399,N_1976,N_1901);
xor U2400 (N_2400,N_1464,N_1863);
or U2401 (N_2401,N_1892,N_1169);
nor U2402 (N_2402,N_1473,N_1117);
or U2403 (N_2403,N_1252,N_1568);
and U2404 (N_2404,N_1461,N_1254);
xor U2405 (N_2405,N_1598,N_1363);
nand U2406 (N_2406,N_1108,N_1092);
and U2407 (N_2407,N_1959,N_1932);
nor U2408 (N_2408,N_1513,N_1179);
and U2409 (N_2409,N_1478,N_1175);
xnor U2410 (N_2410,N_1876,N_1845);
nand U2411 (N_2411,N_1512,N_1051);
or U2412 (N_2412,N_1861,N_1229);
nor U2413 (N_2413,N_1125,N_1484);
and U2414 (N_2414,N_1003,N_1181);
nand U2415 (N_2415,N_1191,N_1326);
and U2416 (N_2416,N_1305,N_1541);
nand U2417 (N_2417,N_1222,N_1244);
or U2418 (N_2418,N_1561,N_1278);
xor U2419 (N_2419,N_1376,N_1676);
nand U2420 (N_2420,N_1720,N_1834);
nand U2421 (N_2421,N_1091,N_1778);
or U2422 (N_2422,N_1026,N_1950);
nor U2423 (N_2423,N_1306,N_1588);
xor U2424 (N_2424,N_1936,N_1112);
nand U2425 (N_2425,N_1972,N_1562);
xnor U2426 (N_2426,N_1889,N_1010);
nor U2427 (N_2427,N_1221,N_1153);
nor U2428 (N_2428,N_1638,N_1494);
or U2429 (N_2429,N_1317,N_1344);
and U2430 (N_2430,N_1531,N_1337);
or U2431 (N_2431,N_1330,N_1273);
xor U2432 (N_2432,N_1312,N_1768);
and U2433 (N_2433,N_1951,N_1284);
nand U2434 (N_2434,N_1040,N_1269);
or U2435 (N_2435,N_1190,N_1498);
and U2436 (N_2436,N_1737,N_1067);
xor U2437 (N_2437,N_1021,N_1038);
nand U2438 (N_2438,N_1925,N_1967);
or U2439 (N_2439,N_1697,N_1636);
or U2440 (N_2440,N_1131,N_1576);
nor U2441 (N_2441,N_1149,N_1578);
nor U2442 (N_2442,N_1114,N_1634);
or U2443 (N_2443,N_1893,N_1853);
xor U2444 (N_2444,N_1193,N_1505);
nor U2445 (N_2445,N_1374,N_1336);
or U2446 (N_2446,N_1991,N_1771);
or U2447 (N_2447,N_1045,N_1391);
or U2448 (N_2448,N_1836,N_1612);
or U2449 (N_2449,N_1629,N_1521);
nor U2450 (N_2450,N_1738,N_1314);
nor U2451 (N_2451,N_1545,N_1329);
or U2452 (N_2452,N_1735,N_1929);
and U2453 (N_2453,N_1324,N_1372);
and U2454 (N_2454,N_1644,N_1014);
xnor U2455 (N_2455,N_1691,N_1481);
xor U2456 (N_2456,N_1467,N_1466);
nor U2457 (N_2457,N_1107,N_1437);
xnor U2458 (N_2458,N_1791,N_1745);
or U2459 (N_2459,N_1263,N_1906);
or U2460 (N_2460,N_1900,N_1209);
nand U2461 (N_2461,N_1740,N_1528);
xor U2462 (N_2462,N_1299,N_1425);
nand U2463 (N_2463,N_1325,N_1407);
or U2464 (N_2464,N_1348,N_1057);
or U2465 (N_2465,N_1916,N_1869);
and U2466 (N_2466,N_1130,N_1965);
nor U2467 (N_2467,N_1948,N_1215);
nor U2468 (N_2468,N_1784,N_1020);
xnor U2469 (N_2469,N_1880,N_1590);
and U2470 (N_2470,N_1236,N_1241);
or U2471 (N_2471,N_1514,N_1015);
and U2472 (N_2472,N_1813,N_1754);
nor U2473 (N_2473,N_1290,N_1809);
nor U2474 (N_2474,N_1409,N_1646);
and U2475 (N_2475,N_1018,N_1989);
and U2476 (N_2476,N_1949,N_1839);
nor U2477 (N_2477,N_1070,N_1571);
and U2478 (N_2478,N_1315,N_1389);
xor U2479 (N_2479,N_1445,N_1184);
or U2480 (N_2480,N_1036,N_1148);
nand U2481 (N_2481,N_1162,N_1786);
xnor U2482 (N_2482,N_1414,N_1100);
xor U2483 (N_2483,N_1062,N_1708);
xnor U2484 (N_2484,N_1451,N_1978);
nor U2485 (N_2485,N_1145,N_1156);
or U2486 (N_2486,N_1961,N_1729);
xor U2487 (N_2487,N_1714,N_1868);
nor U2488 (N_2488,N_1774,N_1957);
nor U2489 (N_2489,N_1243,N_1904);
nor U2490 (N_2490,N_1896,N_1649);
or U2491 (N_2491,N_1923,N_1632);
and U2492 (N_2492,N_1165,N_1025);
xor U2493 (N_2493,N_1518,N_1183);
nand U2494 (N_2494,N_1364,N_1196);
nor U2495 (N_2495,N_1537,N_1824);
xor U2496 (N_2496,N_1201,N_1093);
xor U2497 (N_2497,N_1635,N_1723);
nand U2498 (N_2498,N_1663,N_1981);
or U2499 (N_2499,N_1022,N_1006);
or U2500 (N_2500,N_1779,N_1553);
nand U2501 (N_2501,N_1177,N_1976);
xnor U2502 (N_2502,N_1302,N_1717);
nor U2503 (N_2503,N_1003,N_1507);
or U2504 (N_2504,N_1999,N_1618);
nand U2505 (N_2505,N_1638,N_1753);
and U2506 (N_2506,N_1544,N_1043);
xor U2507 (N_2507,N_1998,N_1492);
nand U2508 (N_2508,N_1733,N_1555);
or U2509 (N_2509,N_1599,N_1232);
nor U2510 (N_2510,N_1327,N_1066);
or U2511 (N_2511,N_1721,N_1132);
nand U2512 (N_2512,N_1077,N_1337);
nand U2513 (N_2513,N_1483,N_1923);
and U2514 (N_2514,N_1873,N_1019);
or U2515 (N_2515,N_1462,N_1141);
or U2516 (N_2516,N_1339,N_1404);
nand U2517 (N_2517,N_1769,N_1930);
xnor U2518 (N_2518,N_1257,N_1584);
and U2519 (N_2519,N_1411,N_1663);
nor U2520 (N_2520,N_1589,N_1970);
nand U2521 (N_2521,N_1843,N_1390);
nor U2522 (N_2522,N_1507,N_1013);
xnor U2523 (N_2523,N_1815,N_1874);
or U2524 (N_2524,N_1033,N_1182);
nand U2525 (N_2525,N_1135,N_1902);
and U2526 (N_2526,N_1800,N_1157);
and U2527 (N_2527,N_1430,N_1118);
xnor U2528 (N_2528,N_1439,N_1575);
nand U2529 (N_2529,N_1258,N_1175);
or U2530 (N_2530,N_1548,N_1945);
xor U2531 (N_2531,N_1344,N_1081);
xnor U2532 (N_2532,N_1292,N_1434);
and U2533 (N_2533,N_1331,N_1673);
nor U2534 (N_2534,N_1932,N_1550);
xnor U2535 (N_2535,N_1311,N_1044);
or U2536 (N_2536,N_1112,N_1305);
xnor U2537 (N_2537,N_1745,N_1362);
nand U2538 (N_2538,N_1582,N_1774);
and U2539 (N_2539,N_1460,N_1759);
xnor U2540 (N_2540,N_1989,N_1973);
nand U2541 (N_2541,N_1473,N_1349);
or U2542 (N_2542,N_1770,N_1966);
nand U2543 (N_2543,N_1039,N_1883);
or U2544 (N_2544,N_1583,N_1119);
xor U2545 (N_2545,N_1028,N_1377);
nand U2546 (N_2546,N_1850,N_1158);
nor U2547 (N_2547,N_1052,N_1929);
or U2548 (N_2548,N_1645,N_1608);
xnor U2549 (N_2549,N_1969,N_1595);
xnor U2550 (N_2550,N_1139,N_1368);
xnor U2551 (N_2551,N_1672,N_1079);
and U2552 (N_2552,N_1739,N_1715);
nand U2553 (N_2553,N_1873,N_1437);
nor U2554 (N_2554,N_1525,N_1412);
nor U2555 (N_2555,N_1381,N_1971);
or U2556 (N_2556,N_1688,N_1946);
or U2557 (N_2557,N_1279,N_1695);
or U2558 (N_2558,N_1457,N_1809);
or U2559 (N_2559,N_1387,N_1822);
nor U2560 (N_2560,N_1824,N_1080);
or U2561 (N_2561,N_1594,N_1567);
nand U2562 (N_2562,N_1789,N_1923);
xnor U2563 (N_2563,N_1027,N_1713);
nand U2564 (N_2564,N_1864,N_1616);
and U2565 (N_2565,N_1844,N_1663);
nand U2566 (N_2566,N_1633,N_1052);
and U2567 (N_2567,N_1935,N_1810);
and U2568 (N_2568,N_1198,N_1460);
nor U2569 (N_2569,N_1439,N_1951);
nand U2570 (N_2570,N_1764,N_1523);
nor U2571 (N_2571,N_1533,N_1981);
nand U2572 (N_2572,N_1288,N_1050);
and U2573 (N_2573,N_1519,N_1665);
nand U2574 (N_2574,N_1656,N_1088);
nand U2575 (N_2575,N_1083,N_1079);
and U2576 (N_2576,N_1358,N_1447);
or U2577 (N_2577,N_1497,N_1001);
xnor U2578 (N_2578,N_1966,N_1412);
and U2579 (N_2579,N_1752,N_1476);
nand U2580 (N_2580,N_1174,N_1222);
or U2581 (N_2581,N_1452,N_1368);
xor U2582 (N_2582,N_1673,N_1460);
or U2583 (N_2583,N_1732,N_1181);
nand U2584 (N_2584,N_1442,N_1439);
and U2585 (N_2585,N_1593,N_1748);
xor U2586 (N_2586,N_1341,N_1176);
nand U2587 (N_2587,N_1800,N_1518);
nor U2588 (N_2588,N_1878,N_1338);
and U2589 (N_2589,N_1880,N_1576);
xnor U2590 (N_2590,N_1819,N_1116);
nor U2591 (N_2591,N_1887,N_1149);
xor U2592 (N_2592,N_1282,N_1335);
xor U2593 (N_2593,N_1514,N_1140);
or U2594 (N_2594,N_1649,N_1638);
and U2595 (N_2595,N_1509,N_1218);
and U2596 (N_2596,N_1023,N_1151);
xnor U2597 (N_2597,N_1287,N_1739);
and U2598 (N_2598,N_1970,N_1797);
and U2599 (N_2599,N_1960,N_1066);
nor U2600 (N_2600,N_1567,N_1503);
xor U2601 (N_2601,N_1488,N_1306);
and U2602 (N_2602,N_1123,N_1267);
nand U2603 (N_2603,N_1167,N_1711);
and U2604 (N_2604,N_1887,N_1530);
and U2605 (N_2605,N_1349,N_1701);
or U2606 (N_2606,N_1133,N_1858);
and U2607 (N_2607,N_1543,N_1754);
nor U2608 (N_2608,N_1015,N_1165);
nand U2609 (N_2609,N_1331,N_1391);
or U2610 (N_2610,N_1482,N_1551);
nand U2611 (N_2611,N_1047,N_1751);
and U2612 (N_2612,N_1033,N_1457);
and U2613 (N_2613,N_1482,N_1299);
nor U2614 (N_2614,N_1957,N_1493);
nor U2615 (N_2615,N_1480,N_1849);
nand U2616 (N_2616,N_1494,N_1315);
nor U2617 (N_2617,N_1463,N_1009);
xnor U2618 (N_2618,N_1939,N_1465);
xor U2619 (N_2619,N_1212,N_1588);
nor U2620 (N_2620,N_1872,N_1236);
nand U2621 (N_2621,N_1809,N_1129);
and U2622 (N_2622,N_1752,N_1589);
or U2623 (N_2623,N_1325,N_1155);
or U2624 (N_2624,N_1341,N_1907);
or U2625 (N_2625,N_1664,N_1060);
and U2626 (N_2626,N_1954,N_1877);
nor U2627 (N_2627,N_1143,N_1597);
nand U2628 (N_2628,N_1771,N_1644);
nor U2629 (N_2629,N_1144,N_1367);
and U2630 (N_2630,N_1905,N_1770);
xor U2631 (N_2631,N_1529,N_1930);
and U2632 (N_2632,N_1479,N_1052);
or U2633 (N_2633,N_1890,N_1024);
xnor U2634 (N_2634,N_1290,N_1192);
and U2635 (N_2635,N_1227,N_1447);
xnor U2636 (N_2636,N_1612,N_1897);
nor U2637 (N_2637,N_1246,N_1173);
and U2638 (N_2638,N_1394,N_1908);
or U2639 (N_2639,N_1934,N_1756);
nand U2640 (N_2640,N_1984,N_1815);
or U2641 (N_2641,N_1498,N_1532);
nand U2642 (N_2642,N_1594,N_1226);
nand U2643 (N_2643,N_1265,N_1747);
and U2644 (N_2644,N_1579,N_1011);
or U2645 (N_2645,N_1131,N_1953);
or U2646 (N_2646,N_1675,N_1935);
xnor U2647 (N_2647,N_1461,N_1776);
nor U2648 (N_2648,N_1480,N_1535);
and U2649 (N_2649,N_1357,N_1084);
nor U2650 (N_2650,N_1752,N_1532);
or U2651 (N_2651,N_1857,N_1736);
xnor U2652 (N_2652,N_1738,N_1300);
and U2653 (N_2653,N_1919,N_1969);
xnor U2654 (N_2654,N_1419,N_1885);
or U2655 (N_2655,N_1307,N_1944);
nand U2656 (N_2656,N_1394,N_1831);
or U2657 (N_2657,N_1140,N_1369);
and U2658 (N_2658,N_1344,N_1297);
xor U2659 (N_2659,N_1650,N_1741);
nand U2660 (N_2660,N_1528,N_1798);
or U2661 (N_2661,N_1617,N_1975);
nor U2662 (N_2662,N_1981,N_1925);
or U2663 (N_2663,N_1437,N_1740);
nor U2664 (N_2664,N_1768,N_1313);
nand U2665 (N_2665,N_1380,N_1769);
or U2666 (N_2666,N_1641,N_1708);
nand U2667 (N_2667,N_1506,N_1298);
or U2668 (N_2668,N_1275,N_1077);
nand U2669 (N_2669,N_1948,N_1222);
xor U2670 (N_2670,N_1586,N_1848);
and U2671 (N_2671,N_1232,N_1540);
xnor U2672 (N_2672,N_1052,N_1860);
or U2673 (N_2673,N_1566,N_1588);
nor U2674 (N_2674,N_1508,N_1017);
nand U2675 (N_2675,N_1363,N_1638);
or U2676 (N_2676,N_1633,N_1463);
or U2677 (N_2677,N_1579,N_1497);
nor U2678 (N_2678,N_1443,N_1588);
nor U2679 (N_2679,N_1174,N_1618);
and U2680 (N_2680,N_1319,N_1049);
nand U2681 (N_2681,N_1113,N_1923);
xnor U2682 (N_2682,N_1438,N_1269);
nor U2683 (N_2683,N_1929,N_1656);
nand U2684 (N_2684,N_1394,N_1738);
xor U2685 (N_2685,N_1272,N_1670);
nor U2686 (N_2686,N_1572,N_1775);
or U2687 (N_2687,N_1234,N_1883);
or U2688 (N_2688,N_1898,N_1273);
xnor U2689 (N_2689,N_1290,N_1131);
and U2690 (N_2690,N_1833,N_1092);
nor U2691 (N_2691,N_1276,N_1851);
nand U2692 (N_2692,N_1830,N_1595);
and U2693 (N_2693,N_1443,N_1999);
or U2694 (N_2694,N_1629,N_1696);
and U2695 (N_2695,N_1833,N_1125);
xor U2696 (N_2696,N_1125,N_1638);
or U2697 (N_2697,N_1133,N_1634);
or U2698 (N_2698,N_1389,N_1848);
or U2699 (N_2699,N_1616,N_1768);
xnor U2700 (N_2700,N_1853,N_1689);
nand U2701 (N_2701,N_1635,N_1088);
nor U2702 (N_2702,N_1143,N_1556);
nand U2703 (N_2703,N_1018,N_1970);
or U2704 (N_2704,N_1223,N_1600);
xnor U2705 (N_2705,N_1127,N_1872);
and U2706 (N_2706,N_1273,N_1394);
and U2707 (N_2707,N_1879,N_1173);
nor U2708 (N_2708,N_1317,N_1881);
nor U2709 (N_2709,N_1270,N_1644);
xnor U2710 (N_2710,N_1822,N_1333);
or U2711 (N_2711,N_1702,N_1457);
xnor U2712 (N_2712,N_1574,N_1197);
nand U2713 (N_2713,N_1612,N_1114);
xor U2714 (N_2714,N_1713,N_1441);
or U2715 (N_2715,N_1295,N_1140);
xor U2716 (N_2716,N_1563,N_1590);
nor U2717 (N_2717,N_1250,N_1097);
nor U2718 (N_2718,N_1000,N_1514);
xor U2719 (N_2719,N_1915,N_1367);
xnor U2720 (N_2720,N_1147,N_1287);
nand U2721 (N_2721,N_1775,N_1179);
and U2722 (N_2722,N_1363,N_1736);
nand U2723 (N_2723,N_1897,N_1252);
and U2724 (N_2724,N_1440,N_1138);
and U2725 (N_2725,N_1499,N_1201);
nor U2726 (N_2726,N_1756,N_1619);
nor U2727 (N_2727,N_1435,N_1803);
nor U2728 (N_2728,N_1763,N_1316);
nor U2729 (N_2729,N_1199,N_1976);
and U2730 (N_2730,N_1756,N_1833);
nand U2731 (N_2731,N_1941,N_1416);
or U2732 (N_2732,N_1526,N_1136);
and U2733 (N_2733,N_1079,N_1088);
nand U2734 (N_2734,N_1778,N_1136);
nor U2735 (N_2735,N_1914,N_1963);
nor U2736 (N_2736,N_1344,N_1340);
nand U2737 (N_2737,N_1291,N_1401);
xor U2738 (N_2738,N_1061,N_1985);
nor U2739 (N_2739,N_1268,N_1069);
and U2740 (N_2740,N_1888,N_1226);
nor U2741 (N_2741,N_1126,N_1916);
or U2742 (N_2742,N_1803,N_1706);
xnor U2743 (N_2743,N_1686,N_1777);
nor U2744 (N_2744,N_1217,N_1308);
or U2745 (N_2745,N_1396,N_1036);
or U2746 (N_2746,N_1609,N_1707);
nor U2747 (N_2747,N_1755,N_1086);
nand U2748 (N_2748,N_1649,N_1696);
and U2749 (N_2749,N_1325,N_1121);
xnor U2750 (N_2750,N_1289,N_1599);
xor U2751 (N_2751,N_1078,N_1374);
nor U2752 (N_2752,N_1596,N_1843);
and U2753 (N_2753,N_1876,N_1732);
or U2754 (N_2754,N_1655,N_1955);
nor U2755 (N_2755,N_1604,N_1087);
and U2756 (N_2756,N_1942,N_1216);
and U2757 (N_2757,N_1279,N_1346);
or U2758 (N_2758,N_1300,N_1905);
or U2759 (N_2759,N_1509,N_1726);
or U2760 (N_2760,N_1504,N_1932);
xnor U2761 (N_2761,N_1661,N_1968);
nand U2762 (N_2762,N_1165,N_1481);
or U2763 (N_2763,N_1665,N_1290);
xnor U2764 (N_2764,N_1122,N_1496);
nor U2765 (N_2765,N_1810,N_1774);
or U2766 (N_2766,N_1380,N_1221);
or U2767 (N_2767,N_1013,N_1177);
nor U2768 (N_2768,N_1795,N_1714);
nand U2769 (N_2769,N_1551,N_1692);
or U2770 (N_2770,N_1294,N_1602);
or U2771 (N_2771,N_1736,N_1679);
xor U2772 (N_2772,N_1686,N_1066);
and U2773 (N_2773,N_1379,N_1146);
or U2774 (N_2774,N_1467,N_1062);
or U2775 (N_2775,N_1496,N_1029);
or U2776 (N_2776,N_1815,N_1387);
and U2777 (N_2777,N_1795,N_1357);
nor U2778 (N_2778,N_1727,N_1349);
nor U2779 (N_2779,N_1732,N_1859);
nand U2780 (N_2780,N_1217,N_1817);
nand U2781 (N_2781,N_1843,N_1733);
or U2782 (N_2782,N_1948,N_1444);
nor U2783 (N_2783,N_1637,N_1113);
xnor U2784 (N_2784,N_1637,N_1018);
nand U2785 (N_2785,N_1233,N_1418);
and U2786 (N_2786,N_1600,N_1392);
nor U2787 (N_2787,N_1449,N_1698);
nand U2788 (N_2788,N_1067,N_1848);
nor U2789 (N_2789,N_1694,N_1636);
nor U2790 (N_2790,N_1802,N_1084);
xor U2791 (N_2791,N_1664,N_1677);
xnor U2792 (N_2792,N_1479,N_1349);
or U2793 (N_2793,N_1729,N_1066);
xor U2794 (N_2794,N_1538,N_1479);
or U2795 (N_2795,N_1814,N_1479);
nand U2796 (N_2796,N_1648,N_1920);
xnor U2797 (N_2797,N_1019,N_1378);
nor U2798 (N_2798,N_1314,N_1417);
nor U2799 (N_2799,N_1988,N_1252);
xor U2800 (N_2800,N_1129,N_1844);
nand U2801 (N_2801,N_1146,N_1967);
nand U2802 (N_2802,N_1118,N_1032);
and U2803 (N_2803,N_1567,N_1147);
and U2804 (N_2804,N_1226,N_1633);
or U2805 (N_2805,N_1846,N_1228);
xor U2806 (N_2806,N_1851,N_1828);
xor U2807 (N_2807,N_1557,N_1871);
nand U2808 (N_2808,N_1166,N_1542);
xnor U2809 (N_2809,N_1566,N_1093);
nor U2810 (N_2810,N_1507,N_1149);
or U2811 (N_2811,N_1031,N_1347);
nor U2812 (N_2812,N_1460,N_1945);
or U2813 (N_2813,N_1298,N_1712);
xnor U2814 (N_2814,N_1962,N_1989);
xor U2815 (N_2815,N_1643,N_1719);
nor U2816 (N_2816,N_1335,N_1200);
and U2817 (N_2817,N_1487,N_1931);
and U2818 (N_2818,N_1613,N_1367);
xor U2819 (N_2819,N_1213,N_1146);
or U2820 (N_2820,N_1197,N_1721);
xnor U2821 (N_2821,N_1015,N_1365);
nand U2822 (N_2822,N_1396,N_1818);
nor U2823 (N_2823,N_1144,N_1541);
nor U2824 (N_2824,N_1804,N_1604);
xor U2825 (N_2825,N_1834,N_1327);
or U2826 (N_2826,N_1517,N_1824);
xnor U2827 (N_2827,N_1381,N_1311);
nand U2828 (N_2828,N_1804,N_1968);
xor U2829 (N_2829,N_1784,N_1703);
nor U2830 (N_2830,N_1179,N_1725);
and U2831 (N_2831,N_1781,N_1804);
and U2832 (N_2832,N_1951,N_1905);
nand U2833 (N_2833,N_1453,N_1066);
and U2834 (N_2834,N_1589,N_1139);
nand U2835 (N_2835,N_1767,N_1094);
xnor U2836 (N_2836,N_1490,N_1177);
nand U2837 (N_2837,N_1810,N_1691);
or U2838 (N_2838,N_1531,N_1559);
or U2839 (N_2839,N_1522,N_1940);
or U2840 (N_2840,N_1016,N_1662);
nor U2841 (N_2841,N_1652,N_1000);
and U2842 (N_2842,N_1430,N_1791);
xor U2843 (N_2843,N_1145,N_1004);
xor U2844 (N_2844,N_1233,N_1391);
nor U2845 (N_2845,N_1176,N_1874);
and U2846 (N_2846,N_1590,N_1959);
xnor U2847 (N_2847,N_1758,N_1347);
xnor U2848 (N_2848,N_1947,N_1491);
or U2849 (N_2849,N_1173,N_1991);
xor U2850 (N_2850,N_1805,N_1718);
nand U2851 (N_2851,N_1025,N_1399);
nand U2852 (N_2852,N_1069,N_1818);
or U2853 (N_2853,N_1396,N_1811);
and U2854 (N_2854,N_1015,N_1800);
or U2855 (N_2855,N_1771,N_1227);
and U2856 (N_2856,N_1175,N_1694);
xor U2857 (N_2857,N_1053,N_1976);
xnor U2858 (N_2858,N_1417,N_1102);
xnor U2859 (N_2859,N_1536,N_1529);
nor U2860 (N_2860,N_1163,N_1692);
or U2861 (N_2861,N_1981,N_1397);
nor U2862 (N_2862,N_1203,N_1758);
and U2863 (N_2863,N_1445,N_1735);
nand U2864 (N_2864,N_1799,N_1013);
or U2865 (N_2865,N_1840,N_1677);
and U2866 (N_2866,N_1976,N_1022);
nand U2867 (N_2867,N_1296,N_1456);
xor U2868 (N_2868,N_1323,N_1765);
or U2869 (N_2869,N_1907,N_1890);
and U2870 (N_2870,N_1754,N_1809);
and U2871 (N_2871,N_1947,N_1143);
and U2872 (N_2872,N_1261,N_1722);
and U2873 (N_2873,N_1654,N_1657);
nand U2874 (N_2874,N_1914,N_1411);
xnor U2875 (N_2875,N_1700,N_1219);
and U2876 (N_2876,N_1360,N_1483);
xor U2877 (N_2877,N_1771,N_1038);
nor U2878 (N_2878,N_1368,N_1809);
nand U2879 (N_2879,N_1652,N_1875);
nand U2880 (N_2880,N_1450,N_1387);
nor U2881 (N_2881,N_1994,N_1845);
xor U2882 (N_2882,N_1250,N_1648);
xor U2883 (N_2883,N_1596,N_1405);
or U2884 (N_2884,N_1618,N_1022);
nor U2885 (N_2885,N_1708,N_1258);
xor U2886 (N_2886,N_1235,N_1978);
nor U2887 (N_2887,N_1112,N_1655);
nor U2888 (N_2888,N_1287,N_1740);
nand U2889 (N_2889,N_1063,N_1543);
nor U2890 (N_2890,N_1597,N_1705);
xor U2891 (N_2891,N_1086,N_1043);
nand U2892 (N_2892,N_1671,N_1940);
nand U2893 (N_2893,N_1895,N_1898);
xnor U2894 (N_2894,N_1792,N_1553);
and U2895 (N_2895,N_1839,N_1553);
nand U2896 (N_2896,N_1555,N_1825);
or U2897 (N_2897,N_1738,N_1742);
xnor U2898 (N_2898,N_1460,N_1575);
nor U2899 (N_2899,N_1814,N_1977);
or U2900 (N_2900,N_1486,N_1603);
and U2901 (N_2901,N_1904,N_1884);
and U2902 (N_2902,N_1574,N_1046);
or U2903 (N_2903,N_1769,N_1790);
and U2904 (N_2904,N_1165,N_1913);
xnor U2905 (N_2905,N_1390,N_1894);
and U2906 (N_2906,N_1147,N_1211);
nand U2907 (N_2907,N_1733,N_1824);
nor U2908 (N_2908,N_1410,N_1198);
and U2909 (N_2909,N_1774,N_1687);
or U2910 (N_2910,N_1282,N_1644);
or U2911 (N_2911,N_1867,N_1000);
xnor U2912 (N_2912,N_1028,N_1064);
nand U2913 (N_2913,N_1838,N_1422);
or U2914 (N_2914,N_1744,N_1756);
nand U2915 (N_2915,N_1468,N_1283);
or U2916 (N_2916,N_1371,N_1206);
nand U2917 (N_2917,N_1247,N_1675);
nand U2918 (N_2918,N_1314,N_1178);
nor U2919 (N_2919,N_1009,N_1596);
or U2920 (N_2920,N_1571,N_1534);
or U2921 (N_2921,N_1095,N_1366);
and U2922 (N_2922,N_1947,N_1418);
nor U2923 (N_2923,N_1752,N_1598);
nand U2924 (N_2924,N_1318,N_1000);
nor U2925 (N_2925,N_1665,N_1645);
nand U2926 (N_2926,N_1423,N_1940);
xor U2927 (N_2927,N_1137,N_1287);
nor U2928 (N_2928,N_1339,N_1818);
nand U2929 (N_2929,N_1159,N_1938);
nand U2930 (N_2930,N_1656,N_1581);
xnor U2931 (N_2931,N_1254,N_1890);
xor U2932 (N_2932,N_1532,N_1276);
and U2933 (N_2933,N_1375,N_1108);
and U2934 (N_2934,N_1099,N_1519);
and U2935 (N_2935,N_1646,N_1099);
nand U2936 (N_2936,N_1116,N_1395);
or U2937 (N_2937,N_1261,N_1568);
and U2938 (N_2938,N_1859,N_1822);
or U2939 (N_2939,N_1964,N_1330);
nor U2940 (N_2940,N_1388,N_1592);
nor U2941 (N_2941,N_1354,N_1299);
nand U2942 (N_2942,N_1325,N_1198);
and U2943 (N_2943,N_1995,N_1052);
xnor U2944 (N_2944,N_1439,N_1433);
xnor U2945 (N_2945,N_1707,N_1914);
nor U2946 (N_2946,N_1266,N_1631);
xor U2947 (N_2947,N_1848,N_1756);
nand U2948 (N_2948,N_1973,N_1916);
or U2949 (N_2949,N_1798,N_1276);
and U2950 (N_2950,N_1204,N_1881);
and U2951 (N_2951,N_1186,N_1264);
or U2952 (N_2952,N_1495,N_1854);
or U2953 (N_2953,N_1889,N_1277);
and U2954 (N_2954,N_1469,N_1941);
and U2955 (N_2955,N_1534,N_1145);
and U2956 (N_2956,N_1826,N_1320);
and U2957 (N_2957,N_1916,N_1698);
nand U2958 (N_2958,N_1258,N_1026);
nor U2959 (N_2959,N_1143,N_1830);
nor U2960 (N_2960,N_1630,N_1921);
nor U2961 (N_2961,N_1483,N_1560);
and U2962 (N_2962,N_1138,N_1926);
xor U2963 (N_2963,N_1368,N_1441);
or U2964 (N_2964,N_1583,N_1527);
or U2965 (N_2965,N_1808,N_1123);
nor U2966 (N_2966,N_1480,N_1775);
or U2967 (N_2967,N_1560,N_1423);
nor U2968 (N_2968,N_1858,N_1897);
nand U2969 (N_2969,N_1123,N_1714);
nor U2970 (N_2970,N_1371,N_1579);
and U2971 (N_2971,N_1062,N_1714);
and U2972 (N_2972,N_1136,N_1509);
xnor U2973 (N_2973,N_1077,N_1442);
nor U2974 (N_2974,N_1715,N_1135);
or U2975 (N_2975,N_1548,N_1955);
and U2976 (N_2976,N_1093,N_1399);
nand U2977 (N_2977,N_1419,N_1308);
or U2978 (N_2978,N_1097,N_1448);
nand U2979 (N_2979,N_1786,N_1246);
or U2980 (N_2980,N_1425,N_1120);
nand U2981 (N_2981,N_1588,N_1087);
and U2982 (N_2982,N_1475,N_1061);
or U2983 (N_2983,N_1411,N_1966);
nand U2984 (N_2984,N_1797,N_1052);
and U2985 (N_2985,N_1757,N_1085);
and U2986 (N_2986,N_1823,N_1285);
and U2987 (N_2987,N_1011,N_1457);
and U2988 (N_2988,N_1862,N_1569);
xnor U2989 (N_2989,N_1512,N_1883);
xor U2990 (N_2990,N_1958,N_1960);
xor U2991 (N_2991,N_1484,N_1294);
and U2992 (N_2992,N_1161,N_1871);
nor U2993 (N_2993,N_1234,N_1002);
nor U2994 (N_2994,N_1372,N_1699);
nand U2995 (N_2995,N_1988,N_1043);
nor U2996 (N_2996,N_1777,N_1107);
xor U2997 (N_2997,N_1054,N_1301);
xnor U2998 (N_2998,N_1550,N_1664);
and U2999 (N_2999,N_1304,N_1011);
xor UO_0 (O_0,N_2808,N_2000);
and UO_1 (O_1,N_2462,N_2694);
nand UO_2 (O_2,N_2554,N_2823);
xnor UO_3 (O_3,N_2116,N_2967);
and UO_4 (O_4,N_2741,N_2849);
and UO_5 (O_5,N_2842,N_2244);
or UO_6 (O_6,N_2128,N_2556);
and UO_7 (O_7,N_2638,N_2494);
xnor UO_8 (O_8,N_2384,N_2342);
and UO_9 (O_9,N_2130,N_2322);
nor UO_10 (O_10,N_2396,N_2492);
nor UO_11 (O_11,N_2773,N_2618);
nand UO_12 (O_12,N_2931,N_2429);
nor UO_13 (O_13,N_2519,N_2856);
nor UO_14 (O_14,N_2250,N_2937);
xor UO_15 (O_15,N_2650,N_2604);
nand UO_16 (O_16,N_2547,N_2348);
or UO_17 (O_17,N_2076,N_2945);
xor UO_18 (O_18,N_2811,N_2804);
nand UO_19 (O_19,N_2932,N_2088);
xnor UO_20 (O_20,N_2413,N_2328);
nor UO_21 (O_21,N_2791,N_2714);
nor UO_22 (O_22,N_2266,N_2057);
and UO_23 (O_23,N_2353,N_2758);
nand UO_24 (O_24,N_2837,N_2537);
nand UO_25 (O_25,N_2767,N_2192);
or UO_26 (O_26,N_2460,N_2739);
or UO_27 (O_27,N_2135,N_2027);
and UO_28 (O_28,N_2038,N_2916);
or UO_29 (O_29,N_2672,N_2805);
or UO_30 (O_30,N_2450,N_2776);
and UO_31 (O_31,N_2892,N_2716);
nand UO_32 (O_32,N_2015,N_2345);
nand UO_33 (O_33,N_2707,N_2898);
nand UO_34 (O_34,N_2184,N_2279);
nor UO_35 (O_35,N_2616,N_2973);
nand UO_36 (O_36,N_2596,N_2398);
nand UO_37 (O_37,N_2676,N_2526);
nor UO_38 (O_38,N_2605,N_2889);
nand UO_39 (O_39,N_2885,N_2026);
or UO_40 (O_40,N_2745,N_2018);
nand UO_41 (O_41,N_2477,N_2882);
or UO_42 (O_42,N_2771,N_2507);
xnor UO_43 (O_43,N_2444,N_2834);
nor UO_44 (O_44,N_2665,N_2032);
nand UO_45 (O_45,N_2341,N_2478);
nor UO_46 (O_46,N_2534,N_2533);
xnor UO_47 (O_47,N_2330,N_2990);
nor UO_48 (O_48,N_2729,N_2818);
xor UO_49 (O_49,N_2235,N_2370);
nand UO_50 (O_50,N_2117,N_2115);
xor UO_51 (O_51,N_2245,N_2439);
xnor UO_52 (O_52,N_2840,N_2911);
nand UO_53 (O_53,N_2590,N_2501);
nand UO_54 (O_54,N_2784,N_2624);
xnor UO_55 (O_55,N_2918,N_2023);
or UO_56 (O_56,N_2021,N_2402);
nand UO_57 (O_57,N_2230,N_2799);
and UO_58 (O_58,N_2742,N_2233);
or UO_59 (O_59,N_2813,N_2265);
and UO_60 (O_60,N_2552,N_2003);
or UO_61 (O_61,N_2428,N_2022);
or UO_62 (O_62,N_2843,N_2409);
and UO_63 (O_63,N_2748,N_2008);
nor UO_64 (O_64,N_2972,N_2603);
nand UO_65 (O_65,N_2613,N_2956);
or UO_66 (O_66,N_2597,N_2194);
or UO_67 (O_67,N_2179,N_2427);
nand UO_68 (O_68,N_2103,N_2900);
nand UO_69 (O_69,N_2254,N_2452);
nor UO_70 (O_70,N_2706,N_2053);
nor UO_71 (O_71,N_2393,N_2642);
and UO_72 (O_72,N_2877,N_2288);
and UO_73 (O_73,N_2327,N_2756);
or UO_74 (O_74,N_2576,N_2903);
nand UO_75 (O_75,N_2123,N_2583);
xnor UO_76 (O_76,N_2432,N_2168);
and UO_77 (O_77,N_2440,N_2311);
nand UO_78 (O_78,N_2326,N_2757);
and UO_79 (O_79,N_2197,N_2518);
or UO_80 (O_80,N_2403,N_2368);
nand UO_81 (O_81,N_2899,N_2559);
or UO_82 (O_82,N_2708,N_2294);
nor UO_83 (O_83,N_2183,N_2521);
nor UO_84 (O_84,N_2270,N_2810);
xnor UO_85 (O_85,N_2530,N_2435);
xor UO_86 (O_86,N_2122,N_2307);
nand UO_87 (O_87,N_2005,N_2713);
nor UO_88 (O_88,N_2912,N_2788);
nand UO_89 (O_89,N_2553,N_2321);
nand UO_90 (O_90,N_2966,N_2221);
or UO_91 (O_91,N_2928,N_2424);
nand UO_92 (O_92,N_2259,N_2723);
nand UO_93 (O_93,N_2062,N_2140);
and UO_94 (O_94,N_2137,N_2175);
nor UO_95 (O_95,N_2880,N_2725);
or UO_96 (O_96,N_2306,N_2142);
nand UO_97 (O_97,N_2861,N_2416);
xnor UO_98 (O_98,N_2679,N_2592);
xor UO_99 (O_99,N_2798,N_2701);
or UO_100 (O_100,N_2352,N_2802);
or UO_101 (O_101,N_2496,N_2119);
or UO_102 (O_102,N_2796,N_2782);
nor UO_103 (O_103,N_2357,N_2981);
xnor UO_104 (O_104,N_2852,N_2129);
or UO_105 (O_105,N_2162,N_2487);
nor UO_106 (O_106,N_2940,N_2565);
nor UO_107 (O_107,N_2464,N_2243);
or UO_108 (O_108,N_2738,N_2278);
nor UO_109 (O_109,N_2905,N_2256);
nand UO_110 (O_110,N_2586,N_2475);
nor UO_111 (O_111,N_2923,N_2505);
xor UO_112 (O_112,N_2835,N_2978);
nand UO_113 (O_113,N_2012,N_2252);
or UO_114 (O_114,N_2848,N_2921);
nor UO_115 (O_115,N_2410,N_2408);
xor UO_116 (O_116,N_2696,N_2317);
nand UO_117 (O_117,N_2608,N_2864);
nor UO_118 (O_118,N_2079,N_2721);
or UO_119 (O_119,N_2793,N_2355);
and UO_120 (O_120,N_2606,N_2759);
or UO_121 (O_121,N_2845,N_2711);
nand UO_122 (O_122,N_2936,N_2871);
and UO_123 (O_123,N_2607,N_2527);
or UO_124 (O_124,N_2684,N_2500);
or UO_125 (O_125,N_2346,N_2289);
xor UO_126 (O_126,N_2447,N_2002);
and UO_127 (O_127,N_2207,N_2068);
nor UO_128 (O_128,N_2036,N_2052);
nand UO_129 (O_129,N_2906,N_2881);
or UO_130 (O_130,N_2013,N_2948);
nand UO_131 (O_131,N_2241,N_2786);
and UO_132 (O_132,N_2663,N_2456);
nor UO_133 (O_133,N_2177,N_2577);
xor UO_134 (O_134,N_2532,N_2872);
or UO_135 (O_135,N_2271,N_2743);
and UO_136 (O_136,N_2640,N_2084);
nor UO_137 (O_137,N_2783,N_2320);
nand UO_138 (O_138,N_2512,N_2910);
or UO_139 (O_139,N_2083,N_2657);
nand UO_140 (O_140,N_2860,N_2132);
or UO_141 (O_141,N_2373,N_2296);
and UO_142 (O_142,N_2314,N_2358);
xor UO_143 (O_143,N_2417,N_2516);
nand UO_144 (O_144,N_2267,N_2111);
and UO_145 (O_145,N_2350,N_2754);
nand UO_146 (O_146,N_2426,N_2147);
nor UO_147 (O_147,N_2213,N_2645);
and UO_148 (O_148,N_2509,N_2564);
xnor UO_149 (O_149,N_2594,N_2089);
and UO_150 (O_150,N_2612,N_2772);
xor UO_151 (O_151,N_2400,N_2205);
or UO_152 (O_152,N_2273,N_2688);
nor UO_153 (O_153,N_2702,N_2572);
nor UO_154 (O_154,N_2765,N_2983);
nand UO_155 (O_155,N_2859,N_2337);
and UO_156 (O_156,N_2755,N_2405);
nor UO_157 (O_157,N_2324,N_2732);
xnor UO_158 (O_158,N_2946,N_2951);
xnor UO_159 (O_159,N_2499,N_2463);
nor UO_160 (O_160,N_2482,N_2020);
nand UO_161 (O_161,N_2007,N_2483);
nor UO_162 (O_162,N_2920,N_2854);
nor UO_163 (O_163,N_2838,N_2704);
or UO_164 (O_164,N_2924,N_2979);
nand UO_165 (O_165,N_2902,N_2588);
nand UO_166 (O_166,N_2391,N_2822);
xnor UO_167 (O_167,N_2568,N_2941);
nor UO_168 (O_168,N_2280,N_2865);
and UO_169 (O_169,N_2367,N_2195);
nand UO_170 (O_170,N_2958,N_2121);
nor UO_171 (O_171,N_2102,N_2883);
nand UO_172 (O_172,N_2141,N_2257);
and UO_173 (O_173,N_2927,N_2231);
or UO_174 (O_174,N_2727,N_2263);
xnor UO_175 (O_175,N_2495,N_2746);
nand UO_176 (O_176,N_2922,N_2453);
xor UO_177 (O_177,N_2987,N_2998);
nor UO_178 (O_178,N_2363,N_2082);
xnor UO_179 (O_179,N_2040,N_2909);
nor UO_180 (O_180,N_2693,N_2430);
nor UO_181 (O_181,N_2770,N_2420);
or UO_182 (O_182,N_2493,N_2692);
or UO_183 (O_183,N_2174,N_2481);
and UO_184 (O_184,N_2646,N_2066);
nor UO_185 (O_185,N_2366,N_2274);
xnor UO_186 (O_186,N_2752,N_2143);
or UO_187 (O_187,N_2044,N_2181);
nand UO_188 (O_188,N_2389,N_2037);
xnor UO_189 (O_189,N_2504,N_2635);
or UO_190 (O_190,N_2726,N_2886);
xor UO_191 (O_191,N_2950,N_2761);
and UO_192 (O_192,N_2208,N_2292);
and UO_193 (O_193,N_2360,N_2960);
nand UO_194 (O_194,N_2826,N_2302);
nor UO_195 (O_195,N_2893,N_2421);
xor UO_196 (O_196,N_2285,N_2001);
and UO_197 (O_197,N_2238,N_2092);
or UO_198 (O_198,N_2098,N_2108);
xnor UO_199 (O_199,N_2331,N_2293);
and UO_200 (O_200,N_2620,N_2217);
nor UO_201 (O_201,N_2789,N_2401);
nand UO_202 (O_202,N_2332,N_2457);
and UO_203 (O_203,N_2844,N_2569);
nand UO_204 (O_204,N_2218,N_2160);
or UO_205 (O_205,N_2514,N_2622);
nand UO_206 (O_206,N_2641,N_2153);
or UO_207 (O_207,N_2340,N_2541);
and UO_208 (O_208,N_2815,N_2077);
xnor UO_209 (O_209,N_2287,N_2709);
or UO_210 (O_210,N_2361,N_2466);
xor UO_211 (O_211,N_2386,N_2609);
nor UO_212 (O_212,N_2744,N_2976);
nor UO_213 (O_213,N_2157,N_2778);
and UO_214 (O_214,N_2919,N_2781);
and UO_215 (O_215,N_2907,N_2310);
nand UO_216 (O_216,N_2281,N_2339);
and UO_217 (O_217,N_2619,N_2884);
nand UO_218 (O_218,N_2644,N_2751);
nor UO_219 (O_219,N_2166,N_2974);
nand UO_220 (O_220,N_2890,N_2485);
xnor UO_221 (O_221,N_2390,N_2938);
and UO_222 (O_222,N_2461,N_2199);
nor UO_223 (O_223,N_2762,N_2561);
nand UO_224 (O_224,N_2853,N_2740);
or UO_225 (O_225,N_2614,N_2993);
nor UO_226 (O_226,N_2343,N_2298);
and UO_227 (O_227,N_2030,N_2867);
or UO_228 (O_228,N_2858,N_2061);
nand UO_229 (O_229,N_2200,N_2049);
nor UO_230 (O_230,N_2387,N_2193);
or UO_231 (O_231,N_2081,N_2961);
or UO_232 (O_232,N_2125,N_2204);
xor UO_233 (O_233,N_2722,N_2520);
nor UO_234 (O_234,N_2009,N_2631);
nor UO_235 (O_235,N_2422,N_2769);
and UO_236 (O_236,N_2570,N_2836);
and UO_237 (O_237,N_2949,N_2582);
or UO_238 (O_238,N_2643,N_2550);
nand UO_239 (O_239,N_2503,N_2627);
and UO_240 (O_240,N_2730,N_2104);
nor UO_241 (O_241,N_2099,N_2043);
and UO_242 (O_242,N_2297,N_2237);
nand UO_243 (O_243,N_2699,N_2623);
and UO_244 (O_244,N_2374,N_2508);
nand UO_245 (O_245,N_2144,N_2551);
and UO_246 (O_246,N_2154,N_2455);
nor UO_247 (O_247,N_2930,N_2107);
xnor UO_248 (O_248,N_2172,N_2803);
xor UO_249 (O_249,N_2965,N_2290);
nand UO_250 (O_250,N_2397,N_2807);
nor UO_251 (O_251,N_2220,N_2656);
nand UO_252 (O_252,N_2134,N_2933);
xor UO_253 (O_253,N_2991,N_2975);
or UO_254 (O_254,N_2375,N_2468);
nand UO_255 (O_255,N_2225,N_2563);
nand UO_256 (O_256,N_2097,N_2513);
and UO_257 (O_257,N_2528,N_2055);
and UO_258 (O_258,N_2029,N_2469);
xor UO_259 (O_259,N_2634,N_2599);
nand UO_260 (O_260,N_2830,N_2666);
and UO_261 (O_261,N_2356,N_2118);
xnor UO_262 (O_262,N_2024,N_2473);
xor UO_263 (O_263,N_2379,N_2774);
and UO_264 (O_264,N_2105,N_2540);
nor UO_265 (O_265,N_2251,N_2498);
or UO_266 (O_266,N_2600,N_2080);
xnor UO_267 (O_267,N_2490,N_2150);
nor UO_268 (O_268,N_2749,N_2735);
nand UO_269 (O_269,N_2598,N_2051);
and UO_270 (O_270,N_2010,N_2847);
nand UO_271 (O_271,N_2070,N_2628);
nand UO_272 (O_272,N_2678,N_2187);
nor UO_273 (O_273,N_2863,N_2698);
nand UO_274 (O_274,N_2249,N_2915);
nor UO_275 (O_275,N_2690,N_2846);
nor UO_276 (O_276,N_2939,N_2303);
nand UO_277 (O_277,N_2214,N_2717);
nand UO_278 (O_278,N_2006,N_2511);
or UO_279 (O_279,N_2575,N_2347);
nand UO_280 (O_280,N_2065,N_2591);
nand UO_281 (O_281,N_2824,N_2056);
and UO_282 (O_282,N_2489,N_2675);
xor UO_283 (O_283,N_2574,N_2146);
nor UO_284 (O_284,N_2674,N_2985);
nand UO_285 (O_285,N_2202,N_2433);
nand UO_286 (O_286,N_2470,N_2325);
nor UO_287 (O_287,N_2747,N_2913);
or UO_288 (O_288,N_2438,N_2067);
or UO_289 (O_289,N_2476,N_2647);
nand UO_290 (O_290,N_2680,N_2219);
xor UO_291 (O_291,N_2904,N_2560);
and UO_292 (O_292,N_2894,N_2106);
nand UO_293 (O_293,N_2887,N_2093);
and UO_294 (O_294,N_2868,N_2284);
nand UO_295 (O_295,N_2159,N_2562);
nor UO_296 (O_296,N_2819,N_2406);
xnor UO_297 (O_297,N_2630,N_2180);
nor UO_298 (O_298,N_2419,N_2649);
xnor UO_299 (O_299,N_2443,N_2779);
xnor UO_300 (O_300,N_2829,N_2720);
nand UO_301 (O_301,N_2203,N_2999);
nand UO_302 (O_302,N_2654,N_2571);
or UO_303 (O_303,N_2545,N_2689);
nand UO_304 (O_304,N_2934,N_2212);
and UO_305 (O_305,N_2874,N_2959);
or UO_306 (O_306,N_2411,N_2377);
or UO_307 (O_307,N_2888,N_2178);
nor UO_308 (O_308,N_2072,N_2228);
or UO_309 (O_309,N_2334,N_2418);
xor UO_310 (O_310,N_2529,N_2486);
or UO_311 (O_311,N_2659,N_2362);
or UO_312 (O_312,N_2794,N_2277);
and UO_313 (O_313,N_2149,N_2268);
nand UO_314 (O_314,N_2611,N_2970);
nand UO_315 (O_315,N_2047,N_2425);
nand UO_316 (O_316,N_2549,N_2766);
xor UO_317 (O_317,N_2392,N_2035);
or UO_318 (O_318,N_2064,N_2996);
or UO_319 (O_319,N_2691,N_2126);
nor UO_320 (O_320,N_2091,N_2349);
nand UO_321 (O_321,N_2138,N_2094);
xnor UO_322 (O_322,N_2929,N_2479);
nand UO_323 (O_323,N_2448,N_2151);
xor UO_324 (O_324,N_2113,N_2777);
and UO_325 (O_325,N_2226,N_2019);
and UO_326 (O_326,N_2982,N_2372);
or UO_327 (O_327,N_2211,N_2261);
and UO_328 (O_328,N_2850,N_2046);
nor UO_329 (O_329,N_2995,N_2045);
or UO_330 (O_330,N_2831,N_2736);
nor UO_331 (O_331,N_2544,N_2371);
xor UO_332 (O_332,N_2812,N_2615);
or UO_333 (O_333,N_2814,N_2626);
nor UO_334 (O_334,N_2917,N_2100);
xor UO_335 (O_335,N_2558,N_2828);
xor UO_336 (O_336,N_2316,N_2120);
xnor UO_337 (O_337,N_2733,N_2087);
nor UO_338 (O_338,N_2388,N_2242);
or UO_339 (O_339,N_2291,N_2039);
nor UO_340 (O_340,N_2060,N_2189);
xnor UO_341 (O_341,N_2472,N_2165);
xor UO_342 (O_342,N_2381,N_2318);
or UO_343 (O_343,N_2336,N_2145);
or UO_344 (O_344,N_2167,N_2797);
nor UO_345 (O_345,N_2954,N_2801);
or UO_346 (O_346,N_2652,N_2697);
nor UO_347 (O_347,N_2997,N_2750);
nor UO_348 (O_348,N_2283,N_2637);
xnor UO_349 (O_349,N_2685,N_2441);
and UO_350 (O_350,N_2412,N_2073);
nor UO_351 (O_351,N_2943,N_2101);
nor UO_352 (O_352,N_2651,N_2870);
xnor UO_353 (O_353,N_2308,N_2668);
and UO_354 (O_354,N_2262,N_2131);
nand UO_355 (O_355,N_2971,N_2191);
nand UO_356 (O_356,N_2633,N_2925);
nand UO_357 (O_357,N_2664,N_2827);
nor UO_358 (O_358,N_2785,N_2133);
and UO_359 (O_359,N_2787,N_2617);
and UO_360 (O_360,N_2977,N_2525);
xor UO_361 (O_361,N_2017,N_2209);
nand UO_362 (O_362,N_2683,N_2869);
or UO_363 (O_363,N_2295,N_2078);
or UO_364 (O_364,N_2096,N_2809);
xor UO_365 (O_365,N_2992,N_2465);
nand UO_366 (O_366,N_2724,N_2260);
or UO_367 (O_367,N_2338,N_2437);
and UO_368 (O_368,N_2703,N_2248);
xor UO_369 (O_369,N_2090,N_2050);
xnor UO_370 (O_370,N_2182,N_2625);
xor UO_371 (O_371,N_2686,N_2344);
and UO_372 (O_372,N_2404,N_2584);
and UO_373 (O_373,N_2124,N_2610);
nand UO_374 (O_374,N_2063,N_2028);
or UO_375 (O_375,N_2232,N_2434);
xor UO_376 (O_376,N_2399,N_2247);
xnor UO_377 (O_377,N_2944,N_2058);
xnor UO_378 (O_378,N_2086,N_2299);
or UO_379 (O_379,N_2670,N_2395);
and UO_380 (O_380,N_2876,N_2719);
nor UO_381 (O_381,N_2156,N_2567);
nand UO_382 (O_382,N_2282,N_2269);
and UO_383 (O_383,N_2313,N_2309);
xor UO_384 (O_384,N_2988,N_2682);
or UO_385 (O_385,N_2947,N_2557);
nor UO_386 (O_386,N_2535,N_2728);
nor UO_387 (O_387,N_2806,N_2258);
nand UO_388 (O_388,N_2671,N_2589);
and UO_389 (O_389,N_2071,N_2775);
nand UO_390 (O_390,N_2382,N_2161);
or UO_391 (O_391,N_2354,N_2994);
nand UO_392 (O_392,N_2768,N_2715);
or UO_393 (O_393,N_2445,N_2196);
nor UO_394 (O_394,N_2169,N_2431);
and UO_395 (O_395,N_2158,N_2595);
nand UO_396 (O_396,N_2112,N_2669);
and UO_397 (O_397,N_2229,N_2908);
nor UO_398 (O_398,N_2579,N_2376);
nand UO_399 (O_399,N_2369,N_2171);
nand UO_400 (O_400,N_2660,N_2968);
or UO_401 (O_401,N_2531,N_2542);
and UO_402 (O_402,N_2127,N_2109);
or UO_403 (O_403,N_2878,N_2335);
xnor UO_404 (O_404,N_2926,N_2255);
nand UO_405 (O_405,N_2378,N_2790);
xor UO_406 (O_406,N_2662,N_2364);
nand UO_407 (O_407,N_2566,N_2655);
nand UO_408 (O_408,N_2446,N_2839);
and UO_409 (O_409,N_2780,N_2069);
nor UO_410 (O_410,N_2234,N_2517);
nand UO_411 (O_411,N_2891,N_2857);
xor UO_412 (O_412,N_2223,N_2901);
nor UO_413 (O_413,N_2710,N_2963);
xor UO_414 (O_414,N_2164,N_2989);
nand UO_415 (O_415,N_2962,N_2048);
or UO_416 (O_416,N_2578,N_2301);
nor UO_417 (O_417,N_2206,N_2155);
nand UO_418 (O_418,N_2190,N_2639);
and UO_419 (O_419,N_2240,N_2188);
and UO_420 (O_420,N_2731,N_2935);
nand UO_421 (O_421,N_2025,N_2955);
nand UO_422 (O_422,N_2895,N_2170);
nand UO_423 (O_423,N_2833,N_2648);
or UO_424 (O_424,N_2873,N_2059);
or UO_425 (O_425,N_2817,N_2186);
nand UO_426 (O_426,N_2276,N_2661);
nor UO_427 (O_427,N_2383,N_2964);
or UO_428 (O_428,N_2969,N_2763);
or UO_429 (O_429,N_2705,N_2862);
xor UO_430 (O_430,N_2380,N_2510);
nand UO_431 (O_431,N_2329,N_2467);
nor UO_432 (O_432,N_2041,N_2074);
or UO_433 (O_433,N_2673,N_2246);
nor UO_434 (O_434,N_2866,N_2451);
and UO_435 (O_435,N_2800,N_2210);
nand UO_436 (O_436,N_2198,N_2152);
and UO_437 (O_437,N_2984,N_2602);
nor UO_438 (O_438,N_2239,N_2095);
nand UO_439 (O_439,N_2524,N_2555);
xnor UO_440 (O_440,N_2832,N_2523);
nand UO_441 (O_441,N_2700,N_2506);
nor UO_442 (O_442,N_2139,N_2695);
or UO_443 (O_443,N_2304,N_2821);
nand UO_444 (O_444,N_2359,N_2820);
nand UO_445 (O_445,N_2459,N_2173);
nand UO_446 (O_446,N_2264,N_2319);
nor UO_447 (O_447,N_2351,N_2952);
and UO_448 (O_448,N_2764,N_2216);
xor UO_449 (O_449,N_2593,N_2734);
or UO_450 (O_450,N_2215,N_2253);
and UO_451 (O_451,N_2687,N_2581);
nor UO_452 (O_452,N_2275,N_2621);
nor UO_453 (O_453,N_2004,N_2491);
nor UO_454 (O_454,N_2031,N_2075);
or UO_455 (O_455,N_2712,N_2636);
nand UO_456 (O_456,N_2488,N_2110);
nor UO_457 (O_457,N_2841,N_2816);
and UO_458 (O_458,N_2224,N_2896);
or UO_459 (O_459,N_2042,N_2737);
and UO_460 (O_460,N_2163,N_2548);
nand UO_461 (O_461,N_2986,N_2658);
and UO_462 (O_462,N_2442,N_2484);
nor UO_463 (O_463,N_2286,N_2365);
nand UO_464 (O_464,N_2471,N_2315);
and UO_465 (O_465,N_2033,N_2629);
nor UO_466 (O_466,N_2323,N_2875);
xor UO_467 (O_467,N_2573,N_2236);
xor UO_468 (O_468,N_2114,N_2415);
nor UO_469 (O_469,N_2385,N_2436);
or UO_470 (O_470,N_2792,N_2632);
and UO_471 (O_471,N_2953,N_2011);
nand UO_472 (O_472,N_2458,N_2855);
or UO_473 (O_473,N_2222,N_2480);
or UO_474 (O_474,N_2054,N_2957);
nor UO_475 (O_475,N_2312,N_2585);
nand UO_476 (O_476,N_2681,N_2185);
nand UO_477 (O_477,N_2016,N_2497);
nor UO_478 (O_478,N_2522,N_2851);
nand UO_479 (O_479,N_2539,N_2300);
xor UO_480 (O_480,N_2449,N_2980);
xnor UO_481 (O_481,N_2538,N_2879);
xnor UO_482 (O_482,N_2795,N_2667);
nor UO_483 (O_483,N_2454,N_2677);
xnor UO_484 (O_484,N_2914,N_2825);
nand UO_485 (O_485,N_2394,N_2333);
and UO_486 (O_486,N_2942,N_2176);
or UO_487 (O_487,N_2753,N_2653);
nand UO_488 (O_488,N_2587,N_2136);
and UO_489 (O_489,N_2897,N_2536);
nor UO_490 (O_490,N_2718,N_2305);
or UO_491 (O_491,N_2407,N_2543);
or UO_492 (O_492,N_2014,N_2201);
nor UO_493 (O_493,N_2034,N_2760);
xor UO_494 (O_494,N_2601,N_2085);
and UO_495 (O_495,N_2515,N_2414);
and UO_496 (O_496,N_2546,N_2423);
xnor UO_497 (O_497,N_2502,N_2272);
nand UO_498 (O_498,N_2148,N_2227);
nand UO_499 (O_499,N_2474,N_2580);
endmodule