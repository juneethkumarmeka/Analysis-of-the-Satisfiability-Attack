module basic_750_5000_1000_2_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2505,N_2507,N_2508,N_2509,N_2510,N_2511,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2524,N_2525,N_2527,N_2528,N_2529,N_2530,N_2531,N_2533,N_2534,N_2536,N_2537,N_2538,N_2540,N_2541,N_2542,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2561,N_2562,N_2563,N_2564,N_2565,N_2567,N_2568,N_2569,N_2574,N_2575,N_2576,N_2577,N_2578,N_2581,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2613,N_2614,N_2615,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2624,N_2626,N_2627,N_2628,N_2630,N_2631,N_2632,N_2633,N_2634,N_2636,N_2637,N_2639,N_2641,N_2642,N_2645,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2659,N_2660,N_2661,N_2662,N_2664,N_2665,N_2666,N_2667,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2687,N_2689,N_2690,N_2691,N_2693,N_2694,N_2695,N_2696,N_2698,N_2699,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2723,N_2724,N_2725,N_2727,N_2728,N_2730,N_2731,N_2732,N_2734,N_2735,N_2736,N_2738,N_2739,N_2740,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2775,N_2776,N_2777,N_2778,N_2780,N_2781,N_2782,N_2785,N_2786,N_2787,N_2788,N_2789,N_2791,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2820,N_2821,N_2823,N_2824,N_2827,N_2829,N_2830,N_2832,N_2833,N_2834,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2847,N_2848,N_2850,N_2851,N_2852,N_2854,N_2856,N_2857,N_2858,N_2859,N_2860,N_2863,N_2864,N_2865,N_2867,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2881,N_2882,N_2884,N_2885,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2906,N_2907,N_2908,N_2909,N_2910,N_2912,N_2913,N_2915,N_2916,N_2917,N_2919,N_2920,N_2921,N_2923,N_2924,N_2925,N_2927,N_2928,N_2929,N_2930,N_2931,N_2933,N_2935,N_2937,N_2938,N_2939,N_2941,N_2942,N_2943,N_2944,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2954,N_2955,N_2956,N_2958,N_2959,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2968,N_2969,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2980,N_2981,N_2982,N_2984,N_2985,N_2988,N_2989,N_2990,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3009,N_3011,N_3013,N_3014,N_3019,N_3020,N_3024,N_3025,N_3026,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3046,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3063,N_3064,N_3065,N_3066,N_3068,N_3069,N_3070,N_3071,N_3074,N_3077,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3088,N_3089,N_3090,N_3091,N_3093,N_3094,N_3096,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3118,N_3119,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3132,N_3133,N_3134,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3152,N_3153,N_3155,N_3156,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3173,N_3174,N_3175,N_3176,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3202,N_3203,N_3205,N_3206,N_3207,N_3208,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3229,N_3230,N_3232,N_3233,N_3234,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3245,N_3246,N_3247,N_3249,N_3250,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3278,N_3279,N_3280,N_3281,N_3283,N_3284,N_3286,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3297,N_3298,N_3299,N_3300,N_3301,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3310,N_3311,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3327,N_3328,N_3330,N_3331,N_3333,N_3334,N_3335,N_3336,N_3337,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3386,N_3389,N_3390,N_3392,N_3395,N_3396,N_3398,N_3399,N_3400,N_3401,N_3402,N_3404,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3425,N_3428,N_3429,N_3430,N_3431,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3443,N_3444,N_3445,N_3446,N_3448,N_3449,N_3450,N_3451,N_3454,N_3455,N_3456,N_3457,N_3459,N_3462,N_3463,N_3464,N_3465,N_3466,N_3468,N_3469,N_3470,N_3473,N_3474,N_3475,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3485,N_3486,N_3487,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3501,N_3502,N_3503,N_3504,N_3507,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3530,N_3531,N_3533,N_3534,N_3536,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3546,N_3547,N_3548,N_3549,N_3550,N_3552,N_3553,N_3555,N_3556,N_3557,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3568,N_3569,N_3570,N_3572,N_3573,N_3575,N_3576,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3627,N_3628,N_3629,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3639,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3651,N_3654,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3666,N_3668,N_3669,N_3671,N_3674,N_3675,N_3676,N_3677,N_3678,N_3680,N_3681,N_3682,N_3683,N_3684,N_3687,N_3688,N_3689,N_3691,N_3693,N_3695,N_3696,N_3697,N_3698,N_3700,N_3701,N_3702,N_3703,N_3704,N_3706,N_3707,N_3708,N_3709,N_3710,N_3712,N_3714,N_3716,N_3717,N_3719,N_3720,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3731,N_3733,N_3734,N_3735,N_3736,N_3737,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3800,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3814,N_3816,N_3817,N_3818,N_3819,N_3820,N_3822,N_3825,N_3827,N_3828,N_3829,N_3830,N_3832,N_3834,N_3835,N_3836,N_3839,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3850,N_3852,N_3853,N_3854,N_3856,N_3857,N_3858,N_3859,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3877,N_3880,N_3881,N_3882,N_3883,N_3884,N_3886,N_3887,N_3888,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3908,N_3909,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3951,N_3955,N_3956,N_3957,N_3958,N_3959,N_3961,N_3962,N_3964,N_3966,N_3969,N_3970,N_3971,N_3972,N_3974,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3993,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4003,N_4004,N_4005,N_4006,N_4009,N_4010,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4021,N_4022,N_4023,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4039,N_4040,N_4042,N_4044,N_4047,N_4048,N_4049,N_4050,N_4052,N_4053,N_4054,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4065,N_4066,N_4068,N_4069,N_4070,N_4072,N_4073,N_4074,N_4076,N_4077,N_4078,N_4079,N_4081,N_4083,N_4084,N_4085,N_4086,N_4088,N_4090,N_4091,N_4093,N_4094,N_4095,N_4096,N_4097,N_4100,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4131,N_4132,N_4133,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4157,N_4158,N_4159,N_4161,N_4162,N_4163,N_4164,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4189,N_4190,N_4192,N_4193,N_4194,N_4196,N_4197,N_4198,N_4199,N_4200,N_4202,N_4203,N_4205,N_4207,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4223,N_4224,N_4225,N_4226,N_4228,N_4229,N_4230,N_4231,N_4233,N_4234,N_4235,N_4239,N_4240,N_4241,N_4242,N_4244,N_4245,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4268,N_4269,N_4270,N_4271,N_4273,N_4276,N_4277,N_4278,N_4279,N_4280,N_4282,N_4283,N_4285,N_4287,N_4290,N_4291,N_4292,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4335,N_4336,N_4337,N_4338,N_4339,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4355,N_4356,N_4357,N_4358,N_4359,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4385,N_4387,N_4388,N_4389,N_4391,N_4392,N_4394,N_4395,N_4396,N_4398,N_4400,N_4401,N_4402,N_4403,N_4404,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4429,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4444,N_4445,N_4448,N_4449,N_4450,N_4451,N_4452,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4461,N_4463,N_4464,N_4466,N_4467,N_4468,N_4469,N_4470,N_4472,N_4473,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4506,N_4507,N_4508,N_4509,N_4510,N_4512,N_4513,N_4514,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4525,N_4527,N_4528,N_4530,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4550,N_4551,N_4553,N_4554,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4563,N_4565,N_4566,N_4568,N_4569,N_4570,N_4571,N_4573,N_4574,N_4575,N_4576,N_4577,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4598,N_4599,N_4600,N_4603,N_4605,N_4606,N_4607,N_4610,N_4611,N_4612,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4667,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4679,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4701,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4723,N_4724,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4737,N_4739,N_4740,N_4742,N_4743,N_4744,N_4745,N_4747,N_4749,N_4750,N_4751,N_4752,N_4753,N_4755,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4772,N_4773,N_4774,N_4775,N_4777,N_4778,N_4780,N_4781,N_4783,N_4784,N_4785,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4803,N_4804,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4814,N_4816,N_4818,N_4819,N_4821,N_4822,N_4823,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4847,N_4850,N_4851,N_4852,N_4853,N_4854,N_4856,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4869,N_4870,N_4872,N_4873,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4891,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4914,N_4916,N_4917,N_4920,N_4921,N_4922,N_4923,N_4926,N_4927,N_4928,N_4931,N_4932,N_4933,N_4935,N_4936,N_4937,N_4938,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4947,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4978,N_4979,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4988,N_4989,N_4990,N_4992,N_4993,N_4994,N_4996,N_4997;
nand U0 (N_0,In_589,In_546);
nand U1 (N_1,In_80,In_490);
nor U2 (N_2,In_729,In_653);
and U3 (N_3,In_498,In_6);
or U4 (N_4,In_15,In_224);
nand U5 (N_5,In_307,In_464);
nor U6 (N_6,In_31,In_372);
nor U7 (N_7,In_209,In_522);
nand U8 (N_8,In_151,In_488);
nand U9 (N_9,In_350,In_302);
nand U10 (N_10,In_555,In_449);
and U11 (N_11,In_171,In_726);
or U12 (N_12,In_698,In_87);
nor U13 (N_13,In_677,In_377);
or U14 (N_14,In_426,In_740);
and U15 (N_15,In_676,In_343);
nor U16 (N_16,In_722,In_651);
nand U17 (N_17,In_406,In_418);
nor U18 (N_18,In_172,In_140);
nor U19 (N_19,In_98,In_571);
nand U20 (N_20,In_413,In_346);
xnor U21 (N_21,In_79,In_491);
nor U22 (N_22,In_743,In_553);
or U23 (N_23,In_8,In_54);
nand U24 (N_24,In_109,In_465);
and U25 (N_25,In_419,In_230);
or U26 (N_26,In_438,In_523);
nor U27 (N_27,In_494,In_430);
nand U28 (N_28,In_388,In_311);
nand U29 (N_29,In_422,In_238);
nand U30 (N_30,In_188,In_431);
nand U31 (N_31,In_414,In_4);
or U32 (N_32,In_310,In_665);
xnor U33 (N_33,In_314,In_683);
xnor U34 (N_34,In_739,In_216);
nor U35 (N_35,In_345,In_349);
and U36 (N_36,In_461,In_253);
nor U37 (N_37,In_301,In_247);
nor U38 (N_38,In_440,In_566);
nor U39 (N_39,In_436,In_703);
and U40 (N_40,In_29,In_374);
nand U41 (N_41,In_549,In_277);
nor U42 (N_42,In_427,In_504);
nor U43 (N_43,In_89,In_381);
and U44 (N_44,In_696,In_386);
nand U45 (N_45,In_398,In_400);
nand U46 (N_46,In_435,In_695);
and U47 (N_47,In_709,In_378);
or U48 (N_48,In_0,In_468);
nand U49 (N_49,In_635,In_579);
nand U50 (N_50,In_68,In_33);
nor U51 (N_51,In_191,In_563);
nand U52 (N_52,In_648,In_126);
or U53 (N_53,In_748,In_691);
nand U54 (N_54,In_46,In_510);
and U55 (N_55,In_581,In_330);
nand U56 (N_56,In_76,In_70);
or U57 (N_57,In_624,In_28);
and U58 (N_58,In_187,In_336);
xor U59 (N_59,In_711,In_530);
nand U60 (N_60,In_533,In_609);
nor U61 (N_61,In_421,In_562);
or U62 (N_62,In_444,In_642);
or U63 (N_63,In_369,In_62);
and U64 (N_64,In_71,In_101);
and U65 (N_65,In_616,In_358);
nand U66 (N_66,In_64,In_282);
or U67 (N_67,In_632,In_316);
xor U68 (N_68,In_652,In_382);
or U69 (N_69,In_561,In_531);
nand U70 (N_70,In_2,In_593);
and U71 (N_71,In_10,In_233);
nor U72 (N_72,In_357,In_700);
nor U73 (N_73,In_161,In_184);
nor U74 (N_74,In_497,In_404);
nor U75 (N_75,In_281,In_737);
and U76 (N_76,In_439,In_567);
xnor U77 (N_77,In_256,In_95);
nand U78 (N_78,In_355,In_99);
nor U79 (N_79,In_305,In_319);
nand U80 (N_80,In_580,In_297);
xnor U81 (N_81,In_170,In_158);
nor U82 (N_82,In_702,In_708);
and U83 (N_83,In_114,In_312);
or U84 (N_84,In_738,In_663);
nand U85 (N_85,In_525,In_644);
or U86 (N_86,In_557,In_452);
and U87 (N_87,In_399,In_543);
nor U88 (N_88,In_218,In_272);
or U89 (N_89,In_463,In_466);
nor U90 (N_90,In_715,In_623);
or U91 (N_91,In_585,In_73);
or U92 (N_92,In_153,In_186);
and U93 (N_93,In_67,In_321);
nand U94 (N_94,In_620,In_239);
xor U95 (N_95,In_598,In_269);
and U96 (N_96,In_385,In_166);
and U97 (N_97,In_617,In_53);
or U98 (N_98,In_169,In_541);
nor U99 (N_99,In_56,In_214);
or U100 (N_100,In_268,In_459);
nand U101 (N_101,In_65,In_469);
or U102 (N_102,In_507,In_627);
nor U103 (N_103,In_621,In_3);
and U104 (N_104,In_402,In_244);
nor U105 (N_105,In_155,In_149);
and U106 (N_106,In_495,In_92);
and U107 (N_107,In_174,In_196);
nor U108 (N_108,In_17,In_118);
and U109 (N_109,In_496,In_123);
nor U110 (N_110,In_606,In_578);
xnor U111 (N_111,In_333,In_594);
and U112 (N_112,In_257,In_403);
nand U113 (N_113,In_441,In_706);
nand U114 (N_114,In_601,In_132);
nand U115 (N_115,In_354,In_394);
and U116 (N_116,In_351,In_639);
or U117 (N_117,In_600,In_163);
nand U118 (N_118,In_285,In_177);
or U119 (N_119,In_237,In_329);
nor U120 (N_120,In_127,In_412);
nor U121 (N_121,In_204,In_542);
and U122 (N_122,In_289,In_582);
nand U123 (N_123,In_707,In_415);
and U124 (N_124,In_667,In_183);
and U125 (N_125,In_456,In_437);
or U126 (N_126,In_339,In_692);
nor U127 (N_127,In_60,In_666);
and U128 (N_128,In_479,In_94);
nor U129 (N_129,In_694,In_558);
and U130 (N_130,In_446,In_270);
nor U131 (N_131,In_524,In_424);
nor U132 (N_132,In_74,In_409);
and U133 (N_133,In_291,In_724);
or U134 (N_134,In_458,In_206);
and U135 (N_135,In_475,In_72);
or U136 (N_136,In_432,In_515);
nor U137 (N_137,In_587,In_150);
and U138 (N_138,In_21,In_656);
nand U139 (N_139,In_210,In_574);
and U140 (N_140,In_408,In_551);
nor U141 (N_141,In_313,In_483);
xnor U142 (N_142,In_117,In_568);
and U143 (N_143,In_411,In_503);
and U144 (N_144,In_128,In_222);
nor U145 (N_145,In_49,In_69);
or U146 (N_146,In_502,In_602);
xor U147 (N_147,In_363,In_19);
nor U148 (N_148,In_539,In_162);
nor U149 (N_149,In_391,In_137);
or U150 (N_150,In_704,In_425);
or U151 (N_151,In_279,In_93);
nand U152 (N_152,In_106,In_520);
or U153 (N_153,In_35,In_607);
xnor U154 (N_154,In_460,In_575);
nand U155 (N_155,In_267,In_544);
nor U156 (N_156,In_716,In_235);
or U157 (N_157,In_178,In_112);
nor U158 (N_158,In_592,In_232);
nor U159 (N_159,In_727,In_489);
and U160 (N_160,In_195,In_241);
xnor U161 (N_161,In_514,In_714);
or U162 (N_162,In_273,In_356);
nand U163 (N_163,In_443,In_130);
nor U164 (N_164,In_323,In_75);
or U165 (N_165,In_455,In_626);
nor U166 (N_166,In_84,In_535);
nand U167 (N_167,In_280,In_110);
and U168 (N_168,In_732,In_608);
or U169 (N_169,In_104,In_517);
or U170 (N_170,In_299,In_344);
and U171 (N_171,In_625,In_317);
or U172 (N_172,In_518,In_143);
or U173 (N_173,In_513,In_682);
and U174 (N_174,In_745,In_529);
nor U175 (N_175,In_451,In_145);
and U176 (N_176,In_293,In_684);
nand U177 (N_177,In_146,In_208);
nor U178 (N_178,In_482,In_560);
or U179 (N_179,In_129,In_105);
or U180 (N_180,In_245,In_227);
nor U181 (N_181,In_338,In_674);
nand U182 (N_182,In_636,In_152);
nand U183 (N_183,In_384,In_261);
or U184 (N_184,In_481,In_113);
nand U185 (N_185,In_348,In_5);
nor U186 (N_186,In_613,In_486);
and U187 (N_187,In_689,In_749);
nor U188 (N_188,In_287,In_182);
nand U189 (N_189,In_295,In_226);
and U190 (N_190,In_326,In_148);
xor U191 (N_191,In_655,In_16);
nand U192 (N_192,In_83,In_645);
nor U193 (N_193,In_243,In_405);
nor U194 (N_194,In_100,In_410);
nand U195 (N_195,In_658,In_20);
and U196 (N_196,In_637,In_548);
nand U197 (N_197,In_618,In_423);
nand U198 (N_198,In_212,In_203);
or U199 (N_199,In_300,In_512);
nand U200 (N_200,In_91,In_526);
nor U201 (N_201,In_612,In_538);
nor U202 (N_202,In_201,In_577);
xor U203 (N_203,In_532,In_379);
nor U204 (N_204,In_116,In_30);
nand U205 (N_205,In_179,In_125);
nand U206 (N_206,In_679,In_556);
nor U207 (N_207,In_559,In_433);
and U208 (N_208,In_198,In_545);
and U209 (N_209,In_688,In_447);
nand U210 (N_210,In_318,In_742);
nand U211 (N_211,In_189,In_131);
or U212 (N_212,In_741,In_687);
nand U213 (N_213,In_366,In_554);
or U214 (N_214,In_629,In_42);
nand U215 (N_215,In_401,In_217);
nor U216 (N_216,In_734,In_485);
nor U217 (N_217,In_640,In_657);
nand U218 (N_218,In_121,In_383);
and U219 (N_219,In_194,In_315);
nor U220 (N_220,In_470,In_678);
or U221 (N_221,In_622,In_120);
or U222 (N_222,In_673,In_202);
and U223 (N_223,In_324,In_133);
or U224 (N_224,In_565,In_111);
nand U225 (N_225,In_180,In_168);
or U226 (N_226,In_597,In_746);
nor U227 (N_227,In_583,In_176);
nor U228 (N_228,In_588,In_511);
nor U229 (N_229,In_659,In_12);
or U230 (N_230,In_25,In_396);
and U231 (N_231,In_649,In_185);
or U232 (N_232,In_51,In_586);
and U233 (N_233,In_86,In_484);
or U234 (N_234,In_718,In_595);
nand U235 (N_235,In_303,In_138);
or U236 (N_236,In_725,In_603);
and U237 (N_237,In_445,In_18);
nor U238 (N_238,In_628,In_521);
and U239 (N_239,In_672,In_50);
nor U240 (N_240,In_24,In_159);
xor U241 (N_241,In_353,In_501);
nand U242 (N_242,In_278,In_453);
and U243 (N_243,In_66,In_1);
or U244 (N_244,In_480,In_611);
or U245 (N_245,In_747,In_728);
and U246 (N_246,In_156,In_699);
or U247 (N_247,In_570,In_175);
and U248 (N_248,In_322,In_154);
or U249 (N_249,In_63,In_685);
and U250 (N_250,In_229,In_646);
and U251 (N_251,In_157,In_32);
nand U252 (N_252,In_610,In_102);
nor U253 (N_253,In_365,In_258);
xnor U254 (N_254,In_442,In_680);
nor U255 (N_255,In_96,In_730);
nor U256 (N_256,In_347,In_368);
xor U257 (N_257,In_234,In_58);
or U258 (N_258,In_454,In_309);
nand U259 (N_259,In_697,In_434);
nand U260 (N_260,In_614,In_670);
nor U261 (N_261,In_228,In_61);
or U262 (N_262,In_360,In_81);
or U263 (N_263,In_219,In_736);
xnor U264 (N_264,In_320,In_527);
nand U265 (N_265,In_342,In_573);
xnor U266 (N_266,In_41,In_43);
xnor U267 (N_267,In_693,In_90);
or U268 (N_268,In_361,In_710);
or U269 (N_269,In_9,In_103);
and U270 (N_270,In_720,In_197);
and U271 (N_271,In_284,In_286);
and U272 (N_272,In_429,In_246);
and U273 (N_273,In_294,In_207);
nand U274 (N_274,In_141,In_599);
nand U275 (N_275,In_242,In_416);
or U276 (N_276,In_373,In_650);
nor U277 (N_277,In_576,In_7);
or U278 (N_278,In_11,In_448);
or U279 (N_279,In_744,In_390);
and U280 (N_280,In_37,In_57);
nor U281 (N_281,In_223,In_263);
or U282 (N_282,In_44,In_248);
and U283 (N_283,In_671,In_662);
or U284 (N_284,In_552,In_370);
xor U285 (N_285,In_254,In_27);
nor U286 (N_286,In_328,In_476);
and U287 (N_287,In_471,In_292);
or U288 (N_288,In_450,In_88);
or U289 (N_289,In_231,In_136);
and U290 (N_290,In_160,In_701);
nor U291 (N_291,In_389,In_251);
and U292 (N_292,In_467,In_547);
and U293 (N_293,In_505,In_509);
xor U294 (N_294,In_135,In_340);
nand U295 (N_295,In_34,In_375);
nor U296 (N_296,In_274,In_306);
nor U297 (N_297,In_55,In_337);
nand U298 (N_298,In_634,In_487);
and U299 (N_299,In_508,In_164);
nor U300 (N_300,In_477,In_221);
nand U301 (N_301,In_631,In_638);
nand U302 (N_302,In_260,In_591);
and U303 (N_303,In_528,In_630);
nand U304 (N_304,In_428,In_265);
nor U305 (N_305,In_516,In_387);
or U306 (N_306,In_457,In_364);
or U307 (N_307,In_534,In_536);
xnor U308 (N_308,In_584,In_499);
xor U309 (N_309,In_376,In_13);
nor U310 (N_310,In_264,In_225);
nand U311 (N_311,In_134,In_647);
or U312 (N_312,In_14,In_52);
nor U313 (N_313,In_167,In_733);
nand U314 (N_314,In_643,In_393);
nand U315 (N_315,In_275,In_712);
and U316 (N_316,In_417,In_331);
nor U317 (N_317,In_619,In_633);
nor U318 (N_318,In_341,In_181);
nand U319 (N_319,In_615,In_537);
nor U320 (N_320,In_38,In_193);
nand U321 (N_321,In_77,In_664);
nand U322 (N_322,In_139,In_142);
or U323 (N_323,In_604,In_669);
or U324 (N_324,In_259,In_407);
nor U325 (N_325,In_641,In_211);
xnor U326 (N_326,In_48,In_506);
and U327 (N_327,In_335,In_500);
nor U328 (N_328,In_271,In_199);
and U329 (N_329,In_173,In_59);
nor U330 (N_330,In_298,In_392);
nand U331 (N_331,In_22,In_240);
nand U332 (N_332,In_283,In_352);
nor U333 (N_333,In_47,In_255);
or U334 (N_334,In_108,In_462);
nand U335 (N_335,In_395,In_540);
nand U336 (N_336,In_200,In_115);
nand U337 (N_337,In_276,In_705);
or U338 (N_338,In_39,In_569);
nor U339 (N_339,In_144,In_367);
nand U340 (N_340,In_721,In_266);
and U341 (N_341,In_23,In_97);
and U342 (N_342,In_686,In_719);
xnor U343 (N_343,In_85,In_107);
and U344 (N_344,In_472,In_735);
and U345 (N_345,In_605,In_675);
nor U346 (N_346,In_36,In_308);
and U347 (N_347,In_288,In_332);
and U348 (N_348,In_474,In_290);
nand U349 (N_349,In_723,In_681);
nor U350 (N_350,In_397,In_717);
and U351 (N_351,In_478,In_78);
nand U352 (N_352,In_190,In_380);
and U353 (N_353,In_250,In_550);
or U354 (N_354,In_492,In_590);
nand U355 (N_355,In_82,In_327);
and U356 (N_356,In_262,In_26);
nand U357 (N_357,In_661,In_147);
or U358 (N_358,In_713,In_124);
xnor U359 (N_359,In_493,In_362);
and U360 (N_360,In_122,In_304);
xor U361 (N_361,In_45,In_473);
and U362 (N_362,In_215,In_420);
xor U363 (N_363,In_296,In_359);
nand U364 (N_364,In_236,In_213);
and U365 (N_365,In_40,In_371);
or U366 (N_366,In_119,In_220);
nand U367 (N_367,In_205,In_192);
or U368 (N_368,In_334,In_564);
nor U369 (N_369,In_654,In_572);
or U370 (N_370,In_690,In_252);
nand U371 (N_371,In_325,In_249);
or U372 (N_372,In_519,In_660);
nand U373 (N_373,In_731,In_668);
and U374 (N_374,In_596,In_165);
nand U375 (N_375,In_541,In_618);
or U376 (N_376,In_394,In_645);
or U377 (N_377,In_422,In_622);
and U378 (N_378,In_135,In_675);
nand U379 (N_379,In_363,In_748);
or U380 (N_380,In_343,In_275);
or U381 (N_381,In_349,In_125);
nor U382 (N_382,In_605,In_698);
nor U383 (N_383,In_191,In_59);
or U384 (N_384,In_507,In_8);
and U385 (N_385,In_284,In_473);
or U386 (N_386,In_338,In_646);
xnor U387 (N_387,In_313,In_726);
and U388 (N_388,In_388,In_316);
xor U389 (N_389,In_378,In_268);
nand U390 (N_390,In_285,In_510);
nor U391 (N_391,In_179,In_581);
and U392 (N_392,In_749,In_550);
and U393 (N_393,In_287,In_738);
nor U394 (N_394,In_507,In_688);
and U395 (N_395,In_526,In_71);
and U396 (N_396,In_366,In_128);
and U397 (N_397,In_531,In_221);
nand U398 (N_398,In_705,In_709);
nor U399 (N_399,In_472,In_24);
nand U400 (N_400,In_79,In_490);
nand U401 (N_401,In_199,In_440);
nor U402 (N_402,In_302,In_0);
and U403 (N_403,In_257,In_276);
and U404 (N_404,In_456,In_749);
nor U405 (N_405,In_482,In_371);
nor U406 (N_406,In_286,In_310);
nor U407 (N_407,In_196,In_360);
xor U408 (N_408,In_393,In_651);
and U409 (N_409,In_704,In_676);
nor U410 (N_410,In_604,In_31);
and U411 (N_411,In_596,In_709);
nor U412 (N_412,In_166,In_105);
or U413 (N_413,In_255,In_96);
nand U414 (N_414,In_41,In_619);
nor U415 (N_415,In_306,In_700);
xnor U416 (N_416,In_573,In_8);
or U417 (N_417,In_360,In_217);
nor U418 (N_418,In_221,In_189);
nor U419 (N_419,In_119,In_724);
nor U420 (N_420,In_665,In_471);
xnor U421 (N_421,In_289,In_732);
and U422 (N_422,In_651,In_605);
nand U423 (N_423,In_530,In_72);
xnor U424 (N_424,In_571,In_485);
and U425 (N_425,In_634,In_655);
nor U426 (N_426,In_151,In_248);
nor U427 (N_427,In_304,In_364);
xnor U428 (N_428,In_541,In_540);
nor U429 (N_429,In_346,In_693);
or U430 (N_430,In_481,In_456);
xnor U431 (N_431,In_241,In_256);
and U432 (N_432,In_74,In_444);
nand U433 (N_433,In_653,In_301);
and U434 (N_434,In_381,In_569);
nor U435 (N_435,In_646,In_748);
or U436 (N_436,In_697,In_109);
and U437 (N_437,In_741,In_306);
and U438 (N_438,In_122,In_187);
nand U439 (N_439,In_119,In_274);
xnor U440 (N_440,In_686,In_348);
and U441 (N_441,In_143,In_636);
nand U442 (N_442,In_4,In_626);
and U443 (N_443,In_513,In_567);
and U444 (N_444,In_4,In_210);
nand U445 (N_445,In_429,In_228);
or U446 (N_446,In_18,In_341);
or U447 (N_447,In_260,In_372);
or U448 (N_448,In_628,In_514);
and U449 (N_449,In_421,In_499);
nor U450 (N_450,In_43,In_438);
nand U451 (N_451,In_386,In_743);
nand U452 (N_452,In_123,In_575);
nand U453 (N_453,In_95,In_449);
and U454 (N_454,In_729,In_436);
or U455 (N_455,In_444,In_78);
and U456 (N_456,In_532,In_428);
or U457 (N_457,In_716,In_144);
nand U458 (N_458,In_602,In_118);
and U459 (N_459,In_342,In_643);
or U460 (N_460,In_11,In_475);
nor U461 (N_461,In_161,In_714);
or U462 (N_462,In_734,In_517);
or U463 (N_463,In_310,In_235);
nand U464 (N_464,In_223,In_520);
or U465 (N_465,In_254,In_216);
or U466 (N_466,In_405,In_481);
nand U467 (N_467,In_112,In_122);
nand U468 (N_468,In_443,In_708);
nor U469 (N_469,In_383,In_478);
or U470 (N_470,In_429,In_284);
xor U471 (N_471,In_483,In_336);
or U472 (N_472,In_323,In_641);
or U473 (N_473,In_616,In_726);
nand U474 (N_474,In_424,In_144);
or U475 (N_475,In_202,In_123);
or U476 (N_476,In_435,In_492);
nand U477 (N_477,In_297,In_285);
or U478 (N_478,In_110,In_667);
xnor U479 (N_479,In_721,In_29);
or U480 (N_480,In_349,In_410);
and U481 (N_481,In_268,In_392);
xnor U482 (N_482,In_357,In_618);
and U483 (N_483,In_233,In_659);
nand U484 (N_484,In_727,In_332);
nor U485 (N_485,In_300,In_749);
nand U486 (N_486,In_365,In_9);
nor U487 (N_487,In_458,In_237);
nand U488 (N_488,In_166,In_612);
nand U489 (N_489,In_745,In_553);
nand U490 (N_490,In_623,In_578);
or U491 (N_491,In_88,In_87);
nor U492 (N_492,In_65,In_112);
and U493 (N_493,In_740,In_385);
and U494 (N_494,In_324,In_190);
nor U495 (N_495,In_327,In_604);
nand U496 (N_496,In_729,In_542);
and U497 (N_497,In_123,In_5);
or U498 (N_498,In_192,In_141);
or U499 (N_499,In_40,In_642);
nor U500 (N_500,In_273,In_77);
xor U501 (N_501,In_671,In_403);
or U502 (N_502,In_416,In_602);
or U503 (N_503,In_412,In_95);
xor U504 (N_504,In_641,In_749);
nor U505 (N_505,In_396,In_403);
nor U506 (N_506,In_168,In_581);
nand U507 (N_507,In_741,In_656);
nand U508 (N_508,In_138,In_132);
and U509 (N_509,In_602,In_739);
and U510 (N_510,In_266,In_533);
and U511 (N_511,In_320,In_285);
and U512 (N_512,In_592,In_746);
nand U513 (N_513,In_141,In_133);
nand U514 (N_514,In_181,In_14);
or U515 (N_515,In_48,In_502);
xor U516 (N_516,In_165,In_427);
nor U517 (N_517,In_228,In_98);
or U518 (N_518,In_667,In_271);
xnor U519 (N_519,In_615,In_8);
or U520 (N_520,In_532,In_435);
and U521 (N_521,In_359,In_32);
nand U522 (N_522,In_247,In_239);
nor U523 (N_523,In_488,In_439);
nor U524 (N_524,In_265,In_75);
or U525 (N_525,In_127,In_337);
nor U526 (N_526,In_745,In_508);
or U527 (N_527,In_356,In_238);
nand U528 (N_528,In_200,In_272);
or U529 (N_529,In_293,In_291);
and U530 (N_530,In_51,In_707);
and U531 (N_531,In_522,In_610);
and U532 (N_532,In_555,In_468);
nand U533 (N_533,In_133,In_169);
nor U534 (N_534,In_115,In_371);
nand U535 (N_535,In_309,In_235);
nand U536 (N_536,In_15,In_232);
or U537 (N_537,In_455,In_505);
or U538 (N_538,In_627,In_85);
nand U539 (N_539,In_97,In_659);
nand U540 (N_540,In_269,In_741);
nor U541 (N_541,In_15,In_41);
or U542 (N_542,In_187,In_519);
nor U543 (N_543,In_306,In_707);
and U544 (N_544,In_676,In_680);
or U545 (N_545,In_357,In_695);
nor U546 (N_546,In_69,In_310);
nor U547 (N_547,In_414,In_619);
and U548 (N_548,In_674,In_408);
nand U549 (N_549,In_118,In_224);
and U550 (N_550,In_180,In_122);
nand U551 (N_551,In_2,In_313);
and U552 (N_552,In_163,In_93);
nand U553 (N_553,In_377,In_655);
or U554 (N_554,In_668,In_392);
xor U555 (N_555,In_333,In_155);
and U556 (N_556,In_744,In_623);
xnor U557 (N_557,In_742,In_353);
and U558 (N_558,In_151,In_67);
nor U559 (N_559,In_249,In_673);
and U560 (N_560,In_519,In_16);
nor U561 (N_561,In_343,In_730);
and U562 (N_562,In_647,In_286);
or U563 (N_563,In_537,In_683);
nand U564 (N_564,In_65,In_257);
nand U565 (N_565,In_311,In_587);
nand U566 (N_566,In_193,In_545);
and U567 (N_567,In_24,In_256);
xnor U568 (N_568,In_561,In_79);
or U569 (N_569,In_434,In_149);
nand U570 (N_570,In_291,In_111);
or U571 (N_571,In_165,In_581);
xnor U572 (N_572,In_742,In_367);
and U573 (N_573,In_599,In_358);
nand U574 (N_574,In_451,In_657);
or U575 (N_575,In_30,In_433);
nand U576 (N_576,In_94,In_292);
and U577 (N_577,In_431,In_455);
xor U578 (N_578,In_679,In_89);
nand U579 (N_579,In_554,In_668);
nor U580 (N_580,In_647,In_45);
or U581 (N_581,In_604,In_243);
and U582 (N_582,In_439,In_572);
nor U583 (N_583,In_552,In_499);
xor U584 (N_584,In_604,In_385);
xnor U585 (N_585,In_692,In_95);
and U586 (N_586,In_321,In_273);
nand U587 (N_587,In_401,In_91);
nand U588 (N_588,In_79,In_173);
nor U589 (N_589,In_259,In_366);
xor U590 (N_590,In_481,In_78);
or U591 (N_591,In_590,In_454);
nor U592 (N_592,In_279,In_439);
or U593 (N_593,In_76,In_410);
nor U594 (N_594,In_616,In_674);
nor U595 (N_595,In_143,In_435);
or U596 (N_596,In_171,In_443);
or U597 (N_597,In_479,In_681);
or U598 (N_598,In_247,In_571);
nor U599 (N_599,In_59,In_732);
or U600 (N_600,In_321,In_557);
nand U601 (N_601,In_15,In_249);
and U602 (N_602,In_572,In_9);
nor U603 (N_603,In_567,In_270);
nand U604 (N_604,In_68,In_736);
or U605 (N_605,In_564,In_558);
or U606 (N_606,In_672,In_400);
and U607 (N_607,In_599,In_662);
and U608 (N_608,In_180,In_251);
nor U609 (N_609,In_719,In_578);
and U610 (N_610,In_502,In_352);
nand U611 (N_611,In_558,In_309);
nand U612 (N_612,In_516,In_329);
or U613 (N_613,In_332,In_411);
and U614 (N_614,In_669,In_565);
nand U615 (N_615,In_714,In_143);
nand U616 (N_616,In_35,In_120);
or U617 (N_617,In_90,In_326);
nor U618 (N_618,In_431,In_89);
or U619 (N_619,In_272,In_38);
xnor U620 (N_620,In_196,In_435);
nor U621 (N_621,In_658,In_687);
nor U622 (N_622,In_652,In_330);
nand U623 (N_623,In_661,In_110);
nand U624 (N_624,In_740,In_450);
and U625 (N_625,In_681,In_637);
nor U626 (N_626,In_663,In_365);
nand U627 (N_627,In_91,In_170);
nand U628 (N_628,In_440,In_187);
nand U629 (N_629,In_714,In_686);
nand U630 (N_630,In_651,In_683);
and U631 (N_631,In_83,In_665);
nor U632 (N_632,In_642,In_677);
nor U633 (N_633,In_588,In_631);
xnor U634 (N_634,In_494,In_100);
and U635 (N_635,In_400,In_582);
nor U636 (N_636,In_507,In_709);
and U637 (N_637,In_411,In_598);
and U638 (N_638,In_477,In_48);
or U639 (N_639,In_636,In_386);
nor U640 (N_640,In_526,In_37);
nor U641 (N_641,In_146,In_42);
or U642 (N_642,In_271,In_15);
nand U643 (N_643,In_489,In_49);
nand U644 (N_644,In_549,In_109);
nand U645 (N_645,In_4,In_427);
nor U646 (N_646,In_600,In_269);
and U647 (N_647,In_652,In_185);
nand U648 (N_648,In_733,In_4);
and U649 (N_649,In_194,In_20);
and U650 (N_650,In_551,In_517);
and U651 (N_651,In_699,In_362);
nor U652 (N_652,In_626,In_59);
or U653 (N_653,In_113,In_287);
nor U654 (N_654,In_651,In_645);
or U655 (N_655,In_551,In_133);
or U656 (N_656,In_328,In_142);
and U657 (N_657,In_310,In_223);
or U658 (N_658,In_669,In_481);
nor U659 (N_659,In_496,In_480);
or U660 (N_660,In_587,In_208);
or U661 (N_661,In_509,In_201);
nor U662 (N_662,In_187,In_735);
nor U663 (N_663,In_501,In_428);
or U664 (N_664,In_115,In_56);
nand U665 (N_665,In_99,In_407);
or U666 (N_666,In_104,In_22);
xnor U667 (N_667,In_620,In_24);
nand U668 (N_668,In_60,In_207);
nand U669 (N_669,In_239,In_263);
nor U670 (N_670,In_198,In_413);
or U671 (N_671,In_351,In_369);
nand U672 (N_672,In_383,In_110);
or U673 (N_673,In_344,In_590);
nor U674 (N_674,In_436,In_480);
or U675 (N_675,In_419,In_675);
nor U676 (N_676,In_737,In_221);
nand U677 (N_677,In_246,In_271);
or U678 (N_678,In_646,In_213);
or U679 (N_679,In_742,In_340);
or U680 (N_680,In_473,In_573);
nand U681 (N_681,In_729,In_274);
or U682 (N_682,In_511,In_550);
or U683 (N_683,In_328,In_96);
nand U684 (N_684,In_586,In_468);
nor U685 (N_685,In_389,In_34);
nor U686 (N_686,In_79,In_700);
or U687 (N_687,In_586,In_448);
nand U688 (N_688,In_398,In_45);
or U689 (N_689,In_200,In_280);
nor U690 (N_690,In_323,In_311);
and U691 (N_691,In_38,In_532);
or U692 (N_692,In_606,In_717);
xnor U693 (N_693,In_172,In_386);
nand U694 (N_694,In_567,In_617);
nand U695 (N_695,In_616,In_509);
and U696 (N_696,In_367,In_136);
or U697 (N_697,In_514,In_612);
xor U698 (N_698,In_192,In_478);
or U699 (N_699,In_702,In_334);
xor U700 (N_700,In_314,In_245);
and U701 (N_701,In_103,In_523);
or U702 (N_702,In_643,In_515);
xor U703 (N_703,In_579,In_667);
and U704 (N_704,In_429,In_83);
nor U705 (N_705,In_513,In_50);
nand U706 (N_706,In_446,In_186);
or U707 (N_707,In_347,In_173);
and U708 (N_708,In_687,In_225);
nor U709 (N_709,In_653,In_484);
xnor U710 (N_710,In_2,In_226);
nor U711 (N_711,In_749,In_568);
and U712 (N_712,In_543,In_305);
or U713 (N_713,In_423,In_295);
or U714 (N_714,In_691,In_428);
xnor U715 (N_715,In_7,In_575);
and U716 (N_716,In_254,In_358);
and U717 (N_717,In_287,In_110);
and U718 (N_718,In_487,In_411);
nor U719 (N_719,In_595,In_636);
nor U720 (N_720,In_723,In_482);
nand U721 (N_721,In_566,In_86);
or U722 (N_722,In_556,In_476);
and U723 (N_723,In_682,In_28);
nor U724 (N_724,In_2,In_330);
or U725 (N_725,In_614,In_348);
nor U726 (N_726,In_269,In_446);
nand U727 (N_727,In_660,In_8);
or U728 (N_728,In_391,In_467);
or U729 (N_729,In_364,In_205);
or U730 (N_730,In_536,In_235);
and U731 (N_731,In_159,In_170);
xor U732 (N_732,In_287,In_640);
or U733 (N_733,In_291,In_81);
nand U734 (N_734,In_246,In_700);
nor U735 (N_735,In_620,In_672);
and U736 (N_736,In_362,In_262);
and U737 (N_737,In_296,In_15);
nor U738 (N_738,In_367,In_476);
nor U739 (N_739,In_508,In_320);
and U740 (N_740,In_56,In_203);
nor U741 (N_741,In_2,In_139);
nor U742 (N_742,In_547,In_447);
and U743 (N_743,In_746,In_344);
nand U744 (N_744,In_375,In_176);
xor U745 (N_745,In_195,In_3);
xor U746 (N_746,In_334,In_441);
and U747 (N_747,In_174,In_388);
nand U748 (N_748,In_649,In_187);
nor U749 (N_749,In_432,In_224);
nand U750 (N_750,In_581,In_118);
nor U751 (N_751,In_146,In_588);
nor U752 (N_752,In_535,In_452);
or U753 (N_753,In_467,In_710);
or U754 (N_754,In_156,In_728);
and U755 (N_755,In_743,In_703);
xnor U756 (N_756,In_430,In_480);
and U757 (N_757,In_222,In_570);
and U758 (N_758,In_194,In_203);
or U759 (N_759,In_43,In_289);
nand U760 (N_760,In_674,In_383);
nor U761 (N_761,In_668,In_80);
nor U762 (N_762,In_595,In_694);
nand U763 (N_763,In_565,In_505);
or U764 (N_764,In_15,In_656);
nor U765 (N_765,In_452,In_134);
and U766 (N_766,In_611,In_106);
nand U767 (N_767,In_500,In_162);
or U768 (N_768,In_514,In_718);
xnor U769 (N_769,In_25,In_747);
or U770 (N_770,In_721,In_296);
or U771 (N_771,In_720,In_614);
nand U772 (N_772,In_677,In_308);
nand U773 (N_773,In_528,In_335);
nand U774 (N_774,In_196,In_564);
and U775 (N_775,In_489,In_633);
nand U776 (N_776,In_509,In_740);
and U777 (N_777,In_743,In_393);
nor U778 (N_778,In_676,In_146);
nand U779 (N_779,In_382,In_179);
or U780 (N_780,In_696,In_246);
and U781 (N_781,In_514,In_9);
and U782 (N_782,In_4,In_550);
and U783 (N_783,In_146,In_240);
nand U784 (N_784,In_53,In_512);
or U785 (N_785,In_417,In_713);
and U786 (N_786,In_348,In_413);
and U787 (N_787,In_119,In_643);
nor U788 (N_788,In_729,In_237);
or U789 (N_789,In_234,In_143);
nand U790 (N_790,In_216,In_267);
and U791 (N_791,In_217,In_33);
nand U792 (N_792,In_351,In_677);
or U793 (N_793,In_109,In_374);
and U794 (N_794,In_189,In_414);
and U795 (N_795,In_293,In_236);
xor U796 (N_796,In_522,In_259);
nor U797 (N_797,In_230,In_560);
and U798 (N_798,In_266,In_59);
nor U799 (N_799,In_306,In_689);
or U800 (N_800,In_56,In_24);
xor U801 (N_801,In_316,In_438);
nor U802 (N_802,In_527,In_196);
or U803 (N_803,In_19,In_247);
or U804 (N_804,In_416,In_269);
or U805 (N_805,In_423,In_619);
and U806 (N_806,In_210,In_265);
or U807 (N_807,In_269,In_721);
or U808 (N_808,In_336,In_689);
nand U809 (N_809,In_397,In_425);
nand U810 (N_810,In_223,In_667);
nand U811 (N_811,In_21,In_379);
nand U812 (N_812,In_470,In_87);
and U813 (N_813,In_236,In_672);
nor U814 (N_814,In_612,In_154);
nor U815 (N_815,In_566,In_127);
or U816 (N_816,In_3,In_121);
or U817 (N_817,In_741,In_59);
nor U818 (N_818,In_695,In_598);
xnor U819 (N_819,In_617,In_315);
nand U820 (N_820,In_161,In_288);
nand U821 (N_821,In_186,In_675);
nor U822 (N_822,In_402,In_516);
nor U823 (N_823,In_722,In_746);
or U824 (N_824,In_624,In_567);
and U825 (N_825,In_716,In_545);
xnor U826 (N_826,In_147,In_167);
and U827 (N_827,In_723,In_85);
nor U828 (N_828,In_503,In_117);
or U829 (N_829,In_644,In_427);
nor U830 (N_830,In_20,In_591);
and U831 (N_831,In_289,In_404);
nand U832 (N_832,In_213,In_707);
or U833 (N_833,In_6,In_287);
nor U834 (N_834,In_699,In_495);
nand U835 (N_835,In_502,In_271);
or U836 (N_836,In_485,In_545);
nor U837 (N_837,In_221,In_281);
nand U838 (N_838,In_632,In_114);
or U839 (N_839,In_370,In_672);
or U840 (N_840,In_638,In_635);
nor U841 (N_841,In_657,In_704);
or U842 (N_842,In_487,In_216);
or U843 (N_843,In_686,In_73);
nand U844 (N_844,In_563,In_124);
xnor U845 (N_845,In_688,In_61);
nor U846 (N_846,In_119,In_621);
nor U847 (N_847,In_491,In_653);
or U848 (N_848,In_357,In_567);
and U849 (N_849,In_266,In_735);
or U850 (N_850,In_183,In_10);
nand U851 (N_851,In_479,In_324);
nand U852 (N_852,In_746,In_602);
or U853 (N_853,In_537,In_653);
or U854 (N_854,In_384,In_220);
nand U855 (N_855,In_465,In_300);
nor U856 (N_856,In_692,In_360);
nor U857 (N_857,In_462,In_638);
and U858 (N_858,In_6,In_699);
nand U859 (N_859,In_680,In_221);
nor U860 (N_860,In_6,In_560);
and U861 (N_861,In_698,In_143);
and U862 (N_862,In_90,In_151);
nand U863 (N_863,In_669,In_733);
or U864 (N_864,In_579,In_664);
nor U865 (N_865,In_644,In_625);
or U866 (N_866,In_570,In_170);
nand U867 (N_867,In_183,In_537);
and U868 (N_868,In_681,In_534);
nor U869 (N_869,In_635,In_132);
and U870 (N_870,In_697,In_253);
nor U871 (N_871,In_341,In_709);
nor U872 (N_872,In_211,In_576);
or U873 (N_873,In_429,In_404);
nor U874 (N_874,In_673,In_595);
or U875 (N_875,In_444,In_55);
and U876 (N_876,In_705,In_564);
nand U877 (N_877,In_225,In_721);
and U878 (N_878,In_75,In_293);
or U879 (N_879,In_708,In_346);
and U880 (N_880,In_94,In_165);
nor U881 (N_881,In_654,In_131);
and U882 (N_882,In_670,In_602);
and U883 (N_883,In_508,In_196);
and U884 (N_884,In_444,In_248);
and U885 (N_885,In_705,In_333);
nand U886 (N_886,In_156,In_52);
and U887 (N_887,In_272,In_706);
or U888 (N_888,In_582,In_288);
and U889 (N_889,In_406,In_350);
and U890 (N_890,In_185,In_319);
nand U891 (N_891,In_37,In_206);
or U892 (N_892,In_51,In_34);
or U893 (N_893,In_663,In_473);
xor U894 (N_894,In_165,In_148);
xnor U895 (N_895,In_300,In_27);
xor U896 (N_896,In_725,In_82);
or U897 (N_897,In_155,In_482);
nand U898 (N_898,In_258,In_59);
or U899 (N_899,In_394,In_484);
nor U900 (N_900,In_489,In_541);
nor U901 (N_901,In_393,In_162);
nor U902 (N_902,In_721,In_604);
or U903 (N_903,In_574,In_625);
nand U904 (N_904,In_682,In_173);
xnor U905 (N_905,In_414,In_250);
and U906 (N_906,In_492,In_108);
and U907 (N_907,In_705,In_463);
nand U908 (N_908,In_394,In_559);
nand U909 (N_909,In_688,In_529);
nand U910 (N_910,In_81,In_562);
xor U911 (N_911,In_494,In_527);
and U912 (N_912,In_203,In_368);
nor U913 (N_913,In_617,In_602);
xnor U914 (N_914,In_620,In_68);
or U915 (N_915,In_75,In_232);
or U916 (N_916,In_539,In_727);
or U917 (N_917,In_304,In_240);
xnor U918 (N_918,In_455,In_232);
nor U919 (N_919,In_462,In_571);
nor U920 (N_920,In_505,In_323);
nor U921 (N_921,In_129,In_23);
and U922 (N_922,In_552,In_411);
xnor U923 (N_923,In_604,In_36);
nor U924 (N_924,In_484,In_734);
and U925 (N_925,In_550,In_117);
or U926 (N_926,In_38,In_637);
nor U927 (N_927,In_638,In_519);
and U928 (N_928,In_7,In_327);
xnor U929 (N_929,In_341,In_95);
nor U930 (N_930,In_674,In_685);
nand U931 (N_931,In_475,In_722);
nor U932 (N_932,In_22,In_228);
nor U933 (N_933,In_215,In_105);
and U934 (N_934,In_641,In_56);
nand U935 (N_935,In_303,In_312);
nand U936 (N_936,In_216,In_544);
and U937 (N_937,In_570,In_711);
nor U938 (N_938,In_485,In_716);
xnor U939 (N_939,In_320,In_350);
nor U940 (N_940,In_227,In_144);
and U941 (N_941,In_265,In_298);
nor U942 (N_942,In_708,In_186);
nor U943 (N_943,In_722,In_358);
nor U944 (N_944,In_146,In_484);
or U945 (N_945,In_132,In_395);
and U946 (N_946,In_500,In_691);
or U947 (N_947,In_600,In_522);
nand U948 (N_948,In_233,In_485);
and U949 (N_949,In_733,In_116);
and U950 (N_950,In_424,In_520);
nand U951 (N_951,In_425,In_536);
or U952 (N_952,In_53,In_151);
nand U953 (N_953,In_681,In_225);
nand U954 (N_954,In_113,In_698);
nor U955 (N_955,In_108,In_113);
nand U956 (N_956,In_661,In_298);
nand U957 (N_957,In_38,In_37);
nand U958 (N_958,In_231,In_266);
or U959 (N_959,In_250,In_381);
and U960 (N_960,In_333,In_540);
nor U961 (N_961,In_667,In_487);
or U962 (N_962,In_664,In_244);
and U963 (N_963,In_468,In_512);
or U964 (N_964,In_208,In_707);
or U965 (N_965,In_387,In_616);
or U966 (N_966,In_708,In_39);
or U967 (N_967,In_436,In_243);
nand U968 (N_968,In_306,In_406);
nand U969 (N_969,In_546,In_681);
or U970 (N_970,In_266,In_503);
xor U971 (N_971,In_46,In_196);
and U972 (N_972,In_527,In_576);
and U973 (N_973,In_27,In_342);
nand U974 (N_974,In_736,In_677);
and U975 (N_975,In_723,In_634);
and U976 (N_976,In_697,In_110);
nand U977 (N_977,In_474,In_372);
or U978 (N_978,In_32,In_396);
nand U979 (N_979,In_289,In_652);
or U980 (N_980,In_193,In_551);
and U981 (N_981,In_562,In_234);
nand U982 (N_982,In_129,In_668);
nand U983 (N_983,In_357,In_148);
nand U984 (N_984,In_281,In_397);
and U985 (N_985,In_657,In_528);
nand U986 (N_986,In_1,In_601);
and U987 (N_987,In_339,In_564);
nand U988 (N_988,In_693,In_511);
or U989 (N_989,In_87,In_271);
or U990 (N_990,In_408,In_403);
and U991 (N_991,In_638,In_228);
nor U992 (N_992,In_6,In_533);
xnor U993 (N_993,In_576,In_640);
or U994 (N_994,In_170,In_39);
nor U995 (N_995,In_42,In_452);
and U996 (N_996,In_451,In_687);
or U997 (N_997,In_532,In_205);
xnor U998 (N_998,In_528,In_512);
or U999 (N_999,In_567,In_482);
or U1000 (N_1000,In_494,In_641);
or U1001 (N_1001,In_642,In_213);
or U1002 (N_1002,In_567,In_479);
nor U1003 (N_1003,In_420,In_560);
or U1004 (N_1004,In_643,In_414);
nand U1005 (N_1005,In_129,In_347);
and U1006 (N_1006,In_677,In_474);
and U1007 (N_1007,In_43,In_681);
or U1008 (N_1008,In_511,In_439);
and U1009 (N_1009,In_32,In_466);
and U1010 (N_1010,In_111,In_733);
nand U1011 (N_1011,In_355,In_687);
nand U1012 (N_1012,In_336,In_105);
or U1013 (N_1013,In_351,In_222);
or U1014 (N_1014,In_505,In_564);
xnor U1015 (N_1015,In_327,In_101);
nor U1016 (N_1016,In_550,In_549);
nor U1017 (N_1017,In_11,In_129);
xor U1018 (N_1018,In_50,In_682);
nor U1019 (N_1019,In_661,In_219);
nor U1020 (N_1020,In_373,In_555);
xor U1021 (N_1021,In_647,In_226);
or U1022 (N_1022,In_98,In_386);
nand U1023 (N_1023,In_475,In_706);
and U1024 (N_1024,In_435,In_202);
nor U1025 (N_1025,In_247,In_13);
and U1026 (N_1026,In_640,In_631);
or U1027 (N_1027,In_682,In_493);
nand U1028 (N_1028,In_106,In_53);
and U1029 (N_1029,In_382,In_129);
nand U1030 (N_1030,In_147,In_169);
xnor U1031 (N_1031,In_93,In_65);
nor U1032 (N_1032,In_650,In_273);
nor U1033 (N_1033,In_654,In_13);
and U1034 (N_1034,In_674,In_668);
nor U1035 (N_1035,In_495,In_477);
and U1036 (N_1036,In_566,In_53);
nor U1037 (N_1037,In_660,In_279);
or U1038 (N_1038,In_237,In_734);
xor U1039 (N_1039,In_202,In_397);
nand U1040 (N_1040,In_443,In_471);
nand U1041 (N_1041,In_48,In_418);
nand U1042 (N_1042,In_482,In_622);
nand U1043 (N_1043,In_288,In_407);
nand U1044 (N_1044,In_417,In_370);
nand U1045 (N_1045,In_120,In_500);
and U1046 (N_1046,In_701,In_133);
and U1047 (N_1047,In_298,In_21);
or U1048 (N_1048,In_688,In_101);
nand U1049 (N_1049,In_183,In_635);
or U1050 (N_1050,In_688,In_745);
nor U1051 (N_1051,In_668,In_316);
or U1052 (N_1052,In_176,In_697);
and U1053 (N_1053,In_384,In_441);
xnor U1054 (N_1054,In_610,In_431);
nand U1055 (N_1055,In_568,In_82);
or U1056 (N_1056,In_291,In_485);
or U1057 (N_1057,In_360,In_393);
or U1058 (N_1058,In_737,In_344);
and U1059 (N_1059,In_595,In_533);
or U1060 (N_1060,In_122,In_459);
nor U1061 (N_1061,In_50,In_345);
or U1062 (N_1062,In_67,In_164);
and U1063 (N_1063,In_120,In_397);
nand U1064 (N_1064,In_206,In_480);
or U1065 (N_1065,In_600,In_744);
nor U1066 (N_1066,In_551,In_613);
nor U1067 (N_1067,In_609,In_486);
nor U1068 (N_1068,In_137,In_56);
nor U1069 (N_1069,In_736,In_731);
and U1070 (N_1070,In_120,In_418);
and U1071 (N_1071,In_549,In_489);
xnor U1072 (N_1072,In_450,In_176);
and U1073 (N_1073,In_222,In_490);
nor U1074 (N_1074,In_489,In_140);
and U1075 (N_1075,In_104,In_140);
xnor U1076 (N_1076,In_511,In_563);
nand U1077 (N_1077,In_143,In_384);
nand U1078 (N_1078,In_573,In_486);
or U1079 (N_1079,In_319,In_174);
xnor U1080 (N_1080,In_548,In_578);
and U1081 (N_1081,In_270,In_22);
and U1082 (N_1082,In_550,In_123);
nor U1083 (N_1083,In_227,In_281);
and U1084 (N_1084,In_332,In_360);
or U1085 (N_1085,In_689,In_61);
nor U1086 (N_1086,In_284,In_305);
and U1087 (N_1087,In_446,In_435);
nand U1088 (N_1088,In_123,In_607);
xor U1089 (N_1089,In_425,In_705);
nand U1090 (N_1090,In_621,In_251);
and U1091 (N_1091,In_643,In_304);
and U1092 (N_1092,In_611,In_114);
and U1093 (N_1093,In_683,In_207);
or U1094 (N_1094,In_520,In_299);
or U1095 (N_1095,In_730,In_398);
nand U1096 (N_1096,In_655,In_8);
nand U1097 (N_1097,In_470,In_54);
or U1098 (N_1098,In_209,In_186);
xor U1099 (N_1099,In_303,In_212);
nand U1100 (N_1100,In_174,In_151);
nor U1101 (N_1101,In_727,In_39);
nand U1102 (N_1102,In_192,In_547);
nand U1103 (N_1103,In_233,In_213);
nor U1104 (N_1104,In_153,In_517);
nor U1105 (N_1105,In_585,In_293);
or U1106 (N_1106,In_279,In_423);
nor U1107 (N_1107,In_658,In_733);
nand U1108 (N_1108,In_89,In_418);
nand U1109 (N_1109,In_551,In_162);
and U1110 (N_1110,In_546,In_257);
nor U1111 (N_1111,In_113,In_400);
nor U1112 (N_1112,In_136,In_515);
or U1113 (N_1113,In_24,In_437);
nor U1114 (N_1114,In_603,In_235);
and U1115 (N_1115,In_494,In_225);
and U1116 (N_1116,In_249,In_715);
or U1117 (N_1117,In_297,In_35);
nand U1118 (N_1118,In_329,In_411);
or U1119 (N_1119,In_410,In_738);
or U1120 (N_1120,In_532,In_617);
nor U1121 (N_1121,In_539,In_550);
nand U1122 (N_1122,In_218,In_520);
or U1123 (N_1123,In_635,In_257);
nor U1124 (N_1124,In_505,In_350);
nand U1125 (N_1125,In_454,In_361);
or U1126 (N_1126,In_532,In_706);
nand U1127 (N_1127,In_202,In_326);
nor U1128 (N_1128,In_410,In_744);
nor U1129 (N_1129,In_352,In_547);
and U1130 (N_1130,In_274,In_531);
nor U1131 (N_1131,In_271,In_467);
and U1132 (N_1132,In_277,In_102);
and U1133 (N_1133,In_268,In_692);
nand U1134 (N_1134,In_80,In_144);
nor U1135 (N_1135,In_176,In_65);
nand U1136 (N_1136,In_582,In_424);
xor U1137 (N_1137,In_516,In_462);
nor U1138 (N_1138,In_602,In_27);
nand U1139 (N_1139,In_722,In_342);
and U1140 (N_1140,In_385,In_159);
and U1141 (N_1141,In_674,In_494);
and U1142 (N_1142,In_332,In_1);
and U1143 (N_1143,In_684,In_342);
and U1144 (N_1144,In_602,In_532);
nand U1145 (N_1145,In_301,In_47);
and U1146 (N_1146,In_203,In_447);
nor U1147 (N_1147,In_265,In_22);
xnor U1148 (N_1148,In_598,In_579);
nand U1149 (N_1149,In_519,In_65);
and U1150 (N_1150,In_208,In_334);
nor U1151 (N_1151,In_578,In_124);
nand U1152 (N_1152,In_338,In_578);
nor U1153 (N_1153,In_164,In_152);
xnor U1154 (N_1154,In_272,In_393);
and U1155 (N_1155,In_580,In_544);
nor U1156 (N_1156,In_32,In_374);
and U1157 (N_1157,In_451,In_101);
or U1158 (N_1158,In_159,In_274);
nand U1159 (N_1159,In_712,In_588);
nand U1160 (N_1160,In_92,In_520);
and U1161 (N_1161,In_544,In_537);
or U1162 (N_1162,In_746,In_496);
or U1163 (N_1163,In_25,In_454);
or U1164 (N_1164,In_460,In_48);
xor U1165 (N_1165,In_632,In_260);
nor U1166 (N_1166,In_93,In_384);
nor U1167 (N_1167,In_377,In_699);
or U1168 (N_1168,In_11,In_337);
or U1169 (N_1169,In_417,In_175);
nand U1170 (N_1170,In_722,In_532);
or U1171 (N_1171,In_283,In_431);
and U1172 (N_1172,In_65,In_742);
or U1173 (N_1173,In_493,In_29);
or U1174 (N_1174,In_385,In_524);
nor U1175 (N_1175,In_654,In_630);
nor U1176 (N_1176,In_213,In_262);
xnor U1177 (N_1177,In_452,In_37);
and U1178 (N_1178,In_39,In_18);
and U1179 (N_1179,In_577,In_419);
nor U1180 (N_1180,In_518,In_94);
and U1181 (N_1181,In_244,In_439);
or U1182 (N_1182,In_629,In_604);
and U1183 (N_1183,In_150,In_517);
and U1184 (N_1184,In_115,In_708);
and U1185 (N_1185,In_129,In_315);
nor U1186 (N_1186,In_92,In_370);
nand U1187 (N_1187,In_465,In_583);
xnor U1188 (N_1188,In_51,In_136);
nor U1189 (N_1189,In_671,In_324);
or U1190 (N_1190,In_400,In_154);
nor U1191 (N_1191,In_438,In_126);
and U1192 (N_1192,In_283,In_712);
and U1193 (N_1193,In_305,In_478);
nand U1194 (N_1194,In_465,In_649);
nor U1195 (N_1195,In_179,In_72);
nor U1196 (N_1196,In_245,In_404);
nand U1197 (N_1197,In_99,In_660);
and U1198 (N_1198,In_204,In_213);
nand U1199 (N_1199,In_233,In_400);
nor U1200 (N_1200,In_339,In_552);
nand U1201 (N_1201,In_14,In_436);
or U1202 (N_1202,In_23,In_405);
and U1203 (N_1203,In_428,In_402);
nor U1204 (N_1204,In_698,In_739);
nor U1205 (N_1205,In_42,In_37);
and U1206 (N_1206,In_293,In_9);
and U1207 (N_1207,In_456,In_391);
or U1208 (N_1208,In_70,In_456);
xor U1209 (N_1209,In_10,In_681);
nand U1210 (N_1210,In_622,In_714);
or U1211 (N_1211,In_68,In_562);
and U1212 (N_1212,In_621,In_589);
xor U1213 (N_1213,In_313,In_577);
or U1214 (N_1214,In_189,In_69);
xnor U1215 (N_1215,In_435,In_53);
or U1216 (N_1216,In_317,In_152);
and U1217 (N_1217,In_221,In_298);
and U1218 (N_1218,In_732,In_22);
nor U1219 (N_1219,In_487,In_297);
nand U1220 (N_1220,In_613,In_257);
nand U1221 (N_1221,In_75,In_694);
or U1222 (N_1222,In_72,In_146);
nand U1223 (N_1223,In_16,In_43);
nand U1224 (N_1224,In_1,In_198);
and U1225 (N_1225,In_122,In_663);
nand U1226 (N_1226,In_119,In_347);
or U1227 (N_1227,In_147,In_5);
nand U1228 (N_1228,In_392,In_150);
nor U1229 (N_1229,In_118,In_429);
nor U1230 (N_1230,In_75,In_515);
or U1231 (N_1231,In_485,In_135);
and U1232 (N_1232,In_513,In_309);
or U1233 (N_1233,In_171,In_366);
or U1234 (N_1234,In_437,In_472);
or U1235 (N_1235,In_197,In_704);
and U1236 (N_1236,In_565,In_429);
or U1237 (N_1237,In_116,In_70);
nand U1238 (N_1238,In_643,In_563);
or U1239 (N_1239,In_568,In_329);
or U1240 (N_1240,In_54,In_150);
nand U1241 (N_1241,In_428,In_128);
xnor U1242 (N_1242,In_719,In_730);
nand U1243 (N_1243,In_604,In_380);
nor U1244 (N_1244,In_687,In_93);
xor U1245 (N_1245,In_698,In_685);
and U1246 (N_1246,In_674,In_598);
nor U1247 (N_1247,In_0,In_74);
or U1248 (N_1248,In_727,In_612);
nor U1249 (N_1249,In_677,In_140);
or U1250 (N_1250,In_241,In_708);
and U1251 (N_1251,In_557,In_519);
nand U1252 (N_1252,In_366,In_677);
or U1253 (N_1253,In_639,In_589);
nor U1254 (N_1254,In_85,In_52);
nor U1255 (N_1255,In_483,In_340);
nand U1256 (N_1256,In_722,In_625);
nand U1257 (N_1257,In_748,In_57);
nor U1258 (N_1258,In_88,In_454);
xor U1259 (N_1259,In_457,In_727);
xnor U1260 (N_1260,In_424,In_369);
xor U1261 (N_1261,In_13,In_547);
and U1262 (N_1262,In_744,In_528);
or U1263 (N_1263,In_652,In_116);
nand U1264 (N_1264,In_7,In_70);
xnor U1265 (N_1265,In_743,In_498);
or U1266 (N_1266,In_32,In_740);
and U1267 (N_1267,In_502,In_54);
and U1268 (N_1268,In_667,In_62);
nand U1269 (N_1269,In_742,In_216);
and U1270 (N_1270,In_486,In_127);
nand U1271 (N_1271,In_538,In_557);
nand U1272 (N_1272,In_541,In_428);
nand U1273 (N_1273,In_692,In_389);
nand U1274 (N_1274,In_442,In_175);
nor U1275 (N_1275,In_501,In_100);
nand U1276 (N_1276,In_432,In_270);
and U1277 (N_1277,In_257,In_116);
xnor U1278 (N_1278,In_601,In_557);
nand U1279 (N_1279,In_741,In_245);
and U1280 (N_1280,In_194,In_351);
nor U1281 (N_1281,In_617,In_640);
nand U1282 (N_1282,In_215,In_460);
and U1283 (N_1283,In_659,In_19);
or U1284 (N_1284,In_129,In_729);
nor U1285 (N_1285,In_137,In_396);
xnor U1286 (N_1286,In_17,In_383);
nor U1287 (N_1287,In_415,In_336);
xor U1288 (N_1288,In_500,In_248);
and U1289 (N_1289,In_390,In_22);
nand U1290 (N_1290,In_135,In_449);
nand U1291 (N_1291,In_670,In_435);
nand U1292 (N_1292,In_523,In_593);
and U1293 (N_1293,In_677,In_131);
nor U1294 (N_1294,In_723,In_430);
xnor U1295 (N_1295,In_566,In_455);
nor U1296 (N_1296,In_255,In_85);
nor U1297 (N_1297,In_330,In_276);
nor U1298 (N_1298,In_725,In_367);
nand U1299 (N_1299,In_197,In_615);
nor U1300 (N_1300,In_40,In_121);
nor U1301 (N_1301,In_629,In_448);
or U1302 (N_1302,In_696,In_711);
or U1303 (N_1303,In_211,In_129);
or U1304 (N_1304,In_65,In_119);
or U1305 (N_1305,In_385,In_509);
and U1306 (N_1306,In_580,In_269);
xor U1307 (N_1307,In_243,In_313);
or U1308 (N_1308,In_616,In_372);
xnor U1309 (N_1309,In_212,In_485);
and U1310 (N_1310,In_123,In_188);
or U1311 (N_1311,In_715,In_556);
nand U1312 (N_1312,In_252,In_579);
and U1313 (N_1313,In_568,In_425);
or U1314 (N_1314,In_535,In_476);
nand U1315 (N_1315,In_302,In_2);
nor U1316 (N_1316,In_528,In_83);
nand U1317 (N_1317,In_742,In_170);
nand U1318 (N_1318,In_118,In_640);
nor U1319 (N_1319,In_112,In_301);
or U1320 (N_1320,In_594,In_739);
and U1321 (N_1321,In_308,In_170);
or U1322 (N_1322,In_167,In_218);
or U1323 (N_1323,In_521,In_680);
or U1324 (N_1324,In_269,In_5);
xor U1325 (N_1325,In_699,In_380);
xnor U1326 (N_1326,In_540,In_253);
and U1327 (N_1327,In_519,In_256);
nand U1328 (N_1328,In_125,In_574);
nor U1329 (N_1329,In_147,In_606);
or U1330 (N_1330,In_552,In_9);
or U1331 (N_1331,In_369,In_598);
xor U1332 (N_1332,In_287,In_540);
nand U1333 (N_1333,In_19,In_693);
or U1334 (N_1334,In_626,In_284);
nand U1335 (N_1335,In_15,In_578);
and U1336 (N_1336,In_229,In_640);
or U1337 (N_1337,In_430,In_261);
nand U1338 (N_1338,In_712,In_499);
xor U1339 (N_1339,In_242,In_256);
nand U1340 (N_1340,In_536,In_582);
nand U1341 (N_1341,In_592,In_342);
nor U1342 (N_1342,In_239,In_443);
nand U1343 (N_1343,In_530,In_83);
nor U1344 (N_1344,In_521,In_232);
or U1345 (N_1345,In_560,In_613);
or U1346 (N_1346,In_78,In_580);
or U1347 (N_1347,In_472,In_285);
and U1348 (N_1348,In_426,In_421);
xor U1349 (N_1349,In_195,In_76);
nor U1350 (N_1350,In_260,In_411);
nand U1351 (N_1351,In_433,In_19);
and U1352 (N_1352,In_516,In_596);
xnor U1353 (N_1353,In_32,In_303);
and U1354 (N_1354,In_90,In_334);
or U1355 (N_1355,In_8,In_643);
and U1356 (N_1356,In_736,In_145);
or U1357 (N_1357,In_727,In_182);
or U1358 (N_1358,In_426,In_463);
nor U1359 (N_1359,In_318,In_2);
nor U1360 (N_1360,In_578,In_188);
or U1361 (N_1361,In_328,In_135);
and U1362 (N_1362,In_242,In_652);
and U1363 (N_1363,In_505,In_334);
xor U1364 (N_1364,In_479,In_116);
xor U1365 (N_1365,In_672,In_300);
and U1366 (N_1366,In_33,In_0);
or U1367 (N_1367,In_176,In_174);
and U1368 (N_1368,In_226,In_373);
or U1369 (N_1369,In_143,In_329);
or U1370 (N_1370,In_346,In_185);
nand U1371 (N_1371,In_603,In_744);
or U1372 (N_1372,In_448,In_51);
or U1373 (N_1373,In_407,In_285);
nor U1374 (N_1374,In_323,In_359);
and U1375 (N_1375,In_736,In_154);
nand U1376 (N_1376,In_329,In_361);
nor U1377 (N_1377,In_330,In_374);
or U1378 (N_1378,In_368,In_317);
and U1379 (N_1379,In_705,In_424);
or U1380 (N_1380,In_129,In_715);
or U1381 (N_1381,In_123,In_86);
and U1382 (N_1382,In_333,In_387);
and U1383 (N_1383,In_709,In_75);
nor U1384 (N_1384,In_97,In_651);
and U1385 (N_1385,In_127,In_339);
xnor U1386 (N_1386,In_11,In_282);
xnor U1387 (N_1387,In_84,In_540);
nand U1388 (N_1388,In_368,In_542);
or U1389 (N_1389,In_95,In_51);
or U1390 (N_1390,In_34,In_377);
and U1391 (N_1391,In_551,In_11);
nand U1392 (N_1392,In_93,In_168);
or U1393 (N_1393,In_227,In_74);
nor U1394 (N_1394,In_269,In_314);
nor U1395 (N_1395,In_380,In_629);
nand U1396 (N_1396,In_194,In_137);
and U1397 (N_1397,In_456,In_439);
and U1398 (N_1398,In_524,In_653);
nand U1399 (N_1399,In_429,In_400);
or U1400 (N_1400,In_188,In_655);
and U1401 (N_1401,In_58,In_230);
or U1402 (N_1402,In_203,In_561);
nand U1403 (N_1403,In_112,In_190);
nor U1404 (N_1404,In_200,In_668);
nand U1405 (N_1405,In_137,In_481);
xnor U1406 (N_1406,In_119,In_0);
and U1407 (N_1407,In_171,In_512);
or U1408 (N_1408,In_267,In_90);
nor U1409 (N_1409,In_478,In_18);
or U1410 (N_1410,In_172,In_358);
nor U1411 (N_1411,In_434,In_592);
xnor U1412 (N_1412,In_83,In_232);
nand U1413 (N_1413,In_252,In_669);
or U1414 (N_1414,In_625,In_473);
nor U1415 (N_1415,In_405,In_63);
nand U1416 (N_1416,In_375,In_211);
xor U1417 (N_1417,In_283,In_540);
nor U1418 (N_1418,In_139,In_482);
nor U1419 (N_1419,In_659,In_361);
nand U1420 (N_1420,In_522,In_345);
or U1421 (N_1421,In_114,In_628);
nand U1422 (N_1422,In_237,In_302);
nor U1423 (N_1423,In_334,In_655);
nor U1424 (N_1424,In_80,In_313);
and U1425 (N_1425,In_358,In_305);
and U1426 (N_1426,In_288,In_238);
nand U1427 (N_1427,In_736,In_167);
nand U1428 (N_1428,In_429,In_421);
nand U1429 (N_1429,In_107,In_669);
nor U1430 (N_1430,In_382,In_301);
and U1431 (N_1431,In_23,In_650);
or U1432 (N_1432,In_211,In_577);
or U1433 (N_1433,In_160,In_569);
and U1434 (N_1434,In_331,In_712);
or U1435 (N_1435,In_516,In_602);
and U1436 (N_1436,In_150,In_318);
or U1437 (N_1437,In_456,In_133);
xor U1438 (N_1438,In_629,In_14);
nand U1439 (N_1439,In_353,In_258);
nand U1440 (N_1440,In_84,In_315);
nand U1441 (N_1441,In_49,In_731);
nor U1442 (N_1442,In_256,In_87);
or U1443 (N_1443,In_257,In_406);
and U1444 (N_1444,In_320,In_333);
or U1445 (N_1445,In_392,In_399);
and U1446 (N_1446,In_134,In_234);
nor U1447 (N_1447,In_643,In_321);
or U1448 (N_1448,In_124,In_477);
xor U1449 (N_1449,In_471,In_175);
xnor U1450 (N_1450,In_5,In_443);
or U1451 (N_1451,In_338,In_154);
nor U1452 (N_1452,In_675,In_696);
nor U1453 (N_1453,In_670,In_223);
and U1454 (N_1454,In_284,In_633);
nand U1455 (N_1455,In_663,In_746);
nor U1456 (N_1456,In_701,In_81);
nand U1457 (N_1457,In_332,In_322);
or U1458 (N_1458,In_549,In_135);
nor U1459 (N_1459,In_467,In_241);
nand U1460 (N_1460,In_689,In_738);
nor U1461 (N_1461,In_167,In_119);
or U1462 (N_1462,In_177,In_135);
nor U1463 (N_1463,In_386,In_1);
nand U1464 (N_1464,In_490,In_423);
or U1465 (N_1465,In_255,In_385);
xnor U1466 (N_1466,In_681,In_620);
xor U1467 (N_1467,In_533,In_238);
nand U1468 (N_1468,In_186,In_130);
nand U1469 (N_1469,In_538,In_687);
or U1470 (N_1470,In_639,In_136);
nor U1471 (N_1471,In_183,In_185);
or U1472 (N_1472,In_421,In_251);
xor U1473 (N_1473,In_453,In_288);
and U1474 (N_1474,In_570,In_34);
and U1475 (N_1475,In_258,In_51);
or U1476 (N_1476,In_729,In_409);
nor U1477 (N_1477,In_577,In_225);
nor U1478 (N_1478,In_255,In_90);
and U1479 (N_1479,In_368,In_455);
nand U1480 (N_1480,In_141,In_444);
or U1481 (N_1481,In_169,In_476);
nand U1482 (N_1482,In_319,In_408);
or U1483 (N_1483,In_193,In_7);
and U1484 (N_1484,In_130,In_609);
and U1485 (N_1485,In_431,In_684);
xnor U1486 (N_1486,In_419,In_469);
nor U1487 (N_1487,In_196,In_237);
and U1488 (N_1488,In_175,In_641);
nand U1489 (N_1489,In_296,In_361);
nand U1490 (N_1490,In_135,In_420);
and U1491 (N_1491,In_6,In_300);
or U1492 (N_1492,In_204,In_6);
xor U1493 (N_1493,In_144,In_483);
xnor U1494 (N_1494,In_426,In_461);
or U1495 (N_1495,In_482,In_358);
and U1496 (N_1496,In_391,In_667);
nor U1497 (N_1497,In_426,In_86);
nand U1498 (N_1498,In_734,In_150);
or U1499 (N_1499,In_469,In_442);
nand U1500 (N_1500,In_20,In_445);
or U1501 (N_1501,In_571,In_327);
nand U1502 (N_1502,In_609,In_496);
and U1503 (N_1503,In_8,In_269);
nor U1504 (N_1504,In_173,In_585);
xnor U1505 (N_1505,In_92,In_175);
or U1506 (N_1506,In_66,In_324);
or U1507 (N_1507,In_72,In_617);
xnor U1508 (N_1508,In_584,In_321);
or U1509 (N_1509,In_125,In_21);
or U1510 (N_1510,In_277,In_236);
and U1511 (N_1511,In_694,In_198);
nand U1512 (N_1512,In_675,In_490);
nor U1513 (N_1513,In_300,In_648);
nand U1514 (N_1514,In_289,In_706);
or U1515 (N_1515,In_34,In_461);
and U1516 (N_1516,In_51,In_399);
nor U1517 (N_1517,In_391,In_220);
or U1518 (N_1518,In_103,In_486);
and U1519 (N_1519,In_77,In_677);
nor U1520 (N_1520,In_403,In_560);
and U1521 (N_1521,In_551,In_272);
and U1522 (N_1522,In_384,In_601);
or U1523 (N_1523,In_680,In_684);
nor U1524 (N_1524,In_328,In_445);
or U1525 (N_1525,In_310,In_698);
or U1526 (N_1526,In_690,In_629);
nor U1527 (N_1527,In_403,In_490);
and U1528 (N_1528,In_697,In_409);
xnor U1529 (N_1529,In_437,In_74);
nor U1530 (N_1530,In_690,In_251);
nor U1531 (N_1531,In_265,In_246);
nand U1532 (N_1532,In_14,In_86);
nand U1533 (N_1533,In_32,In_416);
and U1534 (N_1534,In_275,In_520);
or U1535 (N_1535,In_155,In_164);
and U1536 (N_1536,In_690,In_152);
xor U1537 (N_1537,In_715,In_158);
or U1538 (N_1538,In_311,In_549);
nor U1539 (N_1539,In_441,In_361);
nand U1540 (N_1540,In_539,In_593);
nand U1541 (N_1541,In_374,In_712);
or U1542 (N_1542,In_528,In_124);
and U1543 (N_1543,In_52,In_268);
xor U1544 (N_1544,In_113,In_462);
nand U1545 (N_1545,In_712,In_579);
nor U1546 (N_1546,In_633,In_456);
and U1547 (N_1547,In_375,In_480);
or U1548 (N_1548,In_36,In_535);
or U1549 (N_1549,In_366,In_84);
nor U1550 (N_1550,In_86,In_29);
or U1551 (N_1551,In_465,In_84);
nor U1552 (N_1552,In_160,In_189);
nand U1553 (N_1553,In_238,In_453);
xor U1554 (N_1554,In_493,In_555);
nor U1555 (N_1555,In_693,In_134);
nand U1556 (N_1556,In_738,In_24);
and U1557 (N_1557,In_194,In_612);
or U1558 (N_1558,In_161,In_111);
and U1559 (N_1559,In_689,In_624);
nand U1560 (N_1560,In_423,In_73);
nand U1561 (N_1561,In_641,In_600);
and U1562 (N_1562,In_320,In_636);
nor U1563 (N_1563,In_498,In_463);
and U1564 (N_1564,In_446,In_713);
and U1565 (N_1565,In_52,In_448);
and U1566 (N_1566,In_383,In_13);
and U1567 (N_1567,In_160,In_130);
nor U1568 (N_1568,In_399,In_225);
nand U1569 (N_1569,In_236,In_532);
and U1570 (N_1570,In_624,In_382);
and U1571 (N_1571,In_102,In_72);
or U1572 (N_1572,In_277,In_491);
nand U1573 (N_1573,In_8,In_371);
nor U1574 (N_1574,In_620,In_528);
and U1575 (N_1575,In_740,In_733);
nor U1576 (N_1576,In_388,In_441);
nor U1577 (N_1577,In_284,In_80);
xnor U1578 (N_1578,In_602,In_733);
and U1579 (N_1579,In_450,In_327);
and U1580 (N_1580,In_18,In_637);
nor U1581 (N_1581,In_22,In_180);
or U1582 (N_1582,In_398,In_461);
nor U1583 (N_1583,In_413,In_689);
nor U1584 (N_1584,In_155,In_59);
nor U1585 (N_1585,In_385,In_200);
nor U1586 (N_1586,In_83,In_169);
nand U1587 (N_1587,In_505,In_408);
nor U1588 (N_1588,In_34,In_395);
xor U1589 (N_1589,In_63,In_342);
and U1590 (N_1590,In_420,In_13);
nand U1591 (N_1591,In_176,In_689);
nand U1592 (N_1592,In_74,In_669);
or U1593 (N_1593,In_467,In_199);
nor U1594 (N_1594,In_691,In_734);
or U1595 (N_1595,In_212,In_340);
or U1596 (N_1596,In_690,In_716);
nand U1597 (N_1597,In_197,In_200);
or U1598 (N_1598,In_262,In_75);
or U1599 (N_1599,In_433,In_224);
or U1600 (N_1600,In_578,In_249);
xnor U1601 (N_1601,In_609,In_391);
or U1602 (N_1602,In_267,In_433);
nand U1603 (N_1603,In_334,In_627);
nor U1604 (N_1604,In_202,In_514);
or U1605 (N_1605,In_430,In_82);
nand U1606 (N_1606,In_303,In_98);
nor U1607 (N_1607,In_653,In_597);
or U1608 (N_1608,In_357,In_161);
or U1609 (N_1609,In_549,In_185);
or U1610 (N_1610,In_443,In_676);
and U1611 (N_1611,In_393,In_116);
xnor U1612 (N_1612,In_690,In_425);
nand U1613 (N_1613,In_158,In_212);
and U1614 (N_1614,In_432,In_308);
or U1615 (N_1615,In_317,In_707);
or U1616 (N_1616,In_357,In_10);
or U1617 (N_1617,In_669,In_680);
or U1618 (N_1618,In_136,In_721);
xnor U1619 (N_1619,In_394,In_309);
nand U1620 (N_1620,In_108,In_198);
and U1621 (N_1621,In_576,In_239);
nor U1622 (N_1622,In_29,In_68);
nand U1623 (N_1623,In_282,In_741);
xnor U1624 (N_1624,In_493,In_167);
or U1625 (N_1625,In_571,In_153);
nand U1626 (N_1626,In_677,In_525);
nor U1627 (N_1627,In_212,In_198);
nand U1628 (N_1628,In_290,In_531);
or U1629 (N_1629,In_21,In_401);
and U1630 (N_1630,In_574,In_354);
nand U1631 (N_1631,In_635,In_376);
nand U1632 (N_1632,In_550,In_706);
nor U1633 (N_1633,In_165,In_424);
nor U1634 (N_1634,In_100,In_10);
and U1635 (N_1635,In_116,In_704);
nand U1636 (N_1636,In_749,In_717);
nor U1637 (N_1637,In_649,In_106);
and U1638 (N_1638,In_554,In_674);
and U1639 (N_1639,In_292,In_198);
or U1640 (N_1640,In_224,In_172);
nor U1641 (N_1641,In_54,In_197);
nand U1642 (N_1642,In_28,In_645);
nand U1643 (N_1643,In_557,In_715);
nand U1644 (N_1644,In_65,In_344);
or U1645 (N_1645,In_72,In_327);
nand U1646 (N_1646,In_257,In_170);
nor U1647 (N_1647,In_286,In_402);
nand U1648 (N_1648,In_111,In_652);
xor U1649 (N_1649,In_421,In_147);
and U1650 (N_1650,In_175,In_270);
nor U1651 (N_1651,In_247,In_193);
nor U1652 (N_1652,In_361,In_62);
and U1653 (N_1653,In_348,In_748);
nand U1654 (N_1654,In_58,In_585);
nand U1655 (N_1655,In_598,In_27);
and U1656 (N_1656,In_258,In_150);
and U1657 (N_1657,In_413,In_676);
nor U1658 (N_1658,In_498,In_358);
or U1659 (N_1659,In_75,In_645);
nand U1660 (N_1660,In_350,In_475);
xnor U1661 (N_1661,In_260,In_587);
and U1662 (N_1662,In_239,In_744);
nor U1663 (N_1663,In_104,In_687);
and U1664 (N_1664,In_441,In_516);
or U1665 (N_1665,In_697,In_603);
and U1666 (N_1666,In_350,In_357);
and U1667 (N_1667,In_233,In_335);
xor U1668 (N_1668,In_613,In_192);
nand U1669 (N_1669,In_430,In_558);
nor U1670 (N_1670,In_620,In_183);
nand U1671 (N_1671,In_245,In_61);
nor U1672 (N_1672,In_655,In_488);
and U1673 (N_1673,In_261,In_633);
and U1674 (N_1674,In_469,In_711);
nand U1675 (N_1675,In_415,In_198);
and U1676 (N_1676,In_242,In_714);
nor U1677 (N_1677,In_507,In_406);
nand U1678 (N_1678,In_265,In_659);
or U1679 (N_1679,In_336,In_95);
or U1680 (N_1680,In_127,In_309);
nand U1681 (N_1681,In_93,In_139);
or U1682 (N_1682,In_7,In_110);
and U1683 (N_1683,In_610,In_32);
or U1684 (N_1684,In_696,In_590);
or U1685 (N_1685,In_316,In_354);
and U1686 (N_1686,In_543,In_743);
nand U1687 (N_1687,In_218,In_249);
or U1688 (N_1688,In_710,In_44);
or U1689 (N_1689,In_464,In_508);
or U1690 (N_1690,In_629,In_455);
nor U1691 (N_1691,In_455,In_405);
nand U1692 (N_1692,In_519,In_517);
nor U1693 (N_1693,In_303,In_455);
and U1694 (N_1694,In_171,In_453);
nand U1695 (N_1695,In_276,In_524);
and U1696 (N_1696,In_546,In_132);
or U1697 (N_1697,In_595,In_323);
or U1698 (N_1698,In_304,In_613);
nand U1699 (N_1699,In_31,In_582);
xnor U1700 (N_1700,In_158,In_514);
and U1701 (N_1701,In_46,In_117);
nor U1702 (N_1702,In_264,In_160);
or U1703 (N_1703,In_650,In_172);
and U1704 (N_1704,In_435,In_748);
nand U1705 (N_1705,In_374,In_39);
nor U1706 (N_1706,In_160,In_379);
or U1707 (N_1707,In_302,In_599);
or U1708 (N_1708,In_653,In_677);
nor U1709 (N_1709,In_578,In_324);
or U1710 (N_1710,In_71,In_679);
xor U1711 (N_1711,In_380,In_630);
nor U1712 (N_1712,In_416,In_71);
nor U1713 (N_1713,In_365,In_484);
or U1714 (N_1714,In_18,In_524);
nand U1715 (N_1715,In_665,In_105);
or U1716 (N_1716,In_189,In_165);
nand U1717 (N_1717,In_733,In_495);
and U1718 (N_1718,In_424,In_537);
nand U1719 (N_1719,In_61,In_222);
nand U1720 (N_1720,In_68,In_556);
nor U1721 (N_1721,In_48,In_600);
or U1722 (N_1722,In_373,In_430);
or U1723 (N_1723,In_332,In_745);
nor U1724 (N_1724,In_356,In_233);
or U1725 (N_1725,In_402,In_152);
xnor U1726 (N_1726,In_748,In_133);
nor U1727 (N_1727,In_188,In_545);
nor U1728 (N_1728,In_744,In_573);
nand U1729 (N_1729,In_174,In_668);
nor U1730 (N_1730,In_210,In_195);
nand U1731 (N_1731,In_257,In_173);
nor U1732 (N_1732,In_236,In_261);
and U1733 (N_1733,In_572,In_680);
or U1734 (N_1734,In_54,In_195);
nor U1735 (N_1735,In_132,In_72);
or U1736 (N_1736,In_225,In_528);
and U1737 (N_1737,In_718,In_454);
or U1738 (N_1738,In_270,In_650);
and U1739 (N_1739,In_14,In_280);
nor U1740 (N_1740,In_150,In_358);
nand U1741 (N_1741,In_21,In_93);
or U1742 (N_1742,In_384,In_435);
xnor U1743 (N_1743,In_701,In_468);
and U1744 (N_1744,In_114,In_6);
nand U1745 (N_1745,In_82,In_699);
xor U1746 (N_1746,In_109,In_206);
and U1747 (N_1747,In_554,In_143);
or U1748 (N_1748,In_320,In_108);
nand U1749 (N_1749,In_667,In_658);
nand U1750 (N_1750,In_742,In_286);
and U1751 (N_1751,In_404,In_667);
xor U1752 (N_1752,In_456,In_661);
nor U1753 (N_1753,In_367,In_252);
nand U1754 (N_1754,In_135,In_188);
or U1755 (N_1755,In_70,In_598);
xor U1756 (N_1756,In_407,In_641);
or U1757 (N_1757,In_342,In_411);
and U1758 (N_1758,In_514,In_472);
nor U1759 (N_1759,In_355,In_712);
and U1760 (N_1760,In_233,In_371);
and U1761 (N_1761,In_81,In_715);
nand U1762 (N_1762,In_616,In_17);
nand U1763 (N_1763,In_690,In_538);
xor U1764 (N_1764,In_657,In_186);
and U1765 (N_1765,In_577,In_164);
and U1766 (N_1766,In_260,In_658);
or U1767 (N_1767,In_718,In_544);
or U1768 (N_1768,In_701,In_737);
nor U1769 (N_1769,In_492,In_505);
nor U1770 (N_1770,In_598,In_288);
and U1771 (N_1771,In_227,In_572);
xor U1772 (N_1772,In_157,In_430);
xor U1773 (N_1773,In_528,In_448);
and U1774 (N_1774,In_610,In_92);
or U1775 (N_1775,In_749,In_291);
and U1776 (N_1776,In_194,In_253);
and U1777 (N_1777,In_164,In_692);
nor U1778 (N_1778,In_20,In_601);
and U1779 (N_1779,In_341,In_292);
nand U1780 (N_1780,In_277,In_151);
or U1781 (N_1781,In_297,In_70);
nand U1782 (N_1782,In_460,In_249);
and U1783 (N_1783,In_549,In_373);
or U1784 (N_1784,In_606,In_132);
nor U1785 (N_1785,In_635,In_645);
and U1786 (N_1786,In_389,In_476);
nand U1787 (N_1787,In_702,In_620);
nand U1788 (N_1788,In_214,In_534);
nor U1789 (N_1789,In_338,In_477);
and U1790 (N_1790,In_355,In_498);
and U1791 (N_1791,In_708,In_342);
xnor U1792 (N_1792,In_413,In_361);
xor U1793 (N_1793,In_16,In_456);
nor U1794 (N_1794,In_258,In_309);
or U1795 (N_1795,In_378,In_458);
or U1796 (N_1796,In_507,In_194);
nor U1797 (N_1797,In_435,In_244);
nor U1798 (N_1798,In_687,In_657);
xnor U1799 (N_1799,In_626,In_87);
nand U1800 (N_1800,In_699,In_179);
and U1801 (N_1801,In_353,In_704);
nor U1802 (N_1802,In_460,In_704);
nand U1803 (N_1803,In_660,In_412);
and U1804 (N_1804,In_196,In_253);
or U1805 (N_1805,In_375,In_56);
nor U1806 (N_1806,In_137,In_374);
or U1807 (N_1807,In_521,In_33);
nand U1808 (N_1808,In_658,In_9);
nor U1809 (N_1809,In_396,In_642);
nor U1810 (N_1810,In_309,In_241);
nor U1811 (N_1811,In_148,In_17);
xnor U1812 (N_1812,In_351,In_70);
and U1813 (N_1813,In_190,In_27);
nand U1814 (N_1814,In_661,In_235);
and U1815 (N_1815,In_690,In_660);
xor U1816 (N_1816,In_257,In_66);
and U1817 (N_1817,In_293,In_356);
xnor U1818 (N_1818,In_690,In_151);
nor U1819 (N_1819,In_611,In_189);
nor U1820 (N_1820,In_532,In_201);
nor U1821 (N_1821,In_598,In_591);
and U1822 (N_1822,In_13,In_136);
or U1823 (N_1823,In_8,In_534);
nand U1824 (N_1824,In_683,In_90);
nand U1825 (N_1825,In_730,In_223);
or U1826 (N_1826,In_457,In_612);
nand U1827 (N_1827,In_391,In_566);
and U1828 (N_1828,In_722,In_155);
and U1829 (N_1829,In_379,In_184);
nand U1830 (N_1830,In_556,In_562);
nor U1831 (N_1831,In_345,In_479);
nor U1832 (N_1832,In_232,In_425);
nand U1833 (N_1833,In_196,In_88);
nand U1834 (N_1834,In_712,In_59);
nor U1835 (N_1835,In_397,In_540);
or U1836 (N_1836,In_452,In_743);
or U1837 (N_1837,In_408,In_309);
and U1838 (N_1838,In_250,In_571);
and U1839 (N_1839,In_306,In_426);
and U1840 (N_1840,In_521,In_573);
or U1841 (N_1841,In_402,In_46);
or U1842 (N_1842,In_213,In_359);
nand U1843 (N_1843,In_585,In_620);
or U1844 (N_1844,In_560,In_397);
and U1845 (N_1845,In_73,In_610);
or U1846 (N_1846,In_88,In_695);
nor U1847 (N_1847,In_612,In_103);
or U1848 (N_1848,In_693,In_292);
nor U1849 (N_1849,In_352,In_376);
or U1850 (N_1850,In_619,In_557);
and U1851 (N_1851,In_192,In_357);
nand U1852 (N_1852,In_393,In_65);
nor U1853 (N_1853,In_0,In_520);
nand U1854 (N_1854,In_603,In_687);
or U1855 (N_1855,In_394,In_642);
or U1856 (N_1856,In_651,In_567);
or U1857 (N_1857,In_311,In_371);
or U1858 (N_1858,In_272,In_702);
nor U1859 (N_1859,In_93,In_238);
and U1860 (N_1860,In_3,In_651);
and U1861 (N_1861,In_354,In_341);
nor U1862 (N_1862,In_218,In_340);
nand U1863 (N_1863,In_661,In_379);
nand U1864 (N_1864,In_732,In_646);
or U1865 (N_1865,In_106,In_153);
nand U1866 (N_1866,In_458,In_283);
xor U1867 (N_1867,In_76,In_126);
or U1868 (N_1868,In_44,In_254);
nand U1869 (N_1869,In_7,In_626);
xor U1870 (N_1870,In_729,In_173);
and U1871 (N_1871,In_411,In_355);
and U1872 (N_1872,In_279,In_375);
nand U1873 (N_1873,In_394,In_564);
and U1874 (N_1874,In_260,In_718);
or U1875 (N_1875,In_366,In_209);
and U1876 (N_1876,In_728,In_0);
and U1877 (N_1877,In_246,In_259);
nand U1878 (N_1878,In_365,In_606);
nand U1879 (N_1879,In_510,In_95);
xnor U1880 (N_1880,In_42,In_300);
or U1881 (N_1881,In_394,In_739);
nand U1882 (N_1882,In_351,In_469);
or U1883 (N_1883,In_572,In_384);
and U1884 (N_1884,In_265,In_69);
nor U1885 (N_1885,In_531,In_646);
or U1886 (N_1886,In_547,In_561);
nand U1887 (N_1887,In_694,In_266);
or U1888 (N_1888,In_52,In_513);
and U1889 (N_1889,In_684,In_430);
nand U1890 (N_1890,In_490,In_217);
nand U1891 (N_1891,In_581,In_240);
nor U1892 (N_1892,In_228,In_85);
nand U1893 (N_1893,In_636,In_402);
xnor U1894 (N_1894,In_220,In_202);
and U1895 (N_1895,In_186,In_687);
nor U1896 (N_1896,In_368,In_387);
and U1897 (N_1897,In_393,In_385);
and U1898 (N_1898,In_670,In_93);
or U1899 (N_1899,In_48,In_192);
or U1900 (N_1900,In_300,In_10);
and U1901 (N_1901,In_547,In_253);
nand U1902 (N_1902,In_562,In_366);
or U1903 (N_1903,In_451,In_407);
nor U1904 (N_1904,In_665,In_748);
or U1905 (N_1905,In_85,In_637);
nand U1906 (N_1906,In_116,In_508);
and U1907 (N_1907,In_366,In_573);
or U1908 (N_1908,In_366,In_290);
xnor U1909 (N_1909,In_682,In_542);
or U1910 (N_1910,In_709,In_683);
or U1911 (N_1911,In_622,In_549);
nor U1912 (N_1912,In_159,In_206);
or U1913 (N_1913,In_167,In_685);
or U1914 (N_1914,In_458,In_410);
and U1915 (N_1915,In_45,In_411);
and U1916 (N_1916,In_236,In_4);
nand U1917 (N_1917,In_713,In_650);
nand U1918 (N_1918,In_717,In_152);
or U1919 (N_1919,In_649,In_4);
and U1920 (N_1920,In_37,In_173);
nand U1921 (N_1921,In_44,In_472);
nand U1922 (N_1922,In_397,In_107);
xor U1923 (N_1923,In_48,In_166);
nand U1924 (N_1924,In_324,In_85);
or U1925 (N_1925,In_630,In_412);
nor U1926 (N_1926,In_444,In_126);
and U1927 (N_1927,In_264,In_423);
nor U1928 (N_1928,In_723,In_233);
and U1929 (N_1929,In_559,In_223);
xor U1930 (N_1930,In_520,In_144);
nor U1931 (N_1931,In_631,In_344);
xor U1932 (N_1932,In_285,In_225);
or U1933 (N_1933,In_95,In_132);
nand U1934 (N_1934,In_227,In_168);
xnor U1935 (N_1935,In_116,In_370);
or U1936 (N_1936,In_56,In_242);
and U1937 (N_1937,In_105,In_206);
and U1938 (N_1938,In_286,In_76);
nand U1939 (N_1939,In_147,In_188);
nand U1940 (N_1940,In_178,In_693);
nor U1941 (N_1941,In_20,In_14);
and U1942 (N_1942,In_23,In_153);
xnor U1943 (N_1943,In_46,In_110);
xnor U1944 (N_1944,In_95,In_485);
and U1945 (N_1945,In_583,In_261);
or U1946 (N_1946,In_391,In_285);
and U1947 (N_1947,In_531,In_497);
and U1948 (N_1948,In_615,In_723);
or U1949 (N_1949,In_251,In_143);
and U1950 (N_1950,In_222,In_551);
and U1951 (N_1951,In_568,In_527);
and U1952 (N_1952,In_33,In_326);
and U1953 (N_1953,In_534,In_433);
and U1954 (N_1954,In_148,In_502);
nor U1955 (N_1955,In_61,In_462);
and U1956 (N_1956,In_261,In_559);
and U1957 (N_1957,In_485,In_436);
nor U1958 (N_1958,In_134,In_435);
or U1959 (N_1959,In_372,In_337);
xnor U1960 (N_1960,In_10,In_692);
nor U1961 (N_1961,In_732,In_541);
and U1962 (N_1962,In_478,In_250);
nor U1963 (N_1963,In_103,In_455);
and U1964 (N_1964,In_702,In_188);
or U1965 (N_1965,In_459,In_700);
nor U1966 (N_1966,In_527,In_677);
and U1967 (N_1967,In_427,In_481);
or U1968 (N_1968,In_426,In_456);
and U1969 (N_1969,In_458,In_575);
nor U1970 (N_1970,In_359,In_311);
xor U1971 (N_1971,In_56,In_426);
and U1972 (N_1972,In_376,In_300);
and U1973 (N_1973,In_697,In_6);
and U1974 (N_1974,In_424,In_223);
or U1975 (N_1975,In_8,In_638);
nand U1976 (N_1976,In_475,In_544);
or U1977 (N_1977,In_500,In_362);
nor U1978 (N_1978,In_625,In_28);
xor U1979 (N_1979,In_545,In_462);
nand U1980 (N_1980,In_642,In_636);
nor U1981 (N_1981,In_513,In_286);
nor U1982 (N_1982,In_575,In_262);
nor U1983 (N_1983,In_17,In_161);
nor U1984 (N_1984,In_519,In_615);
nand U1985 (N_1985,In_602,In_166);
nand U1986 (N_1986,In_320,In_488);
nor U1987 (N_1987,In_134,In_623);
and U1988 (N_1988,In_665,In_641);
or U1989 (N_1989,In_545,In_426);
and U1990 (N_1990,In_579,In_192);
and U1991 (N_1991,In_2,In_16);
or U1992 (N_1992,In_573,In_44);
and U1993 (N_1993,In_258,In_646);
or U1994 (N_1994,In_157,In_722);
or U1995 (N_1995,In_385,In_651);
nor U1996 (N_1996,In_604,In_601);
nand U1997 (N_1997,In_69,In_642);
or U1998 (N_1998,In_475,In_512);
xor U1999 (N_1999,In_85,In_459);
or U2000 (N_2000,In_404,In_658);
or U2001 (N_2001,In_222,In_48);
or U2002 (N_2002,In_497,In_108);
nand U2003 (N_2003,In_549,In_228);
or U2004 (N_2004,In_327,In_577);
nand U2005 (N_2005,In_159,In_52);
nor U2006 (N_2006,In_569,In_407);
nor U2007 (N_2007,In_413,In_169);
nor U2008 (N_2008,In_444,In_692);
or U2009 (N_2009,In_548,In_399);
and U2010 (N_2010,In_724,In_27);
xnor U2011 (N_2011,In_367,In_625);
or U2012 (N_2012,In_662,In_625);
nand U2013 (N_2013,In_102,In_300);
nor U2014 (N_2014,In_446,In_449);
xnor U2015 (N_2015,In_359,In_227);
nand U2016 (N_2016,In_58,In_410);
nor U2017 (N_2017,In_475,In_482);
and U2018 (N_2018,In_540,In_678);
nand U2019 (N_2019,In_37,In_251);
or U2020 (N_2020,In_296,In_273);
nor U2021 (N_2021,In_81,In_10);
and U2022 (N_2022,In_328,In_691);
and U2023 (N_2023,In_421,In_351);
xor U2024 (N_2024,In_218,In_296);
nand U2025 (N_2025,In_277,In_211);
and U2026 (N_2026,In_479,In_87);
and U2027 (N_2027,In_566,In_246);
nand U2028 (N_2028,In_567,In_643);
xnor U2029 (N_2029,In_350,In_429);
nor U2030 (N_2030,In_350,In_45);
nor U2031 (N_2031,In_561,In_660);
and U2032 (N_2032,In_414,In_509);
and U2033 (N_2033,In_562,In_600);
nand U2034 (N_2034,In_668,In_649);
or U2035 (N_2035,In_406,In_262);
and U2036 (N_2036,In_544,In_706);
nand U2037 (N_2037,In_519,In_724);
xnor U2038 (N_2038,In_315,In_730);
and U2039 (N_2039,In_704,In_203);
nand U2040 (N_2040,In_69,In_634);
and U2041 (N_2041,In_531,In_83);
nand U2042 (N_2042,In_31,In_672);
nand U2043 (N_2043,In_496,In_305);
and U2044 (N_2044,In_11,In_243);
nand U2045 (N_2045,In_687,In_408);
nand U2046 (N_2046,In_745,In_599);
or U2047 (N_2047,In_564,In_640);
or U2048 (N_2048,In_301,In_251);
xor U2049 (N_2049,In_123,In_401);
nor U2050 (N_2050,In_48,In_313);
or U2051 (N_2051,In_220,In_363);
nand U2052 (N_2052,In_274,In_3);
nor U2053 (N_2053,In_448,In_467);
and U2054 (N_2054,In_526,In_519);
nor U2055 (N_2055,In_110,In_538);
or U2056 (N_2056,In_341,In_37);
nor U2057 (N_2057,In_496,In_182);
and U2058 (N_2058,In_50,In_450);
or U2059 (N_2059,In_680,In_594);
nand U2060 (N_2060,In_302,In_31);
nand U2061 (N_2061,In_534,In_684);
nor U2062 (N_2062,In_258,In_459);
xnor U2063 (N_2063,In_508,In_504);
nor U2064 (N_2064,In_40,In_480);
nor U2065 (N_2065,In_122,In_282);
nor U2066 (N_2066,In_638,In_18);
and U2067 (N_2067,In_400,In_482);
or U2068 (N_2068,In_680,In_399);
and U2069 (N_2069,In_700,In_473);
nor U2070 (N_2070,In_157,In_670);
nand U2071 (N_2071,In_96,In_482);
nor U2072 (N_2072,In_425,In_304);
or U2073 (N_2073,In_709,In_72);
nand U2074 (N_2074,In_3,In_158);
or U2075 (N_2075,In_620,In_679);
nor U2076 (N_2076,In_309,In_78);
or U2077 (N_2077,In_206,In_686);
or U2078 (N_2078,In_355,In_713);
or U2079 (N_2079,In_116,In_224);
or U2080 (N_2080,In_299,In_230);
nand U2081 (N_2081,In_558,In_487);
nor U2082 (N_2082,In_508,In_588);
nor U2083 (N_2083,In_168,In_294);
or U2084 (N_2084,In_153,In_298);
nor U2085 (N_2085,In_635,In_32);
and U2086 (N_2086,In_489,In_333);
nand U2087 (N_2087,In_660,In_49);
and U2088 (N_2088,In_81,In_254);
nand U2089 (N_2089,In_8,In_532);
and U2090 (N_2090,In_579,In_155);
and U2091 (N_2091,In_167,In_511);
nor U2092 (N_2092,In_291,In_662);
nor U2093 (N_2093,In_462,In_112);
or U2094 (N_2094,In_748,In_653);
nor U2095 (N_2095,In_490,In_224);
and U2096 (N_2096,In_89,In_627);
or U2097 (N_2097,In_475,In_436);
and U2098 (N_2098,In_480,In_561);
or U2099 (N_2099,In_548,In_114);
and U2100 (N_2100,In_48,In_182);
and U2101 (N_2101,In_65,In_245);
or U2102 (N_2102,In_576,In_449);
and U2103 (N_2103,In_526,In_227);
nor U2104 (N_2104,In_499,In_190);
or U2105 (N_2105,In_155,In_662);
xnor U2106 (N_2106,In_496,In_536);
nand U2107 (N_2107,In_385,In_554);
or U2108 (N_2108,In_523,In_86);
and U2109 (N_2109,In_576,In_631);
or U2110 (N_2110,In_77,In_305);
or U2111 (N_2111,In_597,In_168);
nand U2112 (N_2112,In_152,In_426);
nand U2113 (N_2113,In_737,In_23);
and U2114 (N_2114,In_368,In_596);
xnor U2115 (N_2115,In_727,In_221);
nand U2116 (N_2116,In_57,In_220);
nor U2117 (N_2117,In_747,In_102);
and U2118 (N_2118,In_272,In_332);
and U2119 (N_2119,In_613,In_458);
or U2120 (N_2120,In_510,In_664);
nor U2121 (N_2121,In_384,In_149);
or U2122 (N_2122,In_663,In_27);
and U2123 (N_2123,In_318,In_540);
or U2124 (N_2124,In_28,In_84);
nor U2125 (N_2125,In_216,In_705);
or U2126 (N_2126,In_591,In_354);
and U2127 (N_2127,In_96,In_342);
nor U2128 (N_2128,In_743,In_429);
or U2129 (N_2129,In_396,In_180);
and U2130 (N_2130,In_165,In_244);
nand U2131 (N_2131,In_623,In_352);
or U2132 (N_2132,In_41,In_539);
nand U2133 (N_2133,In_94,In_195);
xor U2134 (N_2134,In_492,In_227);
nor U2135 (N_2135,In_411,In_736);
nor U2136 (N_2136,In_410,In_26);
nand U2137 (N_2137,In_104,In_341);
xor U2138 (N_2138,In_558,In_520);
and U2139 (N_2139,In_83,In_457);
nor U2140 (N_2140,In_415,In_58);
or U2141 (N_2141,In_234,In_647);
and U2142 (N_2142,In_744,In_642);
and U2143 (N_2143,In_707,In_153);
or U2144 (N_2144,In_339,In_640);
nand U2145 (N_2145,In_645,In_93);
xnor U2146 (N_2146,In_147,In_73);
or U2147 (N_2147,In_521,In_293);
and U2148 (N_2148,In_525,In_711);
or U2149 (N_2149,In_202,In_90);
nand U2150 (N_2150,In_33,In_492);
or U2151 (N_2151,In_466,In_269);
nand U2152 (N_2152,In_374,In_513);
and U2153 (N_2153,In_512,In_377);
xnor U2154 (N_2154,In_5,In_532);
or U2155 (N_2155,In_464,In_671);
nand U2156 (N_2156,In_122,In_129);
nor U2157 (N_2157,In_184,In_403);
nor U2158 (N_2158,In_363,In_367);
nor U2159 (N_2159,In_708,In_29);
or U2160 (N_2160,In_327,In_520);
and U2161 (N_2161,In_140,In_697);
or U2162 (N_2162,In_120,In_736);
xnor U2163 (N_2163,In_80,In_100);
or U2164 (N_2164,In_494,In_323);
xor U2165 (N_2165,In_478,In_133);
nor U2166 (N_2166,In_429,In_478);
xnor U2167 (N_2167,In_229,In_708);
and U2168 (N_2168,In_96,In_655);
or U2169 (N_2169,In_39,In_325);
and U2170 (N_2170,In_442,In_749);
nand U2171 (N_2171,In_186,In_286);
and U2172 (N_2172,In_216,In_464);
nor U2173 (N_2173,In_747,In_540);
and U2174 (N_2174,In_331,In_233);
and U2175 (N_2175,In_741,In_270);
nor U2176 (N_2176,In_692,In_40);
nand U2177 (N_2177,In_107,In_704);
nor U2178 (N_2178,In_447,In_739);
xnor U2179 (N_2179,In_469,In_302);
or U2180 (N_2180,In_633,In_571);
nand U2181 (N_2181,In_423,In_393);
or U2182 (N_2182,In_204,In_163);
and U2183 (N_2183,In_484,In_472);
nand U2184 (N_2184,In_239,In_107);
nor U2185 (N_2185,In_408,In_243);
or U2186 (N_2186,In_515,In_111);
nand U2187 (N_2187,In_338,In_597);
nor U2188 (N_2188,In_19,In_556);
nor U2189 (N_2189,In_621,In_20);
nor U2190 (N_2190,In_567,In_52);
or U2191 (N_2191,In_65,In_10);
xor U2192 (N_2192,In_719,In_617);
nor U2193 (N_2193,In_542,In_499);
or U2194 (N_2194,In_51,In_12);
nor U2195 (N_2195,In_626,In_459);
xor U2196 (N_2196,In_339,In_279);
and U2197 (N_2197,In_163,In_704);
nand U2198 (N_2198,In_384,In_702);
nor U2199 (N_2199,In_467,In_558);
nand U2200 (N_2200,In_117,In_85);
nand U2201 (N_2201,In_511,In_520);
or U2202 (N_2202,In_209,In_70);
nor U2203 (N_2203,In_737,In_6);
nor U2204 (N_2204,In_291,In_736);
nor U2205 (N_2205,In_155,In_475);
nor U2206 (N_2206,In_674,In_545);
and U2207 (N_2207,In_298,In_210);
nor U2208 (N_2208,In_644,In_373);
or U2209 (N_2209,In_227,In_717);
and U2210 (N_2210,In_690,In_109);
nor U2211 (N_2211,In_703,In_318);
or U2212 (N_2212,In_313,In_512);
nand U2213 (N_2213,In_95,In_526);
nand U2214 (N_2214,In_209,In_657);
or U2215 (N_2215,In_643,In_400);
nand U2216 (N_2216,In_29,In_127);
and U2217 (N_2217,In_548,In_13);
or U2218 (N_2218,In_503,In_433);
xor U2219 (N_2219,In_729,In_193);
xor U2220 (N_2220,In_584,In_743);
and U2221 (N_2221,In_47,In_153);
or U2222 (N_2222,In_1,In_27);
nand U2223 (N_2223,In_500,In_666);
or U2224 (N_2224,In_338,In_423);
or U2225 (N_2225,In_623,In_680);
nor U2226 (N_2226,In_678,In_557);
or U2227 (N_2227,In_513,In_672);
and U2228 (N_2228,In_69,In_277);
nand U2229 (N_2229,In_663,In_211);
or U2230 (N_2230,In_482,In_628);
nand U2231 (N_2231,In_452,In_293);
nor U2232 (N_2232,In_526,In_191);
and U2233 (N_2233,In_140,In_384);
nor U2234 (N_2234,In_115,In_216);
nand U2235 (N_2235,In_426,In_358);
or U2236 (N_2236,In_60,In_410);
or U2237 (N_2237,In_602,In_263);
nand U2238 (N_2238,In_240,In_392);
and U2239 (N_2239,In_141,In_14);
or U2240 (N_2240,In_534,In_575);
nand U2241 (N_2241,In_117,In_590);
and U2242 (N_2242,In_241,In_285);
and U2243 (N_2243,In_688,In_75);
and U2244 (N_2244,In_131,In_115);
nand U2245 (N_2245,In_195,In_13);
nand U2246 (N_2246,In_631,In_315);
and U2247 (N_2247,In_648,In_18);
nand U2248 (N_2248,In_396,In_400);
and U2249 (N_2249,In_378,In_277);
nor U2250 (N_2250,In_383,In_720);
xor U2251 (N_2251,In_306,In_349);
or U2252 (N_2252,In_689,In_167);
nand U2253 (N_2253,In_34,In_691);
xnor U2254 (N_2254,In_15,In_551);
xnor U2255 (N_2255,In_202,In_379);
or U2256 (N_2256,In_225,In_205);
nor U2257 (N_2257,In_141,In_189);
or U2258 (N_2258,In_350,In_611);
xnor U2259 (N_2259,In_163,In_368);
or U2260 (N_2260,In_679,In_98);
and U2261 (N_2261,In_25,In_468);
nand U2262 (N_2262,In_471,In_362);
nand U2263 (N_2263,In_356,In_387);
xnor U2264 (N_2264,In_18,In_358);
xnor U2265 (N_2265,In_544,In_128);
nand U2266 (N_2266,In_162,In_688);
and U2267 (N_2267,In_627,In_737);
nand U2268 (N_2268,In_295,In_48);
and U2269 (N_2269,In_647,In_640);
xor U2270 (N_2270,In_585,In_217);
and U2271 (N_2271,In_530,In_302);
nand U2272 (N_2272,In_607,In_445);
nand U2273 (N_2273,In_80,In_119);
nand U2274 (N_2274,In_352,In_113);
nor U2275 (N_2275,In_201,In_678);
and U2276 (N_2276,In_253,In_359);
nor U2277 (N_2277,In_14,In_115);
nor U2278 (N_2278,In_171,In_360);
nand U2279 (N_2279,In_418,In_341);
or U2280 (N_2280,In_598,In_641);
nor U2281 (N_2281,In_487,In_568);
nand U2282 (N_2282,In_96,In_168);
or U2283 (N_2283,In_477,In_30);
nor U2284 (N_2284,In_329,In_413);
and U2285 (N_2285,In_735,In_294);
or U2286 (N_2286,In_290,In_429);
and U2287 (N_2287,In_142,In_432);
nand U2288 (N_2288,In_257,In_135);
xor U2289 (N_2289,In_708,In_247);
or U2290 (N_2290,In_84,In_456);
or U2291 (N_2291,In_499,In_252);
xnor U2292 (N_2292,In_35,In_529);
or U2293 (N_2293,In_486,In_367);
xnor U2294 (N_2294,In_227,In_658);
or U2295 (N_2295,In_568,In_257);
or U2296 (N_2296,In_414,In_267);
xnor U2297 (N_2297,In_153,In_50);
nand U2298 (N_2298,In_33,In_480);
xor U2299 (N_2299,In_331,In_323);
nand U2300 (N_2300,In_506,In_422);
nor U2301 (N_2301,In_275,In_387);
nor U2302 (N_2302,In_79,In_66);
nor U2303 (N_2303,In_43,In_47);
and U2304 (N_2304,In_48,In_621);
or U2305 (N_2305,In_251,In_612);
or U2306 (N_2306,In_602,In_395);
nand U2307 (N_2307,In_559,In_86);
or U2308 (N_2308,In_718,In_85);
nand U2309 (N_2309,In_423,In_688);
nor U2310 (N_2310,In_79,In_202);
and U2311 (N_2311,In_74,In_666);
nor U2312 (N_2312,In_221,In_2);
nor U2313 (N_2313,In_514,In_66);
and U2314 (N_2314,In_176,In_693);
xnor U2315 (N_2315,In_657,In_674);
and U2316 (N_2316,In_65,In_295);
xnor U2317 (N_2317,In_450,In_71);
and U2318 (N_2318,In_548,In_649);
nor U2319 (N_2319,In_556,In_644);
or U2320 (N_2320,In_590,In_388);
or U2321 (N_2321,In_662,In_112);
and U2322 (N_2322,In_328,In_206);
nor U2323 (N_2323,In_384,In_264);
nand U2324 (N_2324,In_456,In_119);
and U2325 (N_2325,In_272,In_321);
xnor U2326 (N_2326,In_405,In_510);
nor U2327 (N_2327,In_726,In_145);
or U2328 (N_2328,In_428,In_569);
xor U2329 (N_2329,In_1,In_657);
xor U2330 (N_2330,In_316,In_540);
and U2331 (N_2331,In_545,In_593);
nor U2332 (N_2332,In_115,In_214);
nand U2333 (N_2333,In_546,In_11);
and U2334 (N_2334,In_310,In_140);
nand U2335 (N_2335,In_573,In_175);
or U2336 (N_2336,In_134,In_590);
nor U2337 (N_2337,In_678,In_558);
or U2338 (N_2338,In_49,In_328);
or U2339 (N_2339,In_160,In_98);
nand U2340 (N_2340,In_116,In_270);
and U2341 (N_2341,In_262,In_447);
and U2342 (N_2342,In_251,In_678);
xnor U2343 (N_2343,In_369,In_295);
or U2344 (N_2344,In_499,In_232);
and U2345 (N_2345,In_528,In_240);
nand U2346 (N_2346,In_121,In_262);
nand U2347 (N_2347,In_467,In_648);
nor U2348 (N_2348,In_76,In_53);
xor U2349 (N_2349,In_539,In_206);
or U2350 (N_2350,In_323,In_197);
or U2351 (N_2351,In_143,In_199);
or U2352 (N_2352,In_603,In_317);
and U2353 (N_2353,In_122,In_370);
and U2354 (N_2354,In_393,In_288);
nand U2355 (N_2355,In_519,In_733);
nand U2356 (N_2356,In_298,In_117);
and U2357 (N_2357,In_118,In_316);
or U2358 (N_2358,In_271,In_67);
xnor U2359 (N_2359,In_38,In_353);
nand U2360 (N_2360,In_350,In_17);
nor U2361 (N_2361,In_92,In_373);
or U2362 (N_2362,In_521,In_298);
nand U2363 (N_2363,In_394,In_384);
and U2364 (N_2364,In_217,In_742);
nand U2365 (N_2365,In_438,In_583);
and U2366 (N_2366,In_407,In_1);
xnor U2367 (N_2367,In_325,In_455);
nand U2368 (N_2368,In_177,In_714);
nor U2369 (N_2369,In_104,In_607);
nand U2370 (N_2370,In_602,In_552);
nand U2371 (N_2371,In_653,In_667);
nand U2372 (N_2372,In_574,In_255);
nor U2373 (N_2373,In_687,In_534);
nand U2374 (N_2374,In_69,In_428);
and U2375 (N_2375,In_290,In_583);
nor U2376 (N_2376,In_667,In_293);
or U2377 (N_2377,In_307,In_252);
nand U2378 (N_2378,In_559,In_699);
nand U2379 (N_2379,In_365,In_403);
and U2380 (N_2380,In_396,In_145);
nand U2381 (N_2381,In_560,In_506);
nor U2382 (N_2382,In_670,In_136);
xnor U2383 (N_2383,In_605,In_88);
and U2384 (N_2384,In_561,In_536);
or U2385 (N_2385,In_315,In_306);
and U2386 (N_2386,In_554,In_84);
nand U2387 (N_2387,In_453,In_243);
xor U2388 (N_2388,In_13,In_717);
nand U2389 (N_2389,In_621,In_547);
nor U2390 (N_2390,In_208,In_220);
and U2391 (N_2391,In_216,In_345);
or U2392 (N_2392,In_618,In_353);
nor U2393 (N_2393,In_608,In_4);
or U2394 (N_2394,In_422,In_544);
and U2395 (N_2395,In_206,In_609);
and U2396 (N_2396,In_155,In_631);
or U2397 (N_2397,In_749,In_346);
or U2398 (N_2398,In_384,In_303);
nor U2399 (N_2399,In_617,In_66);
nor U2400 (N_2400,In_247,In_627);
and U2401 (N_2401,In_8,In_518);
nand U2402 (N_2402,In_112,In_496);
and U2403 (N_2403,In_90,In_294);
xor U2404 (N_2404,In_183,In_149);
nor U2405 (N_2405,In_694,In_99);
xor U2406 (N_2406,In_708,In_357);
and U2407 (N_2407,In_374,In_467);
and U2408 (N_2408,In_656,In_115);
nand U2409 (N_2409,In_248,In_47);
nor U2410 (N_2410,In_86,In_515);
nand U2411 (N_2411,In_239,In_296);
nor U2412 (N_2412,In_365,In_361);
nor U2413 (N_2413,In_4,In_610);
nand U2414 (N_2414,In_502,In_210);
or U2415 (N_2415,In_447,In_127);
and U2416 (N_2416,In_608,In_291);
nand U2417 (N_2417,In_246,In_183);
nor U2418 (N_2418,In_700,In_354);
or U2419 (N_2419,In_308,In_38);
nand U2420 (N_2420,In_663,In_685);
nand U2421 (N_2421,In_607,In_30);
and U2422 (N_2422,In_562,In_510);
nor U2423 (N_2423,In_278,In_495);
and U2424 (N_2424,In_345,In_748);
nand U2425 (N_2425,In_114,In_206);
or U2426 (N_2426,In_28,In_296);
and U2427 (N_2427,In_281,In_730);
xnor U2428 (N_2428,In_231,In_367);
nor U2429 (N_2429,In_660,In_203);
or U2430 (N_2430,In_198,In_18);
nor U2431 (N_2431,In_73,In_540);
or U2432 (N_2432,In_306,In_112);
or U2433 (N_2433,In_264,In_220);
or U2434 (N_2434,In_43,In_446);
xnor U2435 (N_2435,In_170,In_282);
nand U2436 (N_2436,In_220,In_255);
xor U2437 (N_2437,In_59,In_706);
nor U2438 (N_2438,In_83,In_285);
and U2439 (N_2439,In_73,In_313);
nand U2440 (N_2440,In_50,In_341);
or U2441 (N_2441,In_10,In_19);
and U2442 (N_2442,In_147,In_251);
or U2443 (N_2443,In_491,In_290);
xor U2444 (N_2444,In_258,In_736);
nand U2445 (N_2445,In_621,In_488);
xor U2446 (N_2446,In_481,In_150);
nor U2447 (N_2447,In_202,In_62);
nor U2448 (N_2448,In_26,In_349);
and U2449 (N_2449,In_719,In_177);
xnor U2450 (N_2450,In_96,In_383);
xor U2451 (N_2451,In_442,In_159);
nor U2452 (N_2452,In_488,In_533);
or U2453 (N_2453,In_522,In_154);
nor U2454 (N_2454,In_140,In_728);
nand U2455 (N_2455,In_293,In_464);
nand U2456 (N_2456,In_304,In_617);
nand U2457 (N_2457,In_388,In_634);
and U2458 (N_2458,In_488,In_293);
or U2459 (N_2459,In_597,In_126);
and U2460 (N_2460,In_158,In_626);
and U2461 (N_2461,In_237,In_747);
nand U2462 (N_2462,In_691,In_333);
nor U2463 (N_2463,In_9,In_78);
nor U2464 (N_2464,In_121,In_532);
nor U2465 (N_2465,In_641,In_6);
nor U2466 (N_2466,In_594,In_385);
nor U2467 (N_2467,In_443,In_487);
xor U2468 (N_2468,In_280,In_672);
nand U2469 (N_2469,In_166,In_303);
nor U2470 (N_2470,In_260,In_530);
nand U2471 (N_2471,In_440,In_659);
xnor U2472 (N_2472,In_59,In_664);
nand U2473 (N_2473,In_568,In_403);
nor U2474 (N_2474,In_470,In_333);
or U2475 (N_2475,In_286,In_587);
and U2476 (N_2476,In_743,In_348);
and U2477 (N_2477,In_697,In_686);
nor U2478 (N_2478,In_620,In_100);
nor U2479 (N_2479,In_438,In_637);
or U2480 (N_2480,In_97,In_379);
or U2481 (N_2481,In_45,In_22);
nor U2482 (N_2482,In_518,In_451);
and U2483 (N_2483,In_359,In_464);
or U2484 (N_2484,In_505,In_229);
nand U2485 (N_2485,In_341,In_190);
or U2486 (N_2486,In_640,In_343);
nor U2487 (N_2487,In_44,In_114);
xor U2488 (N_2488,In_98,In_51);
or U2489 (N_2489,In_385,In_176);
or U2490 (N_2490,In_226,In_716);
and U2491 (N_2491,In_432,In_470);
or U2492 (N_2492,In_311,In_672);
nand U2493 (N_2493,In_451,In_631);
nand U2494 (N_2494,In_216,In_700);
nand U2495 (N_2495,In_692,In_480);
and U2496 (N_2496,In_170,In_697);
and U2497 (N_2497,In_236,In_496);
or U2498 (N_2498,In_226,In_125);
xor U2499 (N_2499,In_558,In_465);
or U2500 (N_2500,N_2048,N_990);
nor U2501 (N_2501,N_1925,N_1100);
or U2502 (N_2502,N_1782,N_1634);
or U2503 (N_2503,N_847,N_322);
or U2504 (N_2504,N_242,N_1933);
xor U2505 (N_2505,N_1276,N_1238);
nand U2506 (N_2506,N_142,N_2349);
nand U2507 (N_2507,N_736,N_1293);
and U2508 (N_2508,N_385,N_906);
or U2509 (N_2509,N_591,N_1303);
and U2510 (N_2510,N_2463,N_1363);
or U2511 (N_2511,N_860,N_634);
xor U2512 (N_2512,N_1486,N_2232);
and U2513 (N_2513,N_37,N_903);
nand U2514 (N_2514,N_1772,N_840);
xor U2515 (N_2515,N_1991,N_2462);
and U2516 (N_2516,N_1852,N_909);
nand U2517 (N_2517,N_1643,N_1013);
or U2518 (N_2518,N_1329,N_1483);
xnor U2519 (N_2519,N_375,N_2088);
or U2520 (N_2520,N_1855,N_1678);
or U2521 (N_2521,N_1281,N_2243);
nand U2522 (N_2522,N_1858,N_2234);
nor U2523 (N_2523,N_907,N_978);
or U2524 (N_2524,N_1190,N_1155);
nand U2525 (N_2525,N_2411,N_1242);
nor U2526 (N_2526,N_2493,N_1947);
and U2527 (N_2527,N_2062,N_1971);
nand U2528 (N_2528,N_729,N_2258);
or U2529 (N_2529,N_75,N_2076);
and U2530 (N_2530,N_1326,N_1767);
or U2531 (N_2531,N_1975,N_1106);
xnor U2532 (N_2532,N_1628,N_1735);
nor U2533 (N_2533,N_225,N_129);
or U2534 (N_2534,N_2191,N_2229);
xor U2535 (N_2535,N_1224,N_1342);
nor U2536 (N_2536,N_293,N_394);
or U2537 (N_2537,N_2253,N_1951);
and U2538 (N_2538,N_984,N_1079);
or U2539 (N_2539,N_2492,N_198);
or U2540 (N_2540,N_1537,N_122);
and U2541 (N_2541,N_1640,N_1269);
xor U2542 (N_2542,N_2231,N_28);
and U2543 (N_2543,N_2030,N_2302);
and U2544 (N_2544,N_238,N_2329);
nor U2545 (N_2545,N_1567,N_880);
nand U2546 (N_2546,N_1710,N_1532);
or U2547 (N_2547,N_1692,N_557);
or U2548 (N_2548,N_1422,N_1854);
nor U2549 (N_2549,N_703,N_160);
nand U2550 (N_2550,N_698,N_1967);
or U2551 (N_2551,N_1430,N_699);
nand U2552 (N_2552,N_2380,N_27);
nor U2553 (N_2553,N_2063,N_559);
and U2554 (N_2554,N_1774,N_423);
or U2555 (N_2555,N_393,N_71);
nand U2556 (N_2556,N_153,N_1859);
nand U2557 (N_2557,N_945,N_2104);
xnor U2558 (N_2558,N_446,N_1479);
nor U2559 (N_2559,N_1529,N_1445);
xnor U2560 (N_2560,N_1627,N_949);
nand U2561 (N_2561,N_1256,N_959);
and U2562 (N_2562,N_2476,N_10);
nand U2563 (N_2563,N_1139,N_2296);
nand U2564 (N_2564,N_86,N_53);
nor U2565 (N_2565,N_1345,N_60);
and U2566 (N_2566,N_1017,N_392);
nor U2567 (N_2567,N_97,N_1212);
xnor U2568 (N_2568,N_2373,N_2409);
xnor U2569 (N_2569,N_2326,N_1667);
and U2570 (N_2570,N_2321,N_1094);
and U2571 (N_2571,N_124,N_1982);
nand U2572 (N_2572,N_2085,N_1525);
nand U2573 (N_2573,N_1557,N_2135);
or U2574 (N_2574,N_1456,N_606);
nand U2575 (N_2575,N_307,N_994);
and U2576 (N_2576,N_2410,N_2224);
and U2577 (N_2577,N_713,N_2152);
and U2578 (N_2578,N_512,N_756);
nand U2579 (N_2579,N_1372,N_1175);
xor U2580 (N_2580,N_650,N_1336);
or U2581 (N_2581,N_700,N_779);
nor U2582 (N_2582,N_723,N_955);
nor U2583 (N_2583,N_795,N_323);
nor U2584 (N_2584,N_832,N_1516);
xor U2585 (N_2585,N_625,N_731);
or U2586 (N_2586,N_600,N_1332);
and U2587 (N_2587,N_1084,N_2471);
nor U2588 (N_2588,N_962,N_1904);
nor U2589 (N_2589,N_1791,N_2490);
nand U2590 (N_2590,N_883,N_1492);
nand U2591 (N_2591,N_876,N_1434);
nand U2592 (N_2592,N_509,N_1085);
nor U2593 (N_2593,N_2246,N_1458);
or U2594 (N_2594,N_2312,N_1837);
nand U2595 (N_2595,N_2360,N_1821);
nand U2596 (N_2596,N_1878,N_2036);
nand U2597 (N_2597,N_975,N_1810);
or U2598 (N_2598,N_1104,N_2004);
nand U2599 (N_2599,N_1042,N_62);
or U2600 (N_2600,N_1939,N_2173);
nand U2601 (N_2601,N_1273,N_1552);
or U2602 (N_2602,N_1072,N_1311);
or U2603 (N_2603,N_288,N_1550);
nand U2604 (N_2604,N_2215,N_987);
xor U2605 (N_2605,N_867,N_1425);
nand U2606 (N_2606,N_1331,N_2014);
nand U2607 (N_2607,N_2335,N_635);
nor U2608 (N_2608,N_531,N_849);
nor U2609 (N_2609,N_789,N_2041);
nand U2610 (N_2610,N_1760,N_834);
nor U2611 (N_2611,N_1133,N_36);
nor U2612 (N_2612,N_1188,N_735);
nand U2613 (N_2613,N_398,N_1513);
xor U2614 (N_2614,N_1304,N_1615);
nor U2615 (N_2615,N_809,N_105);
nor U2616 (N_2616,N_1356,N_2180);
and U2617 (N_2617,N_1368,N_1503);
and U2618 (N_2618,N_1769,N_1229);
and U2619 (N_2619,N_205,N_672);
or U2620 (N_2620,N_953,N_197);
nor U2621 (N_2621,N_577,N_2415);
xor U2622 (N_2622,N_1301,N_960);
nand U2623 (N_2623,N_1669,N_1547);
and U2624 (N_2624,N_561,N_312);
nor U2625 (N_2625,N_1931,N_2439);
nor U2626 (N_2626,N_2431,N_482);
nand U2627 (N_2627,N_131,N_265);
nand U2628 (N_2628,N_2397,N_988);
or U2629 (N_2629,N_176,N_2128);
nor U2630 (N_2630,N_436,N_985);
nor U2631 (N_2631,N_373,N_245);
nand U2632 (N_2632,N_817,N_1871);
nor U2633 (N_2633,N_1376,N_553);
or U2634 (N_2634,N_275,N_2118);
nand U2635 (N_2635,N_2341,N_718);
nor U2636 (N_2636,N_501,N_1785);
or U2637 (N_2637,N_643,N_1973);
nor U2638 (N_2638,N_1703,N_228);
or U2639 (N_2639,N_2096,N_2137);
and U2640 (N_2640,N_1324,N_355);
and U2641 (N_2641,N_2361,N_280);
nand U2642 (N_2642,N_1839,N_1286);
and U2643 (N_2643,N_1950,N_1515);
or U2644 (N_2644,N_1490,N_1020);
nor U2645 (N_2645,N_2346,N_136);
and U2646 (N_2646,N_51,N_1462);
and U2647 (N_2647,N_2042,N_2115);
or U2648 (N_2648,N_1151,N_497);
or U2649 (N_2649,N_434,N_301);
nand U2650 (N_2650,N_2239,N_1524);
xor U2651 (N_2651,N_1051,N_680);
or U2652 (N_2652,N_1876,N_1637);
or U2653 (N_2653,N_2452,N_399);
nor U2654 (N_2654,N_1087,N_461);
or U2655 (N_2655,N_2130,N_426);
and U2656 (N_2656,N_403,N_1758);
nand U2657 (N_2657,N_1285,N_954);
xnor U2658 (N_2658,N_1246,N_964);
nor U2659 (N_2659,N_976,N_784);
nor U2660 (N_2660,N_1204,N_1375);
nor U2661 (N_2661,N_2363,N_1617);
nand U2662 (N_2662,N_1221,N_2049);
nor U2663 (N_2663,N_266,N_1738);
nand U2664 (N_2664,N_2278,N_2060);
and U2665 (N_2665,N_2156,N_2356);
xor U2666 (N_2666,N_758,N_1753);
and U2667 (N_2667,N_1295,N_585);
nand U2668 (N_2668,N_1977,N_2377);
nand U2669 (N_2669,N_1442,N_421);
and U2670 (N_2670,N_1665,N_708);
and U2671 (N_2671,N_1431,N_1092);
nor U2672 (N_2672,N_31,N_1433);
nand U2673 (N_2673,N_1568,N_2305);
or U2674 (N_2674,N_1834,N_1441);
or U2675 (N_2675,N_1218,N_1943);
and U2676 (N_2676,N_751,N_304);
nor U2677 (N_2677,N_1408,N_739);
and U2678 (N_2678,N_412,N_243);
and U2679 (N_2679,N_41,N_2073);
and U2680 (N_2680,N_2161,N_1327);
or U2681 (N_2681,N_1350,N_1340);
or U2682 (N_2682,N_326,N_939);
nor U2683 (N_2683,N_668,N_294);
nor U2684 (N_2684,N_720,N_2083);
nand U2685 (N_2685,N_530,N_1806);
nor U2686 (N_2686,N_2392,N_2082);
nand U2687 (N_2687,N_1602,N_948);
or U2688 (N_2688,N_1820,N_804);
nand U2689 (N_2689,N_1310,N_2074);
or U2690 (N_2690,N_2008,N_598);
nand U2691 (N_2691,N_231,N_2263);
xor U2692 (N_2692,N_2287,N_1614);
or U2693 (N_2693,N_110,N_802);
nor U2694 (N_2694,N_1842,N_440);
nor U2695 (N_2695,N_1205,N_1621);
nor U2696 (N_2696,N_902,N_1385);
and U2697 (N_2697,N_40,N_15);
xnor U2698 (N_2698,N_2383,N_1118);
nor U2699 (N_2699,N_631,N_678);
nand U2700 (N_2700,N_13,N_193);
nor U2701 (N_2701,N_1805,N_1527);
nand U2702 (N_2702,N_725,N_1910);
and U2703 (N_2703,N_1644,N_661);
xnor U2704 (N_2704,N_1535,N_882);
or U2705 (N_2705,N_647,N_670);
xnor U2706 (N_2706,N_1123,N_574);
xnor U2707 (N_2707,N_646,N_2475);
nand U2708 (N_2708,N_1722,N_16);
and U2709 (N_2709,N_1231,N_2067);
or U2710 (N_2710,N_1704,N_1661);
nand U2711 (N_2711,N_1325,N_2190);
xnor U2712 (N_2712,N_924,N_73);
nand U2713 (N_2713,N_632,N_290);
or U2714 (N_2714,N_2388,N_1193);
or U2715 (N_2715,N_1283,N_1344);
nand U2716 (N_2716,N_582,N_1631);
nand U2717 (N_2717,N_1504,N_32);
or U2718 (N_2718,N_185,N_256);
nand U2719 (N_2719,N_1245,N_68);
or U2720 (N_2720,N_492,N_1194);
nand U2721 (N_2721,N_1500,N_2034);
or U2722 (N_2722,N_523,N_2295);
nor U2723 (N_2723,N_1158,N_732);
nand U2724 (N_2724,N_755,N_207);
or U2725 (N_2725,N_705,N_2252);
xor U2726 (N_2726,N_536,N_1371);
nor U2727 (N_2727,N_1777,N_2017);
or U2728 (N_2728,N_2185,N_1742);
nor U2729 (N_2729,N_586,N_363);
or U2730 (N_2730,N_337,N_1996);
nand U2731 (N_2731,N_1149,N_397);
or U2732 (N_2732,N_2264,N_578);
or U2733 (N_2733,N_2342,N_1401);
nand U2734 (N_2734,N_1400,N_1872);
nor U2735 (N_2735,N_645,N_1302);
nor U2736 (N_2736,N_1157,N_2218);
and U2737 (N_2737,N_1496,N_2106);
and U2738 (N_2738,N_1594,N_109);
nand U2739 (N_2739,N_319,N_1612);
xnor U2740 (N_2740,N_69,N_1195);
nor U2741 (N_2741,N_191,N_2248);
nor U2742 (N_2742,N_730,N_885);
xor U2743 (N_2743,N_360,N_630);
nand U2744 (N_2744,N_212,N_2095);
nand U2745 (N_2745,N_1998,N_1747);
or U2746 (N_2746,N_1506,N_547);
and U2747 (N_2747,N_1688,N_1126);
nor U2748 (N_2748,N_2169,N_338);
nor U2749 (N_2749,N_1217,N_2094);
or U2750 (N_2750,N_1341,N_112);
xor U2751 (N_2751,N_685,N_1952);
nand U2752 (N_2752,N_2027,N_64);
and U2753 (N_2753,N_133,N_659);
nor U2754 (N_2754,N_1768,N_490);
or U2755 (N_2755,N_223,N_590);
xor U2756 (N_2756,N_1618,N_2168);
xnor U2757 (N_2757,N_2434,N_286);
nand U2758 (N_2758,N_1095,N_2407);
xnor U2759 (N_2759,N_1247,N_979);
and U2760 (N_2760,N_2176,N_210);
nor U2761 (N_2761,N_132,N_2100);
nand U2762 (N_2762,N_1163,N_1330);
nor U2763 (N_2763,N_947,N_963);
nand U2764 (N_2764,N_100,N_180);
nor U2765 (N_2765,N_2226,N_2289);
or U2766 (N_2766,N_1891,N_1164);
and U2767 (N_2767,N_2390,N_371);
nand U2768 (N_2768,N_116,N_2480);
xor U2769 (N_2769,N_213,N_1987);
nor U2770 (N_2770,N_1134,N_179);
nand U2771 (N_2771,N_1266,N_1455);
nand U2772 (N_2772,N_820,N_1875);
nor U2773 (N_2773,N_2171,N_734);
and U2774 (N_2774,N_253,N_930);
or U2775 (N_2775,N_1358,N_113);
xor U2776 (N_2776,N_2098,N_1197);
xnor U2777 (N_2777,N_415,N_1160);
or U2778 (N_2778,N_2160,N_727);
nand U2779 (N_2779,N_2102,N_1551);
nand U2780 (N_2780,N_2086,N_749);
or U2781 (N_2781,N_93,N_1646);
and U2782 (N_2782,N_194,N_1071);
and U2783 (N_2783,N_1406,N_858);
and U2784 (N_2784,N_1635,N_1885);
and U2785 (N_2785,N_366,N_2153);
xnor U2786 (N_2786,N_1489,N_701);
and U2787 (N_2787,N_410,N_1869);
and U2788 (N_2788,N_1491,N_236);
nand U2789 (N_2789,N_2270,N_1625);
nor U2790 (N_2790,N_1008,N_1592);
xnor U2791 (N_2791,N_1461,N_2472);
nor U2792 (N_2792,N_527,N_413);
or U2793 (N_2793,N_1879,N_1265);
nor U2794 (N_2794,N_2110,N_2449);
nor U2795 (N_2795,N_824,N_1047);
nand U2796 (N_2796,N_993,N_1314);
nand U2797 (N_2797,N_539,N_2142);
nor U2798 (N_2798,N_409,N_1167);
nand U2799 (N_2799,N_1898,N_447);
nor U2800 (N_2800,N_2369,N_1874);
nor U2801 (N_2801,N_1209,N_2251);
and U2802 (N_2802,N_1979,N_1915);
nand U2803 (N_2803,N_1367,N_619);
xor U2804 (N_2804,N_147,N_1850);
or U2805 (N_2805,N_555,N_794);
and U2806 (N_2806,N_1282,N_311);
nor U2807 (N_2807,N_1705,N_584);
or U2808 (N_2808,N_919,N_2372);
or U2809 (N_2809,N_247,N_216);
nor U2810 (N_2810,N_2491,N_1112);
nand U2811 (N_2811,N_80,N_2365);
nand U2812 (N_2812,N_487,N_1248);
or U2813 (N_2813,N_433,N_2238);
and U2814 (N_2814,N_1029,N_1130);
nand U2815 (N_2815,N_372,N_2453);
and U2816 (N_2816,N_2144,N_1591);
nand U2817 (N_2817,N_1039,N_778);
and U2818 (N_2818,N_2265,N_548);
and U2819 (N_2819,N_277,N_358);
and U2820 (N_2820,N_359,N_1253);
and U2821 (N_2821,N_2136,N_2320);
nor U2822 (N_2822,N_2464,N_1361);
xnor U2823 (N_2823,N_34,N_1143);
nand U2824 (N_2824,N_2023,N_502);
xor U2825 (N_2825,N_932,N_1170);
nor U2826 (N_2826,N_1183,N_1781);
nand U2827 (N_2827,N_1168,N_967);
and U2828 (N_2828,N_1423,N_445);
or U2829 (N_2829,N_335,N_2236);
and U2830 (N_2830,N_1147,N_1860);
nor U2831 (N_2831,N_186,N_856);
nor U2832 (N_2832,N_2366,N_1261);
nand U2833 (N_2833,N_382,N_569);
and U2834 (N_2834,N_2033,N_1630);
and U2835 (N_2835,N_2223,N_515);
and U2836 (N_2836,N_871,N_98);
xnor U2837 (N_2837,N_786,N_1485);
xor U2838 (N_2838,N_1861,N_521);
nor U2839 (N_2839,N_1177,N_981);
and U2840 (N_2840,N_538,N_428);
nand U2841 (N_2841,N_2072,N_1090);
nand U2842 (N_2842,N_320,N_158);
or U2843 (N_2843,N_1714,N_1577);
nand U2844 (N_2844,N_164,N_1558);
and U2845 (N_2845,N_940,N_1351);
or U2846 (N_2846,N_1578,N_1917);
xnor U2847 (N_2847,N_872,N_1011);
or U2848 (N_2848,N_2199,N_361);
and U2849 (N_2849,N_1587,N_2337);
and U2850 (N_2850,N_762,N_2133);
nand U2851 (N_2851,N_2001,N_1409);
nor U2852 (N_2852,N_2007,N_1945);
nand U2853 (N_2853,N_1942,N_2026);
nand U2854 (N_2854,N_298,N_2163);
and U2855 (N_2855,N_268,N_1921);
or U2856 (N_2856,N_777,N_1181);
xnor U2857 (N_2857,N_169,N_922);
nor U2858 (N_2858,N_407,N_904);
and U2859 (N_2859,N_957,N_1001);
and U2860 (N_2860,N_2192,N_55);
or U2861 (N_2861,N_2194,N_1595);
xnor U2862 (N_2862,N_2286,N_2458);
xor U2863 (N_2863,N_696,N_1415);
and U2864 (N_2864,N_1115,N_633);
xor U2865 (N_2865,N_1228,N_90);
nor U2866 (N_2866,N_318,N_263);
nand U2867 (N_2867,N_1546,N_1022);
nand U2868 (N_2868,N_1660,N_1682);
nor U2869 (N_2869,N_914,N_1505);
and U2870 (N_2870,N_1469,N_1420);
and U2871 (N_2871,N_517,N_738);
and U2872 (N_2872,N_2149,N_2276);
and U2873 (N_2873,N_1699,N_1037);
nand U2874 (N_2874,N_1596,N_1294);
nand U2875 (N_2875,N_1866,N_2284);
nand U2876 (N_2876,N_91,N_1521);
nor U2877 (N_2877,N_1729,N_2375);
nor U2878 (N_2878,N_936,N_565);
nand U2879 (N_2879,N_1148,N_1884);
or U2880 (N_2880,N_1339,N_1202);
or U2881 (N_2881,N_781,N_1746);
nor U2882 (N_2882,N_2053,N_1562);
xor U2883 (N_2883,N_893,N_1053);
and U2884 (N_2884,N_343,N_908);
or U2885 (N_2885,N_1452,N_2138);
or U2886 (N_2886,N_336,N_1585);
and U2887 (N_2887,N_261,N_1645);
or U2888 (N_2888,N_2469,N_76);
xor U2889 (N_2889,N_1993,N_1082);
or U2890 (N_2890,N_1284,N_1334);
xnor U2891 (N_2891,N_1225,N_47);
and U2892 (N_2892,N_2131,N_1322);
nor U2893 (N_2893,N_430,N_844);
and U2894 (N_2894,N_1187,N_1739);
and U2895 (N_2895,N_1374,N_1241);
and U2896 (N_2896,N_1033,N_706);
or U2897 (N_2897,N_2396,N_1025);
nor U2898 (N_2898,N_2237,N_195);
nand U2899 (N_2899,N_471,N_1718);
nand U2900 (N_2900,N_588,N_1684);
and U2901 (N_2901,N_1610,N_2241);
nor U2902 (N_2902,N_162,N_2166);
and U2903 (N_2903,N_192,N_101);
and U2904 (N_2904,N_2359,N_2078);
nor U2905 (N_2905,N_230,N_1299);
or U2906 (N_2906,N_1814,N_1240);
nor U2907 (N_2907,N_613,N_2351);
or U2908 (N_2908,N_1905,N_791);
nand U2909 (N_2909,N_1908,N_2268);
nand U2910 (N_2910,N_878,N_1813);
nand U2911 (N_2911,N_839,N_2306);
nand U2912 (N_2912,N_989,N_237);
and U2913 (N_2913,N_2092,N_2101);
nor U2914 (N_2914,N_1156,N_1373);
nor U2915 (N_2915,N_2179,N_1178);
and U2916 (N_2916,N_1320,N_349);
nand U2917 (N_2917,N_1892,N_2440);
nand U2918 (N_2918,N_251,N_1089);
or U2919 (N_2919,N_1726,N_2456);
or U2920 (N_2920,N_383,N_1654);
and U2921 (N_2921,N_1426,N_309);
or U2922 (N_2922,N_2164,N_1648);
nand U2923 (N_2923,N_1459,N_235);
and U2924 (N_2924,N_1763,N_175);
nor U2925 (N_2925,N_2205,N_719);
and U2926 (N_2926,N_119,N_405);
or U2927 (N_2927,N_272,N_1239);
nor U2928 (N_2928,N_1545,N_1709);
or U2929 (N_2929,N_295,N_799);
nand U2930 (N_2930,N_1446,N_1472);
or U2931 (N_2931,N_1399,N_1306);
and U2932 (N_2932,N_641,N_1750);
nor U2933 (N_2933,N_334,N_1838);
nor U2934 (N_2934,N_768,N_1223);
nor U2935 (N_2935,N_388,N_833);
or U2936 (N_2936,N_2266,N_687);
and U2937 (N_2937,N_1882,N_1605);
and U2938 (N_2938,N_1354,N_1257);
and U2939 (N_2939,N_339,N_644);
nand U2940 (N_2940,N_2024,N_1728);
nor U2941 (N_2941,N_1117,N_329);
xnor U2942 (N_2942,N_1288,N_541);
or U2943 (N_2943,N_2057,N_2162);
nor U2944 (N_2944,N_1230,N_1553);
and U2945 (N_2945,N_798,N_1966);
nor U2946 (N_2946,N_890,N_836);
nor U2947 (N_2947,N_1902,N_1538);
nor U2948 (N_2948,N_2386,N_2124);
and U2949 (N_2949,N_1676,N_346);
xnor U2950 (N_2950,N_2277,N_348);
nand U2951 (N_2951,N_823,N_1509);
and U2952 (N_2952,N_594,N_2400);
and U2953 (N_2953,N_1517,N_20);
or U2954 (N_2954,N_1825,N_505);
xnor U2955 (N_2955,N_563,N_693);
nor U2956 (N_2956,N_1036,N_1543);
and U2957 (N_2957,N_604,N_2354);
nand U2958 (N_2958,N_827,N_1641);
nand U2959 (N_2959,N_1141,N_2299);
nor U2960 (N_2960,N_1895,N_760);
or U2961 (N_2961,N_391,N_1833);
nand U2962 (N_2962,N_1903,N_2496);
nand U2963 (N_2963,N_660,N_395);
or U2964 (N_2964,N_362,N_1573);
nor U2965 (N_2965,N_1790,N_252);
or U2966 (N_2966,N_208,N_1108);
and U2967 (N_2967,N_18,N_1508);
or U2968 (N_2968,N_1271,N_1215);
xor U2969 (N_2969,N_1720,N_913);
and U2970 (N_2970,N_2260,N_550);
and U2971 (N_2971,N_365,N_170);
nor U2972 (N_2972,N_658,N_1493);
nand U2973 (N_2973,N_306,N_982);
nand U2974 (N_2974,N_854,N_1063);
nand U2975 (N_2975,N_1279,N_1102);
nand U2976 (N_2976,N_1122,N_1414);
nand U2977 (N_2977,N_2309,N_1407);
nand U2978 (N_2978,N_63,N_1666);
and U2979 (N_2979,N_2466,N_1715);
nor U2980 (N_2980,N_1909,N_1518);
nor U2981 (N_2981,N_2362,N_1800);
and U2982 (N_2982,N_776,N_494);
and U2983 (N_2983,N_797,N_2084);
nand U2984 (N_2984,N_1207,N_2244);
nor U2985 (N_2985,N_42,N_2291);
nand U2986 (N_2986,N_1073,N_1536);
or U2987 (N_2987,N_422,N_2290);
nor U2988 (N_2988,N_161,N_818);
and U2989 (N_2989,N_429,N_1249);
nand U2990 (N_2990,N_1983,N_1685);
nand U2991 (N_2991,N_652,N_2068);
and U2992 (N_2992,N_1632,N_411);
nor U2993 (N_2993,N_579,N_1976);
nand U2994 (N_2994,N_2498,N_1467);
or U2995 (N_2995,N_1989,N_1213);
nor U2996 (N_2996,N_316,N_137);
nor U2997 (N_2997,N_2451,N_287);
nor U2998 (N_2998,N_178,N_1044);
xnor U2999 (N_2999,N_1377,N_544);
and U3000 (N_3000,N_1724,N_1811);
nor U3001 (N_3001,N_499,N_1476);
nand U3002 (N_3002,N_414,N_1475);
or U3003 (N_3003,N_617,N_506);
nor U3004 (N_3004,N_464,N_1883);
and U3005 (N_3005,N_2297,N_1539);
and U3006 (N_3006,N_1817,N_765);
or U3007 (N_3007,N_1783,N_2221);
nand U3008 (N_3008,N_571,N_520);
or U3009 (N_3009,N_2145,N_2447);
nand U3010 (N_3010,N_1347,N_77);
and U3011 (N_3011,N_2435,N_2147);
nor U3012 (N_3012,N_1748,N_1);
xnor U3013 (N_3013,N_1636,N_2184);
nand U3014 (N_3014,N_896,N_742);
nor U3015 (N_3015,N_381,N_1649);
or U3016 (N_3016,N_2097,N_815);
nor U3017 (N_3017,N_2240,N_1992);
xnor U3018 (N_3018,N_886,N_895);
nand U3019 (N_3019,N_486,N_2210);
or U3020 (N_3020,N_115,N_992);
nand U3021 (N_3021,N_2230,N_333);
and U3022 (N_3022,N_1597,N_1323);
nor U3023 (N_3023,N_2433,N_2479);
nand U3024 (N_3024,N_1762,N_1848);
and U3025 (N_3025,N_1877,N_262);
nor U3026 (N_3026,N_2382,N_404);
nand U3027 (N_3027,N_1200,N_504);
nor U3028 (N_3028,N_917,N_2499);
and U3029 (N_3029,N_905,N_1994);
and U3030 (N_3030,N_1574,N_843);
nand U3031 (N_3031,N_968,N_2113);
nand U3032 (N_3032,N_1386,N_2355);
nand U3033 (N_3033,N_1639,N_928);
nand U3034 (N_3034,N_1220,N_1749);
or U3035 (N_3035,N_145,N_855);
or U3036 (N_3036,N_757,N_2140);
nand U3037 (N_3037,N_384,N_1671);
nor U3038 (N_3038,N_1730,N_146);
and U3039 (N_3039,N_1826,N_1383);
nor U3040 (N_3040,N_868,N_1934);
nor U3041 (N_3041,N_2324,N_546);
and U3042 (N_3042,N_828,N_273);
nor U3043 (N_3043,N_884,N_2304);
nand U3044 (N_3044,N_726,N_2141);
nor U3045 (N_3045,N_1424,N_656);
and U3046 (N_3046,N_1963,N_1473);
and U3047 (N_3047,N_1355,N_636);
and U3048 (N_3048,N_188,N_234);
or U3049 (N_3049,N_368,N_481);
xnor U3050 (N_3050,N_2352,N_996);
xor U3051 (N_3051,N_942,N_121);
nand U3052 (N_3052,N_1196,N_803);
and U3053 (N_3053,N_552,N_1978);
and U3054 (N_3054,N_219,N_79);
nor U3055 (N_3055,N_99,N_1651);
and U3056 (N_3056,N_528,N_460);
or U3057 (N_3057,N_717,N_33);
or U3058 (N_3058,N_424,N_1694);
or U3059 (N_3059,N_1566,N_1058);
or U3060 (N_3060,N_278,N_1049);
and U3061 (N_3061,N_1974,N_1731);
or U3062 (N_3062,N_1244,N_2020);
nand U3063 (N_3063,N_1589,N_1270);
nor U3064 (N_3064,N_759,N_853);
xnor U3065 (N_3065,N_1616,N_1721);
nor U3066 (N_3066,N_352,N_1129);
nand U3067 (N_3067,N_1512,N_1926);
and U3068 (N_3068,N_694,N_753);
or U3069 (N_3069,N_830,N_61);
xor U3070 (N_3070,N_2200,N_2436);
and U3071 (N_3071,N_1173,N_747);
nand U3072 (N_3072,N_1432,N_1289);
or U3073 (N_3073,N_941,N_1216);
nand U3074 (N_3074,N_1481,N_1262);
and U3075 (N_3075,N_354,N_87);
nor U3076 (N_3076,N_1064,N_163);
xnor U3077 (N_3077,N_1689,N_1841);
nor U3078 (N_3078,N_12,N_82);
or U3079 (N_3079,N_933,N_1111);
or U3080 (N_3080,N_1482,N_2421);
or U3081 (N_3081,N_614,N_2250);
nand U3082 (N_3082,N_369,N_498);
nor U3083 (N_3083,N_1541,N_465);
nor U3084 (N_3084,N_1474,N_1663);
or U3085 (N_3085,N_2216,N_627);
nor U3086 (N_3086,N_1023,N_291);
or U3087 (N_3087,N_570,N_226);
nand U3088 (N_3088,N_1416,N_638);
xor U3089 (N_3089,N_2059,N_2146);
nor U3090 (N_3090,N_370,N_609);
nor U3091 (N_3091,N_46,N_2148);
nor U3092 (N_3092,N_183,N_2109);
nand U3093 (N_3093,N_901,N_2075);
or U3094 (N_3094,N_24,N_2343);
xor U3095 (N_3095,N_1018,N_1132);
and U3096 (N_3096,N_2267,N_1065);
nand U3097 (N_3097,N_138,N_822);
and U3098 (N_3098,N_740,N_2177);
nand U3099 (N_3099,N_566,N_1815);
and U3100 (N_3100,N_11,N_787);
nor U3101 (N_3101,N_1484,N_1862);
or U3102 (N_3102,N_1795,N_943);
xor U3103 (N_3103,N_1411,N_1349);
and U3104 (N_3104,N_72,N_1480);
or U3105 (N_3105,N_182,N_1227);
nand U3106 (N_3106,N_1608,N_450);
xnor U3107 (N_3107,N_1315,N_918);
and U3108 (N_3108,N_642,N_448);
nor U3109 (N_3109,N_1419,N_1941);
and U3110 (N_3110,N_1812,N_1870);
or U3111 (N_3111,N_244,N_1251);
nand U3112 (N_3112,N_1523,N_1629);
nor U3113 (N_3113,N_1015,N_1972);
xnor U3114 (N_3114,N_1937,N_888);
and U3115 (N_3115,N_1471,N_102);
or U3116 (N_3116,N_1138,N_1944);
nand U3117 (N_3117,N_484,N_1174);
and U3118 (N_3118,N_1754,N_2019);
nor U3119 (N_3119,N_196,N_1888);
and U3120 (N_3120,N_2486,N_865);
and U3121 (N_3121,N_1172,N_141);
nand U3122 (N_3122,N_173,N_1771);
nor U3123 (N_3123,N_419,N_651);
or U3124 (N_3124,N_2214,N_2143);
or U3125 (N_3125,N_248,N_1110);
and U3126 (N_3126,N_728,N_2206);
nor U3127 (N_3127,N_386,N_1165);
nand U3128 (N_3128,N_1236,N_2301);
nor U3129 (N_3129,N_6,N_456);
nand U3130 (N_3130,N_297,N_1275);
nor U3131 (N_3131,N_1924,N_229);
and U3132 (N_3132,N_1274,N_2485);
nand U3133 (N_3133,N_813,N_567);
or U3134 (N_3134,N_1563,N_2430);
nand U3135 (N_3135,N_675,N_1929);
nand U3136 (N_3136,N_2467,N_810);
nor U3137 (N_3137,N_1465,N_1396);
xnor U3138 (N_3138,N_1103,N_140);
or U3139 (N_3139,N_1734,N_2158);
and U3140 (N_3140,N_1598,N_1460);
or U3141 (N_3141,N_282,N_716);
nand U3142 (N_3142,N_1520,N_1725);
or U3143 (N_3143,N_2298,N_526);
nor U3144 (N_3144,N_2065,N_676);
or U3145 (N_3145,N_321,N_25);
nand U3146 (N_3146,N_128,N_1099);
or U3147 (N_3147,N_2381,N_1067);
or U3148 (N_3148,N_1802,N_2121);
nor U3149 (N_3149,N_2000,N_3);
nor U3150 (N_3150,N_1576,N_1312);
xnor U3151 (N_3151,N_325,N_1657);
or U3152 (N_3152,N_1990,N_2254);
and U3153 (N_3153,N_476,N_143);
nand U3154 (N_3154,N_605,N_743);
or U3155 (N_3155,N_1938,N_1613);
or U3156 (N_3156,N_2256,N_1250);
or U3157 (N_3157,N_466,N_1086);
nor U3158 (N_3158,N_1040,N_900);
nand U3159 (N_3159,N_4,N_7);
nand U3160 (N_3160,N_1440,N_2353);
or U3161 (N_3161,N_1041,N_2378);
or U3162 (N_3162,N_862,N_2174);
xnor U3163 (N_3163,N_1291,N_1787);
or U3164 (N_3164,N_628,N_1683);
nand U3165 (N_3165,N_2333,N_811);
nor U3166 (N_3166,N_432,N_249);
nand U3167 (N_3167,N_1068,N_1801);
and U3168 (N_3168,N_1105,N_2047);
nand U3169 (N_3169,N_2457,N_1338);
nor U3170 (N_3170,N_1647,N_1009);
nor U3171 (N_3171,N_2255,N_686);
or U3172 (N_3172,N_23,N_1034);
or U3173 (N_3173,N_1077,N_1873);
or U3174 (N_3174,N_1252,N_2282);
nor U3175 (N_3175,N_2213,N_671);
or U3176 (N_3176,N_543,N_980);
nor U3177 (N_3177,N_773,N_997);
or U3178 (N_3178,N_1590,N_1755);
nor U3179 (N_3179,N_1088,N_95);
or U3180 (N_3180,N_315,N_1201);
and U3181 (N_3181,N_654,N_2125);
nand U3182 (N_3182,N_1380,N_596);
or U3183 (N_3183,N_1693,N_1582);
or U3184 (N_3184,N_2245,N_1447);
nor U3185 (N_3185,N_2370,N_5);
or U3186 (N_3186,N_2235,N_1887);
xnor U3187 (N_3187,N_1192,N_2417);
or U3188 (N_3188,N_969,N_2387);
nor U3189 (N_3189,N_1519,N_1120);
xor U3190 (N_3190,N_488,N_2293);
and U3191 (N_3191,N_54,N_1706);
nand U3192 (N_3192,N_396,N_806);
nor U3193 (N_3193,N_2344,N_1808);
and U3194 (N_3194,N_1317,N_2465);
nand U3195 (N_3195,N_511,N_1161);
nor U3196 (N_3196,N_869,N_1369);
or U3197 (N_3197,N_1364,N_2262);
nand U3198 (N_3198,N_85,N_1836);
or U3199 (N_3199,N_1464,N_2300);
or U3200 (N_3200,N_478,N_2132);
nor U3201 (N_3201,N_525,N_2432);
and U3202 (N_3202,N_971,N_1043);
nand U3203 (N_3203,N_665,N_1162);
and U3204 (N_3204,N_1623,N_715);
and U3205 (N_3205,N_750,N_1154);
nand U3206 (N_3206,N_1548,N_221);
and U3207 (N_3207,N_1136,N_1417);
nor U3208 (N_3208,N_1109,N_2193);
nand U3209 (N_3209,N_209,N_1397);
xor U3210 (N_3210,N_1719,N_1318);
or U3211 (N_3211,N_1540,N_2395);
nand U3212 (N_3212,N_1668,N_801);
or U3213 (N_3213,N_214,N_946);
and U3214 (N_3214,N_2470,N_1564);
nand U3215 (N_3215,N_187,N_1428);
xnor U3216 (N_3216,N_390,N_573);
or U3217 (N_3217,N_202,N_1439);
xnor U3218 (N_3218,N_986,N_2303);
nor U3219 (N_3219,N_2183,N_1186);
and U3220 (N_3220,N_689,N_2099);
or U3221 (N_3221,N_669,N_126);
or U3222 (N_3222,N_1658,N_774);
nand U3223 (N_3223,N_168,N_2317);
or U3224 (N_3224,N_1642,N_2468);
xnor U3225 (N_3225,N_1494,N_785);
and U3226 (N_3226,N_1624,N_467);
and U3227 (N_3227,N_1928,N_1985);
and U3228 (N_3228,N_1856,N_1744);
and U3229 (N_3229,N_1267,N_1970);
nor U3230 (N_3230,N_104,N_622);
or U3231 (N_3231,N_2294,N_1107);
nor U3232 (N_3232,N_1210,N_1410);
or U3233 (N_3233,N_745,N_2055);
and U3234 (N_3234,N_351,N_666);
and U3235 (N_3235,N_1316,N_1664);
nand U3236 (N_3236,N_925,N_123);
and U3237 (N_3237,N_1672,N_667);
xnor U3238 (N_3238,N_1881,N_558);
nand U3239 (N_3239,N_1674,N_21);
and U3240 (N_3240,N_485,N_2376);
nand U3241 (N_3241,N_2310,N_1387);
and U3242 (N_3242,N_1125,N_894);
and U3243 (N_3243,N_1995,N_1074);
nand U3244 (N_3244,N_1559,N_401);
nand U3245 (N_3245,N_1319,N_1752);
xnor U3246 (N_3246,N_130,N_2401);
and U3247 (N_3247,N_1606,N_1030);
nand U3248 (N_3248,N_1443,N_1765);
and U3249 (N_3249,N_1131,N_1370);
nand U3250 (N_3250,N_232,N_829);
nand U3251 (N_3251,N_657,N_1922);
nor U3252 (N_3252,N_1389,N_152);
nor U3253 (N_3253,N_1913,N_1189);
or U3254 (N_3254,N_2077,N_2154);
or U3255 (N_3255,N_1778,N_533);
nand U3256 (N_3256,N_2052,N_1751);
nor U3257 (N_3257,N_2336,N_189);
nor U3258 (N_3258,N_741,N_303);
or U3259 (N_3259,N_1588,N_1280);
and U3260 (N_3260,N_157,N_22);
and U3261 (N_3261,N_1255,N_199);
and U3262 (N_3262,N_2186,N_845);
nor U3263 (N_3263,N_89,N_626);
nand U3264 (N_3264,N_2428,N_489);
or U3265 (N_3265,N_973,N_1712);
or U3266 (N_3266,N_451,N_2116);
nand U3267 (N_3267,N_479,N_560);
and U3268 (N_3268,N_17,N_1427);
and U3269 (N_3269,N_800,N_2348);
nand U3270 (N_3270,N_673,N_1357);
nand U3271 (N_3271,N_2334,N_1384);
and U3272 (N_3272,N_1999,N_562);
nand U3273 (N_3273,N_2340,N_1575);
nand U3274 (N_3274,N_763,N_2454);
nor U3275 (N_3275,N_2165,N_1362);
or U3276 (N_3276,N_1260,N_861);
nand U3277 (N_3277,N_204,N_308);
xnor U3278 (N_3278,N_825,N_1444);
or U3279 (N_3279,N_2091,N_418);
nand U3280 (N_3280,N_1759,N_1137);
xnor U3281 (N_3281,N_14,N_1404);
and U3282 (N_3282,N_2307,N_156);
nand U3283 (N_3283,N_2209,N_1653);
nand U3284 (N_3284,N_1360,N_920);
nand U3285 (N_3285,N_171,N_1736);
and U3286 (N_3286,N_1797,N_50);
and U3287 (N_3287,N_1740,N_2203);
or U3288 (N_3288,N_1569,N_970);
or U3289 (N_3289,N_1702,N_70);
nand U3290 (N_3290,N_1835,N_1868);
nand U3291 (N_3291,N_1889,N_1052);
and U3292 (N_3292,N_892,N_1680);
nand U3293 (N_3293,N_474,N_937);
nor U3294 (N_3294,N_1864,N_1779);
nand U3295 (N_3295,N_1453,N_271);
xnor U3296 (N_3296,N_684,N_875);
or U3297 (N_3297,N_224,N_1337);
nor U3298 (N_3298,N_848,N_1254);
and U3299 (N_3299,N_690,N_2443);
nor U3300 (N_3300,N_2139,N_944);
nand U3301 (N_3301,N_1365,N_1741);
nor U3302 (N_3302,N_48,N_2202);
and U3303 (N_3303,N_1219,N_1984);
nand U3304 (N_3304,N_2064,N_2261);
nand U3305 (N_3305,N_2056,N_927);
nand U3306 (N_3306,N_1932,N_1784);
nor U3307 (N_3307,N_380,N_2012);
nand U3308 (N_3308,N_52,N_2046);
or U3309 (N_3309,N_2249,N_681);
nand U3310 (N_3310,N_264,N_1816);
or U3311 (N_3311,N_1093,N_1832);
xnor U3312 (N_3312,N_1953,N_1214);
nor U3313 (N_3313,N_2427,N_174);
nand U3314 (N_3314,N_1522,N_805);
nor U3315 (N_3315,N_127,N_549);
and U3316 (N_3316,N_1565,N_640);
and U3317 (N_3317,N_1980,N_201);
nand U3318 (N_3318,N_977,N_1531);
nand U3319 (N_3319,N_1146,N_270);
nor U3320 (N_3320,N_607,N_1466);
nor U3321 (N_3321,N_57,N_958);
or U3322 (N_3322,N_1732,N_2122);
xnor U3323 (N_3323,N_664,N_340);
nor U3324 (N_3324,N_790,N_1335);
nand U3325 (N_3325,N_1620,N_1655);
and U3326 (N_3326,N_1691,N_1713);
nor U3327 (N_3327,N_1379,N_356);
and U3328 (N_3328,N_814,N_2280);
nand U3329 (N_3329,N_443,N_712);
nor U3330 (N_3330,N_564,N_864);
and U3331 (N_3331,N_1737,N_43);
xor U3332 (N_3332,N_302,N_851);
xor U3333 (N_3333,N_155,N_2275);
and U3334 (N_3334,N_2281,N_1700);
nand U3335 (N_3335,N_1656,N_983);
nor U3336 (N_3336,N_1792,N_603);
and U3337 (N_3337,N_1145,N_1166);
nor U3338 (N_3338,N_623,N_1586);
xnor U3339 (N_3339,N_2315,N_966);
and U3340 (N_3340,N_200,N_2406);
nand U3341 (N_3341,N_134,N_2482);
xnor U3342 (N_3342,N_682,N_1526);
or U3343 (N_3343,N_1845,N_1819);
or U3344 (N_3344,N_926,N_1695);
and U3345 (N_3345,N_846,N_576);
nand U3346 (N_3346,N_1955,N_792);
and U3347 (N_3347,N_2391,N_378);
and U3348 (N_3348,N_327,N_1421);
nand U3349 (N_3349,N_1788,N_709);
or U3350 (N_3350,N_1457,N_1803);
xnor U3351 (N_3351,N_1914,N_516);
nor U3352 (N_3352,N_2105,N_891);
nand U3353 (N_3353,N_29,N_1846);
nor U3354 (N_3354,N_457,N_2201);
nor U3355 (N_3355,N_2259,N_1448);
xor U3356 (N_3356,N_84,N_1607);
and U3357 (N_3357,N_1583,N_1831);
xor U3358 (N_3358,N_2358,N_475);
and U3359 (N_3359,N_83,N_1857);
or U3360 (N_3360,N_702,N_1723);
nand U3361 (N_3361,N_1199,N_1716);
or U3362 (N_3362,N_1378,N_662);
and U3363 (N_3363,N_1028,N_1776);
and U3364 (N_3364,N_1986,N_222);
and U3365 (N_3365,N_1530,N_1727);
nand U3366 (N_3366,N_258,N_260);
nor U3367 (N_3367,N_1076,N_1662);
or U3368 (N_3368,N_1844,N_556);
and U3369 (N_3369,N_618,N_1057);
nand U3370 (N_3370,N_154,N_1390);
nand U3371 (N_3371,N_203,N_1091);
nor U3372 (N_3372,N_2273,N_350);
or U3373 (N_3373,N_782,N_330);
nor U3374 (N_3374,N_452,N_714);
nor U3375 (N_3375,N_610,N_589);
or U3376 (N_3376,N_96,N_1208);
nand U3377 (N_3377,N_841,N_1798);
nand U3378 (N_3378,N_545,N_2170);
and U3379 (N_3379,N_1853,N_299);
nor U3380 (N_3380,N_695,N_1010);
nand U3381 (N_3381,N_496,N_2119);
nor U3382 (N_3382,N_767,N_444);
and U3383 (N_3383,N_540,N_276);
or U3384 (N_3384,N_463,N_1429);
nand U3385 (N_3385,N_0,N_733);
nand U3386 (N_3386,N_2080,N_1259);
and U3387 (N_3387,N_524,N_754);
nand U3388 (N_3388,N_2134,N_1756);
or U3389 (N_3389,N_532,N_181);
and U3390 (N_3390,N_2332,N_1007);
nor U3391 (N_3391,N_2292,N_217);
nor U3392 (N_3392,N_1488,N_2002);
xor U3393 (N_3393,N_629,N_519);
and U3394 (N_3394,N_2497,N_1059);
nor U3395 (N_3395,N_674,N_227);
or U3396 (N_3396,N_2338,N_279);
nand U3397 (N_3397,N_1002,N_190);
xnor U3398 (N_3398,N_1403,N_965);
nand U3399 (N_3399,N_2043,N_345);
or U3400 (N_3400,N_2429,N_296);
and U3401 (N_3401,N_956,N_593);
nor U3402 (N_3402,N_597,N_324);
nand U3403 (N_3403,N_246,N_897);
and U3404 (N_3404,N_1142,N_30);
and U3405 (N_3405,N_1290,N_1309);
or U3406 (N_3406,N_500,N_437);
nand U3407 (N_3407,N_1775,N_2402);
nor U3408 (N_3408,N_1437,N_807);
nor U3409 (N_3409,N_300,N_877);
nand U3410 (N_3410,N_1743,N_2079);
nor U3411 (N_3411,N_2112,N_1829);
nor U3412 (N_3412,N_254,N_342);
or U3413 (N_3413,N_1054,N_1502);
or U3414 (N_3414,N_2481,N_2403);
and U3415 (N_3415,N_688,N_387);
nor U3416 (N_3416,N_2070,N_2459);
and U3417 (N_3417,N_1032,N_108);
and U3418 (N_3418,N_1681,N_2426);
nand U3419 (N_3419,N_305,N_2357);
nand U3420 (N_3420,N_1061,N_2420);
nand U3421 (N_3421,N_793,N_1935);
or U3422 (N_3422,N_583,N_493);
and U3423 (N_3423,N_1116,N_2418);
nor U3424 (N_3424,N_240,N_2461);
nor U3425 (N_3425,N_2081,N_704);
or U3426 (N_3426,N_2195,N_2172);
nor U3427 (N_3427,N_1675,N_66);
nand U3428 (N_3428,N_1292,N_347);
nand U3429 (N_3429,N_581,N_1346);
and U3430 (N_3430,N_1890,N_1062);
or U3431 (N_3431,N_313,N_1393);
nor U3432 (N_3432,N_455,N_796);
or U3433 (N_3433,N_612,N_211);
or U3434 (N_3434,N_2308,N_2393);
or U3435 (N_3435,N_1101,N_1026);
nand U3436 (N_3436,N_1911,N_710);
or U3437 (N_3437,N_2350,N_972);
and U3438 (N_3438,N_453,N_1930);
nor U3439 (N_3439,N_1333,N_2228);
nand U3440 (N_3440,N_2288,N_1899);
nor U3441 (N_3441,N_1572,N_1004);
and U3442 (N_3442,N_1761,N_999);
and U3443 (N_3443,N_1127,N_950);
xor U3444 (N_3444,N_1060,N_2114);
and U3445 (N_3445,N_2404,N_859);
and U3446 (N_3446,N_961,N_111);
or U3447 (N_3447,N_2155,N_1507);
nor U3448 (N_3448,N_166,N_206);
nor U3449 (N_3449,N_775,N_1823);
xnor U3450 (N_3450,N_1394,N_2414);
xor U3451 (N_3451,N_106,N_364);
nand U3452 (N_3452,N_2040,N_58);
and U3453 (N_3453,N_2187,N_554);
nand U3454 (N_3454,N_1083,N_2371);
nand U3455 (N_3455,N_608,N_1542);
xor U3456 (N_3456,N_2222,N_1222);
nand U3457 (N_3457,N_177,N_1580);
nor U3458 (N_3458,N_2274,N_292);
xor U3459 (N_3459,N_1366,N_899);
nor U3460 (N_3460,N_1822,N_59);
xor U3461 (N_3461,N_1097,N_1690);
or U3462 (N_3462,N_1894,N_2054);
nand U3463 (N_3463,N_107,N_624);
nor U3464 (N_3464,N_2364,N_454);
or U3465 (N_3465,N_1954,N_2483);
nor U3466 (N_3466,N_2032,N_1809);
or U3467 (N_3467,N_1514,N_473);
xor U3468 (N_3468,N_637,N_1016);
nand U3469 (N_3469,N_317,N_1828);
nor U3470 (N_3470,N_1549,N_402);
nor U3471 (N_3471,N_1124,N_1278);
nor U3472 (N_3472,N_2207,N_1843);
nor U3473 (N_3473,N_1328,N_1027);
or U3474 (N_3474,N_374,N_416);
nand U3475 (N_3475,N_2003,N_495);
nor U3476 (N_3476,N_1470,N_595);
nand U3477 (N_3477,N_1003,N_535);
and U3478 (N_3478,N_748,N_1006);
and U3479 (N_3479,N_769,N_746);
nand U3480 (N_3480,N_1560,N_274);
nor U3481 (N_3481,N_469,N_1773);
nand U3482 (N_3482,N_542,N_81);
nor U3483 (N_3483,N_1796,N_78);
nand U3484 (N_3484,N_1277,N_910);
nand U3485 (N_3485,N_722,N_2398);
nor U3486 (N_3486,N_1604,N_2367);
and U3487 (N_3487,N_65,N_1698);
nand U3488 (N_3488,N_2257,N_1055);
xnor U3489 (N_3489,N_1570,N_2384);
and U3490 (N_3490,N_766,N_783);
nand U3491 (N_3491,N_1697,N_2108);
or U3492 (N_3492,N_2413,N_1886);
nand U3493 (N_3493,N_2129,N_148);
xor U3494 (N_3494,N_389,N_239);
or U3495 (N_3495,N_2044,N_2425);
and U3496 (N_3496,N_2368,N_283);
xnor U3497 (N_3497,N_250,N_529);
nor U3498 (N_3498,N_1405,N_863);
nor U3499 (N_3499,N_1268,N_88);
xor U3500 (N_3500,N_2151,N_215);
nand U3501 (N_3501,N_1867,N_2316);
nor U3502 (N_3502,N_44,N_1840);
and U3503 (N_3503,N_938,N_831);
nor U3504 (N_3504,N_1619,N_1150);
nand U3505 (N_3505,N_2182,N_1510);
nand U3506 (N_3506,N_592,N_2477);
nand U3507 (N_3507,N_879,N_289);
or U3508 (N_3508,N_771,N_2045);
and U3509 (N_3509,N_857,N_1554);
nand U3510 (N_3510,N_514,N_911);
or U3511 (N_3511,N_2197,N_1981);
or U3512 (N_3512,N_376,N_2345);
nand U3513 (N_3513,N_1609,N_483);
nand U3514 (N_3514,N_653,N_935);
nor U3515 (N_3515,N_616,N_1463);
and U3516 (N_3516,N_2322,N_74);
nor U3517 (N_3517,N_707,N_2212);
and U3518 (N_3518,N_1659,N_2478);
and U3519 (N_3519,N_2379,N_1847);
or U3520 (N_3520,N_1056,N_679);
nor U3521 (N_3521,N_580,N_1121);
or U3522 (N_3522,N_1533,N_2208);
nand U3523 (N_3523,N_2484,N_2220);
and U3524 (N_3524,N_2385,N_2225);
xnor U3525 (N_3525,N_1381,N_1264);
and U3526 (N_3526,N_991,N_1321);
nor U3527 (N_3527,N_1799,N_2005);
nor U3528 (N_3528,N_2460,N_2127);
nor U3529 (N_3529,N_819,N_1686);
xor U3530 (N_3530,N_1021,N_2242);
and U3531 (N_3531,N_151,N_1031);
xor U3532 (N_3532,N_2445,N_1300);
nor U3533 (N_3533,N_2283,N_1135);
and U3534 (N_3534,N_379,N_1555);
xnor U3535 (N_3535,N_873,N_1912);
nand U3536 (N_3536,N_1793,N_1412);
and U3537 (N_3537,N_1794,N_1733);
or U3538 (N_3538,N_1035,N_1478);
or U3539 (N_3539,N_2150,N_257);
nor U3540 (N_3540,N_1593,N_2178);
nor U3541 (N_3541,N_1184,N_648);
nand U3542 (N_3542,N_255,N_442);
nand U3543 (N_3543,N_94,N_472);
nor U3544 (N_3544,N_328,N_1237);
nand U3545 (N_3545,N_2494,N_1511);
or U3546 (N_3546,N_1708,N_420);
nand U3547 (N_3547,N_2,N_677);
and U3548 (N_3548,N_417,N_761);
nand U3549 (N_3549,N_601,N_400);
nor U3550 (N_3550,N_1096,N_1544);
or U3551 (N_3551,N_2227,N_1851);
nand U3552 (N_3552,N_1968,N_1171);
or U3553 (N_3553,N_2111,N_575);
nor U3554 (N_3554,N_408,N_1232);
and U3555 (N_3555,N_477,N_1046);
nand U3556 (N_3556,N_697,N_912);
and U3557 (N_3557,N_1477,N_788);
or U3558 (N_3558,N_19,N_1965);
and U3559 (N_3559,N_737,N_808);
nor U3560 (N_3560,N_1849,N_241);
xnor U3561 (N_3561,N_1359,N_1297);
nand U3562 (N_3562,N_874,N_1997);
or U3563 (N_3563,N_1000,N_1988);
nand U3564 (N_3564,N_284,N_1807);
nor U3565 (N_3565,N_2090,N_852);
nor U3566 (N_3566,N_2013,N_468);
and U3567 (N_3567,N_1468,N_1180);
xor U3568 (N_3568,N_1701,N_67);
nor U3569 (N_3569,N_2071,N_2058);
nor U3570 (N_3570,N_1962,N_2087);
nor U3571 (N_3571,N_1382,N_1395);
nor U3572 (N_3572,N_1113,N_568);
nand U3573 (N_3573,N_1169,N_281);
or U3574 (N_3574,N_1296,N_1960);
nand U3575 (N_3575,N_491,N_2327);
nor U3576 (N_3576,N_923,N_620);
nor U3577 (N_3577,N_2412,N_1827);
and U3578 (N_3578,N_1398,N_1128);
nand U3579 (N_3579,N_2016,N_2031);
and U3580 (N_3580,N_870,N_2123);
or U3581 (N_3581,N_572,N_2279);
nor U3582 (N_3582,N_2269,N_38);
xnor U3583 (N_3583,N_764,N_1258);
nand U3584 (N_3584,N_1159,N_2015);
and U3585 (N_3585,N_1896,N_1487);
and U3586 (N_3586,N_267,N_1571);
nand U3587 (N_3587,N_1824,N_2189);
nor U3588 (N_3588,N_1946,N_2029);
or U3589 (N_3589,N_118,N_1687);
and U3590 (N_3590,N_2423,N_1182);
xor U3591 (N_3591,N_1498,N_1263);
nand U3592 (N_3592,N_1959,N_1679);
nor U3593 (N_3593,N_1203,N_2389);
xnor U3594 (N_3594,N_103,N_1901);
nand U3595 (N_3595,N_1305,N_1005);
and U3596 (N_3596,N_1343,N_898);
nor U3597 (N_3597,N_39,N_458);
and U3598 (N_3598,N_439,N_259);
nor U3599 (N_3599,N_2311,N_835);
nand U3600 (N_3600,N_135,N_1081);
or U3601 (N_3601,N_931,N_2021);
nand U3602 (N_3602,N_1226,N_470);
nand U3603 (N_3603,N_621,N_1206);
nor U3604 (N_3604,N_26,N_2399);
nand U3605 (N_3605,N_1900,N_2028);
nor U3606 (N_3606,N_462,N_2474);
and U3607 (N_3607,N_2181,N_1413);
nor U3608 (N_3608,N_150,N_285);
or U3609 (N_3609,N_929,N_1307);
xor U3610 (N_3610,N_2437,N_1670);
and U3611 (N_3611,N_1045,N_1352);
and U3612 (N_3612,N_2009,N_1191);
or U3613 (N_3613,N_441,N_1153);
or U3614 (N_3614,N_310,N_1499);
xor U3615 (N_3615,N_692,N_952);
or U3616 (N_3616,N_951,N_663);
or U3617 (N_3617,N_2159,N_889);
nand U3618 (N_3618,N_1152,N_2217);
or U3619 (N_3619,N_2157,N_139);
xnor U3620 (N_3620,N_1652,N_1308);
nor U3621 (N_3621,N_513,N_1633);
xnor U3622 (N_3622,N_1048,N_1418);
nor U3623 (N_3623,N_2089,N_1561);
nor U3624 (N_3624,N_1599,N_1534);
nor U3625 (N_3625,N_1958,N_721);
or U3626 (N_3626,N_1804,N_1436);
or U3627 (N_3627,N_1707,N_2488);
nand U3628 (N_3628,N_9,N_1770);
nor U3629 (N_3629,N_2444,N_1949);
nand U3630 (N_3630,N_2455,N_449);
nor U3631 (N_3631,N_425,N_332);
and U3632 (N_3632,N_2198,N_233);
and U3633 (N_3633,N_1916,N_1114);
nor U3634 (N_3634,N_1501,N_172);
nand U3635 (N_3635,N_842,N_1198);
xor U3636 (N_3636,N_1243,N_2495);
and U3637 (N_3637,N_159,N_2247);
and U3638 (N_3638,N_2330,N_744);
nor U3639 (N_3639,N_2093,N_1235);
nor U3640 (N_3640,N_2219,N_1298);
or U3641 (N_3641,N_1906,N_2339);
and U3642 (N_3642,N_2489,N_683);
nand U3643 (N_3643,N_998,N_1786);
and U3644 (N_3644,N_1584,N_1650);
or U3645 (N_3645,N_1638,N_1388);
and U3646 (N_3646,N_812,N_2050);
or U3647 (N_3647,N_1353,N_837);
or U3648 (N_3648,N_459,N_2066);
or U3649 (N_3649,N_1024,N_1818);
and U3650 (N_3650,N_2422,N_2233);
or U3651 (N_3651,N_377,N_1014);
and U3652 (N_3652,N_2448,N_2473);
nand U3653 (N_3653,N_1038,N_770);
and U3654 (N_3654,N_45,N_2188);
nor U3655 (N_3655,N_1287,N_1272);
and U3656 (N_3656,N_611,N_2196);
nor U3657 (N_3657,N_1144,N_438);
nor U3658 (N_3658,N_2035,N_353);
nand U3659 (N_3659,N_1745,N_1766);
or U3660 (N_3660,N_1964,N_2319);
nor U3661 (N_3661,N_1391,N_2424);
nor U3662 (N_3662,N_1435,N_2167);
or U3663 (N_3663,N_2204,N_1603);
nand U3664 (N_3664,N_1897,N_1711);
and U3665 (N_3665,N_149,N_1893);
and U3666 (N_3666,N_655,N_341);
and U3667 (N_3667,N_35,N_921);
and U3668 (N_3668,N_1234,N_2069);
nor U3669 (N_3669,N_974,N_1830);
or U3670 (N_3670,N_1402,N_2039);
nand U3671 (N_3671,N_1233,N_934);
xor U3672 (N_3672,N_269,N_2331);
and U3673 (N_3673,N_1611,N_1176);
and U3674 (N_3674,N_220,N_724);
and U3675 (N_3675,N_2120,N_1936);
nor U3676 (N_3676,N_2405,N_587);
nand U3677 (N_3677,N_1940,N_1019);
nand U3678 (N_3678,N_2117,N_916);
nor U3679 (N_3679,N_2025,N_1957);
nand U3680 (N_3680,N_1066,N_114);
or U3681 (N_3681,N_826,N_534);
nand U3682 (N_3682,N_537,N_1956);
nand U3683 (N_3683,N_1012,N_2328);
or U3684 (N_3684,N_1601,N_1497);
xnor U3685 (N_3685,N_2211,N_1450);
nor U3686 (N_3686,N_218,N_357);
nor U3687 (N_3687,N_2037,N_331);
and U3688 (N_3688,N_2271,N_1919);
and U3689 (N_3689,N_1717,N_551);
nand U3690 (N_3690,N_881,N_2022);
nand U3691 (N_3691,N_144,N_2314);
nand U3692 (N_3692,N_49,N_2438);
nand U3693 (N_3693,N_2018,N_772);
or U3694 (N_3694,N_1392,N_507);
or U3695 (N_3695,N_1119,N_1185);
or U3696 (N_3696,N_1969,N_1581);
nor U3697 (N_3697,N_1865,N_1069);
nand U3698 (N_3698,N_915,N_1070);
nand U3699 (N_3699,N_92,N_1626);
nor U3700 (N_3700,N_2103,N_816);
and U3701 (N_3701,N_1600,N_1579);
nand U3702 (N_3702,N_2323,N_2416);
nand U3703 (N_3703,N_117,N_367);
nand U3704 (N_3704,N_503,N_1556);
nand U3705 (N_3705,N_2272,N_2374);
or U3706 (N_3706,N_1098,N_314);
or U3707 (N_3707,N_1211,N_711);
or U3708 (N_3708,N_2175,N_1438);
nand U3709 (N_3709,N_522,N_2450);
nor U3710 (N_3710,N_1495,N_2006);
nand U3711 (N_3711,N_866,N_1622);
xor U3712 (N_3712,N_1789,N_1696);
or U3713 (N_3713,N_2107,N_184);
or U3714 (N_3714,N_2325,N_1880);
or U3715 (N_3715,N_1075,N_1673);
xnor U3716 (N_3716,N_995,N_2446);
nor U3717 (N_3717,N_1449,N_1923);
and U3718 (N_3718,N_2347,N_1454);
nand U3719 (N_3719,N_780,N_2010);
nor U3720 (N_3720,N_2313,N_639);
nand U3721 (N_3721,N_1080,N_615);
nand U3722 (N_3722,N_508,N_1348);
nor U3723 (N_3723,N_1528,N_480);
or U3724 (N_3724,N_2441,N_2038);
and U3725 (N_3725,N_599,N_2318);
or U3726 (N_3726,N_431,N_850);
and U3727 (N_3727,N_2419,N_2394);
and U3728 (N_3728,N_125,N_2051);
nor U3729 (N_3729,N_1863,N_1140);
or U3730 (N_3730,N_56,N_2442);
or U3731 (N_3731,N_1907,N_887);
or U3732 (N_3732,N_752,N_1050);
xnor U3733 (N_3733,N_1677,N_1313);
and U3734 (N_3734,N_167,N_1764);
nor U3735 (N_3735,N_344,N_165);
and U3736 (N_3736,N_435,N_2011);
xnor U3737 (N_3737,N_1918,N_518);
or U3738 (N_3738,N_838,N_120);
nand U3739 (N_3739,N_8,N_2285);
nand U3740 (N_3740,N_1780,N_1757);
nand U3741 (N_3741,N_406,N_1920);
and U3742 (N_3742,N_1927,N_821);
or U3743 (N_3743,N_691,N_2061);
and U3744 (N_3744,N_2408,N_649);
or U3745 (N_3745,N_1451,N_602);
and U3746 (N_3746,N_1961,N_427);
nor U3747 (N_3747,N_510,N_1078);
xnor U3748 (N_3748,N_1179,N_2126);
nand U3749 (N_3749,N_2487,N_1948);
and U3750 (N_3750,N_1715,N_1433);
or U3751 (N_3751,N_780,N_2241);
nor U3752 (N_3752,N_1478,N_1200);
and U3753 (N_3753,N_1983,N_688);
nor U3754 (N_3754,N_204,N_2225);
or U3755 (N_3755,N_607,N_411);
or U3756 (N_3756,N_799,N_274);
nor U3757 (N_3757,N_2255,N_1355);
nor U3758 (N_3758,N_1152,N_1151);
nand U3759 (N_3759,N_2415,N_1679);
and U3760 (N_3760,N_1122,N_286);
and U3761 (N_3761,N_845,N_2027);
xnor U3762 (N_3762,N_1657,N_406);
or U3763 (N_3763,N_328,N_368);
and U3764 (N_3764,N_386,N_2475);
and U3765 (N_3765,N_1226,N_738);
or U3766 (N_3766,N_1043,N_1388);
or U3767 (N_3767,N_561,N_111);
xnor U3768 (N_3768,N_2461,N_768);
or U3769 (N_3769,N_1148,N_1579);
or U3770 (N_3770,N_454,N_1154);
and U3771 (N_3771,N_1494,N_1769);
or U3772 (N_3772,N_1300,N_70);
and U3773 (N_3773,N_2159,N_1649);
nor U3774 (N_3774,N_1548,N_1593);
xnor U3775 (N_3775,N_1338,N_2020);
nand U3776 (N_3776,N_2366,N_1105);
nor U3777 (N_3777,N_2165,N_2093);
or U3778 (N_3778,N_563,N_1324);
nand U3779 (N_3779,N_1661,N_1238);
nor U3780 (N_3780,N_2338,N_644);
or U3781 (N_3781,N_1315,N_2297);
nand U3782 (N_3782,N_336,N_2154);
nor U3783 (N_3783,N_1312,N_2136);
xor U3784 (N_3784,N_2241,N_822);
and U3785 (N_3785,N_109,N_1241);
nand U3786 (N_3786,N_272,N_2362);
nor U3787 (N_3787,N_118,N_1538);
nor U3788 (N_3788,N_1618,N_914);
xor U3789 (N_3789,N_312,N_1792);
or U3790 (N_3790,N_2207,N_852);
and U3791 (N_3791,N_520,N_689);
and U3792 (N_3792,N_652,N_411);
and U3793 (N_3793,N_2154,N_180);
or U3794 (N_3794,N_1148,N_1516);
nor U3795 (N_3795,N_224,N_2270);
xnor U3796 (N_3796,N_1025,N_1708);
xnor U3797 (N_3797,N_1093,N_2283);
or U3798 (N_3798,N_1934,N_2150);
nand U3799 (N_3799,N_2169,N_1402);
or U3800 (N_3800,N_1621,N_824);
or U3801 (N_3801,N_2383,N_1272);
nor U3802 (N_3802,N_775,N_889);
or U3803 (N_3803,N_493,N_1308);
nand U3804 (N_3804,N_1169,N_843);
or U3805 (N_3805,N_177,N_1675);
and U3806 (N_3806,N_363,N_274);
nand U3807 (N_3807,N_839,N_2144);
nor U3808 (N_3808,N_2496,N_1880);
or U3809 (N_3809,N_2318,N_2013);
xor U3810 (N_3810,N_1680,N_1895);
nand U3811 (N_3811,N_1346,N_2070);
nand U3812 (N_3812,N_1995,N_2313);
and U3813 (N_3813,N_599,N_450);
nor U3814 (N_3814,N_1762,N_663);
nor U3815 (N_3815,N_1337,N_1726);
or U3816 (N_3816,N_2024,N_1937);
nor U3817 (N_3817,N_2070,N_1252);
nor U3818 (N_3818,N_604,N_1966);
nor U3819 (N_3819,N_1287,N_840);
and U3820 (N_3820,N_732,N_2023);
or U3821 (N_3821,N_920,N_1379);
or U3822 (N_3822,N_1984,N_1708);
and U3823 (N_3823,N_332,N_643);
and U3824 (N_3824,N_591,N_53);
nand U3825 (N_3825,N_2161,N_2364);
nor U3826 (N_3826,N_10,N_1886);
nand U3827 (N_3827,N_2025,N_1343);
and U3828 (N_3828,N_443,N_425);
xnor U3829 (N_3829,N_2112,N_1990);
or U3830 (N_3830,N_1520,N_2303);
or U3831 (N_3831,N_867,N_1947);
nor U3832 (N_3832,N_1971,N_804);
and U3833 (N_3833,N_1100,N_1232);
nor U3834 (N_3834,N_2497,N_81);
and U3835 (N_3835,N_2034,N_1462);
nand U3836 (N_3836,N_1884,N_1351);
nand U3837 (N_3837,N_1785,N_681);
and U3838 (N_3838,N_2385,N_1250);
nand U3839 (N_3839,N_377,N_356);
or U3840 (N_3840,N_2313,N_668);
or U3841 (N_3841,N_855,N_1169);
nor U3842 (N_3842,N_302,N_121);
nor U3843 (N_3843,N_1578,N_653);
nor U3844 (N_3844,N_2460,N_22);
nor U3845 (N_3845,N_2244,N_93);
or U3846 (N_3846,N_1627,N_811);
nand U3847 (N_3847,N_1400,N_1903);
or U3848 (N_3848,N_2432,N_1611);
and U3849 (N_3849,N_628,N_1573);
xnor U3850 (N_3850,N_625,N_204);
and U3851 (N_3851,N_1843,N_645);
nand U3852 (N_3852,N_1211,N_2336);
or U3853 (N_3853,N_1861,N_1770);
nand U3854 (N_3854,N_340,N_812);
nand U3855 (N_3855,N_1157,N_1821);
nand U3856 (N_3856,N_1447,N_198);
nor U3857 (N_3857,N_702,N_887);
and U3858 (N_3858,N_1126,N_1751);
and U3859 (N_3859,N_565,N_1454);
nand U3860 (N_3860,N_809,N_318);
nand U3861 (N_3861,N_1210,N_890);
nand U3862 (N_3862,N_1177,N_100);
xor U3863 (N_3863,N_965,N_2037);
nand U3864 (N_3864,N_887,N_1979);
or U3865 (N_3865,N_752,N_154);
and U3866 (N_3866,N_2103,N_1923);
or U3867 (N_3867,N_588,N_163);
nor U3868 (N_3868,N_2489,N_1134);
nand U3869 (N_3869,N_763,N_1802);
nand U3870 (N_3870,N_629,N_1043);
nor U3871 (N_3871,N_1355,N_2261);
and U3872 (N_3872,N_2288,N_11);
xnor U3873 (N_3873,N_1959,N_912);
and U3874 (N_3874,N_522,N_1073);
or U3875 (N_3875,N_730,N_1889);
xnor U3876 (N_3876,N_1636,N_395);
nor U3877 (N_3877,N_948,N_840);
nor U3878 (N_3878,N_365,N_1558);
nand U3879 (N_3879,N_2010,N_971);
nand U3880 (N_3880,N_87,N_2384);
xnor U3881 (N_3881,N_1977,N_1810);
or U3882 (N_3882,N_1138,N_1981);
nand U3883 (N_3883,N_1736,N_574);
or U3884 (N_3884,N_1223,N_808);
or U3885 (N_3885,N_1504,N_867);
or U3886 (N_3886,N_1684,N_2153);
nor U3887 (N_3887,N_1587,N_949);
and U3888 (N_3888,N_2151,N_743);
nor U3889 (N_3889,N_739,N_1205);
nand U3890 (N_3890,N_276,N_1043);
and U3891 (N_3891,N_597,N_786);
nor U3892 (N_3892,N_2100,N_1925);
nor U3893 (N_3893,N_63,N_1255);
nand U3894 (N_3894,N_1481,N_2482);
nor U3895 (N_3895,N_1820,N_1413);
or U3896 (N_3896,N_949,N_425);
and U3897 (N_3897,N_1279,N_412);
or U3898 (N_3898,N_1410,N_585);
nand U3899 (N_3899,N_1994,N_1236);
nand U3900 (N_3900,N_302,N_1849);
nor U3901 (N_3901,N_1229,N_642);
xor U3902 (N_3902,N_466,N_41);
and U3903 (N_3903,N_2195,N_1086);
nor U3904 (N_3904,N_197,N_2053);
nor U3905 (N_3905,N_2327,N_1728);
nand U3906 (N_3906,N_2027,N_1077);
and U3907 (N_3907,N_2400,N_1562);
nand U3908 (N_3908,N_2059,N_936);
nor U3909 (N_3909,N_1975,N_104);
and U3910 (N_3910,N_1892,N_1001);
nand U3911 (N_3911,N_880,N_611);
nor U3912 (N_3912,N_2316,N_1722);
nor U3913 (N_3913,N_675,N_739);
and U3914 (N_3914,N_960,N_1658);
and U3915 (N_3915,N_2148,N_263);
nand U3916 (N_3916,N_433,N_117);
xor U3917 (N_3917,N_1836,N_220);
and U3918 (N_3918,N_974,N_1374);
nor U3919 (N_3919,N_932,N_1898);
or U3920 (N_3920,N_178,N_625);
and U3921 (N_3921,N_1398,N_1362);
and U3922 (N_3922,N_775,N_509);
and U3923 (N_3923,N_1947,N_1543);
nor U3924 (N_3924,N_583,N_2479);
nor U3925 (N_3925,N_1407,N_1192);
or U3926 (N_3926,N_1306,N_1776);
nand U3927 (N_3927,N_1317,N_1768);
or U3928 (N_3928,N_1542,N_1236);
nand U3929 (N_3929,N_1915,N_562);
nand U3930 (N_3930,N_1574,N_1165);
xnor U3931 (N_3931,N_1360,N_1343);
or U3932 (N_3932,N_1539,N_2117);
nand U3933 (N_3933,N_1529,N_1281);
nand U3934 (N_3934,N_909,N_539);
or U3935 (N_3935,N_794,N_818);
or U3936 (N_3936,N_2011,N_616);
nand U3937 (N_3937,N_2188,N_1130);
xor U3938 (N_3938,N_1196,N_778);
nand U3939 (N_3939,N_949,N_1677);
xnor U3940 (N_3940,N_1174,N_2125);
or U3941 (N_3941,N_255,N_145);
xor U3942 (N_3942,N_1023,N_1429);
xnor U3943 (N_3943,N_2051,N_1760);
xnor U3944 (N_3944,N_1525,N_193);
nor U3945 (N_3945,N_198,N_1208);
or U3946 (N_3946,N_195,N_1516);
nand U3947 (N_3947,N_265,N_1663);
nand U3948 (N_3948,N_600,N_2167);
or U3949 (N_3949,N_1835,N_1189);
or U3950 (N_3950,N_2187,N_331);
nor U3951 (N_3951,N_1954,N_534);
and U3952 (N_3952,N_923,N_499);
xor U3953 (N_3953,N_2250,N_1238);
nor U3954 (N_3954,N_1534,N_1942);
nor U3955 (N_3955,N_1537,N_23);
or U3956 (N_3956,N_1753,N_1472);
nor U3957 (N_3957,N_2436,N_1445);
nor U3958 (N_3958,N_2472,N_1724);
xnor U3959 (N_3959,N_571,N_992);
nand U3960 (N_3960,N_726,N_1545);
nand U3961 (N_3961,N_1846,N_1592);
nor U3962 (N_3962,N_955,N_1482);
or U3963 (N_3963,N_1566,N_918);
nor U3964 (N_3964,N_995,N_845);
nor U3965 (N_3965,N_1242,N_955);
nand U3966 (N_3966,N_1764,N_377);
and U3967 (N_3967,N_1720,N_802);
and U3968 (N_3968,N_2312,N_435);
or U3969 (N_3969,N_91,N_2144);
nor U3970 (N_3970,N_2143,N_1266);
nor U3971 (N_3971,N_2445,N_1576);
nand U3972 (N_3972,N_1686,N_60);
and U3973 (N_3973,N_204,N_884);
nand U3974 (N_3974,N_1890,N_316);
or U3975 (N_3975,N_1762,N_850);
nor U3976 (N_3976,N_715,N_856);
or U3977 (N_3977,N_572,N_1048);
xor U3978 (N_3978,N_2155,N_2167);
and U3979 (N_3979,N_2074,N_1438);
nor U3980 (N_3980,N_728,N_2043);
nand U3981 (N_3981,N_767,N_2104);
or U3982 (N_3982,N_1226,N_342);
or U3983 (N_3983,N_1263,N_1097);
nand U3984 (N_3984,N_2400,N_680);
or U3985 (N_3985,N_526,N_274);
and U3986 (N_3986,N_663,N_2446);
and U3987 (N_3987,N_211,N_2493);
nor U3988 (N_3988,N_713,N_766);
and U3989 (N_3989,N_1670,N_309);
xnor U3990 (N_3990,N_2243,N_1928);
or U3991 (N_3991,N_1584,N_1589);
xor U3992 (N_3992,N_602,N_1628);
nor U3993 (N_3993,N_1971,N_982);
and U3994 (N_3994,N_463,N_2190);
nand U3995 (N_3995,N_282,N_2389);
nor U3996 (N_3996,N_284,N_1346);
nor U3997 (N_3997,N_2394,N_810);
or U3998 (N_3998,N_2107,N_2095);
nand U3999 (N_3999,N_120,N_390);
or U4000 (N_4000,N_2033,N_43);
or U4001 (N_4001,N_2407,N_369);
nand U4002 (N_4002,N_1105,N_313);
or U4003 (N_4003,N_212,N_567);
or U4004 (N_4004,N_1432,N_285);
nand U4005 (N_4005,N_716,N_343);
and U4006 (N_4006,N_1485,N_161);
nand U4007 (N_4007,N_2292,N_503);
nor U4008 (N_4008,N_226,N_869);
xor U4009 (N_4009,N_201,N_1661);
nor U4010 (N_4010,N_2001,N_1697);
nor U4011 (N_4011,N_420,N_1970);
or U4012 (N_4012,N_2364,N_471);
xnor U4013 (N_4013,N_503,N_978);
nand U4014 (N_4014,N_600,N_1199);
or U4015 (N_4015,N_954,N_1951);
or U4016 (N_4016,N_1246,N_374);
or U4017 (N_4017,N_1145,N_1542);
nor U4018 (N_4018,N_1563,N_1135);
or U4019 (N_4019,N_1430,N_89);
and U4020 (N_4020,N_776,N_1226);
nor U4021 (N_4021,N_1214,N_1521);
or U4022 (N_4022,N_902,N_157);
nor U4023 (N_4023,N_934,N_2473);
nor U4024 (N_4024,N_968,N_1234);
or U4025 (N_4025,N_1513,N_1816);
nand U4026 (N_4026,N_1415,N_520);
and U4027 (N_4027,N_1860,N_1279);
nand U4028 (N_4028,N_2225,N_1391);
or U4029 (N_4029,N_680,N_1046);
and U4030 (N_4030,N_2136,N_1065);
and U4031 (N_4031,N_72,N_638);
nor U4032 (N_4032,N_565,N_1943);
and U4033 (N_4033,N_527,N_2220);
nand U4034 (N_4034,N_1981,N_934);
or U4035 (N_4035,N_1724,N_1234);
or U4036 (N_4036,N_339,N_299);
and U4037 (N_4037,N_2408,N_501);
and U4038 (N_4038,N_796,N_1733);
and U4039 (N_4039,N_502,N_1903);
nand U4040 (N_4040,N_2449,N_2411);
or U4041 (N_4041,N_102,N_493);
xnor U4042 (N_4042,N_1436,N_846);
nand U4043 (N_4043,N_1465,N_2144);
and U4044 (N_4044,N_252,N_341);
and U4045 (N_4045,N_235,N_1062);
nor U4046 (N_4046,N_1110,N_659);
nand U4047 (N_4047,N_1674,N_1720);
or U4048 (N_4048,N_1188,N_1893);
or U4049 (N_4049,N_1134,N_503);
nand U4050 (N_4050,N_2029,N_147);
xnor U4051 (N_4051,N_1520,N_1976);
or U4052 (N_4052,N_1319,N_1812);
and U4053 (N_4053,N_1742,N_2261);
and U4054 (N_4054,N_980,N_2109);
nor U4055 (N_4055,N_1699,N_2178);
nor U4056 (N_4056,N_1809,N_1139);
nor U4057 (N_4057,N_530,N_1804);
or U4058 (N_4058,N_1235,N_734);
or U4059 (N_4059,N_2004,N_904);
xor U4060 (N_4060,N_1717,N_2115);
and U4061 (N_4061,N_591,N_799);
xor U4062 (N_4062,N_2091,N_1892);
and U4063 (N_4063,N_278,N_888);
nand U4064 (N_4064,N_602,N_481);
and U4065 (N_4065,N_2495,N_2039);
nand U4066 (N_4066,N_277,N_1308);
nor U4067 (N_4067,N_1801,N_1237);
nand U4068 (N_4068,N_858,N_2449);
nand U4069 (N_4069,N_1276,N_2359);
and U4070 (N_4070,N_1604,N_957);
nand U4071 (N_4071,N_2491,N_922);
nor U4072 (N_4072,N_1580,N_1135);
xnor U4073 (N_4073,N_1720,N_2175);
nand U4074 (N_4074,N_965,N_712);
or U4075 (N_4075,N_1128,N_1555);
and U4076 (N_4076,N_2339,N_571);
and U4077 (N_4077,N_70,N_58);
or U4078 (N_4078,N_834,N_2315);
nand U4079 (N_4079,N_1411,N_1192);
nor U4080 (N_4080,N_1665,N_731);
or U4081 (N_4081,N_1564,N_2112);
or U4082 (N_4082,N_530,N_203);
nand U4083 (N_4083,N_330,N_2341);
and U4084 (N_4084,N_1860,N_1705);
and U4085 (N_4085,N_275,N_30);
nor U4086 (N_4086,N_1317,N_559);
and U4087 (N_4087,N_1655,N_1718);
xor U4088 (N_4088,N_1986,N_748);
or U4089 (N_4089,N_1078,N_517);
nand U4090 (N_4090,N_1042,N_423);
nor U4091 (N_4091,N_2469,N_2063);
xor U4092 (N_4092,N_500,N_2484);
and U4093 (N_4093,N_2184,N_1519);
and U4094 (N_4094,N_1120,N_432);
xor U4095 (N_4095,N_1345,N_649);
nor U4096 (N_4096,N_1414,N_846);
nor U4097 (N_4097,N_1003,N_1379);
and U4098 (N_4098,N_554,N_1538);
or U4099 (N_4099,N_1859,N_357);
and U4100 (N_4100,N_1632,N_1323);
nand U4101 (N_4101,N_756,N_1613);
nand U4102 (N_4102,N_518,N_390);
nor U4103 (N_4103,N_2019,N_2269);
or U4104 (N_4104,N_2290,N_54);
and U4105 (N_4105,N_11,N_2153);
or U4106 (N_4106,N_140,N_910);
nand U4107 (N_4107,N_1128,N_1000);
or U4108 (N_4108,N_88,N_24);
xor U4109 (N_4109,N_2020,N_1213);
nor U4110 (N_4110,N_1147,N_1636);
nor U4111 (N_4111,N_436,N_1585);
nor U4112 (N_4112,N_2210,N_37);
nand U4113 (N_4113,N_2126,N_1975);
or U4114 (N_4114,N_1405,N_460);
nand U4115 (N_4115,N_1319,N_1326);
and U4116 (N_4116,N_581,N_647);
and U4117 (N_4117,N_1910,N_321);
or U4118 (N_4118,N_640,N_2238);
nor U4119 (N_4119,N_771,N_1945);
and U4120 (N_4120,N_1972,N_1780);
nor U4121 (N_4121,N_1011,N_2282);
nor U4122 (N_4122,N_1883,N_1013);
xnor U4123 (N_4123,N_2462,N_146);
or U4124 (N_4124,N_2340,N_1452);
xnor U4125 (N_4125,N_984,N_99);
nor U4126 (N_4126,N_1511,N_989);
or U4127 (N_4127,N_1722,N_1346);
xnor U4128 (N_4128,N_2380,N_1476);
and U4129 (N_4129,N_89,N_880);
or U4130 (N_4130,N_615,N_1672);
nand U4131 (N_4131,N_1288,N_2219);
or U4132 (N_4132,N_1179,N_1983);
nand U4133 (N_4133,N_829,N_2424);
nand U4134 (N_4134,N_1439,N_524);
or U4135 (N_4135,N_1779,N_968);
nor U4136 (N_4136,N_1128,N_1947);
and U4137 (N_4137,N_748,N_905);
nor U4138 (N_4138,N_2190,N_1561);
nor U4139 (N_4139,N_1029,N_1506);
nor U4140 (N_4140,N_1833,N_1731);
and U4141 (N_4141,N_370,N_1782);
nor U4142 (N_4142,N_489,N_600);
nor U4143 (N_4143,N_936,N_1509);
nand U4144 (N_4144,N_2,N_2389);
nor U4145 (N_4145,N_498,N_2023);
and U4146 (N_4146,N_29,N_1417);
and U4147 (N_4147,N_2380,N_1812);
nor U4148 (N_4148,N_711,N_2340);
nor U4149 (N_4149,N_1793,N_210);
or U4150 (N_4150,N_2237,N_1417);
nand U4151 (N_4151,N_1272,N_1455);
nor U4152 (N_4152,N_2306,N_1258);
nor U4153 (N_4153,N_722,N_2058);
xor U4154 (N_4154,N_425,N_1513);
and U4155 (N_4155,N_430,N_1202);
nand U4156 (N_4156,N_158,N_1665);
and U4157 (N_4157,N_2284,N_852);
nand U4158 (N_4158,N_996,N_1183);
or U4159 (N_4159,N_4,N_2136);
xnor U4160 (N_4160,N_1782,N_2306);
or U4161 (N_4161,N_1061,N_260);
nand U4162 (N_4162,N_1161,N_2116);
nor U4163 (N_4163,N_837,N_708);
and U4164 (N_4164,N_820,N_1173);
nand U4165 (N_4165,N_1454,N_165);
xor U4166 (N_4166,N_69,N_719);
and U4167 (N_4167,N_2071,N_2415);
nand U4168 (N_4168,N_462,N_573);
nor U4169 (N_4169,N_890,N_2334);
nor U4170 (N_4170,N_437,N_825);
nor U4171 (N_4171,N_1153,N_261);
nor U4172 (N_4172,N_2190,N_2465);
xnor U4173 (N_4173,N_407,N_141);
or U4174 (N_4174,N_1758,N_2471);
nor U4175 (N_4175,N_670,N_2143);
xor U4176 (N_4176,N_569,N_1274);
or U4177 (N_4177,N_708,N_291);
or U4178 (N_4178,N_2251,N_2232);
or U4179 (N_4179,N_929,N_868);
nor U4180 (N_4180,N_217,N_1805);
nor U4181 (N_4181,N_1284,N_1312);
or U4182 (N_4182,N_1706,N_295);
nor U4183 (N_4183,N_1993,N_105);
nand U4184 (N_4184,N_685,N_1073);
and U4185 (N_4185,N_606,N_882);
and U4186 (N_4186,N_1345,N_1531);
nor U4187 (N_4187,N_1954,N_667);
nor U4188 (N_4188,N_1170,N_984);
and U4189 (N_4189,N_456,N_810);
and U4190 (N_4190,N_1683,N_1786);
nand U4191 (N_4191,N_1198,N_335);
nor U4192 (N_4192,N_159,N_1856);
nand U4193 (N_4193,N_14,N_1874);
xor U4194 (N_4194,N_1689,N_1899);
nand U4195 (N_4195,N_362,N_818);
nand U4196 (N_4196,N_1065,N_419);
xor U4197 (N_4197,N_891,N_1464);
and U4198 (N_4198,N_1679,N_2468);
xor U4199 (N_4199,N_2345,N_1576);
nor U4200 (N_4200,N_930,N_739);
or U4201 (N_4201,N_739,N_1071);
nor U4202 (N_4202,N_1861,N_26);
nor U4203 (N_4203,N_1109,N_642);
or U4204 (N_4204,N_245,N_1461);
and U4205 (N_4205,N_2495,N_328);
nor U4206 (N_4206,N_644,N_2018);
and U4207 (N_4207,N_281,N_918);
nor U4208 (N_4208,N_431,N_134);
nor U4209 (N_4209,N_1988,N_1452);
xnor U4210 (N_4210,N_748,N_2012);
or U4211 (N_4211,N_2356,N_311);
nand U4212 (N_4212,N_2334,N_1439);
nand U4213 (N_4213,N_744,N_175);
nand U4214 (N_4214,N_2244,N_2307);
or U4215 (N_4215,N_424,N_809);
nand U4216 (N_4216,N_1585,N_1359);
or U4217 (N_4217,N_2454,N_325);
or U4218 (N_4218,N_1995,N_33);
xor U4219 (N_4219,N_2292,N_2094);
xnor U4220 (N_4220,N_1031,N_1992);
and U4221 (N_4221,N_1741,N_527);
nor U4222 (N_4222,N_725,N_1609);
and U4223 (N_4223,N_429,N_1356);
and U4224 (N_4224,N_989,N_1358);
nand U4225 (N_4225,N_315,N_748);
nand U4226 (N_4226,N_1120,N_2272);
nand U4227 (N_4227,N_2370,N_2283);
nor U4228 (N_4228,N_991,N_906);
nand U4229 (N_4229,N_1494,N_2310);
nand U4230 (N_4230,N_1578,N_1372);
and U4231 (N_4231,N_389,N_2252);
nor U4232 (N_4232,N_815,N_428);
nor U4233 (N_4233,N_2134,N_2110);
nor U4234 (N_4234,N_90,N_276);
nand U4235 (N_4235,N_538,N_64);
nor U4236 (N_4236,N_546,N_1639);
nor U4237 (N_4237,N_2104,N_7);
xor U4238 (N_4238,N_429,N_2047);
or U4239 (N_4239,N_2086,N_1976);
and U4240 (N_4240,N_125,N_2272);
or U4241 (N_4241,N_1961,N_1892);
or U4242 (N_4242,N_369,N_161);
or U4243 (N_4243,N_1686,N_1401);
and U4244 (N_4244,N_1671,N_2019);
nor U4245 (N_4245,N_1587,N_1799);
xnor U4246 (N_4246,N_558,N_1309);
or U4247 (N_4247,N_1474,N_1636);
nand U4248 (N_4248,N_501,N_1086);
nand U4249 (N_4249,N_1225,N_1817);
or U4250 (N_4250,N_2494,N_1283);
nand U4251 (N_4251,N_963,N_636);
nand U4252 (N_4252,N_2404,N_875);
or U4253 (N_4253,N_1777,N_168);
nand U4254 (N_4254,N_1129,N_1128);
and U4255 (N_4255,N_896,N_1755);
nand U4256 (N_4256,N_79,N_274);
or U4257 (N_4257,N_2235,N_1789);
nor U4258 (N_4258,N_1758,N_1488);
nand U4259 (N_4259,N_2207,N_1011);
nand U4260 (N_4260,N_304,N_1595);
xnor U4261 (N_4261,N_979,N_470);
xnor U4262 (N_4262,N_619,N_1938);
or U4263 (N_4263,N_672,N_347);
and U4264 (N_4264,N_646,N_1227);
and U4265 (N_4265,N_1760,N_638);
or U4266 (N_4266,N_1136,N_1305);
nand U4267 (N_4267,N_1258,N_330);
or U4268 (N_4268,N_1001,N_2255);
nor U4269 (N_4269,N_1424,N_1228);
nor U4270 (N_4270,N_1944,N_1048);
or U4271 (N_4271,N_309,N_1877);
nor U4272 (N_4272,N_364,N_301);
and U4273 (N_4273,N_1293,N_795);
nand U4274 (N_4274,N_2221,N_1716);
and U4275 (N_4275,N_2317,N_1829);
xor U4276 (N_4276,N_1843,N_745);
or U4277 (N_4277,N_2160,N_71);
nor U4278 (N_4278,N_563,N_890);
nand U4279 (N_4279,N_906,N_2094);
and U4280 (N_4280,N_2387,N_341);
or U4281 (N_4281,N_193,N_2009);
and U4282 (N_4282,N_1401,N_1043);
nor U4283 (N_4283,N_159,N_1397);
and U4284 (N_4284,N_1448,N_1567);
and U4285 (N_4285,N_2233,N_1386);
nand U4286 (N_4286,N_1610,N_1855);
nand U4287 (N_4287,N_362,N_846);
or U4288 (N_4288,N_1855,N_444);
nand U4289 (N_4289,N_1449,N_130);
nand U4290 (N_4290,N_1576,N_2310);
xor U4291 (N_4291,N_2077,N_209);
or U4292 (N_4292,N_1846,N_2323);
nand U4293 (N_4293,N_438,N_1430);
and U4294 (N_4294,N_1056,N_2179);
nand U4295 (N_4295,N_1112,N_65);
and U4296 (N_4296,N_319,N_799);
or U4297 (N_4297,N_1303,N_441);
nor U4298 (N_4298,N_1685,N_2236);
nor U4299 (N_4299,N_1744,N_2347);
or U4300 (N_4300,N_1175,N_1004);
nand U4301 (N_4301,N_1674,N_2081);
nor U4302 (N_4302,N_1458,N_2364);
and U4303 (N_4303,N_2011,N_1507);
and U4304 (N_4304,N_258,N_411);
or U4305 (N_4305,N_1646,N_1299);
nand U4306 (N_4306,N_2292,N_297);
nand U4307 (N_4307,N_512,N_1805);
xnor U4308 (N_4308,N_335,N_2392);
or U4309 (N_4309,N_241,N_97);
xor U4310 (N_4310,N_2490,N_175);
xor U4311 (N_4311,N_1320,N_479);
nor U4312 (N_4312,N_2201,N_1563);
or U4313 (N_4313,N_979,N_1767);
and U4314 (N_4314,N_760,N_165);
nor U4315 (N_4315,N_1538,N_2149);
or U4316 (N_4316,N_1973,N_2083);
or U4317 (N_4317,N_1922,N_2119);
or U4318 (N_4318,N_1046,N_236);
nand U4319 (N_4319,N_102,N_2069);
nand U4320 (N_4320,N_847,N_1588);
nand U4321 (N_4321,N_1643,N_397);
nand U4322 (N_4322,N_1864,N_2117);
nor U4323 (N_4323,N_2397,N_1226);
and U4324 (N_4324,N_1416,N_558);
nand U4325 (N_4325,N_1433,N_52);
xnor U4326 (N_4326,N_380,N_580);
or U4327 (N_4327,N_1768,N_830);
nand U4328 (N_4328,N_68,N_734);
and U4329 (N_4329,N_993,N_2362);
and U4330 (N_4330,N_972,N_1238);
or U4331 (N_4331,N_1736,N_2141);
or U4332 (N_4332,N_1217,N_2008);
nor U4333 (N_4333,N_203,N_2034);
and U4334 (N_4334,N_180,N_299);
nor U4335 (N_4335,N_1596,N_1802);
and U4336 (N_4336,N_328,N_1542);
nor U4337 (N_4337,N_642,N_1204);
or U4338 (N_4338,N_720,N_1130);
and U4339 (N_4339,N_2220,N_2304);
and U4340 (N_4340,N_1696,N_1353);
and U4341 (N_4341,N_3,N_1249);
or U4342 (N_4342,N_348,N_710);
and U4343 (N_4343,N_282,N_501);
nor U4344 (N_4344,N_1066,N_476);
nor U4345 (N_4345,N_1308,N_79);
nor U4346 (N_4346,N_171,N_412);
nand U4347 (N_4347,N_1510,N_715);
nand U4348 (N_4348,N_1377,N_976);
nand U4349 (N_4349,N_1073,N_1352);
nand U4350 (N_4350,N_1037,N_2352);
nand U4351 (N_4351,N_430,N_2062);
and U4352 (N_4352,N_1759,N_2057);
and U4353 (N_4353,N_1577,N_569);
and U4354 (N_4354,N_47,N_704);
and U4355 (N_4355,N_1855,N_536);
nand U4356 (N_4356,N_1599,N_1934);
nor U4357 (N_4357,N_1440,N_560);
or U4358 (N_4358,N_542,N_1724);
xor U4359 (N_4359,N_651,N_1238);
and U4360 (N_4360,N_731,N_2095);
nor U4361 (N_4361,N_1412,N_1956);
nor U4362 (N_4362,N_2454,N_774);
and U4363 (N_4363,N_1601,N_571);
nor U4364 (N_4364,N_169,N_468);
nor U4365 (N_4365,N_28,N_415);
nor U4366 (N_4366,N_1893,N_288);
nand U4367 (N_4367,N_178,N_2058);
or U4368 (N_4368,N_1446,N_1024);
or U4369 (N_4369,N_260,N_492);
nand U4370 (N_4370,N_1703,N_961);
and U4371 (N_4371,N_1412,N_185);
xor U4372 (N_4372,N_2134,N_1811);
or U4373 (N_4373,N_1124,N_835);
or U4374 (N_4374,N_1520,N_1197);
and U4375 (N_4375,N_1193,N_280);
or U4376 (N_4376,N_2187,N_1805);
nand U4377 (N_4377,N_1662,N_2321);
and U4378 (N_4378,N_1870,N_1367);
or U4379 (N_4379,N_1684,N_1431);
or U4380 (N_4380,N_225,N_1280);
nor U4381 (N_4381,N_2482,N_372);
nand U4382 (N_4382,N_1716,N_932);
nor U4383 (N_4383,N_391,N_176);
nand U4384 (N_4384,N_2327,N_2262);
xor U4385 (N_4385,N_148,N_1165);
and U4386 (N_4386,N_1919,N_21);
or U4387 (N_4387,N_1455,N_1588);
and U4388 (N_4388,N_1828,N_1331);
or U4389 (N_4389,N_2106,N_78);
or U4390 (N_4390,N_174,N_2257);
nand U4391 (N_4391,N_1911,N_1800);
or U4392 (N_4392,N_412,N_1462);
or U4393 (N_4393,N_702,N_1617);
nor U4394 (N_4394,N_1718,N_1990);
nor U4395 (N_4395,N_2414,N_932);
or U4396 (N_4396,N_739,N_202);
nand U4397 (N_4397,N_1084,N_2007);
xnor U4398 (N_4398,N_1437,N_458);
and U4399 (N_4399,N_787,N_2412);
nor U4400 (N_4400,N_811,N_416);
nor U4401 (N_4401,N_1291,N_960);
and U4402 (N_4402,N_970,N_2468);
and U4403 (N_4403,N_1032,N_989);
or U4404 (N_4404,N_1086,N_1612);
and U4405 (N_4405,N_474,N_1728);
nor U4406 (N_4406,N_2192,N_281);
nand U4407 (N_4407,N_651,N_1686);
and U4408 (N_4408,N_1008,N_508);
nor U4409 (N_4409,N_2132,N_2299);
nor U4410 (N_4410,N_1273,N_772);
nor U4411 (N_4411,N_1483,N_870);
nand U4412 (N_4412,N_1945,N_1941);
or U4413 (N_4413,N_2497,N_1005);
xnor U4414 (N_4414,N_1916,N_1322);
nand U4415 (N_4415,N_1232,N_1077);
or U4416 (N_4416,N_852,N_1941);
nor U4417 (N_4417,N_1736,N_264);
or U4418 (N_4418,N_1875,N_926);
and U4419 (N_4419,N_858,N_1470);
xor U4420 (N_4420,N_432,N_2389);
nor U4421 (N_4421,N_2103,N_1499);
nand U4422 (N_4422,N_869,N_2281);
or U4423 (N_4423,N_2270,N_1561);
or U4424 (N_4424,N_897,N_672);
nand U4425 (N_4425,N_990,N_1610);
or U4426 (N_4426,N_2167,N_1254);
and U4427 (N_4427,N_62,N_75);
nand U4428 (N_4428,N_1126,N_1663);
nand U4429 (N_4429,N_972,N_801);
or U4430 (N_4430,N_337,N_1816);
nor U4431 (N_4431,N_2004,N_2106);
nor U4432 (N_4432,N_1455,N_1614);
or U4433 (N_4433,N_1860,N_1393);
or U4434 (N_4434,N_2113,N_637);
and U4435 (N_4435,N_579,N_1564);
nand U4436 (N_4436,N_1103,N_1693);
nor U4437 (N_4437,N_1619,N_2336);
nand U4438 (N_4438,N_222,N_2237);
and U4439 (N_4439,N_1187,N_771);
xnor U4440 (N_4440,N_685,N_1586);
nand U4441 (N_4441,N_1013,N_1521);
or U4442 (N_4442,N_1505,N_678);
xnor U4443 (N_4443,N_573,N_1588);
xor U4444 (N_4444,N_2332,N_1371);
and U4445 (N_4445,N_1972,N_522);
nand U4446 (N_4446,N_590,N_277);
and U4447 (N_4447,N_2201,N_2352);
or U4448 (N_4448,N_2209,N_1664);
nor U4449 (N_4449,N_1717,N_529);
or U4450 (N_4450,N_1550,N_889);
nand U4451 (N_4451,N_1846,N_1154);
or U4452 (N_4452,N_1219,N_99);
nand U4453 (N_4453,N_1481,N_2309);
and U4454 (N_4454,N_414,N_165);
or U4455 (N_4455,N_1303,N_965);
or U4456 (N_4456,N_1351,N_2320);
nand U4457 (N_4457,N_1186,N_2004);
nor U4458 (N_4458,N_2206,N_2295);
or U4459 (N_4459,N_861,N_1812);
or U4460 (N_4460,N_1773,N_1179);
and U4461 (N_4461,N_586,N_2175);
nor U4462 (N_4462,N_1697,N_1350);
nand U4463 (N_4463,N_2441,N_2166);
or U4464 (N_4464,N_98,N_494);
or U4465 (N_4465,N_2064,N_503);
nor U4466 (N_4466,N_1605,N_140);
or U4467 (N_4467,N_89,N_1214);
xor U4468 (N_4468,N_782,N_226);
or U4469 (N_4469,N_1658,N_1818);
nand U4470 (N_4470,N_766,N_1655);
and U4471 (N_4471,N_1811,N_54);
and U4472 (N_4472,N_2380,N_2012);
and U4473 (N_4473,N_605,N_836);
nor U4474 (N_4474,N_1749,N_2085);
and U4475 (N_4475,N_1190,N_1574);
and U4476 (N_4476,N_1374,N_2283);
nand U4477 (N_4477,N_403,N_1241);
nand U4478 (N_4478,N_615,N_1092);
nand U4479 (N_4479,N_2495,N_278);
nor U4480 (N_4480,N_719,N_1783);
nand U4481 (N_4481,N_487,N_167);
nand U4482 (N_4482,N_2226,N_1164);
nor U4483 (N_4483,N_238,N_1785);
nor U4484 (N_4484,N_1911,N_1736);
xnor U4485 (N_4485,N_683,N_305);
nand U4486 (N_4486,N_1400,N_410);
nor U4487 (N_4487,N_1061,N_1213);
nor U4488 (N_4488,N_2244,N_360);
or U4489 (N_4489,N_126,N_97);
and U4490 (N_4490,N_2458,N_264);
nand U4491 (N_4491,N_1025,N_2309);
or U4492 (N_4492,N_287,N_932);
and U4493 (N_4493,N_1589,N_669);
xor U4494 (N_4494,N_2108,N_80);
nand U4495 (N_4495,N_401,N_311);
and U4496 (N_4496,N_160,N_46);
and U4497 (N_4497,N_2058,N_2180);
nand U4498 (N_4498,N_734,N_485);
or U4499 (N_4499,N_1082,N_2276);
nand U4500 (N_4500,N_2164,N_2285);
xor U4501 (N_4501,N_1704,N_2437);
nor U4502 (N_4502,N_1250,N_1378);
nor U4503 (N_4503,N_1542,N_1113);
or U4504 (N_4504,N_219,N_1159);
and U4505 (N_4505,N_19,N_571);
nand U4506 (N_4506,N_56,N_305);
xnor U4507 (N_4507,N_921,N_2104);
nand U4508 (N_4508,N_1155,N_1607);
nor U4509 (N_4509,N_1225,N_612);
nor U4510 (N_4510,N_329,N_2387);
nand U4511 (N_4511,N_1252,N_2038);
nor U4512 (N_4512,N_1075,N_2360);
and U4513 (N_4513,N_498,N_696);
and U4514 (N_4514,N_1161,N_2232);
nand U4515 (N_4515,N_1310,N_524);
and U4516 (N_4516,N_358,N_1121);
nor U4517 (N_4517,N_1544,N_495);
nor U4518 (N_4518,N_277,N_1819);
and U4519 (N_4519,N_1928,N_384);
or U4520 (N_4520,N_1291,N_984);
xnor U4521 (N_4521,N_808,N_2453);
and U4522 (N_4522,N_1201,N_378);
and U4523 (N_4523,N_431,N_696);
nand U4524 (N_4524,N_736,N_573);
and U4525 (N_4525,N_22,N_2404);
or U4526 (N_4526,N_554,N_1674);
nor U4527 (N_4527,N_531,N_1947);
nand U4528 (N_4528,N_1709,N_1228);
and U4529 (N_4529,N_1459,N_267);
nor U4530 (N_4530,N_104,N_1566);
nand U4531 (N_4531,N_2481,N_2217);
or U4532 (N_4532,N_1459,N_297);
nor U4533 (N_4533,N_107,N_2254);
nor U4534 (N_4534,N_1648,N_257);
or U4535 (N_4535,N_2214,N_1674);
nand U4536 (N_4536,N_214,N_2211);
nor U4537 (N_4537,N_2295,N_1248);
or U4538 (N_4538,N_2034,N_1863);
nand U4539 (N_4539,N_2273,N_767);
and U4540 (N_4540,N_863,N_2277);
or U4541 (N_4541,N_1709,N_178);
or U4542 (N_4542,N_1565,N_247);
nor U4543 (N_4543,N_235,N_142);
nand U4544 (N_4544,N_69,N_1654);
nor U4545 (N_4545,N_596,N_2062);
and U4546 (N_4546,N_1461,N_1908);
nor U4547 (N_4547,N_2151,N_796);
and U4548 (N_4548,N_569,N_2345);
and U4549 (N_4549,N_1151,N_932);
and U4550 (N_4550,N_2067,N_1176);
nand U4551 (N_4551,N_884,N_2368);
and U4552 (N_4552,N_1524,N_1897);
and U4553 (N_4553,N_384,N_815);
or U4554 (N_4554,N_1581,N_1260);
nor U4555 (N_4555,N_1996,N_2416);
nand U4556 (N_4556,N_595,N_2009);
nand U4557 (N_4557,N_2050,N_1549);
xnor U4558 (N_4558,N_27,N_39);
and U4559 (N_4559,N_1819,N_1946);
nor U4560 (N_4560,N_592,N_1282);
nand U4561 (N_4561,N_1619,N_111);
and U4562 (N_4562,N_1596,N_745);
nand U4563 (N_4563,N_1616,N_480);
or U4564 (N_4564,N_227,N_177);
nor U4565 (N_4565,N_1265,N_891);
nand U4566 (N_4566,N_599,N_1894);
or U4567 (N_4567,N_1655,N_1326);
xnor U4568 (N_4568,N_2133,N_192);
or U4569 (N_4569,N_1146,N_717);
nand U4570 (N_4570,N_2058,N_1278);
nand U4571 (N_4571,N_1202,N_1708);
nor U4572 (N_4572,N_1452,N_710);
nor U4573 (N_4573,N_1163,N_783);
nand U4574 (N_4574,N_686,N_71);
and U4575 (N_4575,N_661,N_1779);
or U4576 (N_4576,N_1508,N_1380);
xor U4577 (N_4577,N_477,N_1169);
and U4578 (N_4578,N_666,N_1657);
and U4579 (N_4579,N_2219,N_1343);
nand U4580 (N_4580,N_768,N_109);
or U4581 (N_4581,N_1419,N_929);
nor U4582 (N_4582,N_2083,N_2249);
and U4583 (N_4583,N_666,N_117);
xnor U4584 (N_4584,N_1595,N_984);
nor U4585 (N_4585,N_742,N_1409);
xnor U4586 (N_4586,N_2372,N_1595);
xor U4587 (N_4587,N_1061,N_54);
and U4588 (N_4588,N_2350,N_737);
nand U4589 (N_4589,N_1106,N_1846);
nand U4590 (N_4590,N_574,N_438);
xnor U4591 (N_4591,N_461,N_60);
or U4592 (N_4592,N_1508,N_2175);
nor U4593 (N_4593,N_2389,N_1226);
or U4594 (N_4594,N_900,N_2251);
or U4595 (N_4595,N_935,N_1261);
or U4596 (N_4596,N_1222,N_2432);
or U4597 (N_4597,N_1979,N_721);
xnor U4598 (N_4598,N_2155,N_759);
nor U4599 (N_4599,N_1490,N_1413);
nor U4600 (N_4600,N_2188,N_728);
or U4601 (N_4601,N_798,N_2186);
nand U4602 (N_4602,N_1935,N_1090);
or U4603 (N_4603,N_2300,N_1780);
nor U4604 (N_4604,N_1190,N_1383);
nand U4605 (N_4605,N_571,N_899);
nand U4606 (N_4606,N_492,N_388);
and U4607 (N_4607,N_2007,N_861);
and U4608 (N_4608,N_2464,N_1000);
nand U4609 (N_4609,N_318,N_1180);
and U4610 (N_4610,N_2021,N_1567);
or U4611 (N_4611,N_737,N_726);
nand U4612 (N_4612,N_2026,N_681);
nand U4613 (N_4613,N_2238,N_1125);
nand U4614 (N_4614,N_709,N_2487);
or U4615 (N_4615,N_1974,N_1023);
nor U4616 (N_4616,N_1949,N_1757);
and U4617 (N_4617,N_1521,N_1753);
nand U4618 (N_4618,N_1863,N_770);
or U4619 (N_4619,N_2498,N_2489);
xor U4620 (N_4620,N_1527,N_2464);
xor U4621 (N_4621,N_1232,N_91);
nor U4622 (N_4622,N_2189,N_1718);
or U4623 (N_4623,N_647,N_291);
nand U4624 (N_4624,N_1938,N_158);
and U4625 (N_4625,N_1417,N_852);
and U4626 (N_4626,N_1010,N_826);
and U4627 (N_4627,N_2303,N_1031);
and U4628 (N_4628,N_2117,N_585);
nand U4629 (N_4629,N_881,N_1167);
nor U4630 (N_4630,N_448,N_269);
nor U4631 (N_4631,N_1151,N_333);
and U4632 (N_4632,N_1064,N_1628);
or U4633 (N_4633,N_968,N_1647);
or U4634 (N_4634,N_813,N_1489);
and U4635 (N_4635,N_301,N_1849);
nand U4636 (N_4636,N_418,N_2182);
or U4637 (N_4637,N_641,N_1780);
nor U4638 (N_4638,N_1806,N_1280);
xnor U4639 (N_4639,N_134,N_2351);
or U4640 (N_4640,N_1439,N_422);
or U4641 (N_4641,N_281,N_1721);
or U4642 (N_4642,N_658,N_408);
nor U4643 (N_4643,N_1789,N_2120);
and U4644 (N_4644,N_282,N_1028);
or U4645 (N_4645,N_1348,N_1699);
nand U4646 (N_4646,N_1213,N_1326);
nand U4647 (N_4647,N_1186,N_1782);
and U4648 (N_4648,N_1928,N_316);
and U4649 (N_4649,N_1317,N_1759);
nor U4650 (N_4650,N_2372,N_1006);
nor U4651 (N_4651,N_1957,N_2184);
nand U4652 (N_4652,N_2135,N_1154);
and U4653 (N_4653,N_6,N_2247);
or U4654 (N_4654,N_1302,N_881);
and U4655 (N_4655,N_973,N_1633);
nor U4656 (N_4656,N_1784,N_1688);
nor U4657 (N_4657,N_1150,N_2465);
nand U4658 (N_4658,N_1338,N_585);
nor U4659 (N_4659,N_627,N_999);
and U4660 (N_4660,N_2233,N_739);
or U4661 (N_4661,N_143,N_1573);
nor U4662 (N_4662,N_1656,N_1176);
nand U4663 (N_4663,N_1836,N_1535);
nor U4664 (N_4664,N_1419,N_509);
or U4665 (N_4665,N_2370,N_1709);
nor U4666 (N_4666,N_1587,N_1531);
nand U4667 (N_4667,N_1714,N_959);
nand U4668 (N_4668,N_1218,N_1119);
nor U4669 (N_4669,N_2047,N_2155);
or U4670 (N_4670,N_113,N_1777);
nor U4671 (N_4671,N_2426,N_188);
nor U4672 (N_4672,N_488,N_61);
xnor U4673 (N_4673,N_213,N_665);
nor U4674 (N_4674,N_2185,N_43);
or U4675 (N_4675,N_399,N_1552);
nand U4676 (N_4676,N_268,N_71);
and U4677 (N_4677,N_1448,N_871);
xnor U4678 (N_4678,N_293,N_1717);
nand U4679 (N_4679,N_400,N_976);
nand U4680 (N_4680,N_177,N_198);
or U4681 (N_4681,N_1922,N_419);
or U4682 (N_4682,N_2299,N_1515);
and U4683 (N_4683,N_766,N_2227);
xor U4684 (N_4684,N_358,N_680);
or U4685 (N_4685,N_1027,N_2181);
nand U4686 (N_4686,N_1631,N_1463);
nand U4687 (N_4687,N_473,N_2111);
nor U4688 (N_4688,N_1544,N_1275);
xor U4689 (N_4689,N_1973,N_2415);
and U4690 (N_4690,N_2310,N_2439);
nand U4691 (N_4691,N_943,N_1788);
or U4692 (N_4692,N_1531,N_1281);
nor U4693 (N_4693,N_696,N_595);
and U4694 (N_4694,N_2021,N_545);
nand U4695 (N_4695,N_742,N_237);
nand U4696 (N_4696,N_1122,N_137);
and U4697 (N_4697,N_688,N_1860);
and U4698 (N_4698,N_1086,N_1302);
nor U4699 (N_4699,N_752,N_1868);
nor U4700 (N_4700,N_1440,N_1082);
and U4701 (N_4701,N_64,N_1108);
nor U4702 (N_4702,N_2435,N_396);
or U4703 (N_4703,N_2440,N_1203);
or U4704 (N_4704,N_1918,N_1034);
xor U4705 (N_4705,N_1628,N_296);
and U4706 (N_4706,N_1670,N_2260);
nand U4707 (N_4707,N_976,N_1996);
or U4708 (N_4708,N_810,N_1642);
or U4709 (N_4709,N_1266,N_682);
nor U4710 (N_4710,N_1250,N_1389);
nor U4711 (N_4711,N_282,N_1194);
nand U4712 (N_4712,N_1523,N_1191);
or U4713 (N_4713,N_249,N_1081);
or U4714 (N_4714,N_2061,N_724);
xnor U4715 (N_4715,N_512,N_1745);
nor U4716 (N_4716,N_488,N_44);
nand U4717 (N_4717,N_339,N_864);
nor U4718 (N_4718,N_587,N_245);
xor U4719 (N_4719,N_1049,N_98);
and U4720 (N_4720,N_2231,N_1092);
nand U4721 (N_4721,N_798,N_1362);
and U4722 (N_4722,N_2416,N_1153);
or U4723 (N_4723,N_1287,N_1046);
and U4724 (N_4724,N_353,N_2133);
or U4725 (N_4725,N_822,N_731);
and U4726 (N_4726,N_1708,N_1740);
or U4727 (N_4727,N_2302,N_2172);
and U4728 (N_4728,N_1665,N_2021);
or U4729 (N_4729,N_464,N_2125);
and U4730 (N_4730,N_1198,N_1583);
or U4731 (N_4731,N_709,N_400);
or U4732 (N_4732,N_675,N_1882);
xnor U4733 (N_4733,N_1914,N_521);
and U4734 (N_4734,N_496,N_2038);
nor U4735 (N_4735,N_727,N_2167);
nor U4736 (N_4736,N_983,N_1760);
and U4737 (N_4737,N_1273,N_956);
nand U4738 (N_4738,N_1640,N_417);
nand U4739 (N_4739,N_1867,N_1712);
or U4740 (N_4740,N_1434,N_399);
nand U4741 (N_4741,N_1568,N_471);
or U4742 (N_4742,N_970,N_1968);
nand U4743 (N_4743,N_1042,N_1302);
nand U4744 (N_4744,N_1413,N_409);
xor U4745 (N_4745,N_467,N_191);
nand U4746 (N_4746,N_1533,N_884);
and U4747 (N_4747,N_1993,N_137);
nor U4748 (N_4748,N_2035,N_511);
nand U4749 (N_4749,N_1385,N_1912);
or U4750 (N_4750,N_974,N_2184);
nor U4751 (N_4751,N_695,N_1675);
and U4752 (N_4752,N_1761,N_1882);
nand U4753 (N_4753,N_641,N_248);
nand U4754 (N_4754,N_810,N_2441);
or U4755 (N_4755,N_2113,N_928);
nor U4756 (N_4756,N_1743,N_2360);
nor U4757 (N_4757,N_677,N_740);
or U4758 (N_4758,N_2220,N_2476);
or U4759 (N_4759,N_2048,N_79);
xor U4760 (N_4760,N_702,N_1281);
and U4761 (N_4761,N_492,N_54);
or U4762 (N_4762,N_671,N_1216);
or U4763 (N_4763,N_2387,N_200);
nor U4764 (N_4764,N_1540,N_309);
nor U4765 (N_4765,N_396,N_425);
nand U4766 (N_4766,N_1039,N_627);
nor U4767 (N_4767,N_2379,N_2256);
nor U4768 (N_4768,N_1403,N_849);
or U4769 (N_4769,N_1197,N_816);
nand U4770 (N_4770,N_2290,N_2356);
and U4771 (N_4771,N_159,N_483);
nor U4772 (N_4772,N_2460,N_1134);
nor U4773 (N_4773,N_1357,N_2265);
and U4774 (N_4774,N_791,N_1133);
nor U4775 (N_4775,N_1520,N_1905);
xnor U4776 (N_4776,N_697,N_2124);
or U4777 (N_4777,N_1656,N_139);
nor U4778 (N_4778,N_2178,N_1255);
and U4779 (N_4779,N_398,N_161);
and U4780 (N_4780,N_312,N_2018);
and U4781 (N_4781,N_1743,N_821);
nand U4782 (N_4782,N_2421,N_2228);
xnor U4783 (N_4783,N_223,N_1677);
nor U4784 (N_4784,N_403,N_2163);
and U4785 (N_4785,N_2181,N_1374);
and U4786 (N_4786,N_1268,N_1281);
nand U4787 (N_4787,N_1287,N_1173);
and U4788 (N_4788,N_469,N_1594);
nand U4789 (N_4789,N_2013,N_2109);
and U4790 (N_4790,N_2258,N_545);
nand U4791 (N_4791,N_1328,N_1834);
nor U4792 (N_4792,N_2492,N_1997);
nand U4793 (N_4793,N_930,N_2385);
or U4794 (N_4794,N_1714,N_1644);
or U4795 (N_4795,N_1184,N_1950);
and U4796 (N_4796,N_1785,N_194);
and U4797 (N_4797,N_17,N_1254);
nor U4798 (N_4798,N_1939,N_2115);
nor U4799 (N_4799,N_2185,N_1463);
and U4800 (N_4800,N_2318,N_834);
or U4801 (N_4801,N_839,N_1532);
and U4802 (N_4802,N_2292,N_2320);
and U4803 (N_4803,N_1852,N_979);
and U4804 (N_4804,N_2305,N_989);
nand U4805 (N_4805,N_2212,N_77);
or U4806 (N_4806,N_798,N_2479);
and U4807 (N_4807,N_2313,N_1103);
xor U4808 (N_4808,N_1463,N_546);
and U4809 (N_4809,N_1728,N_2);
or U4810 (N_4810,N_1149,N_2371);
and U4811 (N_4811,N_1833,N_523);
nand U4812 (N_4812,N_1280,N_753);
nor U4813 (N_4813,N_535,N_801);
and U4814 (N_4814,N_719,N_2497);
nand U4815 (N_4815,N_1174,N_2462);
nor U4816 (N_4816,N_1549,N_736);
or U4817 (N_4817,N_629,N_116);
nand U4818 (N_4818,N_897,N_1295);
xor U4819 (N_4819,N_66,N_2200);
or U4820 (N_4820,N_1535,N_959);
or U4821 (N_4821,N_1567,N_1269);
and U4822 (N_4822,N_1412,N_1179);
nand U4823 (N_4823,N_1208,N_1053);
nor U4824 (N_4824,N_1312,N_1849);
nor U4825 (N_4825,N_1983,N_2368);
nor U4826 (N_4826,N_931,N_1696);
nor U4827 (N_4827,N_826,N_1124);
xnor U4828 (N_4828,N_362,N_363);
nand U4829 (N_4829,N_625,N_2345);
nand U4830 (N_4830,N_1409,N_563);
and U4831 (N_4831,N_1307,N_904);
or U4832 (N_4832,N_1310,N_1331);
nand U4833 (N_4833,N_1284,N_1938);
nor U4834 (N_4834,N_64,N_2122);
nor U4835 (N_4835,N_31,N_1730);
nor U4836 (N_4836,N_1466,N_2370);
xor U4837 (N_4837,N_1926,N_1568);
and U4838 (N_4838,N_94,N_1640);
nand U4839 (N_4839,N_1693,N_492);
nand U4840 (N_4840,N_2347,N_74);
nand U4841 (N_4841,N_18,N_240);
nand U4842 (N_4842,N_397,N_2329);
nor U4843 (N_4843,N_2357,N_289);
or U4844 (N_4844,N_620,N_382);
or U4845 (N_4845,N_1134,N_1007);
and U4846 (N_4846,N_865,N_1243);
and U4847 (N_4847,N_104,N_658);
nor U4848 (N_4848,N_1294,N_942);
and U4849 (N_4849,N_1624,N_1376);
or U4850 (N_4850,N_2089,N_2274);
or U4851 (N_4851,N_1356,N_2450);
nor U4852 (N_4852,N_740,N_1244);
and U4853 (N_4853,N_746,N_2087);
and U4854 (N_4854,N_119,N_123);
nand U4855 (N_4855,N_940,N_2312);
nor U4856 (N_4856,N_209,N_689);
xnor U4857 (N_4857,N_19,N_192);
or U4858 (N_4858,N_1085,N_2280);
or U4859 (N_4859,N_718,N_2392);
and U4860 (N_4860,N_1948,N_367);
or U4861 (N_4861,N_1565,N_2150);
nor U4862 (N_4862,N_1173,N_817);
nand U4863 (N_4863,N_1473,N_1951);
or U4864 (N_4864,N_506,N_1103);
or U4865 (N_4865,N_566,N_2368);
nor U4866 (N_4866,N_703,N_696);
or U4867 (N_4867,N_2490,N_886);
nand U4868 (N_4868,N_1291,N_2017);
nor U4869 (N_4869,N_2217,N_1127);
nor U4870 (N_4870,N_2004,N_1011);
or U4871 (N_4871,N_1839,N_1454);
xnor U4872 (N_4872,N_231,N_703);
nor U4873 (N_4873,N_1847,N_1918);
nand U4874 (N_4874,N_525,N_1291);
nand U4875 (N_4875,N_1405,N_42);
xnor U4876 (N_4876,N_2138,N_108);
nor U4877 (N_4877,N_1300,N_1506);
nor U4878 (N_4878,N_1975,N_438);
and U4879 (N_4879,N_1142,N_645);
xnor U4880 (N_4880,N_1248,N_58);
or U4881 (N_4881,N_1880,N_883);
xnor U4882 (N_4882,N_132,N_1762);
nor U4883 (N_4883,N_490,N_1728);
and U4884 (N_4884,N_1797,N_2118);
and U4885 (N_4885,N_962,N_950);
and U4886 (N_4886,N_1431,N_1110);
nand U4887 (N_4887,N_1365,N_2025);
or U4888 (N_4888,N_684,N_883);
or U4889 (N_4889,N_1950,N_624);
nor U4890 (N_4890,N_1694,N_1546);
and U4891 (N_4891,N_260,N_875);
and U4892 (N_4892,N_809,N_771);
nand U4893 (N_4893,N_1319,N_1932);
and U4894 (N_4894,N_1699,N_1474);
and U4895 (N_4895,N_1311,N_413);
and U4896 (N_4896,N_772,N_1743);
or U4897 (N_4897,N_469,N_2394);
and U4898 (N_4898,N_1543,N_1356);
and U4899 (N_4899,N_2104,N_587);
xor U4900 (N_4900,N_262,N_1237);
and U4901 (N_4901,N_423,N_2358);
or U4902 (N_4902,N_1408,N_1983);
or U4903 (N_4903,N_1608,N_1388);
nor U4904 (N_4904,N_1277,N_491);
nand U4905 (N_4905,N_2112,N_2202);
and U4906 (N_4906,N_2217,N_2044);
or U4907 (N_4907,N_1827,N_1328);
nand U4908 (N_4908,N_2477,N_439);
or U4909 (N_4909,N_899,N_1744);
and U4910 (N_4910,N_21,N_2479);
nand U4911 (N_4911,N_1415,N_1681);
or U4912 (N_4912,N_1478,N_1506);
xor U4913 (N_4913,N_2410,N_2213);
and U4914 (N_4914,N_2078,N_936);
or U4915 (N_4915,N_559,N_2333);
nor U4916 (N_4916,N_2299,N_806);
nor U4917 (N_4917,N_1832,N_723);
nand U4918 (N_4918,N_587,N_369);
and U4919 (N_4919,N_1166,N_977);
nor U4920 (N_4920,N_2215,N_1872);
or U4921 (N_4921,N_394,N_1407);
nand U4922 (N_4922,N_472,N_1886);
nor U4923 (N_4923,N_215,N_1355);
nand U4924 (N_4924,N_539,N_2168);
nand U4925 (N_4925,N_41,N_667);
nand U4926 (N_4926,N_2098,N_2240);
nor U4927 (N_4927,N_469,N_2471);
nand U4928 (N_4928,N_796,N_1042);
or U4929 (N_4929,N_1332,N_1141);
nor U4930 (N_4930,N_960,N_604);
nand U4931 (N_4931,N_545,N_566);
nand U4932 (N_4932,N_1092,N_233);
or U4933 (N_4933,N_1710,N_1889);
xor U4934 (N_4934,N_2055,N_2348);
and U4935 (N_4935,N_76,N_218);
and U4936 (N_4936,N_448,N_16);
nand U4937 (N_4937,N_1383,N_1057);
and U4938 (N_4938,N_815,N_1943);
and U4939 (N_4939,N_2089,N_2349);
xor U4940 (N_4940,N_180,N_1905);
nand U4941 (N_4941,N_490,N_1073);
and U4942 (N_4942,N_971,N_344);
or U4943 (N_4943,N_220,N_2116);
and U4944 (N_4944,N_2288,N_749);
nand U4945 (N_4945,N_756,N_1632);
or U4946 (N_4946,N_1644,N_1441);
nor U4947 (N_4947,N_1449,N_1235);
nand U4948 (N_4948,N_2223,N_2282);
xnor U4949 (N_4949,N_1270,N_2170);
nor U4950 (N_4950,N_169,N_621);
xor U4951 (N_4951,N_1197,N_1107);
or U4952 (N_4952,N_2192,N_513);
nand U4953 (N_4953,N_2159,N_873);
nand U4954 (N_4954,N_2413,N_886);
xnor U4955 (N_4955,N_1969,N_1862);
xnor U4956 (N_4956,N_1862,N_630);
nand U4957 (N_4957,N_1467,N_2272);
xor U4958 (N_4958,N_2155,N_1343);
nand U4959 (N_4959,N_59,N_2278);
and U4960 (N_4960,N_1589,N_1995);
nor U4961 (N_4961,N_1231,N_1786);
nor U4962 (N_4962,N_1625,N_596);
nor U4963 (N_4963,N_2016,N_2331);
nor U4964 (N_4964,N_2011,N_1214);
and U4965 (N_4965,N_605,N_2149);
or U4966 (N_4966,N_2021,N_686);
nor U4967 (N_4967,N_797,N_2100);
nor U4968 (N_4968,N_2016,N_1286);
and U4969 (N_4969,N_1840,N_2308);
and U4970 (N_4970,N_1508,N_2457);
or U4971 (N_4971,N_558,N_1766);
nand U4972 (N_4972,N_1038,N_1147);
nand U4973 (N_4973,N_1126,N_2018);
nand U4974 (N_4974,N_15,N_1683);
nor U4975 (N_4975,N_333,N_2422);
nor U4976 (N_4976,N_1092,N_765);
and U4977 (N_4977,N_282,N_542);
nor U4978 (N_4978,N_887,N_1463);
nand U4979 (N_4979,N_1791,N_1305);
nor U4980 (N_4980,N_1416,N_796);
or U4981 (N_4981,N_1988,N_609);
or U4982 (N_4982,N_2255,N_668);
nand U4983 (N_4983,N_669,N_853);
and U4984 (N_4984,N_375,N_1442);
nor U4985 (N_4985,N_1330,N_683);
nand U4986 (N_4986,N_2188,N_14);
and U4987 (N_4987,N_1387,N_1257);
nand U4988 (N_4988,N_1007,N_329);
nand U4989 (N_4989,N_2434,N_2464);
xnor U4990 (N_4990,N_1572,N_1858);
and U4991 (N_4991,N_1870,N_855);
or U4992 (N_4992,N_77,N_1608);
nor U4993 (N_4993,N_1748,N_1861);
or U4994 (N_4994,N_1522,N_380);
and U4995 (N_4995,N_2441,N_761);
and U4996 (N_4996,N_1680,N_1776);
nand U4997 (N_4997,N_767,N_1258);
and U4998 (N_4998,N_72,N_1035);
xor U4999 (N_4999,N_2384,N_1827);
nor UO_0 (O_0,N_3691,N_4029);
nand UO_1 (O_1,N_3422,N_4513);
nand UO_2 (O_2,N_3331,N_3944);
or UO_3 (O_3,N_4900,N_4136);
or UO_4 (O_4,N_2628,N_4822);
and UO_5 (O_5,N_3720,N_3852);
and UO_6 (O_6,N_3829,N_4435);
nand UO_7 (O_7,N_2869,N_3345);
nand UO_8 (O_8,N_3049,N_4303);
nor UO_9 (O_9,N_4944,N_2824);
nand UO_10 (O_10,N_2768,N_3527);
or UO_11 (O_11,N_4797,N_2745);
or UO_12 (O_12,N_4264,N_4642);
or UO_13 (O_13,N_2584,N_4023);
or UO_14 (O_14,N_3734,N_2581);
nand UO_15 (O_15,N_3336,N_4466);
and UO_16 (O_16,N_4844,N_4973);
nor UO_17 (O_17,N_3958,N_4867);
or UO_18 (O_18,N_2653,N_3520);
nand UO_19 (O_19,N_3245,N_3226);
nand UO_20 (O_20,N_3246,N_4840);
nand UO_21 (O_21,N_3369,N_4362);
and UO_22 (O_22,N_3034,N_3714);
nor UO_23 (O_23,N_3024,N_4021);
and UO_24 (O_24,N_4724,N_3409);
nor UO_25 (O_25,N_3623,N_3982);
or UO_26 (O_26,N_3625,N_3269);
xor UO_27 (O_27,N_4637,N_3031);
and UO_28 (O_28,N_4942,N_2931);
and UO_29 (O_29,N_2678,N_3660);
and UO_30 (O_30,N_4184,N_3998);
nor UO_31 (O_31,N_2809,N_4327);
xnor UO_32 (O_32,N_4747,N_3203);
xor UO_33 (O_33,N_3806,N_4713);
or UO_34 (O_34,N_3755,N_2781);
nor UO_35 (O_35,N_3999,N_4054);
nor UO_36 (O_36,N_4076,N_4558);
or UO_37 (O_37,N_4420,N_2780);
or UO_38 (O_38,N_3193,N_3352);
or UO_39 (O_39,N_4798,N_2788);
xor UO_40 (O_40,N_3124,N_3259);
nor UO_41 (O_41,N_2693,N_4108);
nor UO_42 (O_42,N_3457,N_2711);
nor UO_43 (O_43,N_2990,N_3541);
nor UO_44 (O_44,N_3793,N_4200);
xor UO_45 (O_45,N_3753,N_3232);
xnor UO_46 (O_46,N_4727,N_4878);
nand UO_47 (O_47,N_3126,N_2838);
or UO_48 (O_48,N_3192,N_4735);
and UO_49 (O_49,N_3361,N_4147);
and UO_50 (O_50,N_3454,N_2671);
xor UO_51 (O_51,N_3041,N_2910);
nor UO_52 (O_52,N_4945,N_4879);
and UO_53 (O_53,N_4283,N_2734);
nand UO_54 (O_54,N_3693,N_4923);
xor UO_55 (O_55,N_4623,N_4324);
nand UO_56 (O_56,N_3611,N_4158);
or UO_57 (O_57,N_2511,N_4974);
or UO_58 (O_58,N_4116,N_2575);
nor UO_59 (O_59,N_4287,N_4492);
nor UO_60 (O_60,N_4133,N_3328);
or UO_61 (O_61,N_3140,N_3390);
nand UO_62 (O_62,N_3310,N_4203);
nand UO_63 (O_63,N_4534,N_3643);
nand UO_64 (O_64,N_2599,N_3272);
xnor UO_65 (O_65,N_4016,N_4070);
nand UO_66 (O_66,N_3052,N_4792);
nor UO_67 (O_67,N_3538,N_4828);
nor UO_68 (O_68,N_2895,N_4377);
nand UO_69 (O_69,N_2874,N_4926);
nor UO_70 (O_70,N_4898,N_3498);
nor UO_71 (O_71,N_3786,N_4501);
or UO_72 (O_72,N_3182,N_2677);
nor UO_73 (O_73,N_2537,N_2865);
nor UO_74 (O_74,N_3578,N_3706);
nor UO_75 (O_75,N_4419,N_4891);
xor UO_76 (O_76,N_4789,N_3863);
or UO_77 (O_77,N_2769,N_4032);
and UO_78 (O_78,N_2652,N_2544);
nor UO_79 (O_79,N_2715,N_2633);
or UO_80 (O_80,N_4305,N_2634);
and UO_81 (O_81,N_3335,N_4209);
nand UO_82 (O_82,N_4162,N_2577);
and UO_83 (O_83,N_3896,N_3725);
nand UO_84 (O_84,N_4936,N_3901);
nor UO_85 (O_85,N_4731,N_3161);
nand UO_86 (O_86,N_3123,N_4265);
or UO_87 (O_87,N_4808,N_2619);
xor UO_88 (O_88,N_2821,N_2949);
nand UO_89 (O_89,N_3281,N_4211);
or UO_90 (O_90,N_3938,N_3236);
or UO_91 (O_91,N_3857,N_4695);
nor UO_92 (O_92,N_4861,N_3933);
nand UO_93 (O_93,N_4280,N_4291);
nand UO_94 (O_94,N_2705,N_4714);
and UO_95 (O_95,N_3065,N_3115);
and UO_96 (O_96,N_3147,N_3007);
or UO_97 (O_97,N_2515,N_4217);
or UO_98 (O_98,N_4612,N_4566);
nor UO_99 (O_99,N_4996,N_4335);
nand UO_100 (O_100,N_4811,N_4745);
and UO_101 (O_101,N_4744,N_4331);
nor UO_102 (O_102,N_3593,N_4276);
nand UO_103 (O_103,N_3468,N_3241);
and UO_104 (O_104,N_4266,N_3606);
and UO_105 (O_105,N_2534,N_3828);
and UO_106 (O_106,N_3102,N_3544);
nor UO_107 (O_107,N_3977,N_3086);
or UO_108 (O_108,N_2682,N_4883);
nor UO_109 (O_109,N_3628,N_4635);
and UO_110 (O_110,N_2645,N_2830);
xnor UO_111 (O_111,N_4234,N_4819);
or UO_112 (O_112,N_3972,N_4010);
and UO_113 (O_113,N_4641,N_3344);
and UO_114 (O_114,N_3722,N_3239);
and UO_115 (O_115,N_3233,N_3383);
nor UO_116 (O_116,N_4395,N_2561);
or UO_117 (O_117,N_2836,N_2698);
or UO_118 (O_118,N_4825,N_3993);
or UO_119 (O_119,N_4983,N_3723);
nor UO_120 (O_120,N_4235,N_4416);
nand UO_121 (O_121,N_4699,N_4230);
xor UO_122 (O_122,N_4322,N_4297);
nor UO_123 (O_123,N_4074,N_3305);
nand UO_124 (O_124,N_4394,N_3906);
xor UO_125 (O_125,N_3943,N_3278);
nor UO_126 (O_126,N_3313,N_3961);
nor UO_127 (O_127,N_3918,N_3800);
nor UO_128 (O_128,N_3368,N_3249);
and UO_129 (O_129,N_3681,N_4468);
and UO_130 (O_130,N_4489,N_4347);
or UO_131 (O_131,N_2684,N_2680);
xnor UO_132 (O_132,N_4439,N_4730);
and UO_133 (O_133,N_4413,N_4860);
nand UO_134 (O_134,N_3215,N_2548);
nor UO_135 (O_135,N_3780,N_2503);
xor UO_136 (O_136,N_3019,N_4691);
nand UO_137 (O_137,N_2921,N_4311);
or UO_138 (O_138,N_4752,N_4473);
and UO_139 (O_139,N_2969,N_4486);
or UO_140 (O_140,N_4921,N_4421);
or UO_141 (O_141,N_2789,N_4693);
and UO_142 (O_142,N_4940,N_3063);
or UO_143 (O_143,N_3908,N_2636);
and UO_144 (O_144,N_4028,N_2923);
nor UO_145 (O_145,N_3620,N_4319);
or UO_146 (O_146,N_3962,N_4627);
and UO_147 (O_147,N_2917,N_4616);
nor UO_148 (O_148,N_2632,N_4899);
nand UO_149 (O_149,N_4818,N_4762);
nand UO_150 (O_150,N_3139,N_4765);
nand UO_151 (O_151,N_4594,N_2793);
nand UO_152 (O_152,N_4463,N_4794);
nand UO_153 (O_153,N_4990,N_4085);
nor UO_154 (O_154,N_2764,N_4569);
nand UO_155 (O_155,N_3517,N_3661);
nand UO_156 (O_156,N_2777,N_3869);
nand UO_157 (O_157,N_4895,N_3637);
xor UO_158 (O_158,N_4059,N_3599);
nor UO_159 (O_159,N_2980,N_4504);
xor UO_160 (O_160,N_2507,N_2816);
or UO_161 (O_161,N_4120,N_4671);
xor UO_162 (O_162,N_4248,N_4174);
nor UO_163 (O_163,N_3206,N_4452);
xor UO_164 (O_164,N_4259,N_3421);
or UO_165 (O_165,N_4373,N_3046);
nand UO_166 (O_166,N_4650,N_4503);
nand UO_167 (O_167,N_4661,N_4199);
and UO_168 (O_168,N_3787,N_4355);
xor UO_169 (O_169,N_3375,N_2794);
or UO_170 (O_170,N_4649,N_3602);
nand UO_171 (O_171,N_4152,N_2538);
and UO_172 (O_172,N_2525,N_4800);
nor UO_173 (O_173,N_4905,N_4632);
xnor UO_174 (O_174,N_4487,N_4441);
nand UO_175 (O_175,N_3113,N_2811);
and UO_176 (O_176,N_3884,N_2867);
and UO_177 (O_177,N_4494,N_2555);
and UO_178 (O_178,N_4223,N_3893);
nand UO_179 (O_179,N_4807,N_3526);
nand UO_180 (O_180,N_4182,N_2985);
nand UO_181 (O_181,N_3091,N_2942);
xnor UO_182 (O_182,N_4440,N_4884);
nor UO_183 (O_183,N_3428,N_2676);
xor UO_184 (O_184,N_4976,N_2520);
or UO_185 (O_185,N_2912,N_4826);
nand UO_186 (O_186,N_4506,N_4881);
nand UO_187 (O_187,N_3817,N_3084);
nor UO_188 (O_188,N_4270,N_4004);
nand UO_189 (O_189,N_2844,N_2885);
xor UO_190 (O_190,N_4519,N_4520);
nor UO_191 (O_191,N_4845,N_4685);
nor UO_192 (O_192,N_2592,N_4153);
or UO_193 (O_193,N_3229,N_3644);
nand UO_194 (O_194,N_2891,N_2974);
nor UO_195 (O_195,N_3689,N_4717);
and UO_196 (O_196,N_4880,N_2641);
xnor UO_197 (O_197,N_3842,N_3995);
and UO_198 (O_198,N_4068,N_3740);
and UO_199 (O_199,N_2508,N_2630);
xor UO_200 (O_200,N_4037,N_3173);
and UO_201 (O_201,N_3717,N_2510);
and UO_202 (O_202,N_4427,N_3364);
and UO_203 (O_203,N_2755,N_3783);
nor UO_204 (O_204,N_3519,N_4450);
or UO_205 (O_205,N_3440,N_3217);
or UO_206 (O_206,N_4411,N_3353);
and UO_207 (O_207,N_4816,N_3418);
xnor UO_208 (O_208,N_4262,N_4216);
nor UO_209 (O_209,N_4467,N_3210);
nor UO_210 (O_210,N_4885,N_3490);
and UO_211 (O_211,N_3636,N_4034);
or UO_212 (O_212,N_4617,N_3796);
xor UO_213 (O_213,N_3948,N_2742);
and UO_214 (O_214,N_3141,N_2772);
xor UO_215 (O_215,N_3475,N_4306);
nor UO_216 (O_216,N_3219,N_4277);
and UO_217 (O_217,N_4927,N_4433);
and UO_218 (O_218,N_3431,N_3290);
nor UO_219 (O_219,N_3997,N_3039);
xor UO_220 (O_220,N_3479,N_4079);
or UO_221 (O_221,N_4769,N_3396);
or UO_222 (O_222,N_2998,N_4545);
nand UO_223 (O_223,N_4949,N_4061);
or UO_224 (O_224,N_2738,N_4630);
nand UO_225 (O_225,N_3273,N_3002);
or UO_226 (O_226,N_2890,N_4048);
nand UO_227 (O_227,N_4110,N_3784);
and UO_228 (O_228,N_2732,N_4461);
or UO_229 (O_229,N_2603,N_3769);
nor UO_230 (O_230,N_3066,N_4711);
or UO_231 (O_231,N_3565,N_3758);
and UO_232 (O_232,N_3774,N_4901);
or UO_233 (O_233,N_3035,N_3990);
nand UO_234 (O_234,N_4455,N_4090);
nor UO_235 (O_235,N_4829,N_3510);
nand UO_236 (O_236,N_3108,N_4615);
or UO_237 (O_237,N_3128,N_3240);
and UO_238 (O_238,N_3507,N_2568);
or UO_239 (O_239,N_4933,N_3886);
xor UO_240 (O_240,N_3284,N_3365);
nor UO_241 (O_241,N_4655,N_3349);
nand UO_242 (O_242,N_3492,N_4434);
and UO_243 (O_243,N_4304,N_4560);
and UO_244 (O_244,N_2775,N_4823);
or UO_245 (O_245,N_3146,N_2797);
or UO_246 (O_246,N_2884,N_4593);
and UO_247 (O_247,N_3811,N_2767);
nand UO_248 (O_248,N_2748,N_2903);
nor UO_249 (O_249,N_3750,N_2597);
nand UO_250 (O_250,N_4850,N_4273);
nor UO_251 (O_251,N_3540,N_2955);
nand UO_252 (O_252,N_3937,N_3085);
or UO_253 (O_253,N_4172,N_3748);
nand UO_254 (O_254,N_3868,N_4882);
or UO_255 (O_255,N_3727,N_4838);
nor UO_256 (O_256,N_3125,N_4491);
nor UO_257 (O_257,N_4352,N_3562);
nand UO_258 (O_258,N_4620,N_3895);
or UO_259 (O_259,N_4755,N_4220);
or UO_260 (O_260,N_2770,N_4299);
nand UO_261 (O_261,N_4709,N_4796);
nand UO_262 (O_262,N_3225,N_4150);
or UO_263 (O_263,N_2887,N_3595);
nand UO_264 (O_264,N_3742,N_3465);
nand UO_265 (O_265,N_3764,N_4547);
nor UO_266 (O_266,N_3584,N_4718);
and UO_267 (O_267,N_4018,N_3181);
nand UO_268 (O_268,N_3947,N_4167);
or UO_269 (O_269,N_3663,N_3156);
or UO_270 (O_270,N_4626,N_4166);
or UO_271 (O_271,N_3603,N_4228);
nand UO_272 (O_272,N_3770,N_4104);
and UO_273 (O_273,N_4701,N_3978);
and UO_274 (O_274,N_2719,N_3666);
and UO_275 (O_275,N_2857,N_3301);
or UO_276 (O_276,N_2501,N_4025);
nand UO_277 (O_277,N_2751,N_4781);
and UO_278 (O_278,N_4205,N_2876);
and UO_279 (O_279,N_3629,N_3934);
xnor UO_280 (O_280,N_2727,N_3819);
or UO_281 (O_281,N_4683,N_4056);
nand UO_282 (O_282,N_4410,N_3530);
nor UO_283 (O_283,N_4775,N_4047);
or UO_284 (O_284,N_2978,N_2805);
nand UO_285 (O_285,N_2674,N_4571);
or UO_286 (O_286,N_3759,N_3924);
nand UO_287 (O_287,N_3300,N_4645);
xor UO_288 (O_288,N_4245,N_3921);
nor UO_289 (O_289,N_4425,N_4978);
and UO_290 (O_290,N_4662,N_3341);
nand UO_291 (O_291,N_3263,N_4031);
nand UO_292 (O_292,N_4663,N_3931);
and UO_293 (O_293,N_2665,N_3082);
nor UO_294 (O_294,N_3820,N_3822);
and UO_295 (O_295,N_4255,N_3489);
nand UO_296 (O_296,N_3570,N_2588);
or UO_297 (O_297,N_4887,N_4773);
nor UO_298 (O_298,N_3920,N_2661);
nand UO_299 (O_299,N_3148,N_2746);
nor UO_300 (O_300,N_3797,N_3739);
nor UO_301 (O_301,N_3429,N_4062);
or UO_302 (O_302,N_4512,N_2787);
nor UO_303 (O_303,N_3926,N_2820);
and UO_304 (O_304,N_3751,N_4260);
or UO_305 (O_305,N_3928,N_4295);
and UO_306 (O_306,N_3591,N_2915);
or UO_307 (O_307,N_3169,N_2650);
nand UO_308 (O_308,N_4154,N_2516);
or UO_309 (O_309,N_3805,N_3812);
and UO_310 (O_310,N_2908,N_2863);
or UO_311 (O_311,N_2925,N_3726);
and UO_312 (O_312,N_4094,N_3367);
nor UO_313 (O_313,N_4859,N_3729);
nand UO_314 (O_314,N_3903,N_3904);
nand UO_315 (O_315,N_4210,N_3054);
nand UO_316 (O_316,N_4556,N_4852);
and UO_317 (O_317,N_4518,N_2718);
and UO_318 (O_318,N_2892,N_2522);
nand UO_319 (O_319,N_4521,N_4499);
xnor UO_320 (O_320,N_3089,N_4774);
nor UO_321 (O_321,N_3292,N_3466);
xor UO_322 (O_322,N_3747,N_3070);
nand UO_323 (O_323,N_4843,N_3767);
and UO_324 (O_324,N_4833,N_4190);
nor UO_325 (O_325,N_3451,N_4215);
or UO_326 (O_326,N_3274,N_3377);
nand UO_327 (O_327,N_4870,N_4981);
nand UO_328 (O_328,N_2791,N_3112);
and UO_329 (O_329,N_4330,N_2904);
nand UO_330 (O_330,N_3314,N_2968);
nand UO_331 (O_331,N_3163,N_4780);
nor UO_332 (O_332,N_3153,N_3836);
nand UO_333 (O_333,N_3100,N_2801);
nand UO_334 (O_334,N_3700,N_4181);
nor UO_335 (O_335,N_2666,N_2509);
xnor UO_336 (O_336,N_3563,N_3162);
nand UO_337 (O_337,N_3358,N_2556);
nand UO_338 (O_338,N_2889,N_4376);
nand UO_339 (O_339,N_2685,N_4532);
or UO_340 (O_340,N_4464,N_2675);
and UO_341 (O_341,N_4257,N_3197);
or UO_342 (O_342,N_3230,N_3971);
and UO_343 (O_343,N_4993,N_3539);
or UO_344 (O_344,N_2786,N_4586);
and UO_345 (O_345,N_4170,N_4442);
or UO_346 (O_346,N_4126,N_4343);
xor UO_347 (O_347,N_3804,N_3254);
and UO_348 (O_348,N_3376,N_4931);
nand UO_349 (O_349,N_2713,N_4495);
xor UO_350 (O_350,N_4366,N_4398);
nand UO_351 (O_351,N_2704,N_3191);
and UO_352 (O_352,N_3175,N_3974);
and UO_353 (O_353,N_4131,N_4036);
nand UO_354 (O_354,N_2852,N_3835);
nand UO_355 (O_355,N_3627,N_3350);
or UO_356 (O_356,N_4317,N_4516);
nor UO_357 (O_357,N_4920,N_3198);
nor UO_358 (O_358,N_3605,N_3260);
nor UO_359 (O_359,N_3772,N_4757);
and UO_360 (O_360,N_4783,N_3516);
and UO_361 (O_361,N_4862,N_4301);
nor UO_362 (O_362,N_4514,N_4528);
and UO_363 (O_363,N_2993,N_3504);
and UO_364 (O_364,N_3071,N_3487);
xnor UO_365 (O_365,N_3941,N_2973);
or UO_366 (O_366,N_2567,N_3790);
or UO_367 (O_367,N_3058,N_4146);
and UO_368 (O_368,N_4091,N_4239);
nand UO_369 (O_369,N_3132,N_4477);
or UO_370 (O_370,N_4788,N_2513);
xnor UO_371 (O_371,N_2553,N_4278);
nor UO_372 (O_372,N_3386,N_4053);
nor UO_373 (O_373,N_3524,N_3773);
and UO_374 (O_374,N_4965,N_4543);
nor UO_375 (O_375,N_3242,N_2872);
or UO_376 (O_376,N_4194,N_4348);
and UO_377 (O_377,N_2683,N_2771);
or UO_378 (O_378,N_3752,N_3731);
nor UO_379 (O_379,N_3030,N_4734);
nor UO_380 (O_380,N_3709,N_2984);
and UO_381 (O_381,N_2651,N_2730);
or UO_382 (O_382,N_3060,N_2621);
and UO_383 (O_383,N_3411,N_4081);
and UO_384 (O_384,N_2815,N_3261);
and UO_385 (O_385,N_2747,N_3009);
and UO_386 (O_386,N_4873,N_3207);
or UO_387 (O_387,N_3916,N_3159);
or UO_388 (O_388,N_4607,N_4984);
and UO_389 (O_389,N_3107,N_2551);
nor UO_390 (O_390,N_3469,N_2813);
nand UO_391 (O_391,N_3604,N_3378);
nor UO_392 (O_392,N_3315,N_4707);
or UO_393 (O_393,N_4027,N_3213);
xor UO_394 (O_394,N_3915,N_4367);
nor UO_395 (O_395,N_3684,N_2744);
nand UO_396 (O_396,N_2950,N_4431);
and UO_397 (O_397,N_3279,N_2807);
and UO_398 (O_398,N_3875,N_3856);
and UO_399 (O_399,N_3187,N_4574);
nand UO_400 (O_400,N_3659,N_3481);
nor UO_401 (O_401,N_4269,N_4318);
nand UO_402 (O_402,N_4777,N_3395);
xnor UO_403 (O_403,N_3190,N_4705);
and UO_404 (O_404,N_4137,N_4346);
and UO_405 (O_405,N_4122,N_3050);
or UO_406 (O_406,N_4537,N_3515);
nor UO_407 (O_407,N_2589,N_3497);
xor UO_408 (O_408,N_3354,N_4557);
nor UO_409 (O_409,N_2860,N_4896);
nand UO_410 (O_410,N_4533,N_4307);
or UO_411 (O_411,N_4975,N_2907);
or UO_412 (O_412,N_2778,N_3525);
or UO_413 (O_413,N_3196,N_2833);
or UO_414 (O_414,N_3037,N_2785);
xnor UO_415 (O_415,N_2843,N_4353);
nand UO_416 (O_416,N_3608,N_3357);
nand UO_417 (O_417,N_4193,N_4761);
nand UO_418 (O_418,N_2724,N_2947);
or UO_419 (O_419,N_2624,N_4893);
or UO_420 (O_420,N_4665,N_2875);
nor UO_421 (O_421,N_3360,N_4876);
xnor UO_422 (O_422,N_4482,N_3068);
and UO_423 (O_423,N_4903,N_2913);
nor UO_424 (O_424,N_3596,N_3929);
or UO_425 (O_425,N_2604,N_4836);
nand UO_426 (O_426,N_3951,N_3446);
nand UO_427 (O_427,N_4760,N_3503);
nor UO_428 (O_428,N_4737,N_4180);
or UO_429 (O_429,N_3754,N_3905);
or UO_430 (O_430,N_2847,N_3444);
or UO_431 (O_431,N_3178,N_3710);
and UO_432 (O_432,N_4928,N_3621);
nand UO_433 (O_433,N_4856,N_4888);
xor UO_434 (O_434,N_4359,N_3445);
or UO_435 (O_435,N_4723,N_4525);
xnor UO_436 (O_436,N_2552,N_3509);
and UO_437 (O_437,N_2877,N_2901);
and UO_438 (O_438,N_2536,N_3144);
nand UO_439 (O_439,N_2750,N_4559);
nor UO_440 (O_440,N_4498,N_3803);
nor UO_441 (O_441,N_4681,N_4517);
or UO_442 (O_442,N_3435,N_4333);
or UO_443 (O_443,N_2699,N_2966);
nor UO_444 (O_444,N_4957,N_4328);
nand UO_445 (O_445,N_2723,N_3474);
xor UO_446 (O_446,N_3101,N_4035);
or UO_447 (O_447,N_3871,N_2618);
nand UO_448 (O_448,N_2714,N_3841);
nand UO_449 (O_449,N_3576,N_3496);
nand UO_450 (O_450,N_4675,N_3061);
nand UO_451 (O_451,N_3042,N_4916);
nand UO_452 (O_452,N_3981,N_4758);
nand UO_453 (O_453,N_3342,N_2753);
nor UO_454 (O_454,N_3359,N_3398);
nor UO_455 (O_455,N_3013,N_4656);
nor UO_456 (O_456,N_4369,N_4793);
xnor UO_457 (O_457,N_2871,N_3130);
nand UO_458 (O_458,N_3687,N_4982);
and UO_459 (O_459,N_3265,N_4290);
nand UO_460 (O_460,N_2639,N_4698);
and UO_461 (O_461,N_2888,N_2703);
nor UO_462 (O_462,N_2943,N_3216);
nand UO_463 (O_463,N_4344,N_2626);
or UO_464 (O_464,N_3051,N_3164);
and UO_465 (O_465,N_3865,N_2834);
nand UO_466 (O_466,N_4100,N_4603);
nor UO_467 (O_467,N_4357,N_4351);
nor UO_468 (O_468,N_4639,N_3590);
or UO_469 (O_469,N_2758,N_3542);
nor UO_470 (O_470,N_3186,N_3645);
nor UO_471 (O_471,N_3083,N_2878);
and UO_472 (O_472,N_3892,N_2879);
nand UO_473 (O_473,N_2870,N_3976);
or UO_474 (O_474,N_4164,N_4791);
nor UO_475 (O_475,N_4358,N_3791);
xnor UO_476 (O_476,N_4033,N_3202);
nor UO_477 (O_477,N_3588,N_3880);
nand UO_478 (O_478,N_3553,N_3040);
nand UO_479 (O_479,N_2547,N_3294);
or UO_480 (O_480,N_3053,N_4790);
or UO_481 (O_481,N_2600,N_2965);
and UO_482 (O_482,N_2840,N_4247);
nor UO_483 (O_483,N_4125,N_2694);
nor UO_484 (O_484,N_2505,N_3380);
nor UO_485 (O_485,N_4653,N_3160);
nand UO_486 (O_486,N_3408,N_3399);
nand UO_487 (O_487,N_3894,N_4721);
nor UO_488 (O_488,N_3127,N_4422);
nand UO_489 (O_489,N_4941,N_4904);
nand UO_490 (O_490,N_3646,N_3373);
nor UO_491 (O_491,N_4659,N_2550);
or UO_492 (O_492,N_2735,N_4704);
nor UO_493 (O_493,N_2712,N_4821);
nor UO_494 (O_494,N_4488,N_4314);
and UO_495 (O_495,N_4858,N_4140);
nand UO_496 (O_496,N_4454,N_4599);
or UO_497 (O_497,N_4544,N_3379);
nor UO_498 (O_498,N_3317,N_3308);
nor UO_499 (O_499,N_4017,N_2799);
nor UO_500 (O_500,N_2740,N_2627);
xnor UO_501 (O_501,N_3103,N_2851);
nand UO_502 (O_502,N_2832,N_3555);
and UO_503 (O_503,N_4509,N_3478);
nor UO_504 (O_504,N_2972,N_2842);
xor UO_505 (O_505,N_2642,N_4784);
or UO_506 (O_506,N_4404,N_3057);
nand UO_507 (O_507,N_2776,N_3810);
or UO_508 (O_508,N_3522,N_2528);
nand UO_509 (O_509,N_2681,N_4673);
and UO_510 (O_510,N_2982,N_3208);
nor UO_511 (O_511,N_4083,N_4710);
nor UO_512 (O_512,N_3778,N_3321);
and UO_513 (O_513,N_4141,N_4040);
nand UO_514 (O_514,N_2563,N_2924);
or UO_515 (O_515,N_3534,N_3989);
or UO_516 (O_516,N_4143,N_2996);
nand UO_517 (O_517,N_4470,N_4308);
xor UO_518 (O_518,N_3165,N_3888);
xor UO_519 (O_519,N_2930,N_4628);
and UO_520 (O_520,N_4387,N_3195);
xnor UO_521 (O_521,N_3419,N_4298);
xnor UO_522 (O_522,N_4407,N_4953);
or UO_523 (O_523,N_4383,N_3930);
xor UO_524 (O_524,N_2687,N_3942);
nor UO_525 (O_525,N_2602,N_3238);
or UO_526 (O_526,N_4015,N_3406);
xnor UO_527 (O_527,N_4508,N_4827);
or UO_528 (O_528,N_3716,N_4657);
nor UO_529 (O_529,N_3462,N_4368);
or UO_530 (O_530,N_3276,N_2518);
nand UO_531 (O_531,N_3697,N_2800);
and UO_532 (O_532,N_4561,N_3450);
or UO_533 (O_533,N_4565,N_4589);
or UO_534 (O_534,N_2517,N_4197);
xor UO_535 (O_535,N_4138,N_2691);
nand UO_536 (O_536,N_4332,N_4142);
and UO_537 (O_537,N_4233,N_3374);
nor UO_538 (O_538,N_2959,N_4097);
nor UO_539 (O_539,N_3133,N_2669);
nor UO_540 (O_540,N_3789,N_2565);
nor UO_541 (O_541,N_3318,N_2927);
nand UO_542 (O_542,N_2902,N_3703);
nor UO_543 (O_543,N_4251,N_4240);
and UO_544 (O_544,N_2975,N_4767);
xnor UO_545 (O_545,N_3438,N_4282);
or UO_546 (O_546,N_3719,N_3957);
and UO_547 (O_547,N_4189,N_3416);
or UO_548 (O_548,N_3320,N_4510);
nand UO_549 (O_549,N_2873,N_4252);
nand UO_550 (O_550,N_2859,N_4658);
nor UO_551 (O_551,N_4712,N_4244);
nand UO_552 (O_552,N_2672,N_3756);
and UO_553 (O_553,N_4803,N_3807);
and UO_554 (O_554,N_3347,N_3129);
nand UO_555 (O_555,N_4412,N_2995);
nand UO_556 (O_556,N_3741,N_4667);
and UO_557 (O_557,N_3762,N_3439);
nand UO_558 (O_558,N_3081,N_2848);
nor UO_559 (O_559,N_4437,N_3425);
nor UO_560 (O_560,N_4249,N_4073);
or UO_561 (O_561,N_4585,N_3902);
nor UO_562 (O_562,N_3724,N_3702);
nor UO_563 (O_563,N_3964,N_3417);
nand UO_564 (O_564,N_3485,N_3858);
xnor UO_565 (O_565,N_2956,N_2803);
nand UO_566 (O_566,N_3569,N_3275);
xnor UO_567 (O_567,N_4660,N_2845);
and UO_568 (O_568,N_2502,N_4600);
nand UO_569 (O_569,N_3064,N_3323);
or UO_570 (O_570,N_3956,N_3174);
nor UO_571 (O_571,N_2941,N_3832);
or UO_572 (O_572,N_3744,N_4005);
or UO_573 (O_573,N_4742,N_3179);
nand UO_574 (O_574,N_2545,N_4988);
and UO_575 (O_575,N_3619,N_4356);
or UO_576 (O_576,N_3069,N_3184);
nand UO_577 (O_577,N_4575,N_3297);
nor UO_578 (O_578,N_3149,N_4436);
nor UO_579 (O_579,N_4550,N_4636);
nand UO_580 (O_580,N_3000,N_3949);
nor UO_581 (O_581,N_4496,N_4229);
nand UO_582 (O_582,N_2728,N_3733);
or UO_583 (O_583,N_4706,N_3407);
nor UO_584 (O_584,N_2660,N_2614);
nor UO_585 (O_585,N_4484,N_2808);
nand UO_586 (O_586,N_3873,N_2839);
xor UO_587 (O_587,N_3543,N_3150);
nor UO_588 (O_588,N_3970,N_4149);
and UO_589 (O_589,N_4001,N_2928);
and UO_590 (O_590,N_3521,N_2596);
nor UO_591 (O_591,N_3624,N_4728);
and UO_592 (O_592,N_3456,N_2529);
and UO_593 (O_593,N_4992,N_3609);
or UO_594 (O_594,N_4804,N_4271);
and UO_595 (O_595,N_3586,N_2899);
nand UO_596 (O_596,N_3757,N_4581);
and UO_597 (O_597,N_3001,N_4527);
or UO_598 (O_598,N_4392,N_4625);
and UO_599 (O_599,N_3911,N_4321);
or UO_600 (O_600,N_4834,N_3499);
nand UO_601 (O_601,N_3477,N_3582);
or UO_602 (O_602,N_3707,N_4523);
xnor UO_603 (O_603,N_3912,N_4553);
xor UO_604 (O_604,N_3736,N_3909);
or UO_605 (O_605,N_4610,N_3671);
and UO_606 (O_606,N_4084,N_4336);
nand UO_607 (O_607,N_2906,N_4759);
and UO_608 (O_608,N_3612,N_4349);
nand UO_609 (O_609,N_4577,N_4123);
nor UO_610 (O_610,N_3234,N_4093);
nand UO_611 (O_611,N_4592,N_3316);
nor UO_612 (O_612,N_3256,N_4875);
or UO_613 (O_613,N_4866,N_2948);
and UO_614 (O_614,N_4570,N_2702);
nor UO_615 (O_615,N_4716,N_4218);
nand UO_616 (O_616,N_4095,N_3589);
xor UO_617 (O_617,N_4175,N_4606);
and UO_618 (O_618,N_4908,N_2514);
nor UO_619 (O_619,N_2546,N_2541);
nor UO_620 (O_620,N_4379,N_4914);
xor UO_621 (O_621,N_3333,N_4086);
xor UO_622 (O_622,N_4985,N_4872);
or UO_623 (O_623,N_4261,N_2796);
nand UO_624 (O_624,N_4372,N_4444);
or UO_625 (O_625,N_3319,N_4809);
and UO_626 (O_626,N_2569,N_3043);
and UO_627 (O_627,N_3243,N_2601);
or UO_628 (O_628,N_3214,N_4912);
nand UO_629 (O_629,N_2706,N_3420);
nor UO_630 (O_630,N_4584,N_4651);
nand UO_631 (O_631,N_4077,N_3355);
xnor UO_632 (O_632,N_3382,N_4009);
and UO_633 (O_633,N_4350,N_4088);
or UO_634 (O_634,N_4323,N_3463);
nor UO_635 (O_635,N_2954,N_3346);
nor UO_636 (O_636,N_3914,N_4483);
nor UO_637 (O_637,N_4171,N_4670);
and UO_638 (O_638,N_4012,N_4241);
or UO_639 (O_639,N_3531,N_3825);
xnor UO_640 (O_640,N_4638,N_4580);
or UO_641 (O_641,N_4329,N_2812);
and UO_642 (O_642,N_4715,N_4371);
or UO_643 (O_643,N_3105,N_3782);
nor UO_644 (O_644,N_2919,N_3728);
xor UO_645 (O_645,N_4853,N_4644);
nand UO_646 (O_646,N_3987,N_2997);
and UO_647 (O_647,N_2909,N_2762);
nor UO_648 (O_648,N_3996,N_4708);
nor UO_649 (O_649,N_3289,N_2609);
nand UO_650 (O_650,N_3221,N_3511);
xnor UO_651 (O_651,N_3372,N_4854);
nor UO_652 (O_652,N_4943,N_2649);
and UO_653 (O_653,N_2578,N_4102);
nor UO_654 (O_654,N_4363,N_4285);
nor UO_655 (O_655,N_2574,N_3557);
nand UO_656 (O_656,N_2689,N_4864);
nand UO_657 (O_657,N_4114,N_4424);
nor UO_658 (O_658,N_4406,N_2585);
and UO_659 (O_659,N_4155,N_3746);
and UO_660 (O_660,N_3258,N_3984);
nand UO_661 (O_661,N_4733,N_3658);
nand UO_662 (O_662,N_3668,N_3891);
nor UO_663 (O_663,N_3662,N_4720);
nor UO_664 (O_664,N_4751,N_2659);
and UO_665 (O_665,N_4886,N_4922);
nor UO_666 (O_666,N_3592,N_2524);
nor UO_667 (O_667,N_3502,N_4370);
and UO_668 (O_668,N_2829,N_4732);
nor UO_669 (O_669,N_2620,N_2530);
nand UO_670 (O_670,N_4502,N_2654);
xor UO_671 (O_671,N_3194,N_2782);
or UO_672 (O_672,N_2850,N_3991);
nor UO_673 (O_673,N_4341,N_3674);
nand UO_674 (O_674,N_3111,N_4568);
nor UO_675 (O_675,N_4997,N_4296);
xor UO_676 (O_676,N_4739,N_2752);
and UO_677 (O_677,N_3486,N_3006);
xnor UO_678 (O_678,N_4459,N_3074);
or UO_679 (O_679,N_4049,N_4030);
nand UO_680 (O_680,N_3090,N_3776);
and UO_681 (O_681,N_3654,N_2757);
nand UO_682 (O_682,N_3890,N_4633);
nor UO_683 (O_683,N_2590,N_3324);
and UO_684 (O_684,N_3322,N_4316);
nand UO_685 (O_685,N_4445,N_3337);
and UO_686 (O_686,N_4096,N_4263);
nor UO_687 (O_687,N_3032,N_4132);
or UO_688 (O_688,N_2608,N_3632);
and UO_689 (O_689,N_3983,N_4178);
or UO_690 (O_690,N_2754,N_3270);
nand UO_691 (O_691,N_3025,N_3675);
nand UO_692 (O_692,N_2900,N_4400);
or UO_693 (O_693,N_3459,N_4911);
nand UO_694 (O_694,N_3587,N_3222);
or UO_695 (O_695,N_2656,N_4753);
and UO_696 (O_696,N_4841,N_2564);
nor UO_697 (O_697,N_3080,N_2664);
and UO_698 (O_698,N_4423,N_3134);
nand UO_699 (O_699,N_3676,N_4481);
and UO_700 (O_700,N_3271,N_3348);
nand UO_701 (O_701,N_3613,N_2554);
or UO_702 (O_702,N_2944,N_4972);
nand UO_703 (O_703,N_4231,N_2655);
nor UO_704 (O_704,N_4226,N_3622);
nor UO_705 (O_705,N_4458,N_3340);
nor UO_706 (O_706,N_3343,N_4674);
xor UO_707 (O_707,N_3641,N_4057);
xnor UO_708 (O_708,N_2605,N_2743);
and UO_709 (O_709,N_3356,N_2562);
or UO_710 (O_710,N_4989,N_3433);
nand UO_711 (O_711,N_3096,N_3166);
or UO_712 (O_712,N_2731,N_2814);
and UO_713 (O_713,N_4105,N_3585);
or UO_714 (O_714,N_4894,N_3119);
or UO_715 (O_715,N_3859,N_3917);
nand UO_716 (O_716,N_4378,N_3688);
or UO_717 (O_717,N_3137,N_4106);
nand UO_718 (O_718,N_2690,N_3533);
and UO_719 (O_719,N_3038,N_2933);
or UO_720 (O_720,N_4986,N_2893);
and UO_721 (O_721,N_3110,N_3839);
nor UO_722 (O_722,N_4951,N_2533);
or UO_723 (O_723,N_3633,N_3253);
or UO_724 (O_724,N_3616,N_4500);
and UO_725 (O_725,N_4429,N_3980);
nor UO_726 (O_726,N_4448,N_3143);
nor UO_727 (O_727,N_4325,N_3642);
nor UO_728 (O_728,N_3464,N_3003);
nor UO_729 (O_729,N_3985,N_4847);
and UO_730 (O_730,N_3437,N_3712);
xor UO_731 (O_731,N_3872,N_3955);
or UO_732 (O_732,N_3614,N_3775);
and UO_733 (O_733,N_3651,N_4938);
or UO_734 (O_734,N_2810,N_3680);
or UO_735 (O_735,N_3882,N_3704);
nand UO_736 (O_736,N_3152,N_3200);
xnor UO_737 (O_737,N_2716,N_2610);
nand UO_738 (O_738,N_3185,N_4157);
and UO_739 (O_739,N_3299,N_4750);
and UO_740 (O_740,N_3443,N_4339);
nor UO_741 (O_741,N_3601,N_2881);
nor UO_742 (O_742,N_4113,N_2802);
xor UO_743 (O_743,N_2701,N_4242);
and UO_744 (O_744,N_4042,N_2929);
or UO_745 (O_745,N_4365,N_2882);
or UO_746 (O_746,N_3142,N_3389);
nor UO_747 (O_747,N_3325,N_4475);
nor UO_748 (O_748,N_2521,N_3493);
or UO_749 (O_749,N_3946,N_2898);
xor UO_750 (O_750,N_3291,N_4806);
or UO_751 (O_751,N_3639,N_4389);
nand UO_752 (O_752,N_4063,N_3180);
nor UO_753 (O_753,N_3898,N_3877);
or UO_754 (O_754,N_4743,N_4124);
and UO_755 (O_755,N_4478,N_4932);
nor UO_756 (O_756,N_4026,N_4832);
and UO_757 (O_757,N_2773,N_3939);
nor UO_758 (O_758,N_4456,N_2749);
nand UO_759 (O_759,N_4109,N_4168);
nor UO_760 (O_760,N_3925,N_3795);
xnor UO_761 (O_761,N_3870,N_2963);
nand UO_762 (O_762,N_4619,N_4719);
or UO_763 (O_763,N_4337,N_3682);
nand UO_764 (O_764,N_4212,N_3304);
nor UO_765 (O_765,N_2519,N_3695);
nor UO_766 (O_766,N_3827,N_3735);
or UO_767 (O_767,N_4207,N_3737);
nor UO_768 (O_768,N_3850,N_3548);
nand UO_769 (O_769,N_3512,N_4111);
nor UO_770 (O_770,N_2696,N_4013);
or UO_771 (O_771,N_4507,N_3136);
nand UO_772 (O_772,N_4970,N_3552);
xor UO_773 (O_773,N_4485,N_3480);
nor UO_774 (O_774,N_4726,N_3079);
nand UO_775 (O_775,N_4254,N_4686);
nor UO_776 (O_776,N_3247,N_4801);
nor UO_777 (O_777,N_4115,N_3763);
or UO_778 (O_778,N_2841,N_4006);
nor UO_779 (O_779,N_2837,N_4766);
or UO_780 (O_780,N_2759,N_2994);
and UO_781 (O_781,N_3014,N_4740);
or UO_782 (O_782,N_3899,N_4799);
and UO_783 (O_783,N_2709,N_3573);
and UO_784 (O_784,N_3617,N_3568);
or UO_785 (O_785,N_4381,N_3283);
nand UO_786 (O_786,N_4583,N_4183);
and UO_787 (O_787,N_4768,N_4320);
and UO_788 (O_788,N_3945,N_4121);
nand UO_789 (O_789,N_4179,N_3384);
nor UO_790 (O_790,N_3392,N_2795);
nor UO_791 (O_791,N_3366,N_3262);
nand UO_792 (O_792,N_3814,N_3237);
nand UO_793 (O_793,N_3913,N_3171);
and UO_794 (O_794,N_4950,N_4967);
and UO_795 (O_795,N_3311,N_2739);
nand UO_796 (O_796,N_4426,N_3843);
or UO_797 (O_797,N_4472,N_4050);
nand UO_798 (O_798,N_4169,N_4493);
nand UO_799 (O_799,N_4253,N_3205);
and UO_800 (O_800,N_3168,N_2708);
and UO_801 (O_801,N_3556,N_4186);
nand UO_802 (O_802,N_4003,N_3808);
nand UO_803 (O_803,N_3028,N_3600);
nand UO_804 (O_804,N_3250,N_4408);
nand UO_805 (O_805,N_4554,N_3683);
nand UO_806 (O_806,N_4315,N_4388);
nand UO_807 (O_807,N_3029,N_3549);
or UO_808 (O_808,N_3176,N_3809);
xnor UO_809 (O_809,N_3618,N_4968);
and UO_810 (O_810,N_4151,N_4129);
or UO_811 (O_811,N_4072,N_3883);
and UO_812 (O_812,N_4770,N_4579);
nor UO_813 (O_813,N_3594,N_3011);
nor UO_814 (O_814,N_3708,N_4310);
or UO_815 (O_815,N_4438,N_4979);
nand UO_816 (O_816,N_3864,N_3986);
xnor UO_817 (O_817,N_4831,N_4192);
nand UO_818 (O_818,N_3436,N_4646);
and UO_819 (O_819,N_4535,N_4380);
nor UO_820 (O_820,N_4326,N_4402);
or UO_821 (O_821,N_2946,N_3919);
nor UO_822 (O_822,N_4889,N_3109);
nor UO_823 (O_823,N_3227,N_2598);
and UO_824 (O_824,N_4135,N_3761);
nor UO_825 (O_825,N_4994,N_3295);
nand UO_826 (O_826,N_2527,N_3847);
or UO_827 (O_827,N_4576,N_3743);
nand UO_828 (O_828,N_3779,N_3935);
or UO_829 (O_829,N_2583,N_4952);
nor UO_830 (O_830,N_3494,N_3583);
nand UO_831 (O_831,N_2622,N_3482);
or UO_832 (O_832,N_4044,N_3701);
xor UO_833 (O_833,N_4672,N_3610);
nor UO_834 (O_834,N_4112,N_4292);
nor UO_835 (O_835,N_3501,N_2586);
nand UO_836 (O_836,N_4956,N_2670);
xnor UO_837 (O_837,N_2710,N_4684);
nor UO_838 (O_838,N_3288,N_3495);
and UO_839 (O_839,N_4551,N_4161);
or UO_840 (O_840,N_3969,N_3649);
and UO_841 (O_841,N_4624,N_3307);
or UO_842 (O_842,N_3777,N_3430);
nand UO_843 (O_843,N_3634,N_4631);
nor UO_844 (O_844,N_4785,N_2667);
nor UO_845 (O_845,N_4618,N_3404);
xnor UO_846 (O_846,N_3330,N_3854);
nand UO_847 (O_847,N_3255,N_3077);
nand UO_848 (O_848,N_3834,N_4810);
and UO_849 (O_849,N_3223,N_3167);
and UO_850 (O_850,N_3794,N_3400);
or UO_851 (O_851,N_3327,N_3923);
nor UO_852 (O_852,N_4692,N_4842);
xnor UO_853 (O_853,N_4250,N_3059);
nor UO_854 (O_854,N_3293,N_2607);
and UO_855 (O_855,N_4476,N_4652);
nand UO_856 (O_856,N_4345,N_2798);
nand UO_857 (O_857,N_4214,N_2856);
and UO_858 (O_858,N_3874,N_3900);
nand UO_859 (O_859,N_2894,N_3615);
and UO_860 (O_860,N_4185,N_3523);
xnor UO_861 (O_861,N_4268,N_4148);
or UO_862 (O_862,N_4069,N_4591);
or UO_863 (O_863,N_3846,N_3696);
nand UO_864 (O_864,N_4964,N_3199);
nor UO_865 (O_865,N_4947,N_4173);
nand UO_866 (O_866,N_2951,N_3306);
nand UO_867 (O_867,N_3020,N_4910);
or UO_868 (O_868,N_4382,N_2958);
xor UO_869 (O_869,N_4682,N_3635);
and UO_870 (O_870,N_3280,N_2594);
and UO_871 (O_871,N_4338,N_4065);
or UO_872 (O_872,N_2725,N_4696);
nor UO_873 (O_873,N_4764,N_3048);
nor UO_874 (O_874,N_3760,N_3381);
nor UO_875 (O_875,N_4582,N_4676);
nor UO_876 (O_876,N_4902,N_3988);
or UO_877 (O_877,N_4830,N_2981);
nand UO_878 (O_878,N_3932,N_4414);
xnor UO_879 (O_879,N_4342,N_3867);
nand UO_880 (O_880,N_3940,N_4449);
xor UO_881 (O_881,N_3830,N_4469);
or UO_882 (O_882,N_4300,N_2549);
nor UO_883 (O_883,N_3220,N_4536);
nor UO_884 (O_884,N_3434,N_3145);
nand UO_885 (O_885,N_3298,N_2591);
nand UO_886 (O_886,N_4937,N_3402);
nor UO_887 (O_887,N_3897,N_3845);
or UO_888 (O_888,N_4729,N_4479);
or UO_889 (O_889,N_4039,N_3785);
or UO_890 (O_890,N_4225,N_2939);
nand UO_891 (O_891,N_2916,N_3401);
and UO_892 (O_892,N_3004,N_4490);
nor UO_893 (O_893,N_2613,N_4955);
or UO_894 (O_894,N_4689,N_2760);
nor UO_895 (O_895,N_3118,N_2976);
nand UO_896 (O_896,N_3561,N_3979);
xnor UO_897 (O_897,N_2542,N_4432);
nand UO_898 (O_898,N_3579,N_2761);
and UO_899 (O_899,N_4530,N_3218);
nor UO_900 (O_900,N_3094,N_2989);
or UO_901 (O_901,N_4877,N_3765);
xor UO_902 (O_902,N_2804,N_3470);
or UO_903 (O_903,N_3572,N_3455);
or UO_904 (O_904,N_4694,N_3887);
and UO_905 (O_905,N_2576,N_4907);
or UO_906 (O_906,N_4640,N_3669);
or UO_907 (O_907,N_3853,N_4654);
or UO_908 (O_908,N_3881,N_3768);
nor UO_909 (O_909,N_4224,N_2587);
nand UO_910 (O_910,N_4058,N_3550);
xor UO_911 (O_911,N_3371,N_2695);
nor UO_912 (O_912,N_3677,N_4060);
nor UO_913 (O_913,N_3566,N_4595);
or UO_914 (O_914,N_4014,N_3514);
nor UO_915 (O_915,N_3267,N_4000);
nand UO_916 (O_916,N_4451,N_3334);
nor UO_917 (O_917,N_4772,N_3546);
nor UO_918 (O_918,N_3959,N_3792);
nor UO_919 (O_919,N_4690,N_4396);
nand UO_920 (O_920,N_3678,N_3026);
or UO_921 (O_921,N_4022,N_4418);
nor UO_922 (O_922,N_4385,N_4541);
nand UO_923 (O_923,N_4145,N_3093);
nand UO_924 (O_924,N_2595,N_3033);
and UO_925 (O_925,N_2615,N_4679);
and UO_926 (O_926,N_3922,N_4851);
nor UO_927 (O_927,N_3698,N_4374);
nand UO_928 (O_928,N_3189,N_4364);
nor UO_929 (O_929,N_4573,N_3818);
or UO_930 (O_930,N_4643,N_2827);
xor UO_931 (O_931,N_4814,N_3580);
or UO_932 (O_932,N_4127,N_4897);
nand UO_933 (O_933,N_4159,N_3802);
and UO_934 (O_934,N_3268,N_3170);
nand UO_935 (O_935,N_2631,N_3564);
and UO_936 (O_936,N_3491,N_3005);
xnor UO_937 (O_937,N_3257,N_4139);
or UO_938 (O_938,N_4688,N_4611);
nor UO_939 (O_939,N_2964,N_4812);
or UO_940 (O_940,N_4588,N_2606);
or UO_941 (O_941,N_4163,N_2531);
or UO_942 (O_942,N_4697,N_4598);
nor UO_943 (O_943,N_4457,N_2617);
or UO_944 (O_944,N_4778,N_4309);
nor UO_945 (O_945,N_2938,N_2657);
nand UO_946 (O_946,N_3224,N_3866);
and UO_947 (O_947,N_3138,N_4935);
and UO_948 (O_948,N_4909,N_3056);
nand UO_949 (O_949,N_3211,N_4279);
nand UO_950 (O_950,N_4605,N_3536);
nand UO_951 (O_951,N_3104,N_2897);
xnor UO_952 (O_952,N_4409,N_2977);
and UO_953 (O_953,N_3657,N_2673);
xnor UO_954 (O_954,N_2920,N_4294);
or UO_955 (O_955,N_3966,N_2858);
nor UO_956 (O_956,N_3114,N_3771);
xor UO_957 (O_957,N_2935,N_4542);
nor UO_958 (O_958,N_3575,N_4634);
or UO_959 (O_959,N_3518,N_4966);
or UO_960 (O_960,N_2763,N_3212);
nor UO_961 (O_961,N_4971,N_3303);
or UO_962 (O_962,N_4906,N_4863);
nor UO_963 (O_963,N_2557,N_3155);
or UO_964 (O_964,N_4749,N_4078);
and UO_965 (O_965,N_4219,N_3266);
or UO_966 (O_966,N_3055,N_4497);
nand UO_967 (O_967,N_4103,N_4590);
or UO_968 (O_968,N_3862,N_2540);
and UO_969 (O_969,N_4648,N_2937);
nand UO_970 (O_970,N_4202,N_4664);
nor UO_971 (O_971,N_4052,N_4196);
and UO_972 (O_972,N_4522,N_4540);
and UO_973 (O_973,N_4954,N_2500);
xnor UO_974 (O_974,N_4563,N_3844);
nor UO_975 (O_975,N_4066,N_2988);
or UO_976 (O_976,N_4176,N_4763);
or UO_977 (O_977,N_2637,N_3088);
or UO_978 (O_978,N_2717,N_3286);
nand UO_979 (O_979,N_3749,N_2864);
nor UO_980 (O_980,N_3183,N_4391);
nand UO_981 (O_981,N_4958,N_4213);
and UO_982 (O_982,N_4401,N_4546);
or UO_983 (O_983,N_3816,N_3351);
or UO_984 (O_984,N_3581,N_3473);
nand UO_985 (O_985,N_2662,N_3448);
xor UO_986 (O_986,N_4415,N_3547);
nand UO_987 (O_987,N_4869,N_2962);
and UO_988 (O_988,N_4969,N_3528);
and UO_989 (O_989,N_3449,N_3656);
nor UO_990 (O_990,N_2823,N_4403);
nand UO_991 (O_991,N_4107,N_4480);
or UO_992 (O_992,N_4865,N_2961);
or UO_993 (O_993,N_4198,N_4917);
xnor UO_994 (O_994,N_2896,N_3513);
xnor UO_995 (O_995,N_2736,N_4963);
xnor UO_996 (O_996,N_3410,N_4835);
nand UO_997 (O_997,N_2854,N_4837);
or UO_998 (O_998,N_4128,N_3647);
or UO_999 (O_999,N_3648,N_4258);
endmodule