module basic_500_3000_500_3_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_429,In_49);
and U1 (N_1,In_340,In_443);
xor U2 (N_2,In_133,In_334);
nor U3 (N_3,In_281,In_204);
and U4 (N_4,In_75,In_390);
nand U5 (N_5,In_162,In_243);
or U6 (N_6,In_42,In_293);
or U7 (N_7,In_471,In_438);
nor U8 (N_8,In_168,In_160);
or U9 (N_9,In_9,In_86);
nor U10 (N_10,In_360,In_383);
nor U11 (N_11,In_172,In_402);
or U12 (N_12,In_147,In_108);
or U13 (N_13,In_267,In_131);
or U14 (N_14,In_489,In_374);
nand U15 (N_15,In_241,In_183);
and U16 (N_16,In_182,In_109);
or U17 (N_17,In_158,In_128);
nand U18 (N_18,In_240,In_262);
nor U19 (N_19,In_380,In_197);
nor U20 (N_20,In_289,In_40);
or U21 (N_21,In_335,In_487);
or U22 (N_22,In_435,In_413);
and U23 (N_23,In_230,In_244);
nor U24 (N_24,In_364,In_454);
nand U25 (N_25,In_404,In_349);
or U26 (N_26,In_388,In_13);
and U27 (N_27,In_59,In_317);
nor U28 (N_28,In_301,In_92);
or U29 (N_29,In_470,In_365);
and U30 (N_30,In_278,In_210);
or U31 (N_31,In_493,In_137);
or U32 (N_32,In_490,In_94);
and U33 (N_33,In_187,In_494);
and U34 (N_34,In_442,In_163);
and U35 (N_35,In_372,In_408);
or U36 (N_36,In_218,In_273);
nand U37 (N_37,In_248,In_157);
nor U38 (N_38,In_498,In_377);
and U39 (N_39,In_264,In_2);
and U40 (N_40,In_135,In_62);
and U41 (N_41,In_4,In_192);
nand U42 (N_42,In_363,In_252);
nand U43 (N_43,In_444,In_106);
nor U44 (N_44,In_207,In_279);
or U45 (N_45,In_479,In_167);
or U46 (N_46,In_24,In_6);
nand U47 (N_47,In_366,In_72);
nor U48 (N_48,In_419,In_189);
or U49 (N_49,In_330,In_247);
or U50 (N_50,In_292,In_324);
nor U51 (N_51,In_477,In_299);
and U52 (N_52,In_184,In_125);
nand U53 (N_53,In_461,In_394);
and U54 (N_54,In_474,In_190);
nand U55 (N_55,In_65,In_473);
nor U56 (N_56,In_235,In_456);
nor U57 (N_57,In_297,In_356);
and U58 (N_58,In_234,In_307);
or U59 (N_59,In_104,In_126);
and U60 (N_60,In_432,In_123);
and U61 (N_61,In_220,In_97);
or U62 (N_62,In_114,In_336);
or U63 (N_63,In_261,In_180);
and U64 (N_64,In_39,In_451);
and U65 (N_65,In_194,In_395);
and U66 (N_66,In_338,In_358);
nand U67 (N_67,In_132,In_7);
nor U68 (N_68,In_124,In_211);
and U69 (N_69,In_93,In_156);
and U70 (N_70,In_303,In_386);
nand U71 (N_71,In_249,In_339);
nor U72 (N_72,In_313,In_269);
nand U73 (N_73,In_134,In_66);
nor U74 (N_74,In_96,In_239);
or U75 (N_75,In_312,In_164);
nor U76 (N_76,In_369,In_58);
or U77 (N_77,In_393,In_453);
nor U78 (N_78,In_30,In_411);
nor U79 (N_79,In_280,In_286);
nand U80 (N_80,In_226,In_77);
nor U81 (N_81,In_424,In_466);
and U82 (N_82,In_384,In_208);
nor U83 (N_83,In_452,In_397);
nand U84 (N_84,In_344,In_352);
nor U85 (N_85,In_205,In_115);
nor U86 (N_86,In_222,In_354);
nand U87 (N_87,In_326,In_469);
nand U88 (N_88,In_142,In_460);
nor U89 (N_89,In_54,In_351);
and U90 (N_90,In_52,In_50);
and U91 (N_91,In_232,In_271);
nor U92 (N_92,In_57,In_412);
or U93 (N_93,In_159,In_171);
and U94 (N_94,In_136,In_475);
nor U95 (N_95,In_119,In_434);
nor U96 (N_96,In_68,In_329);
and U97 (N_97,In_140,In_485);
and U98 (N_98,In_102,In_311);
nand U99 (N_99,In_256,In_200);
nor U100 (N_100,In_201,In_433);
or U101 (N_101,In_350,In_83);
xnor U102 (N_102,In_316,In_148);
nor U103 (N_103,In_304,In_308);
nand U104 (N_104,In_492,In_467);
nand U105 (N_105,In_224,In_154);
nand U106 (N_106,In_78,In_290);
nor U107 (N_107,In_277,In_254);
and U108 (N_108,In_282,In_80);
or U109 (N_109,In_348,In_87);
or U110 (N_110,In_376,In_191);
and U111 (N_111,In_251,In_99);
nand U112 (N_112,In_310,In_430);
nand U113 (N_113,In_320,In_332);
or U114 (N_114,In_331,In_175);
nand U115 (N_115,In_91,In_300);
or U116 (N_116,In_34,In_382);
nand U117 (N_117,In_143,In_450);
and U118 (N_118,In_245,In_169);
or U119 (N_119,In_8,In_464);
or U120 (N_120,In_69,In_64);
nor U121 (N_121,In_107,In_437);
nand U122 (N_122,In_496,In_19);
nand U123 (N_123,In_228,In_246);
or U124 (N_124,In_353,In_445);
and U125 (N_125,In_459,In_403);
nand U126 (N_126,In_294,In_36);
or U127 (N_127,In_274,In_103);
nand U128 (N_128,In_33,In_321);
nor U129 (N_129,In_355,In_448);
nand U130 (N_130,In_116,In_370);
or U131 (N_131,In_231,In_32);
nor U132 (N_132,In_468,In_275);
nor U133 (N_133,In_499,In_139);
and U134 (N_134,In_37,In_392);
or U135 (N_135,In_298,In_407);
nor U136 (N_136,In_15,In_266);
nor U137 (N_137,In_117,In_56);
or U138 (N_138,In_165,In_43);
or U139 (N_139,In_71,In_458);
nand U140 (N_140,In_122,In_166);
or U141 (N_141,In_414,In_283);
nand U142 (N_142,In_95,In_27);
or U143 (N_143,In_219,In_111);
nand U144 (N_144,In_155,In_90);
and U145 (N_145,In_53,In_127);
nand U146 (N_146,In_185,In_179);
nor U147 (N_147,In_28,In_45);
nor U148 (N_148,In_25,In_447);
nor U149 (N_149,In_21,In_405);
xnor U150 (N_150,In_284,In_409);
and U151 (N_151,In_85,In_225);
nor U152 (N_152,In_476,In_441);
or U153 (N_153,In_378,In_196);
and U154 (N_154,In_359,In_415);
or U155 (N_155,In_150,In_401);
nor U156 (N_156,In_305,In_35);
and U157 (N_157,In_74,In_152);
or U158 (N_158,In_141,In_422);
and U159 (N_159,In_73,In_26);
nand U160 (N_160,In_203,In_209);
nor U161 (N_161,In_12,In_60);
or U162 (N_162,In_181,In_229);
or U163 (N_163,In_257,In_265);
nor U164 (N_164,In_287,In_288);
and U165 (N_165,In_398,In_406);
nand U166 (N_166,In_291,In_215);
and U167 (N_167,In_118,In_236);
and U168 (N_168,In_174,In_144);
nand U169 (N_169,In_391,In_98);
or U170 (N_170,In_112,In_295);
nand U171 (N_171,In_55,In_421);
nand U172 (N_172,In_16,In_10);
nor U173 (N_173,In_51,In_488);
or U174 (N_174,In_345,In_368);
nor U175 (N_175,In_67,In_70);
and U176 (N_176,In_177,In_38);
or U177 (N_177,In_462,In_285);
nand U178 (N_178,In_237,In_253);
and U179 (N_179,In_63,In_100);
and U180 (N_180,In_325,In_121);
or U181 (N_181,In_342,In_199);
nor U182 (N_182,In_88,In_480);
xor U183 (N_183,In_193,In_387);
or U184 (N_184,In_455,In_110);
nand U185 (N_185,In_258,In_11);
nor U186 (N_186,In_385,In_416);
nor U187 (N_187,In_202,In_337);
nand U188 (N_188,In_497,In_431);
or U189 (N_189,In_46,In_161);
and U190 (N_190,In_357,In_268);
or U191 (N_191,In_82,In_449);
nor U192 (N_192,In_176,In_495);
nor U193 (N_193,In_425,In_327);
or U194 (N_194,In_396,In_478);
and U195 (N_195,In_259,In_423);
nand U196 (N_196,In_272,In_212);
and U197 (N_197,In_373,In_206);
and U198 (N_198,In_1,In_347);
nand U199 (N_199,In_44,In_173);
nand U200 (N_200,In_318,In_426);
nor U201 (N_201,In_362,In_436);
nor U202 (N_202,In_195,In_145);
nor U203 (N_203,In_333,In_213);
or U204 (N_204,In_319,In_481);
nor U205 (N_205,In_22,In_260);
nor U206 (N_206,In_483,In_379);
nand U207 (N_207,In_214,In_242);
nor U208 (N_208,In_29,In_361);
nand U209 (N_209,In_418,In_217);
nor U210 (N_210,In_31,In_323);
nand U211 (N_211,In_446,In_328);
nand U212 (N_212,In_491,In_233);
or U213 (N_213,In_216,In_399);
nor U214 (N_214,In_138,In_389);
nor U215 (N_215,In_375,In_186);
nor U216 (N_216,In_120,In_48);
nand U217 (N_217,In_113,In_371);
nand U218 (N_218,In_417,In_41);
or U219 (N_219,In_341,In_81);
nor U220 (N_220,In_343,In_465);
nor U221 (N_221,In_315,In_149);
or U222 (N_222,In_20,In_482);
or U223 (N_223,In_346,In_5);
nand U224 (N_224,In_170,In_101);
nand U225 (N_225,In_3,In_130);
or U226 (N_226,In_129,In_105);
or U227 (N_227,In_428,In_47);
nand U228 (N_228,In_221,In_84);
nor U229 (N_229,In_61,In_188);
and U230 (N_230,In_276,In_79);
nor U231 (N_231,In_367,In_381);
nor U232 (N_232,In_23,In_302);
or U233 (N_233,In_223,In_484);
or U234 (N_234,In_198,In_178);
and U235 (N_235,In_440,In_270);
and U236 (N_236,In_238,In_76);
nand U237 (N_237,In_439,In_0);
nor U238 (N_238,In_151,In_486);
or U239 (N_239,In_296,In_322);
nand U240 (N_240,In_400,In_314);
nand U241 (N_241,In_14,In_153);
and U242 (N_242,In_263,In_463);
or U243 (N_243,In_227,In_420);
and U244 (N_244,In_472,In_309);
or U245 (N_245,In_146,In_18);
nand U246 (N_246,In_250,In_306);
or U247 (N_247,In_89,In_427);
and U248 (N_248,In_255,In_410);
and U249 (N_249,In_457,In_17);
nor U250 (N_250,In_405,In_458);
nand U251 (N_251,In_313,In_355);
and U252 (N_252,In_46,In_39);
nor U253 (N_253,In_199,In_58);
nand U254 (N_254,In_437,In_484);
and U255 (N_255,In_95,In_8);
nor U256 (N_256,In_280,In_208);
and U257 (N_257,In_369,In_153);
and U258 (N_258,In_405,In_1);
and U259 (N_259,In_22,In_131);
nor U260 (N_260,In_494,In_14);
or U261 (N_261,In_464,In_263);
nor U262 (N_262,In_396,In_90);
and U263 (N_263,In_272,In_452);
and U264 (N_264,In_138,In_66);
nand U265 (N_265,In_227,In_129);
xnor U266 (N_266,In_64,In_396);
nand U267 (N_267,In_381,In_15);
nand U268 (N_268,In_249,In_172);
nor U269 (N_269,In_68,In_24);
nor U270 (N_270,In_87,In_59);
nand U271 (N_271,In_470,In_271);
or U272 (N_272,In_17,In_88);
nor U273 (N_273,In_366,In_36);
nand U274 (N_274,In_359,In_113);
nand U275 (N_275,In_281,In_496);
nor U276 (N_276,In_81,In_171);
and U277 (N_277,In_391,In_278);
and U278 (N_278,In_480,In_261);
and U279 (N_279,In_210,In_158);
nor U280 (N_280,In_159,In_471);
nor U281 (N_281,In_39,In_336);
nand U282 (N_282,In_122,In_482);
nand U283 (N_283,In_350,In_23);
and U284 (N_284,In_248,In_50);
and U285 (N_285,In_192,In_363);
and U286 (N_286,In_354,In_342);
nand U287 (N_287,In_424,In_103);
nor U288 (N_288,In_465,In_150);
and U289 (N_289,In_14,In_86);
or U290 (N_290,In_234,In_478);
nor U291 (N_291,In_129,In_215);
and U292 (N_292,In_177,In_65);
nand U293 (N_293,In_296,In_312);
nor U294 (N_294,In_137,In_183);
and U295 (N_295,In_491,In_328);
or U296 (N_296,In_454,In_87);
or U297 (N_297,In_123,In_174);
or U298 (N_298,In_52,In_368);
or U299 (N_299,In_298,In_442);
nor U300 (N_300,In_371,In_274);
nor U301 (N_301,In_174,In_86);
or U302 (N_302,In_135,In_295);
nand U303 (N_303,In_44,In_203);
and U304 (N_304,In_1,In_456);
nand U305 (N_305,In_441,In_337);
or U306 (N_306,In_119,In_399);
nand U307 (N_307,In_261,In_123);
nand U308 (N_308,In_225,In_170);
nand U309 (N_309,In_223,In_205);
nand U310 (N_310,In_56,In_25);
nand U311 (N_311,In_240,In_195);
nor U312 (N_312,In_342,In_267);
nor U313 (N_313,In_113,In_365);
and U314 (N_314,In_361,In_81);
nor U315 (N_315,In_60,In_401);
nand U316 (N_316,In_235,In_452);
and U317 (N_317,In_139,In_424);
and U318 (N_318,In_459,In_4);
or U319 (N_319,In_27,In_320);
nand U320 (N_320,In_400,In_187);
nand U321 (N_321,In_99,In_74);
and U322 (N_322,In_301,In_453);
or U323 (N_323,In_46,In_391);
nor U324 (N_324,In_400,In_336);
or U325 (N_325,In_278,In_84);
nand U326 (N_326,In_365,In_2);
or U327 (N_327,In_352,In_484);
and U328 (N_328,In_314,In_32);
nand U329 (N_329,In_37,In_22);
nand U330 (N_330,In_499,In_328);
nand U331 (N_331,In_43,In_246);
or U332 (N_332,In_182,In_159);
nor U333 (N_333,In_387,In_191);
or U334 (N_334,In_386,In_265);
nor U335 (N_335,In_199,In_497);
nand U336 (N_336,In_96,In_123);
or U337 (N_337,In_82,In_24);
nand U338 (N_338,In_131,In_212);
nand U339 (N_339,In_161,In_286);
and U340 (N_340,In_189,In_208);
nor U341 (N_341,In_280,In_310);
or U342 (N_342,In_212,In_207);
and U343 (N_343,In_257,In_28);
nand U344 (N_344,In_387,In_208);
nand U345 (N_345,In_117,In_333);
and U346 (N_346,In_74,In_389);
nand U347 (N_347,In_312,In_479);
or U348 (N_348,In_351,In_202);
nand U349 (N_349,In_416,In_351);
nor U350 (N_350,In_261,In_140);
nand U351 (N_351,In_346,In_333);
nand U352 (N_352,In_274,In_80);
and U353 (N_353,In_292,In_284);
nor U354 (N_354,In_413,In_91);
and U355 (N_355,In_113,In_132);
and U356 (N_356,In_462,In_293);
nor U357 (N_357,In_155,In_266);
nand U358 (N_358,In_271,In_225);
nor U359 (N_359,In_122,In_356);
or U360 (N_360,In_295,In_493);
and U361 (N_361,In_480,In_356);
nor U362 (N_362,In_217,In_261);
and U363 (N_363,In_220,In_181);
nor U364 (N_364,In_229,In_318);
or U365 (N_365,In_109,In_313);
or U366 (N_366,In_337,In_296);
nand U367 (N_367,In_89,In_489);
and U368 (N_368,In_156,In_29);
and U369 (N_369,In_180,In_416);
nor U370 (N_370,In_308,In_158);
and U371 (N_371,In_73,In_143);
nand U372 (N_372,In_491,In_109);
nor U373 (N_373,In_371,In_446);
nand U374 (N_374,In_79,In_284);
and U375 (N_375,In_182,In_37);
or U376 (N_376,In_97,In_461);
nand U377 (N_377,In_421,In_335);
and U378 (N_378,In_68,In_456);
nor U379 (N_379,In_15,In_342);
and U380 (N_380,In_147,In_246);
or U381 (N_381,In_481,In_86);
and U382 (N_382,In_176,In_276);
nand U383 (N_383,In_337,In_249);
nand U384 (N_384,In_476,In_495);
and U385 (N_385,In_159,In_105);
and U386 (N_386,In_278,In_61);
xnor U387 (N_387,In_377,In_265);
nand U388 (N_388,In_494,In_421);
and U389 (N_389,In_233,In_476);
or U390 (N_390,In_244,In_330);
nand U391 (N_391,In_56,In_153);
nand U392 (N_392,In_168,In_136);
or U393 (N_393,In_174,In_176);
or U394 (N_394,In_466,In_235);
and U395 (N_395,In_245,In_426);
or U396 (N_396,In_266,In_209);
nor U397 (N_397,In_57,In_434);
or U398 (N_398,In_95,In_162);
and U399 (N_399,In_307,In_401);
and U400 (N_400,In_478,In_95);
nand U401 (N_401,In_77,In_463);
or U402 (N_402,In_317,In_328);
and U403 (N_403,In_217,In_123);
nand U404 (N_404,In_487,In_449);
nor U405 (N_405,In_409,In_322);
nand U406 (N_406,In_18,In_329);
or U407 (N_407,In_413,In_150);
or U408 (N_408,In_135,In_331);
or U409 (N_409,In_206,In_372);
and U410 (N_410,In_32,In_18);
nand U411 (N_411,In_49,In_441);
nor U412 (N_412,In_273,In_174);
or U413 (N_413,In_119,In_171);
nand U414 (N_414,In_89,In_368);
and U415 (N_415,In_314,In_315);
nor U416 (N_416,In_452,In_224);
nor U417 (N_417,In_454,In_159);
or U418 (N_418,In_80,In_158);
or U419 (N_419,In_78,In_141);
nor U420 (N_420,In_43,In_492);
or U421 (N_421,In_189,In_118);
nand U422 (N_422,In_303,In_403);
nand U423 (N_423,In_103,In_290);
or U424 (N_424,In_13,In_46);
nand U425 (N_425,In_289,In_318);
or U426 (N_426,In_168,In_214);
and U427 (N_427,In_222,In_281);
nand U428 (N_428,In_153,In_66);
or U429 (N_429,In_172,In_434);
nor U430 (N_430,In_310,In_339);
or U431 (N_431,In_145,In_323);
or U432 (N_432,In_495,In_305);
and U433 (N_433,In_478,In_62);
and U434 (N_434,In_168,In_437);
nand U435 (N_435,In_93,In_343);
and U436 (N_436,In_400,In_467);
nand U437 (N_437,In_71,In_258);
or U438 (N_438,In_191,In_40);
nand U439 (N_439,In_461,In_303);
and U440 (N_440,In_136,In_19);
or U441 (N_441,In_320,In_415);
nor U442 (N_442,In_21,In_303);
nand U443 (N_443,In_359,In_217);
and U444 (N_444,In_248,In_65);
nand U445 (N_445,In_74,In_425);
nand U446 (N_446,In_120,In_268);
and U447 (N_447,In_335,In_367);
nand U448 (N_448,In_369,In_390);
nor U449 (N_449,In_78,In_334);
nor U450 (N_450,In_357,In_258);
or U451 (N_451,In_249,In_170);
or U452 (N_452,In_237,In_140);
nor U453 (N_453,In_220,In_422);
or U454 (N_454,In_460,In_126);
nand U455 (N_455,In_204,In_351);
nor U456 (N_456,In_268,In_420);
nor U457 (N_457,In_465,In_27);
xor U458 (N_458,In_99,In_445);
nor U459 (N_459,In_117,In_441);
and U460 (N_460,In_80,In_447);
or U461 (N_461,In_4,In_294);
and U462 (N_462,In_473,In_23);
nor U463 (N_463,In_215,In_88);
nor U464 (N_464,In_24,In_80);
or U465 (N_465,In_2,In_486);
and U466 (N_466,In_168,In_461);
and U467 (N_467,In_335,In_429);
nand U468 (N_468,In_436,In_118);
or U469 (N_469,In_221,In_467);
nand U470 (N_470,In_429,In_87);
or U471 (N_471,In_170,In_82);
or U472 (N_472,In_213,In_310);
nor U473 (N_473,In_175,In_299);
nor U474 (N_474,In_362,In_409);
nor U475 (N_475,In_99,In_451);
nand U476 (N_476,In_413,In_56);
nand U477 (N_477,In_361,In_384);
nand U478 (N_478,In_17,In_233);
nor U479 (N_479,In_9,In_18);
or U480 (N_480,In_424,In_234);
nor U481 (N_481,In_226,In_467);
nand U482 (N_482,In_6,In_314);
nor U483 (N_483,In_422,In_447);
nor U484 (N_484,In_324,In_187);
or U485 (N_485,In_3,In_267);
and U486 (N_486,In_375,In_241);
nor U487 (N_487,In_460,In_404);
nand U488 (N_488,In_127,In_57);
nand U489 (N_489,In_74,In_66);
nor U490 (N_490,In_480,In_425);
or U491 (N_491,In_125,In_499);
nor U492 (N_492,In_74,In_457);
nor U493 (N_493,In_355,In_15);
or U494 (N_494,In_189,In_344);
or U495 (N_495,In_44,In_370);
nor U496 (N_496,In_41,In_335);
nor U497 (N_497,In_357,In_256);
or U498 (N_498,In_394,In_236);
nand U499 (N_499,In_360,In_31);
nand U500 (N_500,In_365,In_398);
and U501 (N_501,In_384,In_6);
nor U502 (N_502,In_372,In_162);
nand U503 (N_503,In_79,In_101);
nand U504 (N_504,In_92,In_11);
or U505 (N_505,In_280,In_233);
and U506 (N_506,In_237,In_257);
nor U507 (N_507,In_133,In_372);
and U508 (N_508,In_458,In_480);
nand U509 (N_509,In_130,In_348);
and U510 (N_510,In_171,In_499);
nand U511 (N_511,In_296,In_119);
and U512 (N_512,In_38,In_4);
and U513 (N_513,In_108,In_54);
nor U514 (N_514,In_173,In_154);
nor U515 (N_515,In_56,In_132);
nor U516 (N_516,In_255,In_4);
or U517 (N_517,In_28,In_488);
and U518 (N_518,In_192,In_205);
and U519 (N_519,In_360,In_128);
nand U520 (N_520,In_180,In_465);
and U521 (N_521,In_206,In_323);
or U522 (N_522,In_347,In_87);
and U523 (N_523,In_109,In_197);
nor U524 (N_524,In_122,In_340);
nand U525 (N_525,In_427,In_4);
or U526 (N_526,In_164,In_491);
nand U527 (N_527,In_399,In_489);
nor U528 (N_528,In_445,In_211);
and U529 (N_529,In_334,In_288);
nor U530 (N_530,In_254,In_477);
and U531 (N_531,In_317,In_405);
nand U532 (N_532,In_211,In_404);
nand U533 (N_533,In_347,In_204);
or U534 (N_534,In_430,In_396);
and U535 (N_535,In_52,In_374);
and U536 (N_536,In_260,In_395);
nand U537 (N_537,In_455,In_411);
nor U538 (N_538,In_365,In_461);
or U539 (N_539,In_32,In_420);
nand U540 (N_540,In_355,In_426);
or U541 (N_541,In_301,In_209);
and U542 (N_542,In_432,In_150);
or U543 (N_543,In_45,In_433);
nor U544 (N_544,In_25,In_109);
or U545 (N_545,In_416,In_461);
nand U546 (N_546,In_381,In_347);
and U547 (N_547,In_196,In_445);
and U548 (N_548,In_356,In_148);
nand U549 (N_549,In_182,In_244);
nand U550 (N_550,In_159,In_42);
nand U551 (N_551,In_204,In_231);
and U552 (N_552,In_33,In_188);
nand U553 (N_553,In_145,In_377);
nand U554 (N_554,In_162,In_414);
nor U555 (N_555,In_72,In_59);
nand U556 (N_556,In_208,In_33);
nand U557 (N_557,In_107,In_101);
or U558 (N_558,In_431,In_304);
nand U559 (N_559,In_174,In_456);
and U560 (N_560,In_0,In_206);
nor U561 (N_561,In_404,In_327);
and U562 (N_562,In_437,In_93);
nand U563 (N_563,In_448,In_94);
xnor U564 (N_564,In_5,In_320);
nand U565 (N_565,In_103,In_401);
nor U566 (N_566,In_55,In_226);
and U567 (N_567,In_182,In_429);
nand U568 (N_568,In_445,In_175);
or U569 (N_569,In_164,In_420);
or U570 (N_570,In_152,In_305);
or U571 (N_571,In_401,In_373);
xor U572 (N_572,In_187,In_488);
or U573 (N_573,In_402,In_329);
or U574 (N_574,In_465,In_291);
nor U575 (N_575,In_401,In_448);
nand U576 (N_576,In_130,In_265);
nand U577 (N_577,In_453,In_464);
nor U578 (N_578,In_326,In_70);
or U579 (N_579,In_335,In_208);
and U580 (N_580,In_461,In_267);
nand U581 (N_581,In_365,In_299);
and U582 (N_582,In_310,In_259);
or U583 (N_583,In_171,In_370);
and U584 (N_584,In_167,In_405);
and U585 (N_585,In_69,In_144);
or U586 (N_586,In_224,In_447);
nor U587 (N_587,In_241,In_450);
or U588 (N_588,In_256,In_435);
nor U589 (N_589,In_165,In_135);
nor U590 (N_590,In_87,In_372);
nand U591 (N_591,In_115,In_109);
nand U592 (N_592,In_65,In_34);
or U593 (N_593,In_326,In_325);
or U594 (N_594,In_156,In_278);
and U595 (N_595,In_324,In_69);
and U596 (N_596,In_187,In_228);
and U597 (N_597,In_410,In_368);
nand U598 (N_598,In_25,In_170);
nor U599 (N_599,In_172,In_83);
nand U600 (N_600,In_273,In_157);
xor U601 (N_601,In_245,In_237);
or U602 (N_602,In_48,In_449);
nor U603 (N_603,In_453,In_493);
nand U604 (N_604,In_71,In_104);
nor U605 (N_605,In_135,In_179);
or U606 (N_606,In_416,In_380);
nor U607 (N_607,In_218,In_429);
nor U608 (N_608,In_463,In_182);
nor U609 (N_609,In_198,In_237);
and U610 (N_610,In_229,In_430);
or U611 (N_611,In_476,In_39);
and U612 (N_612,In_433,In_353);
nand U613 (N_613,In_62,In_21);
or U614 (N_614,In_194,In_169);
and U615 (N_615,In_146,In_92);
or U616 (N_616,In_337,In_483);
nor U617 (N_617,In_340,In_159);
and U618 (N_618,In_35,In_128);
or U619 (N_619,In_487,In_416);
nor U620 (N_620,In_383,In_367);
or U621 (N_621,In_190,In_360);
or U622 (N_622,In_374,In_125);
nand U623 (N_623,In_245,In_487);
or U624 (N_624,In_130,In_450);
nor U625 (N_625,In_490,In_434);
nand U626 (N_626,In_275,In_466);
or U627 (N_627,In_64,In_90);
nor U628 (N_628,In_72,In_257);
nand U629 (N_629,In_496,In_430);
or U630 (N_630,In_328,In_54);
and U631 (N_631,In_196,In_168);
nand U632 (N_632,In_422,In_197);
and U633 (N_633,In_29,In_281);
and U634 (N_634,In_495,In_301);
or U635 (N_635,In_346,In_36);
and U636 (N_636,In_244,In_319);
or U637 (N_637,In_261,In_418);
or U638 (N_638,In_413,In_307);
nand U639 (N_639,In_176,In_437);
and U640 (N_640,In_13,In_153);
nor U641 (N_641,In_399,In_96);
and U642 (N_642,In_256,In_368);
or U643 (N_643,In_386,In_400);
or U644 (N_644,In_203,In_83);
nor U645 (N_645,In_416,In_285);
and U646 (N_646,In_41,In_163);
or U647 (N_647,In_102,In_476);
or U648 (N_648,In_86,In_60);
or U649 (N_649,In_492,In_33);
and U650 (N_650,In_222,In_282);
and U651 (N_651,In_364,In_300);
and U652 (N_652,In_318,In_411);
or U653 (N_653,In_473,In_248);
or U654 (N_654,In_151,In_472);
nand U655 (N_655,In_267,In_193);
nand U656 (N_656,In_97,In_183);
nand U657 (N_657,In_319,In_448);
nand U658 (N_658,In_67,In_251);
or U659 (N_659,In_436,In_99);
and U660 (N_660,In_7,In_122);
nand U661 (N_661,In_278,In_91);
nor U662 (N_662,In_425,In_51);
nand U663 (N_663,In_427,In_179);
and U664 (N_664,In_379,In_348);
nor U665 (N_665,In_286,In_189);
and U666 (N_666,In_262,In_210);
and U667 (N_667,In_369,In_416);
nand U668 (N_668,In_363,In_247);
nor U669 (N_669,In_197,In_271);
nand U670 (N_670,In_109,In_289);
nor U671 (N_671,In_131,In_194);
and U672 (N_672,In_392,In_388);
or U673 (N_673,In_372,In_98);
or U674 (N_674,In_283,In_217);
nor U675 (N_675,In_400,In_342);
and U676 (N_676,In_393,In_432);
xor U677 (N_677,In_148,In_64);
or U678 (N_678,In_94,In_422);
nor U679 (N_679,In_183,In_151);
nor U680 (N_680,In_239,In_407);
nand U681 (N_681,In_47,In_290);
or U682 (N_682,In_414,In_8);
and U683 (N_683,In_184,In_322);
nor U684 (N_684,In_110,In_429);
or U685 (N_685,In_387,In_268);
nor U686 (N_686,In_306,In_351);
nand U687 (N_687,In_234,In_468);
or U688 (N_688,In_203,In_491);
and U689 (N_689,In_42,In_361);
and U690 (N_690,In_289,In_18);
or U691 (N_691,In_174,In_64);
or U692 (N_692,In_446,In_306);
nand U693 (N_693,In_340,In_394);
or U694 (N_694,In_81,In_47);
and U695 (N_695,In_134,In_30);
or U696 (N_696,In_488,In_324);
and U697 (N_697,In_453,In_127);
nor U698 (N_698,In_367,In_352);
nand U699 (N_699,In_279,In_71);
nor U700 (N_700,In_188,In_172);
nand U701 (N_701,In_74,In_143);
and U702 (N_702,In_264,In_440);
nand U703 (N_703,In_259,In_457);
nor U704 (N_704,In_326,In_161);
and U705 (N_705,In_78,In_153);
nand U706 (N_706,In_98,In_195);
nor U707 (N_707,In_109,In_406);
or U708 (N_708,In_88,In_464);
and U709 (N_709,In_204,In_289);
or U710 (N_710,In_421,In_285);
nand U711 (N_711,In_220,In_58);
or U712 (N_712,In_79,In_378);
nand U713 (N_713,In_262,In_146);
or U714 (N_714,In_278,In_386);
nand U715 (N_715,In_60,In_460);
nand U716 (N_716,In_217,In_78);
nand U717 (N_717,In_352,In_74);
or U718 (N_718,In_258,In_398);
and U719 (N_719,In_247,In_162);
or U720 (N_720,In_307,In_4);
nor U721 (N_721,In_498,In_437);
or U722 (N_722,In_36,In_251);
and U723 (N_723,In_423,In_368);
or U724 (N_724,In_87,In_172);
nand U725 (N_725,In_378,In_199);
and U726 (N_726,In_44,In_402);
or U727 (N_727,In_428,In_465);
and U728 (N_728,In_70,In_250);
nor U729 (N_729,In_9,In_108);
nor U730 (N_730,In_316,In_385);
and U731 (N_731,In_70,In_426);
and U732 (N_732,In_154,In_480);
nor U733 (N_733,In_84,In_489);
nand U734 (N_734,In_186,In_184);
and U735 (N_735,In_98,In_408);
nand U736 (N_736,In_47,In_261);
nor U737 (N_737,In_189,In_16);
and U738 (N_738,In_179,In_279);
nor U739 (N_739,In_490,In_147);
or U740 (N_740,In_261,In_55);
nor U741 (N_741,In_403,In_181);
or U742 (N_742,In_489,In_428);
nor U743 (N_743,In_326,In_385);
nand U744 (N_744,In_350,In_412);
nor U745 (N_745,In_318,In_378);
and U746 (N_746,In_179,In_66);
nor U747 (N_747,In_300,In_278);
or U748 (N_748,In_489,In_326);
or U749 (N_749,In_318,In_28);
or U750 (N_750,In_18,In_163);
nor U751 (N_751,In_283,In_243);
or U752 (N_752,In_128,In_463);
nand U753 (N_753,In_106,In_207);
and U754 (N_754,In_64,In_155);
nand U755 (N_755,In_229,In_163);
nor U756 (N_756,In_345,In_498);
or U757 (N_757,In_359,In_79);
and U758 (N_758,In_33,In_323);
or U759 (N_759,In_156,In_37);
nand U760 (N_760,In_103,In_161);
nor U761 (N_761,In_431,In_439);
xnor U762 (N_762,In_162,In_14);
nand U763 (N_763,In_47,In_145);
nor U764 (N_764,In_228,In_488);
nor U765 (N_765,In_96,In_273);
or U766 (N_766,In_141,In_114);
nor U767 (N_767,In_14,In_320);
and U768 (N_768,In_240,In_323);
nor U769 (N_769,In_72,In_138);
or U770 (N_770,In_319,In_142);
or U771 (N_771,In_87,In_300);
nand U772 (N_772,In_413,In_112);
or U773 (N_773,In_95,In_425);
and U774 (N_774,In_18,In_348);
nand U775 (N_775,In_33,In_497);
or U776 (N_776,In_16,In_333);
and U777 (N_777,In_27,In_311);
and U778 (N_778,In_149,In_386);
nor U779 (N_779,In_478,In_59);
nand U780 (N_780,In_241,In_304);
and U781 (N_781,In_499,In_400);
or U782 (N_782,In_187,In_322);
nand U783 (N_783,In_236,In_416);
or U784 (N_784,In_404,In_59);
or U785 (N_785,In_494,In_402);
nand U786 (N_786,In_336,In_209);
or U787 (N_787,In_361,In_277);
and U788 (N_788,In_50,In_154);
or U789 (N_789,In_227,In_434);
nand U790 (N_790,In_170,In_158);
and U791 (N_791,In_305,In_20);
nor U792 (N_792,In_288,In_14);
nor U793 (N_793,In_52,In_158);
nor U794 (N_794,In_477,In_3);
nand U795 (N_795,In_440,In_346);
and U796 (N_796,In_23,In_58);
nand U797 (N_797,In_183,In_40);
or U798 (N_798,In_321,In_298);
nand U799 (N_799,In_386,In_325);
nor U800 (N_800,In_323,In_128);
nand U801 (N_801,In_303,In_183);
nor U802 (N_802,In_405,In_56);
and U803 (N_803,In_234,In_224);
or U804 (N_804,In_118,In_326);
and U805 (N_805,In_197,In_170);
or U806 (N_806,In_339,In_2);
or U807 (N_807,In_49,In_426);
nor U808 (N_808,In_206,In_24);
nor U809 (N_809,In_128,In_144);
and U810 (N_810,In_70,In_73);
or U811 (N_811,In_57,In_133);
or U812 (N_812,In_83,In_319);
nand U813 (N_813,In_125,In_148);
nor U814 (N_814,In_296,In_272);
nand U815 (N_815,In_151,In_399);
nand U816 (N_816,In_68,In_297);
and U817 (N_817,In_366,In_361);
nand U818 (N_818,In_328,In_309);
nand U819 (N_819,In_454,In_378);
nor U820 (N_820,In_485,In_77);
or U821 (N_821,In_490,In_368);
or U822 (N_822,In_252,In_321);
or U823 (N_823,In_309,In_200);
nor U824 (N_824,In_423,In_311);
or U825 (N_825,In_7,In_461);
nand U826 (N_826,In_378,In_419);
nand U827 (N_827,In_283,In_441);
and U828 (N_828,In_413,In_423);
nor U829 (N_829,In_41,In_402);
and U830 (N_830,In_468,In_439);
or U831 (N_831,In_151,In_268);
nor U832 (N_832,In_203,In_144);
or U833 (N_833,In_279,In_430);
and U834 (N_834,In_209,In_93);
or U835 (N_835,In_37,In_9);
or U836 (N_836,In_109,In_233);
or U837 (N_837,In_217,In_300);
nand U838 (N_838,In_8,In_47);
nor U839 (N_839,In_83,In_35);
and U840 (N_840,In_203,In_283);
or U841 (N_841,In_180,In_330);
and U842 (N_842,In_451,In_389);
nand U843 (N_843,In_349,In_55);
or U844 (N_844,In_79,In_348);
and U845 (N_845,In_480,In_190);
nor U846 (N_846,In_327,In_303);
nor U847 (N_847,In_441,In_93);
nor U848 (N_848,In_395,In_284);
nand U849 (N_849,In_467,In_122);
and U850 (N_850,In_408,In_415);
nand U851 (N_851,In_379,In_9);
nand U852 (N_852,In_133,In_58);
and U853 (N_853,In_462,In_170);
or U854 (N_854,In_268,In_423);
xor U855 (N_855,In_339,In_257);
and U856 (N_856,In_129,In_314);
or U857 (N_857,In_467,In_198);
and U858 (N_858,In_227,In_214);
nand U859 (N_859,In_409,In_264);
and U860 (N_860,In_34,In_182);
and U861 (N_861,In_33,In_177);
or U862 (N_862,In_237,In_415);
and U863 (N_863,In_8,In_401);
and U864 (N_864,In_96,In_80);
nor U865 (N_865,In_368,In_315);
and U866 (N_866,In_158,In_153);
xor U867 (N_867,In_233,In_388);
nor U868 (N_868,In_151,In_105);
nor U869 (N_869,In_79,In_274);
nand U870 (N_870,In_290,In_374);
and U871 (N_871,In_358,In_395);
nand U872 (N_872,In_261,In_442);
or U873 (N_873,In_159,In_461);
and U874 (N_874,In_119,In_484);
nand U875 (N_875,In_346,In_155);
nor U876 (N_876,In_138,In_98);
nor U877 (N_877,In_494,In_310);
or U878 (N_878,In_284,In_381);
and U879 (N_879,In_221,In_41);
nand U880 (N_880,In_434,In_156);
nand U881 (N_881,In_288,In_497);
nand U882 (N_882,In_27,In_272);
nor U883 (N_883,In_317,In_394);
nor U884 (N_884,In_315,In_175);
or U885 (N_885,In_477,In_495);
and U886 (N_886,In_213,In_181);
nand U887 (N_887,In_228,In_99);
nand U888 (N_888,In_274,In_420);
or U889 (N_889,In_337,In_306);
or U890 (N_890,In_41,In_357);
or U891 (N_891,In_279,In_322);
or U892 (N_892,In_355,In_85);
nand U893 (N_893,In_366,In_59);
nor U894 (N_894,In_427,In_90);
or U895 (N_895,In_377,In_384);
nor U896 (N_896,In_441,In_228);
and U897 (N_897,In_53,In_183);
nor U898 (N_898,In_244,In_187);
and U899 (N_899,In_324,In_455);
nor U900 (N_900,In_1,In_262);
xnor U901 (N_901,In_50,In_390);
and U902 (N_902,In_92,In_436);
nor U903 (N_903,In_318,In_321);
nand U904 (N_904,In_378,In_55);
nor U905 (N_905,In_347,In_39);
or U906 (N_906,In_40,In_101);
and U907 (N_907,In_184,In_143);
and U908 (N_908,In_252,In_449);
nand U909 (N_909,In_246,In_210);
nor U910 (N_910,In_194,In_101);
nor U911 (N_911,In_258,In_99);
and U912 (N_912,In_205,In_134);
nor U913 (N_913,In_84,In_330);
nor U914 (N_914,In_8,In_2);
and U915 (N_915,In_229,In_340);
nor U916 (N_916,In_447,In_249);
nor U917 (N_917,In_488,In_56);
or U918 (N_918,In_333,In_250);
nand U919 (N_919,In_13,In_330);
nand U920 (N_920,In_147,In_139);
and U921 (N_921,In_50,In_33);
nor U922 (N_922,In_363,In_386);
nor U923 (N_923,In_390,In_231);
nand U924 (N_924,In_217,In_491);
nand U925 (N_925,In_356,In_473);
nand U926 (N_926,In_120,In_83);
or U927 (N_927,In_446,In_480);
nor U928 (N_928,In_491,In_236);
and U929 (N_929,In_107,In_246);
and U930 (N_930,In_87,In_435);
nor U931 (N_931,In_193,In_316);
nor U932 (N_932,In_448,In_477);
and U933 (N_933,In_442,In_453);
nand U934 (N_934,In_239,In_403);
or U935 (N_935,In_378,In_34);
and U936 (N_936,In_234,In_342);
nor U937 (N_937,In_408,In_119);
nand U938 (N_938,In_462,In_225);
and U939 (N_939,In_458,In_77);
or U940 (N_940,In_71,In_498);
and U941 (N_941,In_223,In_447);
nor U942 (N_942,In_378,In_471);
nor U943 (N_943,In_481,In_427);
nor U944 (N_944,In_448,In_193);
and U945 (N_945,In_55,In_438);
nand U946 (N_946,In_144,In_484);
or U947 (N_947,In_286,In_27);
and U948 (N_948,In_112,In_70);
nor U949 (N_949,In_220,In_59);
and U950 (N_950,In_99,In_418);
or U951 (N_951,In_291,In_403);
or U952 (N_952,In_104,In_481);
nand U953 (N_953,In_282,In_337);
and U954 (N_954,In_46,In_371);
or U955 (N_955,In_190,In_49);
or U956 (N_956,In_65,In_299);
and U957 (N_957,In_200,In_115);
and U958 (N_958,In_217,In_424);
or U959 (N_959,In_433,In_232);
nor U960 (N_960,In_361,In_7);
and U961 (N_961,In_297,In_29);
and U962 (N_962,In_232,In_80);
nand U963 (N_963,In_472,In_170);
and U964 (N_964,In_410,In_101);
nor U965 (N_965,In_171,In_133);
nand U966 (N_966,In_144,In_196);
or U967 (N_967,In_53,In_237);
nand U968 (N_968,In_339,In_100);
nor U969 (N_969,In_137,In_358);
and U970 (N_970,In_124,In_6);
and U971 (N_971,In_263,In_460);
or U972 (N_972,In_85,In_489);
nand U973 (N_973,In_195,In_32);
nand U974 (N_974,In_451,In_292);
nor U975 (N_975,In_351,In_94);
nor U976 (N_976,In_139,In_162);
nor U977 (N_977,In_83,In_215);
nand U978 (N_978,In_90,In_168);
and U979 (N_979,In_34,In_25);
or U980 (N_980,In_76,In_143);
and U981 (N_981,In_115,In_126);
or U982 (N_982,In_338,In_282);
nor U983 (N_983,In_246,In_254);
or U984 (N_984,In_339,In_370);
and U985 (N_985,In_346,In_474);
or U986 (N_986,In_315,In_58);
or U987 (N_987,In_254,In_73);
or U988 (N_988,In_312,In_475);
nor U989 (N_989,In_491,In_6);
nor U990 (N_990,In_359,In_125);
nand U991 (N_991,In_415,In_123);
nor U992 (N_992,In_445,In_110);
or U993 (N_993,In_245,In_33);
or U994 (N_994,In_216,In_354);
nand U995 (N_995,In_311,In_29);
or U996 (N_996,In_350,In_390);
nand U997 (N_997,In_479,In_402);
nor U998 (N_998,In_188,In_370);
nand U999 (N_999,In_50,In_316);
or U1000 (N_1000,N_470,N_315);
and U1001 (N_1001,N_403,N_411);
nor U1002 (N_1002,N_467,N_492);
nand U1003 (N_1003,N_121,N_464);
and U1004 (N_1004,N_225,N_311);
nor U1005 (N_1005,N_985,N_902);
nor U1006 (N_1006,N_772,N_921);
and U1007 (N_1007,N_791,N_124);
nand U1008 (N_1008,N_858,N_859);
nor U1009 (N_1009,N_973,N_759);
nor U1010 (N_1010,N_67,N_175);
nor U1011 (N_1011,N_731,N_254);
and U1012 (N_1012,N_194,N_339);
or U1013 (N_1013,N_473,N_951);
nor U1014 (N_1014,N_910,N_104);
nor U1015 (N_1015,N_689,N_895);
nor U1016 (N_1016,N_610,N_241);
or U1017 (N_1017,N_502,N_647);
nor U1018 (N_1018,N_674,N_372);
nor U1019 (N_1019,N_265,N_938);
and U1020 (N_1020,N_710,N_656);
and U1021 (N_1021,N_586,N_946);
or U1022 (N_1022,N_163,N_595);
nand U1023 (N_1023,N_139,N_440);
nand U1024 (N_1024,N_686,N_916);
and U1025 (N_1025,N_844,N_405);
nor U1026 (N_1026,N_144,N_264);
nor U1027 (N_1027,N_80,N_118);
nor U1028 (N_1028,N_830,N_594);
or U1029 (N_1029,N_739,N_334);
nand U1030 (N_1030,N_606,N_851);
nor U1031 (N_1031,N_833,N_682);
nand U1032 (N_1032,N_788,N_101);
nor U1033 (N_1033,N_857,N_597);
nor U1034 (N_1034,N_335,N_181);
nor U1035 (N_1035,N_977,N_527);
and U1036 (N_1036,N_166,N_439);
and U1037 (N_1037,N_36,N_102);
and U1038 (N_1038,N_716,N_913);
or U1039 (N_1039,N_46,N_683);
and U1040 (N_1040,N_697,N_243);
nand U1041 (N_1041,N_185,N_336);
nand U1042 (N_1042,N_827,N_749);
or U1043 (N_1043,N_915,N_408);
or U1044 (N_1044,N_266,N_74);
and U1045 (N_1045,N_779,N_974);
nand U1046 (N_1046,N_721,N_429);
nand U1047 (N_1047,N_923,N_191);
or U1048 (N_1048,N_126,N_845);
nor U1049 (N_1049,N_333,N_309);
or U1050 (N_1050,N_360,N_249);
and U1051 (N_1051,N_592,N_542);
nand U1052 (N_1052,N_95,N_698);
nand U1053 (N_1053,N_932,N_432);
nand U1054 (N_1054,N_41,N_216);
nand U1055 (N_1055,N_862,N_338);
or U1056 (N_1056,N_744,N_695);
or U1057 (N_1057,N_169,N_217);
or U1058 (N_1058,N_724,N_624);
and U1059 (N_1059,N_110,N_39);
nand U1060 (N_1060,N_981,N_868);
and U1061 (N_1061,N_995,N_584);
nor U1062 (N_1062,N_341,N_846);
nand U1063 (N_1063,N_649,N_61);
and U1064 (N_1064,N_490,N_510);
nand U1065 (N_1065,N_785,N_406);
nor U1066 (N_1066,N_98,N_536);
nor U1067 (N_1067,N_532,N_348);
nor U1068 (N_1068,N_449,N_611);
or U1069 (N_1069,N_222,N_581);
and U1070 (N_1070,N_330,N_461);
or U1071 (N_1071,N_378,N_991);
nand U1072 (N_1072,N_525,N_703);
or U1073 (N_1073,N_706,N_601);
xor U1074 (N_1074,N_108,N_436);
and U1075 (N_1075,N_459,N_969);
nand U1076 (N_1076,N_806,N_795);
nand U1077 (N_1077,N_835,N_94);
and U1078 (N_1078,N_151,N_99);
nor U1079 (N_1079,N_896,N_906);
and U1080 (N_1080,N_920,N_312);
nor U1081 (N_1081,N_13,N_694);
nor U1082 (N_1082,N_741,N_138);
and U1083 (N_1083,N_848,N_219);
nor U1084 (N_1084,N_582,N_297);
nand U1085 (N_1085,N_445,N_456);
or U1086 (N_1086,N_351,N_38);
nand U1087 (N_1087,N_375,N_310);
nand U1088 (N_1088,N_388,N_714);
nand U1089 (N_1089,N_89,N_392);
or U1090 (N_1090,N_887,N_107);
and U1091 (N_1091,N_988,N_953);
and U1092 (N_1092,N_422,N_556);
nor U1093 (N_1093,N_593,N_786);
nor U1094 (N_1094,N_650,N_688);
nor U1095 (N_1095,N_64,N_663);
nor U1096 (N_1096,N_537,N_286);
and U1097 (N_1097,N_911,N_261);
or U1098 (N_1098,N_18,N_47);
or U1099 (N_1099,N_9,N_745);
nor U1100 (N_1100,N_277,N_267);
nor U1101 (N_1101,N_75,N_340);
nor U1102 (N_1102,N_213,N_602);
or U1103 (N_1103,N_96,N_783);
or U1104 (N_1104,N_984,N_8);
nand U1105 (N_1105,N_368,N_442);
nor U1106 (N_1106,N_155,N_454);
and U1107 (N_1107,N_834,N_924);
or U1108 (N_1108,N_979,N_894);
and U1109 (N_1109,N_78,N_416);
nor U1110 (N_1110,N_21,N_996);
nand U1111 (N_1111,N_322,N_904);
nand U1112 (N_1112,N_600,N_382);
nand U1113 (N_1113,N_994,N_162);
and U1114 (N_1114,N_952,N_245);
or U1115 (N_1115,N_747,N_947);
or U1116 (N_1116,N_59,N_573);
nor U1117 (N_1117,N_645,N_725);
or U1118 (N_1118,N_427,N_587);
and U1119 (N_1119,N_123,N_850);
and U1120 (N_1120,N_839,N_70);
or U1121 (N_1121,N_499,N_170);
or U1122 (N_1122,N_736,N_766);
and U1123 (N_1123,N_127,N_253);
or U1124 (N_1124,N_551,N_956);
nand U1125 (N_1125,N_314,N_966);
or U1126 (N_1126,N_302,N_629);
and U1127 (N_1127,N_214,N_304);
or U1128 (N_1128,N_272,N_233);
or U1129 (N_1129,N_120,N_373);
and U1130 (N_1130,N_283,N_733);
or U1131 (N_1131,N_15,N_57);
nor U1132 (N_1132,N_279,N_150);
nor U1133 (N_1133,N_62,N_660);
and U1134 (N_1134,N_521,N_812);
nand U1135 (N_1135,N_450,N_258);
or U1136 (N_1136,N_153,N_135);
or U1137 (N_1137,N_420,N_891);
nor U1138 (N_1138,N_644,N_342);
nand U1139 (N_1139,N_367,N_668);
or U1140 (N_1140,N_329,N_133);
and U1141 (N_1141,N_17,N_908);
or U1142 (N_1142,N_223,N_291);
or U1143 (N_1143,N_631,N_712);
and U1144 (N_1144,N_773,N_928);
nor U1145 (N_1145,N_52,N_705);
nor U1146 (N_1146,N_474,N_49);
nand U1147 (N_1147,N_26,N_221);
nand U1148 (N_1148,N_231,N_672);
or U1149 (N_1149,N_476,N_346);
and U1150 (N_1150,N_643,N_199);
nor U1151 (N_1151,N_805,N_489);
and U1152 (N_1152,N_305,N_798);
and U1153 (N_1153,N_33,N_414);
xor U1154 (N_1154,N_242,N_184);
or U1155 (N_1155,N_147,N_4);
nor U1156 (N_1156,N_662,N_867);
nor U1157 (N_1157,N_145,N_350);
nor U1158 (N_1158,N_178,N_114);
nand U1159 (N_1159,N_524,N_410);
xnor U1160 (N_1160,N_287,N_128);
and U1161 (N_1161,N_999,N_520);
and U1162 (N_1162,N_361,N_616);
and U1163 (N_1163,N_30,N_381);
nor U1164 (N_1164,N_978,N_327);
or U1165 (N_1165,N_929,N_500);
xor U1166 (N_1166,N_715,N_256);
nor U1167 (N_1167,N_353,N_154);
and U1168 (N_1168,N_870,N_412);
nor U1169 (N_1169,N_117,N_722);
or U1170 (N_1170,N_909,N_435);
and U1171 (N_1171,N_383,N_609);
nand U1172 (N_1172,N_797,N_577);
nor U1173 (N_1173,N_905,N_65);
or U1174 (N_1174,N_625,N_230);
nor U1175 (N_1175,N_734,N_24);
and U1176 (N_1176,N_770,N_119);
and U1177 (N_1177,N_260,N_709);
nor U1178 (N_1178,N_418,N_193);
or U1179 (N_1179,N_278,N_681);
or U1180 (N_1180,N_100,N_364);
or U1181 (N_1181,N_320,N_443);
nand U1182 (N_1182,N_5,N_93);
or U1183 (N_1183,N_399,N_822);
or U1184 (N_1184,N_192,N_478);
and U1185 (N_1185,N_83,N_501);
or U1186 (N_1186,N_180,N_452);
nor U1187 (N_1187,N_676,N_651);
and U1188 (N_1188,N_917,N_693);
nor U1189 (N_1189,N_90,N_961);
nand U1190 (N_1190,N_206,N_426);
nor U1191 (N_1191,N_876,N_702);
and U1192 (N_1192,N_247,N_345);
and U1193 (N_1193,N_636,N_479);
and U1194 (N_1194,N_990,N_817);
or U1195 (N_1195,N_972,N_482);
nand U1196 (N_1196,N_884,N_27);
or U1197 (N_1197,N_570,N_893);
nand U1198 (N_1198,N_930,N_40);
and U1199 (N_1199,N_866,N_758);
nand U1200 (N_1200,N_552,N_376);
nor U1201 (N_1201,N_246,N_14);
nand U1202 (N_1202,N_11,N_293);
nor U1203 (N_1203,N_802,N_54);
nand U1204 (N_1204,N_460,N_675);
nor U1205 (N_1205,N_269,N_664);
nor U1206 (N_1206,N_71,N_516);
nand U1207 (N_1207,N_224,N_936);
nor U1208 (N_1208,N_195,N_836);
and U1209 (N_1209,N_738,N_497);
nand U1210 (N_1210,N_438,N_547);
nand U1211 (N_1211,N_66,N_640);
or U1212 (N_1212,N_708,N_687);
and U1213 (N_1213,N_970,N_10);
or U1214 (N_1214,N_496,N_912);
nor U1215 (N_1215,N_677,N_2);
nor U1216 (N_1216,N_273,N_901);
xnor U1217 (N_1217,N_931,N_298);
or U1218 (N_1218,N_652,N_82);
nand U1219 (N_1219,N_628,N_455);
xor U1220 (N_1220,N_960,N_238);
or U1221 (N_1221,N_534,N_282);
and U1222 (N_1222,N_655,N_73);
nor U1223 (N_1223,N_769,N_829);
and U1224 (N_1224,N_183,N_453);
and U1225 (N_1225,N_539,N_630);
and U1226 (N_1226,N_515,N_240);
nand U1227 (N_1227,N_430,N_927);
and U1228 (N_1228,N_385,N_965);
nand U1229 (N_1229,N_485,N_863);
and U1230 (N_1230,N_174,N_574);
nand U1231 (N_1231,N_711,N_533);
or U1232 (N_1232,N_955,N_87);
nand U1233 (N_1233,N_717,N_782);
and U1234 (N_1234,N_255,N_374);
and U1235 (N_1235,N_818,N_634);
nor U1236 (N_1236,N_713,N_771);
and U1237 (N_1237,N_484,N_854);
and U1238 (N_1238,N_993,N_855);
nand U1239 (N_1239,N_226,N_743);
or U1240 (N_1240,N_564,N_997);
or U1241 (N_1241,N_617,N_522);
or U1242 (N_1242,N_434,N_58);
nand U1243 (N_1243,N_604,N_380);
nor U1244 (N_1244,N_718,N_431);
or U1245 (N_1245,N_111,N_641);
nor U1246 (N_1246,N_519,N_692);
nor U1247 (N_1247,N_840,N_356);
nand U1248 (N_1248,N_543,N_28);
or U1249 (N_1249,N_820,N_775);
and U1250 (N_1250,N_560,N_105);
or U1251 (N_1251,N_239,N_428);
or U1252 (N_1252,N_469,N_229);
or U1253 (N_1253,N_989,N_950);
and U1254 (N_1254,N_42,N_513);
and U1255 (N_1255,N_323,N_748);
and U1256 (N_1256,N_578,N_164);
nand U1257 (N_1257,N_419,N_402);
or U1258 (N_1258,N_122,N_842);
and U1259 (N_1259,N_699,N_88);
or U1260 (N_1260,N_136,N_171);
nor U1261 (N_1261,N_648,N_815);
nand U1262 (N_1262,N_451,N_296);
nand U1263 (N_1263,N_638,N_535);
nand U1264 (N_1264,N_826,N_987);
nor U1265 (N_1265,N_319,N_954);
or U1266 (N_1266,N_318,N_746);
nand U1267 (N_1267,N_407,N_400);
nand U1268 (N_1268,N_900,N_251);
nor U1269 (N_1269,N_262,N_415);
and U1270 (N_1270,N_276,N_557);
nor U1271 (N_1271,N_886,N_544);
or U1272 (N_1272,N_813,N_331);
nor U1273 (N_1273,N_158,N_873);
or U1274 (N_1274,N_804,N_579);
or U1275 (N_1275,N_819,N_679);
and U1276 (N_1276,N_566,N_825);
nand U1277 (N_1277,N_761,N_755);
nand U1278 (N_1278,N_131,N_390);
or U1279 (N_1279,N_723,N_498);
nor U1280 (N_1280,N_232,N_22);
nand U1281 (N_1281,N_530,N_892);
nand U1282 (N_1282,N_540,N_856);
nand U1283 (N_1283,N_160,N_665);
and U1284 (N_1284,N_250,N_732);
nor U1285 (N_1285,N_623,N_165);
nor U1286 (N_1286,N_508,N_948);
nand U1287 (N_1287,N_506,N_576);
and U1288 (N_1288,N_307,N_130);
and U1289 (N_1289,N_423,N_325);
nand U1290 (N_1290,N_861,N_349);
and U1291 (N_1291,N_959,N_794);
and U1292 (N_1292,N_37,N_878);
or U1293 (N_1293,N_462,N_409);
and U1294 (N_1294,N_3,N_86);
nand U1295 (N_1295,N_853,N_384);
nand U1296 (N_1296,N_658,N_210);
nand U1297 (N_1297,N_444,N_1);
and U1298 (N_1298,N_907,N_292);
and U1299 (N_1299,N_362,N_555);
or U1300 (N_1300,N_172,N_190);
and U1301 (N_1301,N_860,N_19);
and U1302 (N_1302,N_986,N_227);
and U1303 (N_1303,N_363,N_157);
nor U1304 (N_1304,N_550,N_719);
and U1305 (N_1305,N_531,N_808);
and U1306 (N_1306,N_271,N_754);
and U1307 (N_1307,N_607,N_197);
and U1308 (N_1308,N_899,N_53);
nand U1309 (N_1309,N_796,N_784);
or U1310 (N_1310,N_274,N_507);
and U1311 (N_1311,N_141,N_212);
nand U1312 (N_1312,N_149,N_762);
and U1313 (N_1313,N_202,N_394);
or U1314 (N_1314,N_354,N_620);
nand U1315 (N_1315,N_421,N_55);
and U1316 (N_1316,N_209,N_481);
and U1317 (N_1317,N_992,N_48);
or U1318 (N_1318,N_657,N_188);
nor U1319 (N_1319,N_919,N_34);
nand U1320 (N_1320,N_898,N_401);
and U1321 (N_1321,N_220,N_903);
or U1322 (N_1322,N_832,N_337);
nand U1323 (N_1323,N_945,N_941);
nor U1324 (N_1324,N_168,N_493);
nand U1325 (N_1325,N_182,N_653);
or U1326 (N_1326,N_437,N_847);
nor U1327 (N_1327,N_888,N_204);
or U1328 (N_1328,N_207,N_980);
nand U1329 (N_1329,N_821,N_12);
or U1330 (N_1330,N_940,N_471);
or U1331 (N_1331,N_275,N_236);
or U1332 (N_1332,N_737,N_942);
or U1333 (N_1333,N_763,N_949);
and U1334 (N_1334,N_726,N_727);
and U1335 (N_1335,N_389,N_613);
nand U1336 (N_1336,N_31,N_690);
and U1337 (N_1337,N_637,N_881);
or U1338 (N_1338,N_347,N_300);
and U1339 (N_1339,N_306,N_583);
nand U1340 (N_1340,N_106,N_387);
and U1341 (N_1341,N_205,N_370);
and U1342 (N_1342,N_729,N_523);
nor U1343 (N_1343,N_700,N_838);
or U1344 (N_1344,N_441,N_379);
and U1345 (N_1345,N_463,N_964);
nor U1346 (N_1346,N_200,N_914);
nand U1347 (N_1347,N_567,N_344);
or U1348 (N_1348,N_872,N_807);
nor U1349 (N_1349,N_962,N_377);
nor U1350 (N_1350,N_494,N_659);
and U1351 (N_1351,N_816,N_976);
and U1352 (N_1352,N_109,N_234);
nor U1353 (N_1353,N_646,N_849);
or U1354 (N_1354,N_313,N_789);
xnor U1355 (N_1355,N_303,N_257);
or U1356 (N_1356,N_596,N_397);
and U1357 (N_1357,N_837,N_517);
or U1358 (N_1358,N_684,N_841);
and U1359 (N_1359,N_541,N_7);
nor U1360 (N_1360,N_865,N_875);
nand U1361 (N_1361,N_925,N_777);
and U1362 (N_1362,N_143,N_218);
nor U1363 (N_1363,N_365,N_148);
or U1364 (N_1364,N_963,N_800);
or U1365 (N_1365,N_433,N_918);
or U1366 (N_1366,N_598,N_92);
and U1367 (N_1367,N_803,N_792);
nor U1368 (N_1368,N_186,N_720);
and U1369 (N_1369,N_167,N_572);
and U1370 (N_1370,N_288,N_869);
nor U1371 (N_1371,N_787,N_546);
nand U1372 (N_1372,N_612,N_280);
and U1373 (N_1373,N_299,N_146);
or U1374 (N_1374,N_608,N_666);
and U1375 (N_1375,N_317,N_605);
nor U1376 (N_1376,N_864,N_627);
and U1377 (N_1377,N_159,N_189);
and U1378 (N_1378,N_680,N_161);
and U1379 (N_1379,N_446,N_495);
nand U1380 (N_1380,N_132,N_760);
xor U1381 (N_1381,N_268,N_208);
and U1382 (N_1382,N_569,N_933);
nand U1383 (N_1383,N_228,N_187);
nand U1384 (N_1384,N_685,N_599);
nand U1385 (N_1385,N_44,N_874);
nor U1386 (N_1386,N_528,N_366);
and U1387 (N_1387,N_764,N_505);
and U1388 (N_1388,N_622,N_281);
or U1389 (N_1389,N_357,N_6);
nand U1390 (N_1390,N_480,N_487);
nand U1391 (N_1391,N_529,N_371);
and U1392 (N_1392,N_751,N_998);
or U1393 (N_1393,N_491,N_176);
and U1394 (N_1394,N_799,N_671);
nor U1395 (N_1395,N_369,N_767);
and U1396 (N_1396,N_575,N_558);
or U1397 (N_1397,N_295,N_79);
nor U1398 (N_1398,N_77,N_413);
nand U1399 (N_1399,N_137,N_618);
nor U1400 (N_1400,N_20,N_326);
nand U1401 (N_1401,N_386,N_248);
and U1402 (N_1402,N_880,N_25);
and U1403 (N_1403,N_934,N_824);
or U1404 (N_1404,N_404,N_568);
nand U1405 (N_1405,N_244,N_958);
nor U1406 (N_1406,N_512,N_32);
nor U1407 (N_1407,N_316,N_968);
nand U1408 (N_1408,N_50,N_554);
and U1409 (N_1409,N_526,N_790);
nor U1410 (N_1410,N_701,N_707);
nor U1411 (N_1411,N_943,N_559);
or U1412 (N_1412,N_571,N_81);
and U1413 (N_1413,N_937,N_939);
nand U1414 (N_1414,N_778,N_84);
nand U1415 (N_1415,N_670,N_967);
or U1416 (N_1416,N_425,N_704);
nand U1417 (N_1417,N_639,N_56);
nor U1418 (N_1418,N_177,N_285);
nor U1419 (N_1419,N_179,N_343);
nor U1420 (N_1420,N_774,N_753);
and U1421 (N_1421,N_538,N_63);
or U1422 (N_1422,N_152,N_395);
and U1423 (N_1423,N_211,N_752);
nor U1424 (N_1424,N_294,N_457);
or U1425 (N_1425,N_843,N_926);
nand U1426 (N_1426,N_691,N_877);
or U1427 (N_1427,N_669,N_308);
nand U1428 (N_1428,N_475,N_398);
nand U1429 (N_1429,N_793,N_588);
or U1430 (N_1430,N_140,N_466);
nor U1431 (N_1431,N_352,N_545);
nor U1432 (N_1432,N_518,N_284);
nand U1433 (N_1433,N_831,N_614);
nor U1434 (N_1434,N_673,N_391);
nor U1435 (N_1435,N_129,N_447);
and U1436 (N_1436,N_201,N_68);
nor U1437 (N_1437,N_134,N_615);
nand U1438 (N_1438,N_728,N_603);
or U1439 (N_1439,N_173,N_871);
nand U1440 (N_1440,N_448,N_51);
nand U1441 (N_1441,N_632,N_35);
or U1442 (N_1442,N_944,N_116);
or U1443 (N_1443,N_626,N_621);
or U1444 (N_1444,N_883,N_112);
or U1445 (N_1445,N_971,N_879);
or U1446 (N_1446,N_359,N_811);
nor U1447 (N_1447,N_115,N_355);
nor U1448 (N_1448,N_29,N_503);
nor U1449 (N_1449,N_203,N_424);
nand U1450 (N_1450,N_661,N_321);
or U1451 (N_1451,N_483,N_156);
nor U1452 (N_1452,N_263,N_565);
or U1453 (N_1453,N_982,N_509);
nand U1454 (N_1454,N_468,N_619);
and U1455 (N_1455,N_765,N_562);
or U1456 (N_1456,N_776,N_43);
and U1457 (N_1457,N_215,N_142);
nor U1458 (N_1458,N_72,N_561);
and U1459 (N_1459,N_486,N_514);
and U1460 (N_1460,N_781,N_91);
or U1461 (N_1461,N_125,N_580);
nor U1462 (N_1462,N_548,N_504);
nand U1463 (N_1463,N_259,N_890);
and U1464 (N_1464,N_196,N_740);
and U1465 (N_1465,N_563,N_730);
or U1466 (N_1466,N_957,N_332);
nand U1467 (N_1467,N_16,N_897);
or U1468 (N_1468,N_750,N_678);
and U1469 (N_1469,N_396,N_696);
nor U1470 (N_1470,N_983,N_0);
and U1471 (N_1471,N_809,N_301);
nand U1472 (N_1472,N_654,N_198);
and U1473 (N_1473,N_417,N_103);
or U1474 (N_1474,N_810,N_60);
nand U1475 (N_1475,N_76,N_113);
nor U1476 (N_1476,N_922,N_472);
and U1477 (N_1477,N_828,N_252);
nor U1478 (N_1478,N_289,N_328);
and U1479 (N_1479,N_882,N_590);
nor U1480 (N_1480,N_735,N_801);
nand U1481 (N_1481,N_97,N_235);
nand U1482 (N_1482,N_465,N_756);
or U1483 (N_1483,N_642,N_85);
nor U1484 (N_1484,N_511,N_852);
nor U1485 (N_1485,N_270,N_591);
nand U1486 (N_1486,N_935,N_814);
nand U1487 (N_1487,N_885,N_237);
nor U1488 (N_1488,N_780,N_742);
or U1489 (N_1489,N_458,N_823);
nand U1490 (N_1490,N_69,N_889);
nand U1491 (N_1491,N_488,N_975);
or U1492 (N_1492,N_585,N_633);
and U1493 (N_1493,N_358,N_290);
nand U1494 (N_1494,N_667,N_635);
nand U1495 (N_1495,N_477,N_589);
xnor U1496 (N_1496,N_393,N_549);
nand U1497 (N_1497,N_768,N_553);
nand U1498 (N_1498,N_23,N_45);
nor U1499 (N_1499,N_324,N_757);
nand U1500 (N_1500,N_945,N_519);
nand U1501 (N_1501,N_397,N_873);
nand U1502 (N_1502,N_680,N_281);
nor U1503 (N_1503,N_141,N_423);
or U1504 (N_1504,N_767,N_102);
nor U1505 (N_1505,N_472,N_145);
nor U1506 (N_1506,N_535,N_423);
nor U1507 (N_1507,N_914,N_388);
or U1508 (N_1508,N_351,N_436);
or U1509 (N_1509,N_627,N_391);
nand U1510 (N_1510,N_851,N_272);
or U1511 (N_1511,N_988,N_499);
nor U1512 (N_1512,N_841,N_192);
or U1513 (N_1513,N_784,N_789);
nor U1514 (N_1514,N_399,N_268);
nor U1515 (N_1515,N_994,N_851);
and U1516 (N_1516,N_4,N_764);
and U1517 (N_1517,N_159,N_46);
or U1518 (N_1518,N_452,N_183);
and U1519 (N_1519,N_541,N_677);
and U1520 (N_1520,N_414,N_569);
nand U1521 (N_1521,N_493,N_309);
nand U1522 (N_1522,N_180,N_712);
and U1523 (N_1523,N_453,N_848);
nor U1524 (N_1524,N_953,N_33);
and U1525 (N_1525,N_369,N_779);
nand U1526 (N_1526,N_301,N_929);
and U1527 (N_1527,N_276,N_581);
nor U1528 (N_1528,N_952,N_820);
and U1529 (N_1529,N_182,N_780);
nor U1530 (N_1530,N_912,N_224);
or U1531 (N_1531,N_221,N_134);
or U1532 (N_1532,N_274,N_389);
or U1533 (N_1533,N_642,N_886);
nand U1534 (N_1534,N_125,N_530);
and U1535 (N_1535,N_841,N_354);
and U1536 (N_1536,N_979,N_30);
and U1537 (N_1537,N_809,N_766);
and U1538 (N_1538,N_931,N_35);
or U1539 (N_1539,N_985,N_513);
nor U1540 (N_1540,N_640,N_147);
and U1541 (N_1541,N_20,N_834);
and U1542 (N_1542,N_341,N_704);
nand U1543 (N_1543,N_548,N_675);
or U1544 (N_1544,N_907,N_868);
nor U1545 (N_1545,N_74,N_476);
nand U1546 (N_1546,N_401,N_458);
nand U1547 (N_1547,N_825,N_899);
nor U1548 (N_1548,N_900,N_149);
nor U1549 (N_1549,N_853,N_439);
nor U1550 (N_1550,N_354,N_131);
nand U1551 (N_1551,N_764,N_200);
or U1552 (N_1552,N_509,N_645);
or U1553 (N_1553,N_183,N_473);
and U1554 (N_1554,N_348,N_393);
nor U1555 (N_1555,N_366,N_240);
and U1556 (N_1556,N_562,N_727);
or U1557 (N_1557,N_112,N_167);
or U1558 (N_1558,N_531,N_885);
nor U1559 (N_1559,N_867,N_543);
and U1560 (N_1560,N_129,N_93);
nor U1561 (N_1561,N_657,N_848);
xnor U1562 (N_1562,N_946,N_658);
xor U1563 (N_1563,N_260,N_333);
nor U1564 (N_1564,N_252,N_475);
or U1565 (N_1565,N_457,N_719);
nor U1566 (N_1566,N_388,N_179);
nor U1567 (N_1567,N_909,N_234);
nor U1568 (N_1568,N_35,N_106);
and U1569 (N_1569,N_970,N_609);
or U1570 (N_1570,N_690,N_134);
or U1571 (N_1571,N_387,N_71);
and U1572 (N_1572,N_332,N_135);
and U1573 (N_1573,N_105,N_685);
nand U1574 (N_1574,N_50,N_6);
and U1575 (N_1575,N_564,N_484);
nor U1576 (N_1576,N_182,N_736);
or U1577 (N_1577,N_474,N_545);
and U1578 (N_1578,N_680,N_555);
or U1579 (N_1579,N_519,N_726);
and U1580 (N_1580,N_958,N_632);
or U1581 (N_1581,N_820,N_365);
or U1582 (N_1582,N_335,N_635);
nand U1583 (N_1583,N_284,N_10);
nand U1584 (N_1584,N_104,N_827);
xor U1585 (N_1585,N_136,N_526);
or U1586 (N_1586,N_831,N_53);
or U1587 (N_1587,N_190,N_278);
or U1588 (N_1588,N_660,N_160);
nand U1589 (N_1589,N_708,N_155);
or U1590 (N_1590,N_89,N_337);
and U1591 (N_1591,N_217,N_957);
or U1592 (N_1592,N_777,N_150);
nand U1593 (N_1593,N_882,N_471);
and U1594 (N_1594,N_272,N_402);
or U1595 (N_1595,N_175,N_739);
and U1596 (N_1596,N_784,N_647);
or U1597 (N_1597,N_792,N_708);
and U1598 (N_1598,N_586,N_1);
nor U1599 (N_1599,N_848,N_159);
and U1600 (N_1600,N_854,N_277);
nand U1601 (N_1601,N_235,N_362);
and U1602 (N_1602,N_316,N_224);
or U1603 (N_1603,N_96,N_700);
and U1604 (N_1604,N_813,N_51);
nor U1605 (N_1605,N_128,N_48);
or U1606 (N_1606,N_320,N_822);
and U1607 (N_1607,N_807,N_683);
nand U1608 (N_1608,N_283,N_456);
nand U1609 (N_1609,N_134,N_688);
nor U1610 (N_1610,N_981,N_610);
and U1611 (N_1611,N_767,N_46);
and U1612 (N_1612,N_295,N_637);
xor U1613 (N_1613,N_843,N_421);
nor U1614 (N_1614,N_324,N_368);
nand U1615 (N_1615,N_189,N_559);
and U1616 (N_1616,N_538,N_472);
nand U1617 (N_1617,N_186,N_603);
nand U1618 (N_1618,N_286,N_773);
nand U1619 (N_1619,N_441,N_741);
and U1620 (N_1620,N_293,N_912);
and U1621 (N_1621,N_103,N_421);
or U1622 (N_1622,N_497,N_564);
or U1623 (N_1623,N_177,N_420);
nor U1624 (N_1624,N_519,N_995);
nor U1625 (N_1625,N_585,N_549);
nor U1626 (N_1626,N_770,N_317);
and U1627 (N_1627,N_745,N_830);
nor U1628 (N_1628,N_797,N_885);
or U1629 (N_1629,N_3,N_672);
and U1630 (N_1630,N_44,N_550);
or U1631 (N_1631,N_622,N_790);
and U1632 (N_1632,N_149,N_544);
nor U1633 (N_1633,N_228,N_431);
and U1634 (N_1634,N_386,N_238);
and U1635 (N_1635,N_432,N_785);
nand U1636 (N_1636,N_769,N_15);
nor U1637 (N_1637,N_734,N_105);
nor U1638 (N_1638,N_995,N_293);
nor U1639 (N_1639,N_992,N_136);
or U1640 (N_1640,N_226,N_973);
and U1641 (N_1641,N_575,N_59);
nand U1642 (N_1642,N_134,N_968);
and U1643 (N_1643,N_555,N_662);
and U1644 (N_1644,N_383,N_724);
or U1645 (N_1645,N_662,N_120);
xnor U1646 (N_1646,N_17,N_482);
nand U1647 (N_1647,N_443,N_812);
and U1648 (N_1648,N_5,N_906);
and U1649 (N_1649,N_510,N_93);
nor U1650 (N_1650,N_877,N_398);
nand U1651 (N_1651,N_773,N_851);
or U1652 (N_1652,N_841,N_94);
or U1653 (N_1653,N_260,N_462);
or U1654 (N_1654,N_149,N_538);
nor U1655 (N_1655,N_841,N_138);
nor U1656 (N_1656,N_619,N_623);
nor U1657 (N_1657,N_474,N_723);
or U1658 (N_1658,N_92,N_229);
and U1659 (N_1659,N_479,N_265);
and U1660 (N_1660,N_342,N_758);
nand U1661 (N_1661,N_120,N_917);
and U1662 (N_1662,N_368,N_692);
nor U1663 (N_1663,N_184,N_746);
nand U1664 (N_1664,N_632,N_860);
or U1665 (N_1665,N_643,N_19);
and U1666 (N_1666,N_529,N_906);
nand U1667 (N_1667,N_575,N_911);
nor U1668 (N_1668,N_350,N_279);
or U1669 (N_1669,N_631,N_652);
and U1670 (N_1670,N_851,N_212);
nor U1671 (N_1671,N_874,N_711);
and U1672 (N_1672,N_823,N_95);
and U1673 (N_1673,N_20,N_963);
nand U1674 (N_1674,N_129,N_176);
nand U1675 (N_1675,N_667,N_863);
or U1676 (N_1676,N_566,N_56);
and U1677 (N_1677,N_462,N_723);
or U1678 (N_1678,N_676,N_547);
nand U1679 (N_1679,N_337,N_701);
nor U1680 (N_1680,N_142,N_275);
nor U1681 (N_1681,N_68,N_533);
or U1682 (N_1682,N_803,N_419);
nor U1683 (N_1683,N_793,N_630);
and U1684 (N_1684,N_662,N_615);
nor U1685 (N_1685,N_446,N_110);
nor U1686 (N_1686,N_495,N_223);
nor U1687 (N_1687,N_351,N_286);
and U1688 (N_1688,N_816,N_50);
nand U1689 (N_1689,N_386,N_937);
nor U1690 (N_1690,N_265,N_676);
nand U1691 (N_1691,N_8,N_457);
and U1692 (N_1692,N_585,N_823);
and U1693 (N_1693,N_564,N_730);
and U1694 (N_1694,N_616,N_438);
and U1695 (N_1695,N_779,N_436);
nor U1696 (N_1696,N_327,N_917);
and U1697 (N_1697,N_860,N_375);
or U1698 (N_1698,N_828,N_746);
and U1699 (N_1699,N_688,N_916);
nor U1700 (N_1700,N_538,N_707);
nand U1701 (N_1701,N_729,N_13);
or U1702 (N_1702,N_768,N_6);
nand U1703 (N_1703,N_758,N_339);
or U1704 (N_1704,N_103,N_414);
or U1705 (N_1705,N_50,N_895);
or U1706 (N_1706,N_635,N_56);
and U1707 (N_1707,N_72,N_277);
nand U1708 (N_1708,N_258,N_848);
nor U1709 (N_1709,N_884,N_885);
or U1710 (N_1710,N_167,N_418);
and U1711 (N_1711,N_486,N_672);
and U1712 (N_1712,N_24,N_324);
or U1713 (N_1713,N_627,N_683);
nand U1714 (N_1714,N_861,N_521);
and U1715 (N_1715,N_323,N_35);
nand U1716 (N_1716,N_326,N_31);
and U1717 (N_1717,N_673,N_61);
nor U1718 (N_1718,N_117,N_761);
or U1719 (N_1719,N_521,N_351);
nor U1720 (N_1720,N_266,N_487);
or U1721 (N_1721,N_364,N_797);
and U1722 (N_1722,N_929,N_745);
nor U1723 (N_1723,N_677,N_455);
nor U1724 (N_1724,N_102,N_702);
nor U1725 (N_1725,N_527,N_804);
or U1726 (N_1726,N_566,N_567);
or U1727 (N_1727,N_245,N_232);
nor U1728 (N_1728,N_451,N_419);
nor U1729 (N_1729,N_34,N_24);
nand U1730 (N_1730,N_237,N_324);
or U1731 (N_1731,N_805,N_963);
nor U1732 (N_1732,N_638,N_542);
nand U1733 (N_1733,N_557,N_584);
or U1734 (N_1734,N_178,N_213);
nand U1735 (N_1735,N_69,N_578);
or U1736 (N_1736,N_903,N_890);
or U1737 (N_1737,N_82,N_177);
nand U1738 (N_1738,N_556,N_179);
or U1739 (N_1739,N_30,N_194);
and U1740 (N_1740,N_388,N_639);
or U1741 (N_1741,N_670,N_68);
nand U1742 (N_1742,N_770,N_867);
or U1743 (N_1743,N_653,N_98);
and U1744 (N_1744,N_782,N_722);
or U1745 (N_1745,N_872,N_41);
nand U1746 (N_1746,N_442,N_780);
or U1747 (N_1747,N_169,N_247);
nand U1748 (N_1748,N_579,N_812);
or U1749 (N_1749,N_770,N_953);
xnor U1750 (N_1750,N_576,N_811);
nand U1751 (N_1751,N_603,N_658);
nor U1752 (N_1752,N_566,N_852);
nor U1753 (N_1753,N_20,N_102);
nand U1754 (N_1754,N_226,N_777);
nor U1755 (N_1755,N_337,N_54);
nand U1756 (N_1756,N_638,N_410);
nand U1757 (N_1757,N_429,N_956);
and U1758 (N_1758,N_572,N_785);
nand U1759 (N_1759,N_893,N_378);
nor U1760 (N_1760,N_279,N_467);
nor U1761 (N_1761,N_371,N_848);
nand U1762 (N_1762,N_634,N_606);
or U1763 (N_1763,N_854,N_518);
nor U1764 (N_1764,N_663,N_735);
nor U1765 (N_1765,N_200,N_286);
or U1766 (N_1766,N_354,N_837);
nor U1767 (N_1767,N_849,N_272);
nor U1768 (N_1768,N_632,N_32);
and U1769 (N_1769,N_928,N_869);
and U1770 (N_1770,N_540,N_219);
or U1771 (N_1771,N_922,N_69);
nand U1772 (N_1772,N_582,N_400);
and U1773 (N_1773,N_530,N_262);
nor U1774 (N_1774,N_476,N_392);
and U1775 (N_1775,N_181,N_797);
and U1776 (N_1776,N_555,N_244);
or U1777 (N_1777,N_833,N_119);
nand U1778 (N_1778,N_532,N_323);
nand U1779 (N_1779,N_811,N_850);
nand U1780 (N_1780,N_772,N_304);
nor U1781 (N_1781,N_421,N_25);
or U1782 (N_1782,N_136,N_920);
and U1783 (N_1783,N_181,N_664);
nor U1784 (N_1784,N_521,N_378);
and U1785 (N_1785,N_125,N_897);
nand U1786 (N_1786,N_816,N_946);
or U1787 (N_1787,N_276,N_127);
or U1788 (N_1788,N_649,N_757);
and U1789 (N_1789,N_0,N_714);
and U1790 (N_1790,N_397,N_583);
nand U1791 (N_1791,N_810,N_212);
nand U1792 (N_1792,N_26,N_619);
nor U1793 (N_1793,N_720,N_271);
nor U1794 (N_1794,N_512,N_102);
nand U1795 (N_1795,N_413,N_118);
nand U1796 (N_1796,N_973,N_709);
and U1797 (N_1797,N_282,N_864);
nor U1798 (N_1798,N_464,N_133);
and U1799 (N_1799,N_52,N_922);
nand U1800 (N_1800,N_389,N_621);
nor U1801 (N_1801,N_877,N_881);
nor U1802 (N_1802,N_559,N_326);
or U1803 (N_1803,N_981,N_879);
and U1804 (N_1804,N_792,N_884);
and U1805 (N_1805,N_186,N_77);
or U1806 (N_1806,N_241,N_707);
and U1807 (N_1807,N_507,N_601);
or U1808 (N_1808,N_408,N_486);
nand U1809 (N_1809,N_414,N_963);
nand U1810 (N_1810,N_190,N_697);
and U1811 (N_1811,N_147,N_196);
and U1812 (N_1812,N_579,N_775);
nor U1813 (N_1813,N_510,N_726);
nand U1814 (N_1814,N_788,N_387);
and U1815 (N_1815,N_866,N_294);
or U1816 (N_1816,N_239,N_26);
or U1817 (N_1817,N_636,N_895);
nor U1818 (N_1818,N_304,N_637);
and U1819 (N_1819,N_678,N_933);
nand U1820 (N_1820,N_238,N_442);
and U1821 (N_1821,N_997,N_929);
or U1822 (N_1822,N_347,N_278);
or U1823 (N_1823,N_240,N_269);
or U1824 (N_1824,N_253,N_281);
or U1825 (N_1825,N_68,N_790);
and U1826 (N_1826,N_58,N_680);
nand U1827 (N_1827,N_777,N_996);
or U1828 (N_1828,N_915,N_522);
and U1829 (N_1829,N_519,N_26);
and U1830 (N_1830,N_189,N_400);
nand U1831 (N_1831,N_4,N_260);
or U1832 (N_1832,N_959,N_786);
or U1833 (N_1833,N_555,N_971);
and U1834 (N_1834,N_68,N_83);
and U1835 (N_1835,N_207,N_72);
and U1836 (N_1836,N_723,N_518);
and U1837 (N_1837,N_317,N_84);
and U1838 (N_1838,N_773,N_58);
or U1839 (N_1839,N_215,N_719);
and U1840 (N_1840,N_403,N_705);
nor U1841 (N_1841,N_908,N_621);
or U1842 (N_1842,N_108,N_674);
or U1843 (N_1843,N_384,N_805);
nand U1844 (N_1844,N_832,N_240);
nand U1845 (N_1845,N_609,N_500);
and U1846 (N_1846,N_523,N_583);
and U1847 (N_1847,N_561,N_291);
nor U1848 (N_1848,N_535,N_664);
nor U1849 (N_1849,N_576,N_953);
nor U1850 (N_1850,N_562,N_445);
nand U1851 (N_1851,N_431,N_725);
or U1852 (N_1852,N_473,N_828);
nor U1853 (N_1853,N_357,N_410);
nand U1854 (N_1854,N_904,N_5);
nor U1855 (N_1855,N_946,N_859);
or U1856 (N_1856,N_6,N_848);
nor U1857 (N_1857,N_218,N_735);
nand U1858 (N_1858,N_628,N_939);
nand U1859 (N_1859,N_149,N_976);
nor U1860 (N_1860,N_806,N_369);
and U1861 (N_1861,N_272,N_873);
and U1862 (N_1862,N_975,N_360);
and U1863 (N_1863,N_124,N_359);
nand U1864 (N_1864,N_847,N_701);
nand U1865 (N_1865,N_937,N_421);
or U1866 (N_1866,N_282,N_679);
and U1867 (N_1867,N_216,N_998);
or U1868 (N_1868,N_330,N_592);
nor U1869 (N_1869,N_803,N_696);
nand U1870 (N_1870,N_902,N_409);
xor U1871 (N_1871,N_847,N_664);
and U1872 (N_1872,N_529,N_265);
and U1873 (N_1873,N_566,N_541);
or U1874 (N_1874,N_376,N_616);
nand U1875 (N_1875,N_7,N_880);
nor U1876 (N_1876,N_659,N_165);
nand U1877 (N_1877,N_57,N_981);
and U1878 (N_1878,N_58,N_35);
or U1879 (N_1879,N_358,N_537);
and U1880 (N_1880,N_956,N_7);
nand U1881 (N_1881,N_993,N_518);
nand U1882 (N_1882,N_961,N_434);
nand U1883 (N_1883,N_677,N_327);
or U1884 (N_1884,N_3,N_429);
and U1885 (N_1885,N_632,N_600);
and U1886 (N_1886,N_364,N_433);
nand U1887 (N_1887,N_708,N_866);
nand U1888 (N_1888,N_808,N_569);
nand U1889 (N_1889,N_387,N_315);
nand U1890 (N_1890,N_239,N_643);
nand U1891 (N_1891,N_749,N_382);
nand U1892 (N_1892,N_634,N_771);
nor U1893 (N_1893,N_620,N_206);
or U1894 (N_1894,N_226,N_373);
nand U1895 (N_1895,N_450,N_249);
and U1896 (N_1896,N_507,N_330);
or U1897 (N_1897,N_925,N_179);
nor U1898 (N_1898,N_545,N_661);
or U1899 (N_1899,N_553,N_31);
nor U1900 (N_1900,N_645,N_232);
and U1901 (N_1901,N_141,N_314);
nand U1902 (N_1902,N_490,N_726);
nand U1903 (N_1903,N_850,N_444);
and U1904 (N_1904,N_67,N_860);
nand U1905 (N_1905,N_51,N_399);
or U1906 (N_1906,N_107,N_59);
nor U1907 (N_1907,N_568,N_549);
nand U1908 (N_1908,N_783,N_204);
nand U1909 (N_1909,N_536,N_262);
and U1910 (N_1910,N_492,N_799);
and U1911 (N_1911,N_475,N_325);
and U1912 (N_1912,N_39,N_998);
and U1913 (N_1913,N_501,N_107);
or U1914 (N_1914,N_235,N_424);
and U1915 (N_1915,N_343,N_58);
nand U1916 (N_1916,N_124,N_577);
nor U1917 (N_1917,N_389,N_671);
and U1918 (N_1918,N_417,N_31);
or U1919 (N_1919,N_853,N_885);
or U1920 (N_1920,N_793,N_858);
or U1921 (N_1921,N_809,N_718);
and U1922 (N_1922,N_865,N_985);
and U1923 (N_1923,N_33,N_179);
and U1924 (N_1924,N_652,N_660);
or U1925 (N_1925,N_803,N_555);
nor U1926 (N_1926,N_660,N_784);
nor U1927 (N_1927,N_828,N_713);
nand U1928 (N_1928,N_670,N_339);
nor U1929 (N_1929,N_658,N_75);
or U1930 (N_1930,N_605,N_837);
and U1931 (N_1931,N_314,N_818);
or U1932 (N_1932,N_543,N_203);
or U1933 (N_1933,N_277,N_193);
nand U1934 (N_1934,N_31,N_903);
nand U1935 (N_1935,N_544,N_748);
and U1936 (N_1936,N_291,N_156);
nor U1937 (N_1937,N_157,N_372);
nor U1938 (N_1938,N_1,N_376);
nand U1939 (N_1939,N_236,N_934);
nand U1940 (N_1940,N_958,N_916);
nand U1941 (N_1941,N_682,N_3);
or U1942 (N_1942,N_240,N_697);
or U1943 (N_1943,N_179,N_959);
nand U1944 (N_1944,N_881,N_15);
nor U1945 (N_1945,N_271,N_254);
and U1946 (N_1946,N_197,N_830);
and U1947 (N_1947,N_905,N_350);
nand U1948 (N_1948,N_462,N_922);
or U1949 (N_1949,N_914,N_49);
and U1950 (N_1950,N_902,N_551);
and U1951 (N_1951,N_696,N_722);
and U1952 (N_1952,N_961,N_900);
nor U1953 (N_1953,N_840,N_427);
or U1954 (N_1954,N_247,N_786);
nand U1955 (N_1955,N_709,N_59);
and U1956 (N_1956,N_309,N_216);
nor U1957 (N_1957,N_538,N_286);
nor U1958 (N_1958,N_112,N_8);
nand U1959 (N_1959,N_874,N_700);
nand U1960 (N_1960,N_56,N_781);
or U1961 (N_1961,N_839,N_758);
and U1962 (N_1962,N_462,N_921);
nand U1963 (N_1963,N_309,N_642);
and U1964 (N_1964,N_553,N_933);
nor U1965 (N_1965,N_201,N_943);
nand U1966 (N_1966,N_564,N_411);
nand U1967 (N_1967,N_817,N_627);
nor U1968 (N_1968,N_988,N_320);
and U1969 (N_1969,N_256,N_580);
or U1970 (N_1970,N_614,N_230);
nand U1971 (N_1971,N_824,N_143);
nor U1972 (N_1972,N_798,N_543);
xnor U1973 (N_1973,N_757,N_346);
and U1974 (N_1974,N_977,N_985);
nor U1975 (N_1975,N_381,N_173);
or U1976 (N_1976,N_615,N_343);
nand U1977 (N_1977,N_905,N_229);
and U1978 (N_1978,N_901,N_61);
nor U1979 (N_1979,N_395,N_128);
and U1980 (N_1980,N_180,N_885);
nor U1981 (N_1981,N_359,N_473);
nand U1982 (N_1982,N_651,N_117);
nor U1983 (N_1983,N_795,N_945);
or U1984 (N_1984,N_730,N_614);
and U1985 (N_1985,N_15,N_525);
nor U1986 (N_1986,N_603,N_859);
nand U1987 (N_1987,N_555,N_146);
and U1988 (N_1988,N_830,N_98);
nand U1989 (N_1989,N_788,N_444);
and U1990 (N_1990,N_886,N_990);
and U1991 (N_1991,N_84,N_551);
or U1992 (N_1992,N_450,N_371);
or U1993 (N_1993,N_200,N_795);
and U1994 (N_1994,N_698,N_788);
nor U1995 (N_1995,N_192,N_906);
and U1996 (N_1996,N_906,N_276);
or U1997 (N_1997,N_588,N_707);
and U1998 (N_1998,N_83,N_619);
nand U1999 (N_1999,N_949,N_518);
nor U2000 (N_2000,N_1405,N_1021);
nand U2001 (N_2001,N_1478,N_1709);
nand U2002 (N_2002,N_1221,N_1477);
or U2003 (N_2003,N_1208,N_1545);
nand U2004 (N_2004,N_1307,N_1998);
nor U2005 (N_2005,N_1304,N_1199);
or U2006 (N_2006,N_1329,N_1419);
nor U2007 (N_2007,N_1799,N_1993);
and U2008 (N_2008,N_1507,N_1636);
or U2009 (N_2009,N_1339,N_1809);
nand U2010 (N_2010,N_1785,N_1886);
or U2011 (N_2011,N_1236,N_1291);
nor U2012 (N_2012,N_1510,N_1093);
xor U2013 (N_2013,N_1613,N_1549);
nor U2014 (N_2014,N_1472,N_1318);
xnor U2015 (N_2015,N_1760,N_1125);
and U2016 (N_2016,N_1527,N_1508);
xor U2017 (N_2017,N_1128,N_1045);
nor U2018 (N_2018,N_1495,N_1355);
or U2019 (N_2019,N_1571,N_1747);
or U2020 (N_2020,N_1109,N_1987);
nand U2021 (N_2021,N_1787,N_1780);
or U2022 (N_2022,N_1628,N_1750);
nor U2023 (N_2023,N_1317,N_1281);
nand U2024 (N_2024,N_1248,N_1627);
and U2025 (N_2025,N_1389,N_1937);
nand U2026 (N_2026,N_1845,N_1500);
and U2027 (N_2027,N_1397,N_1222);
nand U2028 (N_2028,N_1270,N_1009);
and U2029 (N_2029,N_1618,N_1438);
nand U2030 (N_2030,N_1942,N_1046);
nor U2031 (N_2031,N_1480,N_1724);
nand U2032 (N_2032,N_1184,N_1385);
or U2033 (N_2033,N_1583,N_1399);
or U2034 (N_2034,N_1548,N_1604);
and U2035 (N_2035,N_1062,N_1080);
or U2036 (N_2036,N_1421,N_1052);
nor U2037 (N_2037,N_1297,N_1567);
and U2038 (N_2038,N_1227,N_1663);
nor U2039 (N_2039,N_1349,N_1955);
and U2040 (N_2040,N_1978,N_1516);
and U2041 (N_2041,N_1686,N_1912);
nor U2042 (N_2042,N_1816,N_1833);
and U2043 (N_2043,N_1773,N_1883);
nor U2044 (N_2044,N_1517,N_1007);
or U2045 (N_2045,N_1559,N_1782);
nand U2046 (N_2046,N_1447,N_1532);
or U2047 (N_2047,N_1884,N_1569);
and U2048 (N_2048,N_1319,N_1084);
nand U2049 (N_2049,N_1757,N_1017);
nor U2050 (N_2050,N_1939,N_1296);
nor U2051 (N_2051,N_1505,N_1759);
or U2052 (N_2052,N_1988,N_1154);
nand U2053 (N_2053,N_1589,N_1908);
nand U2054 (N_2054,N_1336,N_1458);
and U2055 (N_2055,N_1768,N_1704);
nor U2056 (N_2056,N_1441,N_1269);
or U2057 (N_2057,N_1214,N_1538);
nor U2058 (N_2058,N_1829,N_1846);
or U2059 (N_2059,N_1308,N_1578);
nand U2060 (N_2060,N_1032,N_1598);
nor U2061 (N_2061,N_1136,N_1014);
nor U2062 (N_2062,N_1645,N_1177);
and U2063 (N_2063,N_1534,N_1863);
nor U2064 (N_2064,N_1058,N_1079);
and U2065 (N_2065,N_1370,N_1034);
nand U2066 (N_2066,N_1960,N_1675);
nor U2067 (N_2067,N_1376,N_1940);
nor U2068 (N_2068,N_1900,N_1742);
nand U2069 (N_2069,N_1865,N_1762);
nor U2070 (N_2070,N_1387,N_1842);
and U2071 (N_2071,N_1346,N_1660);
nand U2072 (N_2072,N_1999,N_1666);
nor U2073 (N_2073,N_1117,N_1891);
or U2074 (N_2074,N_1005,N_1330);
and U2075 (N_2075,N_1076,N_1374);
or U2076 (N_2076,N_1526,N_1228);
nor U2077 (N_2077,N_1202,N_1022);
nor U2078 (N_2078,N_1655,N_1169);
nor U2079 (N_2079,N_1778,N_1276);
or U2080 (N_2080,N_1909,N_1033);
nand U2081 (N_2081,N_1887,N_1681);
nor U2082 (N_2082,N_1649,N_1662);
nor U2083 (N_2083,N_1607,N_1118);
nor U2084 (N_2084,N_1849,N_1862);
or U2085 (N_2085,N_1588,N_1298);
or U2086 (N_2086,N_1879,N_1889);
or U2087 (N_2087,N_1739,N_1489);
and U2088 (N_2088,N_1707,N_1338);
nand U2089 (N_2089,N_1104,N_1556);
or U2090 (N_2090,N_1257,N_1623);
nand U2091 (N_2091,N_1520,N_1239);
and U2092 (N_2092,N_1486,N_1568);
and U2093 (N_2093,N_1540,N_1688);
and U2094 (N_2094,N_1203,N_1553);
and U2095 (N_2095,N_1935,N_1373);
or U2096 (N_2096,N_1931,N_1929);
nand U2097 (N_2097,N_1766,N_1752);
nor U2098 (N_2098,N_1431,N_1456);
or U2099 (N_2099,N_1087,N_1819);
nand U2100 (N_2100,N_1906,N_1954);
and U2101 (N_2101,N_1643,N_1173);
nand U2102 (N_2102,N_1936,N_1351);
and U2103 (N_2103,N_1753,N_1190);
and U2104 (N_2104,N_1521,N_1689);
nand U2105 (N_2105,N_1619,N_1719);
or U2106 (N_2106,N_1452,N_1947);
and U2107 (N_2107,N_1986,N_1449);
nand U2108 (N_2108,N_1271,N_1562);
nand U2109 (N_2109,N_1915,N_1841);
or U2110 (N_2110,N_1678,N_1745);
and U2111 (N_2111,N_1484,N_1043);
nand U2112 (N_2112,N_1383,N_1606);
nand U2113 (N_2113,N_1275,N_1357);
nand U2114 (N_2114,N_1334,N_1180);
and U2115 (N_2115,N_1566,N_1798);
nor U2116 (N_2116,N_1868,N_1953);
nor U2117 (N_2117,N_1377,N_1610);
and U2118 (N_2118,N_1493,N_1812);
or U2119 (N_2119,N_1916,N_1145);
or U2120 (N_2120,N_1783,N_1235);
or U2121 (N_2121,N_1800,N_1198);
or U2122 (N_2122,N_1866,N_1386);
nand U2123 (N_2123,N_1831,N_1302);
or U2124 (N_2124,N_1337,N_1086);
nor U2125 (N_2125,N_1146,N_1544);
nand U2126 (N_2126,N_1871,N_1226);
nor U2127 (N_2127,N_1167,N_1204);
nor U2128 (N_2128,N_1608,N_1354);
or U2129 (N_2129,N_1706,N_1335);
nor U2130 (N_2130,N_1843,N_1280);
and U2131 (N_2131,N_1633,N_1331);
or U2132 (N_2132,N_1876,N_1844);
and U2133 (N_2133,N_1151,N_1344);
and U2134 (N_2134,N_1153,N_1744);
and U2135 (N_2135,N_1122,N_1168);
nand U2136 (N_2136,N_1856,N_1013);
and U2137 (N_2137,N_1664,N_1127);
nand U2138 (N_2138,N_1702,N_1482);
or U2139 (N_2139,N_1112,N_1300);
and U2140 (N_2140,N_1040,N_1737);
or U2141 (N_2141,N_1027,N_1133);
and U2142 (N_2142,N_1945,N_1362);
nor U2143 (N_2143,N_1769,N_1522);
nor U2144 (N_2144,N_1047,N_1957);
nand U2145 (N_2145,N_1172,N_1944);
or U2146 (N_2146,N_1181,N_1002);
nor U2147 (N_2147,N_1703,N_1801);
nand U2148 (N_2148,N_1767,N_1069);
and U2149 (N_2149,N_1693,N_1488);
nand U2150 (N_2150,N_1342,N_1059);
nor U2151 (N_2151,N_1599,N_1352);
nor U2152 (N_2152,N_1914,N_1984);
nand U2153 (N_2153,N_1754,N_1209);
nand U2154 (N_2154,N_1838,N_1926);
nor U2155 (N_2155,N_1823,N_1267);
nand U2156 (N_2156,N_1810,N_1433);
nor U2157 (N_2157,N_1543,N_1755);
and U2158 (N_2158,N_1904,N_1152);
nor U2159 (N_2159,N_1654,N_1963);
or U2160 (N_2160,N_1605,N_1573);
nor U2161 (N_2161,N_1223,N_1902);
or U2162 (N_2162,N_1730,N_1529);
nor U2163 (N_2163,N_1624,N_1003);
nor U2164 (N_2164,N_1412,N_1313);
nand U2165 (N_2165,N_1322,N_1930);
and U2166 (N_2166,N_1111,N_1347);
or U2167 (N_2167,N_1105,N_1725);
or U2168 (N_2168,N_1746,N_1528);
nand U2169 (N_2169,N_1938,N_1418);
nand U2170 (N_2170,N_1587,N_1282);
and U2171 (N_2171,N_1420,N_1427);
nand U2172 (N_2172,N_1130,N_1743);
and U2173 (N_2173,N_1635,N_1723);
nor U2174 (N_2174,N_1000,N_1827);
nand U2175 (N_2175,N_1969,N_1815);
nor U2176 (N_2176,N_1596,N_1392);
or U2177 (N_2177,N_1614,N_1669);
nand U2178 (N_2178,N_1692,N_1554);
nand U2179 (N_2179,N_1515,N_1758);
or U2180 (N_2180,N_1764,N_1837);
nand U2181 (N_2181,N_1406,N_1314);
and U2182 (N_2182,N_1029,N_1650);
or U2183 (N_2183,N_1924,N_1996);
nand U2184 (N_2184,N_1713,N_1958);
nor U2185 (N_2185,N_1774,N_1364);
and U2186 (N_2186,N_1142,N_1558);
nand U2187 (N_2187,N_1961,N_1309);
and U2188 (N_2188,N_1446,N_1632);
or U2189 (N_2189,N_1789,N_1384);
nand U2190 (N_2190,N_1820,N_1119);
nor U2191 (N_2191,N_1765,N_1592);
or U2192 (N_2192,N_1155,N_1792);
or U2193 (N_2193,N_1892,N_1875);
nand U2194 (N_2194,N_1132,N_1491);
nor U2195 (N_2195,N_1162,N_1840);
or U2196 (N_2196,N_1539,N_1629);
or U2197 (N_2197,N_1665,N_1031);
and U2198 (N_2198,N_1992,N_1455);
or U2199 (N_2199,N_1965,N_1720);
or U2200 (N_2200,N_1115,N_1254);
nand U2201 (N_2201,N_1885,N_1582);
and U2202 (N_2202,N_1671,N_1019);
or U2203 (N_2203,N_1273,N_1325);
and U2204 (N_2204,N_1391,N_1630);
or U2205 (N_2205,N_1514,N_1266);
and U2206 (N_2206,N_1983,N_1575);
nand U2207 (N_2207,N_1247,N_1139);
and U2208 (N_2208,N_1008,N_1343);
and U2209 (N_2209,N_1143,N_1241);
nand U2210 (N_2210,N_1530,N_1525);
and U2211 (N_2211,N_1557,N_1410);
nand U2212 (N_2212,N_1717,N_1847);
or U2213 (N_2213,N_1679,N_1825);
or U2214 (N_2214,N_1292,N_1056);
or U2215 (N_2215,N_1872,N_1905);
nor U2216 (N_2216,N_1416,N_1659);
or U2217 (N_2217,N_1492,N_1020);
nor U2218 (N_2218,N_1380,N_1361);
nand U2219 (N_2219,N_1259,N_1320);
or U2220 (N_2220,N_1928,N_1450);
nor U2221 (N_2221,N_1461,N_1714);
nand U2222 (N_2222,N_1896,N_1805);
or U2223 (N_2223,N_1893,N_1240);
nand U2224 (N_2224,N_1277,N_1733);
and U2225 (N_2225,N_1519,N_1726);
nor U2226 (N_2226,N_1934,N_1877);
nor U2227 (N_2227,N_1030,N_1602);
nor U2228 (N_2228,N_1183,N_1971);
nor U2229 (N_2229,N_1091,N_1170);
nand U2230 (N_2230,N_1159,N_1371);
nand U2231 (N_2231,N_1552,N_1072);
or U2232 (N_2232,N_1771,N_1822);
nor U2233 (N_2233,N_1715,N_1462);
or U2234 (N_2234,N_1301,N_1264);
or U2235 (N_2235,N_1814,N_1791);
or U2236 (N_2236,N_1216,N_1817);
and U2237 (N_2237,N_1708,N_1234);
nor U2238 (N_2238,N_1326,N_1638);
nor U2239 (N_2239,N_1126,N_1150);
nand U2240 (N_2240,N_1718,N_1738);
and U2241 (N_2241,N_1188,N_1191);
or U2242 (N_2242,N_1289,N_1952);
nor U2243 (N_2243,N_1962,N_1581);
nand U2244 (N_2244,N_1262,N_1867);
nand U2245 (N_2245,N_1476,N_1051);
or U2246 (N_2246,N_1981,N_1200);
nor U2247 (N_2247,N_1735,N_1185);
or U2248 (N_2248,N_1206,N_1390);
and U2249 (N_2249,N_1832,N_1473);
or U2250 (N_2250,N_1444,N_1120);
xor U2251 (N_2251,N_1057,N_1727);
nand U2252 (N_2252,N_1751,N_1306);
and U2253 (N_2253,N_1454,N_1970);
or U2254 (N_2254,N_1106,N_1213);
nand U2255 (N_2255,N_1068,N_1796);
or U2256 (N_2256,N_1848,N_1423);
and U2257 (N_2257,N_1511,N_1459);
and U2258 (N_2258,N_1640,N_1580);
nand U2259 (N_2259,N_1415,N_1353);
or U2260 (N_2260,N_1261,N_1137);
or U2261 (N_2261,N_1011,N_1920);
nor U2262 (N_2262,N_1413,N_1836);
and U2263 (N_2263,N_1806,N_1442);
and U2264 (N_2264,N_1859,N_1218);
or U2265 (N_2265,N_1722,N_1616);
nand U2266 (N_2266,N_1481,N_1078);
or U2267 (N_2267,N_1631,N_1586);
nor U2268 (N_2268,N_1542,N_1647);
nand U2269 (N_2269,N_1683,N_1748);
or U2270 (N_2270,N_1363,N_1101);
nor U2271 (N_2271,N_1379,N_1919);
nor U2272 (N_2272,N_1090,N_1479);
nor U2273 (N_2273,N_1600,N_1565);
nor U2274 (N_2274,N_1465,N_1340);
nor U2275 (N_2275,N_1372,N_1285);
nand U2276 (N_2276,N_1657,N_1417);
nor U2277 (N_2277,N_1968,N_1470);
nand U2278 (N_2278,N_1192,N_1049);
nor U2279 (N_2279,N_1359,N_1006);
nand U2280 (N_2280,N_1131,N_1950);
or U2281 (N_2281,N_1332,N_1779);
nor U2282 (N_2282,N_1283,N_1044);
and U2283 (N_2283,N_1601,N_1982);
and U2284 (N_2284,N_1784,N_1927);
or U2285 (N_2285,N_1989,N_1103);
nor U2286 (N_2286,N_1256,N_1010);
or U2287 (N_2287,N_1463,N_1425);
or U2288 (N_2288,N_1639,N_1923);
and U2289 (N_2289,N_1055,N_1158);
nand U2290 (N_2290,N_1595,N_1305);
nor U2291 (N_2291,N_1366,N_1917);
or U2292 (N_2292,N_1288,N_1251);
or U2293 (N_2293,N_1574,N_1878);
and U2294 (N_2294,N_1861,N_1620);
or U2295 (N_2295,N_1585,N_1012);
or U2296 (N_2296,N_1333,N_1365);
or U2297 (N_2297,N_1205,N_1327);
nand U2298 (N_2298,N_1217,N_1852);
or U2299 (N_2299,N_1272,N_1860);
and U2300 (N_2300,N_1697,N_1674);
and U2301 (N_2301,N_1918,N_1096);
or U2302 (N_2302,N_1922,N_1943);
nand U2303 (N_2303,N_1428,N_1134);
and U2304 (N_2304,N_1439,N_1348);
and U2305 (N_2305,N_1187,N_1869);
and U2306 (N_2306,N_1260,N_1626);
and U2307 (N_2307,N_1176,N_1250);
nand U2308 (N_2308,N_1537,N_1258);
nand U2309 (N_2309,N_1411,N_1471);
or U2310 (N_2310,N_1531,N_1547);
or U2311 (N_2311,N_1731,N_1496);
nor U2312 (N_2312,N_1584,N_1881);
or U2313 (N_2313,N_1407,N_1513);
nand U2314 (N_2314,N_1682,N_1839);
and U2315 (N_2315,N_1524,N_1394);
xnor U2316 (N_2316,N_1445,N_1041);
and U2317 (N_2317,N_1037,N_1422);
and U2318 (N_2318,N_1821,N_1375);
and U2319 (N_2319,N_1053,N_1426);
or U2320 (N_2320,N_1207,N_1244);
and U2321 (N_2321,N_1870,N_1498);
nor U2322 (N_2322,N_1432,N_1075);
nand U2323 (N_2323,N_1179,N_1178);
or U2324 (N_2324,N_1523,N_1497);
or U2325 (N_2325,N_1705,N_1253);
and U2326 (N_2326,N_1494,N_1541);
nand U2327 (N_2327,N_1229,N_1360);
or U2328 (N_2328,N_1741,N_1299);
and U2329 (N_2329,N_1368,N_1232);
and U2330 (N_2330,N_1698,N_1138);
nand U2331 (N_2331,N_1701,N_1453);
or U2332 (N_2332,N_1874,N_1967);
nor U2333 (N_2333,N_1356,N_1576);
or U2334 (N_2334,N_1163,N_1564);
nand U2335 (N_2335,N_1911,N_1648);
and U2336 (N_2336,N_1673,N_1503);
nand U2337 (N_2337,N_1156,N_1653);
nor U2338 (N_2338,N_1016,N_1116);
and U2339 (N_2339,N_1546,N_1071);
nand U2340 (N_2340,N_1811,N_1166);
or U2341 (N_2341,N_1182,N_1518);
xnor U2342 (N_2342,N_1894,N_1670);
nand U2343 (N_2343,N_1710,N_1310);
nand U2344 (N_2344,N_1193,N_1129);
and U2345 (N_2345,N_1808,N_1807);
nor U2346 (N_2346,N_1469,N_1061);
nor U2347 (N_2347,N_1393,N_1121);
nor U2348 (N_2348,N_1215,N_1381);
nor U2349 (N_2349,N_1964,N_1550);
or U2350 (N_2350,N_1175,N_1641);
nor U2351 (N_2351,N_1328,N_1123);
or U2352 (N_2352,N_1233,N_1263);
nand U2353 (N_2353,N_1972,N_1265);
nor U2354 (N_2354,N_1023,N_1985);
nand U2355 (N_2355,N_1278,N_1772);
or U2356 (N_2356,N_1858,N_1414);
nand U2357 (N_2357,N_1274,N_1054);
or U2358 (N_2358,N_1436,N_1721);
nor U2359 (N_2359,N_1430,N_1369);
nand U2360 (N_2360,N_1219,N_1144);
or U2361 (N_2361,N_1434,N_1148);
and U2362 (N_2362,N_1404,N_1687);
or U2363 (N_2363,N_1504,N_1082);
nor U2364 (N_2364,N_1695,N_1949);
and U2365 (N_2365,N_1512,N_1312);
nand U2366 (N_2366,N_1835,N_1464);
nand U2367 (N_2367,N_1290,N_1855);
and U2368 (N_2368,N_1490,N_1897);
and U2369 (N_2369,N_1609,N_1658);
nor U2370 (N_2370,N_1063,N_1398);
nand U2371 (N_2371,N_1097,N_1728);
nand U2372 (N_2372,N_1770,N_1311);
nor U2373 (N_2373,N_1475,N_1141);
or U2374 (N_2374,N_1561,N_1316);
and U2375 (N_2375,N_1903,N_1401);
or U2376 (N_2376,N_1321,N_1220);
and U2377 (N_2377,N_1028,N_1776);
and U2378 (N_2378,N_1644,N_1997);
nor U2379 (N_2379,N_1622,N_1979);
or U2380 (N_2380,N_1555,N_1763);
and U2381 (N_2381,N_1857,N_1409);
xor U2382 (N_2382,N_1066,N_1991);
or U2383 (N_2383,N_1994,N_1070);
nand U2384 (N_2384,N_1851,N_1211);
and U2385 (N_2385,N_1976,N_1951);
nand U2386 (N_2386,N_1237,N_1834);
or U2387 (N_2387,N_1245,N_1396);
nor U2388 (N_2388,N_1035,N_1975);
nor U2389 (N_2389,N_1830,N_1388);
or U2390 (N_2390,N_1231,N_1729);
nand U2391 (N_2391,N_1201,N_1165);
and U2392 (N_2392,N_1803,N_1024);
and U2393 (N_2393,N_1015,N_1781);
and U2394 (N_2394,N_1910,N_1637);
nor U2395 (N_2395,N_1933,N_1612);
and U2396 (N_2396,N_1243,N_1590);
or U2397 (N_2397,N_1946,N_1382);
or U2398 (N_2398,N_1898,N_1802);
and U2399 (N_2399,N_1114,N_1048);
or U2400 (N_2400,N_1932,N_1895);
and U2401 (N_2401,N_1225,N_1092);
nand U2402 (N_2402,N_1287,N_1716);
nor U2403 (N_2403,N_1110,N_1295);
or U2404 (N_2404,N_1064,N_1925);
nor U2405 (N_2405,N_1813,N_1597);
nand U2406 (N_2406,N_1873,N_1408);
nor U2407 (N_2407,N_1775,N_1974);
or U2408 (N_2408,N_1824,N_1378);
or U2409 (N_2409,N_1535,N_1980);
and U2410 (N_2410,N_1740,N_1060);
nand U2411 (N_2411,N_1466,N_1468);
nand U2412 (N_2412,N_1826,N_1081);
and U2413 (N_2413,N_1572,N_1790);
nor U2414 (N_2414,N_1113,N_1882);
or U2415 (N_2415,N_1691,N_1621);
and U2416 (N_2416,N_1615,N_1358);
nor U2417 (N_2417,N_1732,N_1424);
or U2418 (N_2418,N_1303,N_1457);
and U2419 (N_2419,N_1651,N_1050);
or U2420 (N_2420,N_1625,N_1094);
or U2421 (N_2421,N_1025,N_1108);
or U2422 (N_2422,N_1966,N_1026);
nand U2423 (N_2423,N_1135,N_1186);
nor U2424 (N_2424,N_1440,N_1777);
or U2425 (N_2425,N_1734,N_1255);
and U2426 (N_2426,N_1102,N_1603);
or U2427 (N_2427,N_1018,N_1324);
nor U2428 (N_2428,N_1077,N_1293);
nor U2429 (N_2429,N_1990,N_1341);
or U2430 (N_2430,N_1350,N_1189);
or U2431 (N_2431,N_1880,N_1443);
nand U2432 (N_2432,N_1073,N_1485);
nand U2433 (N_2433,N_1323,N_1560);
and U2434 (N_2434,N_1437,N_1617);
nor U2435 (N_2435,N_1286,N_1661);
or U2436 (N_2436,N_1948,N_1238);
or U2437 (N_2437,N_1367,N_1451);
nand U2438 (N_2438,N_1095,N_1400);
nand U2439 (N_2439,N_1913,N_1907);
nor U2440 (N_2440,N_1085,N_1249);
nor U2441 (N_2441,N_1536,N_1804);
nand U2442 (N_2442,N_1038,N_1067);
nor U2443 (N_2443,N_1315,N_1956);
or U2444 (N_2444,N_1786,N_1164);
nand U2445 (N_2445,N_1395,N_1004);
nand U2446 (N_2446,N_1579,N_1694);
or U2447 (N_2447,N_1864,N_1345);
nand U2448 (N_2448,N_1149,N_1246);
nor U2449 (N_2449,N_1888,N_1100);
and U2450 (N_2450,N_1570,N_1749);
nor U2451 (N_2451,N_1959,N_1435);
nand U2452 (N_2452,N_1652,N_1088);
and U2453 (N_2453,N_1793,N_1977);
and U2454 (N_2454,N_1854,N_1563);
or U2455 (N_2455,N_1083,N_1696);
and U2456 (N_2456,N_1853,N_1147);
nor U2457 (N_2457,N_1089,N_1001);
nand U2458 (N_2458,N_1761,N_1279);
or U2459 (N_2459,N_1680,N_1501);
nor U2460 (N_2460,N_1157,N_1797);
nor U2461 (N_2461,N_1672,N_1502);
nor U2462 (N_2462,N_1676,N_1699);
nor U2463 (N_2463,N_1467,N_1756);
nand U2464 (N_2464,N_1294,N_1677);
or U2465 (N_2465,N_1593,N_1065);
and U2466 (N_2466,N_1828,N_1995);
nand U2467 (N_2467,N_1642,N_1268);
nor U2468 (N_2468,N_1210,N_1174);
nand U2469 (N_2469,N_1551,N_1700);
or U2470 (N_2470,N_1487,N_1634);
or U2471 (N_2471,N_1212,N_1667);
nor U2472 (N_2472,N_1533,N_1594);
nand U2473 (N_2473,N_1124,N_1850);
and U2474 (N_2474,N_1656,N_1036);
nor U2475 (N_2475,N_1901,N_1252);
or U2476 (N_2476,N_1711,N_1140);
nand U2477 (N_2477,N_1195,N_1196);
nand U2478 (N_2478,N_1795,N_1690);
and U2479 (N_2479,N_1448,N_1224);
nand U2480 (N_2480,N_1074,N_1161);
nand U2481 (N_2481,N_1941,N_1818);
and U2482 (N_2482,N_1099,N_1921);
nand U2483 (N_2483,N_1429,N_1098);
or U2484 (N_2484,N_1042,N_1611);
nor U2485 (N_2485,N_1499,N_1794);
nor U2486 (N_2486,N_1591,N_1577);
and U2487 (N_2487,N_1403,N_1483);
nand U2488 (N_2488,N_1284,N_1788);
nand U2489 (N_2489,N_1899,N_1668);
or U2490 (N_2490,N_1973,N_1684);
nand U2491 (N_2491,N_1039,N_1107);
nor U2492 (N_2492,N_1712,N_1506);
or U2493 (N_2493,N_1194,N_1160);
or U2494 (N_2494,N_1460,N_1509);
or U2495 (N_2495,N_1230,N_1890);
or U2496 (N_2496,N_1402,N_1646);
nor U2497 (N_2497,N_1242,N_1474);
and U2498 (N_2498,N_1197,N_1685);
and U2499 (N_2499,N_1171,N_1736);
or U2500 (N_2500,N_1245,N_1949);
nor U2501 (N_2501,N_1664,N_1090);
nand U2502 (N_2502,N_1094,N_1255);
nor U2503 (N_2503,N_1444,N_1634);
nor U2504 (N_2504,N_1181,N_1518);
nand U2505 (N_2505,N_1184,N_1706);
nor U2506 (N_2506,N_1728,N_1133);
and U2507 (N_2507,N_1507,N_1927);
and U2508 (N_2508,N_1125,N_1887);
and U2509 (N_2509,N_1442,N_1760);
nand U2510 (N_2510,N_1824,N_1558);
nor U2511 (N_2511,N_1149,N_1638);
nor U2512 (N_2512,N_1956,N_1162);
nor U2513 (N_2513,N_1324,N_1040);
or U2514 (N_2514,N_1949,N_1430);
nand U2515 (N_2515,N_1675,N_1215);
and U2516 (N_2516,N_1174,N_1536);
nand U2517 (N_2517,N_1985,N_1641);
and U2518 (N_2518,N_1187,N_1590);
or U2519 (N_2519,N_1156,N_1392);
or U2520 (N_2520,N_1857,N_1954);
and U2521 (N_2521,N_1170,N_1015);
nor U2522 (N_2522,N_1348,N_1835);
or U2523 (N_2523,N_1070,N_1291);
and U2524 (N_2524,N_1648,N_1012);
nand U2525 (N_2525,N_1247,N_1417);
nor U2526 (N_2526,N_1283,N_1747);
or U2527 (N_2527,N_1975,N_1294);
nor U2528 (N_2528,N_1157,N_1953);
or U2529 (N_2529,N_1826,N_1214);
nand U2530 (N_2530,N_1336,N_1386);
and U2531 (N_2531,N_1963,N_1437);
or U2532 (N_2532,N_1464,N_1920);
nand U2533 (N_2533,N_1560,N_1848);
nand U2534 (N_2534,N_1351,N_1790);
nor U2535 (N_2535,N_1636,N_1698);
nand U2536 (N_2536,N_1838,N_1278);
nand U2537 (N_2537,N_1759,N_1805);
nor U2538 (N_2538,N_1324,N_1170);
and U2539 (N_2539,N_1892,N_1409);
nand U2540 (N_2540,N_1680,N_1126);
or U2541 (N_2541,N_1681,N_1958);
nor U2542 (N_2542,N_1953,N_1450);
or U2543 (N_2543,N_1886,N_1233);
or U2544 (N_2544,N_1012,N_1526);
or U2545 (N_2545,N_1736,N_1342);
nand U2546 (N_2546,N_1657,N_1444);
nor U2547 (N_2547,N_1985,N_1983);
nor U2548 (N_2548,N_1303,N_1895);
or U2549 (N_2549,N_1549,N_1312);
and U2550 (N_2550,N_1006,N_1094);
nor U2551 (N_2551,N_1644,N_1170);
nand U2552 (N_2552,N_1462,N_1428);
nor U2553 (N_2553,N_1881,N_1438);
nand U2554 (N_2554,N_1957,N_1763);
nor U2555 (N_2555,N_1047,N_1361);
or U2556 (N_2556,N_1947,N_1112);
nor U2557 (N_2557,N_1976,N_1187);
nand U2558 (N_2558,N_1837,N_1112);
and U2559 (N_2559,N_1587,N_1817);
and U2560 (N_2560,N_1160,N_1365);
nand U2561 (N_2561,N_1885,N_1381);
nor U2562 (N_2562,N_1804,N_1802);
nor U2563 (N_2563,N_1526,N_1889);
nor U2564 (N_2564,N_1890,N_1015);
and U2565 (N_2565,N_1731,N_1587);
nor U2566 (N_2566,N_1426,N_1989);
nor U2567 (N_2567,N_1908,N_1070);
nand U2568 (N_2568,N_1131,N_1457);
nand U2569 (N_2569,N_1120,N_1725);
and U2570 (N_2570,N_1150,N_1121);
or U2571 (N_2571,N_1808,N_1364);
nor U2572 (N_2572,N_1706,N_1077);
and U2573 (N_2573,N_1893,N_1833);
nor U2574 (N_2574,N_1695,N_1251);
or U2575 (N_2575,N_1048,N_1544);
nand U2576 (N_2576,N_1840,N_1760);
or U2577 (N_2577,N_1694,N_1219);
nor U2578 (N_2578,N_1407,N_1473);
nand U2579 (N_2579,N_1597,N_1334);
and U2580 (N_2580,N_1078,N_1069);
and U2581 (N_2581,N_1100,N_1050);
nor U2582 (N_2582,N_1307,N_1441);
nor U2583 (N_2583,N_1509,N_1040);
or U2584 (N_2584,N_1722,N_1036);
nor U2585 (N_2585,N_1723,N_1890);
nor U2586 (N_2586,N_1633,N_1900);
nor U2587 (N_2587,N_1268,N_1953);
nor U2588 (N_2588,N_1269,N_1878);
nor U2589 (N_2589,N_1891,N_1436);
and U2590 (N_2590,N_1739,N_1160);
nor U2591 (N_2591,N_1033,N_1537);
nand U2592 (N_2592,N_1098,N_1373);
or U2593 (N_2593,N_1137,N_1455);
or U2594 (N_2594,N_1826,N_1201);
nor U2595 (N_2595,N_1055,N_1361);
and U2596 (N_2596,N_1169,N_1480);
or U2597 (N_2597,N_1730,N_1026);
nand U2598 (N_2598,N_1320,N_1079);
nand U2599 (N_2599,N_1591,N_1567);
nand U2600 (N_2600,N_1810,N_1466);
and U2601 (N_2601,N_1774,N_1662);
nor U2602 (N_2602,N_1042,N_1875);
xor U2603 (N_2603,N_1273,N_1164);
nor U2604 (N_2604,N_1631,N_1095);
nor U2605 (N_2605,N_1481,N_1816);
or U2606 (N_2606,N_1508,N_1461);
nor U2607 (N_2607,N_1946,N_1576);
nor U2608 (N_2608,N_1299,N_1311);
and U2609 (N_2609,N_1566,N_1222);
nand U2610 (N_2610,N_1072,N_1361);
or U2611 (N_2611,N_1568,N_1416);
or U2612 (N_2612,N_1014,N_1921);
or U2613 (N_2613,N_1444,N_1320);
nor U2614 (N_2614,N_1554,N_1543);
or U2615 (N_2615,N_1176,N_1487);
or U2616 (N_2616,N_1396,N_1829);
and U2617 (N_2617,N_1462,N_1432);
nor U2618 (N_2618,N_1213,N_1569);
and U2619 (N_2619,N_1495,N_1450);
and U2620 (N_2620,N_1732,N_1043);
nand U2621 (N_2621,N_1930,N_1560);
or U2622 (N_2622,N_1794,N_1438);
nand U2623 (N_2623,N_1544,N_1956);
nor U2624 (N_2624,N_1454,N_1220);
nor U2625 (N_2625,N_1537,N_1346);
nand U2626 (N_2626,N_1686,N_1865);
and U2627 (N_2627,N_1259,N_1978);
and U2628 (N_2628,N_1980,N_1445);
nor U2629 (N_2629,N_1392,N_1039);
xor U2630 (N_2630,N_1993,N_1179);
nor U2631 (N_2631,N_1708,N_1204);
xor U2632 (N_2632,N_1703,N_1097);
and U2633 (N_2633,N_1770,N_1404);
nor U2634 (N_2634,N_1869,N_1785);
and U2635 (N_2635,N_1430,N_1317);
or U2636 (N_2636,N_1873,N_1778);
nor U2637 (N_2637,N_1632,N_1831);
and U2638 (N_2638,N_1171,N_1454);
and U2639 (N_2639,N_1485,N_1557);
or U2640 (N_2640,N_1047,N_1683);
or U2641 (N_2641,N_1565,N_1299);
nor U2642 (N_2642,N_1093,N_1657);
or U2643 (N_2643,N_1034,N_1015);
nand U2644 (N_2644,N_1621,N_1807);
nor U2645 (N_2645,N_1264,N_1747);
nor U2646 (N_2646,N_1566,N_1923);
nor U2647 (N_2647,N_1684,N_1220);
nor U2648 (N_2648,N_1251,N_1028);
nand U2649 (N_2649,N_1019,N_1063);
nor U2650 (N_2650,N_1643,N_1185);
or U2651 (N_2651,N_1565,N_1903);
nor U2652 (N_2652,N_1516,N_1672);
nand U2653 (N_2653,N_1200,N_1767);
nor U2654 (N_2654,N_1873,N_1797);
nor U2655 (N_2655,N_1034,N_1356);
nand U2656 (N_2656,N_1985,N_1459);
nor U2657 (N_2657,N_1318,N_1540);
nor U2658 (N_2658,N_1696,N_1114);
nand U2659 (N_2659,N_1515,N_1825);
and U2660 (N_2660,N_1939,N_1958);
nand U2661 (N_2661,N_1138,N_1125);
nand U2662 (N_2662,N_1964,N_1759);
or U2663 (N_2663,N_1098,N_1503);
nand U2664 (N_2664,N_1016,N_1488);
or U2665 (N_2665,N_1861,N_1426);
and U2666 (N_2666,N_1208,N_1408);
and U2667 (N_2667,N_1261,N_1028);
and U2668 (N_2668,N_1702,N_1807);
or U2669 (N_2669,N_1125,N_1290);
and U2670 (N_2670,N_1342,N_1836);
and U2671 (N_2671,N_1930,N_1667);
and U2672 (N_2672,N_1647,N_1792);
nor U2673 (N_2673,N_1443,N_1625);
and U2674 (N_2674,N_1416,N_1363);
and U2675 (N_2675,N_1573,N_1300);
nor U2676 (N_2676,N_1721,N_1550);
or U2677 (N_2677,N_1598,N_1603);
and U2678 (N_2678,N_1358,N_1853);
nand U2679 (N_2679,N_1734,N_1854);
nor U2680 (N_2680,N_1460,N_1145);
or U2681 (N_2681,N_1728,N_1575);
or U2682 (N_2682,N_1176,N_1665);
and U2683 (N_2683,N_1007,N_1750);
or U2684 (N_2684,N_1133,N_1316);
or U2685 (N_2685,N_1444,N_1829);
nor U2686 (N_2686,N_1467,N_1361);
nor U2687 (N_2687,N_1145,N_1961);
and U2688 (N_2688,N_1962,N_1242);
or U2689 (N_2689,N_1533,N_1970);
and U2690 (N_2690,N_1447,N_1418);
and U2691 (N_2691,N_1224,N_1532);
or U2692 (N_2692,N_1008,N_1869);
and U2693 (N_2693,N_1304,N_1958);
nand U2694 (N_2694,N_1722,N_1494);
nor U2695 (N_2695,N_1563,N_1931);
nand U2696 (N_2696,N_1102,N_1414);
nor U2697 (N_2697,N_1818,N_1075);
and U2698 (N_2698,N_1457,N_1235);
and U2699 (N_2699,N_1346,N_1194);
and U2700 (N_2700,N_1633,N_1138);
and U2701 (N_2701,N_1511,N_1807);
and U2702 (N_2702,N_1076,N_1248);
and U2703 (N_2703,N_1297,N_1027);
nand U2704 (N_2704,N_1813,N_1935);
or U2705 (N_2705,N_1321,N_1489);
nor U2706 (N_2706,N_1672,N_1805);
nand U2707 (N_2707,N_1970,N_1043);
and U2708 (N_2708,N_1905,N_1654);
nand U2709 (N_2709,N_1730,N_1472);
and U2710 (N_2710,N_1562,N_1720);
nor U2711 (N_2711,N_1908,N_1867);
or U2712 (N_2712,N_1660,N_1696);
and U2713 (N_2713,N_1171,N_1119);
nand U2714 (N_2714,N_1856,N_1213);
or U2715 (N_2715,N_1149,N_1258);
or U2716 (N_2716,N_1536,N_1596);
and U2717 (N_2717,N_1564,N_1832);
nor U2718 (N_2718,N_1474,N_1637);
or U2719 (N_2719,N_1470,N_1598);
or U2720 (N_2720,N_1574,N_1409);
or U2721 (N_2721,N_1800,N_1901);
nand U2722 (N_2722,N_1518,N_1813);
nor U2723 (N_2723,N_1488,N_1369);
or U2724 (N_2724,N_1740,N_1370);
nor U2725 (N_2725,N_1299,N_1796);
and U2726 (N_2726,N_1937,N_1724);
and U2727 (N_2727,N_1898,N_1611);
nand U2728 (N_2728,N_1509,N_1518);
and U2729 (N_2729,N_1845,N_1672);
or U2730 (N_2730,N_1712,N_1711);
or U2731 (N_2731,N_1101,N_1602);
and U2732 (N_2732,N_1897,N_1327);
or U2733 (N_2733,N_1839,N_1930);
nor U2734 (N_2734,N_1208,N_1893);
or U2735 (N_2735,N_1473,N_1260);
nor U2736 (N_2736,N_1872,N_1248);
nand U2737 (N_2737,N_1571,N_1788);
nor U2738 (N_2738,N_1947,N_1314);
or U2739 (N_2739,N_1243,N_1250);
nor U2740 (N_2740,N_1595,N_1674);
or U2741 (N_2741,N_1097,N_1699);
and U2742 (N_2742,N_1347,N_1682);
nand U2743 (N_2743,N_1595,N_1250);
nand U2744 (N_2744,N_1541,N_1484);
nand U2745 (N_2745,N_1662,N_1532);
nor U2746 (N_2746,N_1160,N_1582);
nor U2747 (N_2747,N_1553,N_1498);
or U2748 (N_2748,N_1026,N_1448);
and U2749 (N_2749,N_1473,N_1507);
or U2750 (N_2750,N_1323,N_1346);
or U2751 (N_2751,N_1589,N_1734);
and U2752 (N_2752,N_1847,N_1070);
nor U2753 (N_2753,N_1426,N_1681);
nand U2754 (N_2754,N_1062,N_1178);
nor U2755 (N_2755,N_1610,N_1353);
nor U2756 (N_2756,N_1777,N_1876);
and U2757 (N_2757,N_1990,N_1815);
nor U2758 (N_2758,N_1880,N_1335);
and U2759 (N_2759,N_1098,N_1260);
and U2760 (N_2760,N_1854,N_1830);
nor U2761 (N_2761,N_1628,N_1253);
nand U2762 (N_2762,N_1579,N_1409);
nand U2763 (N_2763,N_1807,N_1972);
and U2764 (N_2764,N_1599,N_1143);
xor U2765 (N_2765,N_1492,N_1332);
or U2766 (N_2766,N_1053,N_1273);
nor U2767 (N_2767,N_1604,N_1547);
or U2768 (N_2768,N_1072,N_1283);
or U2769 (N_2769,N_1113,N_1599);
and U2770 (N_2770,N_1257,N_1256);
nor U2771 (N_2771,N_1645,N_1017);
or U2772 (N_2772,N_1669,N_1968);
nor U2773 (N_2773,N_1164,N_1704);
nand U2774 (N_2774,N_1186,N_1582);
and U2775 (N_2775,N_1289,N_1818);
and U2776 (N_2776,N_1172,N_1435);
nand U2777 (N_2777,N_1854,N_1412);
or U2778 (N_2778,N_1724,N_1267);
nor U2779 (N_2779,N_1104,N_1343);
nor U2780 (N_2780,N_1860,N_1545);
nand U2781 (N_2781,N_1932,N_1199);
or U2782 (N_2782,N_1777,N_1393);
or U2783 (N_2783,N_1602,N_1140);
nor U2784 (N_2784,N_1875,N_1919);
or U2785 (N_2785,N_1976,N_1597);
and U2786 (N_2786,N_1936,N_1239);
and U2787 (N_2787,N_1296,N_1390);
and U2788 (N_2788,N_1020,N_1386);
or U2789 (N_2789,N_1199,N_1692);
or U2790 (N_2790,N_1476,N_1335);
xor U2791 (N_2791,N_1124,N_1546);
and U2792 (N_2792,N_1336,N_1120);
or U2793 (N_2793,N_1319,N_1649);
and U2794 (N_2794,N_1204,N_1422);
nand U2795 (N_2795,N_1612,N_1788);
and U2796 (N_2796,N_1027,N_1643);
nor U2797 (N_2797,N_1298,N_1592);
and U2798 (N_2798,N_1705,N_1130);
or U2799 (N_2799,N_1005,N_1198);
nor U2800 (N_2800,N_1480,N_1580);
and U2801 (N_2801,N_1498,N_1631);
nor U2802 (N_2802,N_1426,N_1012);
nor U2803 (N_2803,N_1754,N_1025);
nor U2804 (N_2804,N_1644,N_1917);
nand U2805 (N_2805,N_1961,N_1627);
nor U2806 (N_2806,N_1704,N_1465);
nand U2807 (N_2807,N_1527,N_1977);
xnor U2808 (N_2808,N_1922,N_1041);
nor U2809 (N_2809,N_1332,N_1705);
and U2810 (N_2810,N_1535,N_1778);
nand U2811 (N_2811,N_1610,N_1598);
nand U2812 (N_2812,N_1810,N_1851);
nor U2813 (N_2813,N_1823,N_1634);
xor U2814 (N_2814,N_1937,N_1309);
and U2815 (N_2815,N_1168,N_1982);
nand U2816 (N_2816,N_1863,N_1038);
nand U2817 (N_2817,N_1056,N_1646);
and U2818 (N_2818,N_1046,N_1338);
or U2819 (N_2819,N_1790,N_1650);
or U2820 (N_2820,N_1892,N_1001);
nand U2821 (N_2821,N_1975,N_1047);
nand U2822 (N_2822,N_1719,N_1358);
nor U2823 (N_2823,N_1792,N_1967);
nor U2824 (N_2824,N_1639,N_1720);
nand U2825 (N_2825,N_1951,N_1855);
nand U2826 (N_2826,N_1698,N_1198);
nor U2827 (N_2827,N_1619,N_1038);
and U2828 (N_2828,N_1611,N_1286);
or U2829 (N_2829,N_1788,N_1734);
nand U2830 (N_2830,N_1921,N_1361);
and U2831 (N_2831,N_1597,N_1219);
and U2832 (N_2832,N_1951,N_1540);
or U2833 (N_2833,N_1760,N_1653);
nand U2834 (N_2834,N_1797,N_1755);
or U2835 (N_2835,N_1539,N_1006);
or U2836 (N_2836,N_1157,N_1035);
nor U2837 (N_2837,N_1232,N_1065);
nor U2838 (N_2838,N_1587,N_1781);
nor U2839 (N_2839,N_1242,N_1466);
nor U2840 (N_2840,N_1153,N_1180);
nor U2841 (N_2841,N_1241,N_1273);
and U2842 (N_2842,N_1435,N_1883);
or U2843 (N_2843,N_1501,N_1167);
and U2844 (N_2844,N_1041,N_1868);
nor U2845 (N_2845,N_1495,N_1153);
nor U2846 (N_2846,N_1598,N_1183);
and U2847 (N_2847,N_1297,N_1523);
or U2848 (N_2848,N_1369,N_1462);
nor U2849 (N_2849,N_1993,N_1650);
or U2850 (N_2850,N_1398,N_1761);
and U2851 (N_2851,N_1589,N_1717);
nand U2852 (N_2852,N_1557,N_1527);
and U2853 (N_2853,N_1885,N_1177);
and U2854 (N_2854,N_1342,N_1863);
nor U2855 (N_2855,N_1577,N_1568);
nor U2856 (N_2856,N_1972,N_1173);
nand U2857 (N_2857,N_1529,N_1657);
or U2858 (N_2858,N_1870,N_1212);
nand U2859 (N_2859,N_1549,N_1643);
nor U2860 (N_2860,N_1785,N_1377);
nand U2861 (N_2861,N_1494,N_1585);
and U2862 (N_2862,N_1202,N_1527);
nor U2863 (N_2863,N_1602,N_1115);
nand U2864 (N_2864,N_1137,N_1347);
nand U2865 (N_2865,N_1434,N_1259);
nand U2866 (N_2866,N_1327,N_1794);
and U2867 (N_2867,N_1658,N_1655);
or U2868 (N_2868,N_1491,N_1412);
xnor U2869 (N_2869,N_1147,N_1513);
nand U2870 (N_2870,N_1789,N_1562);
nor U2871 (N_2871,N_1186,N_1534);
nand U2872 (N_2872,N_1746,N_1749);
or U2873 (N_2873,N_1354,N_1916);
nor U2874 (N_2874,N_1610,N_1330);
nand U2875 (N_2875,N_1606,N_1465);
and U2876 (N_2876,N_1638,N_1097);
nor U2877 (N_2877,N_1122,N_1616);
and U2878 (N_2878,N_1779,N_1747);
nor U2879 (N_2879,N_1259,N_1449);
nand U2880 (N_2880,N_1904,N_1411);
or U2881 (N_2881,N_1721,N_1183);
nand U2882 (N_2882,N_1658,N_1718);
nand U2883 (N_2883,N_1319,N_1275);
nor U2884 (N_2884,N_1183,N_1570);
nor U2885 (N_2885,N_1274,N_1787);
nand U2886 (N_2886,N_1801,N_1743);
and U2887 (N_2887,N_1740,N_1793);
or U2888 (N_2888,N_1923,N_1622);
nand U2889 (N_2889,N_1712,N_1062);
nor U2890 (N_2890,N_1059,N_1282);
nand U2891 (N_2891,N_1377,N_1667);
nand U2892 (N_2892,N_1861,N_1450);
nor U2893 (N_2893,N_1640,N_1123);
or U2894 (N_2894,N_1799,N_1643);
and U2895 (N_2895,N_1701,N_1646);
and U2896 (N_2896,N_1731,N_1655);
or U2897 (N_2897,N_1011,N_1299);
nor U2898 (N_2898,N_1446,N_1545);
or U2899 (N_2899,N_1605,N_1518);
nor U2900 (N_2900,N_1609,N_1817);
and U2901 (N_2901,N_1299,N_1014);
nand U2902 (N_2902,N_1436,N_1967);
and U2903 (N_2903,N_1248,N_1056);
and U2904 (N_2904,N_1786,N_1494);
and U2905 (N_2905,N_1932,N_1344);
nand U2906 (N_2906,N_1894,N_1822);
nand U2907 (N_2907,N_1362,N_1408);
and U2908 (N_2908,N_1255,N_1469);
nor U2909 (N_2909,N_1626,N_1853);
nor U2910 (N_2910,N_1111,N_1840);
and U2911 (N_2911,N_1971,N_1017);
or U2912 (N_2912,N_1798,N_1752);
nand U2913 (N_2913,N_1608,N_1580);
or U2914 (N_2914,N_1219,N_1099);
or U2915 (N_2915,N_1536,N_1034);
nand U2916 (N_2916,N_1530,N_1237);
nor U2917 (N_2917,N_1440,N_1802);
or U2918 (N_2918,N_1468,N_1458);
nor U2919 (N_2919,N_1602,N_1878);
nand U2920 (N_2920,N_1079,N_1878);
or U2921 (N_2921,N_1923,N_1285);
nor U2922 (N_2922,N_1571,N_1441);
and U2923 (N_2923,N_1117,N_1975);
nor U2924 (N_2924,N_1030,N_1493);
and U2925 (N_2925,N_1047,N_1552);
nand U2926 (N_2926,N_1864,N_1808);
nand U2927 (N_2927,N_1699,N_1264);
nor U2928 (N_2928,N_1590,N_1792);
nor U2929 (N_2929,N_1032,N_1303);
nand U2930 (N_2930,N_1972,N_1356);
or U2931 (N_2931,N_1496,N_1841);
or U2932 (N_2932,N_1826,N_1371);
and U2933 (N_2933,N_1773,N_1337);
or U2934 (N_2934,N_1956,N_1275);
nand U2935 (N_2935,N_1112,N_1516);
nor U2936 (N_2936,N_1252,N_1735);
nand U2937 (N_2937,N_1583,N_1104);
and U2938 (N_2938,N_1155,N_1591);
nand U2939 (N_2939,N_1546,N_1932);
or U2940 (N_2940,N_1428,N_1592);
nor U2941 (N_2941,N_1853,N_1878);
and U2942 (N_2942,N_1081,N_1839);
and U2943 (N_2943,N_1178,N_1803);
or U2944 (N_2944,N_1803,N_1374);
and U2945 (N_2945,N_1807,N_1697);
and U2946 (N_2946,N_1905,N_1912);
and U2947 (N_2947,N_1074,N_1582);
nand U2948 (N_2948,N_1365,N_1334);
or U2949 (N_2949,N_1813,N_1835);
and U2950 (N_2950,N_1184,N_1110);
nor U2951 (N_2951,N_1054,N_1076);
or U2952 (N_2952,N_1167,N_1962);
or U2953 (N_2953,N_1585,N_1258);
and U2954 (N_2954,N_1097,N_1825);
and U2955 (N_2955,N_1771,N_1372);
nor U2956 (N_2956,N_1732,N_1252);
or U2957 (N_2957,N_1452,N_1455);
nor U2958 (N_2958,N_1687,N_1507);
nand U2959 (N_2959,N_1016,N_1551);
nand U2960 (N_2960,N_1214,N_1718);
nand U2961 (N_2961,N_1233,N_1224);
or U2962 (N_2962,N_1208,N_1744);
nand U2963 (N_2963,N_1862,N_1318);
and U2964 (N_2964,N_1384,N_1717);
nor U2965 (N_2965,N_1151,N_1312);
or U2966 (N_2966,N_1454,N_1531);
nand U2967 (N_2967,N_1379,N_1456);
nand U2968 (N_2968,N_1812,N_1374);
and U2969 (N_2969,N_1047,N_1011);
nand U2970 (N_2970,N_1214,N_1668);
and U2971 (N_2971,N_1645,N_1824);
and U2972 (N_2972,N_1343,N_1005);
nor U2973 (N_2973,N_1189,N_1162);
or U2974 (N_2974,N_1478,N_1508);
nand U2975 (N_2975,N_1293,N_1781);
nor U2976 (N_2976,N_1547,N_1432);
nor U2977 (N_2977,N_1142,N_1243);
nand U2978 (N_2978,N_1835,N_1139);
nor U2979 (N_2979,N_1722,N_1948);
and U2980 (N_2980,N_1503,N_1696);
nand U2981 (N_2981,N_1150,N_1369);
or U2982 (N_2982,N_1460,N_1259);
and U2983 (N_2983,N_1690,N_1465);
and U2984 (N_2984,N_1758,N_1016);
nor U2985 (N_2985,N_1025,N_1130);
nand U2986 (N_2986,N_1182,N_1703);
nor U2987 (N_2987,N_1370,N_1956);
or U2988 (N_2988,N_1459,N_1518);
nand U2989 (N_2989,N_1261,N_1088);
nand U2990 (N_2990,N_1354,N_1753);
and U2991 (N_2991,N_1020,N_1877);
and U2992 (N_2992,N_1435,N_1246);
and U2993 (N_2993,N_1639,N_1057);
nor U2994 (N_2994,N_1661,N_1079);
nand U2995 (N_2995,N_1849,N_1856);
and U2996 (N_2996,N_1756,N_1433);
and U2997 (N_2997,N_1479,N_1785);
or U2998 (N_2998,N_1366,N_1198);
and U2999 (N_2999,N_1606,N_1057);
nor UO_0 (O_0,N_2512,N_2802);
and UO_1 (O_1,N_2811,N_2352);
nor UO_2 (O_2,N_2896,N_2147);
or UO_3 (O_3,N_2130,N_2766);
and UO_4 (O_4,N_2342,N_2678);
nor UO_5 (O_5,N_2289,N_2132);
nand UO_6 (O_6,N_2723,N_2041);
nand UO_7 (O_7,N_2333,N_2889);
nor UO_8 (O_8,N_2614,N_2195);
or UO_9 (O_9,N_2984,N_2683);
and UO_10 (O_10,N_2250,N_2929);
nand UO_11 (O_11,N_2098,N_2061);
nor UO_12 (O_12,N_2158,N_2774);
nor UO_13 (O_13,N_2001,N_2297);
nand UO_14 (O_14,N_2496,N_2840);
or UO_15 (O_15,N_2873,N_2134);
nand UO_16 (O_16,N_2861,N_2891);
and UO_17 (O_17,N_2513,N_2322);
and UO_18 (O_18,N_2135,N_2631);
nand UO_19 (O_19,N_2470,N_2318);
or UO_20 (O_20,N_2893,N_2971);
or UO_21 (O_21,N_2137,N_2948);
nand UO_22 (O_22,N_2927,N_2223);
nand UO_23 (O_23,N_2395,N_2643);
nand UO_24 (O_24,N_2939,N_2050);
and UO_25 (O_25,N_2311,N_2899);
nor UO_26 (O_26,N_2445,N_2662);
and UO_27 (O_27,N_2016,N_2721);
xor UO_28 (O_28,N_2313,N_2773);
and UO_29 (O_29,N_2079,N_2031);
and UO_30 (O_30,N_2986,N_2654);
and UO_31 (O_31,N_2995,N_2291);
or UO_32 (O_32,N_2990,N_2494);
and UO_33 (O_33,N_2390,N_2343);
nor UO_34 (O_34,N_2373,N_2262);
and UO_35 (O_35,N_2021,N_2913);
nand UO_36 (O_36,N_2344,N_2882);
nor UO_37 (O_37,N_2286,N_2622);
nand UO_38 (O_38,N_2689,N_2266);
nand UO_39 (O_39,N_2034,N_2430);
or UO_40 (O_40,N_2081,N_2097);
and UO_41 (O_41,N_2007,N_2979);
or UO_42 (O_42,N_2531,N_2303);
and UO_43 (O_43,N_2969,N_2847);
and UO_44 (O_44,N_2642,N_2120);
or UO_45 (O_45,N_2625,N_2363);
and UO_46 (O_46,N_2366,N_2437);
or UO_47 (O_47,N_2183,N_2529);
nor UO_48 (O_48,N_2203,N_2225);
or UO_49 (O_49,N_2434,N_2329);
nor UO_50 (O_50,N_2143,N_2008);
nor UO_51 (O_51,N_2369,N_2900);
nand UO_52 (O_52,N_2895,N_2439);
nor UO_53 (O_53,N_2418,N_2645);
nand UO_54 (O_54,N_2121,N_2327);
or UO_55 (O_55,N_2535,N_2207);
nand UO_56 (O_56,N_2258,N_2566);
and UO_57 (O_57,N_2182,N_2408);
and UO_58 (O_58,N_2825,N_2385);
nand UO_59 (O_59,N_2346,N_2763);
nand UO_60 (O_60,N_2775,N_2644);
nand UO_61 (O_61,N_2960,N_2676);
nor UO_62 (O_62,N_2154,N_2688);
and UO_63 (O_63,N_2658,N_2997);
and UO_64 (O_64,N_2545,N_2166);
and UO_65 (O_65,N_2772,N_2992);
and UO_66 (O_66,N_2181,N_2810);
and UO_67 (O_67,N_2237,N_2010);
nand UO_68 (O_68,N_2495,N_2845);
nand UO_69 (O_69,N_2421,N_2150);
nor UO_70 (O_70,N_2575,N_2484);
nor UO_71 (O_71,N_2768,N_2014);
or UO_72 (O_72,N_2304,N_2024);
nand UO_73 (O_73,N_2393,N_2383);
nand UO_74 (O_74,N_2703,N_2830);
and UO_75 (O_75,N_2353,N_2521);
or UO_76 (O_76,N_2925,N_2320);
nor UO_77 (O_77,N_2454,N_2244);
nor UO_78 (O_78,N_2433,N_2011);
nand UO_79 (O_79,N_2732,N_2488);
and UO_80 (O_80,N_2798,N_2105);
nor UO_81 (O_81,N_2584,N_2469);
and UO_82 (O_82,N_2700,N_2551);
or UO_83 (O_83,N_2075,N_2285);
and UO_84 (O_84,N_2380,N_2035);
nand UO_85 (O_85,N_2485,N_2905);
or UO_86 (O_86,N_2872,N_2954);
and UO_87 (O_87,N_2666,N_2170);
or UO_88 (O_88,N_2582,N_2100);
nor UO_89 (O_89,N_2928,N_2868);
and UO_90 (O_90,N_2414,N_2836);
and UO_91 (O_91,N_2871,N_2853);
and UO_92 (O_92,N_2361,N_2432);
and UO_93 (O_93,N_2860,N_2952);
and UO_94 (O_94,N_2587,N_2419);
or UO_95 (O_95,N_2127,N_2276);
and UO_96 (O_96,N_2885,N_2140);
nand UO_97 (O_97,N_2019,N_2761);
and UO_98 (O_98,N_2719,N_2347);
and UO_99 (O_99,N_2856,N_2538);
and UO_100 (O_100,N_2842,N_2002);
nor UO_101 (O_101,N_2890,N_2686);
nor UO_102 (O_102,N_2123,N_2611);
nor UO_103 (O_103,N_2256,N_2862);
nand UO_104 (O_104,N_2965,N_2918);
and UO_105 (O_105,N_2623,N_2878);
or UO_106 (O_106,N_2606,N_2759);
nor UO_107 (O_107,N_2295,N_2424);
and UO_108 (O_108,N_2886,N_2104);
nor UO_109 (O_109,N_2255,N_2819);
and UO_110 (O_110,N_2152,N_2707);
and UO_111 (O_111,N_2006,N_2942);
or UO_112 (O_112,N_2594,N_2947);
nor UO_113 (O_113,N_2048,N_2278);
nor UO_114 (O_114,N_2972,N_2018);
nand UO_115 (O_115,N_2996,N_2959);
and UO_116 (O_116,N_2086,N_2572);
and UO_117 (O_117,N_2796,N_2530);
nor UO_118 (O_118,N_2377,N_2204);
and UO_119 (O_119,N_2777,N_2471);
or UO_120 (O_120,N_2672,N_2982);
or UO_121 (O_121,N_2839,N_2029);
or UO_122 (O_122,N_2701,N_2804);
nand UO_123 (O_123,N_2934,N_2388);
nand UO_124 (O_124,N_2790,N_2186);
or UO_125 (O_125,N_2157,N_2593);
nand UO_126 (O_126,N_2515,N_2142);
nor UO_127 (O_127,N_2174,N_2341);
or UO_128 (O_128,N_2263,N_2198);
or UO_129 (O_129,N_2667,N_2910);
or UO_130 (O_130,N_2233,N_2765);
nor UO_131 (O_131,N_2074,N_2406);
and UO_132 (O_132,N_2440,N_2312);
nor UO_133 (O_133,N_2659,N_2596);
nand UO_134 (O_134,N_2919,N_2478);
and UO_135 (O_135,N_2957,N_2897);
and UO_136 (O_136,N_2704,N_2724);
nor UO_137 (O_137,N_2630,N_2580);
nand UO_138 (O_138,N_2716,N_2187);
nand UO_139 (O_139,N_2331,N_2624);
nand UO_140 (O_140,N_2036,N_2080);
xor UO_141 (O_141,N_2980,N_2099);
nor UO_142 (O_142,N_2715,N_2475);
nand UO_143 (O_143,N_2820,N_2328);
nand UO_144 (O_144,N_2056,N_2815);
nor UO_145 (O_145,N_2206,N_2326);
and UO_146 (O_146,N_2376,N_2673);
nand UO_147 (O_147,N_2133,N_2556);
nor UO_148 (O_148,N_2310,N_2547);
nor UO_149 (O_149,N_2993,N_2912);
or UO_150 (O_150,N_2917,N_2241);
or UO_151 (O_151,N_2125,N_2946);
nor UO_152 (O_152,N_2898,N_2465);
nor UO_153 (O_153,N_2095,N_2554);
or UO_154 (O_154,N_2785,N_2527);
and UO_155 (O_155,N_2500,N_2473);
and UO_156 (O_156,N_2422,N_2746);
or UO_157 (O_157,N_2938,N_2754);
nand UO_158 (O_158,N_2935,N_2560);
and UO_159 (O_159,N_2637,N_2078);
nand UO_160 (O_160,N_2573,N_2288);
or UO_161 (O_161,N_2141,N_2139);
nor UO_162 (O_162,N_2270,N_2248);
or UO_163 (O_163,N_2949,N_2951);
nor UO_164 (O_164,N_2699,N_2359);
and UO_165 (O_165,N_2146,N_2999);
nor UO_166 (O_166,N_2950,N_2660);
nand UO_167 (O_167,N_2661,N_2641);
and UO_168 (O_168,N_2864,N_2507);
or UO_169 (O_169,N_2742,N_2401);
and UO_170 (O_170,N_2801,N_2827);
nor UO_171 (O_171,N_2536,N_2726);
nand UO_172 (O_172,N_2480,N_2677);
nor UO_173 (O_173,N_2687,N_2524);
nand UO_174 (O_174,N_2570,N_2005);
and UO_175 (O_175,N_2305,N_2583);
nand UO_176 (O_176,N_2601,N_2265);
and UO_177 (O_177,N_2605,N_2378);
nand UO_178 (O_178,N_2438,N_2447);
nand UO_179 (O_179,N_2854,N_2718);
and UO_180 (O_180,N_2943,N_2906);
or UO_181 (O_181,N_2179,N_2273);
nor UO_182 (O_182,N_2755,N_2579);
nand UO_183 (O_183,N_2136,N_2213);
nand UO_184 (O_184,N_2800,N_2160);
nand UO_185 (O_185,N_2032,N_2301);
and UO_186 (O_186,N_2240,N_2602);
or UO_187 (O_187,N_2226,N_2283);
nor UO_188 (O_188,N_2528,N_2932);
nor UO_189 (O_189,N_2298,N_2752);
nor UO_190 (O_190,N_2184,N_2442);
nor UO_191 (O_191,N_2961,N_2115);
and UO_192 (O_192,N_2128,N_2472);
or UO_193 (O_193,N_2537,N_2482);
or UO_194 (O_194,N_2268,N_2067);
nand UO_195 (O_195,N_2619,N_2409);
or UO_196 (O_196,N_2634,N_2849);
or UO_197 (O_197,N_2306,N_2370);
and UO_198 (O_198,N_2981,N_2855);
nand UO_199 (O_199,N_2784,N_2087);
nand UO_200 (O_200,N_2911,N_2779);
xor UO_201 (O_201,N_2745,N_2126);
or UO_202 (O_202,N_2806,N_2783);
nand UO_203 (O_203,N_2316,N_2574);
nor UO_204 (O_204,N_2173,N_2426);
nor UO_205 (O_205,N_2131,N_2546);
and UO_206 (O_206,N_2296,N_2571);
or UO_207 (O_207,N_2112,N_2832);
nand UO_208 (O_208,N_2324,N_2308);
nand UO_209 (O_209,N_2474,N_2835);
or UO_210 (O_210,N_2730,N_2287);
and UO_211 (O_211,N_2568,N_2684);
or UO_212 (O_212,N_2221,N_2915);
nand UO_213 (O_213,N_2931,N_2945);
or UO_214 (O_214,N_2260,N_2211);
and UO_215 (O_215,N_2168,N_2356);
nor UO_216 (O_216,N_2799,N_2358);
or UO_217 (O_217,N_2786,N_2271);
or UO_218 (O_218,N_2503,N_2231);
or UO_219 (O_219,N_2193,N_2216);
or UO_220 (O_220,N_2555,N_2543);
nor UO_221 (O_221,N_2744,N_2200);
and UO_222 (O_222,N_2145,N_2518);
and UO_223 (O_223,N_2588,N_2994);
and UO_224 (O_224,N_2553,N_2501);
nor UO_225 (O_225,N_2238,N_2229);
and UO_226 (O_226,N_2487,N_2787);
nand UO_227 (O_227,N_2397,N_2073);
and UO_228 (O_228,N_2013,N_2251);
nand UO_229 (O_229,N_2065,N_2235);
or UO_230 (O_230,N_2345,N_2788);
and UO_231 (O_231,N_2219,N_2116);
nand UO_232 (O_232,N_2818,N_2481);
and UO_233 (O_233,N_2850,N_2236);
and UO_234 (O_234,N_2043,N_2692);
nand UO_235 (O_235,N_2892,N_2936);
or UO_236 (O_236,N_2567,N_2491);
and UO_237 (O_237,N_2903,N_2817);
and UO_238 (O_238,N_2364,N_2464);
and UO_239 (O_239,N_2398,N_2416);
nand UO_240 (O_240,N_2933,N_2405);
and UO_241 (O_241,N_2693,N_2114);
nand UO_242 (O_242,N_2476,N_2460);
or UO_243 (O_243,N_2640,N_2739);
nor UO_244 (O_244,N_2330,N_2033);
nand UO_245 (O_245,N_2493,N_2793);
xor UO_246 (O_246,N_2698,N_2188);
nor UO_247 (O_247,N_2916,N_2066);
or UO_248 (O_248,N_2884,N_2824);
or UO_249 (O_249,N_2047,N_2350);
nor UO_250 (O_250,N_2646,N_2974);
and UO_251 (O_251,N_2762,N_2671);
and UO_252 (O_252,N_2983,N_2639);
and UO_253 (O_253,N_2246,N_2966);
nor UO_254 (O_254,N_2874,N_2224);
and UO_255 (O_255,N_2710,N_2425);
nand UO_256 (O_256,N_2117,N_2443);
or UO_257 (O_257,N_2448,N_2879);
nor UO_258 (O_258,N_2922,N_2463);
and UO_259 (O_259,N_2004,N_2340);
and UO_260 (O_260,N_2599,N_2563);
or UO_261 (O_261,N_2064,N_2315);
nand UO_262 (O_262,N_2000,N_2791);
nor UO_263 (O_263,N_2795,N_2046);
nand UO_264 (O_264,N_2404,N_2632);
or UO_265 (O_265,N_2412,N_2299);
and UO_266 (O_266,N_2090,N_2944);
xnor UO_267 (O_267,N_2675,N_2550);
nand UO_268 (O_268,N_2148,N_2875);
and UO_269 (O_269,N_2076,N_2321);
nand UO_270 (O_270,N_2489,N_2940);
nand UO_271 (O_271,N_2208,N_2680);
or UO_272 (O_272,N_2375,N_2748);
or UO_273 (O_273,N_2215,N_2586);
and UO_274 (O_274,N_2196,N_2924);
nand UO_275 (O_275,N_2020,N_2778);
and UO_276 (O_276,N_2264,N_2833);
or UO_277 (O_277,N_2411,N_2069);
nand UO_278 (O_278,N_2826,N_2822);
and UO_279 (O_279,N_2520,N_2275);
nand UO_280 (O_280,N_2462,N_2523);
or UO_281 (O_281,N_2807,N_2789);
nand UO_282 (O_282,N_2977,N_2456);
or UO_283 (O_283,N_2068,N_2307);
and UO_284 (O_284,N_2490,N_2539);
nand UO_285 (O_285,N_2743,N_2003);
and UO_286 (O_286,N_2816,N_2022);
nand UO_287 (O_287,N_2725,N_2504);
nor UO_288 (O_288,N_2319,N_2119);
nor UO_289 (O_289,N_2252,N_2272);
and UO_290 (O_290,N_2063,N_2357);
nand UO_291 (O_291,N_2455,N_2909);
and UO_292 (O_292,N_2269,N_2956);
nand UO_293 (O_293,N_2072,N_2055);
nor UO_294 (O_294,N_2467,N_2085);
nor UO_295 (O_295,N_2030,N_2998);
nor UO_296 (O_296,N_2389,N_2869);
or UO_297 (O_297,N_2636,N_2351);
and UO_298 (O_298,N_2760,N_2399);
and UO_299 (O_299,N_2610,N_2082);
and UO_300 (O_300,N_2335,N_2741);
nand UO_301 (O_301,N_2171,N_2505);
nor UO_302 (O_302,N_2650,N_2609);
nand UO_303 (O_303,N_2151,N_2201);
or UO_304 (O_304,N_2023,N_2060);
or UO_305 (O_305,N_2374,N_2461);
nor UO_306 (O_306,N_2348,N_2325);
or UO_307 (O_307,N_2577,N_2647);
or UO_308 (O_308,N_2092,N_2620);
nand UO_309 (O_309,N_2694,N_2058);
and UO_310 (O_310,N_2180,N_2782);
nor UO_311 (O_311,N_2453,N_2604);
nand UO_312 (O_312,N_2598,N_2210);
or UO_313 (O_313,N_2396,N_2300);
and UO_314 (O_314,N_2722,N_2163);
nor UO_315 (O_315,N_2691,N_2040);
and UO_316 (O_316,N_2205,N_2591);
or UO_317 (O_317,N_2852,N_2185);
or UO_318 (O_318,N_2459,N_2243);
nor UO_319 (O_319,N_2441,N_2870);
nand UO_320 (O_320,N_2803,N_2053);
and UO_321 (O_321,N_2449,N_2106);
and UO_322 (O_322,N_2569,N_2901);
nor UO_323 (O_323,N_2192,N_2544);
nor UO_324 (O_324,N_2532,N_2731);
and UO_325 (O_325,N_2165,N_2858);
nor UO_326 (O_326,N_2834,N_2792);
nor UO_327 (O_327,N_2987,N_2394);
nand UO_328 (O_328,N_2967,N_2930);
or UO_329 (O_329,N_2362,N_2057);
nor UO_330 (O_330,N_2403,N_2805);
nand UO_331 (O_331,N_2452,N_2985);
or UO_332 (O_332,N_2209,N_2177);
nand UO_333 (O_333,N_2780,N_2859);
and UO_334 (O_334,N_2212,N_2365);
or UO_335 (O_335,N_2156,N_2978);
or UO_336 (O_336,N_2217,N_2517);
nand UO_337 (O_337,N_2402,N_2733);
nand UO_338 (O_338,N_2338,N_2585);
or UO_339 (O_339,N_2450,N_2712);
nand UO_340 (O_340,N_2561,N_2595);
and UO_341 (O_341,N_2026,N_2410);
nor UO_342 (O_342,N_2093,N_2841);
or UO_343 (O_343,N_2902,N_2877);
nor UO_344 (O_344,N_2111,N_2129);
or UO_345 (O_345,N_2025,N_2914);
or UO_346 (O_346,N_2169,N_2628);
nand UO_347 (O_347,N_2525,N_2823);
nand UO_348 (O_348,N_2510,N_2387);
nand UO_349 (O_349,N_2663,N_2883);
nand UO_350 (O_350,N_2508,N_2468);
or UO_351 (O_351,N_2764,N_2808);
and UO_352 (O_352,N_2533,N_2103);
nand UO_353 (O_353,N_2228,N_2968);
or UO_354 (O_354,N_2565,N_2194);
nor UO_355 (O_355,N_2747,N_2175);
nand UO_356 (O_356,N_2391,N_2626);
or UO_357 (O_357,N_2670,N_2077);
and UO_358 (O_358,N_2102,N_2635);
and UO_359 (O_359,N_2037,N_2355);
nand UO_360 (O_360,N_2592,N_2138);
or UO_361 (O_361,N_2713,N_2757);
nor UO_362 (O_362,N_2540,N_2590);
and UO_363 (O_363,N_2222,N_2379);
nand UO_364 (O_364,N_2638,N_2711);
nand UO_365 (O_365,N_2814,N_2920);
or UO_366 (O_366,N_2557,N_2648);
or UO_367 (O_367,N_2282,N_2894);
nor UO_368 (O_368,N_2242,N_2172);
and UO_369 (O_369,N_2564,N_2696);
and UO_370 (O_370,N_2851,N_2091);
nor UO_371 (O_371,N_2962,N_2697);
nor UO_372 (O_372,N_2429,N_2876);
xor UO_373 (O_373,N_2857,N_2279);
nor UO_374 (O_374,N_2576,N_2973);
nand UO_375 (O_375,N_2039,N_2627);
xor UO_376 (O_376,N_2562,N_2514);
or UO_377 (O_377,N_2431,N_2214);
and UO_378 (O_378,N_2812,N_2578);
or UO_379 (O_379,N_2653,N_2451);
and UO_380 (O_380,N_2124,N_2371);
nor UO_381 (O_381,N_2281,N_2234);
or UO_382 (O_382,N_2109,N_2497);
nand UO_383 (O_383,N_2354,N_2094);
and UO_384 (O_384,N_2734,N_2831);
nand UO_385 (O_385,N_2821,N_2261);
or UO_386 (O_386,N_2277,N_2336);
nand UO_387 (O_387,N_2669,N_2519);
and UO_388 (O_388,N_2436,N_2012);
nor UO_389 (O_389,N_2446,N_2991);
or UO_390 (O_390,N_2809,N_2332);
nand UO_391 (O_391,N_2665,N_2612);
nand UO_392 (O_392,N_2649,N_2413);
or UO_393 (O_393,N_2729,N_2717);
nor UO_394 (O_394,N_2753,N_2400);
and UO_395 (O_395,N_2655,N_2202);
and UO_396 (O_396,N_2613,N_2089);
and UO_397 (O_397,N_2280,N_2552);
nor UO_398 (O_398,N_2907,N_2458);
nor UO_399 (O_399,N_2737,N_2190);
and UO_400 (O_400,N_2964,N_2837);
and UO_401 (O_401,N_2028,N_2045);
and UO_402 (O_402,N_2382,N_2617);
nand UO_403 (O_403,N_2049,N_2958);
nand UO_404 (O_404,N_2110,N_2153);
or UO_405 (O_405,N_2904,N_2302);
nor UO_406 (O_406,N_2600,N_2702);
nor UO_407 (O_407,N_2339,N_2953);
nor UO_408 (O_408,N_2534,N_2071);
and UO_409 (O_409,N_2155,N_2386);
nor UO_410 (O_410,N_2084,N_2674);
and UO_411 (O_411,N_2955,N_2756);
nand UO_412 (O_412,N_2230,N_2970);
and UO_413 (O_413,N_2232,N_2865);
nor UO_414 (O_414,N_2096,N_2027);
or UO_415 (O_415,N_2381,N_2227);
or UO_416 (O_416,N_2257,N_2829);
nand UO_417 (O_417,N_2740,N_2542);
and UO_418 (O_418,N_2923,N_2603);
xor UO_419 (O_419,N_2516,N_2247);
or UO_420 (O_420,N_2477,N_2770);
nand UO_421 (O_421,N_2709,N_2615);
or UO_422 (O_422,N_2976,N_2767);
or UO_423 (O_423,N_2771,N_2334);
nor UO_424 (O_424,N_2813,N_2988);
or UO_425 (O_425,N_2314,N_2368);
and UO_426 (O_426,N_2199,N_2108);
or UO_427 (O_427,N_2652,N_2083);
nor UO_428 (O_428,N_2926,N_2038);
nand UO_429 (O_429,N_2846,N_2616);
and UO_430 (O_430,N_2685,N_2866);
nor UO_431 (O_431,N_2781,N_2867);
nor UO_432 (O_432,N_2618,N_2164);
nand UO_433 (O_433,N_2017,N_2113);
nand UO_434 (O_434,N_2176,N_2526);
nor UO_435 (O_435,N_2118,N_2758);
and UO_436 (O_436,N_2415,N_2509);
and UO_437 (O_437,N_2062,N_2621);
nor UO_438 (O_438,N_2372,N_2690);
nor UO_439 (O_439,N_2597,N_2695);
nor UO_440 (O_440,N_2466,N_2880);
or UO_441 (O_441,N_2292,N_2284);
and UO_442 (O_442,N_2122,N_2502);
nor UO_443 (O_443,N_2054,N_2921);
or UO_444 (O_444,N_2423,N_2738);
and UO_445 (O_445,N_2167,N_2989);
or UO_446 (O_446,N_2706,N_2975);
nand UO_447 (O_447,N_2051,N_2589);
or UO_448 (O_448,N_2349,N_2708);
or UO_449 (O_449,N_2720,N_2681);
nand UO_450 (O_450,N_2189,N_2838);
nand UO_451 (O_451,N_2843,N_2178);
nor UO_452 (O_452,N_2479,N_2161);
nand UO_453 (O_453,N_2052,N_2367);
nor UO_454 (O_454,N_2664,N_2457);
nor UO_455 (O_455,N_2323,N_2267);
nor UO_456 (O_456,N_2444,N_2101);
nor UO_457 (O_457,N_2888,N_2633);
and UO_458 (O_458,N_2254,N_2797);
and UO_459 (O_459,N_2728,N_2548);
nor UO_460 (O_460,N_2218,N_2015);
nand UO_461 (O_461,N_2656,N_2191);
nand UO_462 (O_462,N_2144,N_2435);
or UO_463 (O_463,N_2506,N_2522);
or UO_464 (O_464,N_2417,N_2294);
and UO_465 (O_465,N_2309,N_2149);
and UO_466 (O_466,N_2486,N_2629);
nand UO_467 (O_467,N_2088,N_2274);
or UO_468 (O_468,N_2937,N_2657);
nand UO_469 (O_469,N_2483,N_2751);
nor UO_470 (O_470,N_2668,N_2259);
or UO_471 (O_471,N_2735,N_2608);
and UO_472 (O_472,N_2750,N_2197);
and UO_473 (O_473,N_2941,N_2360);
nand UO_474 (O_474,N_2558,N_2682);
nor UO_475 (O_475,N_2492,N_2290);
xnor UO_476 (O_476,N_2249,N_2392);
nand UO_477 (O_477,N_2863,N_2776);
nor UO_478 (O_478,N_2317,N_2794);
nand UO_479 (O_479,N_2384,N_2337);
nand UO_480 (O_480,N_2651,N_2844);
and UO_481 (O_481,N_2159,N_2407);
nor UO_482 (O_482,N_2559,N_2705);
or UO_483 (O_483,N_2427,N_2511);
nand UO_484 (O_484,N_2428,N_2107);
nor UO_485 (O_485,N_2581,N_2220);
or UO_486 (O_486,N_2679,N_2245);
nor UO_487 (O_487,N_2499,N_2714);
and UO_488 (O_488,N_2239,N_2070);
and UO_489 (O_489,N_2549,N_2420);
or UO_490 (O_490,N_2881,N_2908);
nor UO_491 (O_491,N_2009,N_2498);
nor UO_492 (O_492,N_2044,N_2887);
or UO_493 (O_493,N_2736,N_2828);
nor UO_494 (O_494,N_2293,N_2541);
or UO_495 (O_495,N_2607,N_2253);
and UO_496 (O_496,N_2059,N_2963);
nor UO_497 (O_497,N_2848,N_2749);
nand UO_498 (O_498,N_2162,N_2042);
nor UO_499 (O_499,N_2727,N_2769);
endmodule