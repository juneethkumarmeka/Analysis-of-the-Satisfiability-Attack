module basic_1000_10000_1500_20_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_586,In_549);
and U1 (N_1,In_722,In_627);
and U2 (N_2,In_884,In_705);
or U3 (N_3,In_879,In_874);
nor U4 (N_4,In_995,In_249);
or U5 (N_5,In_297,In_106);
nor U6 (N_6,In_415,In_363);
or U7 (N_7,In_585,In_907);
or U8 (N_8,In_910,In_111);
nand U9 (N_9,In_840,In_308);
and U10 (N_10,In_829,In_669);
nor U11 (N_11,In_851,In_442);
and U12 (N_12,In_554,In_649);
and U13 (N_13,In_285,In_317);
nand U14 (N_14,In_692,In_16);
and U15 (N_15,In_584,In_286);
or U16 (N_16,In_750,In_487);
nor U17 (N_17,In_24,In_519);
nor U18 (N_18,In_524,In_352);
or U19 (N_19,In_839,In_182);
nor U20 (N_20,In_79,In_288);
nor U21 (N_21,In_623,In_136);
xor U22 (N_22,In_609,In_812);
nor U23 (N_23,In_278,In_339);
or U24 (N_24,In_382,In_253);
nand U25 (N_25,In_849,In_837);
and U26 (N_26,In_726,In_731);
or U27 (N_27,In_762,In_915);
nor U28 (N_28,In_872,In_246);
nand U29 (N_29,In_662,In_341);
and U30 (N_30,In_261,In_809);
nand U31 (N_31,In_818,In_203);
or U32 (N_32,In_117,In_282);
nand U33 (N_33,In_606,In_796);
and U34 (N_34,In_979,In_494);
nor U35 (N_35,In_406,In_330);
nor U36 (N_36,In_798,In_174);
nor U37 (N_37,In_362,In_958);
nor U38 (N_38,In_121,In_630);
nand U39 (N_39,In_289,In_758);
nand U40 (N_40,In_313,In_541);
nor U41 (N_41,In_694,In_154);
or U42 (N_42,In_294,In_759);
nor U43 (N_43,In_523,In_999);
nor U44 (N_44,In_882,In_583);
and U45 (N_45,In_336,In_525);
and U46 (N_46,In_27,In_219);
and U47 (N_47,In_160,In_472);
nor U48 (N_48,In_45,In_925);
nand U49 (N_49,In_828,In_986);
nor U50 (N_50,In_903,In_82);
nor U51 (N_51,In_299,In_34);
nand U52 (N_52,In_899,In_187);
nor U53 (N_53,In_582,In_344);
nand U54 (N_54,In_239,In_464);
xor U55 (N_55,In_180,In_469);
nor U56 (N_56,In_949,In_658);
or U57 (N_57,In_384,In_205);
and U58 (N_58,In_67,In_735);
and U59 (N_59,In_431,In_784);
or U60 (N_60,In_416,In_351);
nor U61 (N_61,In_404,In_477);
and U62 (N_62,In_625,In_268);
or U63 (N_63,In_452,In_80);
and U64 (N_64,In_432,In_795);
or U65 (N_65,In_240,In_786);
and U66 (N_66,In_752,In_488);
nand U67 (N_67,In_801,In_982);
and U68 (N_68,In_257,In_28);
nor U69 (N_69,In_624,In_921);
nor U70 (N_70,In_806,In_232);
nand U71 (N_71,In_565,In_230);
or U72 (N_72,In_231,In_610);
and U73 (N_73,In_515,In_139);
and U74 (N_74,In_94,In_573);
and U75 (N_75,In_858,In_763);
nand U76 (N_76,In_14,In_57);
nor U77 (N_77,In_577,In_777);
nand U78 (N_78,In_968,In_667);
nor U79 (N_79,In_683,In_674);
nand U80 (N_80,In_420,In_281);
nand U81 (N_81,In_920,In_428);
nor U82 (N_82,In_615,In_127);
or U83 (N_83,In_888,In_574);
nor U84 (N_84,In_597,In_776);
or U85 (N_85,In_407,In_42);
and U86 (N_86,In_272,In_126);
and U87 (N_87,In_900,In_376);
nand U88 (N_88,In_747,In_811);
nor U89 (N_89,In_755,In_935);
and U90 (N_90,In_846,In_97);
or U91 (N_91,In_275,In_262);
nor U92 (N_92,In_538,In_719);
nand U93 (N_93,In_33,In_697);
nor U94 (N_94,In_419,In_737);
nor U95 (N_95,In_417,In_964);
nand U96 (N_96,In_400,In_62);
nand U97 (N_97,In_401,In_490);
nor U98 (N_98,In_137,In_75);
nand U99 (N_99,In_558,In_41);
nor U100 (N_100,In_173,In_414);
nand U101 (N_101,In_808,In_58);
and U102 (N_102,In_778,In_65);
nor U103 (N_103,In_192,In_242);
or U104 (N_104,In_608,In_591);
nand U105 (N_105,In_437,In_314);
and U106 (N_106,In_581,In_63);
and U107 (N_107,In_244,In_619);
nand U108 (N_108,In_512,In_838);
nand U109 (N_109,In_145,In_571);
nand U110 (N_110,In_875,In_822);
or U111 (N_111,In_652,In_229);
nor U112 (N_112,In_164,In_817);
nor U113 (N_113,In_924,In_596);
nor U114 (N_114,In_491,In_628);
nor U115 (N_115,In_380,In_506);
nor U116 (N_116,In_760,In_265);
nand U117 (N_117,In_302,In_489);
or U118 (N_118,In_73,In_359);
nand U119 (N_119,In_932,In_774);
xnor U120 (N_120,In_883,In_725);
and U121 (N_121,In_396,In_381);
or U122 (N_122,In_251,In_734);
or U123 (N_123,In_871,In_789);
or U124 (N_124,In_35,In_690);
or U125 (N_125,In_592,In_678);
or U126 (N_126,In_657,In_555);
and U127 (N_127,In_587,In_71);
nand U128 (N_128,In_507,In_171);
nor U129 (N_129,In_21,In_181);
nor U130 (N_130,In_948,In_699);
and U131 (N_131,In_805,In_183);
nand U132 (N_132,In_168,In_685);
and U133 (N_133,In_748,In_559);
and U134 (N_134,In_670,In_783);
nand U135 (N_135,In_746,In_112);
nand U136 (N_136,In_594,In_47);
or U137 (N_137,In_455,In_102);
nor U138 (N_138,In_862,In_712);
or U139 (N_139,In_6,In_761);
nand U140 (N_140,In_100,In_859);
xor U141 (N_141,In_751,In_757);
or U142 (N_142,In_354,In_668);
nor U143 (N_143,In_970,In_607);
or U144 (N_144,In_589,In_207);
nor U145 (N_145,In_844,In_482);
and U146 (N_146,In_350,In_315);
nand U147 (N_147,In_312,In_379);
or U148 (N_148,In_61,In_470);
nand U149 (N_149,In_20,In_535);
and U150 (N_150,In_435,In_505);
nor U151 (N_151,In_123,In_894);
nor U152 (N_152,In_377,In_119);
or U153 (N_153,In_998,In_532);
nor U154 (N_154,In_328,In_992);
nand U155 (N_155,In_681,In_409);
or U156 (N_156,In_551,In_850);
and U157 (N_157,In_768,In_296);
nand U158 (N_158,In_572,In_287);
or U159 (N_159,In_638,In_797);
and U160 (N_160,In_516,In_947);
or U161 (N_161,In_614,In_309);
nor U162 (N_162,In_270,In_708);
nand U163 (N_163,In_981,In_247);
or U164 (N_164,In_886,In_601);
nand U165 (N_165,In_238,In_503);
and U166 (N_166,In_468,In_766);
or U167 (N_167,In_660,In_753);
nand U168 (N_168,In_895,In_785);
nor U169 (N_169,In_787,In_855);
nand U170 (N_170,In_646,In_741);
xnor U171 (N_171,In_663,In_353);
and U172 (N_172,In_412,In_700);
nor U173 (N_173,In_7,In_902);
or U174 (N_174,In_526,In_653);
nand U175 (N_175,In_484,In_711);
nor U176 (N_176,In_718,In_984);
nand U177 (N_177,In_953,In_108);
xor U178 (N_178,In_923,In_133);
and U179 (N_179,In_889,In_720);
or U180 (N_180,In_603,In_939);
or U181 (N_181,In_157,In_514);
nand U182 (N_182,In_856,In_233);
xor U183 (N_183,In_178,In_727);
or U184 (N_184,In_337,In_938);
nand U185 (N_185,In_371,In_621);
nand U186 (N_186,In_937,In_418);
nor U187 (N_187,In_590,In_197);
or U188 (N_188,In_733,In_616);
or U189 (N_189,In_989,In_728);
nor U190 (N_190,In_25,In_360);
nand U191 (N_191,In_283,In_633);
nor U192 (N_192,In_854,In_237);
and U193 (N_193,In_322,In_991);
nand U194 (N_194,In_965,In_345);
and U195 (N_195,In_411,In_248);
or U196 (N_196,In_550,In_1);
nand U197 (N_197,In_522,In_451);
xnor U198 (N_198,In_803,In_513);
nand U199 (N_199,In_403,In_676);
and U200 (N_200,In_765,In_185);
nand U201 (N_201,In_501,In_531);
nand U202 (N_202,In_194,In_717);
nor U203 (N_203,In_475,In_366);
or U204 (N_204,In_520,In_905);
and U205 (N_205,In_402,In_880);
nand U206 (N_206,In_511,In_764);
nand U207 (N_207,In_266,In_885);
nand U208 (N_208,In_713,In_26);
nor U209 (N_209,In_413,In_144);
nor U210 (N_210,In_68,In_665);
and U211 (N_211,In_323,In_693);
nor U212 (N_212,In_698,In_456);
or U213 (N_213,In_945,In_51);
nand U214 (N_214,In_466,In_374);
and U215 (N_215,In_710,In_199);
nand U216 (N_216,In_934,In_93);
nand U217 (N_217,In_537,In_952);
or U218 (N_218,In_88,In_729);
nor U219 (N_219,In_426,In_191);
nor U220 (N_220,In_509,In_890);
and U221 (N_221,In_429,In_325);
nand U222 (N_222,In_834,In_162);
nor U223 (N_223,In_825,In_928);
or U224 (N_224,In_504,In_101);
or U225 (N_225,In_643,In_993);
nor U226 (N_226,In_457,In_876);
and U227 (N_227,In_897,In_156);
xnor U228 (N_228,In_129,In_595);
or U229 (N_229,In_664,In_990);
nand U230 (N_230,In_857,In_440);
nand U231 (N_231,In_780,In_405);
nand U232 (N_232,In_90,In_389);
or U233 (N_233,In_629,In_12);
nand U234 (N_234,In_835,In_276);
and U235 (N_235,In_906,In_118);
xor U236 (N_236,In_691,In_175);
nand U237 (N_237,In_357,In_214);
nand U238 (N_238,In_815,In_479);
nor U239 (N_239,In_721,In_96);
xor U240 (N_240,In_454,In_48);
or U241 (N_241,In_974,In_386);
and U242 (N_242,In_116,In_533);
or U243 (N_243,In_518,In_206);
or U244 (N_244,In_4,In_87);
nor U245 (N_245,In_800,In_148);
or U246 (N_246,In_642,In_44);
nand U247 (N_247,In_211,In_320);
or U248 (N_248,In_611,In_226);
and U249 (N_249,In_802,In_893);
nand U250 (N_250,In_770,In_54);
nor U251 (N_251,In_172,In_52);
nand U252 (N_252,In_543,In_866);
nor U253 (N_253,In_19,In_997);
nand U254 (N_254,In_204,In_13);
and U255 (N_255,In_791,In_147);
or U256 (N_256,In_447,In_613);
nand U257 (N_257,In_891,In_213);
nor U258 (N_258,In_43,In_562);
or U259 (N_259,In_749,In_395);
nor U260 (N_260,In_843,In_545);
nand U261 (N_261,In_909,In_686);
nor U262 (N_262,In_2,In_298);
nor U263 (N_263,In_985,In_847);
or U264 (N_264,In_680,In_50);
or U265 (N_265,In_263,In_254);
and U266 (N_266,In_704,In_59);
or U267 (N_267,In_709,In_422);
or U268 (N_268,In_40,In_461);
and U269 (N_269,In_655,In_324);
nand U270 (N_270,In_914,In_159);
nor U271 (N_271,In_772,In_198);
nor U272 (N_272,In_305,In_340);
and U273 (N_273,In_256,In_433);
and U274 (N_274,In_496,In_385);
or U275 (N_275,In_132,In_779);
xor U276 (N_276,In_771,In_95);
nor U277 (N_277,In_332,In_598);
and U278 (N_278,In_140,In_868);
nor U279 (N_279,In_158,In_91);
nor U280 (N_280,In_193,In_579);
nand U281 (N_281,In_845,In_319);
and U282 (N_282,In_439,In_383);
nor U283 (N_283,In_222,In_223);
or U284 (N_284,In_841,In_122);
or U285 (N_285,In_647,In_234);
and U286 (N_286,In_290,In_736);
xnor U287 (N_287,In_284,In_273);
and U288 (N_288,In_936,In_943);
and U289 (N_289,In_146,In_605);
xnor U290 (N_290,In_819,In_84);
and U291 (N_291,In_529,In_955);
nor U292 (N_292,In_602,In_176);
or U293 (N_293,In_863,In_926);
xnor U294 (N_294,In_556,In_218);
xnor U295 (N_295,In_500,In_618);
and U296 (N_296,In_306,In_36);
nand U297 (N_297,In_831,In_311);
nor U298 (N_298,In_166,In_575);
or U299 (N_299,In_696,In_957);
and U300 (N_300,In_987,In_639);
nand U301 (N_301,In_425,In_481);
nor U302 (N_302,In_170,In_620);
and U303 (N_303,In_567,In_980);
nand U304 (N_304,In_155,In_196);
nor U305 (N_305,In_799,In_216);
or U306 (N_306,In_508,In_202);
or U307 (N_307,In_954,In_852);
nand U308 (N_308,In_743,In_944);
nand U309 (N_309,In_347,In_916);
nand U310 (N_310,In_604,In_390);
xnor U311 (N_311,In_378,In_372);
nand U312 (N_312,In_730,In_988);
and U313 (N_313,In_576,In_66);
or U314 (N_314,In_732,In_243);
or U315 (N_315,In_568,In_996);
nor U316 (N_316,In_626,In_521);
nand U317 (N_317,In_274,In_959);
or U318 (N_318,In_271,In_326);
nand U319 (N_319,In_430,In_307);
and U320 (N_320,In_49,In_994);
nor U321 (N_321,In_295,In_460);
nand U322 (N_322,In_17,In_807);
and U323 (N_323,In_373,In_677);
or U324 (N_324,In_0,In_3);
or U325 (N_325,In_612,In_338);
or U326 (N_326,In_105,In_967);
and U327 (N_327,In_972,In_107);
nor U328 (N_328,In_744,In_930);
nand U329 (N_329,In_962,In_637);
or U330 (N_330,In_104,In_640);
nor U331 (N_331,In_177,In_99);
xnor U332 (N_332,In_816,In_528);
nand U333 (N_333,In_31,In_10);
and U334 (N_334,In_189,In_445);
and U335 (N_335,In_53,In_450);
or U336 (N_336,In_634,In_631);
nor U337 (N_337,In_498,In_682);
xor U338 (N_338,In_887,In_22);
xor U339 (N_339,In_277,In_334);
nor U340 (N_340,In_645,In_135);
nand U341 (N_341,In_280,In_865);
or U342 (N_342,In_836,In_740);
xor U343 (N_343,In_536,In_81);
and U344 (N_344,In_570,In_301);
nand U345 (N_345,In_689,In_723);
nand U346 (N_346,In_788,In_349);
and U347 (N_347,In_78,In_901);
and U348 (N_348,In_331,In_599);
xnor U349 (N_349,In_76,In_580);
or U350 (N_350,In_142,In_169);
or U351 (N_351,In_397,In_527);
nor U352 (N_352,In_632,In_410);
nand U353 (N_353,In_37,In_441);
nor U354 (N_354,In_375,In_557);
nor U355 (N_355,In_92,In_898);
or U356 (N_356,In_255,In_85);
nor U357 (N_357,In_224,In_832);
or U358 (N_358,In_421,In_186);
or U359 (N_359,In_961,In_60);
nor U360 (N_360,In_150,In_495);
nand U361 (N_361,In_480,In_814);
nand U362 (N_362,In_120,In_756);
nor U363 (N_363,In_617,In_929);
nor U364 (N_364,In_70,In_424);
nand U365 (N_365,In_911,In_29);
or U366 (N_366,In_208,In_449);
nand U367 (N_367,In_361,In_547);
nor U368 (N_368,In_673,In_473);
and U369 (N_369,In_695,In_963);
nand U370 (N_370,In_179,In_824);
or U371 (N_371,In_392,In_892);
nor U372 (N_372,In_103,In_552);
nor U373 (N_373,In_11,In_217);
or U374 (N_374,In_622,In_861);
and U375 (N_375,In_540,In_56);
or U376 (N_376,In_684,In_259);
nor U377 (N_377,In_399,In_745);
or U378 (N_378,In_942,In_548);
nand U379 (N_379,In_804,In_292);
or U380 (N_380,In_364,In_388);
or U381 (N_381,In_754,In_134);
and U382 (N_382,In_739,In_188);
and U383 (N_383,In_109,In_792);
nor U384 (N_384,In_499,In_195);
or U385 (N_385,In_235,In_827);
and U386 (N_386,In_190,In_453);
nand U387 (N_387,In_293,In_365);
nand U388 (N_388,In_300,In_648);
nand U389 (N_389,In_530,In_842);
or U390 (N_390,In_702,In_114);
nor U391 (N_391,In_333,In_98);
and U392 (N_392,In_877,In_486);
and U393 (N_393,In_544,In_370);
nor U394 (N_394,In_260,In_149);
nor U395 (N_395,In_975,In_252);
nor U396 (N_396,In_654,In_671);
or U397 (N_397,In_342,In_941);
and U398 (N_398,In_201,In_458);
and U399 (N_399,In_769,In_978);
nor U400 (N_400,In_927,In_321);
xnor U401 (N_401,In_553,In_200);
or U402 (N_402,In_343,In_69);
or U403 (N_403,In_74,In_316);
nor U404 (N_404,In_115,In_9);
nand U405 (N_405,In_775,In_912);
or U406 (N_406,In_327,In_656);
xor U407 (N_407,In_356,In_138);
or U408 (N_408,In_55,In_64);
or U409 (N_409,In_641,In_600);
nor U410 (N_410,In_922,In_971);
and U411 (N_411,In_666,In_904);
and U412 (N_412,In_870,In_896);
or U413 (N_413,In_387,In_706);
xnor U414 (N_414,In_933,In_742);
nor U415 (N_415,In_661,In_566);
nor U416 (N_416,In_860,In_210);
xnor U417 (N_417,In_569,In_644);
nand U418 (N_418,In_782,In_434);
or U419 (N_419,In_436,In_77);
nand U420 (N_420,In_83,In_588);
or U421 (N_421,In_30,In_5);
and U422 (N_422,In_820,In_474);
xor U423 (N_423,In_368,In_833);
or U424 (N_424,In_221,In_960);
or U425 (N_425,In_346,In_561);
nand U426 (N_426,In_716,In_908);
and U427 (N_427,In_701,In_534);
and U428 (N_428,In_39,In_335);
nor U429 (N_429,In_355,In_810);
nor U430 (N_430,In_969,In_423);
and U431 (N_431,In_369,In_113);
or U432 (N_432,In_738,In_125);
nand U433 (N_433,In_593,In_636);
and U434 (N_434,In_220,In_279);
nor U435 (N_435,In_258,In_215);
nand U436 (N_436,In_153,In_881);
nor U437 (N_437,In_209,In_241);
and U438 (N_438,In_228,In_560);
nor U439 (N_439,In_715,In_225);
and U440 (N_440,In_651,In_141);
xnor U441 (N_441,In_476,In_869);
and U442 (N_442,In_250,In_227);
and U443 (N_443,In_483,In_86);
or U444 (N_444,In_983,In_635);
and U445 (N_445,In_956,In_165);
nand U446 (N_446,In_950,In_853);
nor U447 (N_447,In_394,In_391);
nand U448 (N_448,In_790,In_448);
xnor U449 (N_449,In_563,In_358);
nand U450 (N_450,In_465,In_767);
nor U451 (N_451,In_38,In_236);
or U452 (N_452,In_46,In_152);
or U453 (N_453,In_269,In_438);
and U454 (N_454,In_781,In_446);
nor U455 (N_455,In_151,In_539);
or U456 (N_456,In_471,In_813);
or U457 (N_457,In_502,In_492);
or U458 (N_458,In_703,In_462);
or U459 (N_459,In_650,In_823);
and U460 (N_460,In_267,In_245);
and U461 (N_461,In_793,In_714);
and U462 (N_462,In_794,In_517);
or U463 (N_463,In_18,In_546);
or U464 (N_464,In_578,In_329);
or U465 (N_465,In_687,In_542);
nand U466 (N_466,In_485,In_675);
nand U467 (N_467,In_163,In_15);
nand U468 (N_468,In_873,In_143);
or U469 (N_469,In_493,In_564);
nand U470 (N_470,In_124,In_72);
nor U471 (N_471,In_848,In_773);
or U472 (N_472,In_478,In_89);
and U473 (N_473,In_303,In_917);
and U474 (N_474,In_348,In_167);
or U475 (N_475,In_32,In_398);
and U476 (N_476,In_212,In_310);
nor U477 (N_477,In_497,In_264);
or U478 (N_478,In_976,In_830);
nor U479 (N_479,In_161,In_688);
and U480 (N_480,In_110,In_966);
and U481 (N_481,In_919,In_443);
nor U482 (N_482,In_973,In_659);
nor U483 (N_483,In_408,In_821);
nand U484 (N_484,In_913,In_940);
or U485 (N_485,In_931,In_444);
nor U486 (N_486,In_724,In_393);
xor U487 (N_487,In_679,In_23);
or U488 (N_488,In_318,In_672);
nand U489 (N_489,In_304,In_878);
nor U490 (N_490,In_427,In_951);
and U491 (N_491,In_128,In_946);
or U492 (N_492,In_291,In_918);
nor U493 (N_493,In_864,In_8);
nor U494 (N_494,In_459,In_367);
and U495 (N_495,In_184,In_867);
or U496 (N_496,In_707,In_977);
nand U497 (N_497,In_510,In_130);
nand U498 (N_498,In_131,In_463);
nor U499 (N_499,In_826,In_467);
and U500 (N_500,N_162,N_51);
nand U501 (N_501,N_155,N_297);
or U502 (N_502,N_475,N_274);
and U503 (N_503,N_181,N_138);
nand U504 (N_504,N_68,N_486);
and U505 (N_505,N_298,N_89);
nand U506 (N_506,N_437,N_380);
nand U507 (N_507,N_344,N_163);
xor U508 (N_508,N_374,N_360);
xor U509 (N_509,N_400,N_407);
nor U510 (N_510,N_498,N_253);
nor U511 (N_511,N_225,N_264);
and U512 (N_512,N_174,N_137);
or U513 (N_513,N_135,N_71);
or U514 (N_514,N_223,N_19);
nor U515 (N_515,N_436,N_122);
nor U516 (N_516,N_247,N_170);
nor U517 (N_517,N_60,N_200);
xor U518 (N_518,N_457,N_58);
and U519 (N_519,N_32,N_289);
or U520 (N_520,N_140,N_364);
nor U521 (N_521,N_202,N_219);
nand U522 (N_522,N_301,N_132);
or U523 (N_523,N_193,N_314);
and U524 (N_524,N_397,N_358);
or U525 (N_525,N_319,N_245);
and U526 (N_526,N_459,N_266);
nand U527 (N_527,N_473,N_487);
nand U528 (N_528,N_418,N_50);
nand U529 (N_529,N_82,N_111);
nor U530 (N_530,N_256,N_139);
and U531 (N_531,N_307,N_496);
or U532 (N_532,N_441,N_405);
nand U533 (N_533,N_377,N_399);
nand U534 (N_534,N_331,N_273);
nand U535 (N_535,N_131,N_294);
nand U536 (N_536,N_218,N_446);
and U537 (N_537,N_56,N_371);
and U538 (N_538,N_101,N_166);
nor U539 (N_539,N_302,N_309);
and U540 (N_540,N_370,N_287);
xnor U541 (N_541,N_185,N_337);
or U542 (N_542,N_291,N_171);
and U543 (N_543,N_278,N_367);
nand U544 (N_544,N_299,N_433);
and U545 (N_545,N_444,N_235);
and U546 (N_546,N_464,N_110);
nand U547 (N_547,N_39,N_308);
nand U548 (N_548,N_17,N_414);
nor U549 (N_549,N_197,N_93);
nor U550 (N_550,N_187,N_366);
or U551 (N_551,N_252,N_312);
or U552 (N_552,N_43,N_25);
and U553 (N_553,N_28,N_73);
and U554 (N_554,N_121,N_44);
or U555 (N_555,N_325,N_488);
nand U556 (N_556,N_124,N_199);
or U557 (N_557,N_410,N_454);
nand U558 (N_558,N_15,N_318);
nor U559 (N_559,N_282,N_64);
nor U560 (N_560,N_396,N_21);
nor U561 (N_561,N_458,N_177);
or U562 (N_562,N_383,N_494);
or U563 (N_563,N_434,N_201);
or U564 (N_564,N_0,N_412);
and U565 (N_565,N_330,N_402);
and U566 (N_566,N_88,N_86);
and U567 (N_567,N_362,N_231);
nand U568 (N_568,N_36,N_455);
xor U569 (N_569,N_203,N_365);
or U570 (N_570,N_161,N_127);
nand U571 (N_571,N_408,N_211);
nor U572 (N_572,N_26,N_246);
nor U573 (N_573,N_279,N_347);
or U574 (N_574,N_439,N_403);
nor U575 (N_575,N_315,N_456);
xnor U576 (N_576,N_61,N_41);
and U577 (N_577,N_34,N_173);
nor U578 (N_578,N_416,N_341);
nor U579 (N_579,N_381,N_428);
nor U580 (N_580,N_189,N_151);
or U581 (N_581,N_244,N_196);
nor U582 (N_582,N_240,N_495);
and U583 (N_583,N_372,N_417);
or U584 (N_584,N_102,N_37);
nand U585 (N_585,N_443,N_76);
xor U586 (N_586,N_492,N_80);
and U587 (N_587,N_157,N_484);
nand U588 (N_588,N_394,N_236);
nand U589 (N_589,N_481,N_250);
and U590 (N_590,N_42,N_438);
nand U591 (N_591,N_263,N_2);
or U592 (N_592,N_213,N_257);
nand U593 (N_593,N_390,N_97);
xor U594 (N_594,N_284,N_237);
or U595 (N_595,N_66,N_106);
xnor U596 (N_596,N_474,N_178);
nand U597 (N_597,N_119,N_316);
nor U598 (N_598,N_207,N_379);
nor U599 (N_599,N_425,N_96);
nand U600 (N_600,N_74,N_99);
nand U601 (N_601,N_69,N_453);
or U602 (N_602,N_483,N_491);
xnor U603 (N_603,N_349,N_313);
nor U604 (N_604,N_206,N_352);
nand U605 (N_605,N_471,N_467);
nand U606 (N_606,N_75,N_345);
nor U607 (N_607,N_415,N_104);
xnor U608 (N_608,N_343,N_290);
nor U609 (N_609,N_227,N_461);
or U610 (N_610,N_241,N_98);
nand U611 (N_611,N_280,N_239);
nor U612 (N_612,N_338,N_270);
and U613 (N_613,N_462,N_62);
nand U614 (N_614,N_259,N_67);
xor U615 (N_615,N_322,N_172);
nor U616 (N_616,N_142,N_375);
nand U617 (N_617,N_215,N_126);
and U618 (N_618,N_490,N_5);
nand U619 (N_619,N_11,N_169);
nand U620 (N_620,N_497,N_499);
or U621 (N_621,N_328,N_6);
and U622 (N_622,N_145,N_160);
nor U623 (N_623,N_478,N_317);
nor U624 (N_624,N_175,N_321);
and U625 (N_625,N_267,N_389);
nand U626 (N_626,N_156,N_342);
nand U627 (N_627,N_233,N_85);
nor U628 (N_628,N_391,N_254);
nand U629 (N_629,N_350,N_9);
nand U630 (N_630,N_183,N_447);
nand U631 (N_631,N_116,N_485);
or U632 (N_632,N_216,N_269);
nor U633 (N_633,N_353,N_30);
and U634 (N_634,N_78,N_288);
nor U635 (N_635,N_329,N_165);
nand U636 (N_636,N_466,N_105);
nor U637 (N_637,N_31,N_188);
and U638 (N_638,N_430,N_123);
nor U639 (N_639,N_84,N_136);
nor U640 (N_640,N_351,N_112);
and U641 (N_641,N_262,N_8);
or U642 (N_642,N_310,N_406);
nand U643 (N_643,N_150,N_260);
nand U644 (N_644,N_452,N_117);
or U645 (N_645,N_335,N_450);
xnor U646 (N_646,N_184,N_45);
and U647 (N_647,N_118,N_369);
nor U648 (N_648,N_376,N_55);
or U649 (N_649,N_432,N_272);
nand U650 (N_650,N_48,N_332);
or U651 (N_651,N_388,N_420);
and U652 (N_652,N_384,N_209);
and U653 (N_653,N_232,N_182);
nand U654 (N_654,N_445,N_482);
or U655 (N_655,N_324,N_361);
nor U656 (N_656,N_354,N_95);
xor U657 (N_657,N_27,N_13);
nor U658 (N_658,N_83,N_275);
nand U659 (N_659,N_24,N_271);
and U660 (N_660,N_210,N_387);
nor U661 (N_661,N_4,N_176);
or U662 (N_662,N_152,N_90);
or U663 (N_663,N_442,N_261);
nand U664 (N_664,N_79,N_293);
and U665 (N_665,N_29,N_186);
and U666 (N_666,N_424,N_285);
or U667 (N_667,N_222,N_295);
and U668 (N_668,N_465,N_1);
nand U669 (N_669,N_40,N_385);
and U670 (N_670,N_224,N_49);
xnor U671 (N_671,N_168,N_133);
or U672 (N_672,N_409,N_336);
or U673 (N_673,N_149,N_228);
nor U674 (N_674,N_248,N_198);
nor U675 (N_675,N_179,N_268);
nand U676 (N_676,N_7,N_423);
nor U677 (N_677,N_386,N_63);
and U678 (N_678,N_469,N_114);
nand U679 (N_679,N_100,N_401);
nand U680 (N_680,N_212,N_449);
or U681 (N_681,N_81,N_300);
nor U682 (N_682,N_363,N_489);
or U683 (N_683,N_12,N_77);
xnor U684 (N_684,N_463,N_143);
nand U685 (N_685,N_217,N_134);
nor U686 (N_686,N_204,N_426);
nand U687 (N_687,N_404,N_440);
xnor U688 (N_688,N_229,N_159);
or U689 (N_689,N_476,N_129);
or U690 (N_690,N_306,N_340);
xor U691 (N_691,N_422,N_339);
and U692 (N_692,N_368,N_255);
or U693 (N_693,N_35,N_57);
nor U694 (N_694,N_10,N_327);
and U695 (N_695,N_92,N_72);
nor U696 (N_696,N_65,N_16);
or U697 (N_697,N_359,N_292);
or U698 (N_698,N_334,N_258);
or U699 (N_699,N_398,N_320);
nand U700 (N_700,N_38,N_348);
and U701 (N_701,N_52,N_33);
and U702 (N_702,N_190,N_109);
or U703 (N_703,N_286,N_113);
or U704 (N_704,N_87,N_230);
nor U705 (N_705,N_303,N_281);
nor U706 (N_706,N_242,N_226);
nand U707 (N_707,N_346,N_125);
nand U708 (N_708,N_192,N_323);
xnor U709 (N_709,N_480,N_249);
and U710 (N_710,N_305,N_146);
or U711 (N_711,N_382,N_20);
and U712 (N_712,N_59,N_431);
nand U713 (N_713,N_421,N_47);
nor U714 (N_714,N_108,N_167);
or U715 (N_715,N_427,N_435);
nor U716 (N_716,N_373,N_46);
nand U717 (N_717,N_205,N_144);
nor U718 (N_718,N_23,N_304);
and U719 (N_719,N_477,N_395);
nand U720 (N_720,N_413,N_153);
nor U721 (N_721,N_392,N_18);
nand U722 (N_722,N_357,N_355);
and U723 (N_723,N_479,N_448);
or U724 (N_724,N_141,N_419);
and U725 (N_725,N_147,N_91);
or U726 (N_726,N_468,N_94);
or U727 (N_727,N_311,N_265);
nand U728 (N_728,N_460,N_164);
and U729 (N_729,N_411,N_393);
or U730 (N_730,N_120,N_243);
nor U731 (N_731,N_493,N_326);
nor U732 (N_732,N_54,N_214);
nand U733 (N_733,N_283,N_296);
and U734 (N_734,N_451,N_115);
nor U735 (N_735,N_128,N_378);
nand U736 (N_736,N_107,N_276);
and U737 (N_737,N_14,N_356);
nor U738 (N_738,N_470,N_22);
xnor U739 (N_739,N_220,N_472);
and U740 (N_740,N_221,N_103);
or U741 (N_741,N_130,N_277);
nor U742 (N_742,N_429,N_53);
or U743 (N_743,N_251,N_3);
or U744 (N_744,N_208,N_234);
nor U745 (N_745,N_195,N_238);
nand U746 (N_746,N_158,N_70);
nor U747 (N_747,N_194,N_148);
nor U748 (N_748,N_154,N_333);
nand U749 (N_749,N_180,N_191);
or U750 (N_750,N_360,N_324);
and U751 (N_751,N_419,N_10);
or U752 (N_752,N_368,N_124);
or U753 (N_753,N_7,N_338);
nand U754 (N_754,N_191,N_326);
and U755 (N_755,N_168,N_192);
nor U756 (N_756,N_76,N_160);
and U757 (N_757,N_343,N_53);
nor U758 (N_758,N_410,N_143);
and U759 (N_759,N_84,N_346);
nand U760 (N_760,N_483,N_498);
nor U761 (N_761,N_83,N_173);
nand U762 (N_762,N_186,N_121);
nand U763 (N_763,N_308,N_67);
nand U764 (N_764,N_486,N_91);
nor U765 (N_765,N_325,N_104);
nor U766 (N_766,N_312,N_433);
xnor U767 (N_767,N_12,N_346);
xnor U768 (N_768,N_165,N_3);
nand U769 (N_769,N_110,N_204);
and U770 (N_770,N_56,N_359);
and U771 (N_771,N_215,N_1);
nor U772 (N_772,N_289,N_347);
xnor U773 (N_773,N_338,N_480);
nor U774 (N_774,N_14,N_205);
and U775 (N_775,N_339,N_303);
xnor U776 (N_776,N_308,N_355);
and U777 (N_777,N_416,N_172);
and U778 (N_778,N_395,N_293);
and U779 (N_779,N_28,N_359);
xnor U780 (N_780,N_95,N_201);
nor U781 (N_781,N_311,N_143);
and U782 (N_782,N_311,N_9);
and U783 (N_783,N_214,N_180);
nor U784 (N_784,N_264,N_462);
xnor U785 (N_785,N_256,N_441);
nor U786 (N_786,N_101,N_146);
and U787 (N_787,N_0,N_134);
or U788 (N_788,N_285,N_389);
nor U789 (N_789,N_446,N_186);
and U790 (N_790,N_28,N_353);
nor U791 (N_791,N_313,N_66);
and U792 (N_792,N_17,N_255);
and U793 (N_793,N_273,N_238);
nand U794 (N_794,N_464,N_226);
nor U795 (N_795,N_31,N_274);
and U796 (N_796,N_120,N_15);
nor U797 (N_797,N_350,N_58);
or U798 (N_798,N_154,N_314);
nand U799 (N_799,N_316,N_229);
nor U800 (N_800,N_184,N_439);
nor U801 (N_801,N_98,N_187);
nand U802 (N_802,N_157,N_262);
and U803 (N_803,N_388,N_115);
or U804 (N_804,N_296,N_87);
nor U805 (N_805,N_127,N_404);
or U806 (N_806,N_251,N_68);
xor U807 (N_807,N_449,N_26);
and U808 (N_808,N_441,N_160);
or U809 (N_809,N_259,N_471);
nand U810 (N_810,N_161,N_186);
nor U811 (N_811,N_453,N_307);
nor U812 (N_812,N_223,N_134);
or U813 (N_813,N_339,N_35);
nand U814 (N_814,N_99,N_212);
nand U815 (N_815,N_222,N_186);
nor U816 (N_816,N_105,N_471);
nor U817 (N_817,N_81,N_464);
or U818 (N_818,N_389,N_430);
nand U819 (N_819,N_186,N_192);
and U820 (N_820,N_332,N_344);
nor U821 (N_821,N_32,N_252);
or U822 (N_822,N_219,N_432);
or U823 (N_823,N_339,N_215);
nor U824 (N_824,N_223,N_345);
nor U825 (N_825,N_227,N_158);
and U826 (N_826,N_371,N_71);
xnor U827 (N_827,N_385,N_291);
nand U828 (N_828,N_291,N_380);
and U829 (N_829,N_134,N_236);
and U830 (N_830,N_297,N_25);
nand U831 (N_831,N_215,N_295);
and U832 (N_832,N_352,N_405);
and U833 (N_833,N_454,N_80);
xor U834 (N_834,N_428,N_464);
or U835 (N_835,N_470,N_109);
xnor U836 (N_836,N_413,N_343);
nand U837 (N_837,N_281,N_227);
nand U838 (N_838,N_326,N_170);
or U839 (N_839,N_233,N_9);
and U840 (N_840,N_401,N_63);
nand U841 (N_841,N_116,N_43);
nor U842 (N_842,N_107,N_492);
or U843 (N_843,N_288,N_331);
nor U844 (N_844,N_273,N_481);
nand U845 (N_845,N_9,N_351);
and U846 (N_846,N_108,N_260);
nand U847 (N_847,N_186,N_204);
and U848 (N_848,N_202,N_231);
and U849 (N_849,N_363,N_59);
nor U850 (N_850,N_442,N_174);
nand U851 (N_851,N_239,N_124);
or U852 (N_852,N_128,N_167);
nor U853 (N_853,N_388,N_175);
or U854 (N_854,N_25,N_308);
nor U855 (N_855,N_437,N_53);
and U856 (N_856,N_368,N_35);
nor U857 (N_857,N_198,N_50);
or U858 (N_858,N_493,N_55);
and U859 (N_859,N_247,N_22);
xor U860 (N_860,N_474,N_173);
and U861 (N_861,N_101,N_248);
or U862 (N_862,N_211,N_4);
nor U863 (N_863,N_114,N_124);
nor U864 (N_864,N_211,N_13);
xor U865 (N_865,N_250,N_246);
nor U866 (N_866,N_237,N_69);
and U867 (N_867,N_381,N_170);
nand U868 (N_868,N_192,N_182);
nand U869 (N_869,N_319,N_214);
and U870 (N_870,N_372,N_98);
nand U871 (N_871,N_493,N_367);
nor U872 (N_872,N_14,N_266);
nor U873 (N_873,N_407,N_466);
nand U874 (N_874,N_460,N_371);
nand U875 (N_875,N_352,N_233);
xor U876 (N_876,N_91,N_152);
nor U877 (N_877,N_194,N_387);
or U878 (N_878,N_499,N_74);
nand U879 (N_879,N_174,N_337);
nor U880 (N_880,N_135,N_220);
or U881 (N_881,N_375,N_417);
nor U882 (N_882,N_263,N_338);
nand U883 (N_883,N_242,N_165);
or U884 (N_884,N_248,N_481);
nand U885 (N_885,N_194,N_417);
and U886 (N_886,N_420,N_57);
nor U887 (N_887,N_338,N_114);
nand U888 (N_888,N_371,N_343);
nand U889 (N_889,N_368,N_20);
nand U890 (N_890,N_457,N_11);
and U891 (N_891,N_155,N_445);
and U892 (N_892,N_407,N_244);
nand U893 (N_893,N_467,N_140);
and U894 (N_894,N_254,N_466);
nor U895 (N_895,N_397,N_84);
or U896 (N_896,N_6,N_326);
xor U897 (N_897,N_388,N_136);
or U898 (N_898,N_497,N_170);
or U899 (N_899,N_68,N_481);
nor U900 (N_900,N_456,N_219);
and U901 (N_901,N_238,N_70);
or U902 (N_902,N_90,N_325);
or U903 (N_903,N_112,N_6);
nand U904 (N_904,N_153,N_377);
nor U905 (N_905,N_414,N_476);
or U906 (N_906,N_73,N_390);
and U907 (N_907,N_458,N_411);
and U908 (N_908,N_369,N_155);
nand U909 (N_909,N_433,N_17);
and U910 (N_910,N_233,N_52);
and U911 (N_911,N_132,N_51);
nor U912 (N_912,N_120,N_402);
and U913 (N_913,N_99,N_35);
and U914 (N_914,N_450,N_154);
nand U915 (N_915,N_155,N_133);
or U916 (N_916,N_424,N_312);
nand U917 (N_917,N_444,N_411);
and U918 (N_918,N_459,N_270);
nor U919 (N_919,N_144,N_150);
nand U920 (N_920,N_162,N_276);
nand U921 (N_921,N_62,N_465);
nor U922 (N_922,N_428,N_159);
or U923 (N_923,N_339,N_24);
nand U924 (N_924,N_421,N_147);
or U925 (N_925,N_107,N_40);
and U926 (N_926,N_175,N_262);
xor U927 (N_927,N_45,N_375);
nand U928 (N_928,N_162,N_16);
xnor U929 (N_929,N_261,N_343);
xnor U930 (N_930,N_317,N_238);
xnor U931 (N_931,N_464,N_265);
nor U932 (N_932,N_477,N_119);
xnor U933 (N_933,N_204,N_207);
nand U934 (N_934,N_232,N_274);
xor U935 (N_935,N_151,N_128);
and U936 (N_936,N_344,N_305);
nor U937 (N_937,N_92,N_269);
nor U938 (N_938,N_142,N_252);
nor U939 (N_939,N_393,N_409);
and U940 (N_940,N_165,N_325);
nor U941 (N_941,N_462,N_374);
or U942 (N_942,N_116,N_149);
or U943 (N_943,N_232,N_496);
nor U944 (N_944,N_387,N_67);
nand U945 (N_945,N_90,N_8);
nand U946 (N_946,N_399,N_26);
or U947 (N_947,N_201,N_480);
nor U948 (N_948,N_214,N_20);
and U949 (N_949,N_318,N_325);
and U950 (N_950,N_25,N_131);
and U951 (N_951,N_61,N_68);
and U952 (N_952,N_336,N_230);
nor U953 (N_953,N_203,N_327);
nor U954 (N_954,N_38,N_252);
or U955 (N_955,N_106,N_492);
nand U956 (N_956,N_219,N_244);
nor U957 (N_957,N_282,N_359);
and U958 (N_958,N_24,N_374);
nor U959 (N_959,N_17,N_60);
or U960 (N_960,N_464,N_287);
nand U961 (N_961,N_182,N_457);
and U962 (N_962,N_401,N_392);
xnor U963 (N_963,N_450,N_454);
nor U964 (N_964,N_425,N_488);
and U965 (N_965,N_129,N_189);
nor U966 (N_966,N_40,N_421);
xnor U967 (N_967,N_138,N_123);
nand U968 (N_968,N_414,N_176);
or U969 (N_969,N_204,N_162);
or U970 (N_970,N_254,N_165);
nor U971 (N_971,N_143,N_394);
and U972 (N_972,N_493,N_243);
or U973 (N_973,N_415,N_81);
and U974 (N_974,N_339,N_220);
nand U975 (N_975,N_287,N_271);
nor U976 (N_976,N_460,N_167);
and U977 (N_977,N_151,N_110);
nor U978 (N_978,N_441,N_410);
nand U979 (N_979,N_224,N_8);
or U980 (N_980,N_204,N_433);
or U981 (N_981,N_50,N_197);
or U982 (N_982,N_320,N_334);
and U983 (N_983,N_311,N_281);
nand U984 (N_984,N_57,N_479);
nor U985 (N_985,N_480,N_361);
and U986 (N_986,N_128,N_426);
or U987 (N_987,N_325,N_317);
and U988 (N_988,N_343,N_403);
nand U989 (N_989,N_390,N_234);
nor U990 (N_990,N_383,N_401);
and U991 (N_991,N_285,N_321);
nor U992 (N_992,N_419,N_153);
or U993 (N_993,N_334,N_34);
nand U994 (N_994,N_450,N_169);
or U995 (N_995,N_373,N_405);
and U996 (N_996,N_131,N_290);
nand U997 (N_997,N_65,N_393);
and U998 (N_998,N_465,N_71);
nand U999 (N_999,N_131,N_320);
xor U1000 (N_1000,N_782,N_603);
nor U1001 (N_1001,N_607,N_592);
xnor U1002 (N_1002,N_569,N_641);
and U1003 (N_1003,N_565,N_899);
nand U1004 (N_1004,N_862,N_551);
or U1005 (N_1005,N_923,N_710);
and U1006 (N_1006,N_672,N_647);
nor U1007 (N_1007,N_785,N_549);
xnor U1008 (N_1008,N_902,N_998);
nor U1009 (N_1009,N_858,N_534);
and U1010 (N_1010,N_810,N_738);
nand U1011 (N_1011,N_966,N_704);
and U1012 (N_1012,N_925,N_876);
or U1013 (N_1013,N_915,N_552);
or U1014 (N_1014,N_624,N_794);
nor U1015 (N_1015,N_575,N_954);
or U1016 (N_1016,N_522,N_508);
nand U1017 (N_1017,N_851,N_669);
or U1018 (N_1018,N_930,N_586);
or U1019 (N_1019,N_688,N_613);
nand U1020 (N_1020,N_676,N_608);
or U1021 (N_1021,N_744,N_511);
nor U1022 (N_1022,N_690,N_536);
nand U1023 (N_1023,N_970,N_720);
nor U1024 (N_1024,N_681,N_708);
xnor U1025 (N_1025,N_771,N_519);
nor U1026 (N_1026,N_849,N_543);
nand U1027 (N_1027,N_820,N_894);
nand U1028 (N_1028,N_531,N_699);
nor U1029 (N_1029,N_996,N_868);
nand U1030 (N_1030,N_595,N_878);
and U1031 (N_1031,N_957,N_756);
or U1032 (N_1032,N_788,N_593);
xnor U1033 (N_1033,N_614,N_768);
nand U1034 (N_1034,N_793,N_917);
nand U1035 (N_1035,N_634,N_955);
nand U1036 (N_1036,N_757,N_786);
nor U1037 (N_1037,N_646,N_594);
or U1038 (N_1038,N_906,N_942);
and U1039 (N_1039,N_843,N_617);
nor U1040 (N_1040,N_960,N_752);
nor U1041 (N_1041,N_736,N_643);
xnor U1042 (N_1042,N_733,N_597);
or U1043 (N_1043,N_784,N_914);
or U1044 (N_1044,N_589,N_761);
nand U1045 (N_1045,N_512,N_934);
nand U1046 (N_1046,N_611,N_668);
and U1047 (N_1047,N_740,N_840);
xor U1048 (N_1048,N_973,N_988);
and U1049 (N_1049,N_572,N_537);
nor U1050 (N_1050,N_836,N_627);
nand U1051 (N_1051,N_853,N_968);
and U1052 (N_1052,N_556,N_891);
nor U1053 (N_1053,N_936,N_818);
and U1054 (N_1054,N_879,N_922);
nand U1055 (N_1055,N_947,N_583);
and U1056 (N_1056,N_510,N_839);
or U1057 (N_1057,N_666,N_846);
or U1058 (N_1058,N_650,N_596);
nor U1059 (N_1059,N_694,N_513);
nand U1060 (N_1060,N_854,N_711);
and U1061 (N_1061,N_911,N_610);
and U1062 (N_1062,N_961,N_566);
nor U1063 (N_1063,N_605,N_937);
or U1064 (N_1064,N_619,N_680);
nor U1065 (N_1065,N_926,N_848);
nand U1066 (N_1066,N_944,N_815);
nor U1067 (N_1067,N_726,N_745);
and U1068 (N_1068,N_995,N_775);
and U1069 (N_1069,N_640,N_866);
xnor U1070 (N_1070,N_938,N_573);
and U1071 (N_1071,N_832,N_692);
nand U1072 (N_1072,N_719,N_675);
or U1073 (N_1073,N_554,N_861);
nor U1074 (N_1074,N_819,N_587);
xor U1075 (N_1075,N_691,N_792);
and U1076 (N_1076,N_881,N_992);
nand U1077 (N_1077,N_791,N_816);
nor U1078 (N_1078,N_542,N_863);
and U1079 (N_1079,N_813,N_558);
or U1080 (N_1080,N_932,N_956);
nand U1081 (N_1081,N_600,N_939);
and U1082 (N_1082,N_940,N_781);
nand U1083 (N_1083,N_532,N_564);
or U1084 (N_1084,N_576,N_987);
nand U1085 (N_1085,N_571,N_770);
or U1086 (N_1086,N_799,N_567);
nand U1087 (N_1087,N_503,N_637);
nand U1088 (N_1088,N_997,N_869);
and U1089 (N_1089,N_527,N_821);
nor U1090 (N_1090,N_974,N_741);
nand U1091 (N_1091,N_962,N_682);
or U1092 (N_1092,N_707,N_765);
nand U1093 (N_1093,N_981,N_528);
and U1094 (N_1094,N_787,N_951);
and U1095 (N_1095,N_919,N_578);
nand U1096 (N_1096,N_969,N_999);
and U1097 (N_1097,N_604,N_993);
or U1098 (N_1098,N_671,N_662);
nand U1099 (N_1099,N_850,N_764);
nor U1100 (N_1100,N_859,N_830);
or U1101 (N_1101,N_801,N_725);
and U1102 (N_1102,N_609,N_827);
xor U1103 (N_1103,N_721,N_847);
or U1104 (N_1104,N_615,N_817);
nor U1105 (N_1105,N_501,N_822);
nand U1106 (N_1106,N_941,N_958);
or U1107 (N_1107,N_730,N_831);
and U1108 (N_1108,N_865,N_842);
and U1109 (N_1109,N_644,N_718);
and U1110 (N_1110,N_625,N_742);
and U1111 (N_1111,N_724,N_588);
or U1112 (N_1112,N_901,N_985);
nor U1113 (N_1113,N_673,N_714);
nor U1114 (N_1114,N_860,N_826);
or U1115 (N_1115,N_766,N_874);
nor U1116 (N_1116,N_715,N_706);
or U1117 (N_1117,N_963,N_924);
nor U1118 (N_1118,N_645,N_778);
and U1119 (N_1119,N_758,N_780);
and U1120 (N_1120,N_547,N_540);
nand U1121 (N_1121,N_553,N_748);
or U1122 (N_1122,N_984,N_732);
and U1123 (N_1123,N_774,N_702);
and U1124 (N_1124,N_579,N_812);
nor U1125 (N_1125,N_628,N_716);
nand U1126 (N_1126,N_769,N_632);
nand U1127 (N_1127,N_977,N_754);
xnor U1128 (N_1128,N_762,N_802);
nor U1129 (N_1129,N_870,N_703);
nand U1130 (N_1130,N_638,N_897);
nand U1131 (N_1131,N_909,N_872);
and U1132 (N_1132,N_633,N_560);
and U1133 (N_1133,N_943,N_877);
and U1134 (N_1134,N_529,N_882);
and U1135 (N_1135,N_746,N_570);
nor U1136 (N_1136,N_642,N_502);
xor U1137 (N_1137,N_743,N_777);
xor U1138 (N_1138,N_798,N_946);
nor U1139 (N_1139,N_857,N_991);
or U1140 (N_1140,N_838,N_659);
nand U1141 (N_1141,N_809,N_749);
or U1142 (N_1142,N_581,N_636);
nand U1143 (N_1143,N_539,N_965);
nor U1144 (N_1144,N_953,N_760);
or U1145 (N_1145,N_883,N_735);
nand U1146 (N_1146,N_773,N_591);
nor U1147 (N_1147,N_750,N_871);
xor U1148 (N_1148,N_814,N_731);
xnor U1149 (N_1149,N_892,N_982);
nand U1150 (N_1150,N_555,N_697);
xor U1151 (N_1151,N_712,N_795);
xnor U1152 (N_1152,N_907,N_890);
nand U1153 (N_1153,N_855,N_622);
or U1154 (N_1154,N_945,N_705);
and U1155 (N_1155,N_626,N_606);
and U1156 (N_1156,N_967,N_811);
nor U1157 (N_1157,N_538,N_563);
or U1158 (N_1158,N_885,N_927);
nor U1159 (N_1159,N_964,N_709);
and U1160 (N_1160,N_678,N_664);
nor U1161 (N_1161,N_582,N_790);
nand U1162 (N_1162,N_621,N_654);
nand U1163 (N_1163,N_796,N_727);
nand U1164 (N_1164,N_935,N_845);
nor U1165 (N_1165,N_910,N_700);
and U1166 (N_1166,N_931,N_722);
or U1167 (N_1167,N_535,N_808);
and U1168 (N_1168,N_844,N_693);
and U1169 (N_1169,N_823,N_585);
and U1170 (N_1170,N_524,N_701);
or U1171 (N_1171,N_639,N_518);
or U1172 (N_1172,N_677,N_759);
and U1173 (N_1173,N_747,N_873);
nor U1174 (N_1174,N_841,N_889);
or U1175 (N_1175,N_978,N_805);
or U1176 (N_1176,N_602,N_667);
nor U1177 (N_1177,N_959,N_695);
nand U1178 (N_1178,N_887,N_949);
or U1179 (N_1179,N_504,N_599);
nand U1180 (N_1180,N_806,N_783);
xnor U1181 (N_1181,N_975,N_655);
nor U1182 (N_1182,N_651,N_656);
nor U1183 (N_1183,N_545,N_729);
nor U1184 (N_1184,N_837,N_896);
nand U1185 (N_1185,N_689,N_568);
or U1186 (N_1186,N_686,N_620);
or U1187 (N_1187,N_674,N_685);
and U1188 (N_1188,N_653,N_557);
or U1189 (N_1189,N_665,N_928);
or U1190 (N_1190,N_630,N_629);
and U1191 (N_1191,N_514,N_893);
nor U1192 (N_1192,N_880,N_670);
and U1193 (N_1193,N_864,N_601);
nand U1194 (N_1194,N_976,N_526);
or U1195 (N_1195,N_523,N_753);
and U1196 (N_1196,N_520,N_658);
nor U1197 (N_1197,N_663,N_679);
nor U1198 (N_1198,N_807,N_833);
xnor U1199 (N_1199,N_717,N_980);
xnor U1200 (N_1200,N_590,N_972);
xnor U1201 (N_1201,N_660,N_776);
or U1202 (N_1202,N_723,N_828);
or U1203 (N_1203,N_867,N_612);
nor U1204 (N_1204,N_971,N_929);
xnor U1205 (N_1205,N_875,N_835);
or U1206 (N_1206,N_506,N_886);
nor U1207 (N_1207,N_541,N_900);
or U1208 (N_1208,N_755,N_684);
or U1209 (N_1209,N_921,N_580);
or U1210 (N_1210,N_661,N_562);
xor U1211 (N_1211,N_948,N_584);
nor U1212 (N_1212,N_623,N_898);
nor U1213 (N_1213,N_912,N_505);
and U1214 (N_1214,N_525,N_648);
and U1215 (N_1215,N_561,N_544);
nor U1216 (N_1216,N_616,N_574);
or U1217 (N_1217,N_952,N_933);
nor U1218 (N_1218,N_635,N_803);
and U1219 (N_1219,N_950,N_546);
nor U1220 (N_1220,N_918,N_804);
and U1221 (N_1221,N_983,N_905);
and U1222 (N_1222,N_657,N_989);
xnor U1223 (N_1223,N_533,N_517);
and U1224 (N_1224,N_767,N_908);
xnor U1225 (N_1225,N_739,N_500);
nand U1226 (N_1226,N_631,N_884);
nand U1227 (N_1227,N_913,N_728);
and U1228 (N_1228,N_903,N_696);
nor U1229 (N_1229,N_530,N_904);
nand U1230 (N_1230,N_687,N_772);
nand U1231 (N_1231,N_797,N_888);
nand U1232 (N_1232,N_652,N_800);
and U1233 (N_1233,N_751,N_829);
xor U1234 (N_1234,N_779,N_789);
or U1235 (N_1235,N_834,N_598);
nand U1236 (N_1236,N_550,N_515);
and U1237 (N_1237,N_734,N_763);
or U1238 (N_1238,N_856,N_559);
nor U1239 (N_1239,N_713,N_895);
or U1240 (N_1240,N_979,N_986);
and U1241 (N_1241,N_509,N_824);
xor U1242 (N_1242,N_548,N_649);
and U1243 (N_1243,N_990,N_994);
nor U1244 (N_1244,N_683,N_920);
and U1245 (N_1245,N_521,N_516);
nor U1246 (N_1246,N_737,N_618);
xnor U1247 (N_1247,N_507,N_852);
nand U1248 (N_1248,N_825,N_577);
or U1249 (N_1249,N_916,N_698);
nand U1250 (N_1250,N_500,N_512);
nor U1251 (N_1251,N_582,N_839);
nand U1252 (N_1252,N_995,N_920);
nand U1253 (N_1253,N_784,N_816);
and U1254 (N_1254,N_699,N_794);
or U1255 (N_1255,N_609,N_865);
nand U1256 (N_1256,N_815,N_600);
nand U1257 (N_1257,N_908,N_783);
and U1258 (N_1258,N_734,N_747);
nor U1259 (N_1259,N_911,N_632);
and U1260 (N_1260,N_814,N_884);
or U1261 (N_1261,N_712,N_967);
xnor U1262 (N_1262,N_622,N_991);
and U1263 (N_1263,N_947,N_529);
nand U1264 (N_1264,N_612,N_792);
nor U1265 (N_1265,N_743,N_926);
nand U1266 (N_1266,N_719,N_999);
or U1267 (N_1267,N_812,N_837);
or U1268 (N_1268,N_642,N_882);
nand U1269 (N_1269,N_658,N_592);
xor U1270 (N_1270,N_618,N_765);
and U1271 (N_1271,N_897,N_664);
and U1272 (N_1272,N_556,N_551);
and U1273 (N_1273,N_622,N_592);
and U1274 (N_1274,N_881,N_620);
nor U1275 (N_1275,N_826,N_861);
nand U1276 (N_1276,N_592,N_544);
and U1277 (N_1277,N_535,N_593);
nand U1278 (N_1278,N_862,N_613);
xnor U1279 (N_1279,N_552,N_555);
or U1280 (N_1280,N_882,N_872);
or U1281 (N_1281,N_538,N_571);
nand U1282 (N_1282,N_846,N_547);
nor U1283 (N_1283,N_669,N_728);
and U1284 (N_1284,N_729,N_787);
xnor U1285 (N_1285,N_534,N_518);
or U1286 (N_1286,N_674,N_502);
nor U1287 (N_1287,N_774,N_594);
and U1288 (N_1288,N_792,N_768);
and U1289 (N_1289,N_891,N_899);
nand U1290 (N_1290,N_689,N_899);
or U1291 (N_1291,N_577,N_699);
xor U1292 (N_1292,N_978,N_773);
or U1293 (N_1293,N_910,N_878);
or U1294 (N_1294,N_618,N_665);
or U1295 (N_1295,N_952,N_852);
or U1296 (N_1296,N_591,N_841);
and U1297 (N_1297,N_997,N_509);
nor U1298 (N_1298,N_858,N_920);
or U1299 (N_1299,N_798,N_869);
nand U1300 (N_1300,N_873,N_753);
nand U1301 (N_1301,N_719,N_607);
nand U1302 (N_1302,N_732,N_743);
nor U1303 (N_1303,N_876,N_549);
nor U1304 (N_1304,N_758,N_556);
nand U1305 (N_1305,N_839,N_561);
xor U1306 (N_1306,N_996,N_582);
or U1307 (N_1307,N_743,N_952);
xor U1308 (N_1308,N_557,N_815);
xnor U1309 (N_1309,N_874,N_795);
nand U1310 (N_1310,N_825,N_514);
or U1311 (N_1311,N_855,N_623);
or U1312 (N_1312,N_900,N_548);
or U1313 (N_1313,N_806,N_883);
nor U1314 (N_1314,N_918,N_791);
nor U1315 (N_1315,N_947,N_964);
nor U1316 (N_1316,N_579,N_520);
or U1317 (N_1317,N_825,N_918);
or U1318 (N_1318,N_951,N_821);
and U1319 (N_1319,N_983,N_752);
nor U1320 (N_1320,N_983,N_783);
nor U1321 (N_1321,N_558,N_632);
or U1322 (N_1322,N_698,N_577);
or U1323 (N_1323,N_611,N_871);
nor U1324 (N_1324,N_504,N_766);
nor U1325 (N_1325,N_766,N_945);
nor U1326 (N_1326,N_955,N_858);
or U1327 (N_1327,N_718,N_889);
nand U1328 (N_1328,N_520,N_583);
xnor U1329 (N_1329,N_781,N_645);
xnor U1330 (N_1330,N_736,N_550);
nor U1331 (N_1331,N_805,N_823);
nor U1332 (N_1332,N_744,N_630);
xnor U1333 (N_1333,N_755,N_829);
nand U1334 (N_1334,N_971,N_738);
and U1335 (N_1335,N_589,N_604);
nor U1336 (N_1336,N_973,N_845);
nand U1337 (N_1337,N_500,N_742);
or U1338 (N_1338,N_806,N_646);
or U1339 (N_1339,N_884,N_955);
nand U1340 (N_1340,N_658,N_949);
nand U1341 (N_1341,N_627,N_984);
nor U1342 (N_1342,N_724,N_682);
or U1343 (N_1343,N_580,N_941);
and U1344 (N_1344,N_706,N_640);
nand U1345 (N_1345,N_756,N_828);
or U1346 (N_1346,N_522,N_690);
nand U1347 (N_1347,N_617,N_853);
or U1348 (N_1348,N_828,N_821);
and U1349 (N_1349,N_843,N_686);
nor U1350 (N_1350,N_920,N_975);
and U1351 (N_1351,N_502,N_992);
or U1352 (N_1352,N_989,N_767);
and U1353 (N_1353,N_828,N_856);
or U1354 (N_1354,N_525,N_506);
or U1355 (N_1355,N_651,N_762);
nor U1356 (N_1356,N_886,N_745);
or U1357 (N_1357,N_552,N_583);
xor U1358 (N_1358,N_504,N_605);
nand U1359 (N_1359,N_568,N_866);
or U1360 (N_1360,N_771,N_973);
and U1361 (N_1361,N_636,N_921);
or U1362 (N_1362,N_648,N_817);
nor U1363 (N_1363,N_760,N_946);
and U1364 (N_1364,N_757,N_892);
and U1365 (N_1365,N_707,N_577);
or U1366 (N_1366,N_715,N_900);
xnor U1367 (N_1367,N_712,N_528);
xnor U1368 (N_1368,N_600,N_590);
and U1369 (N_1369,N_808,N_720);
and U1370 (N_1370,N_910,N_516);
and U1371 (N_1371,N_641,N_943);
and U1372 (N_1372,N_651,N_862);
or U1373 (N_1373,N_547,N_530);
and U1374 (N_1374,N_665,N_921);
and U1375 (N_1375,N_781,N_987);
nand U1376 (N_1376,N_526,N_518);
and U1377 (N_1377,N_888,N_774);
nand U1378 (N_1378,N_784,N_765);
xor U1379 (N_1379,N_968,N_697);
and U1380 (N_1380,N_669,N_859);
nor U1381 (N_1381,N_522,N_882);
xnor U1382 (N_1382,N_603,N_980);
xor U1383 (N_1383,N_664,N_997);
xnor U1384 (N_1384,N_700,N_659);
or U1385 (N_1385,N_789,N_902);
nor U1386 (N_1386,N_923,N_648);
xor U1387 (N_1387,N_683,N_806);
and U1388 (N_1388,N_632,N_677);
nor U1389 (N_1389,N_530,N_855);
and U1390 (N_1390,N_738,N_696);
nor U1391 (N_1391,N_605,N_916);
and U1392 (N_1392,N_890,N_896);
and U1393 (N_1393,N_828,N_937);
nor U1394 (N_1394,N_885,N_782);
nor U1395 (N_1395,N_956,N_860);
and U1396 (N_1396,N_597,N_688);
and U1397 (N_1397,N_839,N_806);
nor U1398 (N_1398,N_593,N_947);
nand U1399 (N_1399,N_904,N_700);
or U1400 (N_1400,N_791,N_539);
and U1401 (N_1401,N_675,N_539);
and U1402 (N_1402,N_845,N_936);
and U1403 (N_1403,N_689,N_720);
and U1404 (N_1404,N_775,N_561);
and U1405 (N_1405,N_525,N_799);
or U1406 (N_1406,N_517,N_914);
nand U1407 (N_1407,N_965,N_845);
or U1408 (N_1408,N_923,N_727);
or U1409 (N_1409,N_861,N_806);
and U1410 (N_1410,N_996,N_785);
nor U1411 (N_1411,N_965,N_881);
and U1412 (N_1412,N_788,N_507);
and U1413 (N_1413,N_701,N_587);
and U1414 (N_1414,N_904,N_814);
or U1415 (N_1415,N_842,N_639);
nand U1416 (N_1416,N_737,N_887);
and U1417 (N_1417,N_500,N_544);
or U1418 (N_1418,N_927,N_752);
nor U1419 (N_1419,N_686,N_772);
and U1420 (N_1420,N_575,N_576);
nor U1421 (N_1421,N_865,N_778);
and U1422 (N_1422,N_747,N_764);
or U1423 (N_1423,N_639,N_649);
nand U1424 (N_1424,N_564,N_953);
or U1425 (N_1425,N_901,N_995);
nand U1426 (N_1426,N_769,N_573);
xor U1427 (N_1427,N_775,N_911);
or U1428 (N_1428,N_519,N_825);
nand U1429 (N_1429,N_965,N_517);
nor U1430 (N_1430,N_808,N_687);
or U1431 (N_1431,N_587,N_785);
xor U1432 (N_1432,N_565,N_983);
nor U1433 (N_1433,N_675,N_784);
or U1434 (N_1434,N_996,N_641);
and U1435 (N_1435,N_629,N_568);
nand U1436 (N_1436,N_510,N_838);
nand U1437 (N_1437,N_612,N_577);
nand U1438 (N_1438,N_677,N_642);
and U1439 (N_1439,N_983,N_540);
or U1440 (N_1440,N_894,N_717);
and U1441 (N_1441,N_982,N_539);
or U1442 (N_1442,N_880,N_825);
and U1443 (N_1443,N_695,N_803);
and U1444 (N_1444,N_607,N_879);
and U1445 (N_1445,N_813,N_979);
xnor U1446 (N_1446,N_650,N_692);
and U1447 (N_1447,N_889,N_918);
or U1448 (N_1448,N_660,N_764);
nand U1449 (N_1449,N_740,N_658);
or U1450 (N_1450,N_528,N_975);
or U1451 (N_1451,N_590,N_887);
and U1452 (N_1452,N_991,N_861);
or U1453 (N_1453,N_984,N_639);
nor U1454 (N_1454,N_661,N_615);
nand U1455 (N_1455,N_609,N_888);
and U1456 (N_1456,N_776,N_741);
nand U1457 (N_1457,N_525,N_902);
xnor U1458 (N_1458,N_771,N_763);
nor U1459 (N_1459,N_710,N_890);
nand U1460 (N_1460,N_960,N_906);
and U1461 (N_1461,N_648,N_694);
and U1462 (N_1462,N_586,N_987);
and U1463 (N_1463,N_675,N_947);
nand U1464 (N_1464,N_929,N_878);
xor U1465 (N_1465,N_999,N_640);
nand U1466 (N_1466,N_525,N_560);
and U1467 (N_1467,N_981,N_594);
or U1468 (N_1468,N_924,N_680);
nand U1469 (N_1469,N_711,N_916);
nor U1470 (N_1470,N_646,N_657);
or U1471 (N_1471,N_939,N_615);
or U1472 (N_1472,N_546,N_843);
nor U1473 (N_1473,N_548,N_518);
nand U1474 (N_1474,N_867,N_917);
and U1475 (N_1475,N_561,N_548);
nand U1476 (N_1476,N_862,N_640);
nand U1477 (N_1477,N_839,N_709);
or U1478 (N_1478,N_951,N_902);
nor U1479 (N_1479,N_937,N_598);
nand U1480 (N_1480,N_696,N_665);
xnor U1481 (N_1481,N_830,N_908);
and U1482 (N_1482,N_590,N_896);
and U1483 (N_1483,N_801,N_712);
nor U1484 (N_1484,N_960,N_972);
nand U1485 (N_1485,N_532,N_886);
nor U1486 (N_1486,N_570,N_738);
or U1487 (N_1487,N_948,N_612);
nand U1488 (N_1488,N_503,N_906);
xnor U1489 (N_1489,N_785,N_579);
nor U1490 (N_1490,N_825,N_898);
nor U1491 (N_1491,N_706,N_525);
nand U1492 (N_1492,N_978,N_743);
xnor U1493 (N_1493,N_533,N_529);
or U1494 (N_1494,N_895,N_944);
nand U1495 (N_1495,N_796,N_754);
or U1496 (N_1496,N_952,N_867);
nand U1497 (N_1497,N_662,N_841);
nand U1498 (N_1498,N_926,N_987);
and U1499 (N_1499,N_639,N_837);
xnor U1500 (N_1500,N_1229,N_1162);
xnor U1501 (N_1501,N_1013,N_1409);
nand U1502 (N_1502,N_1116,N_1087);
xnor U1503 (N_1503,N_1475,N_1105);
or U1504 (N_1504,N_1053,N_1244);
nand U1505 (N_1505,N_1073,N_1478);
and U1506 (N_1506,N_1450,N_1084);
or U1507 (N_1507,N_1265,N_1052);
and U1508 (N_1508,N_1060,N_1304);
or U1509 (N_1509,N_1237,N_1173);
and U1510 (N_1510,N_1449,N_1120);
nor U1511 (N_1511,N_1169,N_1280);
or U1512 (N_1512,N_1296,N_1201);
or U1513 (N_1513,N_1352,N_1108);
or U1514 (N_1514,N_1054,N_1042);
nor U1515 (N_1515,N_1467,N_1132);
or U1516 (N_1516,N_1358,N_1341);
or U1517 (N_1517,N_1092,N_1091);
nor U1518 (N_1518,N_1401,N_1428);
nor U1519 (N_1519,N_1447,N_1346);
and U1520 (N_1520,N_1196,N_1065);
or U1521 (N_1521,N_1184,N_1493);
or U1522 (N_1522,N_1488,N_1474);
or U1523 (N_1523,N_1141,N_1461);
and U1524 (N_1524,N_1000,N_1363);
nand U1525 (N_1525,N_1494,N_1119);
nor U1526 (N_1526,N_1165,N_1199);
nand U1527 (N_1527,N_1011,N_1345);
nor U1528 (N_1528,N_1282,N_1067);
and U1529 (N_1529,N_1342,N_1330);
nor U1530 (N_1530,N_1144,N_1395);
nand U1531 (N_1531,N_1278,N_1227);
nor U1532 (N_1532,N_1321,N_1313);
and U1533 (N_1533,N_1223,N_1406);
nor U1534 (N_1534,N_1248,N_1232);
xnor U1535 (N_1535,N_1347,N_1125);
nor U1536 (N_1536,N_1460,N_1369);
or U1537 (N_1537,N_1365,N_1020);
and U1538 (N_1538,N_1463,N_1036);
nand U1539 (N_1539,N_1202,N_1040);
or U1540 (N_1540,N_1079,N_1086);
xnor U1541 (N_1541,N_1301,N_1076);
or U1542 (N_1542,N_1294,N_1031);
nor U1543 (N_1543,N_1207,N_1016);
and U1544 (N_1544,N_1286,N_1009);
and U1545 (N_1545,N_1057,N_1033);
and U1546 (N_1546,N_1214,N_1434);
nand U1547 (N_1547,N_1143,N_1012);
nor U1548 (N_1548,N_1063,N_1135);
nor U1549 (N_1549,N_1285,N_1198);
nand U1550 (N_1550,N_1161,N_1027);
xnor U1551 (N_1551,N_1459,N_1112);
or U1552 (N_1552,N_1274,N_1097);
or U1553 (N_1553,N_1268,N_1062);
and U1554 (N_1554,N_1149,N_1350);
and U1555 (N_1555,N_1385,N_1208);
or U1556 (N_1556,N_1457,N_1001);
nand U1557 (N_1557,N_1411,N_1498);
and U1558 (N_1558,N_1128,N_1005);
xor U1559 (N_1559,N_1150,N_1239);
xor U1560 (N_1560,N_1405,N_1080);
or U1561 (N_1561,N_1364,N_1098);
nor U1562 (N_1562,N_1034,N_1465);
nor U1563 (N_1563,N_1427,N_1083);
nor U1564 (N_1564,N_1025,N_1315);
and U1565 (N_1565,N_1370,N_1006);
nor U1566 (N_1566,N_1075,N_1220);
nor U1567 (N_1567,N_1295,N_1261);
nand U1568 (N_1568,N_1212,N_1407);
xor U1569 (N_1569,N_1327,N_1418);
nand U1570 (N_1570,N_1382,N_1240);
nor U1571 (N_1571,N_1417,N_1320);
and U1572 (N_1572,N_1335,N_1308);
or U1573 (N_1573,N_1045,N_1484);
nand U1574 (N_1574,N_1311,N_1048);
nand U1575 (N_1575,N_1292,N_1100);
or U1576 (N_1576,N_1153,N_1439);
xor U1577 (N_1577,N_1118,N_1166);
nand U1578 (N_1578,N_1030,N_1233);
or U1579 (N_1579,N_1179,N_1022);
or U1580 (N_1580,N_1154,N_1453);
or U1581 (N_1581,N_1130,N_1055);
or U1582 (N_1582,N_1398,N_1302);
or U1583 (N_1583,N_1152,N_1124);
and U1584 (N_1584,N_1164,N_1456);
and U1585 (N_1585,N_1413,N_1410);
nand U1586 (N_1586,N_1049,N_1200);
nor U1587 (N_1587,N_1085,N_1307);
and U1588 (N_1588,N_1272,N_1387);
and U1589 (N_1589,N_1367,N_1026);
nand U1590 (N_1590,N_1397,N_1176);
nand U1591 (N_1591,N_1246,N_1037);
or U1592 (N_1592,N_1021,N_1414);
nand U1593 (N_1593,N_1117,N_1051);
and U1594 (N_1594,N_1189,N_1448);
nand U1595 (N_1595,N_1127,N_1454);
or U1596 (N_1596,N_1114,N_1276);
and U1597 (N_1597,N_1354,N_1412);
or U1598 (N_1598,N_1194,N_1077);
nor U1599 (N_1599,N_1394,N_1258);
or U1600 (N_1600,N_1247,N_1485);
nand U1601 (N_1601,N_1462,N_1355);
and U1602 (N_1602,N_1445,N_1167);
nor U1603 (N_1603,N_1297,N_1018);
and U1604 (N_1604,N_1017,N_1305);
nand U1605 (N_1605,N_1446,N_1174);
and U1606 (N_1606,N_1339,N_1441);
nor U1607 (N_1607,N_1259,N_1241);
or U1608 (N_1608,N_1181,N_1101);
nor U1609 (N_1609,N_1211,N_1066);
or U1610 (N_1610,N_1380,N_1238);
nand U1611 (N_1611,N_1203,N_1400);
or U1612 (N_1612,N_1050,N_1163);
and U1613 (N_1613,N_1134,N_1399);
nor U1614 (N_1614,N_1175,N_1234);
nor U1615 (N_1615,N_1477,N_1300);
nand U1616 (N_1616,N_1222,N_1046);
and U1617 (N_1617,N_1186,N_1288);
and U1618 (N_1618,N_1182,N_1497);
nand U1619 (N_1619,N_1357,N_1047);
nand U1620 (N_1620,N_1298,N_1333);
nor U1621 (N_1621,N_1121,N_1329);
nor U1622 (N_1622,N_1170,N_1337);
or U1623 (N_1623,N_1139,N_1059);
nor U1624 (N_1624,N_1471,N_1479);
or U1625 (N_1625,N_1317,N_1205);
or U1626 (N_1626,N_1383,N_1002);
or U1627 (N_1627,N_1469,N_1245);
nand U1628 (N_1628,N_1064,N_1160);
or U1629 (N_1629,N_1483,N_1415);
nor U1630 (N_1630,N_1291,N_1224);
nand U1631 (N_1631,N_1041,N_1322);
xnor U1632 (N_1632,N_1107,N_1133);
nand U1633 (N_1633,N_1420,N_1111);
or U1634 (N_1634,N_1072,N_1255);
nor U1635 (N_1635,N_1221,N_1391);
or U1636 (N_1636,N_1374,N_1390);
nand U1637 (N_1637,N_1325,N_1422);
or U1638 (N_1638,N_1106,N_1217);
and U1639 (N_1639,N_1159,N_1252);
and U1640 (N_1640,N_1392,N_1470);
or U1641 (N_1641,N_1340,N_1056);
or U1642 (N_1642,N_1148,N_1082);
nor U1643 (N_1643,N_1426,N_1254);
or U1644 (N_1644,N_1215,N_1180);
xnor U1645 (N_1645,N_1158,N_1023);
and U1646 (N_1646,N_1039,N_1429);
nor U1647 (N_1647,N_1318,N_1271);
nand U1648 (N_1648,N_1102,N_1081);
xnor U1649 (N_1649,N_1284,N_1416);
nand U1650 (N_1650,N_1396,N_1226);
nand U1651 (N_1651,N_1433,N_1142);
and U1652 (N_1652,N_1069,N_1206);
nand U1653 (N_1653,N_1210,N_1443);
nor U1654 (N_1654,N_1424,N_1126);
xor U1655 (N_1655,N_1480,N_1216);
and U1656 (N_1656,N_1468,N_1038);
and U1657 (N_1657,N_1110,N_1476);
xor U1658 (N_1658,N_1193,N_1492);
nand U1659 (N_1659,N_1129,N_1035);
and U1660 (N_1660,N_1310,N_1455);
and U1661 (N_1661,N_1344,N_1332);
or U1662 (N_1662,N_1156,N_1486);
nand U1663 (N_1663,N_1379,N_1338);
and U1664 (N_1664,N_1250,N_1178);
nand U1665 (N_1665,N_1495,N_1078);
nand U1666 (N_1666,N_1482,N_1168);
nor U1667 (N_1667,N_1464,N_1435);
nor U1668 (N_1668,N_1185,N_1360);
and U1669 (N_1669,N_1472,N_1151);
nand U1670 (N_1670,N_1138,N_1177);
nand U1671 (N_1671,N_1442,N_1436);
nor U1672 (N_1672,N_1172,N_1306);
and U1673 (N_1673,N_1458,N_1197);
nor U1674 (N_1674,N_1444,N_1438);
nor U1675 (N_1675,N_1096,N_1290);
nand U1676 (N_1676,N_1195,N_1171);
xnor U1677 (N_1677,N_1491,N_1191);
and U1678 (N_1678,N_1309,N_1334);
nor U1679 (N_1679,N_1499,N_1283);
and U1680 (N_1680,N_1312,N_1043);
and U1681 (N_1681,N_1068,N_1071);
and U1682 (N_1682,N_1366,N_1155);
nand U1683 (N_1683,N_1336,N_1235);
nor U1684 (N_1684,N_1109,N_1319);
nor U1685 (N_1685,N_1122,N_1188);
or U1686 (N_1686,N_1230,N_1281);
nand U1687 (N_1687,N_1431,N_1263);
xnor U1688 (N_1688,N_1377,N_1331);
xnor U1689 (N_1689,N_1279,N_1218);
nand U1690 (N_1690,N_1376,N_1014);
nor U1691 (N_1691,N_1349,N_1253);
and U1692 (N_1692,N_1421,N_1289);
nor U1693 (N_1693,N_1440,N_1389);
or U1694 (N_1694,N_1113,N_1490);
xnor U1695 (N_1695,N_1147,N_1419);
nor U1696 (N_1696,N_1328,N_1140);
or U1697 (N_1697,N_1353,N_1007);
nand U1698 (N_1698,N_1003,N_1190);
nand U1699 (N_1699,N_1362,N_1095);
nor U1700 (N_1700,N_1044,N_1137);
nor U1701 (N_1701,N_1371,N_1204);
nor U1702 (N_1702,N_1004,N_1388);
nand U1703 (N_1703,N_1157,N_1381);
or U1704 (N_1704,N_1316,N_1242);
xnor U1705 (N_1705,N_1088,N_1326);
or U1706 (N_1706,N_1303,N_1032);
nor U1707 (N_1707,N_1093,N_1408);
nand U1708 (N_1708,N_1489,N_1277);
and U1709 (N_1709,N_1187,N_1267);
or U1710 (N_1710,N_1123,N_1131);
or U1711 (N_1711,N_1061,N_1008);
nand U1712 (N_1712,N_1090,N_1228);
nor U1713 (N_1713,N_1293,N_1314);
nor U1714 (N_1714,N_1099,N_1372);
and U1715 (N_1715,N_1386,N_1260);
or U1716 (N_1716,N_1145,N_1209);
or U1717 (N_1717,N_1299,N_1473);
nand U1718 (N_1718,N_1452,N_1146);
nor U1719 (N_1719,N_1324,N_1368);
and U1720 (N_1720,N_1231,N_1423);
nor U1721 (N_1721,N_1356,N_1430);
nand U1722 (N_1722,N_1359,N_1010);
xor U1723 (N_1723,N_1264,N_1192);
or U1724 (N_1724,N_1466,N_1236);
nand U1725 (N_1725,N_1074,N_1273);
xor U1726 (N_1726,N_1058,N_1378);
or U1727 (N_1727,N_1115,N_1343);
and U1728 (N_1728,N_1251,N_1403);
nor U1729 (N_1729,N_1402,N_1425);
nand U1730 (N_1730,N_1219,N_1070);
nor U1731 (N_1731,N_1029,N_1269);
or U1732 (N_1732,N_1257,N_1351);
nand U1733 (N_1733,N_1270,N_1487);
nor U1734 (N_1734,N_1262,N_1104);
or U1735 (N_1735,N_1393,N_1103);
nand U1736 (N_1736,N_1432,N_1256);
nor U1737 (N_1737,N_1384,N_1015);
or U1738 (N_1738,N_1019,N_1266);
nand U1739 (N_1739,N_1249,N_1404);
and U1740 (N_1740,N_1348,N_1375);
nand U1741 (N_1741,N_1361,N_1437);
or U1742 (N_1742,N_1496,N_1243);
nor U1743 (N_1743,N_1287,N_1094);
xor U1744 (N_1744,N_1136,N_1373);
xor U1745 (N_1745,N_1183,N_1213);
or U1746 (N_1746,N_1275,N_1225);
nand U1747 (N_1747,N_1089,N_1028);
nand U1748 (N_1748,N_1481,N_1323);
nor U1749 (N_1749,N_1451,N_1024);
and U1750 (N_1750,N_1300,N_1417);
xnor U1751 (N_1751,N_1064,N_1438);
nor U1752 (N_1752,N_1122,N_1466);
and U1753 (N_1753,N_1202,N_1183);
nor U1754 (N_1754,N_1465,N_1296);
and U1755 (N_1755,N_1320,N_1189);
nor U1756 (N_1756,N_1192,N_1247);
nor U1757 (N_1757,N_1436,N_1045);
nor U1758 (N_1758,N_1421,N_1119);
nor U1759 (N_1759,N_1357,N_1368);
nand U1760 (N_1760,N_1186,N_1488);
nand U1761 (N_1761,N_1087,N_1341);
or U1762 (N_1762,N_1023,N_1141);
or U1763 (N_1763,N_1104,N_1453);
and U1764 (N_1764,N_1216,N_1292);
or U1765 (N_1765,N_1281,N_1452);
and U1766 (N_1766,N_1462,N_1384);
xor U1767 (N_1767,N_1323,N_1434);
nor U1768 (N_1768,N_1120,N_1456);
nand U1769 (N_1769,N_1197,N_1203);
nor U1770 (N_1770,N_1263,N_1284);
nand U1771 (N_1771,N_1279,N_1367);
nand U1772 (N_1772,N_1121,N_1479);
nand U1773 (N_1773,N_1457,N_1015);
nor U1774 (N_1774,N_1147,N_1385);
nand U1775 (N_1775,N_1061,N_1062);
or U1776 (N_1776,N_1278,N_1121);
and U1777 (N_1777,N_1222,N_1348);
xor U1778 (N_1778,N_1000,N_1405);
and U1779 (N_1779,N_1450,N_1159);
nand U1780 (N_1780,N_1201,N_1000);
xnor U1781 (N_1781,N_1006,N_1449);
xor U1782 (N_1782,N_1451,N_1432);
xnor U1783 (N_1783,N_1081,N_1044);
or U1784 (N_1784,N_1234,N_1367);
or U1785 (N_1785,N_1050,N_1494);
nand U1786 (N_1786,N_1121,N_1208);
or U1787 (N_1787,N_1312,N_1332);
nor U1788 (N_1788,N_1224,N_1106);
and U1789 (N_1789,N_1112,N_1056);
nor U1790 (N_1790,N_1224,N_1419);
and U1791 (N_1791,N_1416,N_1400);
or U1792 (N_1792,N_1170,N_1300);
xor U1793 (N_1793,N_1368,N_1214);
nor U1794 (N_1794,N_1338,N_1068);
or U1795 (N_1795,N_1323,N_1291);
nor U1796 (N_1796,N_1059,N_1126);
nand U1797 (N_1797,N_1036,N_1174);
and U1798 (N_1798,N_1349,N_1367);
and U1799 (N_1799,N_1334,N_1000);
and U1800 (N_1800,N_1061,N_1042);
or U1801 (N_1801,N_1155,N_1386);
and U1802 (N_1802,N_1206,N_1267);
nor U1803 (N_1803,N_1061,N_1133);
and U1804 (N_1804,N_1195,N_1188);
nand U1805 (N_1805,N_1305,N_1391);
and U1806 (N_1806,N_1449,N_1368);
or U1807 (N_1807,N_1327,N_1491);
nand U1808 (N_1808,N_1273,N_1423);
nor U1809 (N_1809,N_1110,N_1293);
and U1810 (N_1810,N_1153,N_1446);
nand U1811 (N_1811,N_1281,N_1282);
or U1812 (N_1812,N_1455,N_1079);
and U1813 (N_1813,N_1186,N_1277);
or U1814 (N_1814,N_1354,N_1486);
nor U1815 (N_1815,N_1142,N_1165);
or U1816 (N_1816,N_1330,N_1496);
nand U1817 (N_1817,N_1326,N_1073);
or U1818 (N_1818,N_1225,N_1304);
and U1819 (N_1819,N_1438,N_1197);
and U1820 (N_1820,N_1494,N_1459);
nor U1821 (N_1821,N_1137,N_1057);
xor U1822 (N_1822,N_1031,N_1420);
nand U1823 (N_1823,N_1232,N_1371);
or U1824 (N_1824,N_1043,N_1202);
nand U1825 (N_1825,N_1490,N_1117);
and U1826 (N_1826,N_1286,N_1362);
and U1827 (N_1827,N_1434,N_1178);
nand U1828 (N_1828,N_1450,N_1278);
and U1829 (N_1829,N_1144,N_1452);
nor U1830 (N_1830,N_1242,N_1213);
xnor U1831 (N_1831,N_1059,N_1311);
or U1832 (N_1832,N_1348,N_1457);
xnor U1833 (N_1833,N_1294,N_1386);
and U1834 (N_1834,N_1172,N_1260);
nor U1835 (N_1835,N_1003,N_1185);
or U1836 (N_1836,N_1226,N_1220);
xor U1837 (N_1837,N_1044,N_1388);
nor U1838 (N_1838,N_1011,N_1390);
and U1839 (N_1839,N_1044,N_1060);
or U1840 (N_1840,N_1343,N_1250);
or U1841 (N_1841,N_1100,N_1246);
or U1842 (N_1842,N_1495,N_1374);
or U1843 (N_1843,N_1235,N_1465);
or U1844 (N_1844,N_1326,N_1241);
nand U1845 (N_1845,N_1105,N_1103);
nor U1846 (N_1846,N_1295,N_1103);
and U1847 (N_1847,N_1357,N_1335);
and U1848 (N_1848,N_1318,N_1480);
nand U1849 (N_1849,N_1012,N_1099);
or U1850 (N_1850,N_1077,N_1026);
nor U1851 (N_1851,N_1142,N_1440);
nand U1852 (N_1852,N_1465,N_1383);
or U1853 (N_1853,N_1294,N_1044);
nand U1854 (N_1854,N_1068,N_1145);
and U1855 (N_1855,N_1315,N_1375);
or U1856 (N_1856,N_1102,N_1240);
nand U1857 (N_1857,N_1303,N_1265);
and U1858 (N_1858,N_1022,N_1199);
nor U1859 (N_1859,N_1456,N_1433);
nor U1860 (N_1860,N_1139,N_1321);
nor U1861 (N_1861,N_1308,N_1401);
nand U1862 (N_1862,N_1243,N_1104);
nand U1863 (N_1863,N_1438,N_1138);
or U1864 (N_1864,N_1051,N_1366);
and U1865 (N_1865,N_1358,N_1248);
xor U1866 (N_1866,N_1476,N_1032);
and U1867 (N_1867,N_1083,N_1123);
and U1868 (N_1868,N_1210,N_1188);
nor U1869 (N_1869,N_1114,N_1068);
or U1870 (N_1870,N_1357,N_1026);
xnor U1871 (N_1871,N_1253,N_1194);
and U1872 (N_1872,N_1383,N_1282);
and U1873 (N_1873,N_1239,N_1492);
xor U1874 (N_1874,N_1148,N_1135);
or U1875 (N_1875,N_1334,N_1492);
nor U1876 (N_1876,N_1202,N_1486);
or U1877 (N_1877,N_1130,N_1023);
or U1878 (N_1878,N_1337,N_1277);
or U1879 (N_1879,N_1423,N_1250);
nor U1880 (N_1880,N_1468,N_1153);
or U1881 (N_1881,N_1378,N_1103);
xnor U1882 (N_1882,N_1216,N_1347);
or U1883 (N_1883,N_1416,N_1164);
or U1884 (N_1884,N_1015,N_1233);
or U1885 (N_1885,N_1036,N_1128);
or U1886 (N_1886,N_1380,N_1349);
nand U1887 (N_1887,N_1423,N_1006);
nor U1888 (N_1888,N_1101,N_1068);
nor U1889 (N_1889,N_1033,N_1367);
or U1890 (N_1890,N_1382,N_1163);
and U1891 (N_1891,N_1406,N_1001);
nand U1892 (N_1892,N_1242,N_1335);
and U1893 (N_1893,N_1004,N_1291);
and U1894 (N_1894,N_1270,N_1228);
xor U1895 (N_1895,N_1069,N_1458);
nor U1896 (N_1896,N_1142,N_1092);
or U1897 (N_1897,N_1373,N_1057);
or U1898 (N_1898,N_1113,N_1114);
nor U1899 (N_1899,N_1389,N_1309);
and U1900 (N_1900,N_1427,N_1281);
or U1901 (N_1901,N_1305,N_1176);
or U1902 (N_1902,N_1480,N_1117);
nor U1903 (N_1903,N_1270,N_1133);
nor U1904 (N_1904,N_1146,N_1119);
xnor U1905 (N_1905,N_1358,N_1256);
nor U1906 (N_1906,N_1126,N_1294);
and U1907 (N_1907,N_1000,N_1232);
or U1908 (N_1908,N_1181,N_1187);
or U1909 (N_1909,N_1308,N_1333);
nand U1910 (N_1910,N_1157,N_1238);
nand U1911 (N_1911,N_1332,N_1257);
nor U1912 (N_1912,N_1127,N_1476);
or U1913 (N_1913,N_1118,N_1334);
xnor U1914 (N_1914,N_1371,N_1069);
or U1915 (N_1915,N_1420,N_1195);
nor U1916 (N_1916,N_1210,N_1170);
xnor U1917 (N_1917,N_1484,N_1421);
nand U1918 (N_1918,N_1253,N_1250);
nand U1919 (N_1919,N_1079,N_1375);
or U1920 (N_1920,N_1289,N_1189);
nand U1921 (N_1921,N_1272,N_1132);
nor U1922 (N_1922,N_1258,N_1203);
nor U1923 (N_1923,N_1063,N_1466);
and U1924 (N_1924,N_1410,N_1354);
or U1925 (N_1925,N_1242,N_1249);
or U1926 (N_1926,N_1034,N_1393);
nand U1927 (N_1927,N_1194,N_1116);
nand U1928 (N_1928,N_1372,N_1315);
or U1929 (N_1929,N_1001,N_1332);
or U1930 (N_1930,N_1253,N_1462);
nand U1931 (N_1931,N_1277,N_1411);
or U1932 (N_1932,N_1184,N_1484);
or U1933 (N_1933,N_1155,N_1383);
or U1934 (N_1934,N_1045,N_1004);
nor U1935 (N_1935,N_1364,N_1092);
nor U1936 (N_1936,N_1092,N_1498);
and U1937 (N_1937,N_1091,N_1431);
or U1938 (N_1938,N_1135,N_1071);
or U1939 (N_1939,N_1181,N_1436);
or U1940 (N_1940,N_1458,N_1184);
and U1941 (N_1941,N_1001,N_1419);
or U1942 (N_1942,N_1020,N_1063);
nor U1943 (N_1943,N_1434,N_1061);
nand U1944 (N_1944,N_1288,N_1023);
and U1945 (N_1945,N_1165,N_1184);
nor U1946 (N_1946,N_1185,N_1401);
and U1947 (N_1947,N_1048,N_1180);
xnor U1948 (N_1948,N_1216,N_1105);
or U1949 (N_1949,N_1484,N_1299);
xor U1950 (N_1950,N_1164,N_1437);
nor U1951 (N_1951,N_1021,N_1236);
or U1952 (N_1952,N_1428,N_1285);
or U1953 (N_1953,N_1302,N_1386);
nor U1954 (N_1954,N_1474,N_1193);
xor U1955 (N_1955,N_1246,N_1277);
nor U1956 (N_1956,N_1181,N_1173);
or U1957 (N_1957,N_1458,N_1412);
nand U1958 (N_1958,N_1221,N_1284);
nand U1959 (N_1959,N_1169,N_1194);
nor U1960 (N_1960,N_1374,N_1112);
nand U1961 (N_1961,N_1428,N_1035);
nor U1962 (N_1962,N_1278,N_1345);
or U1963 (N_1963,N_1450,N_1032);
nand U1964 (N_1964,N_1056,N_1164);
nand U1965 (N_1965,N_1299,N_1141);
nor U1966 (N_1966,N_1433,N_1110);
nor U1967 (N_1967,N_1144,N_1062);
nand U1968 (N_1968,N_1245,N_1262);
and U1969 (N_1969,N_1453,N_1387);
xor U1970 (N_1970,N_1454,N_1286);
nand U1971 (N_1971,N_1207,N_1038);
xor U1972 (N_1972,N_1017,N_1089);
xnor U1973 (N_1973,N_1479,N_1334);
nand U1974 (N_1974,N_1089,N_1374);
nand U1975 (N_1975,N_1422,N_1284);
or U1976 (N_1976,N_1454,N_1175);
nor U1977 (N_1977,N_1378,N_1298);
nor U1978 (N_1978,N_1161,N_1486);
and U1979 (N_1979,N_1263,N_1077);
and U1980 (N_1980,N_1360,N_1383);
and U1981 (N_1981,N_1345,N_1209);
nor U1982 (N_1982,N_1336,N_1309);
or U1983 (N_1983,N_1204,N_1157);
or U1984 (N_1984,N_1363,N_1017);
nand U1985 (N_1985,N_1040,N_1062);
nand U1986 (N_1986,N_1055,N_1143);
nor U1987 (N_1987,N_1191,N_1318);
xnor U1988 (N_1988,N_1013,N_1062);
or U1989 (N_1989,N_1422,N_1099);
nor U1990 (N_1990,N_1349,N_1276);
nor U1991 (N_1991,N_1104,N_1050);
nand U1992 (N_1992,N_1363,N_1403);
and U1993 (N_1993,N_1421,N_1100);
nor U1994 (N_1994,N_1178,N_1163);
nand U1995 (N_1995,N_1199,N_1225);
nand U1996 (N_1996,N_1357,N_1118);
nand U1997 (N_1997,N_1138,N_1235);
nor U1998 (N_1998,N_1432,N_1348);
or U1999 (N_1999,N_1084,N_1281);
nand U2000 (N_2000,N_1866,N_1728);
xor U2001 (N_2001,N_1787,N_1687);
and U2002 (N_2002,N_1760,N_1979);
or U2003 (N_2003,N_1905,N_1537);
xnor U2004 (N_2004,N_1689,N_1527);
nand U2005 (N_2005,N_1761,N_1660);
xnor U2006 (N_2006,N_1657,N_1535);
nor U2007 (N_2007,N_1857,N_1950);
nand U2008 (N_2008,N_1526,N_1544);
nor U2009 (N_2009,N_1788,N_1915);
and U2010 (N_2010,N_1700,N_1991);
or U2011 (N_2011,N_1989,N_1503);
nor U2012 (N_2012,N_1607,N_1798);
nand U2013 (N_2013,N_1861,N_1634);
and U2014 (N_2014,N_1724,N_1715);
nor U2015 (N_2015,N_1894,N_1990);
nor U2016 (N_2016,N_1500,N_1834);
nand U2017 (N_2017,N_1563,N_1932);
and U2018 (N_2018,N_1789,N_1704);
and U2019 (N_2019,N_1851,N_1650);
xnor U2020 (N_2020,N_1580,N_1688);
and U2021 (N_2021,N_1868,N_1983);
nor U2022 (N_2022,N_1869,N_1648);
nand U2023 (N_2023,N_1938,N_1890);
and U2024 (N_2024,N_1532,N_1978);
or U2025 (N_2025,N_1848,N_1763);
and U2026 (N_2026,N_1686,N_1737);
nor U2027 (N_2027,N_1792,N_1940);
or U2028 (N_2028,N_1505,N_1923);
or U2029 (N_2029,N_1731,N_1804);
nor U2030 (N_2030,N_1604,N_1546);
and U2031 (N_2031,N_1738,N_1553);
nand U2032 (N_2032,N_1810,N_1528);
nand U2033 (N_2033,N_1930,N_1605);
xor U2034 (N_2034,N_1709,N_1734);
nand U2035 (N_2035,N_1511,N_1720);
or U2036 (N_2036,N_1672,N_1655);
or U2037 (N_2037,N_1741,N_1740);
xor U2038 (N_2038,N_1939,N_1921);
nand U2039 (N_2039,N_1818,N_1632);
or U2040 (N_2040,N_1529,N_1716);
nand U2041 (N_2041,N_1762,N_1576);
nand U2042 (N_2042,N_1730,N_1574);
nand U2043 (N_2043,N_1805,N_1566);
or U2044 (N_2044,N_1729,N_1667);
and U2045 (N_2045,N_1561,N_1562);
xor U2046 (N_2046,N_1901,N_1854);
or U2047 (N_2047,N_1886,N_1876);
or U2048 (N_2048,N_1696,N_1895);
nand U2049 (N_2049,N_1823,N_1897);
nor U2050 (N_2050,N_1556,N_1998);
or U2051 (N_2051,N_1899,N_1530);
xnor U2052 (N_2052,N_1784,N_1839);
xnor U2053 (N_2053,N_1765,N_1969);
nor U2054 (N_2054,N_1985,N_1538);
and U2055 (N_2055,N_1598,N_1555);
nor U2056 (N_2056,N_1842,N_1786);
or U2057 (N_2057,N_1611,N_1705);
and U2058 (N_2058,N_1582,N_1552);
nand U2059 (N_2059,N_1822,N_1852);
or U2060 (N_2060,N_1924,N_1987);
or U2061 (N_2061,N_1508,N_1992);
or U2062 (N_2062,N_1585,N_1577);
and U2063 (N_2063,N_1663,N_1707);
nor U2064 (N_2064,N_1519,N_1695);
nand U2065 (N_2065,N_1829,N_1504);
xor U2066 (N_2066,N_1984,N_1775);
nand U2067 (N_2067,N_1617,N_1692);
nand U2068 (N_2068,N_1942,N_1995);
and U2069 (N_2069,N_1539,N_1898);
nor U2070 (N_2070,N_1652,N_1599);
nand U2071 (N_2071,N_1799,N_1739);
or U2072 (N_2072,N_1625,N_1910);
nor U2073 (N_2073,N_1791,N_1545);
nor U2074 (N_2074,N_1849,N_1759);
and U2075 (N_2075,N_1997,N_1840);
and U2076 (N_2076,N_1690,N_1743);
nor U2077 (N_2077,N_1770,N_1831);
nand U2078 (N_2078,N_1635,N_1571);
or U2079 (N_2079,N_1964,N_1524);
xnor U2080 (N_2080,N_1835,N_1613);
nand U2081 (N_2081,N_1844,N_1664);
nand U2082 (N_2082,N_1683,N_1946);
nand U2083 (N_2083,N_1865,N_1960);
xor U2084 (N_2084,N_1722,N_1879);
and U2085 (N_2085,N_1748,N_1862);
or U2086 (N_2086,N_1751,N_1838);
nand U2087 (N_2087,N_1917,N_1793);
nor U2088 (N_2088,N_1974,N_1907);
nor U2089 (N_2089,N_1887,N_1502);
nand U2090 (N_2090,N_1699,N_1821);
or U2091 (N_2091,N_1712,N_1558);
or U2092 (N_2092,N_1518,N_1806);
nor U2093 (N_2093,N_1883,N_1833);
and U2094 (N_2094,N_1767,N_1994);
nor U2095 (N_2095,N_1808,N_1661);
xnor U2096 (N_2096,N_1976,N_1785);
or U2097 (N_2097,N_1855,N_1903);
nor U2098 (N_2098,N_1579,N_1936);
nand U2099 (N_2099,N_1780,N_1698);
nor U2100 (N_2100,N_1797,N_1628);
or U2101 (N_2101,N_1774,N_1586);
nand U2102 (N_2102,N_1627,N_1515);
and U2103 (N_2103,N_1637,N_1597);
xnor U2104 (N_2104,N_1813,N_1837);
xnor U2105 (N_2105,N_1981,N_1841);
nor U2106 (N_2106,N_1647,N_1856);
and U2107 (N_2107,N_1593,N_1610);
xor U2108 (N_2108,N_1928,N_1509);
nor U2109 (N_2109,N_1522,N_1682);
xor U2110 (N_2110,N_1587,N_1809);
or U2111 (N_2111,N_1825,N_1870);
xnor U2112 (N_2112,N_1764,N_1772);
or U2113 (N_2113,N_1746,N_1807);
and U2114 (N_2114,N_1830,N_1977);
nor U2115 (N_2115,N_1670,N_1570);
nor U2116 (N_2116,N_1754,N_1961);
nand U2117 (N_2117,N_1679,N_1671);
nor U2118 (N_2118,N_1684,N_1711);
xor U2119 (N_2119,N_1814,N_1955);
xor U2120 (N_2120,N_1547,N_1645);
xnor U2121 (N_2121,N_1513,N_1733);
nand U2122 (N_2122,N_1612,N_1567);
or U2123 (N_2123,N_1656,N_1626);
or U2124 (N_2124,N_1512,N_1957);
nand U2125 (N_2125,N_1768,N_1758);
nand U2126 (N_2126,N_1820,N_1859);
or U2127 (N_2127,N_1771,N_1596);
nand U2128 (N_2128,N_1676,N_1536);
or U2129 (N_2129,N_1967,N_1795);
nand U2130 (N_2130,N_1736,N_1615);
and U2131 (N_2131,N_1874,N_1554);
nand U2132 (N_2132,N_1778,N_1678);
or U2133 (N_2133,N_1790,N_1638);
and U2134 (N_2134,N_1581,N_1506);
and U2135 (N_2135,N_1973,N_1846);
nand U2136 (N_2136,N_1871,N_1620);
nor U2137 (N_2137,N_1525,N_1680);
nand U2138 (N_2138,N_1777,N_1944);
nand U2139 (N_2139,N_1710,N_1590);
nor U2140 (N_2140,N_1726,N_1776);
nor U2141 (N_2141,N_1832,N_1675);
or U2142 (N_2142,N_1622,N_1952);
and U2143 (N_2143,N_1920,N_1877);
or U2144 (N_2144,N_1947,N_1937);
or U2145 (N_2145,N_1845,N_1941);
or U2146 (N_2146,N_1640,N_1904);
and U2147 (N_2147,N_1847,N_1623);
or U2148 (N_2148,N_1826,N_1836);
nand U2149 (N_2149,N_1867,N_1551);
and U2150 (N_2150,N_1618,N_1569);
nand U2151 (N_2151,N_1970,N_1589);
xor U2152 (N_2152,N_1636,N_1853);
nand U2153 (N_2153,N_1996,N_1583);
nor U2154 (N_2154,N_1747,N_1673);
nor U2155 (N_2155,N_1662,N_1706);
nor U2156 (N_2156,N_1843,N_1926);
and U2157 (N_2157,N_1616,N_1993);
and U2158 (N_2158,N_1954,N_1919);
nor U2159 (N_2159,N_1510,N_1802);
or U2160 (N_2160,N_1911,N_1828);
nor U2161 (N_2161,N_1742,N_1817);
nor U2162 (N_2162,N_1732,N_1752);
and U2163 (N_2163,N_1864,N_1912);
nand U2164 (N_2164,N_1578,N_1971);
or U2165 (N_2165,N_1816,N_1882);
and U2166 (N_2166,N_1669,N_1630);
and U2167 (N_2167,N_1631,N_1641);
or U2168 (N_2168,N_1697,N_1560);
nand U2169 (N_2169,N_1872,N_1881);
or U2170 (N_2170,N_1665,N_1531);
nor U2171 (N_2171,N_1794,N_1906);
or U2172 (N_2172,N_1727,N_1694);
or U2173 (N_2173,N_1639,N_1773);
nand U2174 (N_2174,N_1934,N_1900);
nand U2175 (N_2175,N_1735,N_1557);
or U2176 (N_2176,N_1933,N_1884);
or U2177 (N_2177,N_1800,N_1540);
nand U2178 (N_2178,N_1668,N_1914);
or U2179 (N_2179,N_1703,N_1542);
nor U2180 (N_2180,N_1931,N_1573);
and U2181 (N_2181,N_1643,N_1507);
or U2182 (N_2182,N_1674,N_1965);
or U2183 (N_2183,N_1811,N_1603);
nand U2184 (N_2184,N_1548,N_1677);
nor U2185 (N_2185,N_1803,N_1781);
and U2186 (N_2186,N_1935,N_1516);
and U2187 (N_2187,N_1922,N_1588);
and U2188 (N_2188,N_1889,N_1606);
and U2189 (N_2189,N_1584,N_1873);
or U2190 (N_2190,N_1602,N_1908);
and U2191 (N_2191,N_1708,N_1609);
or U2192 (N_2192,N_1896,N_1651);
and U2193 (N_2193,N_1949,N_1929);
nor U2194 (N_2194,N_1916,N_1909);
nor U2195 (N_2195,N_1968,N_1719);
nor U2196 (N_2196,N_1723,N_1541);
nor U2197 (N_2197,N_1594,N_1572);
nor U2198 (N_2198,N_1875,N_1959);
nand U2199 (N_2199,N_1501,N_1956);
nor U2200 (N_2200,N_1685,N_1757);
or U2201 (N_2201,N_1953,N_1659);
or U2202 (N_2202,N_1812,N_1714);
and U2203 (N_2203,N_1693,N_1766);
and U2204 (N_2204,N_1963,N_1533);
or U2205 (N_2205,N_1520,N_1559);
nor U2206 (N_2206,N_1815,N_1592);
or U2207 (N_2207,N_1927,N_1943);
or U2208 (N_2208,N_1717,N_1878);
nand U2209 (N_2209,N_1750,N_1591);
nand U2210 (N_2210,N_1608,N_1779);
or U2211 (N_2211,N_1892,N_1575);
nor U2212 (N_2212,N_1796,N_1913);
nand U2213 (N_2213,N_1982,N_1713);
and U2214 (N_2214,N_1918,N_1745);
nor U2215 (N_2215,N_1948,N_1629);
or U2216 (N_2216,N_1782,N_1614);
or U2217 (N_2217,N_1595,N_1749);
nand U2218 (N_2218,N_1653,N_1543);
nor U2219 (N_2219,N_1549,N_1988);
nor U2220 (N_2220,N_1966,N_1858);
or U2221 (N_2221,N_1666,N_1755);
and U2222 (N_2222,N_1521,N_1958);
nor U2223 (N_2223,N_1975,N_1880);
nor U2224 (N_2224,N_1827,N_1621);
xnor U2225 (N_2225,N_1691,N_1951);
and U2226 (N_2226,N_1701,N_1601);
nand U2227 (N_2227,N_1888,N_1925);
nand U2228 (N_2228,N_1624,N_1718);
or U2229 (N_2229,N_1550,N_1769);
nand U2230 (N_2230,N_1517,N_1564);
nor U2231 (N_2231,N_1658,N_1565);
nand U2232 (N_2232,N_1885,N_1783);
nor U2233 (N_2233,N_1753,N_1962);
nor U2234 (N_2234,N_1514,N_1891);
nand U2235 (N_2235,N_1646,N_1568);
nor U2236 (N_2236,N_1619,N_1649);
and U2237 (N_2237,N_1523,N_1893);
and U2238 (N_2238,N_1980,N_1824);
nand U2239 (N_2239,N_1681,N_1902);
and U2240 (N_2240,N_1756,N_1721);
or U2241 (N_2241,N_1654,N_1999);
or U2242 (N_2242,N_1972,N_1863);
and U2243 (N_2243,N_1725,N_1986);
nor U2244 (N_2244,N_1600,N_1633);
nand U2245 (N_2245,N_1644,N_1801);
or U2246 (N_2246,N_1860,N_1850);
nand U2247 (N_2247,N_1534,N_1744);
or U2248 (N_2248,N_1642,N_1819);
and U2249 (N_2249,N_1945,N_1702);
xnor U2250 (N_2250,N_1684,N_1525);
and U2251 (N_2251,N_1566,N_1583);
nand U2252 (N_2252,N_1835,N_1610);
nand U2253 (N_2253,N_1699,N_1883);
xnor U2254 (N_2254,N_1840,N_1749);
nor U2255 (N_2255,N_1888,N_1765);
nor U2256 (N_2256,N_1579,N_1703);
or U2257 (N_2257,N_1653,N_1881);
nor U2258 (N_2258,N_1565,N_1531);
nand U2259 (N_2259,N_1730,N_1530);
xor U2260 (N_2260,N_1859,N_1524);
nor U2261 (N_2261,N_1805,N_1914);
and U2262 (N_2262,N_1834,N_1920);
or U2263 (N_2263,N_1693,N_1858);
or U2264 (N_2264,N_1814,N_1885);
nor U2265 (N_2265,N_1815,N_1727);
or U2266 (N_2266,N_1999,N_1650);
nand U2267 (N_2267,N_1948,N_1851);
and U2268 (N_2268,N_1623,N_1674);
nor U2269 (N_2269,N_1561,N_1573);
or U2270 (N_2270,N_1615,N_1749);
xnor U2271 (N_2271,N_1816,N_1823);
nand U2272 (N_2272,N_1908,N_1856);
and U2273 (N_2273,N_1949,N_1765);
and U2274 (N_2274,N_1777,N_1948);
or U2275 (N_2275,N_1591,N_1782);
and U2276 (N_2276,N_1622,N_1733);
nand U2277 (N_2277,N_1940,N_1728);
nand U2278 (N_2278,N_1547,N_1605);
xnor U2279 (N_2279,N_1677,N_1652);
nand U2280 (N_2280,N_1553,N_1971);
nor U2281 (N_2281,N_1657,N_1722);
and U2282 (N_2282,N_1911,N_1708);
and U2283 (N_2283,N_1814,N_1863);
nand U2284 (N_2284,N_1616,N_1923);
nand U2285 (N_2285,N_1519,N_1846);
xnor U2286 (N_2286,N_1546,N_1588);
nand U2287 (N_2287,N_1642,N_1686);
and U2288 (N_2288,N_1782,N_1754);
xor U2289 (N_2289,N_1768,N_1975);
or U2290 (N_2290,N_1686,N_1553);
and U2291 (N_2291,N_1775,N_1898);
nor U2292 (N_2292,N_1566,N_1844);
nor U2293 (N_2293,N_1709,N_1988);
and U2294 (N_2294,N_1913,N_1633);
or U2295 (N_2295,N_1535,N_1571);
nor U2296 (N_2296,N_1624,N_1766);
or U2297 (N_2297,N_1882,N_1675);
nand U2298 (N_2298,N_1969,N_1708);
nor U2299 (N_2299,N_1619,N_1792);
nor U2300 (N_2300,N_1636,N_1964);
nand U2301 (N_2301,N_1881,N_1839);
xor U2302 (N_2302,N_1589,N_1744);
or U2303 (N_2303,N_1813,N_1515);
nor U2304 (N_2304,N_1557,N_1761);
nand U2305 (N_2305,N_1514,N_1693);
xnor U2306 (N_2306,N_1709,N_1803);
nor U2307 (N_2307,N_1931,N_1790);
and U2308 (N_2308,N_1998,N_1900);
and U2309 (N_2309,N_1894,N_1966);
nand U2310 (N_2310,N_1952,N_1993);
and U2311 (N_2311,N_1989,N_1712);
nor U2312 (N_2312,N_1924,N_1794);
nor U2313 (N_2313,N_1564,N_1914);
xnor U2314 (N_2314,N_1938,N_1617);
and U2315 (N_2315,N_1746,N_1845);
or U2316 (N_2316,N_1545,N_1936);
or U2317 (N_2317,N_1851,N_1790);
nand U2318 (N_2318,N_1963,N_1843);
nand U2319 (N_2319,N_1942,N_1916);
and U2320 (N_2320,N_1946,N_1970);
nand U2321 (N_2321,N_1847,N_1527);
or U2322 (N_2322,N_1525,N_1500);
or U2323 (N_2323,N_1900,N_1536);
and U2324 (N_2324,N_1709,N_1641);
and U2325 (N_2325,N_1681,N_1534);
or U2326 (N_2326,N_1737,N_1523);
or U2327 (N_2327,N_1754,N_1636);
or U2328 (N_2328,N_1853,N_1649);
nand U2329 (N_2329,N_1643,N_1934);
or U2330 (N_2330,N_1614,N_1644);
nor U2331 (N_2331,N_1687,N_1688);
nand U2332 (N_2332,N_1690,N_1874);
nor U2333 (N_2333,N_1562,N_1502);
nor U2334 (N_2334,N_1814,N_1925);
and U2335 (N_2335,N_1683,N_1544);
nor U2336 (N_2336,N_1845,N_1620);
and U2337 (N_2337,N_1535,N_1607);
nand U2338 (N_2338,N_1688,N_1741);
nand U2339 (N_2339,N_1907,N_1599);
and U2340 (N_2340,N_1631,N_1612);
and U2341 (N_2341,N_1656,N_1609);
nand U2342 (N_2342,N_1635,N_1760);
and U2343 (N_2343,N_1956,N_1669);
nor U2344 (N_2344,N_1597,N_1956);
nand U2345 (N_2345,N_1917,N_1979);
nor U2346 (N_2346,N_1714,N_1823);
nor U2347 (N_2347,N_1527,N_1650);
or U2348 (N_2348,N_1716,N_1915);
xnor U2349 (N_2349,N_1604,N_1630);
nand U2350 (N_2350,N_1910,N_1599);
and U2351 (N_2351,N_1969,N_1680);
nor U2352 (N_2352,N_1694,N_1666);
and U2353 (N_2353,N_1587,N_1828);
nor U2354 (N_2354,N_1686,N_1894);
and U2355 (N_2355,N_1954,N_1992);
xnor U2356 (N_2356,N_1741,N_1527);
or U2357 (N_2357,N_1795,N_1514);
xor U2358 (N_2358,N_1746,N_1513);
or U2359 (N_2359,N_1913,N_1979);
or U2360 (N_2360,N_1557,N_1997);
and U2361 (N_2361,N_1842,N_1859);
or U2362 (N_2362,N_1574,N_1630);
or U2363 (N_2363,N_1725,N_1657);
and U2364 (N_2364,N_1853,N_1931);
and U2365 (N_2365,N_1601,N_1891);
and U2366 (N_2366,N_1796,N_1781);
and U2367 (N_2367,N_1578,N_1737);
nand U2368 (N_2368,N_1548,N_1860);
or U2369 (N_2369,N_1562,N_1689);
and U2370 (N_2370,N_1787,N_1679);
or U2371 (N_2371,N_1500,N_1687);
nand U2372 (N_2372,N_1529,N_1834);
and U2373 (N_2373,N_1600,N_1741);
xnor U2374 (N_2374,N_1706,N_1946);
nor U2375 (N_2375,N_1505,N_1530);
or U2376 (N_2376,N_1941,N_1576);
or U2377 (N_2377,N_1990,N_1515);
or U2378 (N_2378,N_1717,N_1616);
or U2379 (N_2379,N_1914,N_1502);
or U2380 (N_2380,N_1935,N_1768);
and U2381 (N_2381,N_1955,N_1767);
or U2382 (N_2382,N_1872,N_1863);
nor U2383 (N_2383,N_1670,N_1960);
nand U2384 (N_2384,N_1604,N_1724);
nor U2385 (N_2385,N_1917,N_1512);
and U2386 (N_2386,N_1577,N_1625);
and U2387 (N_2387,N_1702,N_1555);
nand U2388 (N_2388,N_1552,N_1845);
and U2389 (N_2389,N_1809,N_1834);
nand U2390 (N_2390,N_1800,N_1813);
and U2391 (N_2391,N_1889,N_1699);
nor U2392 (N_2392,N_1570,N_1805);
xor U2393 (N_2393,N_1923,N_1717);
nand U2394 (N_2394,N_1841,N_1774);
xor U2395 (N_2395,N_1892,N_1956);
nor U2396 (N_2396,N_1963,N_1924);
or U2397 (N_2397,N_1643,N_1710);
and U2398 (N_2398,N_1741,N_1554);
nand U2399 (N_2399,N_1501,N_1705);
nor U2400 (N_2400,N_1891,N_1832);
or U2401 (N_2401,N_1858,N_1673);
and U2402 (N_2402,N_1915,N_1760);
or U2403 (N_2403,N_1705,N_1829);
or U2404 (N_2404,N_1766,N_1799);
nand U2405 (N_2405,N_1933,N_1705);
nand U2406 (N_2406,N_1501,N_1813);
xnor U2407 (N_2407,N_1674,N_1991);
or U2408 (N_2408,N_1833,N_1666);
and U2409 (N_2409,N_1615,N_1939);
and U2410 (N_2410,N_1504,N_1597);
and U2411 (N_2411,N_1774,N_1836);
xnor U2412 (N_2412,N_1877,N_1652);
nand U2413 (N_2413,N_1987,N_1797);
and U2414 (N_2414,N_1681,N_1967);
and U2415 (N_2415,N_1879,N_1615);
or U2416 (N_2416,N_1633,N_1779);
nor U2417 (N_2417,N_1765,N_1811);
and U2418 (N_2418,N_1869,N_1515);
and U2419 (N_2419,N_1556,N_1780);
nor U2420 (N_2420,N_1844,N_1636);
and U2421 (N_2421,N_1675,N_1903);
nand U2422 (N_2422,N_1561,N_1934);
nor U2423 (N_2423,N_1822,N_1685);
nand U2424 (N_2424,N_1922,N_1957);
nor U2425 (N_2425,N_1985,N_1541);
nand U2426 (N_2426,N_1680,N_1935);
or U2427 (N_2427,N_1560,N_1877);
or U2428 (N_2428,N_1760,N_1675);
nor U2429 (N_2429,N_1811,N_1624);
nand U2430 (N_2430,N_1895,N_1896);
and U2431 (N_2431,N_1581,N_1950);
or U2432 (N_2432,N_1930,N_1802);
and U2433 (N_2433,N_1659,N_1827);
nand U2434 (N_2434,N_1887,N_1814);
or U2435 (N_2435,N_1929,N_1805);
nor U2436 (N_2436,N_1735,N_1654);
or U2437 (N_2437,N_1641,N_1703);
and U2438 (N_2438,N_1989,N_1816);
xor U2439 (N_2439,N_1805,N_1727);
or U2440 (N_2440,N_1888,N_1621);
or U2441 (N_2441,N_1983,N_1745);
nor U2442 (N_2442,N_1978,N_1652);
and U2443 (N_2443,N_1818,N_1783);
and U2444 (N_2444,N_1602,N_1978);
nand U2445 (N_2445,N_1515,N_1632);
nand U2446 (N_2446,N_1588,N_1808);
and U2447 (N_2447,N_1943,N_1867);
and U2448 (N_2448,N_1724,N_1819);
nand U2449 (N_2449,N_1720,N_1994);
nand U2450 (N_2450,N_1761,N_1576);
xnor U2451 (N_2451,N_1551,N_1614);
nand U2452 (N_2452,N_1883,N_1505);
nand U2453 (N_2453,N_1806,N_1570);
nand U2454 (N_2454,N_1663,N_1712);
nor U2455 (N_2455,N_1901,N_1764);
nand U2456 (N_2456,N_1879,N_1767);
and U2457 (N_2457,N_1656,N_1865);
nand U2458 (N_2458,N_1746,N_1698);
nand U2459 (N_2459,N_1929,N_1800);
xnor U2460 (N_2460,N_1793,N_1538);
or U2461 (N_2461,N_1851,N_1841);
or U2462 (N_2462,N_1866,N_1736);
nand U2463 (N_2463,N_1581,N_1909);
or U2464 (N_2464,N_1899,N_1922);
or U2465 (N_2465,N_1506,N_1939);
nand U2466 (N_2466,N_1951,N_1596);
xnor U2467 (N_2467,N_1877,N_1696);
nand U2468 (N_2468,N_1624,N_1920);
nand U2469 (N_2469,N_1765,N_1553);
and U2470 (N_2470,N_1553,N_1721);
nor U2471 (N_2471,N_1856,N_1534);
nand U2472 (N_2472,N_1771,N_1550);
or U2473 (N_2473,N_1794,N_1567);
or U2474 (N_2474,N_1606,N_1687);
or U2475 (N_2475,N_1937,N_1634);
or U2476 (N_2476,N_1661,N_1908);
xor U2477 (N_2477,N_1961,N_1782);
nand U2478 (N_2478,N_1863,N_1795);
and U2479 (N_2479,N_1513,N_1650);
or U2480 (N_2480,N_1983,N_1655);
and U2481 (N_2481,N_1746,N_1819);
nor U2482 (N_2482,N_1931,N_1778);
and U2483 (N_2483,N_1684,N_1567);
nor U2484 (N_2484,N_1786,N_1665);
or U2485 (N_2485,N_1665,N_1800);
or U2486 (N_2486,N_1621,N_1691);
xor U2487 (N_2487,N_1663,N_1699);
nand U2488 (N_2488,N_1868,N_1907);
nor U2489 (N_2489,N_1870,N_1693);
xnor U2490 (N_2490,N_1774,N_1550);
xor U2491 (N_2491,N_1838,N_1875);
nor U2492 (N_2492,N_1580,N_1625);
nand U2493 (N_2493,N_1676,N_1608);
or U2494 (N_2494,N_1874,N_1903);
or U2495 (N_2495,N_1713,N_1867);
nor U2496 (N_2496,N_1507,N_1670);
and U2497 (N_2497,N_1948,N_1526);
nor U2498 (N_2498,N_1557,N_1829);
nand U2499 (N_2499,N_1881,N_1929);
xnor U2500 (N_2500,N_2314,N_2385);
or U2501 (N_2501,N_2278,N_2174);
and U2502 (N_2502,N_2166,N_2342);
nor U2503 (N_2503,N_2008,N_2115);
nor U2504 (N_2504,N_2212,N_2109);
nor U2505 (N_2505,N_2307,N_2260);
nand U2506 (N_2506,N_2124,N_2226);
nor U2507 (N_2507,N_2257,N_2471);
xor U2508 (N_2508,N_2494,N_2053);
or U2509 (N_2509,N_2203,N_2410);
or U2510 (N_2510,N_2277,N_2335);
nor U2511 (N_2511,N_2327,N_2476);
or U2512 (N_2512,N_2478,N_2297);
xnor U2513 (N_2513,N_2180,N_2369);
nor U2514 (N_2514,N_2444,N_2487);
or U2515 (N_2515,N_2414,N_2113);
or U2516 (N_2516,N_2366,N_2253);
and U2517 (N_2517,N_2001,N_2427);
and U2518 (N_2518,N_2423,N_2356);
and U2519 (N_2519,N_2289,N_2378);
or U2520 (N_2520,N_2035,N_2225);
nand U2521 (N_2521,N_2014,N_2178);
and U2522 (N_2522,N_2400,N_2373);
or U2523 (N_2523,N_2164,N_2172);
or U2524 (N_2524,N_2199,N_2375);
or U2525 (N_2525,N_2310,N_2096);
xor U2526 (N_2526,N_2092,N_2036);
or U2527 (N_2527,N_2029,N_2136);
or U2528 (N_2528,N_2065,N_2102);
nand U2529 (N_2529,N_2087,N_2118);
and U2530 (N_2530,N_2480,N_2252);
or U2531 (N_2531,N_2333,N_2497);
and U2532 (N_2532,N_2493,N_2176);
or U2533 (N_2533,N_2066,N_2192);
nor U2534 (N_2534,N_2391,N_2145);
nand U2535 (N_2535,N_2470,N_2394);
nand U2536 (N_2536,N_2303,N_2147);
and U2537 (N_2537,N_2262,N_2383);
nand U2538 (N_2538,N_2350,N_2439);
and U2539 (N_2539,N_2175,N_2293);
or U2540 (N_2540,N_2355,N_2110);
nand U2541 (N_2541,N_2033,N_2430);
nor U2542 (N_2542,N_2462,N_2438);
nand U2543 (N_2543,N_2059,N_2049);
nor U2544 (N_2544,N_2265,N_2492);
nand U2545 (N_2545,N_2125,N_2422);
xor U2546 (N_2546,N_2085,N_2190);
or U2547 (N_2547,N_2417,N_2481);
and U2548 (N_2548,N_2005,N_2112);
nand U2549 (N_2549,N_2086,N_2041);
nor U2550 (N_2550,N_2181,N_2298);
and U2551 (N_2551,N_2249,N_2283);
nand U2552 (N_2552,N_2149,N_2271);
and U2553 (N_2553,N_2357,N_2047);
or U2554 (N_2554,N_2445,N_2498);
and U2555 (N_2555,N_2062,N_2479);
nor U2556 (N_2556,N_2287,N_2067);
nand U2557 (N_2557,N_2420,N_2093);
or U2558 (N_2558,N_2248,N_2116);
and U2559 (N_2559,N_2339,N_2302);
and U2560 (N_2560,N_2197,N_2456);
and U2561 (N_2561,N_2153,N_2241);
and U2562 (N_2562,N_2240,N_2051);
nor U2563 (N_2563,N_2031,N_2050);
or U2564 (N_2564,N_2448,N_2003);
nor U2565 (N_2565,N_2360,N_2305);
and U2566 (N_2566,N_2021,N_2082);
xnor U2567 (N_2567,N_2043,N_2465);
or U2568 (N_2568,N_2362,N_2200);
nand U2569 (N_2569,N_2274,N_2018);
nand U2570 (N_2570,N_2006,N_2429);
nand U2571 (N_2571,N_2443,N_2434);
xor U2572 (N_2572,N_2080,N_2210);
nand U2573 (N_2573,N_2455,N_2399);
nand U2574 (N_2574,N_2411,N_2209);
nand U2575 (N_2575,N_2388,N_2323);
or U2576 (N_2576,N_2127,N_2398);
nor U2577 (N_2577,N_2030,N_2404);
nand U2578 (N_2578,N_2461,N_2157);
nor U2579 (N_2579,N_2027,N_2010);
or U2580 (N_2580,N_2040,N_2119);
and U2581 (N_2581,N_2464,N_2189);
nand U2582 (N_2582,N_2337,N_2346);
or U2583 (N_2583,N_2348,N_2474);
nor U2584 (N_2584,N_2256,N_2367);
xor U2585 (N_2585,N_2216,N_2143);
and U2586 (N_2586,N_2321,N_2205);
or U2587 (N_2587,N_2340,N_2389);
nor U2588 (N_2588,N_2239,N_2352);
or U2589 (N_2589,N_2120,N_2382);
xor U2590 (N_2590,N_2114,N_2324);
and U2591 (N_2591,N_2467,N_2009);
nor U2592 (N_2592,N_2194,N_2170);
and U2593 (N_2593,N_2242,N_2251);
nor U2594 (N_2594,N_2151,N_2440);
nor U2595 (N_2595,N_2020,N_2351);
or U2596 (N_2596,N_2338,N_2075);
or U2597 (N_2597,N_2048,N_2042);
nor U2598 (N_2598,N_2024,N_2344);
and U2599 (N_2599,N_2246,N_2486);
and U2600 (N_2600,N_2221,N_2215);
nand U2601 (N_2601,N_2140,N_2039);
nor U2602 (N_2602,N_2276,N_2473);
nand U2603 (N_2603,N_2295,N_2095);
or U2604 (N_2604,N_2079,N_2273);
xor U2605 (N_2605,N_2126,N_2211);
or U2606 (N_2606,N_2070,N_2407);
and U2607 (N_2607,N_2488,N_2468);
and U2608 (N_2608,N_2472,N_2223);
nand U2609 (N_2609,N_2122,N_2424);
or U2610 (N_2610,N_2167,N_2182);
nand U2611 (N_2611,N_2466,N_2393);
and U2612 (N_2612,N_2475,N_2090);
xor U2613 (N_2613,N_2421,N_2282);
and U2614 (N_2614,N_2207,N_2158);
or U2615 (N_2615,N_2163,N_2371);
xor U2616 (N_2616,N_2229,N_2368);
or U2617 (N_2617,N_2451,N_2364);
nor U2618 (N_2618,N_2372,N_2442);
nand U2619 (N_2619,N_2330,N_2219);
and U2620 (N_2620,N_2447,N_2272);
and U2621 (N_2621,N_2365,N_2418);
and U2622 (N_2622,N_2435,N_2015);
and U2623 (N_2623,N_2384,N_2098);
nand U2624 (N_2624,N_2237,N_2083);
nor U2625 (N_2625,N_2428,N_2266);
and U2626 (N_2626,N_2173,N_2259);
xor U2627 (N_2627,N_2142,N_2132);
nand U2628 (N_2628,N_2204,N_2325);
and U2629 (N_2629,N_2409,N_2312);
nand U2630 (N_2630,N_2154,N_2416);
and U2631 (N_2631,N_2236,N_2315);
and U2632 (N_2632,N_2381,N_2165);
and U2633 (N_2633,N_2396,N_2458);
nand U2634 (N_2634,N_2477,N_2441);
nor U2635 (N_2635,N_2117,N_2220);
or U2636 (N_2636,N_2074,N_2285);
nand U2637 (N_2637,N_2183,N_2446);
nand U2638 (N_2638,N_2301,N_2206);
nand U2639 (N_2639,N_2485,N_2380);
nor U2640 (N_2640,N_2152,N_2306);
or U2641 (N_2641,N_2160,N_2186);
nand U2642 (N_2642,N_2131,N_2454);
nand U2643 (N_2643,N_2099,N_2234);
nor U2644 (N_2644,N_2012,N_2004);
or U2645 (N_2645,N_2244,N_2291);
and U2646 (N_2646,N_2000,N_2218);
nor U2647 (N_2647,N_2309,N_2491);
nand U2648 (N_2648,N_2290,N_2017);
or U2649 (N_2649,N_2261,N_2308);
nand U2650 (N_2650,N_2247,N_2076);
and U2651 (N_2651,N_2359,N_2425);
nand U2652 (N_2652,N_2134,N_2161);
xor U2653 (N_2653,N_2387,N_2055);
or U2654 (N_2654,N_2453,N_2436);
nor U2655 (N_2655,N_2162,N_2336);
nor U2656 (N_2656,N_2347,N_2452);
xnor U2657 (N_2657,N_2299,N_2402);
nand U2658 (N_2658,N_2353,N_2227);
and U2659 (N_2659,N_2483,N_2184);
and U2660 (N_2660,N_2254,N_2034);
or U2661 (N_2661,N_2077,N_2311);
or U2662 (N_2662,N_2187,N_2135);
or U2663 (N_2663,N_2129,N_2155);
nor U2664 (N_2664,N_2296,N_2103);
xor U2665 (N_2665,N_2361,N_2379);
or U2666 (N_2666,N_2294,N_2171);
nand U2667 (N_2667,N_2072,N_2345);
or U2668 (N_2668,N_2013,N_2358);
and U2669 (N_2669,N_2088,N_2395);
or U2670 (N_2670,N_2270,N_2469);
nand U2671 (N_2671,N_2264,N_2329);
or U2672 (N_2672,N_2107,N_2419);
nand U2673 (N_2673,N_2268,N_2484);
and U2674 (N_2674,N_2354,N_2449);
and U2675 (N_2675,N_2104,N_2332);
nor U2676 (N_2676,N_2032,N_2193);
nand U2677 (N_2677,N_2130,N_2201);
or U2678 (N_2678,N_2097,N_2286);
nand U2679 (N_2679,N_2450,N_2392);
nor U2680 (N_2680,N_2044,N_2284);
and U2681 (N_2681,N_2222,N_2101);
and U2682 (N_2682,N_2046,N_2489);
or U2683 (N_2683,N_2320,N_2026);
nor U2684 (N_2684,N_2144,N_2250);
nand U2685 (N_2685,N_2495,N_2111);
nor U2686 (N_2686,N_2499,N_2137);
xnor U2687 (N_2687,N_2089,N_2401);
nor U2688 (N_2688,N_2023,N_2191);
and U2689 (N_2689,N_2390,N_2150);
or U2690 (N_2690,N_2045,N_2105);
xnor U2691 (N_2691,N_2426,N_2415);
nor U2692 (N_2692,N_2377,N_2007);
or U2693 (N_2693,N_2195,N_2054);
and U2694 (N_2694,N_2100,N_2281);
nor U2695 (N_2695,N_2073,N_2319);
nand U2696 (N_2696,N_2179,N_2185);
nand U2697 (N_2697,N_2094,N_2121);
and U2698 (N_2698,N_2084,N_2224);
xor U2699 (N_2699,N_2138,N_2459);
and U2700 (N_2700,N_2405,N_2016);
nand U2701 (N_2701,N_2349,N_2300);
and U2702 (N_2702,N_2202,N_2437);
nor U2703 (N_2703,N_2235,N_2228);
xor U2704 (N_2704,N_2363,N_2064);
nand U2705 (N_2705,N_2490,N_2217);
or U2706 (N_2706,N_2069,N_2232);
xor U2707 (N_2707,N_2123,N_2128);
and U2708 (N_2708,N_2267,N_2078);
or U2709 (N_2709,N_2322,N_2313);
and U2710 (N_2710,N_2431,N_2208);
nor U2711 (N_2711,N_2275,N_2408);
nand U2712 (N_2712,N_2258,N_2002);
and U2713 (N_2713,N_2060,N_2061);
nor U2714 (N_2714,N_2231,N_2071);
or U2715 (N_2715,N_2386,N_2146);
nand U2716 (N_2716,N_2188,N_2374);
nor U2717 (N_2717,N_2433,N_2156);
and U2718 (N_2718,N_2406,N_2460);
or U2719 (N_2719,N_2022,N_2328);
xor U2720 (N_2720,N_2245,N_2292);
nor U2721 (N_2721,N_2025,N_2019);
nor U2722 (N_2722,N_2230,N_2057);
or U2723 (N_2723,N_2279,N_2343);
nand U2724 (N_2724,N_2028,N_2482);
nor U2725 (N_2725,N_2198,N_2106);
and U2726 (N_2726,N_2376,N_2177);
and U2727 (N_2727,N_2280,N_2334);
xnor U2728 (N_2728,N_2269,N_2068);
or U2729 (N_2729,N_2243,N_2496);
nor U2730 (N_2730,N_2141,N_2432);
nor U2731 (N_2731,N_2255,N_2139);
and U2732 (N_2732,N_2159,N_2081);
or U2733 (N_2733,N_2196,N_2317);
or U2734 (N_2734,N_2058,N_2037);
and U2735 (N_2735,N_2412,N_2316);
and U2736 (N_2736,N_2304,N_2148);
nand U2737 (N_2737,N_2403,N_2413);
nand U2738 (N_2738,N_2370,N_2169);
and U2739 (N_2739,N_2213,N_2063);
nor U2740 (N_2740,N_2108,N_2011);
nor U2741 (N_2741,N_2168,N_2133);
and U2742 (N_2742,N_2238,N_2052);
and U2743 (N_2743,N_2233,N_2326);
or U2744 (N_2744,N_2038,N_2331);
and U2745 (N_2745,N_2341,N_2091);
nor U2746 (N_2746,N_2457,N_2397);
and U2747 (N_2747,N_2263,N_2318);
or U2748 (N_2748,N_2463,N_2056);
and U2749 (N_2749,N_2214,N_2288);
nand U2750 (N_2750,N_2476,N_2239);
nand U2751 (N_2751,N_2446,N_2298);
nand U2752 (N_2752,N_2402,N_2453);
and U2753 (N_2753,N_2414,N_2434);
or U2754 (N_2754,N_2432,N_2252);
nor U2755 (N_2755,N_2120,N_2220);
nand U2756 (N_2756,N_2409,N_2380);
and U2757 (N_2757,N_2453,N_2215);
xor U2758 (N_2758,N_2479,N_2492);
or U2759 (N_2759,N_2198,N_2350);
nor U2760 (N_2760,N_2440,N_2229);
or U2761 (N_2761,N_2291,N_2053);
and U2762 (N_2762,N_2294,N_2318);
and U2763 (N_2763,N_2043,N_2446);
nand U2764 (N_2764,N_2335,N_2400);
nor U2765 (N_2765,N_2421,N_2320);
or U2766 (N_2766,N_2414,N_2348);
nand U2767 (N_2767,N_2079,N_2233);
nor U2768 (N_2768,N_2363,N_2196);
nand U2769 (N_2769,N_2268,N_2328);
xnor U2770 (N_2770,N_2443,N_2157);
nand U2771 (N_2771,N_2103,N_2023);
and U2772 (N_2772,N_2457,N_2400);
nand U2773 (N_2773,N_2215,N_2065);
and U2774 (N_2774,N_2334,N_2406);
or U2775 (N_2775,N_2076,N_2124);
nor U2776 (N_2776,N_2427,N_2376);
or U2777 (N_2777,N_2140,N_2459);
xnor U2778 (N_2778,N_2205,N_2292);
nor U2779 (N_2779,N_2314,N_2019);
or U2780 (N_2780,N_2055,N_2408);
nand U2781 (N_2781,N_2349,N_2342);
xor U2782 (N_2782,N_2461,N_2418);
nand U2783 (N_2783,N_2231,N_2485);
nand U2784 (N_2784,N_2081,N_2244);
nand U2785 (N_2785,N_2112,N_2292);
xnor U2786 (N_2786,N_2390,N_2122);
nand U2787 (N_2787,N_2423,N_2185);
or U2788 (N_2788,N_2495,N_2003);
nor U2789 (N_2789,N_2076,N_2043);
and U2790 (N_2790,N_2272,N_2251);
or U2791 (N_2791,N_2059,N_2153);
and U2792 (N_2792,N_2327,N_2428);
xnor U2793 (N_2793,N_2241,N_2211);
nand U2794 (N_2794,N_2040,N_2359);
and U2795 (N_2795,N_2302,N_2354);
xor U2796 (N_2796,N_2238,N_2478);
or U2797 (N_2797,N_2306,N_2035);
or U2798 (N_2798,N_2457,N_2490);
xor U2799 (N_2799,N_2025,N_2477);
nand U2800 (N_2800,N_2434,N_2212);
nand U2801 (N_2801,N_2161,N_2009);
nand U2802 (N_2802,N_2247,N_2427);
nor U2803 (N_2803,N_2229,N_2226);
xor U2804 (N_2804,N_2010,N_2060);
nand U2805 (N_2805,N_2301,N_2078);
or U2806 (N_2806,N_2403,N_2463);
or U2807 (N_2807,N_2078,N_2190);
nand U2808 (N_2808,N_2235,N_2406);
and U2809 (N_2809,N_2442,N_2252);
nor U2810 (N_2810,N_2410,N_2298);
nor U2811 (N_2811,N_2301,N_2426);
and U2812 (N_2812,N_2265,N_2187);
nor U2813 (N_2813,N_2238,N_2236);
or U2814 (N_2814,N_2452,N_2280);
nand U2815 (N_2815,N_2197,N_2417);
nor U2816 (N_2816,N_2060,N_2160);
or U2817 (N_2817,N_2194,N_2213);
nand U2818 (N_2818,N_2182,N_2459);
or U2819 (N_2819,N_2462,N_2102);
and U2820 (N_2820,N_2345,N_2270);
nand U2821 (N_2821,N_2136,N_2186);
nor U2822 (N_2822,N_2230,N_2050);
or U2823 (N_2823,N_2346,N_2244);
nand U2824 (N_2824,N_2415,N_2380);
and U2825 (N_2825,N_2381,N_2448);
xor U2826 (N_2826,N_2075,N_2086);
xnor U2827 (N_2827,N_2084,N_2195);
and U2828 (N_2828,N_2321,N_2138);
xnor U2829 (N_2829,N_2143,N_2319);
nand U2830 (N_2830,N_2099,N_2102);
and U2831 (N_2831,N_2179,N_2113);
nand U2832 (N_2832,N_2405,N_2071);
nand U2833 (N_2833,N_2132,N_2333);
xor U2834 (N_2834,N_2031,N_2119);
xnor U2835 (N_2835,N_2312,N_2192);
nor U2836 (N_2836,N_2198,N_2398);
nor U2837 (N_2837,N_2095,N_2213);
nand U2838 (N_2838,N_2443,N_2468);
nand U2839 (N_2839,N_2196,N_2284);
nor U2840 (N_2840,N_2157,N_2291);
and U2841 (N_2841,N_2027,N_2464);
nor U2842 (N_2842,N_2257,N_2174);
and U2843 (N_2843,N_2159,N_2154);
xnor U2844 (N_2844,N_2276,N_2441);
nand U2845 (N_2845,N_2152,N_2062);
nand U2846 (N_2846,N_2064,N_2051);
and U2847 (N_2847,N_2385,N_2231);
xnor U2848 (N_2848,N_2101,N_2360);
and U2849 (N_2849,N_2300,N_2245);
and U2850 (N_2850,N_2103,N_2035);
nand U2851 (N_2851,N_2458,N_2185);
nand U2852 (N_2852,N_2102,N_2422);
and U2853 (N_2853,N_2401,N_2009);
nor U2854 (N_2854,N_2360,N_2387);
or U2855 (N_2855,N_2055,N_2288);
xor U2856 (N_2856,N_2470,N_2238);
nand U2857 (N_2857,N_2075,N_2386);
xor U2858 (N_2858,N_2000,N_2107);
and U2859 (N_2859,N_2088,N_2256);
nor U2860 (N_2860,N_2069,N_2014);
nand U2861 (N_2861,N_2467,N_2493);
or U2862 (N_2862,N_2361,N_2045);
nor U2863 (N_2863,N_2060,N_2250);
or U2864 (N_2864,N_2475,N_2455);
or U2865 (N_2865,N_2406,N_2279);
nand U2866 (N_2866,N_2222,N_2278);
nand U2867 (N_2867,N_2111,N_2350);
nor U2868 (N_2868,N_2165,N_2237);
xnor U2869 (N_2869,N_2320,N_2306);
nor U2870 (N_2870,N_2210,N_2248);
nor U2871 (N_2871,N_2036,N_2315);
xor U2872 (N_2872,N_2200,N_2311);
xnor U2873 (N_2873,N_2351,N_2499);
nor U2874 (N_2874,N_2054,N_2369);
nor U2875 (N_2875,N_2166,N_2351);
or U2876 (N_2876,N_2431,N_2090);
nand U2877 (N_2877,N_2122,N_2202);
xnor U2878 (N_2878,N_2096,N_2098);
nor U2879 (N_2879,N_2058,N_2445);
and U2880 (N_2880,N_2281,N_2033);
nor U2881 (N_2881,N_2096,N_2399);
nand U2882 (N_2882,N_2036,N_2173);
nor U2883 (N_2883,N_2012,N_2005);
nor U2884 (N_2884,N_2100,N_2406);
and U2885 (N_2885,N_2407,N_2452);
or U2886 (N_2886,N_2034,N_2491);
and U2887 (N_2887,N_2214,N_2306);
nor U2888 (N_2888,N_2497,N_2369);
nand U2889 (N_2889,N_2375,N_2172);
and U2890 (N_2890,N_2145,N_2289);
nor U2891 (N_2891,N_2121,N_2265);
and U2892 (N_2892,N_2332,N_2164);
nor U2893 (N_2893,N_2082,N_2423);
and U2894 (N_2894,N_2067,N_2143);
or U2895 (N_2895,N_2143,N_2084);
and U2896 (N_2896,N_2140,N_2480);
and U2897 (N_2897,N_2416,N_2471);
and U2898 (N_2898,N_2097,N_2379);
and U2899 (N_2899,N_2134,N_2351);
nand U2900 (N_2900,N_2311,N_2100);
and U2901 (N_2901,N_2097,N_2123);
nand U2902 (N_2902,N_2049,N_2496);
or U2903 (N_2903,N_2445,N_2371);
and U2904 (N_2904,N_2162,N_2140);
nor U2905 (N_2905,N_2064,N_2392);
or U2906 (N_2906,N_2136,N_2392);
or U2907 (N_2907,N_2149,N_2094);
nor U2908 (N_2908,N_2018,N_2428);
or U2909 (N_2909,N_2078,N_2069);
and U2910 (N_2910,N_2096,N_2383);
nand U2911 (N_2911,N_2287,N_2058);
or U2912 (N_2912,N_2232,N_2185);
or U2913 (N_2913,N_2188,N_2205);
nand U2914 (N_2914,N_2252,N_2278);
xor U2915 (N_2915,N_2173,N_2468);
and U2916 (N_2916,N_2275,N_2371);
and U2917 (N_2917,N_2072,N_2289);
and U2918 (N_2918,N_2194,N_2322);
and U2919 (N_2919,N_2092,N_2271);
or U2920 (N_2920,N_2032,N_2392);
nor U2921 (N_2921,N_2008,N_2477);
and U2922 (N_2922,N_2175,N_2262);
nand U2923 (N_2923,N_2060,N_2040);
and U2924 (N_2924,N_2064,N_2373);
and U2925 (N_2925,N_2375,N_2113);
nor U2926 (N_2926,N_2435,N_2197);
nand U2927 (N_2927,N_2138,N_2067);
xnor U2928 (N_2928,N_2010,N_2396);
or U2929 (N_2929,N_2322,N_2273);
nor U2930 (N_2930,N_2164,N_2351);
xnor U2931 (N_2931,N_2370,N_2215);
nand U2932 (N_2932,N_2317,N_2075);
nor U2933 (N_2933,N_2470,N_2343);
nor U2934 (N_2934,N_2477,N_2269);
and U2935 (N_2935,N_2135,N_2085);
nor U2936 (N_2936,N_2400,N_2148);
nor U2937 (N_2937,N_2096,N_2375);
and U2938 (N_2938,N_2005,N_2483);
nand U2939 (N_2939,N_2123,N_2027);
and U2940 (N_2940,N_2362,N_2108);
nand U2941 (N_2941,N_2116,N_2207);
or U2942 (N_2942,N_2246,N_2262);
nand U2943 (N_2943,N_2210,N_2149);
nor U2944 (N_2944,N_2226,N_2281);
xor U2945 (N_2945,N_2145,N_2043);
nor U2946 (N_2946,N_2225,N_2348);
nor U2947 (N_2947,N_2222,N_2410);
or U2948 (N_2948,N_2303,N_2121);
nor U2949 (N_2949,N_2254,N_2141);
and U2950 (N_2950,N_2251,N_2325);
nand U2951 (N_2951,N_2327,N_2223);
and U2952 (N_2952,N_2342,N_2486);
and U2953 (N_2953,N_2414,N_2265);
and U2954 (N_2954,N_2117,N_2229);
and U2955 (N_2955,N_2270,N_2222);
nor U2956 (N_2956,N_2475,N_2110);
and U2957 (N_2957,N_2408,N_2157);
nand U2958 (N_2958,N_2181,N_2331);
or U2959 (N_2959,N_2426,N_2314);
nand U2960 (N_2960,N_2282,N_2233);
or U2961 (N_2961,N_2122,N_2119);
or U2962 (N_2962,N_2090,N_2251);
and U2963 (N_2963,N_2497,N_2391);
or U2964 (N_2964,N_2396,N_2420);
and U2965 (N_2965,N_2241,N_2016);
nor U2966 (N_2966,N_2056,N_2242);
or U2967 (N_2967,N_2226,N_2453);
and U2968 (N_2968,N_2210,N_2478);
or U2969 (N_2969,N_2484,N_2218);
or U2970 (N_2970,N_2190,N_2419);
nand U2971 (N_2971,N_2135,N_2475);
and U2972 (N_2972,N_2352,N_2425);
nand U2973 (N_2973,N_2207,N_2246);
nor U2974 (N_2974,N_2194,N_2352);
nand U2975 (N_2975,N_2486,N_2366);
and U2976 (N_2976,N_2300,N_2400);
nor U2977 (N_2977,N_2106,N_2125);
or U2978 (N_2978,N_2333,N_2054);
or U2979 (N_2979,N_2128,N_2214);
and U2980 (N_2980,N_2078,N_2074);
and U2981 (N_2981,N_2024,N_2139);
or U2982 (N_2982,N_2149,N_2117);
xor U2983 (N_2983,N_2340,N_2418);
and U2984 (N_2984,N_2095,N_2372);
nand U2985 (N_2985,N_2420,N_2054);
or U2986 (N_2986,N_2420,N_2273);
or U2987 (N_2987,N_2344,N_2079);
nor U2988 (N_2988,N_2313,N_2289);
nand U2989 (N_2989,N_2213,N_2416);
or U2990 (N_2990,N_2036,N_2009);
and U2991 (N_2991,N_2028,N_2456);
nand U2992 (N_2992,N_2411,N_2030);
or U2993 (N_2993,N_2127,N_2075);
and U2994 (N_2994,N_2387,N_2410);
nor U2995 (N_2995,N_2179,N_2199);
nand U2996 (N_2996,N_2079,N_2189);
and U2997 (N_2997,N_2107,N_2450);
nand U2998 (N_2998,N_2000,N_2231);
nand U2999 (N_2999,N_2414,N_2254);
and U3000 (N_3000,N_2628,N_2906);
and U3001 (N_3001,N_2884,N_2699);
xor U3002 (N_3002,N_2659,N_2950);
and U3003 (N_3003,N_2820,N_2704);
and U3004 (N_3004,N_2517,N_2814);
xor U3005 (N_3005,N_2744,N_2991);
or U3006 (N_3006,N_2822,N_2911);
nor U3007 (N_3007,N_2904,N_2660);
or U3008 (N_3008,N_2552,N_2637);
or U3009 (N_3009,N_2989,N_2858);
and U3010 (N_3010,N_2752,N_2874);
and U3011 (N_3011,N_2903,N_2706);
nand U3012 (N_3012,N_2936,N_2502);
nand U3013 (N_3013,N_2937,N_2738);
xor U3014 (N_3014,N_2898,N_2784);
nor U3015 (N_3015,N_2540,N_2748);
or U3016 (N_3016,N_2917,N_2916);
or U3017 (N_3017,N_2657,N_2568);
nand U3018 (N_3018,N_2509,N_2798);
nor U3019 (N_3019,N_2598,N_2849);
and U3020 (N_3020,N_2982,N_2740);
nand U3021 (N_3021,N_2875,N_2840);
nor U3022 (N_3022,N_2958,N_2526);
and U3023 (N_3023,N_2632,N_2556);
nor U3024 (N_3024,N_2500,N_2975);
xnor U3025 (N_3025,N_2577,N_2834);
or U3026 (N_3026,N_2787,N_2978);
and U3027 (N_3027,N_2739,N_2501);
xnor U3028 (N_3028,N_2804,N_2909);
or U3029 (N_3029,N_2747,N_2690);
nor U3030 (N_3030,N_2569,N_2731);
or U3031 (N_3031,N_2924,N_2675);
nor U3032 (N_3032,N_2576,N_2710);
or U3033 (N_3033,N_2715,N_2691);
nand U3034 (N_3034,N_2730,N_2801);
nand U3035 (N_3035,N_2671,N_2745);
and U3036 (N_3036,N_2630,N_2932);
nand U3037 (N_3037,N_2976,N_2979);
or U3038 (N_3038,N_2702,N_2639);
and U3039 (N_3039,N_2726,N_2645);
nand U3040 (N_3040,N_2570,N_2993);
nor U3041 (N_3041,N_2929,N_2705);
nor U3042 (N_3042,N_2541,N_2532);
or U3043 (N_3043,N_2995,N_2635);
nor U3044 (N_3044,N_2922,N_2873);
nor U3045 (N_3045,N_2648,N_2537);
nor U3046 (N_3046,N_2890,N_2966);
and U3047 (N_3047,N_2667,N_2942);
or U3048 (N_3048,N_2828,N_2643);
and U3049 (N_3049,N_2689,N_2815);
nor U3050 (N_3050,N_2722,N_2845);
nor U3051 (N_3051,N_2528,N_2714);
nor U3052 (N_3052,N_2848,N_2921);
nor U3053 (N_3053,N_2865,N_2952);
and U3054 (N_3054,N_2510,N_2651);
nor U3055 (N_3055,N_2550,N_2939);
nand U3056 (N_3056,N_2998,N_2817);
and U3057 (N_3057,N_2585,N_2927);
xor U3058 (N_3058,N_2700,N_2616);
or U3059 (N_3059,N_2618,N_2905);
nand U3060 (N_3060,N_2928,N_2818);
nor U3061 (N_3061,N_2683,N_2985);
nand U3062 (N_3062,N_2824,N_2530);
or U3063 (N_3063,N_2833,N_2692);
xor U3064 (N_3064,N_2546,N_2943);
or U3065 (N_3065,N_2572,N_2771);
nand U3066 (N_3066,N_2694,N_2640);
or U3067 (N_3067,N_2767,N_2623);
nand U3068 (N_3068,N_2559,N_2600);
and U3069 (N_3069,N_2518,N_2819);
xor U3070 (N_3070,N_2592,N_2888);
nor U3071 (N_3071,N_2789,N_2987);
nor U3072 (N_3072,N_2565,N_2508);
nand U3073 (N_3073,N_2880,N_2506);
nand U3074 (N_3074,N_2580,N_2946);
nor U3075 (N_3075,N_2972,N_2595);
nor U3076 (N_3076,N_2954,N_2522);
and U3077 (N_3077,N_2653,N_2615);
nand U3078 (N_3078,N_2802,N_2594);
nor U3079 (N_3079,N_2753,N_2588);
and U3080 (N_3080,N_2548,N_2948);
or U3081 (N_3081,N_2586,N_2963);
or U3082 (N_3082,N_2866,N_2887);
nor U3083 (N_3083,N_2750,N_2854);
and U3084 (N_3084,N_2951,N_2792);
nor U3085 (N_3085,N_2727,N_2693);
or U3086 (N_3086,N_2587,N_2621);
or U3087 (N_3087,N_2807,N_2770);
and U3088 (N_3088,N_2918,N_2596);
and U3089 (N_3089,N_2797,N_2581);
and U3090 (N_3090,N_2538,N_2533);
or U3091 (N_3091,N_2733,N_2915);
or U3092 (N_3092,N_2564,N_2677);
nand U3093 (N_3093,N_2647,N_2758);
or U3094 (N_3094,N_2754,N_2799);
and U3095 (N_3095,N_2644,N_2732);
or U3096 (N_3096,N_2925,N_2876);
nor U3097 (N_3097,N_2881,N_2670);
or U3098 (N_3098,N_2949,N_2892);
and U3099 (N_3099,N_2923,N_2878);
and U3100 (N_3100,N_2703,N_2973);
or U3101 (N_3101,N_2725,N_2549);
nor U3102 (N_3102,N_2841,N_2527);
and U3103 (N_3103,N_2934,N_2698);
and U3104 (N_3104,N_2764,N_2761);
nor U3105 (N_3105,N_2786,N_2806);
or U3106 (N_3106,N_2696,N_2762);
xnor U3107 (N_3107,N_2811,N_2713);
nand U3108 (N_3108,N_2859,N_2981);
nor U3109 (N_3109,N_2626,N_2781);
and U3110 (N_3110,N_2553,N_2503);
or U3111 (N_3111,N_2602,N_2894);
and U3112 (N_3112,N_2523,N_2825);
or U3113 (N_3113,N_2955,N_2529);
nor U3114 (N_3114,N_2856,N_2590);
or U3115 (N_3115,N_2908,N_2629);
xnor U3116 (N_3116,N_2558,N_2772);
and U3117 (N_3117,N_2531,N_2913);
nor U3118 (N_3118,N_2920,N_2901);
or U3119 (N_3119,N_2962,N_2869);
or U3120 (N_3120,N_2519,N_2664);
nand U3121 (N_3121,N_2988,N_2777);
nor U3122 (N_3122,N_2843,N_2826);
or U3123 (N_3123,N_2844,N_2575);
nor U3124 (N_3124,N_2662,N_2994);
nor U3125 (N_3125,N_2851,N_2652);
nor U3126 (N_3126,N_2515,N_2610);
and U3127 (N_3127,N_2795,N_2864);
nor U3128 (N_3128,N_2763,N_2545);
or U3129 (N_3129,N_2718,N_2674);
nor U3130 (N_3130,N_2803,N_2885);
or U3131 (N_3131,N_2872,N_2682);
and U3132 (N_3132,N_2769,N_2665);
or U3133 (N_3133,N_2612,N_2709);
nand U3134 (N_3134,N_2959,N_2680);
nor U3135 (N_3135,N_2779,N_2708);
nand U3136 (N_3136,N_2766,N_2658);
nor U3137 (N_3137,N_2684,N_2735);
or U3138 (N_3138,N_2749,N_2614);
nor U3139 (N_3139,N_2810,N_2805);
nor U3140 (N_3140,N_2837,N_2832);
nor U3141 (N_3141,N_2861,N_2900);
or U3142 (N_3142,N_2775,N_2679);
and U3143 (N_3143,N_2571,N_2889);
and U3144 (N_3144,N_2838,N_2964);
nand U3145 (N_3145,N_2977,N_2794);
nor U3146 (N_3146,N_2953,N_2970);
and U3147 (N_3147,N_2721,N_2812);
or U3148 (N_3148,N_2584,N_2631);
xnor U3149 (N_3149,N_2542,N_2741);
and U3150 (N_3150,N_2808,N_2984);
nand U3151 (N_3151,N_2857,N_2839);
nor U3152 (N_3152,N_2716,N_2791);
or U3153 (N_3153,N_2724,N_2980);
or U3154 (N_3154,N_2543,N_2800);
nand U3155 (N_3155,N_2712,N_2609);
or U3156 (N_3156,N_2986,N_2737);
nand U3157 (N_3157,N_2768,N_2656);
nand U3158 (N_3158,N_2672,N_2778);
nor U3159 (N_3159,N_2871,N_2891);
xnor U3160 (N_3160,N_2697,N_2992);
nor U3161 (N_3161,N_2742,N_2863);
nor U3162 (N_3162,N_2646,N_2607);
or U3163 (N_3163,N_2847,N_2967);
or U3164 (N_3164,N_2695,N_2850);
and U3165 (N_3165,N_2926,N_2957);
nand U3166 (N_3166,N_2947,N_2636);
xor U3167 (N_3167,N_2971,N_2678);
nand U3168 (N_3168,N_2551,N_2830);
xnor U3169 (N_3169,N_2743,N_2574);
nor U3170 (N_3170,N_2676,N_2547);
or U3171 (N_3171,N_2886,N_2539);
and U3172 (N_3172,N_2896,N_2511);
nor U3173 (N_3173,N_2512,N_2711);
or U3174 (N_3174,N_2593,N_2617);
nand U3175 (N_3175,N_2835,N_2554);
or U3176 (N_3176,N_2960,N_2757);
nor U3177 (N_3177,N_2831,N_2965);
and U3178 (N_3178,N_2619,N_2782);
or U3179 (N_3179,N_2774,N_2899);
and U3180 (N_3180,N_2627,N_2605);
or U3181 (N_3181,N_2687,N_2686);
nand U3182 (N_3182,N_2821,N_2669);
nor U3183 (N_3183,N_2836,N_2760);
nor U3184 (N_3184,N_2912,N_2685);
xnor U3185 (N_3185,N_2728,N_2759);
nor U3186 (N_3186,N_2723,N_2793);
xnor U3187 (N_3187,N_2513,N_2613);
xor U3188 (N_3188,N_2827,N_2990);
and U3189 (N_3189,N_2666,N_2796);
nand U3190 (N_3190,N_2974,N_2661);
and U3191 (N_3191,N_2868,N_2983);
nand U3192 (N_3192,N_2930,N_2719);
or U3193 (N_3193,N_2536,N_2790);
xor U3194 (N_3194,N_2914,N_2641);
xor U3195 (N_3195,N_2938,N_2736);
nor U3196 (N_3196,N_2720,N_2622);
or U3197 (N_3197,N_2746,N_2562);
nand U3198 (N_3198,N_2624,N_2882);
nand U3199 (N_3199,N_2504,N_2608);
or U3200 (N_3200,N_2603,N_2919);
and U3201 (N_3201,N_2870,N_2582);
xnor U3202 (N_3202,N_2654,N_2649);
or U3203 (N_3203,N_2823,N_2877);
nand U3204 (N_3204,N_2668,N_2566);
and U3205 (N_3205,N_2809,N_2776);
and U3206 (N_3206,N_2935,N_2535);
or U3207 (N_3207,N_2895,N_2544);
or U3208 (N_3208,N_2707,N_2604);
nand U3209 (N_3209,N_2599,N_2583);
or U3210 (N_3210,N_2520,N_2561);
nand U3211 (N_3211,N_2783,N_2996);
or U3212 (N_3212,N_2573,N_2663);
nand U3213 (N_3213,N_2933,N_2852);
and U3214 (N_3214,N_2638,N_2525);
nor U3215 (N_3215,N_2961,N_2813);
or U3216 (N_3216,N_2842,N_2910);
or U3217 (N_3217,N_2944,N_2931);
and U3218 (N_3218,N_2765,N_2907);
or U3219 (N_3219,N_2853,N_2867);
nor U3220 (N_3220,N_2611,N_2557);
or U3221 (N_3221,N_2883,N_2945);
and U3222 (N_3222,N_2524,N_2729);
or U3223 (N_3223,N_2785,N_2507);
nand U3224 (N_3224,N_2620,N_2816);
or U3225 (N_3225,N_2591,N_2534);
and U3226 (N_3226,N_2846,N_2514);
nand U3227 (N_3227,N_2578,N_2999);
and U3228 (N_3228,N_2756,N_2521);
and U3229 (N_3229,N_2681,N_2940);
nand U3230 (N_3230,N_2563,N_2642);
and U3231 (N_3231,N_2941,N_2860);
or U3232 (N_3232,N_2780,N_2968);
and U3233 (N_3233,N_2751,N_2855);
nand U3234 (N_3234,N_2969,N_2893);
or U3235 (N_3235,N_2597,N_2788);
or U3236 (N_3236,N_2734,N_2589);
and U3237 (N_3237,N_2688,N_2634);
or U3238 (N_3238,N_2633,N_2879);
or U3239 (N_3239,N_2701,N_2625);
nor U3240 (N_3240,N_2560,N_2755);
xor U3241 (N_3241,N_2579,N_2601);
and U3242 (N_3242,N_2505,N_2606);
or U3243 (N_3243,N_2997,N_2956);
and U3244 (N_3244,N_2773,N_2673);
nor U3245 (N_3245,N_2902,N_2897);
nand U3246 (N_3246,N_2655,N_2555);
or U3247 (N_3247,N_2829,N_2650);
or U3248 (N_3248,N_2862,N_2516);
and U3249 (N_3249,N_2717,N_2567);
nand U3250 (N_3250,N_2508,N_2520);
xnor U3251 (N_3251,N_2512,N_2634);
nor U3252 (N_3252,N_2796,N_2652);
xnor U3253 (N_3253,N_2549,N_2819);
nor U3254 (N_3254,N_2808,N_2832);
and U3255 (N_3255,N_2622,N_2603);
nor U3256 (N_3256,N_2559,N_2501);
nand U3257 (N_3257,N_2839,N_2643);
or U3258 (N_3258,N_2987,N_2741);
or U3259 (N_3259,N_2845,N_2931);
xor U3260 (N_3260,N_2817,N_2577);
nor U3261 (N_3261,N_2617,N_2521);
and U3262 (N_3262,N_2745,N_2915);
nand U3263 (N_3263,N_2604,N_2834);
or U3264 (N_3264,N_2556,N_2624);
nor U3265 (N_3265,N_2783,N_2976);
or U3266 (N_3266,N_2651,N_2912);
nand U3267 (N_3267,N_2588,N_2952);
or U3268 (N_3268,N_2736,N_2692);
nand U3269 (N_3269,N_2582,N_2961);
and U3270 (N_3270,N_2695,N_2538);
xnor U3271 (N_3271,N_2972,N_2887);
nor U3272 (N_3272,N_2767,N_2608);
and U3273 (N_3273,N_2708,N_2608);
xor U3274 (N_3274,N_2583,N_2915);
or U3275 (N_3275,N_2736,N_2517);
nand U3276 (N_3276,N_2594,N_2670);
and U3277 (N_3277,N_2511,N_2813);
or U3278 (N_3278,N_2956,N_2623);
or U3279 (N_3279,N_2630,N_2825);
nor U3280 (N_3280,N_2715,N_2865);
xor U3281 (N_3281,N_2942,N_2977);
xnor U3282 (N_3282,N_2596,N_2570);
nand U3283 (N_3283,N_2868,N_2518);
xnor U3284 (N_3284,N_2638,N_2690);
and U3285 (N_3285,N_2574,N_2941);
or U3286 (N_3286,N_2597,N_2584);
nor U3287 (N_3287,N_2671,N_2509);
and U3288 (N_3288,N_2588,N_2558);
nand U3289 (N_3289,N_2652,N_2782);
or U3290 (N_3290,N_2678,N_2648);
or U3291 (N_3291,N_2559,N_2745);
and U3292 (N_3292,N_2850,N_2894);
and U3293 (N_3293,N_2743,N_2982);
nor U3294 (N_3294,N_2607,N_2721);
and U3295 (N_3295,N_2785,N_2677);
and U3296 (N_3296,N_2561,N_2867);
and U3297 (N_3297,N_2867,N_2603);
or U3298 (N_3298,N_2640,N_2502);
nand U3299 (N_3299,N_2525,N_2666);
or U3300 (N_3300,N_2579,N_2823);
or U3301 (N_3301,N_2610,N_2548);
and U3302 (N_3302,N_2952,N_2752);
nor U3303 (N_3303,N_2972,N_2590);
or U3304 (N_3304,N_2616,N_2949);
nand U3305 (N_3305,N_2629,N_2682);
or U3306 (N_3306,N_2669,N_2773);
and U3307 (N_3307,N_2809,N_2848);
and U3308 (N_3308,N_2731,N_2953);
and U3309 (N_3309,N_2629,N_2577);
or U3310 (N_3310,N_2631,N_2958);
nor U3311 (N_3311,N_2902,N_2542);
nand U3312 (N_3312,N_2542,N_2921);
nand U3313 (N_3313,N_2992,N_2618);
and U3314 (N_3314,N_2878,N_2638);
nor U3315 (N_3315,N_2518,N_2546);
or U3316 (N_3316,N_2667,N_2775);
and U3317 (N_3317,N_2728,N_2548);
and U3318 (N_3318,N_2516,N_2810);
nand U3319 (N_3319,N_2716,N_2822);
or U3320 (N_3320,N_2752,N_2902);
nand U3321 (N_3321,N_2616,N_2805);
or U3322 (N_3322,N_2942,N_2801);
and U3323 (N_3323,N_2677,N_2986);
nand U3324 (N_3324,N_2796,N_2636);
or U3325 (N_3325,N_2787,N_2908);
xor U3326 (N_3326,N_2993,N_2900);
nor U3327 (N_3327,N_2630,N_2896);
nor U3328 (N_3328,N_2889,N_2732);
and U3329 (N_3329,N_2543,N_2837);
nor U3330 (N_3330,N_2866,N_2847);
and U3331 (N_3331,N_2614,N_2829);
nor U3332 (N_3332,N_2671,N_2778);
or U3333 (N_3333,N_2746,N_2959);
nor U3334 (N_3334,N_2910,N_2505);
and U3335 (N_3335,N_2802,N_2935);
nand U3336 (N_3336,N_2934,N_2547);
or U3337 (N_3337,N_2748,N_2598);
nor U3338 (N_3338,N_2723,N_2855);
or U3339 (N_3339,N_2832,N_2822);
or U3340 (N_3340,N_2557,N_2914);
and U3341 (N_3341,N_2699,N_2986);
nor U3342 (N_3342,N_2629,N_2513);
nand U3343 (N_3343,N_2663,N_2895);
and U3344 (N_3344,N_2803,N_2897);
or U3345 (N_3345,N_2524,N_2736);
and U3346 (N_3346,N_2856,N_2861);
and U3347 (N_3347,N_2526,N_2581);
nor U3348 (N_3348,N_2798,N_2524);
and U3349 (N_3349,N_2732,N_2694);
xor U3350 (N_3350,N_2799,N_2682);
or U3351 (N_3351,N_2733,N_2603);
nand U3352 (N_3352,N_2632,N_2534);
and U3353 (N_3353,N_2567,N_2673);
xnor U3354 (N_3354,N_2787,N_2747);
nand U3355 (N_3355,N_2602,N_2768);
nand U3356 (N_3356,N_2540,N_2681);
and U3357 (N_3357,N_2735,N_2658);
or U3358 (N_3358,N_2955,N_2745);
nand U3359 (N_3359,N_2848,N_2898);
or U3360 (N_3360,N_2857,N_2637);
and U3361 (N_3361,N_2846,N_2760);
nand U3362 (N_3362,N_2674,N_2930);
nor U3363 (N_3363,N_2840,N_2987);
nand U3364 (N_3364,N_2554,N_2514);
or U3365 (N_3365,N_2769,N_2676);
xnor U3366 (N_3366,N_2992,N_2714);
and U3367 (N_3367,N_2545,N_2897);
nand U3368 (N_3368,N_2680,N_2937);
and U3369 (N_3369,N_2621,N_2575);
nand U3370 (N_3370,N_2562,N_2961);
or U3371 (N_3371,N_2701,N_2742);
and U3372 (N_3372,N_2681,N_2828);
xor U3373 (N_3373,N_2858,N_2648);
nor U3374 (N_3374,N_2544,N_2521);
or U3375 (N_3375,N_2608,N_2866);
nor U3376 (N_3376,N_2539,N_2608);
nor U3377 (N_3377,N_2843,N_2834);
nor U3378 (N_3378,N_2819,N_2645);
xor U3379 (N_3379,N_2600,N_2892);
nor U3380 (N_3380,N_2930,N_2871);
or U3381 (N_3381,N_2938,N_2588);
nor U3382 (N_3382,N_2617,N_2691);
or U3383 (N_3383,N_2728,N_2584);
and U3384 (N_3384,N_2622,N_2804);
nor U3385 (N_3385,N_2600,N_2851);
nor U3386 (N_3386,N_2656,N_2594);
nand U3387 (N_3387,N_2706,N_2686);
or U3388 (N_3388,N_2660,N_2790);
and U3389 (N_3389,N_2822,N_2684);
nor U3390 (N_3390,N_2572,N_2848);
or U3391 (N_3391,N_2635,N_2971);
nand U3392 (N_3392,N_2722,N_2775);
nor U3393 (N_3393,N_2717,N_2928);
nand U3394 (N_3394,N_2848,N_2847);
nor U3395 (N_3395,N_2748,N_2807);
nand U3396 (N_3396,N_2759,N_2537);
or U3397 (N_3397,N_2700,N_2580);
or U3398 (N_3398,N_2572,N_2781);
xor U3399 (N_3399,N_2584,N_2735);
nand U3400 (N_3400,N_2728,N_2581);
or U3401 (N_3401,N_2711,N_2515);
or U3402 (N_3402,N_2919,N_2673);
or U3403 (N_3403,N_2569,N_2597);
nor U3404 (N_3404,N_2688,N_2714);
xnor U3405 (N_3405,N_2572,N_2945);
nor U3406 (N_3406,N_2928,N_2588);
nor U3407 (N_3407,N_2997,N_2550);
or U3408 (N_3408,N_2773,N_2924);
xnor U3409 (N_3409,N_2749,N_2622);
nand U3410 (N_3410,N_2978,N_2651);
nand U3411 (N_3411,N_2932,N_2619);
nand U3412 (N_3412,N_2889,N_2549);
nor U3413 (N_3413,N_2902,N_2651);
and U3414 (N_3414,N_2745,N_2506);
nor U3415 (N_3415,N_2860,N_2576);
and U3416 (N_3416,N_2791,N_2719);
and U3417 (N_3417,N_2843,N_2551);
xnor U3418 (N_3418,N_2574,N_2603);
xor U3419 (N_3419,N_2893,N_2620);
or U3420 (N_3420,N_2544,N_2949);
nand U3421 (N_3421,N_2518,N_2931);
and U3422 (N_3422,N_2855,N_2742);
and U3423 (N_3423,N_2535,N_2746);
and U3424 (N_3424,N_2549,N_2751);
or U3425 (N_3425,N_2739,N_2668);
nor U3426 (N_3426,N_2896,N_2639);
or U3427 (N_3427,N_2809,N_2503);
nor U3428 (N_3428,N_2961,N_2579);
nand U3429 (N_3429,N_2816,N_2766);
or U3430 (N_3430,N_2728,N_2872);
or U3431 (N_3431,N_2611,N_2593);
and U3432 (N_3432,N_2809,N_2574);
and U3433 (N_3433,N_2822,N_2904);
nor U3434 (N_3434,N_2594,N_2699);
or U3435 (N_3435,N_2996,N_2507);
xor U3436 (N_3436,N_2822,N_2875);
and U3437 (N_3437,N_2531,N_2896);
xnor U3438 (N_3438,N_2806,N_2622);
or U3439 (N_3439,N_2561,N_2776);
nor U3440 (N_3440,N_2960,N_2696);
and U3441 (N_3441,N_2963,N_2739);
or U3442 (N_3442,N_2624,N_2831);
nor U3443 (N_3443,N_2630,N_2933);
or U3444 (N_3444,N_2886,N_2679);
nand U3445 (N_3445,N_2961,N_2640);
or U3446 (N_3446,N_2984,N_2694);
or U3447 (N_3447,N_2787,N_2911);
nand U3448 (N_3448,N_2700,N_2754);
xor U3449 (N_3449,N_2747,N_2952);
and U3450 (N_3450,N_2833,N_2756);
xnor U3451 (N_3451,N_2924,N_2568);
or U3452 (N_3452,N_2775,N_2964);
nor U3453 (N_3453,N_2818,N_2732);
nor U3454 (N_3454,N_2691,N_2748);
and U3455 (N_3455,N_2714,N_2780);
xnor U3456 (N_3456,N_2796,N_2805);
xnor U3457 (N_3457,N_2522,N_2795);
or U3458 (N_3458,N_2994,N_2651);
or U3459 (N_3459,N_2524,N_2868);
nor U3460 (N_3460,N_2803,N_2550);
and U3461 (N_3461,N_2603,N_2610);
and U3462 (N_3462,N_2883,N_2593);
nand U3463 (N_3463,N_2588,N_2660);
and U3464 (N_3464,N_2688,N_2815);
nand U3465 (N_3465,N_2911,N_2565);
or U3466 (N_3466,N_2537,N_2874);
or U3467 (N_3467,N_2777,N_2674);
nand U3468 (N_3468,N_2726,N_2737);
xor U3469 (N_3469,N_2584,N_2876);
nor U3470 (N_3470,N_2536,N_2781);
xor U3471 (N_3471,N_2704,N_2799);
and U3472 (N_3472,N_2974,N_2920);
or U3473 (N_3473,N_2590,N_2835);
and U3474 (N_3474,N_2581,N_2887);
nand U3475 (N_3475,N_2709,N_2762);
nand U3476 (N_3476,N_2843,N_2521);
and U3477 (N_3477,N_2617,N_2924);
nor U3478 (N_3478,N_2673,N_2690);
and U3479 (N_3479,N_2834,N_2531);
or U3480 (N_3480,N_2924,N_2789);
nor U3481 (N_3481,N_2795,N_2885);
nor U3482 (N_3482,N_2694,N_2724);
and U3483 (N_3483,N_2962,N_2819);
or U3484 (N_3484,N_2860,N_2899);
nor U3485 (N_3485,N_2543,N_2869);
or U3486 (N_3486,N_2978,N_2920);
nand U3487 (N_3487,N_2994,N_2515);
xor U3488 (N_3488,N_2763,N_2857);
nor U3489 (N_3489,N_2928,N_2842);
nand U3490 (N_3490,N_2949,N_2509);
or U3491 (N_3491,N_2510,N_2623);
nor U3492 (N_3492,N_2970,N_2534);
xor U3493 (N_3493,N_2749,N_2906);
nor U3494 (N_3494,N_2751,N_2613);
or U3495 (N_3495,N_2677,N_2532);
xnor U3496 (N_3496,N_2822,N_2611);
or U3497 (N_3497,N_2626,N_2931);
nand U3498 (N_3498,N_2965,N_2744);
and U3499 (N_3499,N_2710,N_2984);
nor U3500 (N_3500,N_3215,N_3264);
or U3501 (N_3501,N_3296,N_3271);
or U3502 (N_3502,N_3431,N_3084);
nor U3503 (N_3503,N_3417,N_3237);
or U3504 (N_3504,N_3437,N_3408);
and U3505 (N_3505,N_3183,N_3198);
or U3506 (N_3506,N_3151,N_3163);
nand U3507 (N_3507,N_3260,N_3282);
nor U3508 (N_3508,N_3203,N_3101);
nand U3509 (N_3509,N_3221,N_3479);
nor U3510 (N_3510,N_3423,N_3470);
nor U3511 (N_3511,N_3441,N_3496);
nor U3512 (N_3512,N_3211,N_3145);
nor U3513 (N_3513,N_3097,N_3251);
xnor U3514 (N_3514,N_3140,N_3193);
nand U3515 (N_3515,N_3029,N_3337);
nor U3516 (N_3516,N_3034,N_3339);
or U3517 (N_3517,N_3332,N_3218);
nor U3518 (N_3518,N_3187,N_3227);
nor U3519 (N_3519,N_3273,N_3338);
or U3520 (N_3520,N_3471,N_3219);
and U3521 (N_3521,N_3000,N_3053);
nand U3522 (N_3522,N_3201,N_3344);
and U3523 (N_3523,N_3306,N_3095);
nor U3524 (N_3524,N_3166,N_3035);
and U3525 (N_3525,N_3388,N_3442);
nor U3526 (N_3526,N_3143,N_3284);
and U3527 (N_3527,N_3397,N_3064);
nor U3528 (N_3528,N_3148,N_3456);
nor U3529 (N_3529,N_3461,N_3204);
nand U3530 (N_3530,N_3077,N_3380);
nor U3531 (N_3531,N_3257,N_3155);
and U3532 (N_3532,N_3321,N_3027);
or U3533 (N_3533,N_3430,N_3214);
xor U3534 (N_3534,N_3454,N_3329);
or U3535 (N_3535,N_3233,N_3241);
and U3536 (N_3536,N_3112,N_3031);
and U3537 (N_3537,N_3007,N_3067);
and U3538 (N_3538,N_3010,N_3424);
or U3539 (N_3539,N_3243,N_3294);
nand U3540 (N_3540,N_3245,N_3407);
xnor U3541 (N_3541,N_3432,N_3150);
and U3542 (N_3542,N_3205,N_3421);
or U3543 (N_3543,N_3017,N_3371);
nor U3544 (N_3544,N_3301,N_3033);
nor U3545 (N_3545,N_3486,N_3307);
nor U3546 (N_3546,N_3037,N_3244);
or U3547 (N_3547,N_3351,N_3063);
nor U3548 (N_3548,N_3169,N_3355);
or U3549 (N_3549,N_3091,N_3116);
xnor U3550 (N_3550,N_3427,N_3314);
nand U3551 (N_3551,N_3179,N_3359);
or U3552 (N_3552,N_3391,N_3178);
and U3553 (N_3553,N_3292,N_3462);
or U3554 (N_3554,N_3360,N_3369);
nor U3555 (N_3555,N_3061,N_3220);
nand U3556 (N_3556,N_3117,N_3209);
nor U3557 (N_3557,N_3399,N_3104);
or U3558 (N_3558,N_3297,N_3485);
or U3559 (N_3559,N_3288,N_3176);
nand U3560 (N_3560,N_3015,N_3045);
xnor U3561 (N_3561,N_3256,N_3448);
nor U3562 (N_3562,N_3390,N_3483);
or U3563 (N_3563,N_3474,N_3457);
nor U3564 (N_3564,N_3139,N_3222);
nor U3565 (N_3565,N_3236,N_3181);
nor U3566 (N_3566,N_3372,N_3170);
or U3567 (N_3567,N_3363,N_3269);
and U3568 (N_3568,N_3270,N_3142);
and U3569 (N_3569,N_3006,N_3113);
nor U3570 (N_3570,N_3239,N_3100);
or U3571 (N_3571,N_3253,N_3223);
and U3572 (N_3572,N_3062,N_3090);
xnor U3573 (N_3573,N_3475,N_3291);
nand U3574 (N_3574,N_3242,N_3103);
or U3575 (N_3575,N_3048,N_3248);
or U3576 (N_3576,N_3184,N_3460);
nor U3577 (N_3577,N_3141,N_3032);
nand U3578 (N_3578,N_3429,N_3370);
nand U3579 (N_3579,N_3463,N_3055);
nand U3580 (N_3580,N_3394,N_3453);
nand U3581 (N_3581,N_3262,N_3386);
or U3582 (N_3582,N_3153,N_3316);
or U3583 (N_3583,N_3348,N_3322);
or U3584 (N_3584,N_3480,N_3309);
nand U3585 (N_3585,N_3452,N_3366);
nor U3586 (N_3586,N_3089,N_3225);
nor U3587 (N_3587,N_3477,N_3247);
nor U3588 (N_3588,N_3107,N_3287);
and U3589 (N_3589,N_3320,N_3347);
xor U3590 (N_3590,N_3235,N_3146);
and U3591 (N_3591,N_3384,N_3088);
and U3592 (N_3592,N_3466,N_3400);
and U3593 (N_3593,N_3435,N_3487);
nand U3594 (N_3594,N_3299,N_3058);
or U3595 (N_3595,N_3488,N_3418);
or U3596 (N_3596,N_3303,N_3134);
or U3597 (N_3597,N_3167,N_3491);
nor U3598 (N_3598,N_3382,N_3357);
and U3599 (N_3599,N_3364,N_3054);
or U3600 (N_3600,N_3272,N_3467);
and U3601 (N_3601,N_3118,N_3081);
nor U3602 (N_3602,N_3298,N_3121);
nor U3603 (N_3603,N_3172,N_3439);
nand U3604 (N_3604,N_3410,N_3376);
and U3605 (N_3605,N_3019,N_3468);
or U3606 (N_3606,N_3440,N_3356);
nor U3607 (N_3607,N_3072,N_3341);
nand U3608 (N_3608,N_3267,N_3494);
nor U3609 (N_3609,N_3276,N_3449);
or U3610 (N_3610,N_3379,N_3005);
or U3611 (N_3611,N_3075,N_3396);
xnor U3612 (N_3612,N_3030,N_3495);
nor U3613 (N_3613,N_3446,N_3459);
nor U3614 (N_3614,N_3076,N_3149);
nand U3615 (N_3615,N_3173,N_3069);
nand U3616 (N_3616,N_3250,N_3231);
nand U3617 (N_3617,N_3484,N_3039);
or U3618 (N_3618,N_3300,N_3229);
nor U3619 (N_3619,N_3174,N_3206);
nor U3620 (N_3620,N_3365,N_3493);
nand U3621 (N_3621,N_3079,N_3008);
nor U3622 (N_3622,N_3001,N_3464);
nor U3623 (N_3623,N_3157,N_3190);
nand U3624 (N_3624,N_3428,N_3336);
and U3625 (N_3625,N_3289,N_3111);
or U3626 (N_3626,N_3123,N_3207);
nand U3627 (N_3627,N_3040,N_3310);
or U3628 (N_3628,N_3425,N_3135);
and U3629 (N_3629,N_3416,N_3028);
nor U3630 (N_3630,N_3346,N_3415);
or U3631 (N_3631,N_3052,N_3189);
nor U3632 (N_3632,N_3185,N_3377);
and U3633 (N_3633,N_3051,N_3278);
nand U3634 (N_3634,N_3144,N_3059);
nor U3635 (N_3635,N_3004,N_3168);
and U3636 (N_3636,N_3354,N_3196);
xnor U3637 (N_3637,N_3108,N_3402);
and U3638 (N_3638,N_3406,N_3312);
xor U3639 (N_3639,N_3383,N_3180);
nand U3640 (N_3640,N_3188,N_3393);
and U3641 (N_3641,N_3258,N_3122);
and U3642 (N_3642,N_3340,N_3110);
nor U3643 (N_3643,N_3124,N_3274);
or U3644 (N_3644,N_3498,N_3451);
nor U3645 (N_3645,N_3130,N_3186);
and U3646 (N_3646,N_3411,N_3327);
nor U3647 (N_3647,N_3162,N_3492);
and U3648 (N_3648,N_3481,N_3044);
or U3649 (N_3649,N_3066,N_3208);
nand U3650 (N_3650,N_3389,N_3182);
or U3651 (N_3651,N_3131,N_3094);
or U3652 (N_3652,N_3458,N_3074);
or U3653 (N_3653,N_3313,N_3216);
nor U3654 (N_3654,N_3362,N_3401);
or U3655 (N_3655,N_3109,N_3436);
nand U3656 (N_3656,N_3318,N_3068);
or U3657 (N_3657,N_3082,N_3246);
and U3658 (N_3658,N_3023,N_3367);
and U3659 (N_3659,N_3129,N_3385);
or U3660 (N_3660,N_3087,N_3102);
nor U3661 (N_3661,N_3345,N_3057);
nor U3662 (N_3662,N_3036,N_3083);
nand U3663 (N_3663,N_3020,N_3434);
xnor U3664 (N_3664,N_3154,N_3137);
nand U3665 (N_3665,N_3445,N_3280);
nor U3666 (N_3666,N_3342,N_3078);
or U3667 (N_3667,N_3330,N_3419);
or U3668 (N_3668,N_3350,N_3002);
xor U3669 (N_3669,N_3093,N_3443);
and U3670 (N_3670,N_3497,N_3240);
nor U3671 (N_3671,N_3455,N_3252);
xor U3672 (N_3672,N_3217,N_3080);
xor U3673 (N_3673,N_3478,N_3197);
and U3674 (N_3674,N_3293,N_3047);
nor U3675 (N_3675,N_3194,N_3343);
nand U3676 (N_3676,N_3210,N_3368);
or U3677 (N_3677,N_3433,N_3473);
nand U3678 (N_3678,N_3404,N_3275);
or U3679 (N_3679,N_3334,N_3073);
xor U3680 (N_3680,N_3331,N_3308);
nand U3681 (N_3681,N_3476,N_3192);
and U3682 (N_3682,N_3147,N_3041);
nand U3683 (N_3683,N_3138,N_3106);
nand U3684 (N_3684,N_3119,N_3302);
nand U3685 (N_3685,N_3200,N_3403);
nor U3686 (N_3686,N_3482,N_3305);
or U3687 (N_3687,N_3114,N_3230);
xor U3688 (N_3688,N_3213,N_3042);
or U3689 (N_3689,N_3447,N_3115);
and U3690 (N_3690,N_3268,N_3426);
and U3691 (N_3691,N_3228,N_3085);
nand U3692 (N_3692,N_3128,N_3286);
nand U3693 (N_3693,N_3013,N_3071);
nor U3694 (N_3694,N_3398,N_3164);
nand U3695 (N_3695,N_3259,N_3158);
nor U3696 (N_3696,N_3304,N_3191);
nand U3697 (N_3697,N_3092,N_3324);
or U3698 (N_3698,N_3490,N_3133);
and U3699 (N_3699,N_3277,N_3352);
and U3700 (N_3700,N_3009,N_3056);
nor U3701 (N_3701,N_3127,N_3249);
and U3702 (N_3702,N_3472,N_3254);
xor U3703 (N_3703,N_3469,N_3171);
or U3704 (N_3704,N_3333,N_3202);
or U3705 (N_3705,N_3387,N_3070);
and U3706 (N_3706,N_3050,N_3226);
nor U3707 (N_3707,N_3049,N_3412);
or U3708 (N_3708,N_3152,N_3358);
nand U3709 (N_3709,N_3317,N_3392);
nor U3710 (N_3710,N_3018,N_3160);
and U3711 (N_3711,N_3136,N_3025);
and U3712 (N_3712,N_3311,N_3420);
and U3713 (N_3713,N_3295,N_3011);
xnor U3714 (N_3714,N_3234,N_3065);
xnor U3715 (N_3715,N_3323,N_3328);
nor U3716 (N_3716,N_3413,N_3465);
xnor U3717 (N_3717,N_3224,N_3098);
and U3718 (N_3718,N_3012,N_3021);
xor U3719 (N_3719,N_3285,N_3026);
or U3720 (N_3720,N_3265,N_3126);
nor U3721 (N_3721,N_3099,N_3444);
nand U3722 (N_3722,N_3279,N_3060);
nand U3723 (N_3723,N_3353,N_3374);
and U3724 (N_3724,N_3014,N_3395);
nand U3725 (N_3725,N_3238,N_3375);
or U3726 (N_3726,N_3232,N_3335);
nor U3727 (N_3727,N_3022,N_3489);
nor U3728 (N_3728,N_3175,N_3038);
xnor U3729 (N_3729,N_3043,N_3016);
nor U3730 (N_3730,N_3105,N_3361);
or U3731 (N_3731,N_3326,N_3261);
and U3732 (N_3732,N_3438,N_3378);
xnor U3733 (N_3733,N_3156,N_3381);
or U3734 (N_3734,N_3281,N_3086);
and U3735 (N_3735,N_3409,N_3125);
nor U3736 (N_3736,N_3263,N_3132);
nand U3737 (N_3737,N_3177,N_3159);
nor U3738 (N_3738,N_3450,N_3414);
nand U3739 (N_3739,N_3195,N_3046);
or U3740 (N_3740,N_3319,N_3255);
and U3741 (N_3741,N_3373,N_3290);
and U3742 (N_3742,N_3499,N_3315);
xor U3743 (N_3743,N_3325,N_3212);
nand U3744 (N_3744,N_3003,N_3120);
nand U3745 (N_3745,N_3199,N_3266);
or U3746 (N_3746,N_3024,N_3405);
and U3747 (N_3747,N_3165,N_3349);
nor U3748 (N_3748,N_3283,N_3422);
nand U3749 (N_3749,N_3161,N_3096);
or U3750 (N_3750,N_3025,N_3081);
or U3751 (N_3751,N_3444,N_3057);
nand U3752 (N_3752,N_3157,N_3098);
nor U3753 (N_3753,N_3491,N_3473);
nor U3754 (N_3754,N_3407,N_3128);
or U3755 (N_3755,N_3083,N_3177);
and U3756 (N_3756,N_3295,N_3202);
and U3757 (N_3757,N_3379,N_3364);
and U3758 (N_3758,N_3326,N_3235);
or U3759 (N_3759,N_3438,N_3103);
or U3760 (N_3760,N_3313,N_3308);
and U3761 (N_3761,N_3304,N_3234);
or U3762 (N_3762,N_3485,N_3325);
or U3763 (N_3763,N_3214,N_3325);
nand U3764 (N_3764,N_3026,N_3212);
nand U3765 (N_3765,N_3409,N_3181);
nand U3766 (N_3766,N_3357,N_3400);
and U3767 (N_3767,N_3359,N_3067);
xnor U3768 (N_3768,N_3196,N_3170);
nor U3769 (N_3769,N_3187,N_3034);
nand U3770 (N_3770,N_3291,N_3270);
and U3771 (N_3771,N_3213,N_3321);
xnor U3772 (N_3772,N_3285,N_3151);
and U3773 (N_3773,N_3407,N_3376);
nand U3774 (N_3774,N_3379,N_3339);
xor U3775 (N_3775,N_3486,N_3095);
nor U3776 (N_3776,N_3012,N_3270);
xor U3777 (N_3777,N_3241,N_3414);
xnor U3778 (N_3778,N_3182,N_3364);
and U3779 (N_3779,N_3355,N_3125);
nor U3780 (N_3780,N_3058,N_3036);
nor U3781 (N_3781,N_3012,N_3314);
nor U3782 (N_3782,N_3443,N_3407);
nor U3783 (N_3783,N_3135,N_3298);
xor U3784 (N_3784,N_3215,N_3277);
nand U3785 (N_3785,N_3220,N_3418);
and U3786 (N_3786,N_3492,N_3409);
nand U3787 (N_3787,N_3415,N_3111);
nand U3788 (N_3788,N_3345,N_3261);
or U3789 (N_3789,N_3161,N_3166);
nor U3790 (N_3790,N_3110,N_3450);
nand U3791 (N_3791,N_3186,N_3305);
nand U3792 (N_3792,N_3461,N_3492);
and U3793 (N_3793,N_3067,N_3152);
nand U3794 (N_3794,N_3281,N_3208);
or U3795 (N_3795,N_3347,N_3496);
or U3796 (N_3796,N_3144,N_3015);
or U3797 (N_3797,N_3265,N_3095);
xnor U3798 (N_3798,N_3143,N_3370);
nand U3799 (N_3799,N_3053,N_3410);
xnor U3800 (N_3800,N_3002,N_3085);
xnor U3801 (N_3801,N_3078,N_3100);
and U3802 (N_3802,N_3198,N_3350);
and U3803 (N_3803,N_3398,N_3178);
nand U3804 (N_3804,N_3483,N_3259);
nor U3805 (N_3805,N_3162,N_3158);
nor U3806 (N_3806,N_3288,N_3399);
and U3807 (N_3807,N_3037,N_3495);
or U3808 (N_3808,N_3242,N_3464);
xnor U3809 (N_3809,N_3140,N_3328);
and U3810 (N_3810,N_3330,N_3283);
nand U3811 (N_3811,N_3147,N_3346);
nor U3812 (N_3812,N_3347,N_3055);
and U3813 (N_3813,N_3412,N_3241);
nor U3814 (N_3814,N_3007,N_3084);
or U3815 (N_3815,N_3247,N_3050);
or U3816 (N_3816,N_3135,N_3000);
and U3817 (N_3817,N_3485,N_3015);
nor U3818 (N_3818,N_3430,N_3443);
or U3819 (N_3819,N_3253,N_3446);
xor U3820 (N_3820,N_3414,N_3294);
nand U3821 (N_3821,N_3256,N_3209);
nor U3822 (N_3822,N_3192,N_3277);
xor U3823 (N_3823,N_3370,N_3202);
or U3824 (N_3824,N_3439,N_3006);
and U3825 (N_3825,N_3438,N_3122);
and U3826 (N_3826,N_3137,N_3499);
and U3827 (N_3827,N_3419,N_3427);
and U3828 (N_3828,N_3451,N_3190);
nand U3829 (N_3829,N_3409,N_3206);
or U3830 (N_3830,N_3395,N_3479);
nor U3831 (N_3831,N_3084,N_3262);
nand U3832 (N_3832,N_3232,N_3401);
xor U3833 (N_3833,N_3086,N_3067);
nand U3834 (N_3834,N_3051,N_3481);
nand U3835 (N_3835,N_3079,N_3412);
or U3836 (N_3836,N_3386,N_3043);
and U3837 (N_3837,N_3349,N_3151);
and U3838 (N_3838,N_3475,N_3084);
nand U3839 (N_3839,N_3019,N_3107);
nor U3840 (N_3840,N_3470,N_3104);
and U3841 (N_3841,N_3219,N_3099);
and U3842 (N_3842,N_3095,N_3020);
nor U3843 (N_3843,N_3169,N_3099);
nor U3844 (N_3844,N_3089,N_3322);
or U3845 (N_3845,N_3106,N_3075);
and U3846 (N_3846,N_3007,N_3311);
and U3847 (N_3847,N_3449,N_3080);
or U3848 (N_3848,N_3021,N_3237);
nor U3849 (N_3849,N_3198,N_3481);
and U3850 (N_3850,N_3342,N_3414);
nand U3851 (N_3851,N_3100,N_3309);
nor U3852 (N_3852,N_3034,N_3214);
xor U3853 (N_3853,N_3132,N_3307);
and U3854 (N_3854,N_3164,N_3086);
and U3855 (N_3855,N_3137,N_3321);
nor U3856 (N_3856,N_3425,N_3363);
nor U3857 (N_3857,N_3044,N_3202);
xnor U3858 (N_3858,N_3379,N_3294);
nor U3859 (N_3859,N_3427,N_3027);
nand U3860 (N_3860,N_3090,N_3350);
nand U3861 (N_3861,N_3439,N_3309);
or U3862 (N_3862,N_3343,N_3240);
nand U3863 (N_3863,N_3326,N_3226);
and U3864 (N_3864,N_3435,N_3040);
nor U3865 (N_3865,N_3097,N_3318);
xor U3866 (N_3866,N_3464,N_3029);
or U3867 (N_3867,N_3381,N_3309);
or U3868 (N_3868,N_3134,N_3343);
nor U3869 (N_3869,N_3004,N_3131);
nor U3870 (N_3870,N_3461,N_3194);
and U3871 (N_3871,N_3049,N_3263);
and U3872 (N_3872,N_3211,N_3428);
or U3873 (N_3873,N_3431,N_3477);
nor U3874 (N_3874,N_3337,N_3382);
xnor U3875 (N_3875,N_3379,N_3332);
xor U3876 (N_3876,N_3219,N_3305);
nor U3877 (N_3877,N_3071,N_3312);
or U3878 (N_3878,N_3137,N_3169);
nor U3879 (N_3879,N_3180,N_3184);
or U3880 (N_3880,N_3320,N_3270);
or U3881 (N_3881,N_3229,N_3385);
and U3882 (N_3882,N_3118,N_3139);
nor U3883 (N_3883,N_3498,N_3232);
nand U3884 (N_3884,N_3193,N_3436);
nor U3885 (N_3885,N_3272,N_3018);
nor U3886 (N_3886,N_3240,N_3265);
nand U3887 (N_3887,N_3475,N_3426);
and U3888 (N_3888,N_3303,N_3239);
or U3889 (N_3889,N_3339,N_3164);
or U3890 (N_3890,N_3352,N_3385);
nand U3891 (N_3891,N_3332,N_3466);
xor U3892 (N_3892,N_3381,N_3124);
nand U3893 (N_3893,N_3176,N_3281);
and U3894 (N_3894,N_3220,N_3469);
nand U3895 (N_3895,N_3414,N_3054);
nor U3896 (N_3896,N_3129,N_3415);
and U3897 (N_3897,N_3354,N_3165);
nor U3898 (N_3898,N_3308,N_3450);
nor U3899 (N_3899,N_3494,N_3473);
or U3900 (N_3900,N_3417,N_3171);
or U3901 (N_3901,N_3366,N_3417);
nand U3902 (N_3902,N_3105,N_3455);
xor U3903 (N_3903,N_3118,N_3255);
and U3904 (N_3904,N_3263,N_3017);
nand U3905 (N_3905,N_3172,N_3424);
nor U3906 (N_3906,N_3481,N_3135);
nand U3907 (N_3907,N_3295,N_3495);
or U3908 (N_3908,N_3259,N_3154);
nand U3909 (N_3909,N_3479,N_3359);
nor U3910 (N_3910,N_3316,N_3367);
and U3911 (N_3911,N_3057,N_3077);
nand U3912 (N_3912,N_3115,N_3181);
nor U3913 (N_3913,N_3493,N_3071);
or U3914 (N_3914,N_3187,N_3237);
or U3915 (N_3915,N_3465,N_3016);
or U3916 (N_3916,N_3323,N_3473);
nor U3917 (N_3917,N_3391,N_3190);
or U3918 (N_3918,N_3456,N_3235);
nor U3919 (N_3919,N_3482,N_3468);
xor U3920 (N_3920,N_3378,N_3299);
or U3921 (N_3921,N_3383,N_3424);
nor U3922 (N_3922,N_3181,N_3481);
nand U3923 (N_3923,N_3183,N_3340);
and U3924 (N_3924,N_3063,N_3289);
nand U3925 (N_3925,N_3486,N_3084);
nor U3926 (N_3926,N_3213,N_3467);
nor U3927 (N_3927,N_3397,N_3255);
nand U3928 (N_3928,N_3460,N_3319);
nand U3929 (N_3929,N_3391,N_3455);
or U3930 (N_3930,N_3310,N_3261);
nand U3931 (N_3931,N_3360,N_3394);
xnor U3932 (N_3932,N_3362,N_3000);
nor U3933 (N_3933,N_3307,N_3320);
and U3934 (N_3934,N_3268,N_3274);
nand U3935 (N_3935,N_3370,N_3351);
and U3936 (N_3936,N_3027,N_3462);
or U3937 (N_3937,N_3493,N_3385);
nand U3938 (N_3938,N_3051,N_3404);
and U3939 (N_3939,N_3368,N_3411);
nand U3940 (N_3940,N_3095,N_3357);
or U3941 (N_3941,N_3313,N_3320);
nor U3942 (N_3942,N_3179,N_3454);
nor U3943 (N_3943,N_3132,N_3195);
nor U3944 (N_3944,N_3400,N_3214);
nand U3945 (N_3945,N_3044,N_3293);
nand U3946 (N_3946,N_3313,N_3018);
or U3947 (N_3947,N_3281,N_3462);
and U3948 (N_3948,N_3121,N_3476);
and U3949 (N_3949,N_3452,N_3464);
or U3950 (N_3950,N_3203,N_3391);
or U3951 (N_3951,N_3214,N_3186);
and U3952 (N_3952,N_3471,N_3018);
nand U3953 (N_3953,N_3323,N_3011);
nor U3954 (N_3954,N_3119,N_3212);
and U3955 (N_3955,N_3180,N_3205);
nor U3956 (N_3956,N_3298,N_3378);
and U3957 (N_3957,N_3344,N_3141);
nor U3958 (N_3958,N_3434,N_3203);
or U3959 (N_3959,N_3174,N_3262);
xnor U3960 (N_3960,N_3232,N_3474);
nor U3961 (N_3961,N_3029,N_3328);
and U3962 (N_3962,N_3353,N_3129);
or U3963 (N_3963,N_3041,N_3405);
nor U3964 (N_3964,N_3053,N_3118);
and U3965 (N_3965,N_3292,N_3158);
nor U3966 (N_3966,N_3224,N_3179);
or U3967 (N_3967,N_3407,N_3222);
nand U3968 (N_3968,N_3446,N_3480);
nand U3969 (N_3969,N_3329,N_3082);
or U3970 (N_3970,N_3004,N_3207);
and U3971 (N_3971,N_3035,N_3247);
or U3972 (N_3972,N_3474,N_3119);
or U3973 (N_3973,N_3302,N_3434);
nor U3974 (N_3974,N_3302,N_3305);
and U3975 (N_3975,N_3309,N_3420);
or U3976 (N_3976,N_3099,N_3081);
or U3977 (N_3977,N_3007,N_3219);
or U3978 (N_3978,N_3183,N_3187);
nor U3979 (N_3979,N_3223,N_3176);
xor U3980 (N_3980,N_3475,N_3360);
and U3981 (N_3981,N_3098,N_3259);
nand U3982 (N_3982,N_3117,N_3326);
nor U3983 (N_3983,N_3038,N_3151);
nor U3984 (N_3984,N_3390,N_3486);
nand U3985 (N_3985,N_3242,N_3366);
nand U3986 (N_3986,N_3222,N_3390);
or U3987 (N_3987,N_3446,N_3193);
nand U3988 (N_3988,N_3251,N_3394);
nor U3989 (N_3989,N_3465,N_3351);
and U3990 (N_3990,N_3269,N_3111);
and U3991 (N_3991,N_3255,N_3355);
nand U3992 (N_3992,N_3352,N_3260);
nand U3993 (N_3993,N_3195,N_3433);
nor U3994 (N_3994,N_3129,N_3322);
or U3995 (N_3995,N_3296,N_3174);
or U3996 (N_3996,N_3220,N_3080);
xnor U3997 (N_3997,N_3191,N_3023);
nor U3998 (N_3998,N_3371,N_3297);
xnor U3999 (N_3999,N_3462,N_3069);
or U4000 (N_4000,N_3558,N_3811);
xor U4001 (N_4001,N_3716,N_3629);
nand U4002 (N_4002,N_3881,N_3595);
and U4003 (N_4003,N_3824,N_3803);
and U4004 (N_4004,N_3760,N_3704);
nand U4005 (N_4005,N_3796,N_3575);
nand U4006 (N_4006,N_3671,N_3653);
nor U4007 (N_4007,N_3984,N_3788);
or U4008 (N_4008,N_3790,N_3622);
and U4009 (N_4009,N_3988,N_3786);
nor U4010 (N_4010,N_3820,N_3714);
or U4011 (N_4011,N_3917,N_3604);
or U4012 (N_4012,N_3530,N_3841);
or U4013 (N_4013,N_3915,N_3855);
or U4014 (N_4014,N_3623,N_3779);
xor U4015 (N_4015,N_3863,N_3983);
nand U4016 (N_4016,N_3734,N_3837);
or U4017 (N_4017,N_3506,N_3905);
and U4018 (N_4018,N_3891,N_3674);
nand U4019 (N_4019,N_3929,N_3541);
and U4020 (N_4020,N_3962,N_3749);
xor U4021 (N_4021,N_3757,N_3675);
or U4022 (N_4022,N_3933,N_3596);
and U4023 (N_4023,N_3975,N_3518);
nand U4024 (N_4024,N_3708,N_3997);
nand U4025 (N_4025,N_3513,N_3569);
or U4026 (N_4026,N_3774,N_3850);
xor U4027 (N_4027,N_3524,N_3885);
and U4028 (N_4028,N_3924,N_3740);
or U4029 (N_4029,N_3587,N_3783);
nor U4030 (N_4030,N_3620,N_3873);
xor U4031 (N_4031,N_3612,N_3735);
nor U4032 (N_4032,N_3738,N_3882);
xnor U4033 (N_4033,N_3900,N_3746);
and U4034 (N_4034,N_3871,N_3744);
nand U4035 (N_4035,N_3679,N_3553);
and U4036 (N_4036,N_3874,N_3998);
and U4037 (N_4037,N_3586,N_3979);
nand U4038 (N_4038,N_3823,N_3694);
nor U4039 (N_4039,N_3659,N_3794);
or U4040 (N_4040,N_3897,N_3951);
nand U4041 (N_4041,N_3764,N_3529);
or U4042 (N_4042,N_3712,N_3732);
nor U4043 (N_4043,N_3718,N_3835);
nand U4044 (N_4044,N_3603,N_3978);
and U4045 (N_4045,N_3948,N_3695);
and U4046 (N_4046,N_3572,N_3822);
or U4047 (N_4047,N_3958,N_3635);
nor U4048 (N_4048,N_3755,N_3789);
nor U4049 (N_4049,N_3836,N_3970);
nor U4050 (N_4050,N_3935,N_3834);
or U4051 (N_4051,N_3560,N_3827);
or U4052 (N_4052,N_3588,N_3793);
and U4053 (N_4053,N_3724,N_3670);
xnor U4054 (N_4054,N_3512,N_3611);
xor U4055 (N_4055,N_3644,N_3767);
or U4056 (N_4056,N_3548,N_3972);
and U4057 (N_4057,N_3550,N_3934);
nand U4058 (N_4058,N_3840,N_3898);
nor U4059 (N_4059,N_3770,N_3643);
and U4060 (N_4060,N_3906,N_3662);
xnor U4061 (N_4061,N_3528,N_3816);
or U4062 (N_4062,N_3943,N_3949);
nand U4063 (N_4063,N_3614,N_3890);
and U4064 (N_4064,N_3814,N_3974);
nor U4065 (N_4065,N_3883,N_3543);
or U4066 (N_4066,N_3856,N_3846);
or U4067 (N_4067,N_3583,N_3886);
or U4068 (N_4068,N_3689,N_3847);
and U4069 (N_4069,N_3830,N_3936);
and U4070 (N_4070,N_3821,N_3812);
and U4071 (N_4071,N_3869,N_3565);
and U4072 (N_4072,N_3778,N_3868);
nand U4073 (N_4073,N_3758,N_3862);
nand U4074 (N_4074,N_3892,N_3564);
and U4075 (N_4075,N_3768,N_3928);
nor U4076 (N_4076,N_3591,N_3792);
and U4077 (N_4077,N_3665,N_3684);
or U4078 (N_4078,N_3660,N_3651);
nand U4079 (N_4079,N_3809,N_3556);
and U4080 (N_4080,N_3706,N_3872);
nand U4081 (N_4081,N_3804,N_3741);
nor U4082 (N_4082,N_3666,N_3580);
nand U4083 (N_4083,N_3516,N_3961);
and U4084 (N_4084,N_3921,N_3508);
or U4085 (N_4085,N_3593,N_3656);
nor U4086 (N_4086,N_3589,N_3826);
xor U4087 (N_4087,N_3567,N_3568);
or U4088 (N_4088,N_3726,N_3960);
xor U4089 (N_4089,N_3663,N_3613);
xor U4090 (N_4090,N_3707,N_3624);
or U4091 (N_4091,N_3813,N_3888);
or U4092 (N_4092,N_3832,N_3545);
or U4093 (N_4093,N_3923,N_3615);
or U4094 (N_4094,N_3537,N_3552);
or U4095 (N_4095,N_3991,N_3599);
or U4096 (N_4096,N_3807,N_3904);
or U4097 (N_4097,N_3861,N_3681);
nor U4098 (N_4098,N_3699,N_3875);
nor U4099 (N_4099,N_3691,N_3715);
nand U4100 (N_4100,N_3838,N_3655);
or U4101 (N_4101,N_3752,N_3722);
xnor U4102 (N_4102,N_3761,N_3747);
or U4103 (N_4103,N_3525,N_3791);
or U4104 (N_4104,N_3954,N_3627);
nor U4105 (N_4105,N_3678,N_3673);
nor U4106 (N_4106,N_3728,N_3831);
nor U4107 (N_4107,N_3621,N_3992);
nor U4108 (N_4108,N_3851,N_3505);
nor U4109 (N_4109,N_3927,N_3668);
nor U4110 (N_4110,N_3787,N_3600);
and U4111 (N_4111,N_3762,N_3798);
nor U4112 (N_4112,N_3579,N_3766);
or U4113 (N_4113,N_3976,N_3852);
xor U4114 (N_4114,N_3562,N_3946);
and U4115 (N_4115,N_3995,N_3605);
and U4116 (N_4116,N_3769,N_3857);
and U4117 (N_4117,N_3980,N_3971);
nor U4118 (N_4118,N_3781,N_3776);
nor U4119 (N_4119,N_3640,N_3842);
and U4120 (N_4120,N_3990,N_3817);
nand U4121 (N_4121,N_3853,N_3602);
or U4122 (N_4122,N_3889,N_3947);
nand U4123 (N_4123,N_3737,N_3815);
and U4124 (N_4124,N_3739,N_3743);
nand U4125 (N_4125,N_3631,N_3843);
or U4126 (N_4126,N_3730,N_3502);
nor U4127 (N_4127,N_3880,N_3711);
and U4128 (N_4128,N_3986,N_3650);
xnor U4129 (N_4129,N_3563,N_3964);
and U4130 (N_4130,N_3866,N_3557);
and U4131 (N_4131,N_3515,N_3633);
nand U4132 (N_4132,N_3982,N_3994);
or U4133 (N_4133,N_3534,N_3683);
nor U4134 (N_4134,N_3672,N_3780);
nand U4135 (N_4135,N_3941,N_3693);
or U4136 (N_4136,N_3899,N_3517);
nor U4137 (N_4137,N_3657,N_3784);
and U4138 (N_4138,N_3953,N_3782);
nor U4139 (N_4139,N_3955,N_3877);
xor U4140 (N_4140,N_3969,N_3700);
or U4141 (N_4141,N_3864,N_3638);
and U4142 (N_4142,N_3725,N_3685);
and U4143 (N_4143,N_3619,N_3802);
and U4144 (N_4144,N_3985,N_3944);
or U4145 (N_4145,N_3561,N_3876);
xnor U4146 (N_4146,N_3532,N_3977);
nand U4147 (N_4147,N_3625,N_3566);
xnor U4148 (N_4148,N_3639,N_3667);
nor U4149 (N_4149,N_3697,N_3542);
nor U4150 (N_4150,N_3647,N_3753);
or U4151 (N_4151,N_3692,N_3884);
nand U4152 (N_4152,N_3521,N_3652);
or U4153 (N_4153,N_3878,N_3894);
or U4154 (N_4154,N_3705,N_3551);
or U4155 (N_4155,N_3800,N_3909);
nand U4156 (N_4156,N_3617,N_3608);
nand U4157 (N_4157,N_3511,N_3854);
nand U4158 (N_4158,N_3993,N_3931);
and U4159 (N_4159,N_3514,N_3733);
and U4160 (N_4160,N_3637,N_3540);
nor U4161 (N_4161,N_3677,N_3696);
and U4162 (N_4162,N_3698,N_3585);
nand U4163 (N_4163,N_3554,N_3573);
nand U4164 (N_4164,N_3938,N_3531);
or U4165 (N_4165,N_3641,N_3680);
or U4166 (N_4166,N_3773,N_3839);
or U4167 (N_4167,N_3818,N_3661);
or U4168 (N_4168,N_3765,N_3559);
nor U4169 (N_4169,N_3544,N_3945);
nand U4170 (N_4170,N_3597,N_3504);
nor U4171 (N_4171,N_3895,N_3632);
nand U4172 (N_4172,N_3916,N_3642);
nand U4173 (N_4173,N_3932,N_3507);
nand U4174 (N_4174,N_3893,N_3785);
nor U4175 (N_4175,N_3669,N_3922);
nor U4176 (N_4176,N_3865,N_3688);
or U4177 (N_4177,N_3717,N_3844);
nand U4178 (N_4178,N_3582,N_3763);
or U4179 (N_4179,N_3501,N_3584);
nor U4180 (N_4180,N_3819,N_3797);
and U4181 (N_4181,N_3859,N_3523);
nor U4182 (N_4182,N_3825,N_3920);
and U4183 (N_4183,N_3759,N_3887);
and U4184 (N_4184,N_3720,N_3925);
or U4185 (N_4185,N_3918,N_3939);
nor U4186 (N_4186,N_3756,N_3845);
or U4187 (N_4187,N_3658,N_3903);
and U4188 (N_4188,N_3594,N_3795);
or U4189 (N_4189,N_3578,N_3701);
and U4190 (N_4190,N_3555,N_3577);
or U4191 (N_4191,N_3729,N_3713);
nand U4192 (N_4192,N_3709,N_3775);
and U4193 (N_4193,N_3930,N_3526);
nand U4194 (N_4194,N_3676,N_3963);
nand U4195 (N_4195,N_3957,N_3828);
and U4196 (N_4196,N_3772,N_3539);
or U4197 (N_4197,N_3648,N_3618);
nor U4198 (N_4198,N_3967,N_3907);
and U4199 (N_4199,N_3912,N_3649);
nor U4200 (N_4200,N_3867,N_3607);
and U4201 (N_4201,N_3959,N_3754);
nand U4202 (N_4202,N_3896,N_3601);
and U4203 (N_4203,N_3500,N_3702);
and U4204 (N_4204,N_3771,N_3549);
and U4205 (N_4205,N_3522,N_3723);
nand U4206 (N_4206,N_3630,N_3808);
nor U4207 (N_4207,N_3833,N_3727);
or U4208 (N_4208,N_3636,N_3721);
and U4209 (N_4209,N_3520,N_3748);
nor U4210 (N_4210,N_3973,N_3799);
or U4211 (N_4211,N_3628,N_3510);
nor U4212 (N_4212,N_3829,N_3879);
nand U4213 (N_4213,N_3731,N_3503);
and U4214 (N_4214,N_3860,N_3848);
nand U4215 (N_4215,N_3519,N_3968);
or U4216 (N_4216,N_3598,N_3858);
xor U4217 (N_4217,N_3509,N_3626);
xor U4218 (N_4218,N_3745,N_3645);
nand U4219 (N_4219,N_3942,N_3940);
or U4220 (N_4220,N_3581,N_3590);
nand U4221 (N_4221,N_3751,N_3571);
and U4222 (N_4222,N_3996,N_3901);
nand U4223 (N_4223,N_3682,N_3914);
nand U4224 (N_4224,N_3736,N_3999);
nor U4225 (N_4225,N_3606,N_3538);
and U4226 (N_4226,N_3646,N_3664);
and U4227 (N_4227,N_3801,N_3849);
or U4228 (N_4228,N_3989,N_3616);
nor U4229 (N_4229,N_3966,N_3806);
nor U4230 (N_4230,N_3952,N_3570);
and U4231 (N_4231,N_3805,N_3913);
nand U4232 (N_4232,N_3911,N_3687);
or U4233 (N_4233,N_3576,N_3908);
nor U4234 (N_4234,N_3634,N_3777);
nand U4235 (N_4235,N_3654,N_3870);
nand U4236 (N_4236,N_3574,N_3810);
or U4237 (N_4237,N_3742,N_3609);
xnor U4238 (N_4238,N_3610,N_3527);
nor U4239 (N_4239,N_3533,N_3546);
nor U4240 (N_4240,N_3686,N_3950);
nor U4241 (N_4241,N_3926,N_3719);
or U4242 (N_4242,N_3987,N_3910);
nand U4243 (N_4243,N_3710,N_3690);
and U4244 (N_4244,N_3547,N_3919);
nor U4245 (N_4245,N_3592,N_3965);
nor U4246 (N_4246,N_3536,N_3750);
nor U4247 (N_4247,N_3535,N_3956);
or U4248 (N_4248,N_3902,N_3937);
xnor U4249 (N_4249,N_3703,N_3981);
nand U4250 (N_4250,N_3847,N_3684);
nand U4251 (N_4251,N_3595,N_3597);
or U4252 (N_4252,N_3945,N_3520);
nand U4253 (N_4253,N_3912,N_3877);
nand U4254 (N_4254,N_3595,N_3865);
nor U4255 (N_4255,N_3535,N_3975);
nand U4256 (N_4256,N_3526,N_3746);
nor U4257 (N_4257,N_3925,N_3787);
xor U4258 (N_4258,N_3501,N_3721);
and U4259 (N_4259,N_3612,N_3639);
or U4260 (N_4260,N_3684,N_3878);
or U4261 (N_4261,N_3836,N_3813);
nand U4262 (N_4262,N_3922,N_3898);
or U4263 (N_4263,N_3831,N_3538);
nor U4264 (N_4264,N_3500,N_3937);
nor U4265 (N_4265,N_3577,N_3613);
nor U4266 (N_4266,N_3910,N_3611);
or U4267 (N_4267,N_3964,N_3531);
nand U4268 (N_4268,N_3887,N_3662);
or U4269 (N_4269,N_3801,N_3807);
or U4270 (N_4270,N_3885,N_3560);
nor U4271 (N_4271,N_3579,N_3577);
or U4272 (N_4272,N_3900,N_3716);
nor U4273 (N_4273,N_3703,N_3670);
and U4274 (N_4274,N_3746,N_3722);
nand U4275 (N_4275,N_3883,N_3800);
or U4276 (N_4276,N_3863,N_3874);
and U4277 (N_4277,N_3614,N_3683);
nand U4278 (N_4278,N_3632,N_3896);
and U4279 (N_4279,N_3873,N_3938);
nor U4280 (N_4280,N_3836,N_3623);
and U4281 (N_4281,N_3609,N_3791);
nor U4282 (N_4282,N_3942,N_3778);
or U4283 (N_4283,N_3822,N_3602);
nand U4284 (N_4284,N_3835,N_3753);
nand U4285 (N_4285,N_3678,N_3548);
nor U4286 (N_4286,N_3603,N_3810);
nor U4287 (N_4287,N_3790,N_3679);
nor U4288 (N_4288,N_3561,N_3570);
and U4289 (N_4289,N_3861,N_3796);
nor U4290 (N_4290,N_3794,N_3776);
and U4291 (N_4291,N_3528,N_3905);
and U4292 (N_4292,N_3766,N_3757);
nor U4293 (N_4293,N_3739,N_3669);
nand U4294 (N_4294,N_3575,N_3812);
nor U4295 (N_4295,N_3804,N_3653);
nor U4296 (N_4296,N_3831,N_3987);
or U4297 (N_4297,N_3536,N_3579);
xor U4298 (N_4298,N_3685,N_3732);
nand U4299 (N_4299,N_3754,N_3970);
or U4300 (N_4300,N_3656,N_3782);
xnor U4301 (N_4301,N_3659,N_3990);
nor U4302 (N_4302,N_3571,N_3734);
or U4303 (N_4303,N_3525,N_3678);
nor U4304 (N_4304,N_3874,N_3942);
and U4305 (N_4305,N_3540,N_3527);
or U4306 (N_4306,N_3758,N_3586);
nor U4307 (N_4307,N_3831,N_3688);
and U4308 (N_4308,N_3975,N_3597);
or U4309 (N_4309,N_3758,N_3844);
xnor U4310 (N_4310,N_3950,N_3507);
xnor U4311 (N_4311,N_3873,N_3755);
or U4312 (N_4312,N_3957,N_3919);
or U4313 (N_4313,N_3992,N_3677);
and U4314 (N_4314,N_3783,N_3901);
and U4315 (N_4315,N_3701,N_3979);
or U4316 (N_4316,N_3820,N_3826);
and U4317 (N_4317,N_3770,N_3980);
or U4318 (N_4318,N_3579,N_3811);
or U4319 (N_4319,N_3944,N_3529);
nand U4320 (N_4320,N_3584,N_3909);
or U4321 (N_4321,N_3567,N_3678);
or U4322 (N_4322,N_3824,N_3740);
nor U4323 (N_4323,N_3934,N_3601);
or U4324 (N_4324,N_3757,N_3798);
nand U4325 (N_4325,N_3636,N_3916);
or U4326 (N_4326,N_3844,N_3847);
nand U4327 (N_4327,N_3922,N_3980);
xor U4328 (N_4328,N_3501,N_3871);
and U4329 (N_4329,N_3567,N_3921);
nand U4330 (N_4330,N_3693,N_3819);
and U4331 (N_4331,N_3622,N_3509);
or U4332 (N_4332,N_3535,N_3997);
nor U4333 (N_4333,N_3749,N_3651);
and U4334 (N_4334,N_3853,N_3574);
and U4335 (N_4335,N_3735,N_3852);
nand U4336 (N_4336,N_3600,N_3676);
and U4337 (N_4337,N_3903,N_3879);
and U4338 (N_4338,N_3523,N_3803);
and U4339 (N_4339,N_3518,N_3968);
and U4340 (N_4340,N_3635,N_3679);
nor U4341 (N_4341,N_3576,N_3672);
or U4342 (N_4342,N_3803,N_3909);
and U4343 (N_4343,N_3915,N_3615);
nor U4344 (N_4344,N_3724,N_3806);
nor U4345 (N_4345,N_3816,N_3956);
nor U4346 (N_4346,N_3715,N_3828);
nand U4347 (N_4347,N_3891,N_3754);
nor U4348 (N_4348,N_3917,N_3829);
or U4349 (N_4349,N_3624,N_3901);
or U4350 (N_4350,N_3758,N_3793);
and U4351 (N_4351,N_3950,N_3723);
nand U4352 (N_4352,N_3695,N_3799);
nor U4353 (N_4353,N_3645,N_3689);
nand U4354 (N_4354,N_3777,N_3705);
nand U4355 (N_4355,N_3832,N_3603);
and U4356 (N_4356,N_3809,N_3884);
and U4357 (N_4357,N_3914,N_3797);
and U4358 (N_4358,N_3508,N_3857);
nand U4359 (N_4359,N_3500,N_3893);
or U4360 (N_4360,N_3886,N_3544);
nor U4361 (N_4361,N_3885,N_3993);
or U4362 (N_4362,N_3543,N_3500);
or U4363 (N_4363,N_3585,N_3940);
nor U4364 (N_4364,N_3875,N_3634);
and U4365 (N_4365,N_3511,N_3729);
or U4366 (N_4366,N_3639,N_3560);
nor U4367 (N_4367,N_3722,N_3723);
and U4368 (N_4368,N_3756,N_3769);
and U4369 (N_4369,N_3509,N_3933);
nor U4370 (N_4370,N_3942,N_3695);
xnor U4371 (N_4371,N_3888,N_3640);
nor U4372 (N_4372,N_3704,N_3778);
or U4373 (N_4373,N_3646,N_3791);
nand U4374 (N_4374,N_3544,N_3546);
and U4375 (N_4375,N_3984,N_3550);
nor U4376 (N_4376,N_3982,N_3592);
nor U4377 (N_4377,N_3513,N_3886);
and U4378 (N_4378,N_3741,N_3582);
nor U4379 (N_4379,N_3792,N_3976);
and U4380 (N_4380,N_3648,N_3833);
nor U4381 (N_4381,N_3663,N_3745);
nor U4382 (N_4382,N_3992,N_3771);
xnor U4383 (N_4383,N_3568,N_3555);
nor U4384 (N_4384,N_3855,N_3816);
nor U4385 (N_4385,N_3788,N_3576);
or U4386 (N_4386,N_3525,N_3875);
nor U4387 (N_4387,N_3910,N_3735);
nor U4388 (N_4388,N_3726,N_3623);
nand U4389 (N_4389,N_3963,N_3688);
or U4390 (N_4390,N_3805,N_3699);
or U4391 (N_4391,N_3806,N_3803);
or U4392 (N_4392,N_3756,N_3714);
or U4393 (N_4393,N_3824,N_3617);
or U4394 (N_4394,N_3979,N_3755);
or U4395 (N_4395,N_3512,N_3722);
or U4396 (N_4396,N_3843,N_3636);
xor U4397 (N_4397,N_3840,N_3800);
nand U4398 (N_4398,N_3704,N_3640);
nand U4399 (N_4399,N_3915,N_3758);
nor U4400 (N_4400,N_3512,N_3651);
or U4401 (N_4401,N_3572,N_3941);
or U4402 (N_4402,N_3833,N_3730);
nor U4403 (N_4403,N_3816,N_3797);
nand U4404 (N_4404,N_3555,N_3710);
nand U4405 (N_4405,N_3967,N_3846);
nor U4406 (N_4406,N_3899,N_3846);
nand U4407 (N_4407,N_3861,N_3868);
or U4408 (N_4408,N_3808,N_3748);
and U4409 (N_4409,N_3576,N_3929);
xnor U4410 (N_4410,N_3706,N_3993);
and U4411 (N_4411,N_3932,N_3906);
nor U4412 (N_4412,N_3675,N_3992);
xnor U4413 (N_4413,N_3921,N_3886);
nand U4414 (N_4414,N_3633,N_3529);
nor U4415 (N_4415,N_3850,N_3621);
nand U4416 (N_4416,N_3978,N_3836);
or U4417 (N_4417,N_3809,N_3673);
and U4418 (N_4418,N_3974,N_3529);
nand U4419 (N_4419,N_3519,N_3589);
nor U4420 (N_4420,N_3790,N_3649);
nand U4421 (N_4421,N_3517,N_3877);
and U4422 (N_4422,N_3695,N_3520);
nand U4423 (N_4423,N_3556,N_3877);
or U4424 (N_4424,N_3826,N_3825);
or U4425 (N_4425,N_3796,N_3747);
nand U4426 (N_4426,N_3988,N_3921);
xnor U4427 (N_4427,N_3714,N_3884);
or U4428 (N_4428,N_3538,N_3852);
xnor U4429 (N_4429,N_3730,N_3644);
nor U4430 (N_4430,N_3734,N_3578);
and U4431 (N_4431,N_3732,N_3744);
or U4432 (N_4432,N_3885,N_3721);
or U4433 (N_4433,N_3858,N_3619);
and U4434 (N_4434,N_3752,N_3931);
and U4435 (N_4435,N_3923,N_3765);
or U4436 (N_4436,N_3760,N_3802);
or U4437 (N_4437,N_3997,N_3828);
xor U4438 (N_4438,N_3559,N_3741);
nand U4439 (N_4439,N_3817,N_3769);
and U4440 (N_4440,N_3955,N_3796);
and U4441 (N_4441,N_3512,N_3917);
nand U4442 (N_4442,N_3739,N_3927);
nor U4443 (N_4443,N_3967,N_3652);
nor U4444 (N_4444,N_3527,N_3546);
nand U4445 (N_4445,N_3920,N_3803);
nand U4446 (N_4446,N_3541,N_3689);
nand U4447 (N_4447,N_3645,N_3632);
nand U4448 (N_4448,N_3995,N_3840);
and U4449 (N_4449,N_3829,N_3726);
xnor U4450 (N_4450,N_3713,N_3920);
xnor U4451 (N_4451,N_3533,N_3569);
or U4452 (N_4452,N_3744,N_3931);
xnor U4453 (N_4453,N_3962,N_3928);
or U4454 (N_4454,N_3670,N_3905);
and U4455 (N_4455,N_3552,N_3705);
nand U4456 (N_4456,N_3780,N_3921);
or U4457 (N_4457,N_3619,N_3825);
and U4458 (N_4458,N_3537,N_3539);
xnor U4459 (N_4459,N_3780,N_3851);
or U4460 (N_4460,N_3959,N_3869);
nor U4461 (N_4461,N_3874,N_3558);
and U4462 (N_4462,N_3562,N_3805);
xnor U4463 (N_4463,N_3529,N_3787);
nand U4464 (N_4464,N_3830,N_3774);
nor U4465 (N_4465,N_3745,N_3573);
xor U4466 (N_4466,N_3760,N_3873);
xnor U4467 (N_4467,N_3503,N_3641);
nor U4468 (N_4468,N_3926,N_3949);
and U4469 (N_4469,N_3756,N_3720);
nor U4470 (N_4470,N_3805,N_3557);
and U4471 (N_4471,N_3936,N_3945);
and U4472 (N_4472,N_3544,N_3731);
and U4473 (N_4473,N_3815,N_3653);
xnor U4474 (N_4474,N_3574,N_3880);
nand U4475 (N_4475,N_3785,N_3570);
xnor U4476 (N_4476,N_3505,N_3519);
and U4477 (N_4477,N_3690,N_3754);
or U4478 (N_4478,N_3551,N_3516);
or U4479 (N_4479,N_3900,N_3526);
nand U4480 (N_4480,N_3676,N_3507);
or U4481 (N_4481,N_3998,N_3773);
and U4482 (N_4482,N_3710,N_3850);
xor U4483 (N_4483,N_3896,N_3666);
or U4484 (N_4484,N_3930,N_3771);
and U4485 (N_4485,N_3590,N_3981);
or U4486 (N_4486,N_3508,N_3716);
nand U4487 (N_4487,N_3612,N_3743);
and U4488 (N_4488,N_3740,N_3611);
or U4489 (N_4489,N_3941,N_3604);
or U4490 (N_4490,N_3969,N_3767);
or U4491 (N_4491,N_3772,N_3824);
nand U4492 (N_4492,N_3753,N_3943);
xor U4493 (N_4493,N_3663,N_3537);
nor U4494 (N_4494,N_3680,N_3779);
or U4495 (N_4495,N_3766,N_3887);
xnor U4496 (N_4496,N_3926,N_3852);
nor U4497 (N_4497,N_3763,N_3738);
xor U4498 (N_4498,N_3599,N_3856);
nand U4499 (N_4499,N_3647,N_3655);
nand U4500 (N_4500,N_4380,N_4228);
nand U4501 (N_4501,N_4344,N_4077);
nor U4502 (N_4502,N_4140,N_4249);
nand U4503 (N_4503,N_4285,N_4186);
xnor U4504 (N_4504,N_4447,N_4289);
or U4505 (N_4505,N_4423,N_4343);
nand U4506 (N_4506,N_4340,N_4378);
or U4507 (N_4507,N_4113,N_4133);
or U4508 (N_4508,N_4466,N_4135);
nand U4509 (N_4509,N_4170,N_4111);
and U4510 (N_4510,N_4411,N_4109);
or U4511 (N_4511,N_4098,N_4345);
or U4512 (N_4512,N_4335,N_4421);
xnor U4513 (N_4513,N_4040,N_4292);
or U4514 (N_4514,N_4000,N_4174);
and U4515 (N_4515,N_4473,N_4153);
xnor U4516 (N_4516,N_4264,N_4161);
and U4517 (N_4517,N_4189,N_4350);
xnor U4518 (N_4518,N_4367,N_4014);
nor U4519 (N_4519,N_4015,N_4461);
or U4520 (N_4520,N_4169,N_4194);
or U4521 (N_4521,N_4406,N_4073);
or U4522 (N_4522,N_4079,N_4360);
nor U4523 (N_4523,N_4104,N_4469);
nor U4524 (N_4524,N_4474,N_4400);
and U4525 (N_4525,N_4033,N_4084);
or U4526 (N_4526,N_4148,N_4349);
nand U4527 (N_4527,N_4041,N_4106);
and U4528 (N_4528,N_4201,N_4067);
or U4529 (N_4529,N_4375,N_4499);
or U4530 (N_4530,N_4200,N_4222);
or U4531 (N_4531,N_4008,N_4063);
and U4532 (N_4532,N_4171,N_4483);
or U4533 (N_4533,N_4205,N_4495);
and U4534 (N_4534,N_4308,N_4478);
nor U4535 (N_4535,N_4432,N_4385);
nand U4536 (N_4536,N_4456,N_4341);
or U4537 (N_4537,N_4134,N_4187);
and U4538 (N_4538,N_4061,N_4017);
nor U4539 (N_4539,N_4379,N_4229);
xnor U4540 (N_4540,N_4177,N_4271);
nand U4541 (N_4541,N_4108,N_4147);
or U4542 (N_4542,N_4458,N_4368);
xnor U4543 (N_4543,N_4465,N_4353);
and U4544 (N_4544,N_4481,N_4317);
nand U4545 (N_4545,N_4139,N_4355);
or U4546 (N_4546,N_4386,N_4418);
nor U4547 (N_4547,N_4371,N_4300);
nand U4548 (N_4548,N_4298,N_4036);
nor U4549 (N_4549,N_4444,N_4382);
nor U4550 (N_4550,N_4373,N_4198);
or U4551 (N_4551,N_4269,N_4088);
nand U4552 (N_4552,N_4207,N_4052);
and U4553 (N_4553,N_4286,N_4120);
and U4554 (N_4554,N_4283,N_4241);
nand U4555 (N_4555,N_4393,N_4125);
nor U4556 (N_4556,N_4438,N_4116);
and U4557 (N_4557,N_4152,N_4055);
xor U4558 (N_4558,N_4351,N_4107);
nor U4559 (N_4559,N_4457,N_4387);
or U4560 (N_4560,N_4306,N_4346);
nand U4561 (N_4561,N_4434,N_4081);
nand U4562 (N_4562,N_4415,N_4244);
xnor U4563 (N_4563,N_4414,N_4058);
or U4564 (N_4564,N_4488,N_4131);
nor U4565 (N_4565,N_4181,N_4090);
and U4566 (N_4566,N_4020,N_4333);
nand U4567 (N_4567,N_4272,N_4007);
and U4568 (N_4568,N_4004,N_4236);
nor U4569 (N_4569,N_4195,N_4326);
xor U4570 (N_4570,N_4093,N_4383);
and U4571 (N_4571,N_4476,N_4211);
and U4572 (N_4572,N_4295,N_4384);
xnor U4573 (N_4573,N_4451,N_4489);
and U4574 (N_4574,N_4167,N_4149);
or U4575 (N_4575,N_4193,N_4394);
nand U4576 (N_4576,N_4275,N_4239);
and U4577 (N_4577,N_4471,N_4254);
xor U4578 (N_4578,N_4137,N_4316);
nand U4579 (N_4579,N_4190,N_4182);
nor U4580 (N_4580,N_4376,N_4206);
or U4581 (N_4581,N_4409,N_4462);
nand U4582 (N_4582,N_4163,N_4321);
xnor U4583 (N_4583,N_4362,N_4218);
or U4584 (N_4584,N_4401,N_4331);
xor U4585 (N_4585,N_4196,N_4112);
xor U4586 (N_4586,N_4043,N_4310);
and U4587 (N_4587,N_4035,N_4010);
nand U4588 (N_4588,N_4332,N_4048);
and U4589 (N_4589,N_4012,N_4099);
xor U4590 (N_4590,N_4365,N_4301);
nor U4591 (N_4591,N_4407,N_4215);
nand U4592 (N_4592,N_4482,N_4097);
nor U4593 (N_4593,N_4044,N_4138);
nand U4594 (N_4594,N_4188,N_4083);
or U4595 (N_4595,N_4220,N_4213);
and U4596 (N_4596,N_4297,N_4042);
xnor U4597 (N_4597,N_4389,N_4231);
or U4598 (N_4598,N_4202,N_4026);
or U4599 (N_4599,N_4240,N_4075);
and U4600 (N_4600,N_4381,N_4025);
or U4601 (N_4601,N_4277,N_4255);
xor U4602 (N_4602,N_4160,N_4024);
or U4603 (N_4603,N_4094,N_4175);
and U4604 (N_4604,N_4404,N_4433);
and U4605 (N_4605,N_4288,N_4467);
nand U4606 (N_4606,N_4027,N_4136);
and U4607 (N_4607,N_4183,N_4173);
nor U4608 (N_4608,N_4494,N_4266);
nand U4609 (N_4609,N_4251,N_4060);
or U4610 (N_4610,N_4477,N_4492);
or U4611 (N_4611,N_4057,N_4263);
or U4612 (N_4612,N_4029,N_4059);
or U4613 (N_4613,N_4180,N_4356);
xnor U4614 (N_4614,N_4219,N_4031);
or U4615 (N_4615,N_4006,N_4037);
or U4616 (N_4616,N_4118,N_4459);
nor U4617 (N_4617,N_4224,N_4009);
and U4618 (N_4618,N_4399,N_4439);
nand U4619 (N_4619,N_4357,N_4290);
and U4620 (N_4620,N_4150,N_4078);
nor U4621 (N_4621,N_4080,N_4179);
nor U4622 (N_4622,N_4309,N_4337);
nor U4623 (N_4623,N_4436,N_4199);
nand U4624 (N_4624,N_4440,N_4420);
or U4625 (N_4625,N_4330,N_4273);
nor U4626 (N_4626,N_4416,N_4145);
xnor U4627 (N_4627,N_4156,N_4247);
nand U4628 (N_4628,N_4463,N_4311);
and U4629 (N_4629,N_4287,N_4279);
or U4630 (N_4630,N_4486,N_4305);
and U4631 (N_4631,N_4086,N_4257);
or U4632 (N_4632,N_4424,N_4313);
and U4633 (N_4633,N_4450,N_4100);
and U4634 (N_4634,N_4221,N_4270);
nor U4635 (N_4635,N_4066,N_4312);
and U4636 (N_4636,N_4105,N_4338);
or U4637 (N_4637,N_4296,N_4028);
and U4638 (N_4638,N_4324,N_4455);
nor U4639 (N_4639,N_4342,N_4437);
nand U4640 (N_4640,N_4267,N_4413);
nand U4641 (N_4641,N_4051,N_4019);
and U4642 (N_4642,N_4070,N_4121);
or U4643 (N_4643,N_4082,N_4352);
nand U4644 (N_4644,N_4262,N_4216);
and U4645 (N_4645,N_4128,N_4155);
or U4646 (N_4646,N_4119,N_4475);
and U4647 (N_4647,N_4126,N_4226);
and U4648 (N_4648,N_4261,N_4274);
xor U4649 (N_4649,N_4363,N_4322);
nor U4650 (N_4650,N_4197,N_4364);
xor U4651 (N_4651,N_4302,N_4103);
or U4652 (N_4652,N_4192,N_4168);
and U4653 (N_4653,N_4038,N_4178);
xor U4654 (N_4654,N_4238,N_4243);
and U4655 (N_4655,N_4130,N_4165);
or U4656 (N_4656,N_4101,N_4422);
and U4657 (N_4657,N_4203,N_4252);
and U4658 (N_4658,N_4487,N_4282);
nand U4659 (N_4659,N_4072,N_4154);
or U4660 (N_4660,N_4314,N_4242);
nor U4661 (N_4661,N_4230,N_4303);
and U4662 (N_4662,N_4054,N_4110);
nand U4663 (N_4663,N_4122,N_4001);
and U4664 (N_4664,N_4348,N_4491);
nor U4665 (N_4665,N_4425,N_4472);
xor U4666 (N_4666,N_4428,N_4497);
or U4667 (N_4667,N_4347,N_4032);
nor U4668 (N_4668,N_4328,N_4443);
or U4669 (N_4669,N_4291,N_4396);
or U4670 (N_4670,N_4498,N_4064);
or U4671 (N_4671,N_4071,N_4370);
or U4672 (N_4672,N_4184,N_4265);
nand U4673 (N_4673,N_4076,N_4325);
nand U4674 (N_4674,N_4448,N_4430);
nor U4675 (N_4675,N_4039,N_4449);
nand U4676 (N_4676,N_4369,N_4320);
or U4677 (N_4677,N_4127,N_4096);
xor U4678 (N_4678,N_4095,N_4157);
nand U4679 (N_4679,N_4278,N_4315);
or U4680 (N_4680,N_4217,N_4294);
or U4681 (N_4681,N_4208,N_4388);
nor U4682 (N_4682,N_4237,N_4258);
or U4683 (N_4683,N_4452,N_4016);
nor U4684 (N_4684,N_4377,N_4276);
or U4685 (N_4685,N_4429,N_4062);
or U4686 (N_4686,N_4256,N_4018);
or U4687 (N_4687,N_4232,N_4246);
nand U4688 (N_4688,N_4124,N_4453);
and U4689 (N_4689,N_4435,N_4468);
nor U4690 (N_4690,N_4132,N_4210);
or U4691 (N_4691,N_4490,N_4403);
and U4692 (N_4692,N_4299,N_4069);
nor U4693 (N_4693,N_4053,N_4446);
nand U4694 (N_4694,N_4336,N_4454);
nor U4695 (N_4695,N_4390,N_4144);
nor U4696 (N_4696,N_4253,N_4307);
nand U4697 (N_4697,N_4158,N_4259);
nand U4698 (N_4698,N_4002,N_4260);
nor U4699 (N_4699,N_4123,N_4146);
nor U4700 (N_4700,N_4049,N_4493);
and U4701 (N_4701,N_4402,N_4023);
or U4702 (N_4702,N_4003,N_4092);
nor U4703 (N_4703,N_4176,N_4392);
or U4704 (N_4704,N_4479,N_4085);
and U4705 (N_4705,N_4227,N_4426);
xor U4706 (N_4706,N_4047,N_4419);
nand U4707 (N_4707,N_4089,N_4159);
or U4708 (N_4708,N_4225,N_4074);
or U4709 (N_4709,N_4021,N_4166);
nor U4710 (N_4710,N_4114,N_4372);
and U4711 (N_4711,N_4318,N_4204);
and U4712 (N_4712,N_4046,N_4212);
or U4713 (N_4713,N_4485,N_4065);
and U4714 (N_4714,N_4172,N_4366);
and U4715 (N_4715,N_4034,N_4293);
and U4716 (N_4716,N_4143,N_4405);
xor U4717 (N_4717,N_4470,N_4398);
xor U4718 (N_4718,N_4408,N_4091);
nor U4719 (N_4719,N_4395,N_4056);
or U4720 (N_4720,N_4191,N_4087);
nand U4721 (N_4721,N_4068,N_4235);
or U4722 (N_4722,N_4268,N_4011);
or U4723 (N_4723,N_4445,N_4129);
or U4724 (N_4724,N_4248,N_4361);
xnor U4725 (N_4725,N_4359,N_4339);
and U4726 (N_4726,N_4374,N_4329);
and U4727 (N_4727,N_4304,N_4005);
and U4728 (N_4728,N_4045,N_4151);
nor U4729 (N_4729,N_4233,N_4480);
or U4730 (N_4730,N_4464,N_4334);
nor U4731 (N_4731,N_4431,N_4442);
nor U4732 (N_4732,N_4117,N_4484);
nand U4733 (N_4733,N_4164,N_4460);
xor U4734 (N_4734,N_4417,N_4427);
and U4735 (N_4735,N_4115,N_4250);
nand U4736 (N_4736,N_4141,N_4142);
and U4737 (N_4737,N_4354,N_4162);
or U4738 (N_4738,N_4185,N_4013);
and U4739 (N_4739,N_4102,N_4358);
nand U4740 (N_4740,N_4412,N_4280);
and U4741 (N_4741,N_4030,N_4397);
and U4742 (N_4742,N_4323,N_4391);
and U4743 (N_4743,N_4050,N_4245);
nand U4744 (N_4744,N_4281,N_4327);
and U4745 (N_4745,N_4496,N_4022);
and U4746 (N_4746,N_4441,N_4410);
and U4747 (N_4747,N_4284,N_4319);
nand U4748 (N_4748,N_4209,N_4214);
nor U4749 (N_4749,N_4223,N_4234);
nand U4750 (N_4750,N_4037,N_4127);
xnor U4751 (N_4751,N_4339,N_4077);
nor U4752 (N_4752,N_4285,N_4488);
or U4753 (N_4753,N_4029,N_4101);
xnor U4754 (N_4754,N_4002,N_4258);
nand U4755 (N_4755,N_4354,N_4336);
and U4756 (N_4756,N_4276,N_4249);
or U4757 (N_4757,N_4290,N_4005);
nand U4758 (N_4758,N_4310,N_4366);
nor U4759 (N_4759,N_4031,N_4086);
and U4760 (N_4760,N_4422,N_4121);
nor U4761 (N_4761,N_4483,N_4429);
xnor U4762 (N_4762,N_4207,N_4372);
nor U4763 (N_4763,N_4262,N_4100);
nand U4764 (N_4764,N_4357,N_4031);
nand U4765 (N_4765,N_4047,N_4253);
nand U4766 (N_4766,N_4253,N_4163);
and U4767 (N_4767,N_4305,N_4389);
nor U4768 (N_4768,N_4131,N_4307);
and U4769 (N_4769,N_4129,N_4443);
and U4770 (N_4770,N_4166,N_4450);
and U4771 (N_4771,N_4101,N_4332);
nand U4772 (N_4772,N_4049,N_4089);
and U4773 (N_4773,N_4124,N_4423);
xnor U4774 (N_4774,N_4053,N_4137);
and U4775 (N_4775,N_4492,N_4440);
nand U4776 (N_4776,N_4369,N_4127);
nand U4777 (N_4777,N_4460,N_4101);
and U4778 (N_4778,N_4393,N_4442);
nor U4779 (N_4779,N_4260,N_4464);
nand U4780 (N_4780,N_4087,N_4156);
or U4781 (N_4781,N_4150,N_4300);
or U4782 (N_4782,N_4068,N_4315);
nand U4783 (N_4783,N_4199,N_4401);
nand U4784 (N_4784,N_4465,N_4166);
and U4785 (N_4785,N_4434,N_4208);
nor U4786 (N_4786,N_4398,N_4268);
nor U4787 (N_4787,N_4195,N_4029);
xnor U4788 (N_4788,N_4103,N_4049);
or U4789 (N_4789,N_4077,N_4361);
nand U4790 (N_4790,N_4452,N_4342);
and U4791 (N_4791,N_4077,N_4107);
or U4792 (N_4792,N_4401,N_4378);
or U4793 (N_4793,N_4022,N_4155);
nor U4794 (N_4794,N_4015,N_4292);
nand U4795 (N_4795,N_4205,N_4044);
nor U4796 (N_4796,N_4251,N_4247);
and U4797 (N_4797,N_4032,N_4180);
or U4798 (N_4798,N_4130,N_4309);
or U4799 (N_4799,N_4429,N_4393);
nor U4800 (N_4800,N_4167,N_4380);
nor U4801 (N_4801,N_4213,N_4339);
nand U4802 (N_4802,N_4385,N_4152);
nand U4803 (N_4803,N_4314,N_4131);
nand U4804 (N_4804,N_4175,N_4019);
or U4805 (N_4805,N_4113,N_4382);
or U4806 (N_4806,N_4150,N_4183);
nand U4807 (N_4807,N_4358,N_4158);
and U4808 (N_4808,N_4274,N_4368);
or U4809 (N_4809,N_4408,N_4122);
and U4810 (N_4810,N_4096,N_4315);
nand U4811 (N_4811,N_4171,N_4137);
and U4812 (N_4812,N_4327,N_4347);
or U4813 (N_4813,N_4293,N_4462);
and U4814 (N_4814,N_4400,N_4259);
or U4815 (N_4815,N_4031,N_4300);
nor U4816 (N_4816,N_4455,N_4421);
nor U4817 (N_4817,N_4019,N_4179);
and U4818 (N_4818,N_4128,N_4466);
and U4819 (N_4819,N_4165,N_4079);
nand U4820 (N_4820,N_4334,N_4116);
nand U4821 (N_4821,N_4094,N_4152);
nor U4822 (N_4822,N_4225,N_4022);
xor U4823 (N_4823,N_4119,N_4230);
or U4824 (N_4824,N_4191,N_4336);
xor U4825 (N_4825,N_4260,N_4080);
nor U4826 (N_4826,N_4393,N_4499);
and U4827 (N_4827,N_4271,N_4065);
nor U4828 (N_4828,N_4260,N_4219);
and U4829 (N_4829,N_4078,N_4095);
nor U4830 (N_4830,N_4148,N_4229);
nand U4831 (N_4831,N_4340,N_4022);
or U4832 (N_4832,N_4361,N_4317);
nand U4833 (N_4833,N_4129,N_4336);
or U4834 (N_4834,N_4151,N_4492);
nand U4835 (N_4835,N_4450,N_4248);
xnor U4836 (N_4836,N_4333,N_4171);
or U4837 (N_4837,N_4339,N_4033);
or U4838 (N_4838,N_4116,N_4371);
nand U4839 (N_4839,N_4157,N_4477);
nand U4840 (N_4840,N_4117,N_4396);
or U4841 (N_4841,N_4038,N_4324);
nor U4842 (N_4842,N_4155,N_4390);
or U4843 (N_4843,N_4114,N_4455);
nand U4844 (N_4844,N_4138,N_4249);
and U4845 (N_4845,N_4140,N_4320);
and U4846 (N_4846,N_4486,N_4450);
xor U4847 (N_4847,N_4272,N_4237);
nand U4848 (N_4848,N_4434,N_4438);
and U4849 (N_4849,N_4250,N_4292);
or U4850 (N_4850,N_4134,N_4412);
xor U4851 (N_4851,N_4184,N_4178);
nand U4852 (N_4852,N_4037,N_4227);
nand U4853 (N_4853,N_4348,N_4127);
nand U4854 (N_4854,N_4405,N_4149);
nand U4855 (N_4855,N_4088,N_4498);
or U4856 (N_4856,N_4048,N_4146);
or U4857 (N_4857,N_4486,N_4281);
nand U4858 (N_4858,N_4412,N_4052);
or U4859 (N_4859,N_4274,N_4205);
nor U4860 (N_4860,N_4441,N_4390);
or U4861 (N_4861,N_4418,N_4034);
nor U4862 (N_4862,N_4284,N_4377);
nand U4863 (N_4863,N_4060,N_4174);
nor U4864 (N_4864,N_4131,N_4478);
or U4865 (N_4865,N_4037,N_4433);
and U4866 (N_4866,N_4379,N_4331);
and U4867 (N_4867,N_4348,N_4471);
nand U4868 (N_4868,N_4391,N_4189);
or U4869 (N_4869,N_4185,N_4263);
nand U4870 (N_4870,N_4133,N_4365);
xnor U4871 (N_4871,N_4243,N_4140);
and U4872 (N_4872,N_4331,N_4304);
nand U4873 (N_4873,N_4246,N_4432);
nor U4874 (N_4874,N_4451,N_4039);
nand U4875 (N_4875,N_4385,N_4356);
or U4876 (N_4876,N_4049,N_4124);
or U4877 (N_4877,N_4491,N_4415);
and U4878 (N_4878,N_4016,N_4424);
nor U4879 (N_4879,N_4200,N_4003);
or U4880 (N_4880,N_4490,N_4330);
nand U4881 (N_4881,N_4312,N_4212);
or U4882 (N_4882,N_4118,N_4414);
and U4883 (N_4883,N_4017,N_4307);
and U4884 (N_4884,N_4344,N_4454);
or U4885 (N_4885,N_4139,N_4362);
xor U4886 (N_4886,N_4415,N_4199);
or U4887 (N_4887,N_4132,N_4187);
nand U4888 (N_4888,N_4107,N_4159);
and U4889 (N_4889,N_4381,N_4037);
nor U4890 (N_4890,N_4164,N_4186);
xor U4891 (N_4891,N_4208,N_4039);
or U4892 (N_4892,N_4148,N_4266);
and U4893 (N_4893,N_4248,N_4269);
and U4894 (N_4894,N_4352,N_4223);
or U4895 (N_4895,N_4339,N_4036);
and U4896 (N_4896,N_4157,N_4088);
nor U4897 (N_4897,N_4174,N_4493);
nor U4898 (N_4898,N_4391,N_4438);
nand U4899 (N_4899,N_4421,N_4278);
and U4900 (N_4900,N_4473,N_4388);
nor U4901 (N_4901,N_4299,N_4490);
or U4902 (N_4902,N_4096,N_4080);
nor U4903 (N_4903,N_4047,N_4019);
or U4904 (N_4904,N_4219,N_4023);
and U4905 (N_4905,N_4039,N_4431);
nand U4906 (N_4906,N_4496,N_4124);
nor U4907 (N_4907,N_4179,N_4227);
and U4908 (N_4908,N_4150,N_4427);
nand U4909 (N_4909,N_4017,N_4284);
nand U4910 (N_4910,N_4391,N_4345);
nand U4911 (N_4911,N_4070,N_4156);
nand U4912 (N_4912,N_4483,N_4261);
xnor U4913 (N_4913,N_4035,N_4227);
nand U4914 (N_4914,N_4118,N_4471);
and U4915 (N_4915,N_4265,N_4075);
and U4916 (N_4916,N_4467,N_4305);
nor U4917 (N_4917,N_4220,N_4385);
or U4918 (N_4918,N_4307,N_4256);
nand U4919 (N_4919,N_4316,N_4270);
or U4920 (N_4920,N_4004,N_4058);
or U4921 (N_4921,N_4230,N_4080);
nor U4922 (N_4922,N_4355,N_4361);
nand U4923 (N_4923,N_4040,N_4078);
nand U4924 (N_4924,N_4365,N_4315);
or U4925 (N_4925,N_4101,N_4055);
or U4926 (N_4926,N_4217,N_4033);
nor U4927 (N_4927,N_4202,N_4132);
nor U4928 (N_4928,N_4301,N_4040);
and U4929 (N_4929,N_4220,N_4359);
nor U4930 (N_4930,N_4260,N_4436);
and U4931 (N_4931,N_4397,N_4165);
xnor U4932 (N_4932,N_4378,N_4273);
and U4933 (N_4933,N_4215,N_4023);
nor U4934 (N_4934,N_4337,N_4008);
or U4935 (N_4935,N_4054,N_4470);
xor U4936 (N_4936,N_4187,N_4094);
or U4937 (N_4937,N_4146,N_4283);
nor U4938 (N_4938,N_4196,N_4158);
and U4939 (N_4939,N_4298,N_4037);
nor U4940 (N_4940,N_4071,N_4204);
nand U4941 (N_4941,N_4244,N_4133);
xnor U4942 (N_4942,N_4207,N_4399);
and U4943 (N_4943,N_4019,N_4458);
and U4944 (N_4944,N_4466,N_4403);
nor U4945 (N_4945,N_4138,N_4072);
or U4946 (N_4946,N_4047,N_4106);
or U4947 (N_4947,N_4362,N_4456);
nor U4948 (N_4948,N_4131,N_4248);
nand U4949 (N_4949,N_4056,N_4306);
nand U4950 (N_4950,N_4014,N_4352);
or U4951 (N_4951,N_4368,N_4336);
or U4952 (N_4952,N_4193,N_4025);
and U4953 (N_4953,N_4405,N_4319);
nor U4954 (N_4954,N_4028,N_4081);
nor U4955 (N_4955,N_4217,N_4377);
and U4956 (N_4956,N_4272,N_4051);
nor U4957 (N_4957,N_4245,N_4466);
and U4958 (N_4958,N_4238,N_4192);
nor U4959 (N_4959,N_4030,N_4273);
nor U4960 (N_4960,N_4083,N_4389);
nor U4961 (N_4961,N_4364,N_4092);
or U4962 (N_4962,N_4328,N_4055);
or U4963 (N_4963,N_4268,N_4354);
or U4964 (N_4964,N_4297,N_4493);
and U4965 (N_4965,N_4239,N_4493);
nor U4966 (N_4966,N_4250,N_4473);
nor U4967 (N_4967,N_4077,N_4340);
nor U4968 (N_4968,N_4264,N_4069);
nor U4969 (N_4969,N_4215,N_4381);
nor U4970 (N_4970,N_4176,N_4224);
nor U4971 (N_4971,N_4252,N_4039);
and U4972 (N_4972,N_4056,N_4222);
xor U4973 (N_4973,N_4355,N_4098);
nor U4974 (N_4974,N_4007,N_4300);
and U4975 (N_4975,N_4266,N_4428);
xor U4976 (N_4976,N_4225,N_4425);
and U4977 (N_4977,N_4269,N_4404);
xor U4978 (N_4978,N_4449,N_4348);
nand U4979 (N_4979,N_4205,N_4136);
and U4980 (N_4980,N_4002,N_4060);
or U4981 (N_4981,N_4271,N_4021);
xnor U4982 (N_4982,N_4102,N_4432);
xnor U4983 (N_4983,N_4217,N_4442);
xnor U4984 (N_4984,N_4304,N_4241);
and U4985 (N_4985,N_4292,N_4382);
and U4986 (N_4986,N_4127,N_4314);
or U4987 (N_4987,N_4099,N_4036);
nor U4988 (N_4988,N_4045,N_4223);
and U4989 (N_4989,N_4490,N_4022);
or U4990 (N_4990,N_4285,N_4133);
and U4991 (N_4991,N_4055,N_4385);
xnor U4992 (N_4992,N_4099,N_4245);
or U4993 (N_4993,N_4045,N_4327);
nor U4994 (N_4994,N_4237,N_4384);
nand U4995 (N_4995,N_4003,N_4492);
xnor U4996 (N_4996,N_4313,N_4146);
nor U4997 (N_4997,N_4337,N_4129);
nor U4998 (N_4998,N_4333,N_4383);
and U4999 (N_4999,N_4395,N_4116);
or U5000 (N_5000,N_4902,N_4558);
and U5001 (N_5001,N_4709,N_4614);
nor U5002 (N_5002,N_4972,N_4710);
nor U5003 (N_5003,N_4875,N_4579);
or U5004 (N_5004,N_4743,N_4873);
nand U5005 (N_5005,N_4629,N_4949);
or U5006 (N_5006,N_4944,N_4570);
nand U5007 (N_5007,N_4728,N_4714);
or U5008 (N_5008,N_4699,N_4560);
nand U5009 (N_5009,N_4762,N_4565);
nand U5010 (N_5010,N_4853,N_4918);
nand U5011 (N_5011,N_4670,N_4954);
and U5012 (N_5012,N_4581,N_4755);
nor U5013 (N_5013,N_4955,N_4617);
and U5014 (N_5014,N_4790,N_4915);
and U5015 (N_5015,N_4910,N_4795);
and U5016 (N_5016,N_4635,N_4865);
or U5017 (N_5017,N_4885,N_4829);
nand U5018 (N_5018,N_4843,N_4845);
and U5019 (N_5019,N_4633,N_4940);
nor U5020 (N_5020,N_4807,N_4870);
xnor U5021 (N_5021,N_4936,N_4983);
or U5022 (N_5022,N_4832,N_4914);
or U5023 (N_5023,N_4527,N_4691);
nor U5024 (N_5024,N_4749,N_4968);
and U5025 (N_5025,N_4981,N_4596);
nor U5026 (N_5026,N_4545,N_4549);
nand U5027 (N_5027,N_4591,N_4592);
xnor U5028 (N_5028,N_4759,N_4995);
or U5029 (N_5029,N_4757,N_4788);
or U5030 (N_5030,N_4585,N_4830);
or U5031 (N_5031,N_4847,N_4530);
or U5032 (N_5032,N_4980,N_4756);
and U5033 (N_5033,N_4953,N_4882);
nor U5034 (N_5034,N_4842,N_4599);
or U5035 (N_5035,N_4645,N_4779);
nor U5036 (N_5036,N_4874,N_4838);
and U5037 (N_5037,N_4905,N_4957);
nor U5038 (N_5038,N_4822,N_4605);
nand U5039 (N_5039,N_4646,N_4977);
or U5040 (N_5040,N_4576,N_4719);
and U5041 (N_5041,N_4781,N_4868);
nand U5042 (N_5042,N_4886,N_4777);
nand U5043 (N_5043,N_4774,N_4741);
and U5044 (N_5044,N_4609,N_4907);
nor U5045 (N_5045,N_4583,N_4960);
xor U5046 (N_5046,N_4770,N_4990);
nor U5047 (N_5047,N_4715,N_4852);
nor U5048 (N_5048,N_4884,N_4809);
or U5049 (N_5049,N_4982,N_4651);
or U5050 (N_5050,N_4932,N_4831);
nor U5051 (N_5051,N_4751,N_4880);
nor U5052 (N_5052,N_4825,N_4567);
and U5053 (N_5053,N_4791,N_4950);
and U5054 (N_5054,N_4561,N_4912);
nor U5055 (N_5055,N_4978,N_4604);
and U5056 (N_5056,N_4523,N_4803);
nand U5057 (N_5057,N_4542,N_4533);
nand U5058 (N_5058,N_4712,N_4909);
nor U5059 (N_5059,N_4817,N_4679);
nor U5060 (N_5060,N_4696,N_4532);
nor U5061 (N_5061,N_4804,N_4575);
nor U5062 (N_5062,N_4922,N_4738);
xnor U5063 (N_5063,N_4761,N_4685);
nor U5064 (N_5064,N_4616,N_4716);
xor U5065 (N_5065,N_4623,N_4535);
xor U5066 (N_5066,N_4725,N_4971);
nand U5067 (N_5067,N_4890,N_4858);
or U5068 (N_5068,N_4962,N_4703);
nand U5069 (N_5069,N_4734,N_4956);
or U5070 (N_5070,N_4638,N_4811);
and U5071 (N_5071,N_4826,N_4684);
nor U5072 (N_5072,N_4720,N_4776);
nor U5073 (N_5073,N_4548,N_4833);
nor U5074 (N_5074,N_4933,N_4640);
nor U5075 (N_5075,N_4667,N_4601);
xnor U5076 (N_5076,N_4666,N_4544);
nor U5077 (N_5077,N_4913,N_4669);
nand U5078 (N_5078,N_4677,N_4692);
and U5079 (N_5079,N_4773,N_4924);
nand U5080 (N_5080,N_4554,N_4893);
nand U5081 (N_5081,N_4784,N_4694);
xnor U5082 (N_5082,N_4767,N_4552);
and U5083 (N_5083,N_4577,N_4597);
or U5084 (N_5084,N_4979,N_4615);
and U5085 (N_5085,N_4816,N_4919);
and U5086 (N_5086,N_4578,N_4580);
nand U5087 (N_5087,N_4555,N_4920);
or U5088 (N_5088,N_4938,N_4763);
nor U5089 (N_5089,N_4840,N_4587);
or U5090 (N_5090,N_4753,N_4937);
nand U5091 (N_5091,N_4985,N_4780);
nor U5092 (N_5092,N_4748,N_4705);
xnor U5093 (N_5093,N_4974,N_4557);
or U5094 (N_5094,N_4624,N_4721);
and U5095 (N_5095,N_4675,N_4904);
or U5096 (N_5096,N_4765,N_4808);
or U5097 (N_5097,N_4824,N_4900);
xnor U5098 (N_5098,N_4989,N_4518);
or U5099 (N_5099,N_4752,N_4665);
nand U5100 (N_5100,N_4819,N_4908);
or U5101 (N_5101,N_4639,N_4512);
nor U5102 (N_5102,N_4730,N_4772);
or U5103 (N_5103,N_4986,N_4903);
nor U5104 (N_5104,N_4792,N_4859);
and U5105 (N_5105,N_4998,N_4747);
nand U5106 (N_5106,N_4637,N_4655);
and U5107 (N_5107,N_4556,N_4939);
nor U5108 (N_5108,N_4931,N_4887);
and U5109 (N_5109,N_4879,N_4595);
nand U5110 (N_5110,N_4851,N_4671);
or U5111 (N_5111,N_4872,N_4727);
nor U5112 (N_5112,N_4511,N_4729);
nand U5113 (N_5113,N_4706,N_4610);
or U5114 (N_5114,N_4618,N_4657);
and U5115 (N_5115,N_4997,N_4783);
nand U5116 (N_5116,N_4820,N_4628);
nor U5117 (N_5117,N_4963,N_4547);
and U5118 (N_5118,N_4634,N_4625);
nand U5119 (N_5119,N_4508,N_4534);
or U5120 (N_5120,N_4967,N_4891);
xnor U5121 (N_5121,N_4786,N_4854);
nand U5122 (N_5122,N_4863,N_4877);
xor U5123 (N_5123,N_4517,N_4794);
nand U5124 (N_5124,N_4674,N_4844);
nand U5125 (N_5125,N_4976,N_4500);
and U5126 (N_5126,N_4573,N_4531);
or U5127 (N_5127,N_4515,N_4975);
nand U5128 (N_5128,N_4505,N_4641);
nand U5129 (N_5129,N_4537,N_4805);
nand U5130 (N_5130,N_4564,N_4810);
and U5131 (N_5131,N_4524,N_4590);
xor U5132 (N_5132,N_4529,N_4574);
or U5133 (N_5133,N_4526,N_4506);
and U5134 (N_5134,N_4946,N_4837);
nor U5135 (N_5135,N_4821,N_4588);
and U5136 (N_5136,N_4806,N_4660);
and U5137 (N_5137,N_4562,N_4966);
nand U5138 (N_5138,N_4627,N_4622);
xor U5139 (N_5139,N_4649,N_4855);
or U5140 (N_5140,N_4673,N_4503);
nand U5141 (N_5141,N_4563,N_4881);
nor U5142 (N_5142,N_4945,N_4961);
and U5143 (N_5143,N_4815,N_4582);
nand U5144 (N_5144,N_4690,N_4536);
or U5145 (N_5145,N_4896,N_4841);
and U5146 (N_5146,N_4867,N_4906);
nor U5147 (N_5147,N_4718,N_4839);
nand U5148 (N_5148,N_4735,N_4688);
nor U5149 (N_5149,N_4731,N_4593);
nand U5150 (N_5150,N_4869,N_4540);
nand U5151 (N_5151,N_4658,N_4823);
nor U5152 (N_5152,N_4519,N_4711);
nor U5153 (N_5153,N_4857,N_4899);
nand U5154 (N_5154,N_4764,N_4916);
or U5155 (N_5155,N_4636,N_4994);
and U5156 (N_5156,N_4693,N_4668);
nor U5157 (N_5157,N_4796,N_4828);
and U5158 (N_5158,N_4894,N_4612);
or U5159 (N_5159,N_4987,N_4594);
and U5160 (N_5160,N_4513,N_4921);
or U5161 (N_5161,N_4850,N_4964);
or U5162 (N_5162,N_4521,N_4745);
nand U5163 (N_5163,N_4686,N_4750);
nor U5164 (N_5164,N_4608,N_4754);
nor U5165 (N_5165,N_4586,N_4959);
nor U5166 (N_5166,N_4736,N_4947);
and U5167 (N_5167,N_4973,N_4943);
or U5168 (N_5168,N_4510,N_4771);
nor U5169 (N_5169,N_4680,N_4801);
nand U5170 (N_5170,N_4707,N_4871);
nand U5171 (N_5171,N_4895,N_4621);
or U5172 (N_5172,N_4861,N_4572);
or U5173 (N_5173,N_4584,N_4571);
and U5174 (N_5174,N_4948,N_4889);
nand U5175 (N_5175,N_4704,N_4930);
nand U5176 (N_5176,N_4659,N_4897);
or U5177 (N_5177,N_4793,N_4901);
or U5178 (N_5178,N_4746,N_4952);
nor U5179 (N_5179,N_4923,N_4726);
or U5180 (N_5180,N_4797,N_4543);
nand U5181 (N_5181,N_4864,N_4768);
and U5182 (N_5182,N_4883,N_4514);
and U5183 (N_5183,N_4769,N_4662);
or U5184 (N_5184,N_4802,N_4520);
or U5185 (N_5185,N_4509,N_4969);
and U5186 (N_5186,N_4708,N_4700);
and U5187 (N_5187,N_4999,N_4733);
and U5188 (N_5188,N_4856,N_4800);
nor U5189 (N_5189,N_4559,N_4606);
nor U5190 (N_5190,N_4501,N_4504);
or U5191 (N_5191,N_4528,N_4935);
and U5192 (N_5192,N_4663,N_4713);
or U5193 (N_5193,N_4525,N_4647);
or U5194 (N_5194,N_4502,N_4568);
nor U5195 (N_5195,N_4775,N_4827);
or U5196 (N_5196,N_4553,N_4516);
nor U5197 (N_5197,N_4611,N_4744);
nand U5198 (N_5198,N_4522,N_4598);
nand U5199 (N_5199,N_4507,N_4613);
and U5200 (N_5200,N_4834,N_4818);
nand U5201 (N_5201,N_4812,N_4551);
xor U5202 (N_5202,N_4654,N_4782);
nor U5203 (N_5203,N_4607,N_4799);
and U5204 (N_5204,N_4742,N_4992);
and U5205 (N_5205,N_4724,N_4689);
or U5206 (N_5206,N_4603,N_4723);
nand U5207 (N_5207,N_4630,N_4911);
or U5208 (N_5208,N_4737,N_4653);
nand U5209 (N_5209,N_4626,N_4740);
nor U5210 (N_5210,N_4789,N_4766);
nor U5211 (N_5211,N_4546,N_4785);
nor U5212 (N_5212,N_4849,N_4569);
and U5213 (N_5213,N_4717,N_4848);
nand U5214 (N_5214,N_4778,N_4566);
and U5215 (N_5215,N_4701,N_4928);
and U5216 (N_5216,N_4996,N_4836);
or U5217 (N_5217,N_4652,N_4951);
or U5218 (N_5218,N_4958,N_4934);
and U5219 (N_5219,N_4929,N_4732);
and U5220 (N_5220,N_4642,N_4619);
xnor U5221 (N_5221,N_4620,N_4683);
and U5222 (N_5222,N_4602,N_4860);
or U5223 (N_5223,N_4664,N_4862);
xnor U5224 (N_5224,N_4697,N_4702);
nor U5225 (N_5225,N_4917,N_4682);
or U5226 (N_5226,N_4927,N_4991);
nor U5227 (N_5227,N_4984,N_4835);
or U5228 (N_5228,N_4876,N_4589);
and U5229 (N_5229,N_4941,N_4798);
nor U5230 (N_5230,N_4787,N_4550);
or U5231 (N_5231,N_4648,N_4925);
or U5232 (N_5232,N_4878,N_4988);
and U5233 (N_5233,N_4898,N_4993);
xor U5234 (N_5234,N_4539,N_4676);
and U5235 (N_5235,N_4866,N_4698);
nor U5236 (N_5236,N_4965,N_4695);
xnor U5237 (N_5237,N_4644,N_4631);
and U5238 (N_5238,N_4681,N_4650);
or U5239 (N_5239,N_4632,N_4926);
or U5240 (N_5240,N_4656,N_4678);
nor U5241 (N_5241,N_4760,N_4814);
and U5242 (N_5242,N_4600,N_4538);
nand U5243 (N_5243,N_4687,N_4892);
and U5244 (N_5244,N_4722,N_4541);
nor U5245 (N_5245,N_4758,N_4739);
or U5246 (N_5246,N_4643,N_4672);
and U5247 (N_5247,N_4888,N_4970);
nand U5248 (N_5248,N_4813,N_4942);
nand U5249 (N_5249,N_4661,N_4846);
or U5250 (N_5250,N_4590,N_4545);
and U5251 (N_5251,N_4620,N_4950);
nor U5252 (N_5252,N_4888,N_4960);
or U5253 (N_5253,N_4848,N_4982);
nor U5254 (N_5254,N_4513,N_4851);
nor U5255 (N_5255,N_4651,N_4532);
and U5256 (N_5256,N_4858,N_4839);
or U5257 (N_5257,N_4667,N_4876);
nand U5258 (N_5258,N_4810,N_4768);
nor U5259 (N_5259,N_4606,N_4777);
and U5260 (N_5260,N_4700,N_4772);
and U5261 (N_5261,N_4986,N_4621);
nand U5262 (N_5262,N_4919,N_4819);
nand U5263 (N_5263,N_4813,N_4827);
or U5264 (N_5264,N_4961,N_4646);
nor U5265 (N_5265,N_4500,N_4734);
or U5266 (N_5266,N_4629,N_4988);
nor U5267 (N_5267,N_4926,N_4895);
xnor U5268 (N_5268,N_4642,N_4723);
nand U5269 (N_5269,N_4776,N_4524);
nand U5270 (N_5270,N_4982,N_4877);
nor U5271 (N_5271,N_4886,N_4783);
nor U5272 (N_5272,N_4887,N_4658);
or U5273 (N_5273,N_4722,N_4735);
nand U5274 (N_5274,N_4566,N_4711);
nand U5275 (N_5275,N_4942,N_4599);
nor U5276 (N_5276,N_4912,N_4960);
and U5277 (N_5277,N_4541,N_4947);
nor U5278 (N_5278,N_4847,N_4571);
and U5279 (N_5279,N_4608,N_4520);
nor U5280 (N_5280,N_4826,N_4914);
nor U5281 (N_5281,N_4576,N_4749);
nor U5282 (N_5282,N_4618,N_4671);
and U5283 (N_5283,N_4891,N_4766);
xnor U5284 (N_5284,N_4598,N_4874);
nand U5285 (N_5285,N_4607,N_4646);
and U5286 (N_5286,N_4837,N_4674);
and U5287 (N_5287,N_4967,N_4775);
nor U5288 (N_5288,N_4805,N_4698);
or U5289 (N_5289,N_4512,N_4606);
nand U5290 (N_5290,N_4746,N_4908);
or U5291 (N_5291,N_4898,N_4907);
nor U5292 (N_5292,N_4849,N_4697);
nand U5293 (N_5293,N_4744,N_4678);
nor U5294 (N_5294,N_4916,N_4897);
or U5295 (N_5295,N_4561,N_4513);
xor U5296 (N_5296,N_4938,N_4936);
nand U5297 (N_5297,N_4547,N_4654);
nand U5298 (N_5298,N_4671,N_4705);
nor U5299 (N_5299,N_4958,N_4776);
nand U5300 (N_5300,N_4721,N_4762);
nor U5301 (N_5301,N_4846,N_4921);
or U5302 (N_5302,N_4779,N_4531);
or U5303 (N_5303,N_4623,N_4916);
and U5304 (N_5304,N_4866,N_4977);
nor U5305 (N_5305,N_4875,N_4962);
xnor U5306 (N_5306,N_4906,N_4730);
and U5307 (N_5307,N_4567,N_4629);
nand U5308 (N_5308,N_4608,N_4750);
and U5309 (N_5309,N_4899,N_4720);
xor U5310 (N_5310,N_4616,N_4775);
nand U5311 (N_5311,N_4737,N_4986);
or U5312 (N_5312,N_4859,N_4505);
and U5313 (N_5313,N_4746,N_4519);
and U5314 (N_5314,N_4865,N_4711);
or U5315 (N_5315,N_4635,N_4531);
nand U5316 (N_5316,N_4772,N_4643);
nor U5317 (N_5317,N_4672,N_4698);
and U5318 (N_5318,N_4699,N_4773);
nor U5319 (N_5319,N_4661,N_4504);
and U5320 (N_5320,N_4761,N_4756);
or U5321 (N_5321,N_4941,N_4853);
nand U5322 (N_5322,N_4651,N_4629);
nor U5323 (N_5323,N_4985,N_4581);
or U5324 (N_5324,N_4862,N_4984);
or U5325 (N_5325,N_4538,N_4598);
and U5326 (N_5326,N_4699,N_4656);
nand U5327 (N_5327,N_4902,N_4747);
and U5328 (N_5328,N_4785,N_4833);
or U5329 (N_5329,N_4952,N_4540);
or U5330 (N_5330,N_4546,N_4566);
xnor U5331 (N_5331,N_4774,N_4876);
xnor U5332 (N_5332,N_4799,N_4836);
nor U5333 (N_5333,N_4813,N_4859);
or U5334 (N_5334,N_4768,N_4609);
nand U5335 (N_5335,N_4673,N_4603);
and U5336 (N_5336,N_4994,N_4787);
or U5337 (N_5337,N_4510,N_4866);
xor U5338 (N_5338,N_4920,N_4830);
and U5339 (N_5339,N_4806,N_4994);
nor U5340 (N_5340,N_4709,N_4618);
nor U5341 (N_5341,N_4626,N_4714);
nor U5342 (N_5342,N_4714,N_4974);
nand U5343 (N_5343,N_4735,N_4632);
xor U5344 (N_5344,N_4722,N_4942);
nor U5345 (N_5345,N_4710,N_4786);
and U5346 (N_5346,N_4502,N_4746);
and U5347 (N_5347,N_4958,N_4896);
or U5348 (N_5348,N_4721,N_4583);
nor U5349 (N_5349,N_4596,N_4649);
xnor U5350 (N_5350,N_4814,N_4970);
nor U5351 (N_5351,N_4828,N_4721);
or U5352 (N_5352,N_4578,N_4872);
and U5353 (N_5353,N_4554,N_4626);
or U5354 (N_5354,N_4585,N_4551);
and U5355 (N_5355,N_4725,N_4765);
nor U5356 (N_5356,N_4559,N_4519);
and U5357 (N_5357,N_4925,N_4778);
or U5358 (N_5358,N_4918,N_4779);
and U5359 (N_5359,N_4513,N_4896);
nand U5360 (N_5360,N_4580,N_4647);
and U5361 (N_5361,N_4787,N_4841);
xor U5362 (N_5362,N_4968,N_4931);
nor U5363 (N_5363,N_4806,N_4815);
and U5364 (N_5364,N_4758,N_4859);
nand U5365 (N_5365,N_4975,N_4745);
and U5366 (N_5366,N_4744,N_4880);
xnor U5367 (N_5367,N_4891,N_4636);
nand U5368 (N_5368,N_4578,N_4597);
nand U5369 (N_5369,N_4638,N_4597);
nand U5370 (N_5370,N_4594,N_4542);
or U5371 (N_5371,N_4980,N_4644);
xor U5372 (N_5372,N_4957,N_4550);
and U5373 (N_5373,N_4639,N_4973);
or U5374 (N_5374,N_4518,N_4626);
nand U5375 (N_5375,N_4806,N_4778);
nand U5376 (N_5376,N_4858,N_4738);
xnor U5377 (N_5377,N_4933,N_4835);
and U5378 (N_5378,N_4722,N_4743);
and U5379 (N_5379,N_4699,N_4635);
nand U5380 (N_5380,N_4702,N_4650);
or U5381 (N_5381,N_4770,N_4975);
or U5382 (N_5382,N_4948,N_4731);
nor U5383 (N_5383,N_4770,N_4900);
xnor U5384 (N_5384,N_4808,N_4905);
xor U5385 (N_5385,N_4878,N_4915);
nand U5386 (N_5386,N_4741,N_4955);
nand U5387 (N_5387,N_4689,N_4815);
nand U5388 (N_5388,N_4743,N_4574);
nor U5389 (N_5389,N_4764,N_4720);
nor U5390 (N_5390,N_4867,N_4972);
and U5391 (N_5391,N_4747,N_4549);
nand U5392 (N_5392,N_4927,N_4701);
nand U5393 (N_5393,N_4510,N_4621);
and U5394 (N_5394,N_4649,N_4922);
xnor U5395 (N_5395,N_4704,N_4654);
and U5396 (N_5396,N_4745,N_4814);
nor U5397 (N_5397,N_4594,N_4856);
or U5398 (N_5398,N_4845,N_4991);
nand U5399 (N_5399,N_4529,N_4692);
nand U5400 (N_5400,N_4888,N_4988);
nand U5401 (N_5401,N_4871,N_4559);
or U5402 (N_5402,N_4973,N_4805);
nand U5403 (N_5403,N_4829,N_4679);
nor U5404 (N_5404,N_4941,N_4925);
nor U5405 (N_5405,N_4627,N_4824);
nand U5406 (N_5406,N_4937,N_4665);
nor U5407 (N_5407,N_4880,N_4872);
and U5408 (N_5408,N_4674,N_4805);
nor U5409 (N_5409,N_4761,N_4949);
nor U5410 (N_5410,N_4564,N_4700);
nand U5411 (N_5411,N_4973,N_4662);
nor U5412 (N_5412,N_4602,N_4552);
nor U5413 (N_5413,N_4889,N_4596);
nand U5414 (N_5414,N_4930,N_4586);
nand U5415 (N_5415,N_4813,N_4596);
and U5416 (N_5416,N_4828,N_4540);
or U5417 (N_5417,N_4525,N_4966);
or U5418 (N_5418,N_4742,N_4573);
nand U5419 (N_5419,N_4852,N_4565);
nor U5420 (N_5420,N_4758,N_4672);
nand U5421 (N_5421,N_4766,N_4778);
nor U5422 (N_5422,N_4645,N_4825);
and U5423 (N_5423,N_4931,N_4609);
and U5424 (N_5424,N_4825,N_4694);
nor U5425 (N_5425,N_4585,N_4664);
nand U5426 (N_5426,N_4657,N_4856);
nor U5427 (N_5427,N_4603,N_4706);
and U5428 (N_5428,N_4795,N_4640);
xor U5429 (N_5429,N_4958,N_4654);
nand U5430 (N_5430,N_4600,N_4648);
and U5431 (N_5431,N_4704,N_4510);
nor U5432 (N_5432,N_4584,N_4802);
or U5433 (N_5433,N_4948,N_4961);
nor U5434 (N_5434,N_4816,N_4700);
nor U5435 (N_5435,N_4920,N_4671);
nor U5436 (N_5436,N_4667,N_4856);
and U5437 (N_5437,N_4745,N_4882);
or U5438 (N_5438,N_4803,N_4948);
and U5439 (N_5439,N_4915,N_4798);
nand U5440 (N_5440,N_4720,N_4725);
and U5441 (N_5441,N_4854,N_4771);
and U5442 (N_5442,N_4832,N_4801);
or U5443 (N_5443,N_4799,N_4677);
nor U5444 (N_5444,N_4838,N_4505);
and U5445 (N_5445,N_4627,N_4936);
or U5446 (N_5446,N_4987,N_4778);
and U5447 (N_5447,N_4542,N_4655);
nor U5448 (N_5448,N_4968,N_4897);
nor U5449 (N_5449,N_4756,N_4864);
xnor U5450 (N_5450,N_4603,N_4620);
and U5451 (N_5451,N_4794,N_4519);
and U5452 (N_5452,N_4809,N_4881);
and U5453 (N_5453,N_4644,N_4592);
or U5454 (N_5454,N_4629,N_4799);
or U5455 (N_5455,N_4979,N_4818);
xnor U5456 (N_5456,N_4520,N_4623);
nor U5457 (N_5457,N_4598,N_4648);
nand U5458 (N_5458,N_4677,N_4602);
xnor U5459 (N_5459,N_4880,N_4732);
or U5460 (N_5460,N_4668,N_4896);
nand U5461 (N_5461,N_4562,N_4761);
or U5462 (N_5462,N_4735,N_4640);
or U5463 (N_5463,N_4865,N_4966);
and U5464 (N_5464,N_4847,N_4792);
nor U5465 (N_5465,N_4678,N_4971);
and U5466 (N_5466,N_4828,N_4557);
xor U5467 (N_5467,N_4933,N_4728);
nor U5468 (N_5468,N_4734,N_4982);
xor U5469 (N_5469,N_4587,N_4855);
and U5470 (N_5470,N_4802,N_4852);
and U5471 (N_5471,N_4986,N_4796);
nor U5472 (N_5472,N_4720,N_4607);
and U5473 (N_5473,N_4921,N_4733);
xor U5474 (N_5474,N_4772,N_4726);
nor U5475 (N_5475,N_4797,N_4574);
nand U5476 (N_5476,N_4815,N_4520);
nand U5477 (N_5477,N_4686,N_4730);
nor U5478 (N_5478,N_4925,N_4773);
nor U5479 (N_5479,N_4693,N_4948);
and U5480 (N_5480,N_4800,N_4783);
nor U5481 (N_5481,N_4965,N_4822);
or U5482 (N_5482,N_4987,N_4985);
nor U5483 (N_5483,N_4513,N_4969);
nor U5484 (N_5484,N_4621,N_4912);
xnor U5485 (N_5485,N_4513,N_4987);
nand U5486 (N_5486,N_4717,N_4720);
and U5487 (N_5487,N_4833,N_4764);
xor U5488 (N_5488,N_4791,N_4639);
and U5489 (N_5489,N_4583,N_4534);
or U5490 (N_5490,N_4851,N_4782);
nand U5491 (N_5491,N_4819,N_4886);
nor U5492 (N_5492,N_4826,N_4832);
nor U5493 (N_5493,N_4730,N_4629);
or U5494 (N_5494,N_4710,N_4686);
nor U5495 (N_5495,N_4652,N_4782);
or U5496 (N_5496,N_4609,N_4631);
nor U5497 (N_5497,N_4905,N_4700);
xnor U5498 (N_5498,N_4924,N_4919);
and U5499 (N_5499,N_4846,N_4752);
nand U5500 (N_5500,N_5238,N_5357);
nand U5501 (N_5501,N_5099,N_5186);
nor U5502 (N_5502,N_5430,N_5338);
and U5503 (N_5503,N_5497,N_5282);
and U5504 (N_5504,N_5489,N_5008);
nor U5505 (N_5505,N_5457,N_5261);
or U5506 (N_5506,N_5265,N_5244);
nand U5507 (N_5507,N_5358,N_5406);
or U5508 (N_5508,N_5336,N_5355);
or U5509 (N_5509,N_5475,N_5060);
and U5510 (N_5510,N_5254,N_5288);
and U5511 (N_5511,N_5450,N_5108);
and U5512 (N_5512,N_5226,N_5204);
and U5513 (N_5513,N_5347,N_5296);
xnor U5514 (N_5514,N_5456,N_5028);
nor U5515 (N_5515,N_5268,N_5441);
nand U5516 (N_5516,N_5321,N_5319);
or U5517 (N_5517,N_5427,N_5266);
or U5518 (N_5518,N_5216,N_5146);
xor U5519 (N_5519,N_5317,N_5198);
and U5520 (N_5520,N_5148,N_5245);
or U5521 (N_5521,N_5260,N_5182);
nor U5522 (N_5522,N_5122,N_5371);
or U5523 (N_5523,N_5442,N_5435);
xor U5524 (N_5524,N_5169,N_5256);
and U5525 (N_5525,N_5144,N_5119);
nand U5526 (N_5526,N_5200,N_5395);
or U5527 (N_5527,N_5318,N_5123);
nor U5528 (N_5528,N_5249,N_5298);
nor U5529 (N_5529,N_5454,N_5076);
nor U5530 (N_5530,N_5209,N_5440);
or U5531 (N_5531,N_5025,N_5384);
xor U5532 (N_5532,N_5356,N_5477);
nor U5533 (N_5533,N_5412,N_5041);
nor U5534 (N_5534,N_5037,N_5488);
and U5535 (N_5535,N_5141,N_5227);
nor U5536 (N_5536,N_5402,N_5349);
and U5537 (N_5537,N_5431,N_5313);
xor U5538 (N_5538,N_5149,N_5071);
or U5539 (N_5539,N_5068,N_5368);
and U5540 (N_5540,N_5409,N_5214);
nand U5541 (N_5541,N_5029,N_5424);
xor U5542 (N_5542,N_5417,N_5155);
nor U5543 (N_5543,N_5063,N_5210);
nor U5544 (N_5544,N_5075,N_5309);
nor U5545 (N_5545,N_5375,N_5276);
and U5546 (N_5546,N_5138,N_5414);
or U5547 (N_5547,N_5135,N_5040);
and U5548 (N_5548,N_5125,N_5228);
and U5549 (N_5549,N_5251,N_5449);
or U5550 (N_5550,N_5102,N_5364);
nor U5551 (N_5551,N_5096,N_5013);
and U5552 (N_5552,N_5308,N_5429);
nor U5553 (N_5553,N_5280,N_5448);
nand U5554 (N_5554,N_5085,N_5324);
nand U5555 (N_5555,N_5295,N_5039);
and U5556 (N_5556,N_5016,N_5460);
nor U5557 (N_5557,N_5162,N_5258);
and U5558 (N_5558,N_5496,N_5436);
nor U5559 (N_5559,N_5378,N_5354);
or U5560 (N_5560,N_5168,N_5001);
or U5561 (N_5561,N_5136,N_5049);
xnor U5562 (N_5562,N_5199,N_5161);
and U5563 (N_5563,N_5381,N_5328);
nand U5564 (N_5564,N_5474,N_5084);
nor U5565 (N_5565,N_5118,N_5332);
nand U5566 (N_5566,N_5438,N_5339);
and U5567 (N_5567,N_5337,N_5445);
and U5568 (N_5568,N_5444,N_5153);
nand U5569 (N_5569,N_5274,N_5187);
xor U5570 (N_5570,N_5472,N_5181);
or U5571 (N_5571,N_5425,N_5124);
nor U5572 (N_5572,N_5294,N_5112);
and U5573 (N_5573,N_5150,N_5326);
or U5574 (N_5574,N_5064,N_5189);
nand U5575 (N_5575,N_5252,N_5396);
and U5576 (N_5576,N_5233,N_5316);
nand U5577 (N_5577,N_5281,N_5463);
or U5578 (N_5578,N_5493,N_5062);
or U5579 (N_5579,N_5273,N_5481);
or U5580 (N_5580,N_5482,N_5270);
and U5581 (N_5581,N_5272,N_5009);
nor U5582 (N_5582,N_5163,N_5320);
nand U5583 (N_5583,N_5301,N_5439);
xor U5584 (N_5584,N_5152,N_5235);
xor U5585 (N_5585,N_5134,N_5107);
or U5586 (N_5586,N_5139,N_5348);
nor U5587 (N_5587,N_5290,N_5340);
and U5588 (N_5588,N_5329,N_5092);
or U5589 (N_5589,N_5042,N_5361);
nand U5590 (N_5590,N_5129,N_5079);
nand U5591 (N_5591,N_5059,N_5106);
xor U5592 (N_5592,N_5372,N_5394);
or U5593 (N_5593,N_5377,N_5302);
and U5594 (N_5594,N_5350,N_5014);
or U5595 (N_5595,N_5067,N_5094);
and U5596 (N_5596,N_5154,N_5173);
or U5597 (N_5597,N_5243,N_5022);
and U5598 (N_5598,N_5021,N_5159);
nor U5599 (N_5599,N_5185,N_5048);
nand U5600 (N_5600,N_5027,N_5393);
nor U5601 (N_5601,N_5432,N_5299);
and U5602 (N_5602,N_5117,N_5101);
and U5603 (N_5603,N_5081,N_5002);
or U5604 (N_5604,N_5277,N_5495);
and U5605 (N_5605,N_5083,N_5053);
or U5606 (N_5606,N_5422,N_5470);
and U5607 (N_5607,N_5334,N_5434);
nand U5608 (N_5608,N_5240,N_5116);
nor U5609 (N_5609,N_5088,N_5137);
and U5610 (N_5610,N_5271,N_5351);
and U5611 (N_5611,N_5065,N_5177);
and U5612 (N_5612,N_5145,N_5360);
or U5613 (N_5613,N_5423,N_5160);
nor U5614 (N_5614,N_5213,N_5056);
and U5615 (N_5615,N_5373,N_5218);
nor U5616 (N_5616,N_5389,N_5201);
nand U5617 (N_5617,N_5484,N_5415);
nor U5618 (N_5618,N_5003,N_5476);
or U5619 (N_5619,N_5247,N_5283);
xnor U5620 (N_5620,N_5379,N_5366);
or U5621 (N_5621,N_5494,N_5212);
nand U5622 (N_5622,N_5090,N_5312);
or U5623 (N_5623,N_5420,N_5012);
or U5624 (N_5624,N_5109,N_5115);
nand U5625 (N_5625,N_5050,N_5365);
or U5626 (N_5626,N_5331,N_5073);
nor U5627 (N_5627,N_5284,N_5446);
nor U5628 (N_5628,N_5239,N_5230);
or U5629 (N_5629,N_5246,N_5253);
nand U5630 (N_5630,N_5224,N_5074);
nand U5631 (N_5631,N_5262,N_5275);
and U5632 (N_5632,N_5399,N_5492);
and U5633 (N_5633,N_5468,N_5353);
nand U5634 (N_5634,N_5297,N_5419);
xor U5635 (N_5635,N_5188,N_5404);
nand U5636 (N_5636,N_5370,N_5121);
nand U5637 (N_5637,N_5411,N_5172);
or U5638 (N_5638,N_5267,N_5405);
nand U5639 (N_5639,N_5443,N_5259);
nor U5640 (N_5640,N_5231,N_5057);
or U5641 (N_5641,N_5487,N_5447);
nor U5642 (N_5642,N_5176,N_5195);
or U5643 (N_5643,N_5193,N_5359);
nand U5644 (N_5644,N_5385,N_5098);
nand U5645 (N_5645,N_5292,N_5498);
and U5646 (N_5646,N_5306,N_5089);
xnor U5647 (N_5647,N_5220,N_5343);
xnor U5648 (N_5648,N_5207,N_5352);
and U5649 (N_5649,N_5234,N_5410);
or U5650 (N_5650,N_5369,N_5325);
xnor U5651 (N_5651,N_5330,N_5208);
xnor U5652 (N_5652,N_5196,N_5026);
or U5653 (N_5653,N_5458,N_5314);
or U5654 (N_5654,N_5077,N_5278);
nor U5655 (N_5655,N_5011,N_5263);
nor U5656 (N_5656,N_5491,N_5054);
nand U5657 (N_5657,N_5024,N_5130);
xnor U5658 (N_5658,N_5034,N_5390);
nand U5659 (N_5659,N_5175,N_5030);
or U5660 (N_5660,N_5225,N_5242);
nand U5661 (N_5661,N_5382,N_5191);
nand U5662 (N_5662,N_5279,N_5202);
and U5663 (N_5663,N_5052,N_5408);
and U5664 (N_5664,N_5205,N_5156);
nand U5665 (N_5665,N_5069,N_5322);
or U5666 (N_5666,N_5327,N_5237);
nand U5667 (N_5667,N_5223,N_5221);
nand U5668 (N_5668,N_5416,N_5219);
or U5669 (N_5669,N_5113,N_5418);
and U5670 (N_5670,N_5211,N_5180);
nor U5671 (N_5671,N_5206,N_5407);
nand U5672 (N_5672,N_5105,N_5104);
nand U5673 (N_5673,N_5035,N_5392);
and U5674 (N_5674,N_5165,N_5248);
nand U5675 (N_5675,N_5362,N_5315);
nand U5676 (N_5676,N_5387,N_5033);
nand U5677 (N_5677,N_5401,N_5044);
nor U5678 (N_5678,N_5192,N_5335);
xnor U5679 (N_5679,N_5000,N_5178);
nand U5680 (N_5680,N_5143,N_5363);
and U5681 (N_5681,N_5421,N_5131);
and U5682 (N_5682,N_5391,N_5015);
nand U5683 (N_5683,N_5197,N_5342);
and U5684 (N_5684,N_5264,N_5287);
nor U5685 (N_5685,N_5157,N_5045);
nor U5686 (N_5686,N_5483,N_5166);
and U5687 (N_5687,N_5344,N_5170);
and U5688 (N_5688,N_5469,N_5091);
nand U5689 (N_5689,N_5017,N_5473);
or U5690 (N_5690,N_5093,N_5183);
nand U5691 (N_5691,N_5459,N_5031);
xnor U5692 (N_5692,N_5451,N_5462);
nand U5693 (N_5693,N_5479,N_5023);
or U5694 (N_5694,N_5464,N_5303);
nor U5695 (N_5695,N_5043,N_5367);
and U5696 (N_5696,N_5386,N_5127);
and U5697 (N_5697,N_5466,N_5413);
nor U5698 (N_5698,N_5380,N_5285);
and U5699 (N_5699,N_5100,N_5304);
or U5700 (N_5700,N_5151,N_5307);
or U5701 (N_5701,N_5480,N_5485);
xor U5702 (N_5702,N_5293,N_5341);
nand U5703 (N_5703,N_5215,N_5465);
nand U5704 (N_5704,N_5478,N_5499);
nand U5705 (N_5705,N_5428,N_5066);
xor U5706 (N_5706,N_5374,N_5055);
nor U5707 (N_5707,N_5376,N_5158);
and U5708 (N_5708,N_5222,N_5019);
and U5709 (N_5709,N_5147,N_5010);
nor U5710 (N_5710,N_5020,N_5467);
nor U5711 (N_5711,N_5036,N_5250);
xnor U5712 (N_5712,N_5080,N_5490);
and U5713 (N_5713,N_5078,N_5046);
or U5714 (N_5714,N_5142,N_5236);
or U5715 (N_5715,N_5133,N_5400);
nand U5716 (N_5716,N_5171,N_5452);
and U5717 (N_5717,N_5126,N_5005);
and U5718 (N_5718,N_5110,N_5286);
and U5719 (N_5719,N_5061,N_5289);
and U5720 (N_5720,N_5241,N_5403);
or U5721 (N_5721,N_5132,N_5194);
nand U5722 (N_5722,N_5203,N_5257);
nand U5723 (N_5723,N_5453,N_5310);
or U5724 (N_5724,N_5111,N_5388);
or U5725 (N_5725,N_5007,N_5140);
or U5726 (N_5726,N_5051,N_5269);
and U5727 (N_5727,N_5174,N_5006);
nand U5728 (N_5728,N_5311,N_5217);
nand U5729 (N_5729,N_5082,N_5333);
nor U5730 (N_5730,N_5167,N_5486);
nor U5731 (N_5731,N_5072,N_5103);
and U5732 (N_5732,N_5461,N_5164);
nor U5733 (N_5733,N_5179,N_5433);
nand U5734 (N_5734,N_5232,N_5426);
nand U5735 (N_5735,N_5004,N_5097);
and U5736 (N_5736,N_5087,N_5455);
xor U5737 (N_5737,N_5190,N_5305);
nor U5738 (N_5738,N_5058,N_5255);
nand U5739 (N_5739,N_5398,N_5095);
nand U5740 (N_5740,N_5128,N_5114);
nand U5741 (N_5741,N_5437,N_5383);
or U5742 (N_5742,N_5346,N_5471);
and U5743 (N_5743,N_5032,N_5323);
or U5744 (N_5744,N_5120,N_5184);
xnor U5745 (N_5745,N_5300,N_5397);
nor U5746 (N_5746,N_5038,N_5229);
and U5747 (N_5747,N_5086,N_5018);
nor U5748 (N_5748,N_5345,N_5047);
nor U5749 (N_5749,N_5291,N_5070);
or U5750 (N_5750,N_5487,N_5449);
nand U5751 (N_5751,N_5303,N_5224);
nor U5752 (N_5752,N_5225,N_5231);
nand U5753 (N_5753,N_5279,N_5324);
nand U5754 (N_5754,N_5468,N_5335);
and U5755 (N_5755,N_5098,N_5333);
or U5756 (N_5756,N_5435,N_5481);
or U5757 (N_5757,N_5397,N_5013);
nand U5758 (N_5758,N_5455,N_5145);
and U5759 (N_5759,N_5198,N_5025);
nor U5760 (N_5760,N_5279,N_5451);
or U5761 (N_5761,N_5329,N_5343);
and U5762 (N_5762,N_5025,N_5298);
and U5763 (N_5763,N_5182,N_5348);
nand U5764 (N_5764,N_5028,N_5158);
nor U5765 (N_5765,N_5286,N_5495);
and U5766 (N_5766,N_5181,N_5292);
and U5767 (N_5767,N_5449,N_5268);
nor U5768 (N_5768,N_5263,N_5300);
nand U5769 (N_5769,N_5310,N_5029);
nand U5770 (N_5770,N_5228,N_5430);
xnor U5771 (N_5771,N_5163,N_5491);
or U5772 (N_5772,N_5493,N_5031);
and U5773 (N_5773,N_5045,N_5287);
nor U5774 (N_5774,N_5105,N_5495);
nand U5775 (N_5775,N_5280,N_5313);
nor U5776 (N_5776,N_5455,N_5187);
nand U5777 (N_5777,N_5036,N_5372);
and U5778 (N_5778,N_5379,N_5497);
or U5779 (N_5779,N_5083,N_5273);
and U5780 (N_5780,N_5336,N_5216);
nor U5781 (N_5781,N_5253,N_5334);
or U5782 (N_5782,N_5304,N_5298);
nor U5783 (N_5783,N_5245,N_5174);
nand U5784 (N_5784,N_5344,N_5331);
nand U5785 (N_5785,N_5450,N_5046);
or U5786 (N_5786,N_5257,N_5371);
nor U5787 (N_5787,N_5260,N_5336);
nor U5788 (N_5788,N_5198,N_5024);
or U5789 (N_5789,N_5372,N_5278);
nor U5790 (N_5790,N_5371,N_5148);
xor U5791 (N_5791,N_5163,N_5166);
and U5792 (N_5792,N_5055,N_5435);
or U5793 (N_5793,N_5331,N_5176);
nand U5794 (N_5794,N_5053,N_5374);
and U5795 (N_5795,N_5016,N_5088);
xnor U5796 (N_5796,N_5369,N_5031);
or U5797 (N_5797,N_5237,N_5070);
and U5798 (N_5798,N_5306,N_5209);
and U5799 (N_5799,N_5385,N_5069);
nand U5800 (N_5800,N_5054,N_5116);
or U5801 (N_5801,N_5218,N_5107);
nor U5802 (N_5802,N_5462,N_5200);
nor U5803 (N_5803,N_5474,N_5195);
or U5804 (N_5804,N_5466,N_5087);
and U5805 (N_5805,N_5293,N_5246);
or U5806 (N_5806,N_5390,N_5202);
nor U5807 (N_5807,N_5032,N_5400);
nor U5808 (N_5808,N_5357,N_5342);
or U5809 (N_5809,N_5464,N_5382);
nor U5810 (N_5810,N_5401,N_5485);
or U5811 (N_5811,N_5101,N_5426);
nor U5812 (N_5812,N_5028,N_5269);
and U5813 (N_5813,N_5145,N_5068);
nor U5814 (N_5814,N_5288,N_5418);
or U5815 (N_5815,N_5017,N_5364);
nand U5816 (N_5816,N_5012,N_5075);
or U5817 (N_5817,N_5281,N_5347);
nor U5818 (N_5818,N_5228,N_5212);
nor U5819 (N_5819,N_5418,N_5332);
nand U5820 (N_5820,N_5006,N_5191);
nand U5821 (N_5821,N_5045,N_5096);
or U5822 (N_5822,N_5468,N_5028);
nor U5823 (N_5823,N_5384,N_5332);
and U5824 (N_5824,N_5016,N_5271);
or U5825 (N_5825,N_5472,N_5073);
or U5826 (N_5826,N_5273,N_5049);
nor U5827 (N_5827,N_5123,N_5208);
or U5828 (N_5828,N_5497,N_5271);
nor U5829 (N_5829,N_5212,N_5195);
or U5830 (N_5830,N_5281,N_5249);
and U5831 (N_5831,N_5294,N_5203);
xor U5832 (N_5832,N_5021,N_5322);
nand U5833 (N_5833,N_5459,N_5229);
or U5834 (N_5834,N_5208,N_5076);
nor U5835 (N_5835,N_5439,N_5021);
nor U5836 (N_5836,N_5119,N_5332);
and U5837 (N_5837,N_5021,N_5098);
nand U5838 (N_5838,N_5163,N_5058);
nand U5839 (N_5839,N_5350,N_5048);
nor U5840 (N_5840,N_5151,N_5284);
nor U5841 (N_5841,N_5454,N_5032);
nor U5842 (N_5842,N_5032,N_5161);
nand U5843 (N_5843,N_5257,N_5351);
or U5844 (N_5844,N_5498,N_5456);
xor U5845 (N_5845,N_5258,N_5317);
nor U5846 (N_5846,N_5149,N_5140);
nor U5847 (N_5847,N_5156,N_5001);
or U5848 (N_5848,N_5151,N_5437);
nand U5849 (N_5849,N_5177,N_5156);
or U5850 (N_5850,N_5127,N_5013);
nand U5851 (N_5851,N_5367,N_5007);
nand U5852 (N_5852,N_5044,N_5209);
nor U5853 (N_5853,N_5134,N_5210);
nand U5854 (N_5854,N_5224,N_5075);
nand U5855 (N_5855,N_5104,N_5288);
nor U5856 (N_5856,N_5219,N_5201);
and U5857 (N_5857,N_5175,N_5061);
or U5858 (N_5858,N_5246,N_5009);
and U5859 (N_5859,N_5279,N_5116);
and U5860 (N_5860,N_5498,N_5192);
and U5861 (N_5861,N_5428,N_5126);
or U5862 (N_5862,N_5389,N_5436);
nor U5863 (N_5863,N_5143,N_5013);
nand U5864 (N_5864,N_5320,N_5094);
nor U5865 (N_5865,N_5156,N_5382);
nand U5866 (N_5866,N_5162,N_5173);
and U5867 (N_5867,N_5067,N_5463);
or U5868 (N_5868,N_5368,N_5111);
or U5869 (N_5869,N_5215,N_5036);
nand U5870 (N_5870,N_5469,N_5147);
nand U5871 (N_5871,N_5167,N_5091);
xnor U5872 (N_5872,N_5004,N_5422);
or U5873 (N_5873,N_5246,N_5439);
or U5874 (N_5874,N_5178,N_5399);
nor U5875 (N_5875,N_5198,N_5367);
or U5876 (N_5876,N_5271,N_5419);
nor U5877 (N_5877,N_5265,N_5210);
nand U5878 (N_5878,N_5161,N_5357);
and U5879 (N_5879,N_5154,N_5198);
nor U5880 (N_5880,N_5456,N_5287);
nand U5881 (N_5881,N_5241,N_5442);
or U5882 (N_5882,N_5344,N_5246);
nand U5883 (N_5883,N_5124,N_5063);
nor U5884 (N_5884,N_5420,N_5010);
nand U5885 (N_5885,N_5210,N_5259);
nand U5886 (N_5886,N_5176,N_5383);
and U5887 (N_5887,N_5313,N_5156);
nand U5888 (N_5888,N_5347,N_5414);
xnor U5889 (N_5889,N_5036,N_5266);
or U5890 (N_5890,N_5241,N_5191);
xor U5891 (N_5891,N_5285,N_5098);
nor U5892 (N_5892,N_5410,N_5005);
or U5893 (N_5893,N_5090,N_5437);
nand U5894 (N_5894,N_5185,N_5425);
and U5895 (N_5895,N_5140,N_5278);
xor U5896 (N_5896,N_5385,N_5026);
nor U5897 (N_5897,N_5267,N_5021);
nor U5898 (N_5898,N_5302,N_5470);
nor U5899 (N_5899,N_5312,N_5298);
or U5900 (N_5900,N_5011,N_5287);
nor U5901 (N_5901,N_5322,N_5271);
xnor U5902 (N_5902,N_5405,N_5276);
nor U5903 (N_5903,N_5144,N_5430);
nand U5904 (N_5904,N_5465,N_5018);
nor U5905 (N_5905,N_5021,N_5259);
nand U5906 (N_5906,N_5116,N_5266);
or U5907 (N_5907,N_5114,N_5204);
nand U5908 (N_5908,N_5062,N_5184);
nor U5909 (N_5909,N_5265,N_5305);
nor U5910 (N_5910,N_5195,N_5145);
xor U5911 (N_5911,N_5172,N_5410);
xnor U5912 (N_5912,N_5087,N_5166);
nor U5913 (N_5913,N_5185,N_5261);
or U5914 (N_5914,N_5151,N_5221);
or U5915 (N_5915,N_5085,N_5146);
or U5916 (N_5916,N_5022,N_5472);
nor U5917 (N_5917,N_5100,N_5285);
and U5918 (N_5918,N_5010,N_5378);
and U5919 (N_5919,N_5048,N_5025);
nor U5920 (N_5920,N_5460,N_5001);
nand U5921 (N_5921,N_5464,N_5304);
xor U5922 (N_5922,N_5138,N_5159);
or U5923 (N_5923,N_5072,N_5173);
or U5924 (N_5924,N_5386,N_5240);
and U5925 (N_5925,N_5258,N_5239);
or U5926 (N_5926,N_5496,N_5482);
or U5927 (N_5927,N_5336,N_5191);
nand U5928 (N_5928,N_5037,N_5175);
nor U5929 (N_5929,N_5143,N_5235);
xor U5930 (N_5930,N_5010,N_5158);
xnor U5931 (N_5931,N_5365,N_5208);
or U5932 (N_5932,N_5395,N_5209);
or U5933 (N_5933,N_5017,N_5107);
or U5934 (N_5934,N_5242,N_5312);
nor U5935 (N_5935,N_5491,N_5261);
nand U5936 (N_5936,N_5346,N_5430);
nand U5937 (N_5937,N_5323,N_5118);
nor U5938 (N_5938,N_5100,N_5484);
and U5939 (N_5939,N_5156,N_5168);
or U5940 (N_5940,N_5445,N_5146);
nand U5941 (N_5941,N_5456,N_5006);
or U5942 (N_5942,N_5037,N_5058);
and U5943 (N_5943,N_5433,N_5403);
nor U5944 (N_5944,N_5130,N_5033);
nand U5945 (N_5945,N_5312,N_5156);
nor U5946 (N_5946,N_5105,N_5297);
nor U5947 (N_5947,N_5106,N_5484);
nor U5948 (N_5948,N_5460,N_5347);
nor U5949 (N_5949,N_5162,N_5081);
and U5950 (N_5950,N_5409,N_5286);
nand U5951 (N_5951,N_5126,N_5186);
nand U5952 (N_5952,N_5145,N_5255);
and U5953 (N_5953,N_5035,N_5107);
or U5954 (N_5954,N_5033,N_5061);
and U5955 (N_5955,N_5239,N_5040);
nor U5956 (N_5956,N_5477,N_5376);
nor U5957 (N_5957,N_5401,N_5125);
or U5958 (N_5958,N_5440,N_5413);
nor U5959 (N_5959,N_5445,N_5159);
or U5960 (N_5960,N_5436,N_5250);
and U5961 (N_5961,N_5048,N_5002);
nand U5962 (N_5962,N_5057,N_5405);
nand U5963 (N_5963,N_5403,N_5170);
or U5964 (N_5964,N_5499,N_5190);
or U5965 (N_5965,N_5155,N_5169);
nand U5966 (N_5966,N_5239,N_5337);
and U5967 (N_5967,N_5368,N_5009);
or U5968 (N_5968,N_5213,N_5493);
and U5969 (N_5969,N_5230,N_5168);
and U5970 (N_5970,N_5182,N_5347);
or U5971 (N_5971,N_5285,N_5106);
nand U5972 (N_5972,N_5469,N_5473);
nand U5973 (N_5973,N_5153,N_5195);
or U5974 (N_5974,N_5474,N_5156);
nand U5975 (N_5975,N_5051,N_5379);
and U5976 (N_5976,N_5498,N_5179);
nand U5977 (N_5977,N_5081,N_5143);
and U5978 (N_5978,N_5403,N_5297);
xor U5979 (N_5979,N_5108,N_5392);
and U5980 (N_5980,N_5044,N_5087);
or U5981 (N_5981,N_5364,N_5047);
or U5982 (N_5982,N_5398,N_5256);
or U5983 (N_5983,N_5390,N_5101);
xnor U5984 (N_5984,N_5140,N_5154);
or U5985 (N_5985,N_5408,N_5272);
xor U5986 (N_5986,N_5434,N_5069);
or U5987 (N_5987,N_5172,N_5059);
nor U5988 (N_5988,N_5496,N_5125);
nand U5989 (N_5989,N_5069,N_5460);
and U5990 (N_5990,N_5214,N_5399);
nand U5991 (N_5991,N_5262,N_5250);
nor U5992 (N_5992,N_5431,N_5290);
or U5993 (N_5993,N_5236,N_5220);
or U5994 (N_5994,N_5155,N_5086);
or U5995 (N_5995,N_5318,N_5015);
nor U5996 (N_5996,N_5262,N_5473);
or U5997 (N_5997,N_5081,N_5020);
and U5998 (N_5998,N_5406,N_5159);
and U5999 (N_5999,N_5122,N_5221);
nand U6000 (N_6000,N_5603,N_5660);
or U6001 (N_6001,N_5577,N_5697);
nor U6002 (N_6002,N_5525,N_5662);
and U6003 (N_6003,N_5788,N_5838);
nand U6004 (N_6004,N_5574,N_5916);
nor U6005 (N_6005,N_5804,N_5686);
xor U6006 (N_6006,N_5598,N_5817);
xor U6007 (N_6007,N_5856,N_5815);
or U6008 (N_6008,N_5573,N_5701);
or U6009 (N_6009,N_5555,N_5732);
nand U6010 (N_6010,N_5721,N_5944);
nand U6011 (N_6011,N_5772,N_5535);
nand U6012 (N_6012,N_5830,N_5570);
or U6013 (N_6013,N_5735,N_5629);
and U6014 (N_6014,N_5738,N_5962);
or U6015 (N_6015,N_5814,N_5726);
or U6016 (N_6016,N_5582,N_5786);
nand U6017 (N_6017,N_5544,N_5587);
nand U6018 (N_6018,N_5632,N_5554);
and U6019 (N_6019,N_5842,N_5831);
or U6020 (N_6020,N_5910,N_5876);
nor U6021 (N_6021,N_5595,N_5988);
nand U6022 (N_6022,N_5578,N_5779);
or U6023 (N_6023,N_5941,N_5930);
or U6024 (N_6024,N_5547,N_5989);
and U6025 (N_6025,N_5783,N_5503);
nor U6026 (N_6026,N_5625,N_5947);
nor U6027 (N_6027,N_5889,N_5537);
and U6028 (N_6028,N_5714,N_5911);
or U6029 (N_6029,N_5657,N_5664);
or U6030 (N_6030,N_5972,N_5608);
xor U6031 (N_6031,N_5542,N_5997);
or U6032 (N_6032,N_5763,N_5920);
and U6033 (N_6033,N_5516,N_5514);
and U6034 (N_6034,N_5954,N_5965);
nand U6035 (N_6035,N_5648,N_5995);
nor U6036 (N_6036,N_5899,N_5593);
nand U6037 (N_6037,N_5794,N_5541);
and U6038 (N_6038,N_5727,N_5986);
nand U6039 (N_6039,N_5543,N_5613);
nand U6040 (N_6040,N_5583,N_5680);
or U6041 (N_6041,N_5705,N_5650);
or U6042 (N_6042,N_5840,N_5870);
nor U6043 (N_6043,N_5746,N_5903);
xor U6044 (N_6044,N_5631,N_5971);
and U6045 (N_6045,N_5681,N_5756);
nor U6046 (N_6046,N_5599,N_5633);
nor U6047 (N_6047,N_5642,N_5862);
and U6048 (N_6048,N_5741,N_5579);
nand U6049 (N_6049,N_5908,N_5679);
or U6050 (N_6050,N_5517,N_5791);
and U6051 (N_6051,N_5829,N_5925);
and U6052 (N_6052,N_5687,N_5961);
nor U6053 (N_6053,N_5668,N_5959);
xor U6054 (N_6054,N_5528,N_5742);
or U6055 (N_6055,N_5766,N_5833);
nor U6056 (N_6056,N_5622,N_5875);
and U6057 (N_6057,N_5912,N_5855);
nand U6058 (N_6058,N_5940,N_5767);
nand U6059 (N_6059,N_5983,N_5931);
nand U6060 (N_6060,N_5684,N_5708);
xor U6061 (N_6061,N_5782,N_5780);
nand U6062 (N_6062,N_5607,N_5592);
nor U6063 (N_6063,N_5611,N_5576);
xnor U6064 (N_6064,N_5745,N_5935);
xor U6065 (N_6065,N_5702,N_5803);
xor U6066 (N_6066,N_5581,N_5623);
nor U6067 (N_6067,N_5801,N_5755);
nand U6068 (N_6068,N_5851,N_5627);
nor U6069 (N_6069,N_5649,N_5774);
nor U6070 (N_6070,N_5868,N_5723);
or U6071 (N_6071,N_5764,N_5644);
and U6072 (N_6072,N_5952,N_5559);
nand U6073 (N_6073,N_5634,N_5594);
or U6074 (N_6074,N_5653,N_5597);
nor U6075 (N_6075,N_5770,N_5784);
xnor U6076 (N_6076,N_5874,N_5575);
or U6077 (N_6077,N_5993,N_5926);
xor U6078 (N_6078,N_5663,N_5567);
nand U6079 (N_6079,N_5850,N_5877);
and U6080 (N_6080,N_5975,N_5685);
nand U6081 (N_6081,N_5809,N_5904);
and U6082 (N_6082,N_5945,N_5504);
and U6083 (N_6083,N_5812,N_5754);
and U6084 (N_6084,N_5566,N_5897);
or U6085 (N_6085,N_5557,N_5957);
or U6086 (N_6086,N_5729,N_5713);
or U6087 (N_6087,N_5939,N_5951);
xor U6088 (N_6088,N_5928,N_5602);
nand U6089 (N_6089,N_5606,N_5518);
nor U6090 (N_6090,N_5731,N_5658);
xor U6091 (N_6091,N_5506,N_5591);
nor U6092 (N_6092,N_5892,N_5641);
nor U6093 (N_6093,N_5869,N_5884);
nand U6094 (N_6094,N_5715,N_5548);
xor U6095 (N_6095,N_5698,N_5747);
nor U6096 (N_6096,N_5848,N_5672);
and U6097 (N_6097,N_5502,N_5725);
xor U6098 (N_6098,N_5828,N_5762);
or U6099 (N_6099,N_5707,N_5820);
and U6100 (N_6100,N_5530,N_5560);
and U6101 (N_6101,N_5861,N_5895);
nor U6102 (N_6102,N_5968,N_5849);
nor U6103 (N_6103,N_5666,N_5550);
and U6104 (N_6104,N_5656,N_5781);
and U6105 (N_6105,N_5757,N_5847);
xnor U6106 (N_6106,N_5963,N_5621);
or U6107 (N_6107,N_5775,N_5647);
nor U6108 (N_6108,N_5969,N_5758);
nand U6109 (N_6109,N_5932,N_5618);
nand U6110 (N_6110,N_5695,N_5860);
xor U6111 (N_6111,N_5998,N_5545);
nand U6112 (N_6112,N_5825,N_5584);
and U6113 (N_6113,N_5752,N_5948);
nor U6114 (N_6114,N_5790,N_5906);
nor U6115 (N_6115,N_5515,N_5845);
nand U6116 (N_6116,N_5964,N_5933);
nor U6117 (N_6117,N_5846,N_5551);
and U6118 (N_6118,N_5643,N_5915);
nor U6119 (N_6119,N_5572,N_5612);
nor U6120 (N_6120,N_5521,N_5802);
nor U6121 (N_6121,N_5859,N_5991);
nor U6122 (N_6122,N_5615,N_5938);
nand U6123 (N_6123,N_5696,N_5999);
nor U6124 (N_6124,N_5854,N_5953);
xor U6125 (N_6125,N_5785,N_5917);
nand U6126 (N_6126,N_5743,N_5558);
or U6127 (N_6127,N_5748,N_5699);
or U6128 (N_6128,N_5946,N_5778);
nand U6129 (N_6129,N_5671,N_5553);
nand U6130 (N_6130,N_5863,N_5994);
nor U6131 (N_6131,N_5977,N_5624);
nor U6132 (N_6132,N_5604,N_5609);
or U6133 (N_6133,N_5682,N_5841);
nand U6134 (N_6134,N_5898,N_5793);
nor U6135 (N_6135,N_5835,N_5956);
nor U6136 (N_6136,N_5880,N_5981);
and U6137 (N_6137,N_5588,N_5694);
or U6138 (N_6138,N_5651,N_5510);
and U6139 (N_6139,N_5990,N_5885);
nor U6140 (N_6140,N_5524,N_5822);
nand U6141 (N_6141,N_5980,N_5564);
nor U6142 (N_6142,N_5585,N_5960);
nor U6143 (N_6143,N_5508,N_5894);
nor U6144 (N_6144,N_5692,N_5569);
or U6145 (N_6145,N_5659,N_5601);
xnor U6146 (N_6146,N_5792,N_5500);
xor U6147 (N_6147,N_5922,N_5561);
or U6148 (N_6148,N_5873,N_5882);
or U6149 (N_6149,N_5966,N_5777);
and U6150 (N_6150,N_5832,N_5739);
xor U6151 (N_6151,N_5942,N_5638);
or U6152 (N_6152,N_5901,N_5676);
nand U6153 (N_6153,N_5529,N_5761);
nand U6154 (N_6154,N_5556,N_5798);
nand U6155 (N_6155,N_5526,N_5827);
or U6156 (N_6156,N_5534,N_5867);
and U6157 (N_6157,N_5652,N_5967);
xnor U6158 (N_6158,N_5523,N_5883);
and U6159 (N_6159,N_5736,N_5900);
or U6160 (N_6160,N_5734,N_5987);
nor U6161 (N_6161,N_5670,N_5807);
nand U6162 (N_6162,N_5985,N_5744);
or U6163 (N_6163,N_5620,N_5843);
and U6164 (N_6164,N_5984,N_5700);
nor U6165 (N_6165,N_5886,N_5816);
and U6166 (N_6166,N_5808,N_5619);
nor U6167 (N_6167,N_5586,N_5799);
nand U6168 (N_6168,N_5974,N_5691);
and U6169 (N_6169,N_5605,N_5858);
or U6170 (N_6170,N_5532,N_5538);
nor U6171 (N_6171,N_5639,N_5728);
or U6172 (N_6172,N_5918,N_5501);
nor U6173 (N_6173,N_5724,N_5852);
xnor U6174 (N_6174,N_5710,N_5864);
and U6175 (N_6175,N_5646,N_5513);
and U6176 (N_6176,N_5890,N_5665);
or U6177 (N_6177,N_5704,N_5776);
nand U6178 (N_6178,N_5865,N_5552);
nand U6179 (N_6179,N_5718,N_5914);
or U6180 (N_6180,N_5719,N_5887);
or U6181 (N_6181,N_5678,N_5511);
and U6182 (N_6182,N_5531,N_5590);
nor U6183 (N_6183,N_5789,N_5507);
xnor U6184 (N_6184,N_5949,N_5539);
or U6185 (N_6185,N_5805,N_5667);
and U6186 (N_6186,N_5982,N_5669);
nand U6187 (N_6187,N_5936,N_5893);
or U6188 (N_6188,N_5645,N_5536);
or U6189 (N_6189,N_5654,N_5636);
nand U6190 (N_6190,N_5675,N_5703);
or U6191 (N_6191,N_5673,N_5834);
nand U6192 (N_6192,N_5902,N_5637);
or U6193 (N_6193,N_5811,N_5768);
nand U6194 (N_6194,N_5796,N_5549);
xnor U6195 (N_6195,N_5913,N_5810);
nand U6196 (N_6196,N_5709,N_5616);
or U6197 (N_6197,N_5923,N_5787);
or U6198 (N_6198,N_5565,N_5821);
or U6199 (N_6199,N_5853,N_5600);
nor U6200 (N_6200,N_5765,N_5519);
nand U6201 (N_6201,N_5857,N_5753);
xnor U6202 (N_6202,N_5872,N_5527);
and U6203 (N_6203,N_5563,N_5836);
and U6204 (N_6204,N_5806,N_5771);
xor U6205 (N_6205,N_5509,N_5505);
or U6206 (N_6206,N_5750,N_5824);
xor U6207 (N_6207,N_5929,N_5773);
and U6208 (N_6208,N_5819,N_5866);
or U6209 (N_6209,N_5888,N_5655);
and U6210 (N_6210,N_5717,N_5562);
xnor U6211 (N_6211,N_5795,N_5958);
nand U6212 (N_6212,N_5891,N_5818);
and U6213 (N_6213,N_5759,N_5826);
and U6214 (N_6214,N_5711,N_5749);
xor U6215 (N_6215,N_5937,N_5823);
or U6216 (N_6216,N_5924,N_5979);
nor U6217 (N_6217,N_5706,N_5896);
nand U6218 (N_6218,N_5733,N_5540);
and U6219 (N_6219,N_5976,N_5740);
nand U6220 (N_6220,N_5722,N_5907);
xor U6221 (N_6221,N_5813,N_5878);
nor U6222 (N_6222,N_5690,N_5992);
nand U6223 (N_6223,N_5760,N_5512);
or U6224 (N_6224,N_5589,N_5533);
nor U6225 (N_6225,N_5769,N_5844);
and U6226 (N_6226,N_5596,N_5628);
nor U6227 (N_6227,N_5970,N_5716);
nor U6228 (N_6228,N_5905,N_5879);
nor U6229 (N_6229,N_5683,N_5919);
xnor U6230 (N_6230,N_5689,N_5800);
or U6231 (N_6231,N_5978,N_5568);
nand U6232 (N_6232,N_5614,N_5571);
and U6233 (N_6233,N_5546,N_5693);
and U6234 (N_6234,N_5943,N_5520);
nand U6235 (N_6235,N_5626,N_5837);
or U6236 (N_6236,N_5839,N_5934);
or U6237 (N_6237,N_5996,N_5751);
and U6238 (N_6238,N_5688,N_5677);
or U6239 (N_6239,N_5640,N_5580);
and U6240 (N_6240,N_5950,N_5674);
xor U6241 (N_6241,N_5720,N_5635);
or U6242 (N_6242,N_5712,N_5522);
and U6243 (N_6243,N_5661,N_5881);
xnor U6244 (N_6244,N_5797,N_5737);
or U6245 (N_6245,N_5610,N_5730);
or U6246 (N_6246,N_5921,N_5927);
xnor U6247 (N_6247,N_5630,N_5909);
xor U6248 (N_6248,N_5973,N_5617);
and U6249 (N_6249,N_5871,N_5955);
nor U6250 (N_6250,N_5734,N_5617);
nand U6251 (N_6251,N_5599,N_5780);
nand U6252 (N_6252,N_5812,N_5939);
nand U6253 (N_6253,N_5559,N_5657);
nand U6254 (N_6254,N_5900,N_5877);
or U6255 (N_6255,N_5528,N_5514);
and U6256 (N_6256,N_5963,N_5854);
and U6257 (N_6257,N_5828,N_5579);
xnor U6258 (N_6258,N_5557,N_5891);
xor U6259 (N_6259,N_5918,N_5763);
and U6260 (N_6260,N_5571,N_5930);
and U6261 (N_6261,N_5810,N_5847);
xnor U6262 (N_6262,N_5557,N_5639);
nor U6263 (N_6263,N_5812,N_5661);
or U6264 (N_6264,N_5549,N_5756);
nor U6265 (N_6265,N_5571,N_5638);
or U6266 (N_6266,N_5995,N_5590);
nor U6267 (N_6267,N_5600,N_5573);
nand U6268 (N_6268,N_5804,N_5852);
nor U6269 (N_6269,N_5871,N_5908);
or U6270 (N_6270,N_5531,N_5918);
nand U6271 (N_6271,N_5709,N_5532);
and U6272 (N_6272,N_5561,N_5870);
and U6273 (N_6273,N_5761,N_5909);
and U6274 (N_6274,N_5987,N_5615);
xnor U6275 (N_6275,N_5919,N_5747);
and U6276 (N_6276,N_5789,N_5796);
and U6277 (N_6277,N_5886,N_5577);
or U6278 (N_6278,N_5735,N_5532);
nand U6279 (N_6279,N_5687,N_5606);
nand U6280 (N_6280,N_5779,N_5995);
nand U6281 (N_6281,N_5768,N_5828);
and U6282 (N_6282,N_5986,N_5565);
and U6283 (N_6283,N_5964,N_5542);
xnor U6284 (N_6284,N_5935,N_5725);
nand U6285 (N_6285,N_5551,N_5824);
nor U6286 (N_6286,N_5694,N_5968);
nand U6287 (N_6287,N_5567,N_5998);
nor U6288 (N_6288,N_5541,N_5604);
or U6289 (N_6289,N_5843,N_5842);
and U6290 (N_6290,N_5509,N_5762);
xnor U6291 (N_6291,N_5785,N_5548);
nor U6292 (N_6292,N_5567,N_5596);
and U6293 (N_6293,N_5562,N_5525);
or U6294 (N_6294,N_5611,N_5772);
nand U6295 (N_6295,N_5545,N_5973);
nand U6296 (N_6296,N_5514,N_5753);
nand U6297 (N_6297,N_5638,N_5764);
or U6298 (N_6298,N_5650,N_5515);
nand U6299 (N_6299,N_5831,N_5908);
and U6300 (N_6300,N_5671,N_5842);
nor U6301 (N_6301,N_5847,N_5928);
nor U6302 (N_6302,N_5960,N_5777);
and U6303 (N_6303,N_5589,N_5643);
nand U6304 (N_6304,N_5864,N_5714);
nor U6305 (N_6305,N_5927,N_5778);
nor U6306 (N_6306,N_5672,N_5709);
nor U6307 (N_6307,N_5578,N_5731);
nor U6308 (N_6308,N_5592,N_5990);
nor U6309 (N_6309,N_5671,N_5697);
or U6310 (N_6310,N_5886,N_5920);
or U6311 (N_6311,N_5591,N_5894);
or U6312 (N_6312,N_5948,N_5676);
and U6313 (N_6313,N_5562,N_5500);
nor U6314 (N_6314,N_5948,N_5913);
nand U6315 (N_6315,N_5883,N_5923);
and U6316 (N_6316,N_5594,N_5923);
or U6317 (N_6317,N_5568,N_5770);
and U6318 (N_6318,N_5529,N_5922);
and U6319 (N_6319,N_5867,N_5994);
nand U6320 (N_6320,N_5902,N_5770);
xnor U6321 (N_6321,N_5642,N_5957);
or U6322 (N_6322,N_5563,N_5670);
and U6323 (N_6323,N_5782,N_5561);
nand U6324 (N_6324,N_5906,N_5910);
nor U6325 (N_6325,N_5984,N_5543);
xnor U6326 (N_6326,N_5736,N_5723);
and U6327 (N_6327,N_5944,N_5982);
and U6328 (N_6328,N_5521,N_5792);
and U6329 (N_6329,N_5733,N_5722);
nand U6330 (N_6330,N_5685,N_5848);
or U6331 (N_6331,N_5910,N_5505);
and U6332 (N_6332,N_5590,N_5568);
or U6333 (N_6333,N_5511,N_5856);
nor U6334 (N_6334,N_5832,N_5669);
nand U6335 (N_6335,N_5895,N_5734);
or U6336 (N_6336,N_5608,N_5891);
and U6337 (N_6337,N_5735,N_5585);
or U6338 (N_6338,N_5729,N_5945);
nor U6339 (N_6339,N_5890,N_5762);
and U6340 (N_6340,N_5605,N_5550);
nor U6341 (N_6341,N_5600,N_5899);
xor U6342 (N_6342,N_5955,N_5721);
and U6343 (N_6343,N_5522,N_5698);
and U6344 (N_6344,N_5893,N_5956);
or U6345 (N_6345,N_5845,N_5854);
nand U6346 (N_6346,N_5608,N_5823);
and U6347 (N_6347,N_5957,N_5906);
and U6348 (N_6348,N_5711,N_5894);
and U6349 (N_6349,N_5635,N_5772);
nand U6350 (N_6350,N_5784,N_5500);
xor U6351 (N_6351,N_5576,N_5997);
nor U6352 (N_6352,N_5944,N_5868);
or U6353 (N_6353,N_5816,N_5903);
or U6354 (N_6354,N_5957,N_5952);
or U6355 (N_6355,N_5511,N_5679);
and U6356 (N_6356,N_5906,N_5660);
xnor U6357 (N_6357,N_5598,N_5964);
xnor U6358 (N_6358,N_5761,N_5746);
or U6359 (N_6359,N_5629,N_5598);
or U6360 (N_6360,N_5616,N_5761);
or U6361 (N_6361,N_5970,N_5924);
nand U6362 (N_6362,N_5583,N_5677);
nand U6363 (N_6363,N_5829,N_5580);
nand U6364 (N_6364,N_5774,N_5839);
and U6365 (N_6365,N_5515,N_5571);
nand U6366 (N_6366,N_5930,N_5724);
nand U6367 (N_6367,N_5644,N_5555);
and U6368 (N_6368,N_5931,N_5833);
or U6369 (N_6369,N_5948,N_5784);
nor U6370 (N_6370,N_5602,N_5521);
nand U6371 (N_6371,N_5948,N_5746);
nand U6372 (N_6372,N_5759,N_5935);
and U6373 (N_6373,N_5647,N_5568);
nor U6374 (N_6374,N_5905,N_5941);
nor U6375 (N_6375,N_5715,N_5771);
nand U6376 (N_6376,N_5824,N_5533);
and U6377 (N_6377,N_5987,N_5949);
nor U6378 (N_6378,N_5824,N_5754);
or U6379 (N_6379,N_5877,N_5805);
and U6380 (N_6380,N_5572,N_5963);
and U6381 (N_6381,N_5887,N_5895);
or U6382 (N_6382,N_5667,N_5727);
nor U6383 (N_6383,N_5816,N_5950);
xor U6384 (N_6384,N_5741,N_5547);
and U6385 (N_6385,N_5897,N_5737);
or U6386 (N_6386,N_5923,N_5531);
or U6387 (N_6387,N_5818,N_5949);
nand U6388 (N_6388,N_5624,N_5752);
and U6389 (N_6389,N_5833,N_5810);
or U6390 (N_6390,N_5749,N_5978);
or U6391 (N_6391,N_5781,N_5734);
nand U6392 (N_6392,N_5740,N_5600);
and U6393 (N_6393,N_5884,N_5674);
nor U6394 (N_6394,N_5952,N_5595);
nor U6395 (N_6395,N_5563,N_5528);
and U6396 (N_6396,N_5608,N_5868);
xor U6397 (N_6397,N_5555,N_5973);
nor U6398 (N_6398,N_5821,N_5512);
nand U6399 (N_6399,N_5743,N_5553);
nor U6400 (N_6400,N_5657,N_5963);
nor U6401 (N_6401,N_5839,N_5677);
or U6402 (N_6402,N_5682,N_5517);
nand U6403 (N_6403,N_5567,N_5783);
nor U6404 (N_6404,N_5949,N_5773);
nor U6405 (N_6405,N_5875,N_5578);
nor U6406 (N_6406,N_5599,N_5888);
and U6407 (N_6407,N_5593,N_5690);
and U6408 (N_6408,N_5730,N_5773);
xnor U6409 (N_6409,N_5877,N_5544);
nand U6410 (N_6410,N_5624,N_5702);
or U6411 (N_6411,N_5752,N_5818);
or U6412 (N_6412,N_5787,N_5560);
or U6413 (N_6413,N_5577,N_5660);
or U6414 (N_6414,N_5945,N_5733);
nor U6415 (N_6415,N_5998,N_5556);
nor U6416 (N_6416,N_5734,N_5712);
and U6417 (N_6417,N_5890,N_5691);
and U6418 (N_6418,N_5687,N_5509);
or U6419 (N_6419,N_5634,N_5549);
or U6420 (N_6420,N_5778,N_5743);
nand U6421 (N_6421,N_5722,N_5536);
nand U6422 (N_6422,N_5527,N_5657);
and U6423 (N_6423,N_5594,N_5571);
xnor U6424 (N_6424,N_5546,N_5826);
xor U6425 (N_6425,N_5514,N_5986);
nand U6426 (N_6426,N_5545,N_5660);
nand U6427 (N_6427,N_5809,N_5520);
xnor U6428 (N_6428,N_5856,N_5644);
and U6429 (N_6429,N_5661,N_5715);
and U6430 (N_6430,N_5804,N_5619);
xnor U6431 (N_6431,N_5917,N_5790);
or U6432 (N_6432,N_5657,N_5682);
xnor U6433 (N_6433,N_5552,N_5964);
xnor U6434 (N_6434,N_5836,N_5940);
or U6435 (N_6435,N_5534,N_5503);
or U6436 (N_6436,N_5611,N_5599);
nor U6437 (N_6437,N_5765,N_5728);
and U6438 (N_6438,N_5572,N_5925);
nand U6439 (N_6439,N_5651,N_5722);
or U6440 (N_6440,N_5533,N_5925);
or U6441 (N_6441,N_5607,N_5734);
and U6442 (N_6442,N_5942,N_5903);
nor U6443 (N_6443,N_5507,N_5851);
nor U6444 (N_6444,N_5669,N_5957);
and U6445 (N_6445,N_5831,N_5529);
nand U6446 (N_6446,N_5914,N_5595);
or U6447 (N_6447,N_5935,N_5514);
nand U6448 (N_6448,N_5818,N_5857);
and U6449 (N_6449,N_5730,N_5625);
nand U6450 (N_6450,N_5599,N_5718);
nand U6451 (N_6451,N_5746,N_5536);
or U6452 (N_6452,N_5886,N_5602);
and U6453 (N_6453,N_5517,N_5796);
or U6454 (N_6454,N_5819,N_5911);
nand U6455 (N_6455,N_5545,N_5733);
or U6456 (N_6456,N_5938,N_5557);
or U6457 (N_6457,N_5892,N_5920);
or U6458 (N_6458,N_5840,N_5818);
nand U6459 (N_6459,N_5932,N_5600);
nor U6460 (N_6460,N_5803,N_5680);
nor U6461 (N_6461,N_5793,N_5822);
xor U6462 (N_6462,N_5602,N_5887);
nor U6463 (N_6463,N_5646,N_5594);
or U6464 (N_6464,N_5554,N_5685);
and U6465 (N_6465,N_5899,N_5517);
nor U6466 (N_6466,N_5857,N_5528);
nor U6467 (N_6467,N_5655,N_5995);
nor U6468 (N_6468,N_5759,N_5769);
nor U6469 (N_6469,N_5828,N_5522);
or U6470 (N_6470,N_5564,N_5924);
nand U6471 (N_6471,N_5954,N_5625);
and U6472 (N_6472,N_5744,N_5899);
nor U6473 (N_6473,N_5567,N_5939);
or U6474 (N_6474,N_5904,N_5565);
or U6475 (N_6475,N_5841,N_5835);
or U6476 (N_6476,N_5598,N_5967);
nand U6477 (N_6477,N_5566,N_5806);
and U6478 (N_6478,N_5628,N_5969);
and U6479 (N_6479,N_5583,N_5778);
or U6480 (N_6480,N_5833,N_5895);
nand U6481 (N_6481,N_5731,N_5839);
and U6482 (N_6482,N_5817,N_5815);
or U6483 (N_6483,N_5542,N_5557);
nand U6484 (N_6484,N_5880,N_5839);
nor U6485 (N_6485,N_5805,N_5838);
and U6486 (N_6486,N_5609,N_5880);
and U6487 (N_6487,N_5935,N_5851);
and U6488 (N_6488,N_5950,N_5608);
nand U6489 (N_6489,N_5652,N_5805);
and U6490 (N_6490,N_5681,N_5855);
or U6491 (N_6491,N_5574,N_5797);
or U6492 (N_6492,N_5957,N_5798);
nand U6493 (N_6493,N_5722,N_5883);
nor U6494 (N_6494,N_5730,N_5567);
and U6495 (N_6495,N_5782,N_5515);
xnor U6496 (N_6496,N_5575,N_5537);
and U6497 (N_6497,N_5768,N_5693);
nand U6498 (N_6498,N_5563,N_5900);
nor U6499 (N_6499,N_5837,N_5590);
nor U6500 (N_6500,N_6183,N_6418);
and U6501 (N_6501,N_6011,N_6133);
or U6502 (N_6502,N_6036,N_6128);
nand U6503 (N_6503,N_6097,N_6182);
or U6504 (N_6504,N_6433,N_6157);
or U6505 (N_6505,N_6226,N_6338);
and U6506 (N_6506,N_6363,N_6320);
and U6507 (N_6507,N_6148,N_6449);
xor U6508 (N_6508,N_6172,N_6118);
nor U6509 (N_6509,N_6101,N_6303);
xor U6510 (N_6510,N_6178,N_6120);
nand U6511 (N_6511,N_6307,N_6170);
and U6512 (N_6512,N_6187,N_6197);
nor U6513 (N_6513,N_6089,N_6115);
and U6514 (N_6514,N_6305,N_6437);
nor U6515 (N_6515,N_6162,N_6137);
nand U6516 (N_6516,N_6211,N_6257);
nand U6517 (N_6517,N_6213,N_6090);
and U6518 (N_6518,N_6264,N_6436);
and U6519 (N_6519,N_6049,N_6136);
xor U6520 (N_6520,N_6311,N_6399);
nand U6521 (N_6521,N_6330,N_6027);
and U6522 (N_6522,N_6283,N_6252);
xor U6523 (N_6523,N_6383,N_6122);
xnor U6524 (N_6524,N_6143,N_6452);
nand U6525 (N_6525,N_6254,N_6222);
or U6526 (N_6526,N_6343,N_6072);
and U6527 (N_6527,N_6054,N_6432);
and U6528 (N_6528,N_6391,N_6159);
xnor U6529 (N_6529,N_6411,N_6439);
xnor U6530 (N_6530,N_6160,N_6488);
and U6531 (N_6531,N_6123,N_6308);
and U6532 (N_6532,N_6209,N_6400);
nand U6533 (N_6533,N_6359,N_6313);
or U6534 (N_6534,N_6013,N_6316);
nand U6535 (N_6535,N_6425,N_6212);
nand U6536 (N_6536,N_6484,N_6131);
nand U6537 (N_6537,N_6253,N_6245);
or U6538 (N_6538,N_6181,N_6002);
nand U6539 (N_6539,N_6427,N_6053);
xnor U6540 (N_6540,N_6294,N_6219);
nand U6541 (N_6541,N_6358,N_6328);
or U6542 (N_6542,N_6149,N_6227);
and U6543 (N_6543,N_6239,N_6063);
nor U6544 (N_6544,N_6085,N_6349);
or U6545 (N_6545,N_6348,N_6016);
nand U6546 (N_6546,N_6247,N_6228);
and U6547 (N_6547,N_6326,N_6472);
and U6548 (N_6548,N_6024,N_6015);
nand U6549 (N_6549,N_6074,N_6420);
nor U6550 (N_6550,N_6234,N_6055);
or U6551 (N_6551,N_6144,N_6280);
or U6552 (N_6552,N_6084,N_6007);
or U6553 (N_6553,N_6435,N_6289);
nand U6554 (N_6554,N_6417,N_6052);
nand U6555 (N_6555,N_6481,N_6447);
or U6556 (N_6556,N_6493,N_6302);
nand U6557 (N_6557,N_6265,N_6448);
or U6558 (N_6558,N_6116,N_6486);
or U6559 (N_6559,N_6106,N_6379);
nor U6560 (N_6560,N_6281,N_6384);
nand U6561 (N_6561,N_6017,N_6478);
nand U6562 (N_6562,N_6499,N_6366);
nor U6563 (N_6563,N_6362,N_6155);
or U6564 (N_6564,N_6029,N_6340);
or U6565 (N_6565,N_6385,N_6457);
and U6566 (N_6566,N_6445,N_6467);
or U6567 (N_6567,N_6475,N_6415);
nor U6568 (N_6568,N_6071,N_6355);
nand U6569 (N_6569,N_6390,N_6235);
nand U6570 (N_6570,N_6494,N_6010);
nor U6571 (N_6571,N_6025,N_6271);
nor U6572 (N_6572,N_6476,N_6306);
or U6573 (N_6573,N_6060,N_6008);
nor U6574 (N_6574,N_6082,N_6310);
nand U6575 (N_6575,N_6040,N_6407);
and U6576 (N_6576,N_6471,N_6266);
nand U6577 (N_6577,N_6288,N_6180);
and U6578 (N_6578,N_6272,N_6332);
nand U6579 (N_6579,N_6466,N_6496);
or U6580 (N_6580,N_6165,N_6361);
xnor U6581 (N_6581,N_6026,N_6173);
nand U6582 (N_6582,N_6477,N_6167);
nand U6583 (N_6583,N_6102,N_6263);
and U6584 (N_6584,N_6278,N_6479);
and U6585 (N_6585,N_6387,N_6189);
nor U6586 (N_6586,N_6158,N_6062);
nand U6587 (N_6587,N_6166,N_6031);
nand U6588 (N_6588,N_6462,N_6012);
nand U6589 (N_6589,N_6103,N_6000);
and U6590 (N_6590,N_6039,N_6346);
nor U6591 (N_6591,N_6421,N_6438);
xnor U6592 (N_6592,N_6414,N_6230);
and U6593 (N_6593,N_6386,N_6270);
or U6594 (N_6594,N_6057,N_6075);
xor U6595 (N_6595,N_6339,N_6048);
nand U6596 (N_6596,N_6256,N_6091);
nand U6597 (N_6597,N_6498,N_6287);
nor U6598 (N_6598,N_6217,N_6333);
nor U6599 (N_6599,N_6004,N_6380);
and U6600 (N_6600,N_6369,N_6111);
or U6601 (N_6601,N_6161,N_6375);
or U6602 (N_6602,N_6087,N_6056);
or U6603 (N_6603,N_6315,N_6196);
or U6604 (N_6604,N_6020,N_6125);
or U6605 (N_6605,N_6274,N_6184);
xor U6606 (N_6606,N_6403,N_6037);
nand U6607 (N_6607,N_6487,N_6237);
or U6608 (N_6608,N_6463,N_6443);
or U6609 (N_6609,N_6273,N_6454);
and U6610 (N_6610,N_6188,N_6460);
nand U6611 (N_6611,N_6322,N_6080);
and U6612 (N_6612,N_6114,N_6474);
or U6613 (N_6613,N_6350,N_6014);
xor U6614 (N_6614,N_6318,N_6042);
nor U6615 (N_6615,N_6099,N_6216);
and U6616 (N_6616,N_6392,N_6461);
nand U6617 (N_6617,N_6317,N_6351);
and U6618 (N_6618,N_6088,N_6334);
nor U6619 (N_6619,N_6223,N_6325);
and U6620 (N_6620,N_6110,N_6431);
xor U6621 (N_6621,N_6490,N_6200);
or U6622 (N_6622,N_6360,N_6297);
and U6623 (N_6623,N_6497,N_6480);
nand U6624 (N_6624,N_6352,N_6067);
nand U6625 (N_6625,N_6127,N_6290);
xor U6626 (N_6626,N_6112,N_6098);
nand U6627 (N_6627,N_6168,N_6107);
or U6628 (N_6628,N_6413,N_6176);
nand U6629 (N_6629,N_6489,N_6347);
nand U6630 (N_6630,N_6203,N_6201);
or U6631 (N_6631,N_6299,N_6259);
or U6632 (N_6632,N_6204,N_6251);
nor U6633 (N_6633,N_6374,N_6022);
nand U6634 (N_6634,N_6105,N_6373);
and U6635 (N_6635,N_6073,N_6190);
and U6636 (N_6636,N_6255,N_6150);
nand U6637 (N_6637,N_6066,N_6376);
and U6638 (N_6638,N_6426,N_6336);
xnor U6639 (N_6639,N_6070,N_6059);
nor U6640 (N_6640,N_6241,N_6469);
nor U6641 (N_6641,N_6249,N_6248);
nand U6642 (N_6642,N_6006,N_6277);
or U6643 (N_6643,N_6221,N_6065);
nor U6644 (N_6644,N_6142,N_6381);
nor U6645 (N_6645,N_6129,N_6378);
or U6646 (N_6646,N_6191,N_6416);
xnor U6647 (N_6647,N_6304,N_6455);
nor U6648 (N_6648,N_6243,N_6398);
nand U6649 (N_6649,N_6081,N_6430);
xnor U6650 (N_6650,N_6092,N_6312);
or U6651 (N_6651,N_6260,N_6423);
and U6652 (N_6652,N_6045,N_6458);
and U6653 (N_6653,N_6193,N_6077);
or U6654 (N_6654,N_6079,N_6083);
nor U6655 (N_6655,N_6268,N_6152);
xor U6656 (N_6656,N_6335,N_6422);
nand U6657 (N_6657,N_6001,N_6371);
or U6658 (N_6658,N_6210,N_6061);
or U6659 (N_6659,N_6175,N_6282);
or U6660 (N_6660,N_6406,N_6396);
nand U6661 (N_6661,N_6286,N_6215);
nor U6662 (N_6662,N_6470,N_6370);
nand U6663 (N_6663,N_6284,N_6309);
or U6664 (N_6664,N_6229,N_6327);
nor U6665 (N_6665,N_6169,N_6300);
nand U6666 (N_6666,N_6291,N_6195);
nand U6667 (N_6667,N_6394,N_6242);
or U6668 (N_6668,N_6258,N_6434);
nand U6669 (N_6669,N_6344,N_6078);
and U6670 (N_6670,N_6473,N_6202);
nor U6671 (N_6671,N_6404,N_6064);
xnor U6672 (N_6672,N_6408,N_6468);
nand U6673 (N_6673,N_6035,N_6261);
nor U6674 (N_6674,N_6321,N_6113);
or U6675 (N_6675,N_6207,N_6285);
nor U6676 (N_6676,N_6319,N_6206);
nand U6677 (N_6677,N_6185,N_6232);
or U6678 (N_6678,N_6108,N_6147);
nor U6679 (N_6679,N_6096,N_6041);
nand U6680 (N_6680,N_6446,N_6492);
and U6681 (N_6681,N_6208,N_6341);
nor U6682 (N_6682,N_6104,N_6134);
nand U6683 (N_6683,N_6086,N_6068);
or U6684 (N_6684,N_6388,N_6246);
or U6685 (N_6685,N_6238,N_6402);
and U6686 (N_6686,N_6323,N_6028);
or U6687 (N_6687,N_6199,N_6395);
and U6688 (N_6688,N_6124,N_6353);
nand U6689 (N_6689,N_6132,N_6051);
or U6690 (N_6690,N_6009,N_6262);
or U6691 (N_6691,N_6043,N_6450);
and U6692 (N_6692,N_6186,N_6058);
nor U6693 (N_6693,N_6032,N_6044);
and U6694 (N_6694,N_6331,N_6046);
nor U6695 (N_6695,N_6214,N_6365);
nor U6696 (N_6696,N_6356,N_6459);
nor U6697 (N_6697,N_6109,N_6177);
nor U6698 (N_6698,N_6174,N_6192);
and U6699 (N_6699,N_6440,N_6126);
or U6700 (N_6700,N_6018,N_6050);
and U6701 (N_6701,N_6019,N_6441);
nand U6702 (N_6702,N_6357,N_6412);
and U6703 (N_6703,N_6179,N_6231);
nand U6704 (N_6704,N_6034,N_6377);
nor U6705 (N_6705,N_6093,N_6156);
nand U6706 (N_6706,N_6151,N_6389);
and U6707 (N_6707,N_6047,N_6003);
xnor U6708 (N_6708,N_6153,N_6135);
xor U6709 (N_6709,N_6139,N_6023);
nor U6710 (N_6710,N_6419,N_6205);
or U6711 (N_6711,N_6424,N_6224);
nand U6712 (N_6712,N_6405,N_6292);
nand U6713 (N_6713,N_6121,N_6117);
and U6714 (N_6714,N_6464,N_6364);
and U6715 (N_6715,N_6119,N_6410);
nor U6716 (N_6716,N_6094,N_6456);
and U6717 (N_6717,N_6295,N_6146);
or U6718 (N_6718,N_6337,N_6465);
nor U6719 (N_6719,N_6267,N_6030);
xor U6720 (N_6720,N_6276,N_6453);
or U6721 (N_6721,N_6485,N_6038);
or U6722 (N_6722,N_6095,N_6368);
nor U6723 (N_6723,N_6401,N_6138);
nand U6724 (N_6724,N_6451,N_6269);
or U6725 (N_6725,N_6495,N_6301);
xor U6726 (N_6726,N_6240,N_6069);
xor U6727 (N_6727,N_6296,N_6005);
nor U6728 (N_6728,N_6298,N_6428);
or U6729 (N_6729,N_6130,N_6367);
xnor U6730 (N_6730,N_6244,N_6382);
xor U6731 (N_6731,N_6314,N_6491);
nand U6732 (N_6732,N_6409,N_6393);
and U6733 (N_6733,N_6342,N_6397);
nor U6734 (N_6734,N_6236,N_6154);
and U6735 (N_6735,N_6076,N_6198);
nand U6736 (N_6736,N_6140,N_6250);
nand U6737 (N_6737,N_6163,N_6354);
nor U6738 (N_6738,N_6329,N_6141);
or U6739 (N_6739,N_6279,N_6225);
or U6740 (N_6740,N_6429,N_6345);
or U6741 (N_6741,N_6033,N_6233);
and U6742 (N_6742,N_6164,N_6275);
nand U6743 (N_6743,N_6483,N_6482);
or U6744 (N_6744,N_6218,N_6220);
or U6745 (N_6745,N_6444,N_6293);
or U6746 (N_6746,N_6194,N_6100);
and U6747 (N_6747,N_6324,N_6021);
nand U6748 (N_6748,N_6171,N_6442);
xnor U6749 (N_6749,N_6145,N_6372);
nor U6750 (N_6750,N_6334,N_6075);
or U6751 (N_6751,N_6157,N_6162);
nor U6752 (N_6752,N_6378,N_6280);
or U6753 (N_6753,N_6235,N_6340);
nand U6754 (N_6754,N_6339,N_6384);
nand U6755 (N_6755,N_6420,N_6235);
or U6756 (N_6756,N_6385,N_6296);
nor U6757 (N_6757,N_6216,N_6487);
nand U6758 (N_6758,N_6348,N_6035);
nor U6759 (N_6759,N_6184,N_6341);
nor U6760 (N_6760,N_6242,N_6009);
and U6761 (N_6761,N_6139,N_6286);
xnor U6762 (N_6762,N_6404,N_6173);
and U6763 (N_6763,N_6091,N_6259);
nand U6764 (N_6764,N_6134,N_6037);
nand U6765 (N_6765,N_6103,N_6321);
nor U6766 (N_6766,N_6203,N_6288);
nor U6767 (N_6767,N_6239,N_6153);
and U6768 (N_6768,N_6156,N_6443);
xnor U6769 (N_6769,N_6115,N_6053);
or U6770 (N_6770,N_6065,N_6381);
or U6771 (N_6771,N_6374,N_6355);
nor U6772 (N_6772,N_6091,N_6437);
nor U6773 (N_6773,N_6495,N_6442);
or U6774 (N_6774,N_6200,N_6173);
xnor U6775 (N_6775,N_6450,N_6000);
nor U6776 (N_6776,N_6045,N_6400);
nand U6777 (N_6777,N_6008,N_6479);
xnor U6778 (N_6778,N_6262,N_6345);
nor U6779 (N_6779,N_6243,N_6450);
or U6780 (N_6780,N_6418,N_6443);
and U6781 (N_6781,N_6455,N_6416);
xnor U6782 (N_6782,N_6225,N_6334);
or U6783 (N_6783,N_6179,N_6393);
and U6784 (N_6784,N_6159,N_6464);
or U6785 (N_6785,N_6104,N_6484);
and U6786 (N_6786,N_6289,N_6192);
or U6787 (N_6787,N_6441,N_6364);
nor U6788 (N_6788,N_6144,N_6374);
or U6789 (N_6789,N_6006,N_6478);
and U6790 (N_6790,N_6341,N_6312);
nor U6791 (N_6791,N_6287,N_6429);
nand U6792 (N_6792,N_6124,N_6469);
and U6793 (N_6793,N_6104,N_6127);
nor U6794 (N_6794,N_6246,N_6252);
nand U6795 (N_6795,N_6424,N_6100);
or U6796 (N_6796,N_6426,N_6055);
and U6797 (N_6797,N_6197,N_6464);
nor U6798 (N_6798,N_6415,N_6039);
and U6799 (N_6799,N_6009,N_6454);
or U6800 (N_6800,N_6313,N_6026);
nor U6801 (N_6801,N_6468,N_6313);
nand U6802 (N_6802,N_6480,N_6034);
and U6803 (N_6803,N_6106,N_6300);
nor U6804 (N_6804,N_6170,N_6385);
nand U6805 (N_6805,N_6046,N_6459);
nand U6806 (N_6806,N_6026,N_6107);
nand U6807 (N_6807,N_6318,N_6092);
nor U6808 (N_6808,N_6122,N_6465);
nor U6809 (N_6809,N_6092,N_6256);
nor U6810 (N_6810,N_6196,N_6402);
or U6811 (N_6811,N_6399,N_6165);
and U6812 (N_6812,N_6382,N_6024);
or U6813 (N_6813,N_6189,N_6375);
nor U6814 (N_6814,N_6320,N_6025);
xnor U6815 (N_6815,N_6251,N_6381);
nand U6816 (N_6816,N_6066,N_6347);
nor U6817 (N_6817,N_6137,N_6241);
nand U6818 (N_6818,N_6003,N_6065);
nand U6819 (N_6819,N_6068,N_6296);
nor U6820 (N_6820,N_6338,N_6486);
nor U6821 (N_6821,N_6269,N_6489);
and U6822 (N_6822,N_6489,N_6009);
nand U6823 (N_6823,N_6077,N_6032);
nand U6824 (N_6824,N_6366,N_6162);
xnor U6825 (N_6825,N_6483,N_6018);
xnor U6826 (N_6826,N_6475,N_6018);
or U6827 (N_6827,N_6480,N_6461);
xor U6828 (N_6828,N_6001,N_6096);
xnor U6829 (N_6829,N_6109,N_6154);
nor U6830 (N_6830,N_6372,N_6373);
nor U6831 (N_6831,N_6157,N_6075);
and U6832 (N_6832,N_6303,N_6263);
nor U6833 (N_6833,N_6464,N_6292);
or U6834 (N_6834,N_6225,N_6214);
or U6835 (N_6835,N_6373,N_6321);
or U6836 (N_6836,N_6072,N_6021);
nand U6837 (N_6837,N_6373,N_6468);
and U6838 (N_6838,N_6357,N_6259);
nand U6839 (N_6839,N_6169,N_6405);
or U6840 (N_6840,N_6226,N_6255);
or U6841 (N_6841,N_6096,N_6061);
nor U6842 (N_6842,N_6180,N_6119);
xor U6843 (N_6843,N_6436,N_6277);
nor U6844 (N_6844,N_6075,N_6200);
or U6845 (N_6845,N_6346,N_6298);
nor U6846 (N_6846,N_6240,N_6288);
nor U6847 (N_6847,N_6054,N_6419);
nand U6848 (N_6848,N_6322,N_6252);
nor U6849 (N_6849,N_6143,N_6117);
or U6850 (N_6850,N_6282,N_6207);
nor U6851 (N_6851,N_6445,N_6477);
nor U6852 (N_6852,N_6243,N_6152);
and U6853 (N_6853,N_6348,N_6383);
or U6854 (N_6854,N_6383,N_6004);
nor U6855 (N_6855,N_6052,N_6090);
and U6856 (N_6856,N_6241,N_6087);
and U6857 (N_6857,N_6169,N_6190);
and U6858 (N_6858,N_6299,N_6271);
nor U6859 (N_6859,N_6083,N_6011);
or U6860 (N_6860,N_6208,N_6467);
nor U6861 (N_6861,N_6471,N_6272);
or U6862 (N_6862,N_6454,N_6060);
or U6863 (N_6863,N_6118,N_6113);
or U6864 (N_6864,N_6443,N_6498);
nor U6865 (N_6865,N_6023,N_6212);
or U6866 (N_6866,N_6071,N_6408);
nand U6867 (N_6867,N_6045,N_6384);
xor U6868 (N_6868,N_6069,N_6477);
or U6869 (N_6869,N_6154,N_6090);
nand U6870 (N_6870,N_6077,N_6242);
nor U6871 (N_6871,N_6283,N_6456);
and U6872 (N_6872,N_6231,N_6472);
nor U6873 (N_6873,N_6473,N_6128);
nand U6874 (N_6874,N_6278,N_6089);
or U6875 (N_6875,N_6102,N_6245);
and U6876 (N_6876,N_6404,N_6422);
and U6877 (N_6877,N_6130,N_6485);
and U6878 (N_6878,N_6052,N_6179);
nor U6879 (N_6879,N_6000,N_6214);
nand U6880 (N_6880,N_6237,N_6414);
or U6881 (N_6881,N_6269,N_6223);
and U6882 (N_6882,N_6436,N_6421);
nor U6883 (N_6883,N_6369,N_6074);
or U6884 (N_6884,N_6240,N_6187);
and U6885 (N_6885,N_6469,N_6029);
and U6886 (N_6886,N_6231,N_6143);
or U6887 (N_6887,N_6367,N_6246);
or U6888 (N_6888,N_6216,N_6238);
or U6889 (N_6889,N_6202,N_6282);
and U6890 (N_6890,N_6218,N_6356);
nor U6891 (N_6891,N_6434,N_6225);
xor U6892 (N_6892,N_6203,N_6431);
xor U6893 (N_6893,N_6356,N_6483);
or U6894 (N_6894,N_6363,N_6389);
and U6895 (N_6895,N_6192,N_6488);
nand U6896 (N_6896,N_6191,N_6432);
and U6897 (N_6897,N_6195,N_6006);
and U6898 (N_6898,N_6125,N_6210);
and U6899 (N_6899,N_6451,N_6241);
nor U6900 (N_6900,N_6278,N_6242);
nand U6901 (N_6901,N_6294,N_6056);
and U6902 (N_6902,N_6121,N_6339);
nor U6903 (N_6903,N_6358,N_6113);
and U6904 (N_6904,N_6160,N_6448);
or U6905 (N_6905,N_6161,N_6322);
xnor U6906 (N_6906,N_6102,N_6170);
nand U6907 (N_6907,N_6174,N_6267);
or U6908 (N_6908,N_6420,N_6428);
nand U6909 (N_6909,N_6257,N_6041);
and U6910 (N_6910,N_6090,N_6393);
or U6911 (N_6911,N_6323,N_6008);
and U6912 (N_6912,N_6132,N_6477);
nand U6913 (N_6913,N_6091,N_6112);
nand U6914 (N_6914,N_6091,N_6153);
or U6915 (N_6915,N_6389,N_6399);
or U6916 (N_6916,N_6343,N_6400);
or U6917 (N_6917,N_6066,N_6116);
or U6918 (N_6918,N_6454,N_6310);
nand U6919 (N_6919,N_6062,N_6300);
nor U6920 (N_6920,N_6353,N_6400);
nand U6921 (N_6921,N_6493,N_6388);
and U6922 (N_6922,N_6477,N_6499);
or U6923 (N_6923,N_6115,N_6166);
and U6924 (N_6924,N_6238,N_6291);
nor U6925 (N_6925,N_6295,N_6250);
nand U6926 (N_6926,N_6420,N_6411);
nor U6927 (N_6927,N_6310,N_6408);
or U6928 (N_6928,N_6490,N_6271);
or U6929 (N_6929,N_6460,N_6338);
xor U6930 (N_6930,N_6368,N_6042);
nor U6931 (N_6931,N_6392,N_6112);
nand U6932 (N_6932,N_6492,N_6451);
and U6933 (N_6933,N_6259,N_6159);
nor U6934 (N_6934,N_6039,N_6063);
xnor U6935 (N_6935,N_6101,N_6119);
xor U6936 (N_6936,N_6228,N_6224);
nand U6937 (N_6937,N_6193,N_6417);
nand U6938 (N_6938,N_6476,N_6058);
nor U6939 (N_6939,N_6445,N_6278);
nor U6940 (N_6940,N_6137,N_6148);
and U6941 (N_6941,N_6199,N_6095);
xnor U6942 (N_6942,N_6463,N_6462);
and U6943 (N_6943,N_6032,N_6021);
or U6944 (N_6944,N_6336,N_6129);
or U6945 (N_6945,N_6190,N_6212);
nand U6946 (N_6946,N_6168,N_6065);
or U6947 (N_6947,N_6187,N_6253);
nor U6948 (N_6948,N_6382,N_6125);
nand U6949 (N_6949,N_6411,N_6106);
or U6950 (N_6950,N_6181,N_6021);
xnor U6951 (N_6951,N_6274,N_6287);
nor U6952 (N_6952,N_6267,N_6305);
nand U6953 (N_6953,N_6150,N_6483);
or U6954 (N_6954,N_6493,N_6489);
nor U6955 (N_6955,N_6185,N_6428);
and U6956 (N_6956,N_6465,N_6093);
or U6957 (N_6957,N_6185,N_6037);
xor U6958 (N_6958,N_6465,N_6424);
xor U6959 (N_6959,N_6242,N_6025);
nor U6960 (N_6960,N_6079,N_6097);
nor U6961 (N_6961,N_6245,N_6402);
xor U6962 (N_6962,N_6046,N_6265);
xor U6963 (N_6963,N_6115,N_6020);
nand U6964 (N_6964,N_6181,N_6466);
or U6965 (N_6965,N_6379,N_6265);
or U6966 (N_6966,N_6116,N_6314);
and U6967 (N_6967,N_6349,N_6090);
nor U6968 (N_6968,N_6160,N_6450);
or U6969 (N_6969,N_6452,N_6298);
xor U6970 (N_6970,N_6313,N_6462);
nand U6971 (N_6971,N_6318,N_6422);
xor U6972 (N_6972,N_6041,N_6226);
and U6973 (N_6973,N_6137,N_6009);
nor U6974 (N_6974,N_6034,N_6001);
nor U6975 (N_6975,N_6447,N_6397);
xnor U6976 (N_6976,N_6242,N_6020);
and U6977 (N_6977,N_6392,N_6062);
or U6978 (N_6978,N_6046,N_6272);
nand U6979 (N_6979,N_6121,N_6478);
nor U6980 (N_6980,N_6365,N_6390);
or U6981 (N_6981,N_6311,N_6046);
nor U6982 (N_6982,N_6131,N_6143);
nor U6983 (N_6983,N_6184,N_6369);
or U6984 (N_6984,N_6056,N_6096);
nand U6985 (N_6985,N_6126,N_6290);
nand U6986 (N_6986,N_6246,N_6414);
nand U6987 (N_6987,N_6344,N_6181);
nor U6988 (N_6988,N_6053,N_6232);
nand U6989 (N_6989,N_6371,N_6446);
nand U6990 (N_6990,N_6259,N_6397);
nand U6991 (N_6991,N_6123,N_6413);
nand U6992 (N_6992,N_6189,N_6326);
nor U6993 (N_6993,N_6107,N_6146);
and U6994 (N_6994,N_6026,N_6274);
nand U6995 (N_6995,N_6380,N_6427);
or U6996 (N_6996,N_6051,N_6100);
xor U6997 (N_6997,N_6193,N_6152);
nor U6998 (N_6998,N_6140,N_6370);
or U6999 (N_6999,N_6288,N_6124);
nor U7000 (N_7000,N_6947,N_6847);
or U7001 (N_7001,N_6906,N_6727);
xor U7002 (N_7002,N_6602,N_6842);
or U7003 (N_7003,N_6944,N_6566);
nand U7004 (N_7004,N_6525,N_6781);
nand U7005 (N_7005,N_6757,N_6739);
or U7006 (N_7006,N_6966,N_6932);
or U7007 (N_7007,N_6865,N_6586);
xnor U7008 (N_7008,N_6854,N_6989);
nand U7009 (N_7009,N_6667,N_6876);
or U7010 (N_7010,N_6861,N_6829);
xor U7011 (N_7011,N_6941,N_6538);
and U7012 (N_7012,N_6509,N_6970);
or U7013 (N_7013,N_6780,N_6617);
nor U7014 (N_7014,N_6974,N_6799);
nand U7015 (N_7015,N_6576,N_6807);
nor U7016 (N_7016,N_6852,N_6565);
nor U7017 (N_7017,N_6720,N_6637);
nor U7018 (N_7018,N_6598,N_6850);
nor U7019 (N_7019,N_6964,N_6649);
or U7020 (N_7020,N_6918,N_6791);
nand U7021 (N_7021,N_6759,N_6857);
nand U7022 (N_7022,N_6962,N_6561);
nor U7023 (N_7023,N_6661,N_6597);
nand U7024 (N_7024,N_6976,N_6978);
and U7025 (N_7025,N_6644,N_6969);
xor U7026 (N_7026,N_6764,N_6680);
nand U7027 (N_7027,N_6736,N_6646);
nand U7028 (N_7028,N_6758,N_6638);
or U7029 (N_7029,N_6864,N_6582);
nor U7030 (N_7030,N_6685,N_6578);
nor U7031 (N_7031,N_6772,N_6543);
nor U7032 (N_7032,N_6882,N_6802);
nand U7033 (N_7033,N_6684,N_6705);
nor U7034 (N_7034,N_6777,N_6907);
nand U7035 (N_7035,N_6963,N_6831);
and U7036 (N_7036,N_6501,N_6760);
nor U7037 (N_7037,N_6620,N_6670);
nand U7038 (N_7038,N_6821,N_6827);
xor U7039 (N_7039,N_6635,N_6722);
or U7040 (N_7040,N_6783,N_6689);
and U7041 (N_7041,N_6625,N_6936);
xor U7042 (N_7042,N_6693,N_6912);
or U7043 (N_7043,N_6539,N_6933);
nor U7044 (N_7044,N_6993,N_6623);
or U7045 (N_7045,N_6871,N_6826);
xnor U7046 (N_7046,N_6800,N_6778);
nand U7047 (N_7047,N_6817,N_6948);
nand U7048 (N_7048,N_6508,N_6731);
and U7049 (N_7049,N_6511,N_6603);
and U7050 (N_7050,N_6557,N_6591);
nand U7051 (N_7051,N_6558,N_6610);
nor U7052 (N_7052,N_6564,N_6665);
nor U7053 (N_7053,N_6837,N_6931);
xnor U7054 (N_7054,N_6686,N_6812);
nor U7055 (N_7055,N_6929,N_6880);
nor U7056 (N_7056,N_6896,N_6740);
nor U7057 (N_7057,N_6940,N_6529);
or U7058 (N_7058,N_6658,N_6587);
nand U7059 (N_7059,N_6921,N_6694);
xor U7060 (N_7060,N_6755,N_6518);
and U7061 (N_7061,N_6650,N_6814);
or U7062 (N_7062,N_6984,N_6920);
xor U7063 (N_7063,N_6887,N_6741);
or U7064 (N_7064,N_6553,N_6572);
and U7065 (N_7065,N_6700,N_6725);
nand U7066 (N_7066,N_6999,N_6728);
or U7067 (N_7067,N_6743,N_6830);
nor U7068 (N_7068,N_6593,N_6765);
xnor U7069 (N_7069,N_6951,N_6784);
nand U7070 (N_7070,N_6890,N_6698);
or U7071 (N_7071,N_6721,N_6884);
xnor U7072 (N_7072,N_6943,N_6959);
and U7073 (N_7073,N_6704,N_6879);
nand U7074 (N_7074,N_6626,N_6897);
nor U7075 (N_7075,N_6633,N_6872);
and U7076 (N_7076,N_6788,N_6604);
and U7077 (N_7077,N_6517,N_6647);
nand U7078 (N_7078,N_6971,N_6713);
xor U7079 (N_7079,N_6779,N_6859);
nor U7080 (N_7080,N_6608,N_6595);
nor U7081 (N_7081,N_6675,N_6874);
xnor U7082 (N_7082,N_6832,N_6592);
or U7083 (N_7083,N_6664,N_6526);
and U7084 (N_7084,N_6752,N_6523);
nor U7085 (N_7085,N_6917,N_6856);
nand U7086 (N_7086,N_6775,N_6886);
nand U7087 (N_7087,N_6891,N_6889);
nor U7088 (N_7088,N_6810,N_6998);
xor U7089 (N_7089,N_6581,N_6589);
or U7090 (N_7090,N_6733,N_6979);
nand U7091 (N_7091,N_6819,N_6546);
nor U7092 (N_7092,N_6697,N_6945);
and U7093 (N_7093,N_6988,N_6512);
nand U7094 (N_7094,N_6734,N_6688);
nor U7095 (N_7095,N_6678,N_6866);
and U7096 (N_7096,N_6513,N_6629);
or U7097 (N_7097,N_6754,N_6824);
nor U7098 (N_7098,N_6977,N_6957);
or U7099 (N_7099,N_6766,N_6939);
and U7100 (N_7100,N_6611,N_6510);
and U7101 (N_7101,N_6952,N_6596);
nand U7102 (N_7102,N_6796,N_6701);
nor U7103 (N_7103,N_6719,N_6858);
nand U7104 (N_7104,N_6574,N_6848);
and U7105 (N_7105,N_6937,N_6750);
or U7106 (N_7106,N_6537,N_6909);
xnor U7107 (N_7107,N_6738,N_6823);
and U7108 (N_7108,N_6811,N_6682);
nand U7109 (N_7109,N_6716,N_6655);
nand U7110 (N_7110,N_6562,N_6803);
and U7111 (N_7111,N_6973,N_6540);
xor U7112 (N_7112,N_6885,N_6900);
nor U7113 (N_7113,N_6541,N_6605);
or U7114 (N_7114,N_6691,N_6818);
nor U7115 (N_7115,N_6908,N_6601);
xor U7116 (N_7116,N_6676,N_6606);
nand U7117 (N_7117,N_6516,N_6875);
or U7118 (N_7118,N_6913,N_6514);
and U7119 (N_7119,N_6749,N_6753);
and U7120 (N_7120,N_6652,N_6965);
and U7121 (N_7121,N_6901,N_6816);
xnor U7122 (N_7122,N_6938,N_6982);
nand U7123 (N_7123,N_6881,N_6748);
nand U7124 (N_7124,N_6699,N_6506);
nand U7125 (N_7125,N_6668,N_6527);
and U7126 (N_7126,N_6924,N_6552);
nor U7127 (N_7127,N_6782,N_6946);
and U7128 (N_7128,N_6789,N_6899);
or U7129 (N_7129,N_6735,N_6573);
or U7130 (N_7130,N_6949,N_6806);
nor U7131 (N_7131,N_6869,N_6773);
nand U7132 (N_7132,N_6567,N_6961);
and U7133 (N_7133,N_6990,N_6922);
nand U7134 (N_7134,N_6996,N_6547);
nand U7135 (N_7135,N_6762,N_6744);
nor U7136 (N_7136,N_6895,N_6709);
xnor U7137 (N_7137,N_6795,N_6883);
and U7138 (N_7138,N_6645,N_6528);
nor U7139 (N_7139,N_6769,N_6981);
nand U7140 (N_7140,N_6532,N_6563);
nand U7141 (N_7141,N_6968,N_6870);
and U7142 (N_7142,N_6651,N_6588);
nor U7143 (N_7143,N_6535,N_6843);
and U7144 (N_7144,N_6956,N_6787);
nand U7145 (N_7145,N_6808,N_6571);
nand U7146 (N_7146,N_6640,N_6695);
and U7147 (N_7147,N_6726,N_6534);
and U7148 (N_7148,N_6706,N_6515);
and U7149 (N_7149,N_6844,N_6729);
or U7150 (N_7150,N_6530,N_6533);
nor U7151 (N_7151,N_6504,N_6923);
nor U7152 (N_7152,N_6860,N_6925);
or U7153 (N_7153,N_6991,N_6828);
nor U7154 (N_7154,N_6853,N_6621);
or U7155 (N_7155,N_6916,N_6544);
or U7156 (N_7156,N_6618,N_6556);
and U7157 (N_7157,N_6849,N_6672);
nand U7158 (N_7158,N_6607,N_6724);
and U7159 (N_7159,N_6833,N_6894);
nand U7160 (N_7160,N_6717,N_6584);
nand U7161 (N_7161,N_6730,N_6792);
nor U7162 (N_7162,N_6711,N_6793);
and U7163 (N_7163,N_6960,N_6980);
nand U7164 (N_7164,N_6674,N_6707);
nor U7165 (N_7165,N_6804,N_6953);
nand U7166 (N_7166,N_6545,N_6585);
and U7167 (N_7167,N_6522,N_6851);
nor U7168 (N_7168,N_6888,N_6656);
nand U7169 (N_7169,N_6955,N_6703);
and U7170 (N_7170,N_6659,N_6632);
nor U7171 (N_7171,N_6500,N_6642);
nand U7172 (N_7172,N_6867,N_6590);
nand U7173 (N_7173,N_6663,N_6519);
xnor U7174 (N_7174,N_6505,N_6737);
xnor U7175 (N_7175,N_6846,N_6628);
nand U7176 (N_7176,N_6942,N_6580);
or U7177 (N_7177,N_6502,N_6654);
nand U7178 (N_7178,N_6873,N_6614);
or U7179 (N_7179,N_6771,N_6863);
nand U7180 (N_7180,N_6554,N_6718);
nand U7181 (N_7181,N_6926,N_6776);
nand U7182 (N_7182,N_6579,N_6542);
and U7183 (N_7183,N_6641,N_6636);
nor U7184 (N_7184,N_6822,N_6615);
nor U7185 (N_7185,N_6631,N_6613);
or U7186 (N_7186,N_6967,N_6774);
and U7187 (N_7187,N_6935,N_6761);
xor U7188 (N_7188,N_6904,N_6845);
and U7189 (N_7189,N_6594,N_6815);
nor U7190 (N_7190,N_6855,N_6609);
nor U7191 (N_7191,N_6622,N_6751);
xor U7192 (N_7192,N_6627,N_6696);
nor U7193 (N_7193,N_6805,N_6555);
or U7194 (N_7194,N_6507,N_6732);
xor U7195 (N_7195,N_6930,N_6767);
nor U7196 (N_7196,N_6919,N_6985);
or U7197 (N_7197,N_6570,N_6928);
or U7198 (N_7198,N_6673,N_6549);
and U7199 (N_7199,N_6653,N_6836);
nand U7200 (N_7200,N_6994,N_6868);
or U7201 (N_7201,N_6524,N_6747);
nand U7202 (N_7202,N_6905,N_6708);
nand U7203 (N_7203,N_6839,N_6634);
or U7204 (N_7204,N_6893,N_6657);
and U7205 (N_7205,N_6715,N_6834);
and U7206 (N_7206,N_6862,N_6997);
or U7207 (N_7207,N_6575,N_6648);
and U7208 (N_7208,N_6841,N_6521);
nor U7209 (N_7209,N_6995,N_6798);
or U7210 (N_7210,N_6531,N_6548);
and U7211 (N_7211,N_6577,N_6568);
and U7212 (N_7212,N_6702,N_6742);
nor U7213 (N_7213,N_6550,N_6559);
xnor U7214 (N_7214,N_6786,N_6878);
nand U7215 (N_7215,N_6662,N_6583);
and U7216 (N_7216,N_6745,N_6972);
nor U7217 (N_7217,N_6820,N_6690);
nor U7218 (N_7218,N_6975,N_6987);
nor U7219 (N_7219,N_6958,N_6619);
or U7220 (N_7220,N_6677,N_6910);
or U7221 (N_7221,N_6746,N_6630);
or U7222 (N_7222,N_6838,N_6756);
and U7223 (N_7223,N_6660,N_6877);
xor U7224 (N_7224,N_6624,N_6914);
and U7225 (N_7225,N_6616,N_6520);
nor U7226 (N_7226,N_6892,N_6669);
and U7227 (N_7227,N_6794,N_6643);
nor U7228 (N_7228,N_6954,N_6712);
nand U7229 (N_7229,N_6911,N_6934);
xnor U7230 (N_7230,N_6679,N_6950);
or U7231 (N_7231,N_6770,N_6560);
or U7232 (N_7232,N_6903,N_6992);
xnor U7233 (N_7233,N_6986,N_6666);
or U7234 (N_7234,N_6790,N_6915);
or U7235 (N_7235,N_6671,N_6813);
or U7236 (N_7236,N_6569,N_6612);
and U7237 (N_7237,N_6768,N_6983);
nor U7238 (N_7238,N_6710,N_6825);
and U7239 (N_7239,N_6763,N_6902);
or U7240 (N_7240,N_6503,N_6692);
xor U7241 (N_7241,N_6723,N_6801);
or U7242 (N_7242,N_6599,N_6551);
nor U7243 (N_7243,N_6536,N_6840);
nor U7244 (N_7244,N_6714,N_6683);
nor U7245 (N_7245,N_6927,N_6687);
xnor U7246 (N_7246,N_6797,N_6809);
nand U7247 (N_7247,N_6898,N_6600);
nand U7248 (N_7248,N_6835,N_6681);
nor U7249 (N_7249,N_6785,N_6639);
and U7250 (N_7250,N_6772,N_6967);
nor U7251 (N_7251,N_6993,N_6744);
nor U7252 (N_7252,N_6689,N_6672);
and U7253 (N_7253,N_6515,N_6617);
xnor U7254 (N_7254,N_6847,N_6825);
nand U7255 (N_7255,N_6834,N_6838);
and U7256 (N_7256,N_6707,N_6522);
or U7257 (N_7257,N_6708,N_6520);
and U7258 (N_7258,N_6798,N_6687);
xnor U7259 (N_7259,N_6605,N_6715);
or U7260 (N_7260,N_6992,N_6680);
nor U7261 (N_7261,N_6732,N_6560);
nor U7262 (N_7262,N_6897,N_6630);
nor U7263 (N_7263,N_6890,N_6978);
nand U7264 (N_7264,N_6586,N_6667);
or U7265 (N_7265,N_6559,N_6718);
xnor U7266 (N_7266,N_6888,N_6690);
or U7267 (N_7267,N_6950,N_6656);
nand U7268 (N_7268,N_6989,N_6517);
nand U7269 (N_7269,N_6813,N_6854);
nand U7270 (N_7270,N_6967,N_6861);
nor U7271 (N_7271,N_6684,N_6652);
nand U7272 (N_7272,N_6674,N_6727);
nand U7273 (N_7273,N_6811,N_6892);
and U7274 (N_7274,N_6551,N_6724);
and U7275 (N_7275,N_6901,N_6712);
or U7276 (N_7276,N_6536,N_6950);
nand U7277 (N_7277,N_6776,N_6690);
nand U7278 (N_7278,N_6794,N_6896);
and U7279 (N_7279,N_6985,N_6802);
nand U7280 (N_7280,N_6672,N_6564);
nand U7281 (N_7281,N_6633,N_6592);
or U7282 (N_7282,N_6714,N_6839);
nand U7283 (N_7283,N_6893,N_6654);
nand U7284 (N_7284,N_6623,N_6575);
nor U7285 (N_7285,N_6892,N_6904);
nor U7286 (N_7286,N_6636,N_6629);
or U7287 (N_7287,N_6783,N_6736);
or U7288 (N_7288,N_6910,N_6619);
and U7289 (N_7289,N_6897,N_6808);
and U7290 (N_7290,N_6555,N_6852);
nand U7291 (N_7291,N_6617,N_6730);
nor U7292 (N_7292,N_6760,N_6910);
nand U7293 (N_7293,N_6506,N_6524);
or U7294 (N_7294,N_6642,N_6815);
and U7295 (N_7295,N_6604,N_6731);
or U7296 (N_7296,N_6563,N_6880);
or U7297 (N_7297,N_6986,N_6856);
or U7298 (N_7298,N_6780,N_6758);
nand U7299 (N_7299,N_6637,N_6745);
xnor U7300 (N_7300,N_6608,N_6789);
and U7301 (N_7301,N_6805,N_6925);
and U7302 (N_7302,N_6611,N_6601);
and U7303 (N_7303,N_6622,N_6616);
nand U7304 (N_7304,N_6843,N_6689);
nand U7305 (N_7305,N_6837,N_6597);
nand U7306 (N_7306,N_6514,N_6520);
and U7307 (N_7307,N_6955,N_6862);
nor U7308 (N_7308,N_6741,N_6721);
nor U7309 (N_7309,N_6682,N_6560);
or U7310 (N_7310,N_6553,N_6920);
xor U7311 (N_7311,N_6618,N_6792);
xor U7312 (N_7312,N_6940,N_6772);
nand U7313 (N_7313,N_6989,N_6608);
and U7314 (N_7314,N_6554,N_6556);
or U7315 (N_7315,N_6544,N_6782);
nand U7316 (N_7316,N_6841,N_6700);
nand U7317 (N_7317,N_6831,N_6979);
nand U7318 (N_7318,N_6553,N_6596);
or U7319 (N_7319,N_6665,N_6595);
and U7320 (N_7320,N_6921,N_6722);
or U7321 (N_7321,N_6865,N_6663);
nand U7322 (N_7322,N_6974,N_6590);
nand U7323 (N_7323,N_6719,N_6773);
nor U7324 (N_7324,N_6556,N_6920);
nand U7325 (N_7325,N_6600,N_6616);
nand U7326 (N_7326,N_6697,N_6850);
or U7327 (N_7327,N_6792,N_6766);
nand U7328 (N_7328,N_6684,N_6604);
and U7329 (N_7329,N_6877,N_6766);
nor U7330 (N_7330,N_6807,N_6929);
nand U7331 (N_7331,N_6910,N_6743);
nand U7332 (N_7332,N_6635,N_6761);
nor U7333 (N_7333,N_6917,N_6509);
nand U7334 (N_7334,N_6922,N_6999);
nand U7335 (N_7335,N_6801,N_6655);
or U7336 (N_7336,N_6871,N_6644);
and U7337 (N_7337,N_6582,N_6620);
nand U7338 (N_7338,N_6786,N_6664);
or U7339 (N_7339,N_6632,N_6906);
xnor U7340 (N_7340,N_6998,N_6555);
and U7341 (N_7341,N_6927,N_6982);
nand U7342 (N_7342,N_6550,N_6548);
nor U7343 (N_7343,N_6786,N_6954);
nor U7344 (N_7344,N_6542,N_6661);
and U7345 (N_7345,N_6771,N_6554);
or U7346 (N_7346,N_6629,N_6913);
and U7347 (N_7347,N_6936,N_6553);
nor U7348 (N_7348,N_6895,N_6780);
and U7349 (N_7349,N_6707,N_6696);
nand U7350 (N_7350,N_6706,N_6611);
nand U7351 (N_7351,N_6977,N_6775);
or U7352 (N_7352,N_6966,N_6820);
nand U7353 (N_7353,N_6934,N_6977);
or U7354 (N_7354,N_6560,N_6518);
nor U7355 (N_7355,N_6823,N_6548);
and U7356 (N_7356,N_6910,N_6508);
nand U7357 (N_7357,N_6738,N_6964);
nand U7358 (N_7358,N_6973,N_6924);
and U7359 (N_7359,N_6869,N_6517);
or U7360 (N_7360,N_6829,N_6526);
xnor U7361 (N_7361,N_6569,N_6756);
or U7362 (N_7362,N_6997,N_6609);
and U7363 (N_7363,N_6957,N_6941);
nand U7364 (N_7364,N_6670,N_6626);
nand U7365 (N_7365,N_6534,N_6550);
or U7366 (N_7366,N_6521,N_6910);
and U7367 (N_7367,N_6647,N_6725);
nand U7368 (N_7368,N_6948,N_6615);
and U7369 (N_7369,N_6879,N_6667);
nand U7370 (N_7370,N_6836,N_6808);
and U7371 (N_7371,N_6911,N_6807);
or U7372 (N_7372,N_6771,N_6860);
or U7373 (N_7373,N_6916,N_6612);
nor U7374 (N_7374,N_6642,N_6651);
nor U7375 (N_7375,N_6626,N_6660);
or U7376 (N_7376,N_6663,N_6817);
and U7377 (N_7377,N_6852,N_6965);
and U7378 (N_7378,N_6528,N_6517);
or U7379 (N_7379,N_6771,N_6687);
and U7380 (N_7380,N_6520,N_6959);
or U7381 (N_7381,N_6672,N_6709);
nand U7382 (N_7382,N_6725,N_6667);
nand U7383 (N_7383,N_6910,N_6993);
or U7384 (N_7384,N_6598,N_6715);
xnor U7385 (N_7385,N_6957,N_6927);
and U7386 (N_7386,N_6919,N_6840);
or U7387 (N_7387,N_6861,N_6961);
nand U7388 (N_7388,N_6850,N_6915);
nand U7389 (N_7389,N_6705,N_6829);
and U7390 (N_7390,N_6985,N_6953);
nor U7391 (N_7391,N_6575,N_6656);
nor U7392 (N_7392,N_6811,N_6861);
nand U7393 (N_7393,N_6919,N_6903);
and U7394 (N_7394,N_6962,N_6964);
nand U7395 (N_7395,N_6597,N_6764);
or U7396 (N_7396,N_6669,N_6752);
nand U7397 (N_7397,N_6515,N_6841);
nor U7398 (N_7398,N_6725,N_6833);
or U7399 (N_7399,N_6966,N_6653);
or U7400 (N_7400,N_6945,N_6666);
and U7401 (N_7401,N_6734,N_6941);
xor U7402 (N_7402,N_6930,N_6800);
nand U7403 (N_7403,N_6508,N_6673);
nor U7404 (N_7404,N_6924,N_6606);
nand U7405 (N_7405,N_6958,N_6859);
nand U7406 (N_7406,N_6646,N_6822);
nor U7407 (N_7407,N_6555,N_6888);
nand U7408 (N_7408,N_6589,N_6615);
or U7409 (N_7409,N_6964,N_6697);
nand U7410 (N_7410,N_6773,N_6861);
nand U7411 (N_7411,N_6808,N_6615);
nand U7412 (N_7412,N_6722,N_6523);
xor U7413 (N_7413,N_6847,N_6676);
nor U7414 (N_7414,N_6924,N_6510);
and U7415 (N_7415,N_6666,N_6888);
nor U7416 (N_7416,N_6700,N_6569);
or U7417 (N_7417,N_6801,N_6677);
xor U7418 (N_7418,N_6667,N_6803);
or U7419 (N_7419,N_6772,N_6616);
nor U7420 (N_7420,N_6924,N_6513);
xor U7421 (N_7421,N_6806,N_6561);
xor U7422 (N_7422,N_6520,N_6962);
nand U7423 (N_7423,N_6515,N_6994);
nor U7424 (N_7424,N_6991,N_6607);
nand U7425 (N_7425,N_6606,N_6516);
nor U7426 (N_7426,N_6531,N_6966);
nor U7427 (N_7427,N_6565,N_6521);
nand U7428 (N_7428,N_6894,N_6754);
and U7429 (N_7429,N_6651,N_6806);
nor U7430 (N_7430,N_6827,N_6510);
nor U7431 (N_7431,N_6863,N_6948);
and U7432 (N_7432,N_6514,N_6693);
or U7433 (N_7433,N_6935,N_6892);
xor U7434 (N_7434,N_6972,N_6978);
and U7435 (N_7435,N_6666,N_6507);
and U7436 (N_7436,N_6695,N_6883);
and U7437 (N_7437,N_6689,N_6892);
nand U7438 (N_7438,N_6990,N_6898);
or U7439 (N_7439,N_6570,N_6944);
and U7440 (N_7440,N_6639,N_6850);
nand U7441 (N_7441,N_6589,N_6971);
or U7442 (N_7442,N_6624,N_6575);
and U7443 (N_7443,N_6806,N_6772);
and U7444 (N_7444,N_6530,N_6895);
and U7445 (N_7445,N_6509,N_6740);
nor U7446 (N_7446,N_6842,N_6959);
xnor U7447 (N_7447,N_6662,N_6707);
nor U7448 (N_7448,N_6880,N_6584);
or U7449 (N_7449,N_6940,N_6810);
and U7450 (N_7450,N_6597,N_6610);
and U7451 (N_7451,N_6589,N_6551);
nand U7452 (N_7452,N_6829,N_6666);
or U7453 (N_7453,N_6817,N_6767);
nand U7454 (N_7454,N_6966,N_6660);
nand U7455 (N_7455,N_6553,N_6852);
nand U7456 (N_7456,N_6626,N_6989);
or U7457 (N_7457,N_6650,N_6640);
nor U7458 (N_7458,N_6976,N_6531);
xor U7459 (N_7459,N_6687,N_6611);
and U7460 (N_7460,N_6519,N_6922);
or U7461 (N_7461,N_6695,N_6843);
or U7462 (N_7462,N_6669,N_6821);
nor U7463 (N_7463,N_6788,N_6597);
nand U7464 (N_7464,N_6904,N_6940);
nor U7465 (N_7465,N_6520,N_6785);
nor U7466 (N_7466,N_6520,N_6948);
nor U7467 (N_7467,N_6957,N_6654);
or U7468 (N_7468,N_6643,N_6630);
nor U7469 (N_7469,N_6538,N_6935);
or U7470 (N_7470,N_6628,N_6660);
or U7471 (N_7471,N_6656,N_6823);
or U7472 (N_7472,N_6530,N_6827);
nor U7473 (N_7473,N_6904,N_6928);
nand U7474 (N_7474,N_6872,N_6866);
nand U7475 (N_7475,N_6914,N_6863);
nand U7476 (N_7476,N_6642,N_6925);
and U7477 (N_7477,N_6732,N_6914);
or U7478 (N_7478,N_6948,N_6844);
nand U7479 (N_7479,N_6990,N_6889);
nor U7480 (N_7480,N_6931,N_6923);
nand U7481 (N_7481,N_6523,N_6622);
or U7482 (N_7482,N_6616,N_6501);
nand U7483 (N_7483,N_6977,N_6701);
nor U7484 (N_7484,N_6702,N_6733);
or U7485 (N_7485,N_6721,N_6822);
and U7486 (N_7486,N_6722,N_6950);
and U7487 (N_7487,N_6976,N_6699);
and U7488 (N_7488,N_6967,N_6541);
xor U7489 (N_7489,N_6939,N_6827);
and U7490 (N_7490,N_6549,N_6954);
nand U7491 (N_7491,N_6779,N_6577);
or U7492 (N_7492,N_6546,N_6608);
nor U7493 (N_7493,N_6686,N_6991);
nand U7494 (N_7494,N_6887,N_6779);
or U7495 (N_7495,N_6761,N_6590);
or U7496 (N_7496,N_6602,N_6914);
nor U7497 (N_7497,N_6675,N_6955);
nor U7498 (N_7498,N_6853,N_6789);
xnor U7499 (N_7499,N_6995,N_6850);
and U7500 (N_7500,N_7121,N_7286);
nor U7501 (N_7501,N_7188,N_7157);
nand U7502 (N_7502,N_7104,N_7031);
nor U7503 (N_7503,N_7006,N_7111);
nand U7504 (N_7504,N_7219,N_7255);
nand U7505 (N_7505,N_7159,N_7493);
nor U7506 (N_7506,N_7181,N_7138);
nor U7507 (N_7507,N_7236,N_7002);
or U7508 (N_7508,N_7357,N_7471);
nor U7509 (N_7509,N_7217,N_7205);
nand U7510 (N_7510,N_7402,N_7048);
nor U7511 (N_7511,N_7132,N_7320);
or U7512 (N_7512,N_7478,N_7208);
or U7513 (N_7513,N_7338,N_7095);
xnor U7514 (N_7514,N_7023,N_7393);
xor U7515 (N_7515,N_7271,N_7253);
or U7516 (N_7516,N_7124,N_7430);
nor U7517 (N_7517,N_7274,N_7462);
nor U7518 (N_7518,N_7213,N_7116);
and U7519 (N_7519,N_7364,N_7339);
xnor U7520 (N_7520,N_7428,N_7375);
and U7521 (N_7521,N_7042,N_7449);
nor U7522 (N_7522,N_7491,N_7414);
nand U7523 (N_7523,N_7486,N_7399);
nand U7524 (N_7524,N_7390,N_7293);
nand U7525 (N_7525,N_7052,N_7066);
and U7526 (N_7526,N_7228,N_7030);
nand U7527 (N_7527,N_7018,N_7056);
and U7528 (N_7528,N_7404,N_7251);
xnor U7529 (N_7529,N_7101,N_7283);
nand U7530 (N_7530,N_7290,N_7352);
nand U7531 (N_7531,N_7200,N_7322);
and U7532 (N_7532,N_7452,N_7191);
nand U7533 (N_7533,N_7425,N_7222);
or U7534 (N_7534,N_7093,N_7445);
nor U7535 (N_7535,N_7440,N_7315);
and U7536 (N_7536,N_7300,N_7298);
or U7537 (N_7537,N_7496,N_7137);
or U7538 (N_7538,N_7483,N_7131);
nor U7539 (N_7539,N_7108,N_7078);
or U7540 (N_7540,N_7372,N_7426);
nor U7541 (N_7541,N_7017,N_7475);
nand U7542 (N_7542,N_7340,N_7058);
and U7543 (N_7543,N_7015,N_7317);
or U7544 (N_7544,N_7127,N_7079);
or U7545 (N_7545,N_7266,N_7203);
nand U7546 (N_7546,N_7480,N_7029);
nor U7547 (N_7547,N_7419,N_7256);
nand U7548 (N_7548,N_7162,N_7140);
or U7549 (N_7549,N_7073,N_7223);
and U7550 (N_7550,N_7163,N_7099);
and U7551 (N_7551,N_7190,N_7450);
nor U7552 (N_7552,N_7201,N_7392);
nor U7553 (N_7553,N_7246,N_7244);
or U7554 (N_7554,N_7453,N_7403);
nor U7555 (N_7555,N_7362,N_7242);
or U7556 (N_7556,N_7479,N_7154);
or U7557 (N_7557,N_7356,N_7458);
nand U7558 (N_7558,N_7128,N_7368);
nor U7559 (N_7559,N_7265,N_7463);
nor U7560 (N_7560,N_7423,N_7313);
and U7561 (N_7561,N_7305,N_7335);
and U7562 (N_7562,N_7468,N_7429);
or U7563 (N_7563,N_7182,N_7459);
nor U7564 (N_7564,N_7366,N_7355);
nor U7565 (N_7565,N_7091,N_7443);
and U7566 (N_7566,N_7169,N_7295);
or U7567 (N_7567,N_7331,N_7025);
or U7568 (N_7568,N_7276,N_7278);
or U7569 (N_7569,N_7050,N_7319);
nand U7570 (N_7570,N_7466,N_7420);
nor U7571 (N_7571,N_7062,N_7408);
nand U7572 (N_7572,N_7460,N_7032);
or U7573 (N_7573,N_7397,N_7324);
or U7574 (N_7574,N_7406,N_7282);
or U7575 (N_7575,N_7467,N_7326);
nand U7576 (N_7576,N_7381,N_7387);
or U7577 (N_7577,N_7446,N_7036);
and U7578 (N_7578,N_7046,N_7084);
nand U7579 (N_7579,N_7220,N_7080);
or U7580 (N_7580,N_7092,N_7343);
or U7581 (N_7581,N_7325,N_7369);
and U7582 (N_7582,N_7260,N_7151);
xnor U7583 (N_7583,N_7008,N_7411);
nand U7584 (N_7584,N_7301,N_7198);
xor U7585 (N_7585,N_7035,N_7060);
nor U7586 (N_7586,N_7410,N_7027);
nor U7587 (N_7587,N_7299,N_7363);
nand U7588 (N_7588,N_7371,N_7413);
nor U7589 (N_7589,N_7102,N_7409);
and U7590 (N_7590,N_7441,N_7344);
or U7591 (N_7591,N_7185,N_7373);
and U7592 (N_7592,N_7226,N_7388);
or U7593 (N_7593,N_7168,N_7361);
and U7594 (N_7594,N_7125,N_7037);
nor U7595 (N_7595,N_7360,N_7234);
nand U7596 (N_7596,N_7156,N_7418);
or U7597 (N_7597,N_7396,N_7476);
nand U7598 (N_7598,N_7119,N_7342);
nor U7599 (N_7599,N_7051,N_7438);
and U7600 (N_7600,N_7382,N_7248);
or U7601 (N_7601,N_7264,N_7164);
and U7602 (N_7602,N_7341,N_7176);
nor U7603 (N_7603,N_7321,N_7126);
and U7604 (N_7604,N_7421,N_7351);
nand U7605 (N_7605,N_7327,N_7153);
nand U7606 (N_7606,N_7063,N_7416);
nor U7607 (N_7607,N_7498,N_7395);
nor U7608 (N_7608,N_7249,N_7318);
and U7609 (N_7609,N_7113,N_7141);
nand U7610 (N_7610,N_7149,N_7383);
or U7611 (N_7611,N_7225,N_7405);
nor U7612 (N_7612,N_7165,N_7235);
or U7613 (N_7613,N_7385,N_7435);
xor U7614 (N_7614,N_7207,N_7232);
and U7615 (N_7615,N_7391,N_7177);
and U7616 (N_7616,N_7328,N_7152);
nand U7617 (N_7617,N_7484,N_7014);
xnor U7618 (N_7618,N_7133,N_7199);
nor U7619 (N_7619,N_7145,N_7353);
or U7620 (N_7620,N_7069,N_7401);
xor U7621 (N_7621,N_7304,N_7136);
or U7622 (N_7622,N_7214,N_7332);
nor U7623 (N_7623,N_7323,N_7001);
or U7624 (N_7624,N_7227,N_7433);
and U7625 (N_7625,N_7389,N_7270);
or U7626 (N_7626,N_7284,N_7489);
or U7627 (N_7627,N_7469,N_7081);
and U7628 (N_7628,N_7100,N_7252);
nand U7629 (N_7629,N_7071,N_7034);
nand U7630 (N_7630,N_7494,N_7146);
or U7631 (N_7631,N_7041,N_7129);
and U7632 (N_7632,N_7365,N_7135);
nor U7633 (N_7633,N_7285,N_7412);
xnor U7634 (N_7634,N_7134,N_7336);
nand U7635 (N_7635,N_7189,N_7019);
or U7636 (N_7636,N_7005,N_7011);
nor U7637 (N_7637,N_7296,N_7292);
or U7638 (N_7638,N_7142,N_7055);
nand U7639 (N_7639,N_7487,N_7122);
and U7640 (N_7640,N_7022,N_7485);
and U7641 (N_7641,N_7139,N_7044);
xor U7642 (N_7642,N_7279,N_7209);
and U7643 (N_7643,N_7334,N_7302);
nor U7644 (N_7644,N_7345,N_7273);
nor U7645 (N_7645,N_7247,N_7170);
or U7646 (N_7646,N_7243,N_7378);
nand U7647 (N_7647,N_7086,N_7202);
nand U7648 (N_7648,N_7431,N_7075);
nor U7649 (N_7649,N_7269,N_7085);
nor U7650 (N_7650,N_7303,N_7377);
nand U7651 (N_7651,N_7310,N_7258);
nand U7652 (N_7652,N_7474,N_7171);
or U7653 (N_7653,N_7239,N_7180);
and U7654 (N_7654,N_7061,N_7077);
xor U7655 (N_7655,N_7206,N_7497);
nor U7656 (N_7656,N_7442,N_7280);
nor U7657 (N_7657,N_7106,N_7120);
nor U7658 (N_7658,N_7007,N_7059);
or U7659 (N_7659,N_7354,N_7367);
xor U7660 (N_7660,N_7407,N_7291);
or U7661 (N_7661,N_7178,N_7472);
nand U7662 (N_7662,N_7499,N_7175);
nand U7663 (N_7663,N_7043,N_7233);
nor U7664 (N_7664,N_7263,N_7094);
or U7665 (N_7665,N_7337,N_7481);
and U7666 (N_7666,N_7039,N_7314);
nor U7667 (N_7667,N_7147,N_7144);
and U7668 (N_7668,N_7238,N_7155);
nor U7669 (N_7669,N_7434,N_7229);
nor U7670 (N_7670,N_7461,N_7312);
and U7671 (N_7671,N_7384,N_7187);
or U7672 (N_7672,N_7281,N_7398);
or U7673 (N_7673,N_7422,N_7103);
nor U7674 (N_7674,N_7415,N_7306);
xor U7675 (N_7675,N_7148,N_7473);
or U7676 (N_7676,N_7218,N_7432);
nor U7677 (N_7677,N_7150,N_7192);
or U7678 (N_7678,N_7427,N_7386);
and U7679 (N_7679,N_7010,N_7183);
nor U7680 (N_7680,N_7329,N_7020);
and U7681 (N_7681,N_7262,N_7068);
nand U7682 (N_7682,N_7359,N_7216);
nand U7683 (N_7683,N_7289,N_7437);
nor U7684 (N_7684,N_7455,N_7003);
or U7685 (N_7685,N_7464,N_7424);
and U7686 (N_7686,N_7047,N_7013);
or U7687 (N_7687,N_7240,N_7370);
or U7688 (N_7688,N_7307,N_7117);
or U7689 (N_7689,N_7114,N_7297);
and U7690 (N_7690,N_7211,N_7186);
nor U7691 (N_7691,N_7349,N_7105);
xnor U7692 (N_7692,N_7465,N_7087);
nor U7693 (N_7693,N_7064,N_7118);
nand U7694 (N_7694,N_7330,N_7143);
or U7695 (N_7695,N_7495,N_7110);
xor U7696 (N_7696,N_7254,N_7000);
nand U7697 (N_7697,N_7374,N_7259);
and U7698 (N_7698,N_7076,N_7012);
nand U7699 (N_7699,N_7350,N_7089);
nand U7700 (N_7700,N_7161,N_7309);
or U7701 (N_7701,N_7123,N_7166);
or U7702 (N_7702,N_7028,N_7346);
nand U7703 (N_7703,N_7492,N_7275);
nor U7704 (N_7704,N_7221,N_7488);
nor U7705 (N_7705,N_7130,N_7268);
nor U7706 (N_7706,N_7380,N_7054);
nor U7707 (N_7707,N_7287,N_7237);
nor U7708 (N_7708,N_7158,N_7444);
and U7709 (N_7709,N_7311,N_7067);
and U7710 (N_7710,N_7033,N_7272);
and U7711 (N_7711,N_7195,N_7204);
nor U7712 (N_7712,N_7482,N_7447);
nor U7713 (N_7713,N_7115,N_7004);
and U7714 (N_7714,N_7016,N_7172);
xor U7715 (N_7715,N_7184,N_7107);
nor U7716 (N_7716,N_7477,N_7070);
and U7717 (N_7717,N_7112,N_7090);
nor U7718 (N_7718,N_7316,N_7417);
nand U7719 (N_7719,N_7379,N_7457);
nand U7720 (N_7720,N_7294,N_7210);
nand U7721 (N_7721,N_7333,N_7057);
and U7722 (N_7722,N_7261,N_7038);
nor U7723 (N_7723,N_7096,N_7308);
or U7724 (N_7724,N_7045,N_7267);
nor U7725 (N_7725,N_7215,N_7024);
or U7726 (N_7726,N_7490,N_7009);
or U7727 (N_7727,N_7348,N_7470);
or U7728 (N_7728,N_7196,N_7212);
and U7729 (N_7729,N_7098,N_7241);
xnor U7730 (N_7730,N_7082,N_7358);
nand U7731 (N_7731,N_7021,N_7167);
nand U7732 (N_7732,N_7088,N_7193);
or U7733 (N_7733,N_7097,N_7230);
or U7734 (N_7734,N_7454,N_7347);
nor U7735 (N_7735,N_7074,N_7288);
or U7736 (N_7736,N_7456,N_7053);
or U7737 (N_7737,N_7376,N_7194);
or U7738 (N_7738,N_7065,N_7394);
nand U7739 (N_7739,N_7245,N_7109);
or U7740 (N_7740,N_7174,N_7179);
or U7741 (N_7741,N_7224,N_7026);
and U7742 (N_7742,N_7160,N_7083);
and U7743 (N_7743,N_7049,N_7451);
nor U7744 (N_7744,N_7439,N_7277);
and U7745 (N_7745,N_7250,N_7040);
nor U7746 (N_7746,N_7257,N_7400);
xnor U7747 (N_7747,N_7436,N_7173);
nor U7748 (N_7748,N_7448,N_7231);
or U7749 (N_7749,N_7072,N_7197);
nor U7750 (N_7750,N_7034,N_7243);
or U7751 (N_7751,N_7134,N_7402);
nor U7752 (N_7752,N_7213,N_7143);
nor U7753 (N_7753,N_7079,N_7097);
nand U7754 (N_7754,N_7449,N_7092);
nand U7755 (N_7755,N_7245,N_7296);
xnor U7756 (N_7756,N_7488,N_7451);
or U7757 (N_7757,N_7333,N_7365);
and U7758 (N_7758,N_7317,N_7452);
or U7759 (N_7759,N_7204,N_7160);
nand U7760 (N_7760,N_7460,N_7428);
nor U7761 (N_7761,N_7321,N_7264);
xor U7762 (N_7762,N_7488,N_7436);
and U7763 (N_7763,N_7208,N_7248);
and U7764 (N_7764,N_7469,N_7023);
and U7765 (N_7765,N_7213,N_7367);
or U7766 (N_7766,N_7488,N_7490);
nand U7767 (N_7767,N_7261,N_7470);
xor U7768 (N_7768,N_7353,N_7497);
xnor U7769 (N_7769,N_7240,N_7475);
nand U7770 (N_7770,N_7379,N_7030);
xor U7771 (N_7771,N_7474,N_7466);
and U7772 (N_7772,N_7468,N_7345);
nor U7773 (N_7773,N_7149,N_7419);
and U7774 (N_7774,N_7290,N_7004);
or U7775 (N_7775,N_7088,N_7271);
and U7776 (N_7776,N_7257,N_7439);
nand U7777 (N_7777,N_7122,N_7085);
and U7778 (N_7778,N_7248,N_7213);
or U7779 (N_7779,N_7145,N_7305);
xor U7780 (N_7780,N_7232,N_7179);
nand U7781 (N_7781,N_7073,N_7142);
and U7782 (N_7782,N_7494,N_7099);
nand U7783 (N_7783,N_7478,N_7393);
xnor U7784 (N_7784,N_7107,N_7484);
nor U7785 (N_7785,N_7089,N_7463);
nor U7786 (N_7786,N_7115,N_7353);
or U7787 (N_7787,N_7108,N_7439);
nor U7788 (N_7788,N_7307,N_7224);
and U7789 (N_7789,N_7043,N_7405);
or U7790 (N_7790,N_7437,N_7134);
xnor U7791 (N_7791,N_7389,N_7252);
nand U7792 (N_7792,N_7299,N_7002);
or U7793 (N_7793,N_7358,N_7135);
or U7794 (N_7794,N_7414,N_7033);
nor U7795 (N_7795,N_7140,N_7079);
or U7796 (N_7796,N_7259,N_7257);
nor U7797 (N_7797,N_7097,N_7396);
nand U7798 (N_7798,N_7478,N_7085);
xnor U7799 (N_7799,N_7097,N_7414);
and U7800 (N_7800,N_7065,N_7142);
or U7801 (N_7801,N_7357,N_7389);
and U7802 (N_7802,N_7035,N_7420);
and U7803 (N_7803,N_7306,N_7397);
nor U7804 (N_7804,N_7134,N_7330);
nand U7805 (N_7805,N_7056,N_7307);
nand U7806 (N_7806,N_7173,N_7479);
xnor U7807 (N_7807,N_7066,N_7391);
and U7808 (N_7808,N_7138,N_7041);
and U7809 (N_7809,N_7217,N_7315);
nand U7810 (N_7810,N_7082,N_7417);
nand U7811 (N_7811,N_7021,N_7456);
or U7812 (N_7812,N_7029,N_7274);
and U7813 (N_7813,N_7439,N_7220);
nand U7814 (N_7814,N_7143,N_7184);
and U7815 (N_7815,N_7072,N_7487);
nand U7816 (N_7816,N_7003,N_7085);
and U7817 (N_7817,N_7428,N_7247);
nor U7818 (N_7818,N_7121,N_7077);
nor U7819 (N_7819,N_7328,N_7223);
nor U7820 (N_7820,N_7480,N_7475);
or U7821 (N_7821,N_7252,N_7276);
nor U7822 (N_7822,N_7230,N_7294);
or U7823 (N_7823,N_7355,N_7338);
nand U7824 (N_7824,N_7181,N_7498);
and U7825 (N_7825,N_7309,N_7292);
nor U7826 (N_7826,N_7149,N_7045);
nand U7827 (N_7827,N_7032,N_7112);
nor U7828 (N_7828,N_7156,N_7427);
and U7829 (N_7829,N_7305,N_7249);
nand U7830 (N_7830,N_7265,N_7184);
nor U7831 (N_7831,N_7021,N_7365);
and U7832 (N_7832,N_7365,N_7023);
and U7833 (N_7833,N_7011,N_7424);
and U7834 (N_7834,N_7289,N_7065);
nand U7835 (N_7835,N_7132,N_7017);
nor U7836 (N_7836,N_7389,N_7088);
xor U7837 (N_7837,N_7153,N_7080);
nor U7838 (N_7838,N_7189,N_7229);
nand U7839 (N_7839,N_7396,N_7110);
or U7840 (N_7840,N_7439,N_7003);
or U7841 (N_7841,N_7282,N_7403);
nand U7842 (N_7842,N_7375,N_7095);
and U7843 (N_7843,N_7483,N_7253);
and U7844 (N_7844,N_7448,N_7118);
nand U7845 (N_7845,N_7465,N_7002);
nor U7846 (N_7846,N_7426,N_7216);
nand U7847 (N_7847,N_7145,N_7198);
xnor U7848 (N_7848,N_7009,N_7007);
or U7849 (N_7849,N_7108,N_7397);
xnor U7850 (N_7850,N_7062,N_7419);
nor U7851 (N_7851,N_7470,N_7472);
nand U7852 (N_7852,N_7206,N_7180);
nand U7853 (N_7853,N_7442,N_7092);
nor U7854 (N_7854,N_7485,N_7009);
nor U7855 (N_7855,N_7441,N_7397);
and U7856 (N_7856,N_7040,N_7134);
or U7857 (N_7857,N_7149,N_7173);
xor U7858 (N_7858,N_7176,N_7042);
nand U7859 (N_7859,N_7039,N_7485);
nand U7860 (N_7860,N_7309,N_7412);
nor U7861 (N_7861,N_7472,N_7247);
nand U7862 (N_7862,N_7335,N_7477);
nor U7863 (N_7863,N_7240,N_7472);
and U7864 (N_7864,N_7345,N_7389);
or U7865 (N_7865,N_7296,N_7077);
nand U7866 (N_7866,N_7235,N_7098);
or U7867 (N_7867,N_7031,N_7120);
or U7868 (N_7868,N_7229,N_7235);
and U7869 (N_7869,N_7040,N_7387);
nand U7870 (N_7870,N_7136,N_7282);
nor U7871 (N_7871,N_7201,N_7285);
nor U7872 (N_7872,N_7265,N_7113);
or U7873 (N_7873,N_7131,N_7352);
nor U7874 (N_7874,N_7317,N_7228);
or U7875 (N_7875,N_7205,N_7219);
or U7876 (N_7876,N_7381,N_7096);
and U7877 (N_7877,N_7277,N_7290);
nand U7878 (N_7878,N_7108,N_7232);
nor U7879 (N_7879,N_7359,N_7483);
nor U7880 (N_7880,N_7187,N_7191);
nor U7881 (N_7881,N_7425,N_7201);
or U7882 (N_7882,N_7316,N_7110);
or U7883 (N_7883,N_7428,N_7317);
xnor U7884 (N_7884,N_7392,N_7098);
nand U7885 (N_7885,N_7248,N_7230);
and U7886 (N_7886,N_7180,N_7087);
nor U7887 (N_7887,N_7361,N_7414);
and U7888 (N_7888,N_7471,N_7203);
nor U7889 (N_7889,N_7180,N_7103);
and U7890 (N_7890,N_7290,N_7282);
nor U7891 (N_7891,N_7004,N_7118);
xor U7892 (N_7892,N_7040,N_7106);
and U7893 (N_7893,N_7331,N_7493);
and U7894 (N_7894,N_7355,N_7367);
nand U7895 (N_7895,N_7320,N_7019);
nand U7896 (N_7896,N_7089,N_7162);
and U7897 (N_7897,N_7285,N_7349);
nor U7898 (N_7898,N_7405,N_7206);
nand U7899 (N_7899,N_7220,N_7236);
nand U7900 (N_7900,N_7298,N_7257);
nor U7901 (N_7901,N_7155,N_7286);
xnor U7902 (N_7902,N_7103,N_7371);
nand U7903 (N_7903,N_7222,N_7484);
xor U7904 (N_7904,N_7381,N_7211);
xor U7905 (N_7905,N_7264,N_7480);
or U7906 (N_7906,N_7101,N_7225);
or U7907 (N_7907,N_7060,N_7392);
xor U7908 (N_7908,N_7384,N_7206);
nor U7909 (N_7909,N_7067,N_7090);
nor U7910 (N_7910,N_7299,N_7355);
or U7911 (N_7911,N_7156,N_7446);
and U7912 (N_7912,N_7286,N_7461);
nand U7913 (N_7913,N_7382,N_7197);
and U7914 (N_7914,N_7478,N_7316);
xnor U7915 (N_7915,N_7391,N_7004);
or U7916 (N_7916,N_7412,N_7019);
and U7917 (N_7917,N_7264,N_7348);
nor U7918 (N_7918,N_7349,N_7358);
nand U7919 (N_7919,N_7041,N_7018);
nor U7920 (N_7920,N_7204,N_7485);
or U7921 (N_7921,N_7100,N_7367);
nand U7922 (N_7922,N_7058,N_7247);
nand U7923 (N_7923,N_7289,N_7390);
nand U7924 (N_7924,N_7264,N_7313);
nor U7925 (N_7925,N_7348,N_7334);
nor U7926 (N_7926,N_7033,N_7099);
and U7927 (N_7927,N_7432,N_7043);
nor U7928 (N_7928,N_7439,N_7475);
or U7929 (N_7929,N_7031,N_7231);
nor U7930 (N_7930,N_7394,N_7308);
nor U7931 (N_7931,N_7228,N_7234);
or U7932 (N_7932,N_7048,N_7346);
and U7933 (N_7933,N_7065,N_7022);
and U7934 (N_7934,N_7310,N_7465);
nor U7935 (N_7935,N_7260,N_7140);
nand U7936 (N_7936,N_7456,N_7328);
nor U7937 (N_7937,N_7429,N_7061);
nand U7938 (N_7938,N_7287,N_7109);
nor U7939 (N_7939,N_7086,N_7204);
and U7940 (N_7940,N_7118,N_7057);
nor U7941 (N_7941,N_7384,N_7420);
and U7942 (N_7942,N_7332,N_7122);
nand U7943 (N_7943,N_7465,N_7071);
nor U7944 (N_7944,N_7168,N_7287);
nor U7945 (N_7945,N_7459,N_7140);
nor U7946 (N_7946,N_7261,N_7112);
nor U7947 (N_7947,N_7270,N_7328);
or U7948 (N_7948,N_7357,N_7452);
xnor U7949 (N_7949,N_7429,N_7268);
nand U7950 (N_7950,N_7439,N_7495);
nand U7951 (N_7951,N_7317,N_7352);
nand U7952 (N_7952,N_7050,N_7210);
nand U7953 (N_7953,N_7325,N_7073);
or U7954 (N_7954,N_7465,N_7297);
xor U7955 (N_7955,N_7437,N_7266);
and U7956 (N_7956,N_7409,N_7273);
nand U7957 (N_7957,N_7081,N_7400);
and U7958 (N_7958,N_7279,N_7122);
nand U7959 (N_7959,N_7266,N_7229);
or U7960 (N_7960,N_7048,N_7184);
nand U7961 (N_7961,N_7467,N_7454);
nor U7962 (N_7962,N_7366,N_7276);
xnor U7963 (N_7963,N_7314,N_7422);
or U7964 (N_7964,N_7454,N_7073);
or U7965 (N_7965,N_7377,N_7422);
or U7966 (N_7966,N_7226,N_7204);
nand U7967 (N_7967,N_7243,N_7310);
and U7968 (N_7968,N_7079,N_7442);
nand U7969 (N_7969,N_7091,N_7458);
nor U7970 (N_7970,N_7014,N_7024);
nand U7971 (N_7971,N_7012,N_7348);
and U7972 (N_7972,N_7215,N_7133);
nand U7973 (N_7973,N_7472,N_7035);
xnor U7974 (N_7974,N_7095,N_7101);
nor U7975 (N_7975,N_7488,N_7119);
xor U7976 (N_7976,N_7273,N_7489);
and U7977 (N_7977,N_7345,N_7410);
or U7978 (N_7978,N_7402,N_7131);
or U7979 (N_7979,N_7301,N_7261);
and U7980 (N_7980,N_7486,N_7078);
and U7981 (N_7981,N_7006,N_7407);
nand U7982 (N_7982,N_7267,N_7113);
or U7983 (N_7983,N_7421,N_7429);
nor U7984 (N_7984,N_7324,N_7482);
or U7985 (N_7985,N_7330,N_7358);
or U7986 (N_7986,N_7034,N_7185);
xnor U7987 (N_7987,N_7365,N_7234);
xnor U7988 (N_7988,N_7329,N_7017);
nand U7989 (N_7989,N_7420,N_7045);
or U7990 (N_7990,N_7301,N_7022);
nor U7991 (N_7991,N_7164,N_7456);
xor U7992 (N_7992,N_7043,N_7497);
nor U7993 (N_7993,N_7479,N_7247);
and U7994 (N_7994,N_7027,N_7335);
or U7995 (N_7995,N_7340,N_7400);
and U7996 (N_7996,N_7003,N_7069);
and U7997 (N_7997,N_7160,N_7494);
or U7998 (N_7998,N_7272,N_7382);
and U7999 (N_7999,N_7053,N_7303);
nand U8000 (N_8000,N_7583,N_7932);
nor U8001 (N_8001,N_7980,N_7720);
nor U8002 (N_8002,N_7505,N_7902);
nand U8003 (N_8003,N_7629,N_7983);
or U8004 (N_8004,N_7817,N_7652);
and U8005 (N_8005,N_7595,N_7634);
nor U8006 (N_8006,N_7805,N_7935);
and U8007 (N_8007,N_7685,N_7815);
xor U8008 (N_8008,N_7764,N_7984);
nor U8009 (N_8009,N_7526,N_7787);
and U8010 (N_8010,N_7694,N_7898);
nand U8011 (N_8011,N_7551,N_7524);
nor U8012 (N_8012,N_7995,N_7577);
nor U8013 (N_8013,N_7920,N_7534);
or U8014 (N_8014,N_7573,N_7814);
and U8015 (N_8015,N_7574,N_7942);
nand U8016 (N_8016,N_7769,N_7934);
nand U8017 (N_8017,N_7851,N_7861);
nor U8018 (N_8018,N_7758,N_7530);
nand U8019 (N_8019,N_7722,N_7788);
or U8020 (N_8020,N_7614,N_7841);
or U8021 (N_8021,N_7716,N_7775);
nand U8022 (N_8022,N_7850,N_7559);
nand U8023 (N_8023,N_7963,N_7907);
and U8024 (N_8024,N_7818,N_7992);
or U8025 (N_8025,N_7514,N_7681);
nand U8026 (N_8026,N_7831,N_7964);
nor U8027 (N_8027,N_7522,N_7721);
nor U8028 (N_8028,N_7585,N_7656);
or U8029 (N_8029,N_7823,N_7800);
nand U8030 (N_8030,N_7771,N_7881);
nor U8031 (N_8031,N_7858,N_7579);
xor U8032 (N_8032,N_7550,N_7874);
and U8033 (N_8033,N_7885,N_7693);
xor U8034 (N_8034,N_7873,N_7682);
nand U8035 (N_8035,N_7708,N_7811);
and U8036 (N_8036,N_7589,N_7677);
or U8037 (N_8037,N_7588,N_7752);
nor U8038 (N_8038,N_7894,N_7649);
or U8039 (N_8039,N_7944,N_7864);
and U8040 (N_8040,N_7508,N_7690);
nor U8041 (N_8041,N_7616,N_7725);
nor U8042 (N_8042,N_7926,N_7836);
nand U8043 (N_8043,N_7840,N_7949);
or U8044 (N_8044,N_7987,N_7698);
or U8045 (N_8045,N_7795,N_7611);
nor U8046 (N_8046,N_7901,N_7896);
and U8047 (N_8047,N_7950,N_7511);
and U8048 (N_8048,N_7968,N_7679);
nand U8049 (N_8049,N_7986,N_7596);
nand U8050 (N_8050,N_7643,N_7994);
xnor U8051 (N_8051,N_7518,N_7878);
xor U8052 (N_8052,N_7726,N_7739);
or U8053 (N_8053,N_7691,N_7832);
nand U8054 (N_8054,N_7804,N_7504);
nor U8055 (N_8055,N_7566,N_7843);
nor U8056 (N_8056,N_7922,N_7662);
nand U8057 (N_8057,N_7871,N_7625);
nor U8058 (N_8058,N_7711,N_7848);
or U8059 (N_8059,N_7765,N_7704);
nand U8060 (N_8060,N_7658,N_7970);
or U8061 (N_8061,N_7978,N_7819);
and U8062 (N_8062,N_7971,N_7664);
xnor U8063 (N_8063,N_7906,N_7736);
nand U8064 (N_8064,N_7703,N_7740);
nor U8065 (N_8065,N_7510,N_7745);
nor U8066 (N_8066,N_7558,N_7809);
nand U8067 (N_8067,N_7731,N_7977);
or U8068 (N_8068,N_7692,N_7940);
nor U8069 (N_8069,N_7607,N_7673);
nor U8070 (N_8070,N_7501,N_7748);
and U8071 (N_8071,N_7939,N_7960);
nor U8072 (N_8072,N_7821,N_7737);
and U8073 (N_8073,N_7762,N_7751);
and U8074 (N_8074,N_7816,N_7536);
nor U8075 (N_8075,N_7976,N_7930);
nand U8076 (N_8076,N_7908,N_7569);
xnor U8077 (N_8077,N_7863,N_7601);
xnor U8078 (N_8078,N_7602,N_7715);
or U8079 (N_8079,N_7648,N_7827);
nand U8080 (N_8080,N_7888,N_7810);
and U8081 (N_8081,N_7791,N_7660);
or U8082 (N_8082,N_7626,N_7644);
and U8083 (N_8083,N_7729,N_7519);
xor U8084 (N_8084,N_7928,N_7772);
or U8085 (N_8085,N_7785,N_7697);
nor U8086 (N_8086,N_7639,N_7610);
and U8087 (N_8087,N_7892,N_7780);
nand U8088 (N_8088,N_7512,N_7724);
or U8089 (N_8089,N_7806,N_7824);
nor U8090 (N_8090,N_7886,N_7853);
nand U8091 (N_8091,N_7661,N_7909);
or U8092 (N_8092,N_7860,N_7502);
and U8093 (N_8093,N_7592,N_7520);
and U8094 (N_8094,N_7947,N_7604);
xnor U8095 (N_8095,N_7856,N_7855);
nor U8096 (N_8096,N_7621,N_7707);
nand U8097 (N_8097,N_7647,N_7717);
nand U8098 (N_8098,N_7666,N_7945);
nand U8099 (N_8099,N_7783,N_7700);
or U8100 (N_8100,N_7706,N_7884);
and U8101 (N_8101,N_7955,N_7958);
nor U8102 (N_8102,N_7535,N_7867);
and U8103 (N_8103,N_7865,N_7587);
and U8104 (N_8104,N_7567,N_7774);
and U8105 (N_8105,N_7870,N_7619);
or U8106 (N_8106,N_7883,N_7628);
nand U8107 (N_8107,N_7575,N_7719);
and U8108 (N_8108,N_7913,N_7889);
nand U8109 (N_8109,N_7744,N_7770);
or U8110 (N_8110,N_7555,N_7852);
xnor U8111 (N_8111,N_7600,N_7796);
or U8112 (N_8112,N_7747,N_7859);
nand U8113 (N_8113,N_7957,N_7582);
and U8114 (N_8114,N_7710,N_7797);
or U8115 (N_8115,N_7993,N_7733);
and U8116 (N_8116,N_7572,N_7571);
or U8117 (N_8117,N_7833,N_7544);
or U8118 (N_8118,N_7672,N_7651);
or U8119 (N_8119,N_7830,N_7869);
nand U8120 (N_8120,N_7838,N_7631);
nand U8121 (N_8121,N_7576,N_7828);
nand U8122 (N_8122,N_7956,N_7835);
nor U8123 (N_8123,N_7515,N_7713);
and U8124 (N_8124,N_7542,N_7659);
nand U8125 (N_8125,N_7546,N_7862);
nand U8126 (N_8126,N_7812,N_7842);
or U8127 (N_8127,N_7645,N_7777);
xnor U8128 (N_8128,N_7979,N_7702);
nor U8129 (N_8129,N_7829,N_7820);
nor U8130 (N_8130,N_7872,N_7781);
nand U8131 (N_8131,N_7635,N_7590);
xnor U8132 (N_8132,N_7734,N_7766);
nor U8133 (N_8133,N_7521,N_7917);
nand U8134 (N_8134,N_7997,N_7844);
nand U8135 (N_8135,N_7728,N_7529);
nor U8136 (N_8136,N_7689,N_7539);
xnor U8137 (N_8137,N_7880,N_7756);
nand U8138 (N_8138,N_7517,N_7825);
and U8139 (N_8139,N_7578,N_7793);
or U8140 (N_8140,N_7834,N_7620);
and U8141 (N_8141,N_7537,N_7742);
or U8142 (N_8142,N_7877,N_7549);
nand U8143 (N_8143,N_7623,N_7650);
and U8144 (N_8144,N_7563,N_7750);
or U8145 (N_8145,N_7973,N_7857);
and U8146 (N_8146,N_7790,N_7591);
nor U8147 (N_8147,N_7799,N_7921);
nand U8148 (N_8148,N_7669,N_7594);
nand U8149 (N_8149,N_7723,N_7761);
or U8150 (N_8150,N_7826,N_7789);
and U8151 (N_8151,N_7568,N_7794);
nor U8152 (N_8152,N_7753,N_7670);
and U8153 (N_8153,N_7738,N_7718);
or U8154 (N_8154,N_7532,N_7500);
nand U8155 (N_8155,N_7943,N_7974);
and U8156 (N_8156,N_7784,N_7895);
nand U8157 (N_8157,N_7768,N_7674);
nand U8158 (N_8158,N_7543,N_7959);
or U8159 (N_8159,N_7686,N_7646);
nand U8160 (N_8160,N_7699,N_7887);
nand U8161 (N_8161,N_7509,N_7547);
xor U8162 (N_8162,N_7931,N_7605);
and U8163 (N_8163,N_7961,N_7813);
nand U8164 (N_8164,N_7680,N_7581);
or U8165 (N_8165,N_7714,N_7545);
or U8166 (N_8166,N_7641,N_7919);
and U8167 (N_8167,N_7910,N_7755);
nand U8168 (N_8168,N_7507,N_7760);
nand U8169 (N_8169,N_7802,N_7732);
or U8170 (N_8170,N_7675,N_7642);
xnor U8171 (N_8171,N_7952,N_7754);
xor U8172 (N_8172,N_7924,N_7655);
nor U8173 (N_8173,N_7786,N_7845);
nand U8174 (N_8174,N_7808,N_7759);
nor U8175 (N_8175,N_7560,N_7933);
and U8176 (N_8176,N_7846,N_7962);
and U8177 (N_8177,N_7696,N_7773);
or U8178 (N_8178,N_7903,N_7570);
nand U8179 (N_8179,N_7527,N_7606);
nand U8180 (N_8180,N_7876,N_7678);
nand U8181 (N_8181,N_7941,N_7683);
and U8182 (N_8182,N_7911,N_7528);
and U8183 (N_8183,N_7905,N_7951);
or U8184 (N_8184,N_7598,N_7554);
nor U8185 (N_8185,N_7929,N_7868);
and U8186 (N_8186,N_7757,N_7667);
nor U8187 (N_8187,N_7741,N_7556);
nor U8188 (N_8188,N_7712,N_7875);
and U8189 (N_8189,N_7565,N_7792);
xnor U8190 (N_8190,N_7687,N_7705);
nand U8191 (N_8191,N_7916,N_7513);
or U8192 (N_8192,N_7969,N_7915);
nor U8193 (N_8193,N_7900,N_7531);
and U8194 (N_8194,N_7632,N_7541);
or U8195 (N_8195,N_7608,N_7798);
nor U8196 (N_8196,N_7676,N_7612);
nor U8197 (N_8197,N_7540,N_7599);
nand U8198 (N_8198,N_7636,N_7552);
nor U8199 (N_8199,N_7584,N_7613);
or U8200 (N_8200,N_7640,N_7914);
nand U8201 (N_8201,N_7990,N_7657);
nor U8202 (N_8202,N_7893,N_7562);
and U8203 (N_8203,N_7918,N_7633);
nand U8204 (N_8204,N_7782,N_7839);
or U8205 (N_8205,N_7912,N_7927);
and U8206 (N_8206,N_7897,N_7982);
or U8207 (N_8207,N_7779,N_7991);
and U8208 (N_8208,N_7965,N_7776);
or U8209 (N_8209,N_7624,N_7561);
or U8210 (N_8210,N_7688,N_7763);
nand U8211 (N_8211,N_7597,N_7822);
and U8212 (N_8212,N_7925,N_7988);
nand U8213 (N_8213,N_7730,N_7701);
and U8214 (N_8214,N_7807,N_7890);
xor U8215 (N_8215,N_7999,N_7953);
nand U8216 (N_8216,N_7735,N_7954);
nor U8217 (N_8217,N_7654,N_7665);
and U8218 (N_8218,N_7746,N_7557);
nand U8219 (N_8219,N_7671,N_7975);
nand U8220 (N_8220,N_7630,N_7866);
nor U8221 (N_8221,N_7996,N_7989);
and U8222 (N_8222,N_7891,N_7603);
and U8223 (N_8223,N_7533,N_7749);
and U8224 (N_8224,N_7923,N_7948);
nand U8225 (N_8225,N_7609,N_7627);
and U8226 (N_8226,N_7966,N_7516);
and U8227 (N_8227,N_7553,N_7998);
or U8228 (N_8228,N_7936,N_7854);
xor U8229 (N_8229,N_7663,N_7622);
nor U8230 (N_8230,N_7593,N_7727);
or U8231 (N_8231,N_7849,N_7503);
nor U8232 (N_8232,N_7523,N_7981);
or U8233 (N_8233,N_7972,N_7778);
and U8234 (N_8234,N_7617,N_7684);
nand U8235 (N_8235,N_7638,N_7882);
nor U8236 (N_8236,N_7767,N_7803);
and U8237 (N_8237,N_7548,N_7564);
or U8238 (N_8238,N_7743,N_7653);
and U8239 (N_8239,N_7985,N_7580);
nor U8240 (N_8240,N_7837,N_7937);
nor U8241 (N_8241,N_7801,N_7668);
nor U8242 (N_8242,N_7946,N_7615);
nand U8243 (N_8243,N_7709,N_7847);
xnor U8244 (N_8244,N_7967,N_7899);
nand U8245 (N_8245,N_7506,N_7618);
xnor U8246 (N_8246,N_7586,N_7695);
and U8247 (N_8247,N_7637,N_7938);
xnor U8248 (N_8248,N_7904,N_7538);
and U8249 (N_8249,N_7879,N_7525);
nand U8250 (N_8250,N_7799,N_7894);
nor U8251 (N_8251,N_7647,N_7520);
or U8252 (N_8252,N_7904,N_7900);
nor U8253 (N_8253,N_7627,N_7636);
and U8254 (N_8254,N_7975,N_7701);
or U8255 (N_8255,N_7511,N_7522);
xor U8256 (N_8256,N_7847,N_7913);
nor U8257 (N_8257,N_7741,N_7935);
nand U8258 (N_8258,N_7565,N_7972);
nor U8259 (N_8259,N_7700,N_7747);
and U8260 (N_8260,N_7622,N_7926);
and U8261 (N_8261,N_7938,N_7583);
nand U8262 (N_8262,N_7656,N_7500);
nand U8263 (N_8263,N_7610,N_7839);
nor U8264 (N_8264,N_7601,N_7925);
nor U8265 (N_8265,N_7713,N_7640);
or U8266 (N_8266,N_7753,N_7709);
xnor U8267 (N_8267,N_7538,N_7780);
nand U8268 (N_8268,N_7632,N_7931);
nand U8269 (N_8269,N_7954,N_7811);
and U8270 (N_8270,N_7518,N_7984);
nor U8271 (N_8271,N_7980,N_7560);
nor U8272 (N_8272,N_7830,N_7517);
nor U8273 (N_8273,N_7597,N_7911);
and U8274 (N_8274,N_7984,N_7996);
or U8275 (N_8275,N_7911,N_7672);
xnor U8276 (N_8276,N_7934,N_7911);
nand U8277 (N_8277,N_7869,N_7849);
xor U8278 (N_8278,N_7828,N_7798);
nor U8279 (N_8279,N_7829,N_7953);
or U8280 (N_8280,N_7794,N_7719);
nand U8281 (N_8281,N_7678,N_7794);
and U8282 (N_8282,N_7873,N_7706);
or U8283 (N_8283,N_7751,N_7847);
or U8284 (N_8284,N_7740,N_7693);
nand U8285 (N_8285,N_7964,N_7958);
nand U8286 (N_8286,N_7966,N_7663);
or U8287 (N_8287,N_7830,N_7936);
and U8288 (N_8288,N_7896,N_7702);
and U8289 (N_8289,N_7743,N_7502);
and U8290 (N_8290,N_7968,N_7730);
or U8291 (N_8291,N_7510,N_7555);
or U8292 (N_8292,N_7757,N_7973);
nand U8293 (N_8293,N_7741,N_7675);
nor U8294 (N_8294,N_7536,N_7792);
nor U8295 (N_8295,N_7908,N_7590);
and U8296 (N_8296,N_7583,N_7961);
and U8297 (N_8297,N_7701,N_7934);
nor U8298 (N_8298,N_7724,N_7650);
or U8299 (N_8299,N_7926,N_7892);
nor U8300 (N_8300,N_7944,N_7790);
xnor U8301 (N_8301,N_7810,N_7949);
or U8302 (N_8302,N_7767,N_7998);
xnor U8303 (N_8303,N_7769,N_7831);
xor U8304 (N_8304,N_7901,N_7626);
nand U8305 (N_8305,N_7972,N_7751);
nor U8306 (N_8306,N_7789,N_7725);
nor U8307 (N_8307,N_7809,N_7912);
or U8308 (N_8308,N_7508,N_7599);
or U8309 (N_8309,N_7923,N_7633);
nand U8310 (N_8310,N_7745,N_7603);
nor U8311 (N_8311,N_7929,N_7853);
nor U8312 (N_8312,N_7650,N_7561);
or U8313 (N_8313,N_7715,N_7981);
and U8314 (N_8314,N_7920,N_7935);
or U8315 (N_8315,N_7721,N_7714);
and U8316 (N_8316,N_7927,N_7551);
nor U8317 (N_8317,N_7970,N_7992);
or U8318 (N_8318,N_7656,N_7732);
xor U8319 (N_8319,N_7702,N_7562);
or U8320 (N_8320,N_7724,N_7828);
nand U8321 (N_8321,N_7742,N_7604);
nor U8322 (N_8322,N_7942,N_7924);
and U8323 (N_8323,N_7633,N_7712);
and U8324 (N_8324,N_7928,N_7974);
nand U8325 (N_8325,N_7563,N_7624);
or U8326 (N_8326,N_7727,N_7913);
xor U8327 (N_8327,N_7769,N_7511);
nor U8328 (N_8328,N_7615,N_7854);
and U8329 (N_8329,N_7693,N_7526);
and U8330 (N_8330,N_7718,N_7804);
or U8331 (N_8331,N_7711,N_7816);
nor U8332 (N_8332,N_7823,N_7993);
or U8333 (N_8333,N_7806,N_7600);
or U8334 (N_8334,N_7513,N_7830);
nand U8335 (N_8335,N_7563,N_7920);
nor U8336 (N_8336,N_7941,N_7612);
and U8337 (N_8337,N_7928,N_7972);
xor U8338 (N_8338,N_7949,N_7747);
nand U8339 (N_8339,N_7773,N_7852);
nor U8340 (N_8340,N_7985,N_7971);
and U8341 (N_8341,N_7827,N_7622);
and U8342 (N_8342,N_7538,N_7706);
nor U8343 (N_8343,N_7709,N_7751);
and U8344 (N_8344,N_7583,N_7534);
nor U8345 (N_8345,N_7577,N_7584);
and U8346 (N_8346,N_7923,N_7733);
or U8347 (N_8347,N_7808,N_7769);
nor U8348 (N_8348,N_7941,N_7557);
nor U8349 (N_8349,N_7641,N_7642);
nand U8350 (N_8350,N_7720,N_7575);
nand U8351 (N_8351,N_7708,N_7817);
and U8352 (N_8352,N_7544,N_7566);
or U8353 (N_8353,N_7540,N_7611);
nand U8354 (N_8354,N_7735,N_7730);
and U8355 (N_8355,N_7793,N_7561);
nor U8356 (N_8356,N_7950,N_7925);
or U8357 (N_8357,N_7572,N_7752);
and U8358 (N_8358,N_7936,N_7793);
or U8359 (N_8359,N_7876,N_7930);
xor U8360 (N_8360,N_7891,N_7741);
and U8361 (N_8361,N_7840,N_7649);
nor U8362 (N_8362,N_7918,N_7833);
or U8363 (N_8363,N_7671,N_7714);
or U8364 (N_8364,N_7979,N_7680);
or U8365 (N_8365,N_7964,N_7529);
nor U8366 (N_8366,N_7548,N_7595);
and U8367 (N_8367,N_7793,N_7848);
and U8368 (N_8368,N_7929,N_7592);
nand U8369 (N_8369,N_7891,N_7957);
nor U8370 (N_8370,N_7978,N_7732);
nand U8371 (N_8371,N_7564,N_7970);
nand U8372 (N_8372,N_7875,N_7957);
nor U8373 (N_8373,N_7779,N_7939);
or U8374 (N_8374,N_7545,N_7732);
nand U8375 (N_8375,N_7609,N_7833);
and U8376 (N_8376,N_7624,N_7607);
and U8377 (N_8377,N_7949,N_7817);
or U8378 (N_8378,N_7847,N_7770);
or U8379 (N_8379,N_7587,N_7715);
nor U8380 (N_8380,N_7516,N_7576);
nand U8381 (N_8381,N_7521,N_7627);
nand U8382 (N_8382,N_7597,N_7990);
nand U8383 (N_8383,N_7522,N_7750);
nand U8384 (N_8384,N_7867,N_7500);
or U8385 (N_8385,N_7521,N_7690);
or U8386 (N_8386,N_7621,N_7862);
or U8387 (N_8387,N_7714,N_7980);
and U8388 (N_8388,N_7559,N_7842);
nor U8389 (N_8389,N_7699,N_7713);
xor U8390 (N_8390,N_7569,N_7619);
and U8391 (N_8391,N_7588,N_7811);
and U8392 (N_8392,N_7531,N_7865);
nor U8393 (N_8393,N_7824,N_7625);
nor U8394 (N_8394,N_7990,N_7953);
xor U8395 (N_8395,N_7730,N_7616);
nor U8396 (N_8396,N_7619,N_7644);
nand U8397 (N_8397,N_7814,N_7969);
nand U8398 (N_8398,N_7739,N_7828);
or U8399 (N_8399,N_7783,N_7591);
and U8400 (N_8400,N_7578,N_7517);
nor U8401 (N_8401,N_7840,N_7639);
or U8402 (N_8402,N_7971,N_7774);
and U8403 (N_8403,N_7732,N_7731);
and U8404 (N_8404,N_7599,N_7641);
xor U8405 (N_8405,N_7618,N_7743);
and U8406 (N_8406,N_7874,N_7797);
or U8407 (N_8407,N_7995,N_7923);
or U8408 (N_8408,N_7879,N_7698);
or U8409 (N_8409,N_7833,N_7786);
and U8410 (N_8410,N_7655,N_7734);
nand U8411 (N_8411,N_7608,N_7751);
and U8412 (N_8412,N_7567,N_7696);
nor U8413 (N_8413,N_7710,N_7942);
nor U8414 (N_8414,N_7713,N_7721);
nand U8415 (N_8415,N_7619,N_7701);
nor U8416 (N_8416,N_7955,N_7718);
and U8417 (N_8417,N_7514,N_7971);
or U8418 (N_8418,N_7551,N_7577);
nand U8419 (N_8419,N_7862,N_7615);
and U8420 (N_8420,N_7639,N_7563);
or U8421 (N_8421,N_7525,N_7869);
nor U8422 (N_8422,N_7770,N_7928);
nor U8423 (N_8423,N_7529,N_7655);
or U8424 (N_8424,N_7521,N_7520);
nor U8425 (N_8425,N_7909,N_7875);
nor U8426 (N_8426,N_7684,N_7702);
nand U8427 (N_8427,N_7761,N_7751);
nor U8428 (N_8428,N_7507,N_7677);
and U8429 (N_8429,N_7508,N_7695);
xnor U8430 (N_8430,N_7513,N_7511);
and U8431 (N_8431,N_7831,N_7868);
xor U8432 (N_8432,N_7533,N_7576);
nand U8433 (N_8433,N_7749,N_7659);
nand U8434 (N_8434,N_7915,N_7600);
nor U8435 (N_8435,N_7532,N_7986);
nand U8436 (N_8436,N_7884,N_7686);
xnor U8437 (N_8437,N_7590,N_7688);
nor U8438 (N_8438,N_7879,N_7815);
or U8439 (N_8439,N_7756,N_7743);
nor U8440 (N_8440,N_7549,N_7781);
or U8441 (N_8441,N_7929,N_7849);
or U8442 (N_8442,N_7689,N_7549);
and U8443 (N_8443,N_7942,N_7709);
nand U8444 (N_8444,N_7609,N_7983);
and U8445 (N_8445,N_7555,N_7761);
nand U8446 (N_8446,N_7679,N_7999);
nor U8447 (N_8447,N_7790,N_7873);
or U8448 (N_8448,N_7538,N_7796);
and U8449 (N_8449,N_7605,N_7595);
nand U8450 (N_8450,N_7617,N_7966);
nor U8451 (N_8451,N_7739,N_7592);
nand U8452 (N_8452,N_7974,N_7758);
or U8453 (N_8453,N_7630,N_7518);
or U8454 (N_8454,N_7795,N_7915);
or U8455 (N_8455,N_7884,N_7939);
xor U8456 (N_8456,N_7653,N_7592);
nand U8457 (N_8457,N_7693,N_7981);
nor U8458 (N_8458,N_7946,N_7844);
and U8459 (N_8459,N_7943,N_7818);
nor U8460 (N_8460,N_7863,N_7987);
nor U8461 (N_8461,N_7728,N_7647);
nand U8462 (N_8462,N_7965,N_7610);
nand U8463 (N_8463,N_7894,N_7519);
or U8464 (N_8464,N_7563,N_7676);
nand U8465 (N_8465,N_7994,N_7934);
or U8466 (N_8466,N_7978,N_7880);
nand U8467 (N_8467,N_7957,N_7679);
nand U8468 (N_8468,N_7909,N_7655);
and U8469 (N_8469,N_7650,N_7779);
nor U8470 (N_8470,N_7960,N_7616);
and U8471 (N_8471,N_7758,N_7731);
nor U8472 (N_8472,N_7869,N_7938);
and U8473 (N_8473,N_7583,N_7622);
nor U8474 (N_8474,N_7502,N_7951);
or U8475 (N_8475,N_7947,N_7560);
and U8476 (N_8476,N_7850,N_7814);
or U8477 (N_8477,N_7871,N_7649);
or U8478 (N_8478,N_7671,N_7928);
or U8479 (N_8479,N_7910,N_7695);
nor U8480 (N_8480,N_7673,N_7805);
nand U8481 (N_8481,N_7851,N_7986);
or U8482 (N_8482,N_7684,N_7878);
and U8483 (N_8483,N_7620,N_7706);
and U8484 (N_8484,N_7501,N_7984);
nand U8485 (N_8485,N_7558,N_7835);
or U8486 (N_8486,N_7523,N_7930);
or U8487 (N_8487,N_7565,N_7786);
xor U8488 (N_8488,N_7899,N_7652);
nand U8489 (N_8489,N_7859,N_7502);
xor U8490 (N_8490,N_7933,N_7839);
nor U8491 (N_8491,N_7721,N_7768);
nor U8492 (N_8492,N_7750,N_7963);
or U8493 (N_8493,N_7729,N_7887);
or U8494 (N_8494,N_7829,N_7752);
and U8495 (N_8495,N_7984,N_7818);
and U8496 (N_8496,N_7922,N_7719);
and U8497 (N_8497,N_7690,N_7626);
and U8498 (N_8498,N_7614,N_7987);
and U8499 (N_8499,N_7848,N_7620);
or U8500 (N_8500,N_8492,N_8463);
nand U8501 (N_8501,N_8167,N_8471);
nor U8502 (N_8502,N_8147,N_8429);
and U8503 (N_8503,N_8187,N_8390);
nor U8504 (N_8504,N_8459,N_8410);
and U8505 (N_8505,N_8242,N_8485);
nor U8506 (N_8506,N_8134,N_8046);
or U8507 (N_8507,N_8286,N_8338);
nand U8508 (N_8508,N_8297,N_8073);
nand U8509 (N_8509,N_8274,N_8316);
nand U8510 (N_8510,N_8189,N_8218);
or U8511 (N_8511,N_8498,N_8044);
or U8512 (N_8512,N_8381,N_8141);
and U8513 (N_8513,N_8118,N_8301);
nand U8514 (N_8514,N_8422,N_8039);
nor U8515 (N_8515,N_8121,N_8092);
nor U8516 (N_8516,N_8020,N_8227);
and U8517 (N_8517,N_8369,N_8409);
nor U8518 (N_8518,N_8013,N_8331);
nand U8519 (N_8519,N_8193,N_8220);
xor U8520 (N_8520,N_8265,N_8451);
nand U8521 (N_8521,N_8483,N_8185);
and U8522 (N_8522,N_8088,N_8418);
and U8523 (N_8523,N_8486,N_8241);
nand U8524 (N_8524,N_8181,N_8027);
nand U8525 (N_8525,N_8403,N_8380);
and U8526 (N_8526,N_8008,N_8499);
nor U8527 (N_8527,N_8014,N_8068);
xor U8528 (N_8528,N_8329,N_8405);
or U8529 (N_8529,N_8096,N_8466);
nand U8530 (N_8530,N_8469,N_8462);
or U8531 (N_8531,N_8011,N_8006);
nor U8532 (N_8532,N_8036,N_8294);
and U8533 (N_8533,N_8320,N_8079);
and U8534 (N_8534,N_8195,N_8012);
xnor U8535 (N_8535,N_8365,N_8256);
nand U8536 (N_8536,N_8076,N_8382);
nor U8537 (N_8537,N_8360,N_8254);
or U8538 (N_8538,N_8427,N_8154);
nand U8539 (N_8539,N_8392,N_8041);
and U8540 (N_8540,N_8186,N_8133);
and U8541 (N_8541,N_8450,N_8002);
nor U8542 (N_8542,N_8445,N_8435);
nand U8543 (N_8543,N_8055,N_8484);
nor U8544 (N_8544,N_8176,N_8225);
nor U8545 (N_8545,N_8414,N_8206);
nand U8546 (N_8546,N_8489,N_8053);
or U8547 (N_8547,N_8072,N_8109);
and U8548 (N_8548,N_8355,N_8430);
and U8549 (N_8549,N_8040,N_8395);
and U8550 (N_8550,N_8077,N_8091);
nor U8551 (N_8551,N_8303,N_8424);
or U8552 (N_8552,N_8122,N_8363);
and U8553 (N_8553,N_8477,N_8437);
nand U8554 (N_8554,N_8051,N_8143);
and U8555 (N_8555,N_8283,N_8070);
nand U8556 (N_8556,N_8413,N_8100);
and U8557 (N_8557,N_8065,N_8099);
or U8558 (N_8558,N_8194,N_8284);
xnor U8559 (N_8559,N_8362,N_8421);
nand U8560 (N_8560,N_8244,N_8131);
xor U8561 (N_8561,N_8114,N_8043);
and U8562 (N_8562,N_8037,N_8179);
nor U8563 (N_8563,N_8003,N_8416);
and U8564 (N_8564,N_8059,N_8432);
nor U8565 (N_8565,N_8084,N_8157);
and U8566 (N_8566,N_8064,N_8042);
nor U8567 (N_8567,N_8123,N_8394);
or U8568 (N_8568,N_8074,N_8191);
or U8569 (N_8569,N_8139,N_8386);
and U8570 (N_8570,N_8314,N_8032);
nand U8571 (N_8571,N_8080,N_8106);
nor U8572 (N_8572,N_8262,N_8232);
nand U8573 (N_8573,N_8278,N_8155);
nand U8574 (N_8574,N_8488,N_8052);
or U8575 (N_8575,N_8095,N_8023);
nor U8576 (N_8576,N_8468,N_8457);
or U8577 (N_8577,N_8183,N_8145);
and U8578 (N_8578,N_8368,N_8307);
nand U8579 (N_8579,N_8190,N_8067);
or U8580 (N_8580,N_8196,N_8018);
nand U8581 (N_8581,N_8169,N_8470);
or U8582 (N_8582,N_8302,N_8247);
nor U8583 (N_8583,N_8211,N_8366);
nand U8584 (N_8584,N_8340,N_8028);
nor U8585 (N_8585,N_8407,N_8330);
nor U8586 (N_8586,N_8325,N_8458);
or U8587 (N_8587,N_8175,N_8045);
or U8588 (N_8588,N_8280,N_8214);
and U8589 (N_8589,N_8226,N_8162);
nor U8590 (N_8590,N_8184,N_8022);
or U8591 (N_8591,N_8347,N_8357);
and U8592 (N_8592,N_8085,N_8015);
and U8593 (N_8593,N_8149,N_8017);
nor U8594 (N_8594,N_8370,N_8377);
xnor U8595 (N_8595,N_8354,N_8257);
nand U8596 (N_8596,N_8465,N_8245);
nand U8597 (N_8597,N_8219,N_8078);
nand U8598 (N_8598,N_8446,N_8229);
or U8599 (N_8599,N_8476,N_8481);
xnor U8600 (N_8600,N_8246,N_8269);
nor U8601 (N_8601,N_8361,N_8495);
nor U8602 (N_8602,N_8060,N_8066);
xnor U8603 (N_8603,N_8172,N_8038);
nor U8604 (N_8604,N_8127,N_8261);
xor U8605 (N_8605,N_8001,N_8397);
nand U8606 (N_8606,N_8019,N_8433);
nand U8607 (N_8607,N_8200,N_8428);
nor U8608 (N_8608,N_8393,N_8454);
nand U8609 (N_8609,N_8115,N_8335);
and U8610 (N_8610,N_8479,N_8299);
nand U8611 (N_8611,N_8308,N_8375);
nor U8612 (N_8612,N_8238,N_8062);
nand U8613 (N_8613,N_8102,N_8034);
or U8614 (N_8614,N_8310,N_8058);
nand U8615 (N_8615,N_8222,N_8097);
nand U8616 (N_8616,N_8388,N_8290);
xnor U8617 (N_8617,N_8321,N_8332);
nand U8618 (N_8618,N_8268,N_8341);
nand U8619 (N_8619,N_8272,N_8048);
and U8620 (N_8620,N_8164,N_8082);
and U8621 (N_8621,N_8137,N_8306);
and U8622 (N_8622,N_8103,N_8083);
and U8623 (N_8623,N_8236,N_8209);
nor U8624 (N_8624,N_8152,N_8231);
nand U8625 (N_8625,N_8266,N_8442);
or U8626 (N_8626,N_8417,N_8174);
or U8627 (N_8627,N_8420,N_8075);
xor U8628 (N_8628,N_8201,N_8258);
nor U8629 (N_8629,N_8124,N_8161);
and U8630 (N_8630,N_8087,N_8223);
nand U8631 (N_8631,N_8431,N_8300);
nor U8632 (N_8632,N_8318,N_8259);
nand U8633 (N_8633,N_8260,N_8192);
and U8634 (N_8634,N_8163,N_8344);
or U8635 (N_8635,N_8132,N_8090);
and U8636 (N_8636,N_8173,N_8285);
or U8637 (N_8637,N_8293,N_8452);
nor U8638 (N_8638,N_8271,N_8342);
or U8639 (N_8639,N_8309,N_8210);
or U8640 (N_8640,N_8276,N_8061);
or U8641 (N_8641,N_8251,N_8408);
nor U8642 (N_8642,N_8202,N_8295);
or U8643 (N_8643,N_8093,N_8383);
or U8644 (N_8644,N_8205,N_8021);
xnor U8645 (N_8645,N_8033,N_8472);
nor U8646 (N_8646,N_8497,N_8116);
nor U8647 (N_8647,N_8277,N_8327);
and U8648 (N_8648,N_8402,N_8024);
and U8649 (N_8649,N_8108,N_8343);
or U8650 (N_8650,N_8009,N_8352);
nor U8651 (N_8651,N_8279,N_8156);
nor U8652 (N_8652,N_8140,N_8292);
nand U8653 (N_8653,N_8030,N_8004);
xor U8654 (N_8654,N_8168,N_8112);
nor U8655 (N_8655,N_8107,N_8010);
or U8656 (N_8656,N_8081,N_8025);
nand U8657 (N_8657,N_8119,N_8101);
nand U8658 (N_8658,N_8399,N_8204);
or U8659 (N_8659,N_8224,N_8166);
nand U8660 (N_8660,N_8125,N_8425);
xor U8661 (N_8661,N_8339,N_8304);
and U8662 (N_8662,N_8456,N_8197);
nand U8663 (N_8663,N_8056,N_8263);
nand U8664 (N_8664,N_8412,N_8391);
and U8665 (N_8665,N_8270,N_8378);
nor U8666 (N_8666,N_8207,N_8250);
nor U8667 (N_8667,N_8372,N_8171);
nor U8668 (N_8668,N_8319,N_8094);
or U8669 (N_8669,N_8221,N_8291);
and U8670 (N_8670,N_8135,N_8128);
or U8671 (N_8671,N_8063,N_8473);
nand U8672 (N_8672,N_8358,N_8120);
xor U8673 (N_8673,N_8373,N_8482);
nand U8674 (N_8674,N_8117,N_8016);
or U8675 (N_8675,N_8349,N_8239);
or U8676 (N_8676,N_8324,N_8203);
and U8677 (N_8677,N_8089,N_8346);
nor U8678 (N_8678,N_8364,N_8404);
nor U8679 (N_8679,N_8480,N_8000);
nor U8680 (N_8680,N_8490,N_8287);
nand U8681 (N_8681,N_8423,N_8475);
nand U8682 (N_8682,N_8144,N_8252);
nor U8683 (N_8683,N_8031,N_8464);
nand U8684 (N_8684,N_8129,N_8275);
nand U8685 (N_8685,N_8182,N_8448);
and U8686 (N_8686,N_8359,N_8379);
nor U8687 (N_8687,N_8385,N_8345);
or U8688 (N_8688,N_8105,N_8350);
nor U8689 (N_8689,N_8281,N_8406);
or U8690 (N_8690,N_8426,N_8334);
or U8691 (N_8691,N_8353,N_8216);
nor U8692 (N_8692,N_8026,N_8213);
xnor U8693 (N_8693,N_8142,N_8496);
xnor U8694 (N_8694,N_8313,N_8315);
nand U8695 (N_8695,N_8312,N_8057);
nand U8696 (N_8696,N_8208,N_8180);
and U8697 (N_8697,N_8071,N_8323);
and U8698 (N_8698,N_8461,N_8449);
or U8699 (N_8699,N_8151,N_8298);
xnor U8700 (N_8700,N_8326,N_8438);
nand U8701 (N_8701,N_8444,N_8411);
nand U8702 (N_8702,N_8237,N_8165);
or U8703 (N_8703,N_8153,N_8282);
nand U8704 (N_8704,N_8337,N_8367);
xnor U8705 (N_8705,N_8267,N_8170);
nand U8706 (N_8706,N_8086,N_8047);
xor U8707 (N_8707,N_8126,N_8098);
or U8708 (N_8708,N_8374,N_8460);
nand U8709 (N_8709,N_8322,N_8371);
or U8710 (N_8710,N_8493,N_8264);
or U8711 (N_8711,N_8248,N_8328);
and U8712 (N_8712,N_8387,N_8447);
or U8713 (N_8713,N_8443,N_8400);
or U8714 (N_8714,N_8138,N_8249);
nor U8715 (N_8715,N_8178,N_8401);
and U8716 (N_8716,N_8255,N_8240);
nand U8717 (N_8717,N_8069,N_8376);
nand U8718 (N_8718,N_8351,N_8029);
or U8719 (N_8719,N_8317,N_8113);
nor U8720 (N_8720,N_8333,N_8305);
nand U8721 (N_8721,N_8441,N_8478);
and U8722 (N_8722,N_8289,N_8136);
and U8723 (N_8723,N_8311,N_8158);
and U8724 (N_8724,N_8288,N_8440);
nand U8725 (N_8725,N_8160,N_8111);
and U8726 (N_8726,N_8348,N_8198);
and U8727 (N_8727,N_8035,N_8110);
nand U8728 (N_8728,N_8230,N_8336);
and U8729 (N_8729,N_8217,N_8007);
or U8730 (N_8730,N_8296,N_8474);
nor U8731 (N_8731,N_8273,N_8235);
or U8732 (N_8732,N_8491,N_8243);
xnor U8733 (N_8733,N_8054,N_8455);
or U8734 (N_8734,N_8005,N_8439);
nand U8735 (N_8735,N_8253,N_8228);
nor U8736 (N_8736,N_8130,N_8050);
nor U8737 (N_8737,N_8159,N_8396);
nand U8738 (N_8738,N_8215,N_8419);
nand U8739 (N_8739,N_8199,N_8467);
nand U8740 (N_8740,N_8487,N_8177);
nor U8741 (N_8741,N_8494,N_8234);
or U8742 (N_8742,N_8146,N_8233);
nand U8743 (N_8743,N_8389,N_8212);
or U8744 (N_8744,N_8415,N_8148);
and U8745 (N_8745,N_8104,N_8150);
nor U8746 (N_8746,N_8398,N_8356);
xnor U8747 (N_8747,N_8384,N_8188);
and U8748 (N_8748,N_8436,N_8434);
and U8749 (N_8749,N_8049,N_8453);
nor U8750 (N_8750,N_8422,N_8341);
nor U8751 (N_8751,N_8294,N_8020);
or U8752 (N_8752,N_8025,N_8252);
and U8753 (N_8753,N_8233,N_8204);
nor U8754 (N_8754,N_8138,N_8489);
and U8755 (N_8755,N_8028,N_8097);
or U8756 (N_8756,N_8466,N_8157);
and U8757 (N_8757,N_8032,N_8113);
nor U8758 (N_8758,N_8048,N_8119);
and U8759 (N_8759,N_8111,N_8479);
nor U8760 (N_8760,N_8396,N_8499);
and U8761 (N_8761,N_8056,N_8395);
or U8762 (N_8762,N_8130,N_8128);
nor U8763 (N_8763,N_8214,N_8483);
nor U8764 (N_8764,N_8468,N_8209);
nor U8765 (N_8765,N_8110,N_8332);
and U8766 (N_8766,N_8347,N_8166);
nand U8767 (N_8767,N_8227,N_8358);
and U8768 (N_8768,N_8274,N_8009);
nand U8769 (N_8769,N_8472,N_8332);
and U8770 (N_8770,N_8323,N_8077);
or U8771 (N_8771,N_8270,N_8430);
or U8772 (N_8772,N_8284,N_8034);
and U8773 (N_8773,N_8076,N_8249);
or U8774 (N_8774,N_8461,N_8211);
and U8775 (N_8775,N_8245,N_8118);
and U8776 (N_8776,N_8169,N_8187);
nand U8777 (N_8777,N_8026,N_8465);
or U8778 (N_8778,N_8314,N_8394);
xor U8779 (N_8779,N_8394,N_8102);
nor U8780 (N_8780,N_8408,N_8000);
or U8781 (N_8781,N_8200,N_8138);
nand U8782 (N_8782,N_8244,N_8453);
nor U8783 (N_8783,N_8447,N_8108);
nor U8784 (N_8784,N_8217,N_8198);
or U8785 (N_8785,N_8161,N_8113);
and U8786 (N_8786,N_8217,N_8077);
nor U8787 (N_8787,N_8162,N_8211);
nor U8788 (N_8788,N_8311,N_8473);
nor U8789 (N_8789,N_8345,N_8078);
xor U8790 (N_8790,N_8252,N_8096);
or U8791 (N_8791,N_8360,N_8151);
and U8792 (N_8792,N_8364,N_8139);
nand U8793 (N_8793,N_8109,N_8187);
nor U8794 (N_8794,N_8113,N_8200);
nor U8795 (N_8795,N_8352,N_8482);
or U8796 (N_8796,N_8424,N_8339);
or U8797 (N_8797,N_8445,N_8084);
nand U8798 (N_8798,N_8066,N_8009);
and U8799 (N_8799,N_8194,N_8174);
or U8800 (N_8800,N_8047,N_8114);
or U8801 (N_8801,N_8452,N_8378);
nor U8802 (N_8802,N_8002,N_8098);
nand U8803 (N_8803,N_8444,N_8182);
and U8804 (N_8804,N_8283,N_8393);
or U8805 (N_8805,N_8188,N_8028);
nand U8806 (N_8806,N_8387,N_8068);
xor U8807 (N_8807,N_8172,N_8174);
and U8808 (N_8808,N_8239,N_8460);
nor U8809 (N_8809,N_8470,N_8163);
nor U8810 (N_8810,N_8001,N_8498);
or U8811 (N_8811,N_8008,N_8030);
xnor U8812 (N_8812,N_8071,N_8017);
nor U8813 (N_8813,N_8091,N_8454);
nand U8814 (N_8814,N_8055,N_8342);
nor U8815 (N_8815,N_8225,N_8491);
xor U8816 (N_8816,N_8365,N_8484);
nor U8817 (N_8817,N_8076,N_8332);
nand U8818 (N_8818,N_8095,N_8363);
nand U8819 (N_8819,N_8035,N_8037);
and U8820 (N_8820,N_8234,N_8086);
xnor U8821 (N_8821,N_8086,N_8287);
and U8822 (N_8822,N_8434,N_8471);
and U8823 (N_8823,N_8217,N_8058);
or U8824 (N_8824,N_8279,N_8177);
or U8825 (N_8825,N_8151,N_8356);
or U8826 (N_8826,N_8450,N_8144);
nand U8827 (N_8827,N_8154,N_8305);
nand U8828 (N_8828,N_8135,N_8295);
and U8829 (N_8829,N_8182,N_8280);
nand U8830 (N_8830,N_8017,N_8356);
or U8831 (N_8831,N_8379,N_8490);
or U8832 (N_8832,N_8338,N_8434);
nand U8833 (N_8833,N_8158,N_8288);
and U8834 (N_8834,N_8425,N_8333);
nand U8835 (N_8835,N_8074,N_8143);
nand U8836 (N_8836,N_8397,N_8010);
nor U8837 (N_8837,N_8043,N_8268);
nand U8838 (N_8838,N_8258,N_8316);
or U8839 (N_8839,N_8094,N_8449);
and U8840 (N_8840,N_8101,N_8422);
nand U8841 (N_8841,N_8267,N_8425);
nand U8842 (N_8842,N_8123,N_8230);
and U8843 (N_8843,N_8192,N_8080);
and U8844 (N_8844,N_8483,N_8320);
and U8845 (N_8845,N_8393,N_8338);
and U8846 (N_8846,N_8453,N_8364);
and U8847 (N_8847,N_8041,N_8160);
nor U8848 (N_8848,N_8069,N_8253);
nand U8849 (N_8849,N_8449,N_8230);
and U8850 (N_8850,N_8307,N_8430);
and U8851 (N_8851,N_8382,N_8142);
nor U8852 (N_8852,N_8154,N_8315);
nor U8853 (N_8853,N_8442,N_8213);
nand U8854 (N_8854,N_8036,N_8184);
nand U8855 (N_8855,N_8174,N_8474);
nand U8856 (N_8856,N_8378,N_8039);
or U8857 (N_8857,N_8028,N_8181);
nand U8858 (N_8858,N_8445,N_8346);
or U8859 (N_8859,N_8278,N_8223);
or U8860 (N_8860,N_8145,N_8297);
nor U8861 (N_8861,N_8115,N_8189);
nor U8862 (N_8862,N_8479,N_8180);
and U8863 (N_8863,N_8009,N_8425);
or U8864 (N_8864,N_8035,N_8303);
nand U8865 (N_8865,N_8311,N_8174);
nor U8866 (N_8866,N_8280,N_8069);
or U8867 (N_8867,N_8339,N_8338);
nor U8868 (N_8868,N_8446,N_8120);
and U8869 (N_8869,N_8440,N_8418);
and U8870 (N_8870,N_8319,N_8375);
or U8871 (N_8871,N_8498,N_8256);
nor U8872 (N_8872,N_8058,N_8463);
nor U8873 (N_8873,N_8095,N_8146);
xor U8874 (N_8874,N_8165,N_8344);
nor U8875 (N_8875,N_8422,N_8277);
or U8876 (N_8876,N_8425,N_8318);
and U8877 (N_8877,N_8342,N_8224);
and U8878 (N_8878,N_8022,N_8476);
nand U8879 (N_8879,N_8181,N_8095);
nor U8880 (N_8880,N_8445,N_8234);
or U8881 (N_8881,N_8390,N_8477);
nor U8882 (N_8882,N_8339,N_8075);
or U8883 (N_8883,N_8415,N_8419);
nand U8884 (N_8884,N_8128,N_8283);
or U8885 (N_8885,N_8052,N_8172);
nor U8886 (N_8886,N_8390,N_8108);
and U8887 (N_8887,N_8340,N_8196);
or U8888 (N_8888,N_8101,N_8133);
nand U8889 (N_8889,N_8474,N_8277);
nand U8890 (N_8890,N_8226,N_8137);
xnor U8891 (N_8891,N_8072,N_8038);
xor U8892 (N_8892,N_8276,N_8458);
or U8893 (N_8893,N_8096,N_8168);
nor U8894 (N_8894,N_8233,N_8033);
and U8895 (N_8895,N_8062,N_8245);
nand U8896 (N_8896,N_8261,N_8385);
nand U8897 (N_8897,N_8033,N_8481);
nand U8898 (N_8898,N_8009,N_8251);
and U8899 (N_8899,N_8004,N_8375);
nor U8900 (N_8900,N_8113,N_8310);
nand U8901 (N_8901,N_8040,N_8343);
xor U8902 (N_8902,N_8302,N_8423);
nor U8903 (N_8903,N_8175,N_8144);
nor U8904 (N_8904,N_8052,N_8142);
nor U8905 (N_8905,N_8066,N_8236);
nor U8906 (N_8906,N_8031,N_8366);
nor U8907 (N_8907,N_8331,N_8433);
or U8908 (N_8908,N_8122,N_8316);
and U8909 (N_8909,N_8466,N_8128);
nand U8910 (N_8910,N_8108,N_8311);
nor U8911 (N_8911,N_8217,N_8169);
or U8912 (N_8912,N_8494,N_8114);
nor U8913 (N_8913,N_8238,N_8317);
nor U8914 (N_8914,N_8312,N_8442);
or U8915 (N_8915,N_8479,N_8400);
or U8916 (N_8916,N_8115,N_8183);
xnor U8917 (N_8917,N_8428,N_8256);
nor U8918 (N_8918,N_8293,N_8154);
and U8919 (N_8919,N_8354,N_8015);
xnor U8920 (N_8920,N_8474,N_8178);
xnor U8921 (N_8921,N_8480,N_8256);
nand U8922 (N_8922,N_8458,N_8314);
nor U8923 (N_8923,N_8484,N_8139);
nand U8924 (N_8924,N_8127,N_8072);
xor U8925 (N_8925,N_8280,N_8025);
nand U8926 (N_8926,N_8341,N_8221);
and U8927 (N_8927,N_8114,N_8361);
nand U8928 (N_8928,N_8084,N_8325);
nand U8929 (N_8929,N_8343,N_8332);
nor U8930 (N_8930,N_8312,N_8002);
xor U8931 (N_8931,N_8353,N_8245);
xnor U8932 (N_8932,N_8271,N_8402);
or U8933 (N_8933,N_8145,N_8036);
xor U8934 (N_8934,N_8115,N_8205);
nor U8935 (N_8935,N_8149,N_8099);
or U8936 (N_8936,N_8449,N_8161);
nand U8937 (N_8937,N_8391,N_8124);
nand U8938 (N_8938,N_8075,N_8252);
or U8939 (N_8939,N_8035,N_8308);
nand U8940 (N_8940,N_8161,N_8294);
nor U8941 (N_8941,N_8442,N_8062);
and U8942 (N_8942,N_8053,N_8327);
nor U8943 (N_8943,N_8437,N_8087);
or U8944 (N_8944,N_8287,N_8128);
nor U8945 (N_8945,N_8439,N_8207);
xor U8946 (N_8946,N_8282,N_8184);
nor U8947 (N_8947,N_8467,N_8205);
nand U8948 (N_8948,N_8377,N_8371);
or U8949 (N_8949,N_8057,N_8439);
nor U8950 (N_8950,N_8029,N_8253);
nor U8951 (N_8951,N_8139,N_8109);
and U8952 (N_8952,N_8120,N_8323);
nand U8953 (N_8953,N_8475,N_8155);
and U8954 (N_8954,N_8232,N_8431);
and U8955 (N_8955,N_8482,N_8349);
and U8956 (N_8956,N_8339,N_8260);
nor U8957 (N_8957,N_8157,N_8484);
nand U8958 (N_8958,N_8358,N_8392);
and U8959 (N_8959,N_8114,N_8363);
xor U8960 (N_8960,N_8014,N_8016);
nand U8961 (N_8961,N_8082,N_8260);
or U8962 (N_8962,N_8204,N_8140);
nand U8963 (N_8963,N_8119,N_8478);
and U8964 (N_8964,N_8195,N_8015);
xor U8965 (N_8965,N_8268,N_8132);
nand U8966 (N_8966,N_8499,N_8181);
and U8967 (N_8967,N_8414,N_8471);
xnor U8968 (N_8968,N_8036,N_8108);
and U8969 (N_8969,N_8410,N_8009);
xor U8970 (N_8970,N_8412,N_8294);
or U8971 (N_8971,N_8260,N_8281);
nand U8972 (N_8972,N_8276,N_8309);
nand U8973 (N_8973,N_8289,N_8176);
nand U8974 (N_8974,N_8330,N_8372);
nor U8975 (N_8975,N_8393,N_8199);
or U8976 (N_8976,N_8364,N_8279);
and U8977 (N_8977,N_8311,N_8334);
and U8978 (N_8978,N_8061,N_8143);
and U8979 (N_8979,N_8069,N_8334);
nand U8980 (N_8980,N_8336,N_8173);
and U8981 (N_8981,N_8164,N_8239);
or U8982 (N_8982,N_8261,N_8303);
nor U8983 (N_8983,N_8124,N_8142);
or U8984 (N_8984,N_8191,N_8026);
nor U8985 (N_8985,N_8048,N_8339);
nor U8986 (N_8986,N_8493,N_8247);
nor U8987 (N_8987,N_8006,N_8195);
and U8988 (N_8988,N_8498,N_8209);
nor U8989 (N_8989,N_8468,N_8185);
nor U8990 (N_8990,N_8073,N_8027);
and U8991 (N_8991,N_8221,N_8239);
nand U8992 (N_8992,N_8181,N_8458);
nand U8993 (N_8993,N_8484,N_8111);
nor U8994 (N_8994,N_8131,N_8304);
and U8995 (N_8995,N_8455,N_8092);
xnor U8996 (N_8996,N_8087,N_8352);
or U8997 (N_8997,N_8419,N_8388);
or U8998 (N_8998,N_8425,N_8355);
nor U8999 (N_8999,N_8137,N_8345);
or U9000 (N_9000,N_8670,N_8547);
nor U9001 (N_9001,N_8521,N_8714);
nand U9002 (N_9002,N_8910,N_8921);
and U9003 (N_9003,N_8880,N_8848);
nor U9004 (N_9004,N_8805,N_8631);
nor U9005 (N_9005,N_8620,N_8876);
nor U9006 (N_9006,N_8702,N_8622);
nor U9007 (N_9007,N_8500,N_8685);
or U9008 (N_9008,N_8992,N_8891);
or U9009 (N_9009,N_8802,N_8801);
xnor U9010 (N_9010,N_8882,N_8942);
nor U9011 (N_9011,N_8937,N_8572);
or U9012 (N_9012,N_8540,N_8683);
nor U9013 (N_9013,N_8774,N_8995);
and U9014 (N_9014,N_8971,N_8728);
or U9015 (N_9015,N_8958,N_8528);
nand U9016 (N_9016,N_8633,N_8546);
and U9017 (N_9017,N_8564,N_8752);
nand U9018 (N_9018,N_8798,N_8954);
and U9019 (N_9019,N_8539,N_8931);
and U9020 (N_9020,N_8713,N_8721);
nor U9021 (N_9021,N_8626,N_8587);
xor U9022 (N_9022,N_8803,N_8689);
nand U9023 (N_9023,N_8775,N_8696);
nand U9024 (N_9024,N_8823,N_8748);
nand U9025 (N_9025,N_8691,N_8744);
nand U9026 (N_9026,N_8705,N_8613);
and U9027 (N_9027,N_8973,N_8753);
or U9028 (N_9028,N_8665,N_8844);
and U9029 (N_9029,N_8680,N_8514);
and U9030 (N_9030,N_8896,N_8727);
or U9031 (N_9031,N_8655,N_8778);
nor U9032 (N_9032,N_8706,N_8825);
nand U9033 (N_9033,N_8980,N_8584);
or U9034 (N_9034,N_8981,N_8818);
or U9035 (N_9035,N_8535,N_8901);
and U9036 (N_9036,N_8905,N_8555);
nand U9037 (N_9037,N_8678,N_8758);
nand U9038 (N_9038,N_8791,N_8720);
and U9039 (N_9039,N_8501,N_8715);
or U9040 (N_9040,N_8976,N_8984);
nand U9041 (N_9041,N_8811,N_8900);
nand U9042 (N_9042,N_8765,N_8747);
xor U9043 (N_9043,N_8915,N_8703);
nor U9044 (N_9044,N_8993,N_8759);
nor U9045 (N_9045,N_8904,N_8754);
nor U9046 (N_9046,N_8527,N_8830);
xor U9047 (N_9047,N_8756,N_8847);
nor U9048 (N_9048,N_8570,N_8968);
nor U9049 (N_9049,N_8790,N_8870);
nand U9050 (N_9050,N_8855,N_8762);
and U9051 (N_9051,N_8615,N_8682);
nand U9052 (N_9052,N_8810,N_8813);
nand U9053 (N_9053,N_8738,N_8837);
nand U9054 (N_9054,N_8635,N_8533);
and U9055 (N_9055,N_8600,N_8530);
xnor U9056 (N_9056,N_8771,N_8663);
or U9057 (N_9057,N_8551,N_8578);
or U9058 (N_9058,N_8700,N_8939);
nor U9059 (N_9059,N_8671,N_8959);
nor U9060 (N_9060,N_8519,N_8918);
xor U9061 (N_9061,N_8674,N_8913);
nor U9062 (N_9062,N_8881,N_8781);
nor U9063 (N_9063,N_8977,N_8623);
nor U9064 (N_9064,N_8602,N_8567);
or U9065 (N_9065,N_8629,N_8816);
and U9066 (N_9066,N_8854,N_8831);
or U9067 (N_9067,N_8525,N_8941);
or U9068 (N_9068,N_8660,N_8757);
nand U9069 (N_9069,N_8554,N_8808);
xnor U9070 (N_9070,N_8944,N_8741);
nor U9071 (N_9071,N_8907,N_8859);
or U9072 (N_9072,N_8743,N_8897);
nor U9073 (N_9073,N_8725,N_8614);
nand U9074 (N_9074,N_8920,N_8645);
nand U9075 (N_9075,N_8783,N_8787);
and U9076 (N_9076,N_8866,N_8888);
nor U9077 (N_9077,N_8928,N_8822);
or U9078 (N_9078,N_8639,N_8940);
nand U9079 (N_9079,N_8863,N_8932);
and U9080 (N_9080,N_8961,N_8707);
or U9081 (N_9081,N_8693,N_8580);
nor U9082 (N_9082,N_8761,N_8886);
or U9083 (N_9083,N_8594,N_8768);
nor U9084 (N_9084,N_8731,N_8925);
nor U9085 (N_9085,N_8878,N_8826);
and U9086 (N_9086,N_8522,N_8652);
and U9087 (N_9087,N_8719,N_8601);
nand U9088 (N_9088,N_8688,N_8986);
nor U9089 (N_9089,N_8677,N_8617);
and U9090 (N_9090,N_8974,N_8767);
nand U9091 (N_9091,N_8516,N_8653);
nand U9092 (N_9092,N_8914,N_8618);
nand U9093 (N_9093,N_8573,N_8553);
nand U9094 (N_9094,N_8681,N_8972);
nand U9095 (N_9095,N_8912,N_8637);
nand U9096 (N_9096,N_8679,N_8899);
and U9097 (N_9097,N_8926,N_8951);
nand U9098 (N_9098,N_8793,N_8651);
and U9099 (N_9099,N_8504,N_8605);
nand U9100 (N_9100,N_8698,N_8890);
nor U9101 (N_9101,N_8979,N_8952);
and U9102 (N_9102,N_8934,N_8569);
nand U9103 (N_9103,N_8773,N_8879);
nor U9104 (N_9104,N_8789,N_8667);
nor U9105 (N_9105,N_8732,N_8656);
nor U9106 (N_9106,N_8794,N_8510);
xnor U9107 (N_9107,N_8591,N_8557);
nor U9108 (N_9108,N_8585,N_8887);
nor U9109 (N_9109,N_8627,N_8675);
nand U9110 (N_9110,N_8709,N_8566);
nor U9111 (N_9111,N_8865,N_8505);
nand U9112 (N_9112,N_8740,N_8832);
and U9113 (N_9113,N_8695,N_8529);
nor U9114 (N_9114,N_8745,N_8630);
or U9115 (N_9115,N_8593,N_8936);
nand U9116 (N_9116,N_8953,N_8603);
and U9117 (N_9117,N_8869,N_8735);
or U9118 (N_9118,N_8746,N_8697);
nand U9119 (N_9119,N_8838,N_8526);
or U9120 (N_9120,N_8909,N_8503);
xor U9121 (N_9121,N_8769,N_8906);
and U9122 (N_9122,N_8917,N_8710);
nand U9123 (N_9123,N_8807,N_8659);
xor U9124 (N_9124,N_8733,N_8842);
xnor U9125 (N_9125,N_8902,N_8970);
xnor U9126 (N_9126,N_8819,N_8956);
xnor U9127 (N_9127,N_8788,N_8922);
or U9128 (N_9128,N_8989,N_8895);
or U9129 (N_9129,N_8786,N_8898);
nand U9130 (N_9130,N_8751,N_8549);
nand U9131 (N_9131,N_8628,N_8829);
nand U9132 (N_9132,N_8929,N_8606);
and U9133 (N_9133,N_8843,N_8916);
nor U9134 (N_9134,N_8619,N_8571);
nand U9135 (N_9135,N_8556,N_8662);
nand U9136 (N_9136,N_8817,N_8650);
xnor U9137 (N_9137,N_8784,N_8574);
nor U9138 (N_9138,N_8550,N_8766);
xnor U9139 (N_9139,N_8581,N_8841);
nor U9140 (N_9140,N_8692,N_8647);
xnor U9141 (N_9141,N_8861,N_8779);
or U9142 (N_9142,N_8945,N_8795);
or U9143 (N_9143,N_8884,N_8845);
nand U9144 (N_9144,N_8800,N_8853);
and U9145 (N_9145,N_8799,N_8985);
nand U9146 (N_9146,N_8508,N_8621);
nand U9147 (N_9147,N_8770,N_8796);
nor U9148 (N_9148,N_8666,N_8988);
nor U9149 (N_9149,N_8634,N_8722);
or U9150 (N_9150,N_8777,N_8996);
xnor U9151 (N_9151,N_8669,N_8577);
nor U9152 (N_9152,N_8560,N_8576);
or U9153 (N_9153,N_8998,N_8860);
and U9154 (N_9154,N_8736,N_8946);
nor U9155 (N_9155,N_8718,N_8668);
nor U9156 (N_9156,N_8641,N_8792);
and U9157 (N_9157,N_8568,N_8604);
nor U9158 (N_9158,N_8924,N_8903);
or U9159 (N_9159,N_8933,N_8856);
nor U9160 (N_9160,N_8846,N_8563);
xor U9161 (N_9161,N_8644,N_8962);
nand U9162 (N_9162,N_8990,N_8542);
nor U9163 (N_9163,N_8686,N_8558);
nand U9164 (N_9164,N_8649,N_8515);
nand U9165 (N_9165,N_8820,N_8642);
nand U9166 (N_9166,N_8967,N_8726);
nand U9167 (N_9167,N_8716,N_8764);
nor U9168 (N_9168,N_8755,N_8955);
nor U9169 (N_9169,N_8923,N_8548);
and U9170 (N_9170,N_8852,N_8687);
xnor U9171 (N_9171,N_8894,N_8850);
nand U9172 (N_9172,N_8836,N_8908);
and U9173 (N_9173,N_8868,N_8699);
or U9174 (N_9174,N_8760,N_8780);
and U9175 (N_9175,N_8772,N_8930);
and U9176 (N_9176,N_8565,N_8885);
and U9177 (N_9177,N_8661,N_8763);
nand U9178 (N_9178,N_8806,N_8969);
and U9179 (N_9179,N_8724,N_8947);
or U9180 (N_9180,N_8911,N_8654);
or U9181 (N_9181,N_8561,N_8948);
or U9182 (N_9182,N_8867,N_8949);
or U9183 (N_9183,N_8541,N_8590);
xnor U9184 (N_9184,N_8597,N_8711);
nand U9185 (N_9185,N_8609,N_8610);
or U9186 (N_9186,N_8513,N_8797);
nand U9187 (N_9187,N_8592,N_8935);
or U9188 (N_9188,N_8632,N_8927);
or U9189 (N_9189,N_8648,N_8520);
nand U9190 (N_9190,N_8704,N_8809);
xnor U9191 (N_9191,N_8595,N_8730);
and U9192 (N_9192,N_8658,N_8717);
nor U9193 (N_9193,N_8750,N_8840);
xnor U9194 (N_9194,N_8994,N_8690);
and U9195 (N_9195,N_8858,N_8518);
and U9196 (N_9196,N_8776,N_8739);
nand U9197 (N_9197,N_8982,N_8512);
nor U9198 (N_9198,N_8599,N_8835);
nand U9199 (N_9199,N_8506,N_8643);
or U9200 (N_9200,N_8701,N_8749);
and U9201 (N_9201,N_8734,N_8598);
and U9202 (N_9202,N_8625,N_8960);
and U9203 (N_9203,N_8507,N_8544);
and U9204 (N_9204,N_8511,N_8532);
or U9205 (N_9205,N_8987,N_8943);
nand U9206 (N_9206,N_8871,N_8883);
or U9207 (N_9207,N_8536,N_8785);
or U9208 (N_9208,N_8729,N_8965);
nor U9209 (N_9209,N_8583,N_8531);
nor U9210 (N_9210,N_8607,N_8815);
nand U9211 (N_9211,N_8938,N_8638);
nand U9212 (N_9212,N_8657,N_8664);
nor U9213 (N_9213,N_8964,N_8684);
or U9214 (N_9214,N_8517,N_8646);
or U9215 (N_9215,N_8608,N_8636);
nand U9216 (N_9216,N_8824,N_8708);
nor U9217 (N_9217,N_8509,N_8712);
nor U9218 (N_9218,N_8849,N_8966);
nand U9219 (N_9219,N_8827,N_8534);
nor U9220 (N_9220,N_8812,N_8997);
or U9221 (N_9221,N_8611,N_8588);
xor U9222 (N_9222,N_8640,N_8804);
or U9223 (N_9223,N_8545,N_8612);
xor U9224 (N_9224,N_8596,N_8673);
or U9225 (N_9225,N_8872,N_8862);
nor U9226 (N_9226,N_8857,N_8502);
or U9227 (N_9227,N_8537,N_8991);
nand U9228 (N_9228,N_8828,N_8834);
and U9229 (N_9229,N_8983,N_8889);
nor U9230 (N_9230,N_8737,N_8851);
nor U9231 (N_9231,N_8833,N_8538);
or U9232 (N_9232,N_8575,N_8582);
nor U9233 (N_9233,N_8814,N_8742);
and U9234 (N_9234,N_8919,N_8579);
xnor U9235 (N_9235,N_8950,N_8893);
or U9236 (N_9236,N_8624,N_8978);
nand U9237 (N_9237,N_8975,N_8963);
or U9238 (N_9238,N_8723,N_8523);
xor U9239 (N_9239,N_8676,N_8874);
nand U9240 (N_9240,N_8864,N_8892);
and U9241 (N_9241,N_8821,N_8589);
nor U9242 (N_9242,N_8616,N_8957);
and U9243 (N_9243,N_8873,N_8694);
or U9244 (N_9244,N_8999,N_8559);
nor U9245 (N_9245,N_8524,N_8552);
nand U9246 (N_9246,N_8877,N_8562);
or U9247 (N_9247,N_8543,N_8586);
and U9248 (N_9248,N_8672,N_8839);
nand U9249 (N_9249,N_8875,N_8782);
or U9250 (N_9250,N_8729,N_8870);
and U9251 (N_9251,N_8602,N_8541);
nor U9252 (N_9252,N_8904,N_8660);
nor U9253 (N_9253,N_8991,N_8787);
nor U9254 (N_9254,N_8768,N_8837);
nor U9255 (N_9255,N_8938,N_8633);
or U9256 (N_9256,N_8955,N_8725);
nor U9257 (N_9257,N_8727,N_8761);
xor U9258 (N_9258,N_8556,N_8543);
nor U9259 (N_9259,N_8606,N_8850);
nor U9260 (N_9260,N_8513,N_8646);
or U9261 (N_9261,N_8936,N_8652);
nor U9262 (N_9262,N_8728,N_8752);
nor U9263 (N_9263,N_8718,N_8914);
or U9264 (N_9264,N_8518,N_8962);
or U9265 (N_9265,N_8786,N_8724);
or U9266 (N_9266,N_8525,N_8862);
or U9267 (N_9267,N_8718,N_8817);
xnor U9268 (N_9268,N_8886,N_8875);
or U9269 (N_9269,N_8845,N_8790);
and U9270 (N_9270,N_8707,N_8743);
nand U9271 (N_9271,N_8581,N_8617);
nor U9272 (N_9272,N_8643,N_8827);
xor U9273 (N_9273,N_8665,N_8694);
or U9274 (N_9274,N_8567,N_8970);
nand U9275 (N_9275,N_8504,N_8646);
nand U9276 (N_9276,N_8760,N_8706);
or U9277 (N_9277,N_8879,N_8651);
nand U9278 (N_9278,N_8776,N_8908);
and U9279 (N_9279,N_8902,N_8523);
nand U9280 (N_9280,N_8837,N_8870);
nor U9281 (N_9281,N_8673,N_8566);
and U9282 (N_9282,N_8896,N_8557);
nor U9283 (N_9283,N_8814,N_8651);
xnor U9284 (N_9284,N_8702,N_8874);
and U9285 (N_9285,N_8511,N_8935);
or U9286 (N_9286,N_8923,N_8542);
nor U9287 (N_9287,N_8728,N_8753);
nand U9288 (N_9288,N_8972,N_8574);
and U9289 (N_9289,N_8594,N_8562);
and U9290 (N_9290,N_8575,N_8946);
and U9291 (N_9291,N_8904,N_8921);
nand U9292 (N_9292,N_8633,N_8556);
nand U9293 (N_9293,N_8948,N_8595);
nand U9294 (N_9294,N_8616,N_8567);
nand U9295 (N_9295,N_8823,N_8955);
nand U9296 (N_9296,N_8825,N_8536);
nor U9297 (N_9297,N_8885,N_8519);
nand U9298 (N_9298,N_8692,N_8976);
xnor U9299 (N_9299,N_8516,N_8669);
xnor U9300 (N_9300,N_8935,N_8777);
nor U9301 (N_9301,N_8901,N_8602);
nand U9302 (N_9302,N_8643,N_8588);
and U9303 (N_9303,N_8944,N_8906);
nand U9304 (N_9304,N_8688,N_8944);
nand U9305 (N_9305,N_8598,N_8700);
nand U9306 (N_9306,N_8817,N_8531);
nor U9307 (N_9307,N_8999,N_8746);
and U9308 (N_9308,N_8683,N_8808);
nand U9309 (N_9309,N_8695,N_8577);
nor U9310 (N_9310,N_8888,N_8848);
nor U9311 (N_9311,N_8669,N_8744);
and U9312 (N_9312,N_8660,N_8900);
nor U9313 (N_9313,N_8962,N_8991);
and U9314 (N_9314,N_8880,N_8712);
or U9315 (N_9315,N_8642,N_8628);
nand U9316 (N_9316,N_8745,N_8652);
or U9317 (N_9317,N_8790,N_8862);
nor U9318 (N_9318,N_8621,N_8655);
nor U9319 (N_9319,N_8987,N_8721);
and U9320 (N_9320,N_8726,N_8596);
and U9321 (N_9321,N_8635,N_8683);
or U9322 (N_9322,N_8754,N_8966);
xor U9323 (N_9323,N_8664,N_8509);
or U9324 (N_9324,N_8503,N_8845);
nor U9325 (N_9325,N_8963,N_8709);
nor U9326 (N_9326,N_8723,N_8958);
xor U9327 (N_9327,N_8598,N_8502);
and U9328 (N_9328,N_8649,N_8845);
or U9329 (N_9329,N_8624,N_8787);
or U9330 (N_9330,N_8530,N_8755);
nand U9331 (N_9331,N_8776,N_8655);
nor U9332 (N_9332,N_8517,N_8624);
and U9333 (N_9333,N_8942,N_8900);
xor U9334 (N_9334,N_8592,N_8513);
and U9335 (N_9335,N_8984,N_8546);
or U9336 (N_9336,N_8623,N_8790);
and U9337 (N_9337,N_8864,N_8883);
and U9338 (N_9338,N_8640,N_8667);
and U9339 (N_9339,N_8994,N_8612);
or U9340 (N_9340,N_8513,N_8685);
nor U9341 (N_9341,N_8559,N_8752);
nor U9342 (N_9342,N_8991,N_8648);
nor U9343 (N_9343,N_8811,N_8625);
and U9344 (N_9344,N_8584,N_8714);
and U9345 (N_9345,N_8529,N_8885);
nand U9346 (N_9346,N_8624,N_8844);
and U9347 (N_9347,N_8692,N_8827);
nand U9348 (N_9348,N_8586,N_8768);
and U9349 (N_9349,N_8561,N_8963);
nand U9350 (N_9350,N_8976,N_8900);
nand U9351 (N_9351,N_8603,N_8963);
nor U9352 (N_9352,N_8699,N_8724);
and U9353 (N_9353,N_8938,N_8804);
nand U9354 (N_9354,N_8719,N_8568);
or U9355 (N_9355,N_8532,N_8843);
or U9356 (N_9356,N_8578,N_8985);
nand U9357 (N_9357,N_8989,N_8707);
xor U9358 (N_9358,N_8558,N_8530);
or U9359 (N_9359,N_8939,N_8758);
or U9360 (N_9360,N_8979,N_8627);
and U9361 (N_9361,N_8520,N_8769);
nor U9362 (N_9362,N_8548,N_8896);
nor U9363 (N_9363,N_8875,N_8768);
nor U9364 (N_9364,N_8619,N_8799);
nand U9365 (N_9365,N_8516,N_8531);
nor U9366 (N_9366,N_8794,N_8886);
and U9367 (N_9367,N_8802,N_8523);
nor U9368 (N_9368,N_8842,N_8896);
and U9369 (N_9369,N_8567,N_8874);
nor U9370 (N_9370,N_8858,N_8661);
nor U9371 (N_9371,N_8559,N_8799);
nor U9372 (N_9372,N_8562,N_8709);
nor U9373 (N_9373,N_8569,N_8709);
nor U9374 (N_9374,N_8560,N_8664);
xor U9375 (N_9375,N_8502,N_8630);
nand U9376 (N_9376,N_8725,N_8951);
nor U9377 (N_9377,N_8570,N_8913);
nor U9378 (N_9378,N_8901,N_8778);
nor U9379 (N_9379,N_8879,N_8580);
nand U9380 (N_9380,N_8855,N_8728);
nor U9381 (N_9381,N_8722,N_8647);
nand U9382 (N_9382,N_8569,N_8809);
or U9383 (N_9383,N_8992,N_8957);
or U9384 (N_9384,N_8885,N_8811);
nor U9385 (N_9385,N_8896,N_8866);
or U9386 (N_9386,N_8889,N_8652);
nand U9387 (N_9387,N_8607,N_8998);
nor U9388 (N_9388,N_8779,N_8797);
nand U9389 (N_9389,N_8940,N_8578);
or U9390 (N_9390,N_8909,N_8877);
nor U9391 (N_9391,N_8582,N_8978);
or U9392 (N_9392,N_8783,N_8702);
nand U9393 (N_9393,N_8781,N_8778);
or U9394 (N_9394,N_8971,N_8621);
nand U9395 (N_9395,N_8889,N_8966);
or U9396 (N_9396,N_8567,N_8969);
xnor U9397 (N_9397,N_8986,N_8927);
xor U9398 (N_9398,N_8870,N_8855);
and U9399 (N_9399,N_8667,N_8715);
nand U9400 (N_9400,N_8507,N_8840);
or U9401 (N_9401,N_8501,N_8675);
nand U9402 (N_9402,N_8641,N_8844);
nor U9403 (N_9403,N_8846,N_8721);
xnor U9404 (N_9404,N_8618,N_8611);
and U9405 (N_9405,N_8804,N_8829);
nand U9406 (N_9406,N_8506,N_8919);
or U9407 (N_9407,N_8571,N_8702);
xnor U9408 (N_9408,N_8739,N_8549);
or U9409 (N_9409,N_8884,N_8957);
and U9410 (N_9410,N_8977,N_8711);
nand U9411 (N_9411,N_8592,N_8611);
or U9412 (N_9412,N_8721,N_8637);
or U9413 (N_9413,N_8854,N_8567);
and U9414 (N_9414,N_8621,N_8862);
or U9415 (N_9415,N_8765,N_8866);
or U9416 (N_9416,N_8737,N_8642);
nand U9417 (N_9417,N_8874,N_8798);
xnor U9418 (N_9418,N_8968,N_8935);
and U9419 (N_9419,N_8634,N_8736);
or U9420 (N_9420,N_8833,N_8984);
xnor U9421 (N_9421,N_8593,N_8545);
nand U9422 (N_9422,N_8945,N_8825);
and U9423 (N_9423,N_8654,N_8811);
xor U9424 (N_9424,N_8915,N_8677);
nor U9425 (N_9425,N_8671,N_8523);
xnor U9426 (N_9426,N_8569,N_8746);
or U9427 (N_9427,N_8785,N_8974);
nand U9428 (N_9428,N_8760,N_8886);
nand U9429 (N_9429,N_8736,N_8783);
xor U9430 (N_9430,N_8570,N_8881);
and U9431 (N_9431,N_8772,N_8752);
or U9432 (N_9432,N_8668,N_8566);
and U9433 (N_9433,N_8662,N_8813);
or U9434 (N_9434,N_8690,N_8817);
or U9435 (N_9435,N_8659,N_8574);
nand U9436 (N_9436,N_8610,N_8894);
nor U9437 (N_9437,N_8783,N_8514);
or U9438 (N_9438,N_8947,N_8983);
or U9439 (N_9439,N_8902,N_8610);
nand U9440 (N_9440,N_8959,N_8967);
nor U9441 (N_9441,N_8562,N_8578);
or U9442 (N_9442,N_8846,N_8601);
xor U9443 (N_9443,N_8546,N_8900);
and U9444 (N_9444,N_8538,N_8872);
and U9445 (N_9445,N_8997,N_8946);
nand U9446 (N_9446,N_8966,N_8847);
xor U9447 (N_9447,N_8755,N_8922);
nand U9448 (N_9448,N_8863,N_8574);
and U9449 (N_9449,N_8750,N_8876);
and U9450 (N_9450,N_8604,N_8628);
nand U9451 (N_9451,N_8564,N_8810);
xnor U9452 (N_9452,N_8671,N_8921);
xnor U9453 (N_9453,N_8846,N_8805);
or U9454 (N_9454,N_8770,N_8861);
nand U9455 (N_9455,N_8628,N_8814);
nand U9456 (N_9456,N_8857,N_8587);
nor U9457 (N_9457,N_8891,N_8677);
nand U9458 (N_9458,N_8668,N_8689);
nor U9459 (N_9459,N_8829,N_8510);
or U9460 (N_9460,N_8605,N_8622);
or U9461 (N_9461,N_8672,N_8925);
and U9462 (N_9462,N_8526,N_8865);
and U9463 (N_9463,N_8592,N_8665);
and U9464 (N_9464,N_8542,N_8658);
nand U9465 (N_9465,N_8644,N_8747);
nand U9466 (N_9466,N_8967,N_8792);
nor U9467 (N_9467,N_8777,N_8500);
nand U9468 (N_9468,N_8710,N_8961);
xor U9469 (N_9469,N_8957,N_8805);
and U9470 (N_9470,N_8983,N_8603);
nand U9471 (N_9471,N_8974,N_8506);
and U9472 (N_9472,N_8702,N_8962);
or U9473 (N_9473,N_8786,N_8972);
and U9474 (N_9474,N_8681,N_8965);
or U9475 (N_9475,N_8571,N_8716);
nand U9476 (N_9476,N_8812,N_8742);
and U9477 (N_9477,N_8562,N_8502);
or U9478 (N_9478,N_8999,N_8759);
or U9479 (N_9479,N_8643,N_8850);
and U9480 (N_9480,N_8620,N_8892);
nand U9481 (N_9481,N_8585,N_8528);
nand U9482 (N_9482,N_8818,N_8940);
nor U9483 (N_9483,N_8944,N_8897);
nand U9484 (N_9484,N_8532,N_8589);
and U9485 (N_9485,N_8871,N_8873);
or U9486 (N_9486,N_8683,N_8902);
and U9487 (N_9487,N_8871,N_8789);
or U9488 (N_9488,N_8615,N_8900);
nor U9489 (N_9489,N_8883,N_8796);
xnor U9490 (N_9490,N_8684,N_8827);
nor U9491 (N_9491,N_8874,N_8805);
nand U9492 (N_9492,N_8779,N_8777);
nand U9493 (N_9493,N_8924,N_8624);
and U9494 (N_9494,N_8842,N_8501);
nor U9495 (N_9495,N_8670,N_8574);
nand U9496 (N_9496,N_8555,N_8893);
or U9497 (N_9497,N_8832,N_8906);
nor U9498 (N_9498,N_8620,N_8769);
and U9499 (N_9499,N_8556,N_8911);
and U9500 (N_9500,N_9044,N_9009);
nand U9501 (N_9501,N_9281,N_9033);
xnor U9502 (N_9502,N_9200,N_9302);
nor U9503 (N_9503,N_9499,N_9307);
nor U9504 (N_9504,N_9114,N_9139);
and U9505 (N_9505,N_9346,N_9251);
or U9506 (N_9506,N_9424,N_9075);
nor U9507 (N_9507,N_9154,N_9193);
nor U9508 (N_9508,N_9072,N_9460);
and U9509 (N_9509,N_9431,N_9481);
nor U9510 (N_9510,N_9282,N_9110);
nor U9511 (N_9511,N_9276,N_9048);
nand U9512 (N_9512,N_9096,N_9131);
or U9513 (N_9513,N_9464,N_9037);
and U9514 (N_9514,N_9190,N_9456);
nand U9515 (N_9515,N_9393,N_9268);
nor U9516 (N_9516,N_9375,N_9252);
nand U9517 (N_9517,N_9026,N_9250);
and U9518 (N_9518,N_9471,N_9201);
xnor U9519 (N_9519,N_9247,N_9449);
or U9520 (N_9520,N_9391,N_9183);
nor U9521 (N_9521,N_9034,N_9377);
nor U9522 (N_9522,N_9204,N_9416);
nor U9523 (N_9523,N_9434,N_9153);
nor U9524 (N_9524,N_9219,N_9477);
or U9525 (N_9525,N_9487,N_9148);
nor U9526 (N_9526,N_9236,N_9345);
nor U9527 (N_9527,N_9127,N_9203);
or U9528 (N_9528,N_9165,N_9334);
and U9529 (N_9529,N_9383,N_9237);
nand U9530 (N_9530,N_9270,N_9141);
and U9531 (N_9531,N_9397,N_9340);
nand U9532 (N_9532,N_9043,N_9001);
xnor U9533 (N_9533,N_9032,N_9476);
nand U9534 (N_9534,N_9292,N_9374);
and U9535 (N_9535,N_9233,N_9196);
nand U9536 (N_9536,N_9261,N_9197);
or U9537 (N_9537,N_9028,N_9243);
nor U9538 (N_9538,N_9145,N_9007);
nor U9539 (N_9539,N_9485,N_9064);
xnor U9540 (N_9540,N_9408,N_9163);
or U9541 (N_9541,N_9315,N_9494);
nand U9542 (N_9542,N_9318,N_9308);
or U9543 (N_9543,N_9419,N_9228);
or U9544 (N_9544,N_9128,N_9003);
nor U9545 (N_9545,N_9355,N_9194);
and U9546 (N_9546,N_9202,N_9150);
or U9547 (N_9547,N_9070,N_9327);
or U9548 (N_9548,N_9339,N_9267);
xnor U9549 (N_9549,N_9351,N_9293);
or U9550 (N_9550,N_9303,N_9239);
or U9551 (N_9551,N_9223,N_9294);
nor U9552 (N_9552,N_9211,N_9323);
nor U9553 (N_9553,N_9452,N_9160);
xnor U9554 (N_9554,N_9002,N_9467);
nand U9555 (N_9555,N_9184,N_9210);
and U9556 (N_9556,N_9269,N_9212);
nand U9557 (N_9557,N_9395,N_9229);
and U9558 (N_9558,N_9429,N_9112);
xnor U9559 (N_9559,N_9142,N_9344);
nand U9560 (N_9560,N_9102,N_9284);
nor U9561 (N_9561,N_9135,N_9271);
or U9562 (N_9562,N_9017,N_9177);
and U9563 (N_9563,N_9496,N_9086);
and U9564 (N_9564,N_9483,N_9093);
and U9565 (N_9565,N_9046,N_9491);
and U9566 (N_9566,N_9192,N_9301);
nand U9567 (N_9567,N_9011,N_9451);
nor U9568 (N_9568,N_9242,N_9309);
nor U9569 (N_9569,N_9446,N_9062);
nor U9570 (N_9570,N_9372,N_9101);
nand U9571 (N_9571,N_9328,N_9061);
and U9572 (N_9572,N_9480,N_9295);
nor U9573 (N_9573,N_9352,N_9258);
xnor U9574 (N_9574,N_9156,N_9079);
and U9575 (N_9575,N_9240,N_9207);
or U9576 (N_9576,N_9018,N_9461);
and U9577 (N_9577,N_9423,N_9470);
or U9578 (N_9578,N_9151,N_9117);
and U9579 (N_9579,N_9244,N_9306);
or U9580 (N_9580,N_9299,N_9472);
nand U9581 (N_9581,N_9359,N_9132);
and U9582 (N_9582,N_9362,N_9364);
nand U9583 (N_9583,N_9254,N_9035);
xor U9584 (N_9584,N_9067,N_9134);
nand U9585 (N_9585,N_9298,N_9126);
nand U9586 (N_9586,N_9417,N_9222);
and U9587 (N_9587,N_9332,N_9158);
or U9588 (N_9588,N_9052,N_9189);
and U9589 (N_9589,N_9272,N_9418);
or U9590 (N_9590,N_9389,N_9369);
and U9591 (N_9591,N_9444,N_9263);
nand U9592 (N_9592,N_9209,N_9342);
and U9593 (N_9593,N_9278,N_9232);
or U9594 (N_9594,N_9162,N_9285);
and U9595 (N_9595,N_9199,N_9103);
and U9596 (N_9596,N_9166,N_9071);
nor U9597 (N_9597,N_9104,N_9379);
and U9598 (N_9598,N_9113,N_9404);
nor U9599 (N_9599,N_9358,N_9171);
nand U9600 (N_9600,N_9231,N_9310);
and U9601 (N_9601,N_9325,N_9498);
and U9602 (N_9602,N_9347,N_9300);
nand U9603 (N_9603,N_9195,N_9324);
or U9604 (N_9604,N_9257,N_9394);
or U9605 (N_9605,N_9349,N_9279);
and U9606 (N_9606,N_9405,N_9290);
and U9607 (N_9607,N_9403,N_9462);
nand U9608 (N_9608,N_9187,N_9024);
or U9609 (N_9609,N_9454,N_9466);
nor U9610 (N_9610,N_9036,N_9433);
and U9611 (N_9611,N_9450,N_9140);
and U9612 (N_9612,N_9225,N_9085);
or U9613 (N_9613,N_9100,N_9245);
and U9614 (N_9614,N_9121,N_9060);
nand U9615 (N_9615,N_9387,N_9287);
nor U9616 (N_9616,N_9410,N_9057);
nor U9617 (N_9617,N_9084,N_9095);
nor U9618 (N_9618,N_9343,N_9421);
or U9619 (N_9619,N_9384,N_9008);
nand U9620 (N_9620,N_9123,N_9159);
and U9621 (N_9621,N_9049,N_9216);
nand U9622 (N_9622,N_9092,N_9053);
and U9623 (N_9623,N_9333,N_9320);
nand U9624 (N_9624,N_9442,N_9412);
and U9625 (N_9625,N_9164,N_9068);
or U9626 (N_9626,N_9365,N_9356);
and U9627 (N_9627,N_9174,N_9275);
nor U9628 (N_9628,N_9492,N_9063);
nor U9629 (N_9629,N_9178,N_9413);
nor U9630 (N_9630,N_9118,N_9181);
and U9631 (N_9631,N_9371,N_9213);
nand U9632 (N_9632,N_9425,N_9437);
nand U9633 (N_9633,N_9330,N_9169);
or U9634 (N_9634,N_9042,N_9221);
or U9635 (N_9635,N_9055,N_9090);
nor U9636 (N_9636,N_9406,N_9399);
and U9637 (N_9637,N_9482,N_9291);
and U9638 (N_9638,N_9208,N_9056);
nor U9639 (N_9639,N_9381,N_9361);
xor U9640 (N_9640,N_9445,N_9255);
xnor U9641 (N_9641,N_9441,N_9326);
and U9642 (N_9642,N_9014,N_9360);
xor U9643 (N_9643,N_9206,N_9402);
nor U9644 (N_9644,N_9137,N_9463);
nor U9645 (N_9645,N_9266,N_9478);
nand U9646 (N_9646,N_9493,N_9115);
nor U9647 (N_9647,N_9336,N_9474);
and U9648 (N_9648,N_9317,N_9396);
or U9649 (N_9649,N_9180,N_9378);
and U9650 (N_9650,N_9296,N_9021);
and U9651 (N_9651,N_9373,N_9099);
or U9652 (N_9652,N_9138,N_9168);
and U9653 (N_9653,N_9186,N_9338);
or U9654 (N_9654,N_9205,N_9078);
or U9655 (N_9655,N_9319,N_9265);
or U9656 (N_9656,N_9022,N_9227);
nor U9657 (N_9657,N_9226,N_9077);
and U9658 (N_9658,N_9447,N_9286);
or U9659 (N_9659,N_9337,N_9312);
and U9660 (N_9660,N_9191,N_9149);
xor U9661 (N_9661,N_9106,N_9124);
nand U9662 (N_9662,N_9439,N_9039);
or U9663 (N_9663,N_9422,N_9025);
and U9664 (N_9664,N_9031,N_9217);
nand U9665 (N_9665,N_9047,N_9288);
and U9666 (N_9666,N_9479,N_9004);
or U9667 (N_9667,N_9438,N_9176);
and U9668 (N_9668,N_9074,N_9069);
and U9669 (N_9669,N_9440,N_9430);
or U9670 (N_9670,N_9277,N_9392);
nand U9671 (N_9671,N_9054,N_9260);
and U9672 (N_9672,N_9458,N_9133);
or U9673 (N_9673,N_9019,N_9157);
xor U9674 (N_9674,N_9185,N_9311);
xor U9675 (N_9675,N_9170,N_9427);
nand U9676 (N_9676,N_9420,N_9367);
and U9677 (N_9677,N_9220,N_9182);
nor U9678 (N_9678,N_9144,N_9407);
and U9679 (N_9679,N_9188,N_9256);
xnor U9680 (N_9680,N_9146,N_9322);
nor U9681 (N_9681,N_9076,N_9348);
or U9682 (N_9682,N_9366,N_9283);
nand U9683 (N_9683,N_9111,N_9475);
or U9684 (N_9684,N_9274,N_9262);
or U9685 (N_9685,N_9030,N_9119);
and U9686 (N_9686,N_9058,N_9414);
nand U9687 (N_9687,N_9313,N_9214);
and U9688 (N_9688,N_9167,N_9050);
nor U9689 (N_9689,N_9125,N_9426);
xnor U9690 (N_9690,N_9495,N_9108);
nand U9691 (N_9691,N_9215,N_9297);
nand U9692 (N_9692,N_9235,N_9273);
nand U9693 (N_9693,N_9136,N_9341);
or U9694 (N_9694,N_9155,N_9013);
or U9695 (N_9695,N_9038,N_9304);
nor U9696 (N_9696,N_9143,N_9289);
or U9697 (N_9697,N_9027,N_9314);
and U9698 (N_9698,N_9073,N_9172);
xnor U9699 (N_9699,N_9249,N_9241);
nor U9700 (N_9700,N_9329,N_9147);
and U9701 (N_9701,N_9059,N_9122);
or U9702 (N_9702,N_9457,N_9370);
or U9703 (N_9703,N_9094,N_9097);
and U9704 (N_9704,N_9488,N_9246);
xnor U9705 (N_9705,N_9029,N_9224);
and U9706 (N_9706,N_9468,N_9040);
nand U9707 (N_9707,N_9321,N_9259);
nor U9708 (N_9708,N_9116,N_9489);
and U9709 (N_9709,N_9152,N_9305);
nor U9710 (N_9710,N_9015,N_9051);
nand U9711 (N_9711,N_9486,N_9473);
nand U9712 (N_9712,N_9428,N_9091);
nand U9713 (N_9713,N_9218,N_9382);
nand U9714 (N_9714,N_9253,N_9080);
nand U9715 (N_9715,N_9436,N_9198);
xnor U9716 (N_9716,N_9083,N_9000);
nor U9717 (N_9717,N_9082,N_9497);
nand U9718 (N_9718,N_9087,N_9088);
and U9719 (N_9719,N_9005,N_9129);
nand U9720 (N_9720,N_9175,N_9443);
or U9721 (N_9721,N_9012,N_9484);
and U9722 (N_9722,N_9105,N_9130);
nor U9723 (N_9723,N_9459,N_9435);
nor U9724 (N_9724,N_9161,N_9264);
and U9725 (N_9725,N_9066,N_9006);
nor U9726 (N_9726,N_9385,N_9109);
and U9727 (N_9727,N_9081,N_9173);
nand U9728 (N_9728,N_9388,N_9120);
and U9729 (N_9729,N_9353,N_9230);
and U9730 (N_9730,N_9248,N_9401);
nor U9731 (N_9731,N_9400,N_9354);
nand U9732 (N_9732,N_9415,N_9380);
and U9733 (N_9733,N_9010,N_9107);
nor U9734 (N_9734,N_9179,N_9363);
and U9735 (N_9735,N_9453,N_9386);
nand U9736 (N_9736,N_9023,N_9016);
nor U9737 (N_9737,N_9469,N_9350);
and U9738 (N_9738,N_9234,N_9335);
nand U9739 (N_9739,N_9280,N_9357);
nand U9740 (N_9740,N_9411,N_9390);
and U9741 (N_9741,N_9490,N_9316);
nor U9742 (N_9742,N_9098,N_9020);
or U9743 (N_9743,N_9331,N_9238);
nor U9744 (N_9744,N_9448,N_9376);
xnor U9745 (N_9745,N_9065,N_9465);
or U9746 (N_9746,N_9432,N_9398);
nor U9747 (N_9747,N_9089,N_9368);
xor U9748 (N_9748,N_9045,N_9455);
or U9749 (N_9749,N_9409,N_9041);
or U9750 (N_9750,N_9379,N_9019);
or U9751 (N_9751,N_9267,N_9026);
nor U9752 (N_9752,N_9032,N_9481);
and U9753 (N_9753,N_9222,N_9362);
nor U9754 (N_9754,N_9355,N_9204);
or U9755 (N_9755,N_9481,N_9171);
nor U9756 (N_9756,N_9284,N_9271);
and U9757 (N_9757,N_9139,N_9296);
and U9758 (N_9758,N_9094,N_9203);
nor U9759 (N_9759,N_9348,N_9454);
nor U9760 (N_9760,N_9073,N_9316);
nand U9761 (N_9761,N_9000,N_9362);
nor U9762 (N_9762,N_9396,N_9046);
nand U9763 (N_9763,N_9040,N_9318);
xnor U9764 (N_9764,N_9326,N_9257);
and U9765 (N_9765,N_9307,N_9002);
xnor U9766 (N_9766,N_9421,N_9449);
xnor U9767 (N_9767,N_9231,N_9068);
nor U9768 (N_9768,N_9394,N_9377);
or U9769 (N_9769,N_9139,N_9037);
nor U9770 (N_9770,N_9411,N_9143);
nor U9771 (N_9771,N_9331,N_9398);
nor U9772 (N_9772,N_9283,N_9001);
nand U9773 (N_9773,N_9255,N_9345);
or U9774 (N_9774,N_9116,N_9183);
nor U9775 (N_9775,N_9228,N_9262);
or U9776 (N_9776,N_9421,N_9194);
nor U9777 (N_9777,N_9172,N_9275);
or U9778 (N_9778,N_9114,N_9045);
nand U9779 (N_9779,N_9163,N_9153);
nand U9780 (N_9780,N_9178,N_9005);
and U9781 (N_9781,N_9094,N_9181);
nand U9782 (N_9782,N_9001,N_9377);
nand U9783 (N_9783,N_9081,N_9470);
and U9784 (N_9784,N_9128,N_9111);
nor U9785 (N_9785,N_9441,N_9005);
nand U9786 (N_9786,N_9499,N_9441);
nand U9787 (N_9787,N_9168,N_9055);
and U9788 (N_9788,N_9039,N_9124);
and U9789 (N_9789,N_9320,N_9048);
and U9790 (N_9790,N_9199,N_9247);
nand U9791 (N_9791,N_9040,N_9313);
nand U9792 (N_9792,N_9389,N_9348);
and U9793 (N_9793,N_9488,N_9170);
or U9794 (N_9794,N_9435,N_9253);
and U9795 (N_9795,N_9497,N_9389);
nand U9796 (N_9796,N_9269,N_9428);
and U9797 (N_9797,N_9324,N_9161);
xor U9798 (N_9798,N_9493,N_9262);
nand U9799 (N_9799,N_9016,N_9127);
nand U9800 (N_9800,N_9470,N_9116);
nand U9801 (N_9801,N_9484,N_9035);
nand U9802 (N_9802,N_9349,N_9343);
nor U9803 (N_9803,N_9133,N_9244);
nor U9804 (N_9804,N_9356,N_9241);
and U9805 (N_9805,N_9469,N_9172);
or U9806 (N_9806,N_9200,N_9395);
nor U9807 (N_9807,N_9463,N_9433);
nor U9808 (N_9808,N_9456,N_9245);
or U9809 (N_9809,N_9148,N_9322);
xnor U9810 (N_9810,N_9119,N_9292);
and U9811 (N_9811,N_9114,N_9212);
and U9812 (N_9812,N_9471,N_9163);
nand U9813 (N_9813,N_9294,N_9052);
nand U9814 (N_9814,N_9483,N_9466);
nor U9815 (N_9815,N_9481,N_9094);
nor U9816 (N_9816,N_9274,N_9401);
nor U9817 (N_9817,N_9410,N_9331);
nand U9818 (N_9818,N_9058,N_9015);
nand U9819 (N_9819,N_9018,N_9390);
nor U9820 (N_9820,N_9050,N_9152);
xor U9821 (N_9821,N_9487,N_9186);
or U9822 (N_9822,N_9141,N_9139);
and U9823 (N_9823,N_9223,N_9387);
or U9824 (N_9824,N_9120,N_9289);
and U9825 (N_9825,N_9338,N_9046);
or U9826 (N_9826,N_9336,N_9162);
or U9827 (N_9827,N_9227,N_9319);
nor U9828 (N_9828,N_9234,N_9356);
nor U9829 (N_9829,N_9058,N_9176);
and U9830 (N_9830,N_9409,N_9228);
nor U9831 (N_9831,N_9325,N_9423);
or U9832 (N_9832,N_9213,N_9429);
xor U9833 (N_9833,N_9207,N_9433);
nor U9834 (N_9834,N_9236,N_9470);
nor U9835 (N_9835,N_9034,N_9357);
xor U9836 (N_9836,N_9448,N_9355);
nor U9837 (N_9837,N_9053,N_9081);
nand U9838 (N_9838,N_9435,N_9369);
nor U9839 (N_9839,N_9472,N_9139);
or U9840 (N_9840,N_9338,N_9453);
xnor U9841 (N_9841,N_9488,N_9126);
and U9842 (N_9842,N_9448,N_9149);
and U9843 (N_9843,N_9003,N_9373);
nand U9844 (N_9844,N_9389,N_9214);
nor U9845 (N_9845,N_9415,N_9046);
nor U9846 (N_9846,N_9476,N_9202);
xor U9847 (N_9847,N_9340,N_9339);
nand U9848 (N_9848,N_9399,N_9194);
xor U9849 (N_9849,N_9019,N_9015);
and U9850 (N_9850,N_9274,N_9318);
or U9851 (N_9851,N_9044,N_9005);
nor U9852 (N_9852,N_9128,N_9118);
nor U9853 (N_9853,N_9075,N_9357);
or U9854 (N_9854,N_9333,N_9136);
nand U9855 (N_9855,N_9141,N_9275);
xor U9856 (N_9856,N_9324,N_9213);
nand U9857 (N_9857,N_9185,N_9280);
nor U9858 (N_9858,N_9308,N_9206);
or U9859 (N_9859,N_9311,N_9187);
nand U9860 (N_9860,N_9019,N_9156);
nor U9861 (N_9861,N_9018,N_9255);
nand U9862 (N_9862,N_9285,N_9153);
or U9863 (N_9863,N_9036,N_9374);
nand U9864 (N_9864,N_9171,N_9002);
nor U9865 (N_9865,N_9330,N_9005);
and U9866 (N_9866,N_9190,N_9284);
nand U9867 (N_9867,N_9306,N_9293);
nor U9868 (N_9868,N_9443,N_9196);
or U9869 (N_9869,N_9205,N_9363);
nor U9870 (N_9870,N_9241,N_9424);
nor U9871 (N_9871,N_9259,N_9287);
and U9872 (N_9872,N_9273,N_9060);
and U9873 (N_9873,N_9310,N_9108);
and U9874 (N_9874,N_9115,N_9467);
or U9875 (N_9875,N_9402,N_9234);
nor U9876 (N_9876,N_9431,N_9281);
nand U9877 (N_9877,N_9011,N_9278);
or U9878 (N_9878,N_9296,N_9450);
or U9879 (N_9879,N_9051,N_9080);
nand U9880 (N_9880,N_9087,N_9396);
nor U9881 (N_9881,N_9384,N_9106);
nand U9882 (N_9882,N_9270,N_9205);
nand U9883 (N_9883,N_9430,N_9246);
nand U9884 (N_9884,N_9316,N_9301);
nor U9885 (N_9885,N_9351,N_9200);
and U9886 (N_9886,N_9201,N_9216);
nand U9887 (N_9887,N_9299,N_9040);
nor U9888 (N_9888,N_9056,N_9097);
or U9889 (N_9889,N_9078,N_9397);
nand U9890 (N_9890,N_9437,N_9174);
or U9891 (N_9891,N_9170,N_9372);
nor U9892 (N_9892,N_9017,N_9203);
nor U9893 (N_9893,N_9448,N_9205);
and U9894 (N_9894,N_9419,N_9402);
or U9895 (N_9895,N_9004,N_9117);
nor U9896 (N_9896,N_9282,N_9041);
nand U9897 (N_9897,N_9268,N_9367);
or U9898 (N_9898,N_9214,N_9085);
nand U9899 (N_9899,N_9015,N_9228);
or U9900 (N_9900,N_9309,N_9143);
and U9901 (N_9901,N_9189,N_9370);
and U9902 (N_9902,N_9413,N_9258);
or U9903 (N_9903,N_9380,N_9411);
nand U9904 (N_9904,N_9294,N_9330);
or U9905 (N_9905,N_9433,N_9055);
and U9906 (N_9906,N_9049,N_9057);
nand U9907 (N_9907,N_9350,N_9251);
xnor U9908 (N_9908,N_9386,N_9423);
nor U9909 (N_9909,N_9374,N_9149);
nand U9910 (N_9910,N_9004,N_9470);
xor U9911 (N_9911,N_9482,N_9457);
and U9912 (N_9912,N_9072,N_9412);
nor U9913 (N_9913,N_9399,N_9035);
and U9914 (N_9914,N_9266,N_9279);
nor U9915 (N_9915,N_9019,N_9283);
nor U9916 (N_9916,N_9485,N_9454);
nand U9917 (N_9917,N_9481,N_9293);
and U9918 (N_9918,N_9134,N_9331);
and U9919 (N_9919,N_9187,N_9419);
nand U9920 (N_9920,N_9169,N_9336);
and U9921 (N_9921,N_9369,N_9283);
nor U9922 (N_9922,N_9328,N_9376);
nand U9923 (N_9923,N_9375,N_9236);
and U9924 (N_9924,N_9030,N_9113);
nand U9925 (N_9925,N_9391,N_9027);
nor U9926 (N_9926,N_9338,N_9009);
and U9927 (N_9927,N_9438,N_9246);
nor U9928 (N_9928,N_9005,N_9248);
and U9929 (N_9929,N_9288,N_9057);
or U9930 (N_9930,N_9224,N_9379);
nand U9931 (N_9931,N_9494,N_9263);
and U9932 (N_9932,N_9056,N_9403);
or U9933 (N_9933,N_9321,N_9283);
or U9934 (N_9934,N_9382,N_9120);
xor U9935 (N_9935,N_9004,N_9073);
or U9936 (N_9936,N_9242,N_9046);
and U9937 (N_9937,N_9102,N_9013);
or U9938 (N_9938,N_9384,N_9118);
xor U9939 (N_9939,N_9025,N_9185);
nand U9940 (N_9940,N_9035,N_9483);
or U9941 (N_9941,N_9386,N_9483);
or U9942 (N_9942,N_9083,N_9182);
or U9943 (N_9943,N_9376,N_9280);
and U9944 (N_9944,N_9391,N_9194);
nor U9945 (N_9945,N_9442,N_9124);
nor U9946 (N_9946,N_9227,N_9049);
and U9947 (N_9947,N_9148,N_9467);
nor U9948 (N_9948,N_9233,N_9095);
or U9949 (N_9949,N_9079,N_9132);
nand U9950 (N_9950,N_9407,N_9107);
xnor U9951 (N_9951,N_9240,N_9123);
nor U9952 (N_9952,N_9397,N_9034);
or U9953 (N_9953,N_9294,N_9029);
or U9954 (N_9954,N_9019,N_9086);
or U9955 (N_9955,N_9387,N_9426);
nor U9956 (N_9956,N_9015,N_9417);
and U9957 (N_9957,N_9387,N_9190);
nor U9958 (N_9958,N_9169,N_9180);
nor U9959 (N_9959,N_9051,N_9103);
or U9960 (N_9960,N_9138,N_9162);
nor U9961 (N_9961,N_9277,N_9139);
and U9962 (N_9962,N_9189,N_9272);
and U9963 (N_9963,N_9042,N_9440);
and U9964 (N_9964,N_9378,N_9245);
nor U9965 (N_9965,N_9304,N_9041);
and U9966 (N_9966,N_9124,N_9009);
and U9967 (N_9967,N_9260,N_9331);
nand U9968 (N_9968,N_9489,N_9255);
nor U9969 (N_9969,N_9009,N_9347);
xnor U9970 (N_9970,N_9282,N_9022);
xnor U9971 (N_9971,N_9089,N_9341);
nor U9972 (N_9972,N_9090,N_9479);
nand U9973 (N_9973,N_9366,N_9088);
nor U9974 (N_9974,N_9173,N_9339);
nor U9975 (N_9975,N_9208,N_9105);
nand U9976 (N_9976,N_9430,N_9462);
and U9977 (N_9977,N_9432,N_9325);
nor U9978 (N_9978,N_9189,N_9150);
xnor U9979 (N_9979,N_9469,N_9007);
or U9980 (N_9980,N_9340,N_9484);
nor U9981 (N_9981,N_9035,N_9032);
nand U9982 (N_9982,N_9358,N_9157);
and U9983 (N_9983,N_9225,N_9000);
xnor U9984 (N_9984,N_9275,N_9051);
and U9985 (N_9985,N_9134,N_9447);
or U9986 (N_9986,N_9211,N_9053);
nand U9987 (N_9987,N_9189,N_9051);
and U9988 (N_9988,N_9264,N_9168);
or U9989 (N_9989,N_9308,N_9358);
nand U9990 (N_9990,N_9348,N_9267);
and U9991 (N_9991,N_9447,N_9168);
xnor U9992 (N_9992,N_9039,N_9480);
nand U9993 (N_9993,N_9334,N_9250);
nand U9994 (N_9994,N_9425,N_9443);
and U9995 (N_9995,N_9427,N_9402);
or U9996 (N_9996,N_9337,N_9150);
and U9997 (N_9997,N_9129,N_9359);
xnor U9998 (N_9998,N_9011,N_9267);
nand U9999 (N_9999,N_9355,N_9450);
xnor UO_0 (O_0,N_9872,N_9514);
xnor UO_1 (O_1,N_9586,N_9766);
or UO_2 (O_2,N_9581,N_9575);
nand UO_3 (O_3,N_9897,N_9844);
nand UO_4 (O_4,N_9672,N_9749);
nor UO_5 (O_5,N_9772,N_9989);
or UO_6 (O_6,N_9781,N_9795);
nor UO_7 (O_7,N_9674,N_9942);
or UO_8 (O_8,N_9995,N_9652);
and UO_9 (O_9,N_9682,N_9697);
and UO_10 (O_10,N_9861,N_9667);
or UO_11 (O_11,N_9547,N_9822);
nand UO_12 (O_12,N_9912,N_9585);
and UO_13 (O_13,N_9531,N_9792);
nand UO_14 (O_14,N_9618,N_9933);
and UO_15 (O_15,N_9638,N_9837);
or UO_16 (O_16,N_9563,N_9768);
or UO_17 (O_17,N_9759,N_9883);
nor UO_18 (O_18,N_9594,N_9946);
nand UO_19 (O_19,N_9587,N_9863);
or UO_20 (O_20,N_9911,N_9501);
and UO_21 (O_21,N_9906,N_9655);
nor UO_22 (O_22,N_9903,N_9802);
and UO_23 (O_23,N_9633,N_9976);
nand UO_24 (O_24,N_9612,N_9789);
nand UO_25 (O_25,N_9829,N_9687);
or UO_26 (O_26,N_9816,N_9647);
or UO_27 (O_27,N_9967,N_9701);
and UO_28 (O_28,N_9523,N_9584);
nor UO_29 (O_29,N_9666,N_9710);
and UO_30 (O_30,N_9824,N_9814);
and UO_31 (O_31,N_9509,N_9573);
nand UO_32 (O_32,N_9916,N_9922);
nand UO_33 (O_33,N_9656,N_9538);
nand UO_34 (O_34,N_9699,N_9893);
xor UO_35 (O_35,N_9676,N_9619);
nand UO_36 (O_36,N_9705,N_9843);
and UO_37 (O_37,N_9924,N_9854);
and UO_38 (O_38,N_9606,N_9935);
or UO_39 (O_39,N_9921,N_9529);
and UO_40 (O_40,N_9970,N_9838);
nand UO_41 (O_41,N_9600,N_9831);
or UO_42 (O_42,N_9777,N_9929);
or UO_43 (O_43,N_9823,N_9557);
nand UO_44 (O_44,N_9537,N_9566);
nor UO_45 (O_45,N_9974,N_9668);
nand UO_46 (O_46,N_9930,N_9971);
and UO_47 (O_47,N_9920,N_9728);
or UO_48 (O_48,N_9830,N_9966);
nand UO_49 (O_49,N_9570,N_9712);
nand UO_50 (O_50,N_9720,N_9568);
nand UO_51 (O_51,N_9702,N_9528);
nand UO_52 (O_52,N_9640,N_9776);
and UO_53 (O_53,N_9960,N_9887);
nand UO_54 (O_54,N_9654,N_9956);
nor UO_55 (O_55,N_9669,N_9534);
nor UO_56 (O_56,N_9583,N_9630);
nor UO_57 (O_57,N_9907,N_9909);
nor UO_58 (O_58,N_9622,N_9972);
nor UO_59 (O_59,N_9836,N_9686);
nand UO_60 (O_60,N_9646,N_9740);
and UO_61 (O_61,N_9842,N_9592);
xnor UO_62 (O_62,N_9992,N_9828);
nor UO_63 (O_63,N_9695,N_9516);
nor UO_64 (O_64,N_9550,N_9939);
nor UO_65 (O_65,N_9827,N_9614);
or UO_66 (O_66,N_9867,N_9671);
and UO_67 (O_67,N_9503,N_9886);
nor UO_68 (O_68,N_9898,N_9752);
nor UO_69 (O_69,N_9505,N_9554);
or UO_70 (O_70,N_9940,N_9582);
nand UO_71 (O_71,N_9821,N_9859);
or UO_72 (O_72,N_9748,N_9965);
or UO_73 (O_73,N_9603,N_9799);
xor UO_74 (O_74,N_9739,N_9810);
xnor UO_75 (O_75,N_9502,N_9951);
nand UO_76 (O_76,N_9657,N_9663);
nand UO_77 (O_77,N_9724,N_9678);
nor UO_78 (O_78,N_9910,N_9524);
and UO_79 (O_79,N_9977,N_9665);
or UO_80 (O_80,N_9741,N_9987);
and UO_81 (O_81,N_9527,N_9609);
nand UO_82 (O_82,N_9913,N_9934);
and UO_83 (O_83,N_9707,N_9990);
xnor UO_84 (O_84,N_9545,N_9574);
and UO_85 (O_85,N_9706,N_9716);
nand UO_86 (O_86,N_9690,N_9508);
nand UO_87 (O_87,N_9525,N_9868);
nand UO_88 (O_88,N_9847,N_9954);
nand UO_89 (O_89,N_9878,N_9994);
and UO_90 (O_90,N_9653,N_9693);
or UO_91 (O_91,N_9778,N_9597);
and UO_92 (O_92,N_9708,N_9961);
or UO_93 (O_93,N_9700,N_9988);
nand UO_94 (O_94,N_9756,N_9753);
nand UO_95 (O_95,N_9698,N_9985);
nand UO_96 (O_96,N_9571,N_9876);
nand UO_97 (O_97,N_9993,N_9873);
nor UO_98 (O_98,N_9986,N_9797);
and UO_99 (O_99,N_9905,N_9670);
or UO_100 (O_100,N_9798,N_9629);
xor UO_101 (O_101,N_9635,N_9894);
nand UO_102 (O_102,N_9780,N_9659);
nand UO_103 (O_103,N_9813,N_9532);
or UO_104 (O_104,N_9628,N_9714);
or UO_105 (O_105,N_9950,N_9561);
or UO_106 (O_106,N_9602,N_9808);
nand UO_107 (O_107,N_9504,N_9978);
nand UO_108 (O_108,N_9650,N_9998);
nand UO_109 (O_109,N_9641,N_9945);
nor UO_110 (O_110,N_9996,N_9809);
nand UO_111 (O_111,N_9806,N_9895);
or UO_112 (O_112,N_9569,N_9560);
and UO_113 (O_113,N_9729,N_9825);
and UO_114 (O_114,N_9599,N_9999);
xnor UO_115 (O_115,N_9851,N_9757);
nand UO_116 (O_116,N_9888,N_9555);
nand UO_117 (O_117,N_9937,N_9725);
and UO_118 (O_118,N_9746,N_9984);
or UO_119 (O_119,N_9535,N_9662);
nor UO_120 (O_120,N_9673,N_9551);
nand UO_121 (O_121,N_9846,N_9623);
nand UO_122 (O_122,N_9848,N_9621);
and UO_123 (O_123,N_9896,N_9925);
and UO_124 (O_124,N_9579,N_9926);
nand UO_125 (O_125,N_9533,N_9747);
or UO_126 (O_126,N_9860,N_9723);
or UO_127 (O_127,N_9730,N_9593);
nor UO_128 (O_128,N_9608,N_9796);
and UO_129 (O_129,N_9879,N_9811);
or UO_130 (O_130,N_9677,N_9648);
nand UO_131 (O_131,N_9691,N_9625);
nor UO_132 (O_132,N_9807,N_9949);
or UO_133 (O_133,N_9639,N_9783);
nor UO_134 (O_134,N_9862,N_9649);
or UO_135 (O_135,N_9882,N_9855);
nand UO_136 (O_136,N_9578,N_9884);
nor UO_137 (O_137,N_9959,N_9856);
or UO_138 (O_138,N_9680,N_9745);
and UO_139 (O_139,N_9644,N_9694);
xor UO_140 (O_140,N_9890,N_9773);
nand UO_141 (O_141,N_9704,N_9803);
nand UO_142 (O_142,N_9834,N_9715);
nand UO_143 (O_143,N_9519,N_9590);
nand UO_144 (O_144,N_9565,N_9785);
or UO_145 (O_145,N_9958,N_9932);
xor UO_146 (O_146,N_9923,N_9761);
nand UO_147 (O_147,N_9900,N_9791);
and UO_148 (O_148,N_9679,N_9651);
or UO_149 (O_149,N_9731,N_9553);
and UO_150 (O_150,N_9727,N_9526);
or UO_151 (O_151,N_9709,N_9908);
or UO_152 (O_152,N_9564,N_9786);
xor UO_153 (O_153,N_9904,N_9952);
xor UO_154 (O_154,N_9589,N_9871);
and UO_155 (O_155,N_9763,N_9964);
and UO_156 (O_156,N_9675,N_9562);
and UO_157 (O_157,N_9507,N_9760);
and UO_158 (O_158,N_9552,N_9610);
nor UO_159 (O_159,N_9917,N_9634);
and UO_160 (O_160,N_9758,N_9853);
nor UO_161 (O_161,N_9626,N_9643);
nor UO_162 (O_162,N_9751,N_9518);
xor UO_163 (O_163,N_9901,N_9632);
nor UO_164 (O_164,N_9559,N_9767);
xor UO_165 (O_165,N_9953,N_9688);
nand UO_166 (O_166,N_9591,N_9931);
nor UO_167 (O_167,N_9735,N_9975);
nand UO_168 (O_168,N_9963,N_9510);
nand UO_169 (O_169,N_9750,N_9820);
or UO_170 (O_170,N_9755,N_9849);
nand UO_171 (O_171,N_9793,N_9616);
or UO_172 (O_172,N_9733,N_9536);
or UO_173 (O_173,N_9637,N_9962);
nor UO_174 (O_174,N_9892,N_9541);
and UO_175 (O_175,N_9779,N_9736);
and UO_176 (O_176,N_9889,N_9815);
nand UO_177 (O_177,N_9968,N_9515);
or UO_178 (O_178,N_9645,N_9875);
or UO_179 (O_179,N_9620,N_9684);
nor UO_180 (O_180,N_9734,N_9919);
nor UO_181 (O_181,N_9580,N_9784);
nor UO_182 (O_182,N_9558,N_9717);
or UO_183 (O_183,N_9611,N_9850);
nor UO_184 (O_184,N_9607,N_9754);
nor UO_185 (O_185,N_9549,N_9627);
nand UO_186 (O_186,N_9601,N_9774);
nor UO_187 (O_187,N_9718,N_9979);
nand UO_188 (O_188,N_9540,N_9790);
or UO_189 (O_189,N_9839,N_9530);
or UO_190 (O_190,N_9511,N_9969);
nand UO_191 (O_191,N_9744,N_9506);
or UO_192 (O_192,N_9770,N_9865);
nor UO_193 (O_193,N_9689,N_9835);
nor UO_194 (O_194,N_9983,N_9845);
nand UO_195 (O_195,N_9500,N_9520);
xnor UO_196 (O_196,N_9726,N_9765);
nor UO_197 (O_197,N_9885,N_9864);
or UO_198 (O_198,N_9818,N_9928);
and UO_199 (O_199,N_9874,N_9775);
nand UO_200 (O_200,N_9521,N_9771);
or UO_201 (O_201,N_9902,N_9936);
or UO_202 (O_202,N_9703,N_9713);
or UO_203 (O_203,N_9881,N_9567);
nand UO_204 (O_204,N_9826,N_9548);
or UO_205 (O_205,N_9943,N_9721);
xor UO_206 (O_206,N_9683,N_9915);
or UO_207 (O_207,N_9660,N_9743);
and UO_208 (O_208,N_9941,N_9877);
nor UO_209 (O_209,N_9696,N_9512);
nand UO_210 (O_210,N_9615,N_9613);
nand UO_211 (O_211,N_9738,N_9782);
nand UO_212 (O_212,N_9817,N_9546);
nor UO_213 (O_213,N_9819,N_9517);
or UO_214 (O_214,N_9572,N_9711);
nor UO_215 (O_215,N_9880,N_9891);
nand UO_216 (O_216,N_9732,N_9857);
or UO_217 (O_217,N_9631,N_9764);
nor UO_218 (O_218,N_9604,N_9596);
nor UO_219 (O_219,N_9801,N_9769);
or UO_220 (O_220,N_9858,N_9658);
nor UO_221 (O_221,N_9914,N_9852);
and UO_222 (O_222,N_9598,N_9539);
or UO_223 (O_223,N_9692,N_9991);
or UO_224 (O_224,N_9588,N_9542);
nor UO_225 (O_225,N_9955,N_9664);
and UO_226 (O_226,N_9681,N_9522);
nand UO_227 (O_227,N_9737,N_9617);
or UO_228 (O_228,N_9870,N_9899);
xnor UO_229 (O_229,N_9981,N_9812);
nand UO_230 (O_230,N_9719,N_9577);
nor UO_231 (O_231,N_9556,N_9661);
xor UO_232 (O_232,N_9636,N_9980);
nand UO_233 (O_233,N_9642,N_9840);
xor UO_234 (O_234,N_9685,N_9833);
nor UO_235 (O_235,N_9927,N_9805);
and UO_236 (O_236,N_9869,N_9973);
and UO_237 (O_237,N_9918,N_9794);
nor UO_238 (O_238,N_9742,N_9948);
and UO_239 (O_239,N_9804,N_9722);
or UO_240 (O_240,N_9595,N_9832);
nor UO_241 (O_241,N_9624,N_9788);
nand UO_242 (O_242,N_9944,N_9576);
and UO_243 (O_243,N_9787,N_9762);
or UO_244 (O_244,N_9866,N_9997);
nor UO_245 (O_245,N_9513,N_9841);
nand UO_246 (O_246,N_9543,N_9544);
nand UO_247 (O_247,N_9800,N_9938);
or UO_248 (O_248,N_9982,N_9947);
or UO_249 (O_249,N_9605,N_9957);
nand UO_250 (O_250,N_9921,N_9950);
nor UO_251 (O_251,N_9512,N_9580);
nand UO_252 (O_252,N_9684,N_9936);
and UO_253 (O_253,N_9506,N_9991);
nand UO_254 (O_254,N_9513,N_9576);
or UO_255 (O_255,N_9573,N_9646);
or UO_256 (O_256,N_9643,N_9824);
or UO_257 (O_257,N_9798,N_9710);
nor UO_258 (O_258,N_9894,N_9566);
or UO_259 (O_259,N_9924,N_9541);
or UO_260 (O_260,N_9971,N_9940);
nand UO_261 (O_261,N_9822,N_9693);
and UO_262 (O_262,N_9744,N_9570);
xnor UO_263 (O_263,N_9520,N_9749);
nor UO_264 (O_264,N_9674,N_9556);
nor UO_265 (O_265,N_9705,N_9636);
and UO_266 (O_266,N_9600,N_9677);
nor UO_267 (O_267,N_9574,N_9914);
nor UO_268 (O_268,N_9885,N_9921);
nor UO_269 (O_269,N_9697,N_9684);
nor UO_270 (O_270,N_9735,N_9708);
nand UO_271 (O_271,N_9818,N_9881);
and UO_272 (O_272,N_9777,N_9939);
xnor UO_273 (O_273,N_9842,N_9686);
or UO_274 (O_274,N_9785,N_9726);
nand UO_275 (O_275,N_9800,N_9511);
nand UO_276 (O_276,N_9745,N_9800);
nor UO_277 (O_277,N_9880,N_9821);
and UO_278 (O_278,N_9599,N_9593);
and UO_279 (O_279,N_9674,N_9776);
or UO_280 (O_280,N_9786,N_9906);
and UO_281 (O_281,N_9825,N_9865);
or UO_282 (O_282,N_9908,N_9792);
xnor UO_283 (O_283,N_9746,N_9951);
nand UO_284 (O_284,N_9917,N_9933);
nand UO_285 (O_285,N_9678,N_9801);
xor UO_286 (O_286,N_9888,N_9672);
or UO_287 (O_287,N_9865,N_9929);
and UO_288 (O_288,N_9922,N_9829);
or UO_289 (O_289,N_9694,N_9946);
and UO_290 (O_290,N_9600,N_9594);
nor UO_291 (O_291,N_9726,N_9719);
nand UO_292 (O_292,N_9661,N_9561);
or UO_293 (O_293,N_9614,N_9665);
or UO_294 (O_294,N_9590,N_9953);
nand UO_295 (O_295,N_9770,N_9775);
nand UO_296 (O_296,N_9587,N_9818);
and UO_297 (O_297,N_9561,N_9721);
or UO_298 (O_298,N_9875,N_9539);
or UO_299 (O_299,N_9880,N_9720);
or UO_300 (O_300,N_9992,N_9596);
or UO_301 (O_301,N_9630,N_9568);
nor UO_302 (O_302,N_9625,N_9734);
nand UO_303 (O_303,N_9896,N_9910);
nor UO_304 (O_304,N_9992,N_9537);
or UO_305 (O_305,N_9964,N_9663);
and UO_306 (O_306,N_9627,N_9953);
nand UO_307 (O_307,N_9650,N_9676);
nor UO_308 (O_308,N_9500,N_9883);
or UO_309 (O_309,N_9558,N_9609);
nor UO_310 (O_310,N_9512,N_9915);
nand UO_311 (O_311,N_9860,N_9907);
nor UO_312 (O_312,N_9998,N_9945);
xnor UO_313 (O_313,N_9907,N_9929);
nand UO_314 (O_314,N_9501,N_9796);
and UO_315 (O_315,N_9686,N_9984);
or UO_316 (O_316,N_9917,N_9858);
or UO_317 (O_317,N_9802,N_9917);
nor UO_318 (O_318,N_9637,N_9680);
nor UO_319 (O_319,N_9775,N_9733);
nor UO_320 (O_320,N_9961,N_9812);
nand UO_321 (O_321,N_9932,N_9618);
and UO_322 (O_322,N_9627,N_9623);
nor UO_323 (O_323,N_9995,N_9538);
nand UO_324 (O_324,N_9727,N_9997);
nor UO_325 (O_325,N_9638,N_9622);
or UO_326 (O_326,N_9956,N_9533);
xnor UO_327 (O_327,N_9784,N_9621);
nand UO_328 (O_328,N_9553,N_9803);
or UO_329 (O_329,N_9974,N_9564);
and UO_330 (O_330,N_9529,N_9824);
or UO_331 (O_331,N_9866,N_9545);
nor UO_332 (O_332,N_9613,N_9654);
and UO_333 (O_333,N_9609,N_9985);
and UO_334 (O_334,N_9619,N_9684);
and UO_335 (O_335,N_9541,N_9683);
nor UO_336 (O_336,N_9748,N_9849);
and UO_337 (O_337,N_9645,N_9762);
and UO_338 (O_338,N_9719,N_9781);
or UO_339 (O_339,N_9553,N_9593);
xor UO_340 (O_340,N_9539,N_9746);
or UO_341 (O_341,N_9733,N_9502);
and UO_342 (O_342,N_9723,N_9561);
and UO_343 (O_343,N_9967,N_9544);
xor UO_344 (O_344,N_9861,N_9856);
nor UO_345 (O_345,N_9968,N_9611);
nand UO_346 (O_346,N_9935,N_9687);
and UO_347 (O_347,N_9571,N_9570);
xnor UO_348 (O_348,N_9857,N_9852);
nor UO_349 (O_349,N_9788,N_9720);
nand UO_350 (O_350,N_9801,N_9916);
nand UO_351 (O_351,N_9512,N_9506);
and UO_352 (O_352,N_9817,N_9968);
or UO_353 (O_353,N_9959,N_9777);
nor UO_354 (O_354,N_9672,N_9617);
nor UO_355 (O_355,N_9753,N_9742);
nor UO_356 (O_356,N_9945,N_9920);
or UO_357 (O_357,N_9742,N_9915);
nand UO_358 (O_358,N_9526,N_9719);
or UO_359 (O_359,N_9628,N_9669);
and UO_360 (O_360,N_9998,N_9816);
nand UO_361 (O_361,N_9889,N_9845);
xnor UO_362 (O_362,N_9957,N_9594);
nand UO_363 (O_363,N_9964,N_9594);
and UO_364 (O_364,N_9809,N_9717);
and UO_365 (O_365,N_9556,N_9853);
nor UO_366 (O_366,N_9693,N_9533);
and UO_367 (O_367,N_9705,N_9517);
or UO_368 (O_368,N_9636,N_9658);
nor UO_369 (O_369,N_9734,N_9659);
nor UO_370 (O_370,N_9811,N_9807);
and UO_371 (O_371,N_9838,N_9607);
or UO_372 (O_372,N_9930,N_9562);
and UO_373 (O_373,N_9835,N_9555);
nor UO_374 (O_374,N_9557,N_9658);
or UO_375 (O_375,N_9630,N_9948);
nand UO_376 (O_376,N_9598,N_9601);
nand UO_377 (O_377,N_9723,N_9914);
and UO_378 (O_378,N_9622,N_9534);
nor UO_379 (O_379,N_9536,N_9523);
and UO_380 (O_380,N_9601,N_9917);
nand UO_381 (O_381,N_9990,N_9631);
or UO_382 (O_382,N_9959,N_9743);
nor UO_383 (O_383,N_9953,N_9576);
or UO_384 (O_384,N_9959,N_9659);
or UO_385 (O_385,N_9575,N_9957);
nand UO_386 (O_386,N_9876,N_9658);
and UO_387 (O_387,N_9803,N_9993);
and UO_388 (O_388,N_9518,N_9504);
or UO_389 (O_389,N_9961,N_9896);
and UO_390 (O_390,N_9723,N_9548);
nor UO_391 (O_391,N_9689,N_9927);
and UO_392 (O_392,N_9579,N_9503);
xnor UO_393 (O_393,N_9558,N_9744);
nor UO_394 (O_394,N_9802,N_9548);
and UO_395 (O_395,N_9590,N_9827);
nand UO_396 (O_396,N_9807,N_9642);
nand UO_397 (O_397,N_9516,N_9514);
or UO_398 (O_398,N_9954,N_9910);
nor UO_399 (O_399,N_9886,N_9825);
or UO_400 (O_400,N_9901,N_9651);
xor UO_401 (O_401,N_9968,N_9608);
nor UO_402 (O_402,N_9896,N_9921);
xnor UO_403 (O_403,N_9944,N_9821);
nand UO_404 (O_404,N_9941,N_9799);
nand UO_405 (O_405,N_9609,N_9617);
and UO_406 (O_406,N_9522,N_9642);
nand UO_407 (O_407,N_9886,N_9646);
and UO_408 (O_408,N_9577,N_9667);
and UO_409 (O_409,N_9911,N_9813);
or UO_410 (O_410,N_9643,N_9780);
or UO_411 (O_411,N_9503,N_9820);
nor UO_412 (O_412,N_9530,N_9993);
nand UO_413 (O_413,N_9653,N_9594);
nand UO_414 (O_414,N_9600,N_9718);
or UO_415 (O_415,N_9636,N_9569);
nand UO_416 (O_416,N_9755,N_9863);
and UO_417 (O_417,N_9683,N_9826);
and UO_418 (O_418,N_9868,N_9778);
or UO_419 (O_419,N_9737,N_9716);
nand UO_420 (O_420,N_9696,N_9551);
nor UO_421 (O_421,N_9966,N_9842);
and UO_422 (O_422,N_9942,N_9564);
nor UO_423 (O_423,N_9728,N_9713);
or UO_424 (O_424,N_9579,N_9731);
or UO_425 (O_425,N_9636,N_9790);
nor UO_426 (O_426,N_9834,N_9630);
or UO_427 (O_427,N_9878,N_9868);
and UO_428 (O_428,N_9741,N_9856);
and UO_429 (O_429,N_9984,N_9531);
nand UO_430 (O_430,N_9746,N_9634);
and UO_431 (O_431,N_9605,N_9727);
or UO_432 (O_432,N_9977,N_9995);
nand UO_433 (O_433,N_9949,N_9953);
xor UO_434 (O_434,N_9602,N_9839);
and UO_435 (O_435,N_9736,N_9813);
and UO_436 (O_436,N_9921,N_9887);
xor UO_437 (O_437,N_9718,N_9646);
nor UO_438 (O_438,N_9638,N_9556);
and UO_439 (O_439,N_9690,N_9622);
nand UO_440 (O_440,N_9649,N_9808);
nor UO_441 (O_441,N_9787,N_9942);
nor UO_442 (O_442,N_9616,N_9514);
or UO_443 (O_443,N_9677,N_9855);
or UO_444 (O_444,N_9936,N_9595);
nor UO_445 (O_445,N_9503,N_9658);
nor UO_446 (O_446,N_9733,N_9643);
nor UO_447 (O_447,N_9523,N_9500);
xnor UO_448 (O_448,N_9706,N_9571);
nor UO_449 (O_449,N_9791,N_9965);
xor UO_450 (O_450,N_9540,N_9595);
and UO_451 (O_451,N_9681,N_9964);
and UO_452 (O_452,N_9611,N_9846);
and UO_453 (O_453,N_9610,N_9633);
nor UO_454 (O_454,N_9767,N_9541);
nand UO_455 (O_455,N_9840,N_9846);
nand UO_456 (O_456,N_9522,N_9914);
nand UO_457 (O_457,N_9525,N_9651);
nand UO_458 (O_458,N_9511,N_9723);
and UO_459 (O_459,N_9552,N_9989);
xor UO_460 (O_460,N_9559,N_9850);
nand UO_461 (O_461,N_9767,N_9708);
and UO_462 (O_462,N_9974,N_9910);
and UO_463 (O_463,N_9885,N_9733);
nor UO_464 (O_464,N_9694,N_9697);
nor UO_465 (O_465,N_9607,N_9855);
or UO_466 (O_466,N_9999,N_9899);
nand UO_467 (O_467,N_9969,N_9590);
nor UO_468 (O_468,N_9678,N_9957);
nand UO_469 (O_469,N_9556,N_9766);
nor UO_470 (O_470,N_9658,N_9975);
nor UO_471 (O_471,N_9785,N_9939);
xnor UO_472 (O_472,N_9963,N_9587);
nor UO_473 (O_473,N_9979,N_9969);
and UO_474 (O_474,N_9840,N_9514);
nand UO_475 (O_475,N_9611,N_9555);
xnor UO_476 (O_476,N_9815,N_9868);
nand UO_477 (O_477,N_9819,N_9505);
nand UO_478 (O_478,N_9660,N_9681);
or UO_479 (O_479,N_9781,N_9928);
xnor UO_480 (O_480,N_9728,N_9752);
nor UO_481 (O_481,N_9827,N_9627);
or UO_482 (O_482,N_9667,N_9972);
and UO_483 (O_483,N_9917,N_9510);
and UO_484 (O_484,N_9901,N_9707);
nor UO_485 (O_485,N_9973,N_9953);
or UO_486 (O_486,N_9800,N_9823);
and UO_487 (O_487,N_9854,N_9857);
xnor UO_488 (O_488,N_9562,N_9946);
nor UO_489 (O_489,N_9880,N_9789);
nand UO_490 (O_490,N_9722,N_9724);
and UO_491 (O_491,N_9928,N_9544);
and UO_492 (O_492,N_9615,N_9695);
and UO_493 (O_493,N_9898,N_9500);
or UO_494 (O_494,N_9774,N_9851);
nor UO_495 (O_495,N_9707,N_9847);
nor UO_496 (O_496,N_9870,N_9880);
nor UO_497 (O_497,N_9744,N_9888);
xnor UO_498 (O_498,N_9721,N_9812);
or UO_499 (O_499,N_9708,N_9998);
or UO_500 (O_500,N_9942,N_9580);
or UO_501 (O_501,N_9711,N_9769);
and UO_502 (O_502,N_9909,N_9895);
and UO_503 (O_503,N_9677,N_9700);
xnor UO_504 (O_504,N_9918,N_9944);
nand UO_505 (O_505,N_9685,N_9895);
and UO_506 (O_506,N_9846,N_9602);
nand UO_507 (O_507,N_9548,N_9894);
nor UO_508 (O_508,N_9535,N_9598);
nand UO_509 (O_509,N_9813,N_9967);
or UO_510 (O_510,N_9722,N_9781);
nand UO_511 (O_511,N_9706,N_9803);
nor UO_512 (O_512,N_9510,N_9782);
and UO_513 (O_513,N_9693,N_9630);
or UO_514 (O_514,N_9829,N_9991);
nor UO_515 (O_515,N_9737,N_9618);
nand UO_516 (O_516,N_9737,N_9651);
nand UO_517 (O_517,N_9628,N_9506);
nor UO_518 (O_518,N_9938,N_9579);
nor UO_519 (O_519,N_9873,N_9892);
xor UO_520 (O_520,N_9839,N_9726);
or UO_521 (O_521,N_9607,N_9885);
and UO_522 (O_522,N_9809,N_9902);
or UO_523 (O_523,N_9514,N_9727);
and UO_524 (O_524,N_9948,N_9860);
or UO_525 (O_525,N_9855,N_9568);
nand UO_526 (O_526,N_9827,N_9833);
xnor UO_527 (O_527,N_9802,N_9954);
xnor UO_528 (O_528,N_9555,N_9653);
and UO_529 (O_529,N_9502,N_9611);
xor UO_530 (O_530,N_9732,N_9693);
nand UO_531 (O_531,N_9743,N_9623);
nand UO_532 (O_532,N_9770,N_9574);
or UO_533 (O_533,N_9510,N_9634);
and UO_534 (O_534,N_9979,N_9746);
and UO_535 (O_535,N_9992,N_9658);
nand UO_536 (O_536,N_9946,N_9701);
nand UO_537 (O_537,N_9581,N_9586);
nor UO_538 (O_538,N_9802,N_9556);
nand UO_539 (O_539,N_9921,N_9586);
nor UO_540 (O_540,N_9898,N_9534);
nor UO_541 (O_541,N_9677,N_9569);
xor UO_542 (O_542,N_9627,N_9710);
and UO_543 (O_543,N_9567,N_9697);
and UO_544 (O_544,N_9522,N_9769);
nand UO_545 (O_545,N_9941,N_9842);
nand UO_546 (O_546,N_9715,N_9853);
xor UO_547 (O_547,N_9969,N_9578);
nand UO_548 (O_548,N_9810,N_9640);
xor UO_549 (O_549,N_9899,N_9564);
nand UO_550 (O_550,N_9548,N_9732);
xor UO_551 (O_551,N_9997,N_9823);
or UO_552 (O_552,N_9650,N_9633);
or UO_553 (O_553,N_9675,N_9957);
nor UO_554 (O_554,N_9757,N_9904);
nor UO_555 (O_555,N_9654,N_9799);
or UO_556 (O_556,N_9573,N_9858);
and UO_557 (O_557,N_9611,N_9735);
or UO_558 (O_558,N_9754,N_9597);
or UO_559 (O_559,N_9875,N_9593);
nand UO_560 (O_560,N_9972,N_9845);
and UO_561 (O_561,N_9537,N_9839);
and UO_562 (O_562,N_9752,N_9981);
xnor UO_563 (O_563,N_9968,N_9588);
and UO_564 (O_564,N_9892,N_9867);
or UO_565 (O_565,N_9994,N_9915);
nand UO_566 (O_566,N_9594,N_9916);
or UO_567 (O_567,N_9670,N_9580);
nor UO_568 (O_568,N_9640,N_9977);
nor UO_569 (O_569,N_9764,N_9991);
xor UO_570 (O_570,N_9608,N_9697);
nor UO_571 (O_571,N_9949,N_9675);
and UO_572 (O_572,N_9698,N_9814);
or UO_573 (O_573,N_9674,N_9891);
xor UO_574 (O_574,N_9640,N_9535);
and UO_575 (O_575,N_9786,N_9677);
or UO_576 (O_576,N_9931,N_9958);
or UO_577 (O_577,N_9618,N_9515);
and UO_578 (O_578,N_9544,N_9942);
and UO_579 (O_579,N_9980,N_9826);
and UO_580 (O_580,N_9513,N_9958);
nand UO_581 (O_581,N_9598,N_9733);
or UO_582 (O_582,N_9983,N_9970);
nand UO_583 (O_583,N_9991,N_9835);
and UO_584 (O_584,N_9557,N_9755);
or UO_585 (O_585,N_9742,N_9545);
and UO_586 (O_586,N_9519,N_9961);
or UO_587 (O_587,N_9526,N_9691);
and UO_588 (O_588,N_9768,N_9713);
and UO_589 (O_589,N_9677,N_9580);
nand UO_590 (O_590,N_9712,N_9520);
or UO_591 (O_591,N_9672,N_9629);
nor UO_592 (O_592,N_9679,N_9533);
xnor UO_593 (O_593,N_9530,N_9791);
and UO_594 (O_594,N_9623,N_9719);
or UO_595 (O_595,N_9699,N_9693);
nand UO_596 (O_596,N_9717,N_9886);
nor UO_597 (O_597,N_9547,N_9802);
nand UO_598 (O_598,N_9990,N_9811);
or UO_599 (O_599,N_9765,N_9566);
nand UO_600 (O_600,N_9532,N_9699);
and UO_601 (O_601,N_9852,N_9944);
or UO_602 (O_602,N_9589,N_9615);
or UO_603 (O_603,N_9828,N_9926);
nor UO_604 (O_604,N_9741,N_9868);
and UO_605 (O_605,N_9743,N_9703);
and UO_606 (O_606,N_9849,N_9553);
and UO_607 (O_607,N_9984,N_9899);
nor UO_608 (O_608,N_9977,N_9592);
nand UO_609 (O_609,N_9986,N_9700);
and UO_610 (O_610,N_9873,N_9668);
and UO_611 (O_611,N_9773,N_9571);
or UO_612 (O_612,N_9847,N_9756);
nor UO_613 (O_613,N_9581,N_9693);
and UO_614 (O_614,N_9568,N_9554);
nand UO_615 (O_615,N_9831,N_9666);
or UO_616 (O_616,N_9963,N_9855);
nor UO_617 (O_617,N_9634,N_9782);
nand UO_618 (O_618,N_9960,N_9723);
and UO_619 (O_619,N_9693,N_9648);
nand UO_620 (O_620,N_9514,N_9723);
nand UO_621 (O_621,N_9532,N_9627);
xnor UO_622 (O_622,N_9823,N_9810);
and UO_623 (O_623,N_9633,N_9733);
and UO_624 (O_624,N_9741,N_9527);
nor UO_625 (O_625,N_9944,N_9961);
and UO_626 (O_626,N_9696,N_9614);
or UO_627 (O_627,N_9951,N_9522);
nor UO_628 (O_628,N_9725,N_9613);
and UO_629 (O_629,N_9835,N_9827);
or UO_630 (O_630,N_9569,N_9578);
and UO_631 (O_631,N_9540,N_9527);
and UO_632 (O_632,N_9657,N_9508);
nand UO_633 (O_633,N_9642,N_9526);
and UO_634 (O_634,N_9609,N_9897);
or UO_635 (O_635,N_9952,N_9916);
or UO_636 (O_636,N_9561,N_9727);
nor UO_637 (O_637,N_9683,N_9746);
nor UO_638 (O_638,N_9735,N_9562);
and UO_639 (O_639,N_9508,N_9777);
nand UO_640 (O_640,N_9892,N_9600);
or UO_641 (O_641,N_9679,N_9600);
and UO_642 (O_642,N_9959,N_9732);
xnor UO_643 (O_643,N_9803,N_9901);
nor UO_644 (O_644,N_9565,N_9961);
nand UO_645 (O_645,N_9597,N_9984);
and UO_646 (O_646,N_9583,N_9906);
or UO_647 (O_647,N_9589,N_9984);
or UO_648 (O_648,N_9639,N_9981);
and UO_649 (O_649,N_9858,N_9730);
nor UO_650 (O_650,N_9631,N_9858);
nor UO_651 (O_651,N_9988,N_9875);
nor UO_652 (O_652,N_9522,N_9623);
nand UO_653 (O_653,N_9500,N_9577);
nand UO_654 (O_654,N_9889,N_9536);
nand UO_655 (O_655,N_9663,N_9719);
xnor UO_656 (O_656,N_9550,N_9728);
nand UO_657 (O_657,N_9772,N_9762);
and UO_658 (O_658,N_9643,N_9554);
nand UO_659 (O_659,N_9687,N_9973);
and UO_660 (O_660,N_9587,N_9677);
xor UO_661 (O_661,N_9970,N_9694);
nand UO_662 (O_662,N_9742,N_9506);
and UO_663 (O_663,N_9640,N_9547);
nor UO_664 (O_664,N_9850,N_9711);
or UO_665 (O_665,N_9695,N_9710);
or UO_666 (O_666,N_9803,N_9544);
and UO_667 (O_667,N_9574,N_9678);
and UO_668 (O_668,N_9901,N_9617);
and UO_669 (O_669,N_9812,N_9833);
and UO_670 (O_670,N_9817,N_9763);
or UO_671 (O_671,N_9598,N_9532);
and UO_672 (O_672,N_9839,N_9714);
nor UO_673 (O_673,N_9771,N_9545);
or UO_674 (O_674,N_9922,N_9924);
and UO_675 (O_675,N_9654,N_9571);
nand UO_676 (O_676,N_9757,N_9918);
and UO_677 (O_677,N_9511,N_9813);
nor UO_678 (O_678,N_9926,N_9943);
and UO_679 (O_679,N_9973,N_9694);
nand UO_680 (O_680,N_9553,N_9537);
nand UO_681 (O_681,N_9578,N_9547);
nor UO_682 (O_682,N_9711,N_9773);
or UO_683 (O_683,N_9511,N_9809);
nand UO_684 (O_684,N_9882,N_9677);
nand UO_685 (O_685,N_9531,N_9634);
nand UO_686 (O_686,N_9732,N_9781);
and UO_687 (O_687,N_9666,N_9526);
or UO_688 (O_688,N_9992,N_9855);
and UO_689 (O_689,N_9524,N_9755);
nor UO_690 (O_690,N_9663,N_9883);
and UO_691 (O_691,N_9923,N_9962);
or UO_692 (O_692,N_9531,N_9986);
xor UO_693 (O_693,N_9619,N_9866);
xnor UO_694 (O_694,N_9859,N_9588);
nand UO_695 (O_695,N_9857,N_9989);
nor UO_696 (O_696,N_9937,N_9902);
nand UO_697 (O_697,N_9650,N_9954);
and UO_698 (O_698,N_9897,N_9697);
nand UO_699 (O_699,N_9688,N_9597);
xor UO_700 (O_700,N_9804,N_9884);
or UO_701 (O_701,N_9824,N_9670);
nand UO_702 (O_702,N_9777,N_9502);
nor UO_703 (O_703,N_9889,N_9907);
and UO_704 (O_704,N_9548,N_9557);
or UO_705 (O_705,N_9900,N_9668);
or UO_706 (O_706,N_9516,N_9693);
nor UO_707 (O_707,N_9930,N_9861);
nand UO_708 (O_708,N_9630,N_9726);
nor UO_709 (O_709,N_9592,N_9777);
nor UO_710 (O_710,N_9868,N_9629);
nor UO_711 (O_711,N_9546,N_9976);
and UO_712 (O_712,N_9876,N_9848);
or UO_713 (O_713,N_9819,N_9965);
nor UO_714 (O_714,N_9610,N_9915);
and UO_715 (O_715,N_9866,N_9912);
nor UO_716 (O_716,N_9767,N_9851);
and UO_717 (O_717,N_9597,N_9526);
or UO_718 (O_718,N_9748,N_9559);
or UO_719 (O_719,N_9587,N_9966);
xnor UO_720 (O_720,N_9701,N_9813);
and UO_721 (O_721,N_9705,N_9655);
xnor UO_722 (O_722,N_9659,N_9664);
and UO_723 (O_723,N_9607,N_9536);
or UO_724 (O_724,N_9846,N_9576);
nor UO_725 (O_725,N_9842,N_9955);
nand UO_726 (O_726,N_9905,N_9934);
nor UO_727 (O_727,N_9739,N_9543);
and UO_728 (O_728,N_9561,N_9949);
or UO_729 (O_729,N_9964,N_9548);
nor UO_730 (O_730,N_9666,N_9556);
nand UO_731 (O_731,N_9800,N_9580);
and UO_732 (O_732,N_9542,N_9939);
nand UO_733 (O_733,N_9832,N_9547);
and UO_734 (O_734,N_9632,N_9614);
and UO_735 (O_735,N_9508,N_9972);
nor UO_736 (O_736,N_9607,N_9783);
and UO_737 (O_737,N_9857,N_9717);
nand UO_738 (O_738,N_9787,N_9684);
nand UO_739 (O_739,N_9708,N_9586);
and UO_740 (O_740,N_9655,N_9636);
nor UO_741 (O_741,N_9600,N_9963);
or UO_742 (O_742,N_9761,N_9954);
nor UO_743 (O_743,N_9764,N_9856);
xor UO_744 (O_744,N_9840,N_9999);
or UO_745 (O_745,N_9757,N_9574);
nand UO_746 (O_746,N_9644,N_9625);
nand UO_747 (O_747,N_9585,N_9916);
nor UO_748 (O_748,N_9832,N_9731);
nand UO_749 (O_749,N_9553,N_9811);
and UO_750 (O_750,N_9694,N_9531);
nor UO_751 (O_751,N_9516,N_9877);
nand UO_752 (O_752,N_9908,N_9972);
nand UO_753 (O_753,N_9808,N_9560);
or UO_754 (O_754,N_9679,N_9738);
nor UO_755 (O_755,N_9806,N_9505);
or UO_756 (O_756,N_9623,N_9735);
or UO_757 (O_757,N_9689,N_9511);
and UO_758 (O_758,N_9768,N_9735);
and UO_759 (O_759,N_9714,N_9809);
xnor UO_760 (O_760,N_9762,N_9973);
and UO_761 (O_761,N_9726,N_9584);
or UO_762 (O_762,N_9764,N_9508);
nor UO_763 (O_763,N_9944,N_9775);
nor UO_764 (O_764,N_9854,N_9642);
and UO_765 (O_765,N_9911,N_9688);
or UO_766 (O_766,N_9549,N_9761);
and UO_767 (O_767,N_9776,N_9716);
or UO_768 (O_768,N_9925,N_9669);
nor UO_769 (O_769,N_9995,N_9757);
nand UO_770 (O_770,N_9962,N_9953);
and UO_771 (O_771,N_9754,N_9805);
xor UO_772 (O_772,N_9706,N_9832);
or UO_773 (O_773,N_9872,N_9819);
and UO_774 (O_774,N_9818,N_9966);
or UO_775 (O_775,N_9791,N_9637);
xnor UO_776 (O_776,N_9902,N_9870);
nor UO_777 (O_777,N_9726,N_9993);
nand UO_778 (O_778,N_9646,N_9501);
or UO_779 (O_779,N_9588,N_9604);
nor UO_780 (O_780,N_9628,N_9670);
or UO_781 (O_781,N_9754,N_9599);
or UO_782 (O_782,N_9802,N_9546);
nor UO_783 (O_783,N_9663,N_9894);
and UO_784 (O_784,N_9965,N_9848);
or UO_785 (O_785,N_9691,N_9990);
or UO_786 (O_786,N_9850,N_9766);
xor UO_787 (O_787,N_9556,N_9612);
nor UO_788 (O_788,N_9875,N_9917);
and UO_789 (O_789,N_9865,N_9615);
nor UO_790 (O_790,N_9787,N_9945);
nor UO_791 (O_791,N_9951,N_9668);
or UO_792 (O_792,N_9606,N_9515);
or UO_793 (O_793,N_9646,N_9864);
nor UO_794 (O_794,N_9766,N_9510);
or UO_795 (O_795,N_9600,N_9689);
xnor UO_796 (O_796,N_9683,N_9824);
nand UO_797 (O_797,N_9728,N_9810);
and UO_798 (O_798,N_9987,N_9703);
nand UO_799 (O_799,N_9820,N_9886);
and UO_800 (O_800,N_9849,N_9692);
nor UO_801 (O_801,N_9552,N_9713);
or UO_802 (O_802,N_9930,N_9981);
and UO_803 (O_803,N_9722,N_9663);
nor UO_804 (O_804,N_9854,N_9526);
nand UO_805 (O_805,N_9873,N_9900);
nor UO_806 (O_806,N_9658,N_9621);
xor UO_807 (O_807,N_9545,N_9685);
xnor UO_808 (O_808,N_9533,N_9889);
or UO_809 (O_809,N_9992,N_9818);
nand UO_810 (O_810,N_9803,N_9561);
nor UO_811 (O_811,N_9807,N_9998);
or UO_812 (O_812,N_9835,N_9995);
and UO_813 (O_813,N_9655,N_9738);
and UO_814 (O_814,N_9906,N_9983);
or UO_815 (O_815,N_9745,N_9970);
nor UO_816 (O_816,N_9739,N_9559);
and UO_817 (O_817,N_9933,N_9851);
or UO_818 (O_818,N_9869,N_9844);
and UO_819 (O_819,N_9769,N_9690);
and UO_820 (O_820,N_9786,N_9718);
and UO_821 (O_821,N_9931,N_9512);
or UO_822 (O_822,N_9617,N_9990);
nand UO_823 (O_823,N_9642,N_9665);
nand UO_824 (O_824,N_9662,N_9717);
nor UO_825 (O_825,N_9561,N_9562);
or UO_826 (O_826,N_9924,N_9971);
and UO_827 (O_827,N_9905,N_9605);
or UO_828 (O_828,N_9825,N_9884);
nand UO_829 (O_829,N_9886,N_9655);
and UO_830 (O_830,N_9729,N_9627);
nor UO_831 (O_831,N_9748,N_9922);
nand UO_832 (O_832,N_9935,N_9891);
xor UO_833 (O_833,N_9540,N_9892);
nor UO_834 (O_834,N_9667,N_9765);
nand UO_835 (O_835,N_9781,N_9734);
xnor UO_836 (O_836,N_9782,N_9879);
or UO_837 (O_837,N_9558,N_9538);
and UO_838 (O_838,N_9569,N_9894);
nor UO_839 (O_839,N_9604,N_9841);
or UO_840 (O_840,N_9657,N_9541);
xor UO_841 (O_841,N_9674,N_9700);
and UO_842 (O_842,N_9706,N_9737);
or UO_843 (O_843,N_9585,N_9940);
or UO_844 (O_844,N_9509,N_9887);
nand UO_845 (O_845,N_9951,N_9848);
nor UO_846 (O_846,N_9743,N_9513);
or UO_847 (O_847,N_9698,N_9544);
nor UO_848 (O_848,N_9717,N_9913);
and UO_849 (O_849,N_9757,N_9776);
and UO_850 (O_850,N_9549,N_9623);
xnor UO_851 (O_851,N_9889,N_9724);
nand UO_852 (O_852,N_9513,N_9527);
and UO_853 (O_853,N_9695,N_9613);
or UO_854 (O_854,N_9666,N_9601);
nor UO_855 (O_855,N_9887,N_9586);
or UO_856 (O_856,N_9989,N_9569);
and UO_857 (O_857,N_9567,N_9502);
or UO_858 (O_858,N_9899,N_9561);
xnor UO_859 (O_859,N_9795,N_9866);
and UO_860 (O_860,N_9928,N_9776);
nand UO_861 (O_861,N_9980,N_9962);
or UO_862 (O_862,N_9881,N_9940);
or UO_863 (O_863,N_9952,N_9849);
nand UO_864 (O_864,N_9671,N_9873);
nand UO_865 (O_865,N_9692,N_9809);
and UO_866 (O_866,N_9731,N_9523);
or UO_867 (O_867,N_9810,N_9775);
nand UO_868 (O_868,N_9912,N_9785);
nand UO_869 (O_869,N_9725,N_9877);
nor UO_870 (O_870,N_9923,N_9850);
or UO_871 (O_871,N_9965,N_9812);
and UO_872 (O_872,N_9851,N_9700);
xor UO_873 (O_873,N_9568,N_9957);
nand UO_874 (O_874,N_9534,N_9620);
and UO_875 (O_875,N_9969,N_9580);
or UO_876 (O_876,N_9904,N_9693);
or UO_877 (O_877,N_9857,N_9741);
nand UO_878 (O_878,N_9999,N_9723);
xor UO_879 (O_879,N_9721,N_9645);
nand UO_880 (O_880,N_9848,N_9769);
nand UO_881 (O_881,N_9865,N_9872);
or UO_882 (O_882,N_9581,N_9520);
or UO_883 (O_883,N_9777,N_9833);
xor UO_884 (O_884,N_9812,N_9694);
nand UO_885 (O_885,N_9552,N_9580);
or UO_886 (O_886,N_9858,N_9871);
or UO_887 (O_887,N_9725,N_9850);
nor UO_888 (O_888,N_9556,N_9826);
and UO_889 (O_889,N_9929,N_9984);
and UO_890 (O_890,N_9613,N_9784);
and UO_891 (O_891,N_9864,N_9824);
nand UO_892 (O_892,N_9546,N_9890);
or UO_893 (O_893,N_9908,N_9699);
or UO_894 (O_894,N_9584,N_9665);
or UO_895 (O_895,N_9572,N_9612);
nor UO_896 (O_896,N_9941,N_9530);
nor UO_897 (O_897,N_9878,N_9575);
and UO_898 (O_898,N_9978,N_9920);
nand UO_899 (O_899,N_9606,N_9599);
or UO_900 (O_900,N_9935,N_9729);
or UO_901 (O_901,N_9566,N_9853);
or UO_902 (O_902,N_9573,N_9520);
nand UO_903 (O_903,N_9912,N_9536);
and UO_904 (O_904,N_9966,N_9762);
and UO_905 (O_905,N_9971,N_9537);
or UO_906 (O_906,N_9681,N_9667);
and UO_907 (O_907,N_9727,N_9816);
and UO_908 (O_908,N_9959,N_9799);
nor UO_909 (O_909,N_9906,N_9777);
nor UO_910 (O_910,N_9776,N_9778);
and UO_911 (O_911,N_9732,N_9897);
or UO_912 (O_912,N_9750,N_9960);
and UO_913 (O_913,N_9690,N_9781);
or UO_914 (O_914,N_9935,N_9886);
or UO_915 (O_915,N_9746,N_9635);
nor UO_916 (O_916,N_9687,N_9692);
or UO_917 (O_917,N_9893,N_9975);
nand UO_918 (O_918,N_9735,N_9984);
and UO_919 (O_919,N_9862,N_9927);
and UO_920 (O_920,N_9895,N_9619);
or UO_921 (O_921,N_9622,N_9572);
nand UO_922 (O_922,N_9505,N_9955);
xor UO_923 (O_923,N_9610,N_9592);
nand UO_924 (O_924,N_9628,N_9574);
nand UO_925 (O_925,N_9832,N_9519);
nor UO_926 (O_926,N_9733,N_9599);
or UO_927 (O_927,N_9712,N_9915);
nor UO_928 (O_928,N_9692,N_9660);
or UO_929 (O_929,N_9778,N_9818);
nand UO_930 (O_930,N_9688,N_9852);
xor UO_931 (O_931,N_9837,N_9787);
and UO_932 (O_932,N_9576,N_9965);
nor UO_933 (O_933,N_9622,N_9506);
nor UO_934 (O_934,N_9779,N_9630);
nand UO_935 (O_935,N_9620,N_9927);
or UO_936 (O_936,N_9870,N_9708);
or UO_937 (O_937,N_9517,N_9589);
nand UO_938 (O_938,N_9950,N_9851);
or UO_939 (O_939,N_9550,N_9693);
or UO_940 (O_940,N_9692,N_9502);
and UO_941 (O_941,N_9986,N_9966);
and UO_942 (O_942,N_9529,N_9751);
or UO_943 (O_943,N_9713,N_9558);
nor UO_944 (O_944,N_9824,N_9792);
and UO_945 (O_945,N_9614,N_9957);
and UO_946 (O_946,N_9667,N_9896);
and UO_947 (O_947,N_9753,N_9900);
nand UO_948 (O_948,N_9902,N_9979);
nor UO_949 (O_949,N_9643,N_9903);
nor UO_950 (O_950,N_9504,N_9662);
nor UO_951 (O_951,N_9673,N_9670);
or UO_952 (O_952,N_9949,N_9987);
or UO_953 (O_953,N_9512,N_9841);
xnor UO_954 (O_954,N_9537,N_9949);
and UO_955 (O_955,N_9907,N_9614);
nor UO_956 (O_956,N_9777,N_9519);
nor UO_957 (O_957,N_9959,N_9656);
nor UO_958 (O_958,N_9696,N_9687);
or UO_959 (O_959,N_9696,N_9626);
nor UO_960 (O_960,N_9877,N_9513);
and UO_961 (O_961,N_9976,N_9715);
xor UO_962 (O_962,N_9976,N_9905);
or UO_963 (O_963,N_9671,N_9517);
and UO_964 (O_964,N_9629,N_9741);
xnor UO_965 (O_965,N_9597,N_9900);
nand UO_966 (O_966,N_9739,N_9847);
or UO_967 (O_967,N_9791,N_9735);
or UO_968 (O_968,N_9668,N_9563);
nor UO_969 (O_969,N_9528,N_9991);
or UO_970 (O_970,N_9627,N_9711);
and UO_971 (O_971,N_9702,N_9876);
nor UO_972 (O_972,N_9542,N_9756);
or UO_973 (O_973,N_9653,N_9695);
or UO_974 (O_974,N_9741,N_9528);
xnor UO_975 (O_975,N_9580,N_9950);
nor UO_976 (O_976,N_9919,N_9996);
and UO_977 (O_977,N_9858,N_9583);
and UO_978 (O_978,N_9525,N_9871);
or UO_979 (O_979,N_9703,N_9898);
nand UO_980 (O_980,N_9804,N_9816);
xnor UO_981 (O_981,N_9887,N_9780);
and UO_982 (O_982,N_9655,N_9610);
nand UO_983 (O_983,N_9724,N_9796);
nand UO_984 (O_984,N_9629,N_9758);
and UO_985 (O_985,N_9803,N_9765);
nand UO_986 (O_986,N_9838,N_9708);
nor UO_987 (O_987,N_9745,N_9655);
xor UO_988 (O_988,N_9814,N_9584);
nand UO_989 (O_989,N_9845,N_9753);
and UO_990 (O_990,N_9715,N_9726);
and UO_991 (O_991,N_9862,N_9891);
nor UO_992 (O_992,N_9689,N_9681);
nor UO_993 (O_993,N_9835,N_9917);
or UO_994 (O_994,N_9982,N_9687);
nand UO_995 (O_995,N_9990,N_9598);
xnor UO_996 (O_996,N_9961,N_9697);
and UO_997 (O_997,N_9794,N_9510);
or UO_998 (O_998,N_9572,N_9615);
and UO_999 (O_999,N_9608,N_9506);
xor UO_1000 (O_1000,N_9549,N_9567);
nand UO_1001 (O_1001,N_9943,N_9557);
nor UO_1002 (O_1002,N_9926,N_9537);
nand UO_1003 (O_1003,N_9733,N_9932);
and UO_1004 (O_1004,N_9575,N_9671);
and UO_1005 (O_1005,N_9692,N_9705);
xnor UO_1006 (O_1006,N_9585,N_9512);
and UO_1007 (O_1007,N_9991,N_9538);
nand UO_1008 (O_1008,N_9619,N_9704);
nor UO_1009 (O_1009,N_9778,N_9530);
or UO_1010 (O_1010,N_9965,N_9529);
nor UO_1011 (O_1011,N_9671,N_9936);
nor UO_1012 (O_1012,N_9506,N_9777);
nor UO_1013 (O_1013,N_9584,N_9711);
nand UO_1014 (O_1014,N_9523,N_9767);
nand UO_1015 (O_1015,N_9910,N_9865);
nor UO_1016 (O_1016,N_9700,N_9953);
nand UO_1017 (O_1017,N_9637,N_9745);
nor UO_1018 (O_1018,N_9990,N_9915);
nor UO_1019 (O_1019,N_9573,N_9599);
or UO_1020 (O_1020,N_9879,N_9532);
or UO_1021 (O_1021,N_9868,N_9527);
nor UO_1022 (O_1022,N_9681,N_9852);
nor UO_1023 (O_1023,N_9611,N_9865);
nand UO_1024 (O_1024,N_9728,N_9890);
nor UO_1025 (O_1025,N_9969,N_9960);
nor UO_1026 (O_1026,N_9636,N_9796);
nand UO_1027 (O_1027,N_9635,N_9948);
nor UO_1028 (O_1028,N_9672,N_9625);
and UO_1029 (O_1029,N_9699,N_9613);
and UO_1030 (O_1030,N_9719,N_9706);
xor UO_1031 (O_1031,N_9808,N_9915);
nor UO_1032 (O_1032,N_9523,N_9544);
and UO_1033 (O_1033,N_9779,N_9599);
or UO_1034 (O_1034,N_9970,N_9973);
nor UO_1035 (O_1035,N_9703,N_9890);
or UO_1036 (O_1036,N_9729,N_9663);
nand UO_1037 (O_1037,N_9612,N_9585);
nor UO_1038 (O_1038,N_9976,N_9843);
nand UO_1039 (O_1039,N_9741,N_9676);
and UO_1040 (O_1040,N_9819,N_9746);
or UO_1041 (O_1041,N_9515,N_9676);
or UO_1042 (O_1042,N_9953,N_9826);
and UO_1043 (O_1043,N_9926,N_9938);
and UO_1044 (O_1044,N_9634,N_9747);
and UO_1045 (O_1045,N_9662,N_9553);
nor UO_1046 (O_1046,N_9696,N_9724);
and UO_1047 (O_1047,N_9905,N_9619);
nand UO_1048 (O_1048,N_9739,N_9873);
nand UO_1049 (O_1049,N_9740,N_9517);
and UO_1050 (O_1050,N_9917,N_9641);
or UO_1051 (O_1051,N_9635,N_9826);
nor UO_1052 (O_1052,N_9659,N_9723);
and UO_1053 (O_1053,N_9601,N_9769);
and UO_1054 (O_1054,N_9705,N_9990);
nand UO_1055 (O_1055,N_9753,N_9959);
or UO_1056 (O_1056,N_9577,N_9506);
nor UO_1057 (O_1057,N_9620,N_9731);
nand UO_1058 (O_1058,N_9801,N_9633);
nand UO_1059 (O_1059,N_9855,N_9500);
and UO_1060 (O_1060,N_9940,N_9911);
nor UO_1061 (O_1061,N_9979,N_9948);
nor UO_1062 (O_1062,N_9704,N_9807);
and UO_1063 (O_1063,N_9683,N_9799);
or UO_1064 (O_1064,N_9739,N_9901);
nand UO_1065 (O_1065,N_9601,N_9874);
or UO_1066 (O_1066,N_9743,N_9541);
or UO_1067 (O_1067,N_9745,N_9754);
or UO_1068 (O_1068,N_9532,N_9800);
nor UO_1069 (O_1069,N_9608,N_9823);
or UO_1070 (O_1070,N_9796,N_9881);
or UO_1071 (O_1071,N_9793,N_9879);
nor UO_1072 (O_1072,N_9862,N_9867);
nor UO_1073 (O_1073,N_9810,N_9523);
nor UO_1074 (O_1074,N_9604,N_9918);
nand UO_1075 (O_1075,N_9905,N_9998);
or UO_1076 (O_1076,N_9595,N_9808);
and UO_1077 (O_1077,N_9579,N_9822);
or UO_1078 (O_1078,N_9690,N_9888);
and UO_1079 (O_1079,N_9592,N_9946);
and UO_1080 (O_1080,N_9955,N_9665);
nor UO_1081 (O_1081,N_9773,N_9892);
and UO_1082 (O_1082,N_9913,N_9968);
nand UO_1083 (O_1083,N_9672,N_9780);
xnor UO_1084 (O_1084,N_9733,N_9948);
and UO_1085 (O_1085,N_9606,N_9924);
or UO_1086 (O_1086,N_9862,N_9629);
nor UO_1087 (O_1087,N_9894,N_9949);
nand UO_1088 (O_1088,N_9763,N_9775);
nor UO_1089 (O_1089,N_9660,N_9944);
and UO_1090 (O_1090,N_9835,N_9767);
nand UO_1091 (O_1091,N_9943,N_9832);
or UO_1092 (O_1092,N_9576,N_9517);
xnor UO_1093 (O_1093,N_9934,N_9552);
nor UO_1094 (O_1094,N_9687,N_9821);
or UO_1095 (O_1095,N_9947,N_9714);
xnor UO_1096 (O_1096,N_9538,N_9742);
nor UO_1097 (O_1097,N_9803,N_9705);
nor UO_1098 (O_1098,N_9954,N_9553);
or UO_1099 (O_1099,N_9695,N_9560);
nor UO_1100 (O_1100,N_9888,N_9790);
or UO_1101 (O_1101,N_9875,N_9772);
nand UO_1102 (O_1102,N_9731,N_9658);
nand UO_1103 (O_1103,N_9697,N_9586);
nor UO_1104 (O_1104,N_9503,N_9809);
nor UO_1105 (O_1105,N_9987,N_9695);
or UO_1106 (O_1106,N_9817,N_9791);
nand UO_1107 (O_1107,N_9968,N_9841);
or UO_1108 (O_1108,N_9650,N_9589);
xnor UO_1109 (O_1109,N_9919,N_9922);
nor UO_1110 (O_1110,N_9843,N_9910);
nor UO_1111 (O_1111,N_9854,N_9709);
xnor UO_1112 (O_1112,N_9833,N_9601);
nand UO_1113 (O_1113,N_9508,N_9512);
nor UO_1114 (O_1114,N_9825,N_9882);
or UO_1115 (O_1115,N_9760,N_9719);
and UO_1116 (O_1116,N_9828,N_9693);
or UO_1117 (O_1117,N_9613,N_9794);
nand UO_1118 (O_1118,N_9937,N_9897);
xnor UO_1119 (O_1119,N_9818,N_9815);
nor UO_1120 (O_1120,N_9830,N_9942);
nor UO_1121 (O_1121,N_9814,N_9632);
nor UO_1122 (O_1122,N_9823,N_9937);
and UO_1123 (O_1123,N_9787,N_9964);
or UO_1124 (O_1124,N_9679,N_9823);
nor UO_1125 (O_1125,N_9782,N_9842);
and UO_1126 (O_1126,N_9989,N_9793);
nand UO_1127 (O_1127,N_9934,N_9517);
nand UO_1128 (O_1128,N_9556,N_9838);
or UO_1129 (O_1129,N_9551,N_9916);
or UO_1130 (O_1130,N_9658,N_9799);
and UO_1131 (O_1131,N_9782,N_9583);
nor UO_1132 (O_1132,N_9830,N_9598);
or UO_1133 (O_1133,N_9813,N_9832);
nand UO_1134 (O_1134,N_9634,N_9502);
nor UO_1135 (O_1135,N_9586,N_9915);
and UO_1136 (O_1136,N_9651,N_9678);
xor UO_1137 (O_1137,N_9684,N_9695);
nor UO_1138 (O_1138,N_9745,N_9626);
or UO_1139 (O_1139,N_9719,N_9991);
and UO_1140 (O_1140,N_9501,N_9605);
nand UO_1141 (O_1141,N_9708,N_9810);
and UO_1142 (O_1142,N_9565,N_9733);
and UO_1143 (O_1143,N_9765,N_9939);
or UO_1144 (O_1144,N_9831,N_9888);
nand UO_1145 (O_1145,N_9961,N_9915);
or UO_1146 (O_1146,N_9764,N_9580);
nor UO_1147 (O_1147,N_9531,N_9605);
nand UO_1148 (O_1148,N_9587,N_9945);
and UO_1149 (O_1149,N_9779,N_9634);
or UO_1150 (O_1150,N_9931,N_9537);
or UO_1151 (O_1151,N_9785,N_9721);
nand UO_1152 (O_1152,N_9703,N_9995);
xnor UO_1153 (O_1153,N_9871,N_9990);
and UO_1154 (O_1154,N_9654,N_9534);
nor UO_1155 (O_1155,N_9689,N_9731);
or UO_1156 (O_1156,N_9805,N_9708);
nand UO_1157 (O_1157,N_9747,N_9502);
nand UO_1158 (O_1158,N_9634,N_9653);
nand UO_1159 (O_1159,N_9869,N_9769);
or UO_1160 (O_1160,N_9872,N_9843);
and UO_1161 (O_1161,N_9926,N_9687);
xor UO_1162 (O_1162,N_9732,N_9606);
nand UO_1163 (O_1163,N_9840,N_9865);
nand UO_1164 (O_1164,N_9764,N_9506);
nor UO_1165 (O_1165,N_9914,N_9790);
and UO_1166 (O_1166,N_9681,N_9612);
and UO_1167 (O_1167,N_9961,N_9761);
or UO_1168 (O_1168,N_9955,N_9535);
nor UO_1169 (O_1169,N_9880,N_9524);
or UO_1170 (O_1170,N_9515,N_9597);
nand UO_1171 (O_1171,N_9512,N_9567);
or UO_1172 (O_1172,N_9582,N_9995);
nor UO_1173 (O_1173,N_9640,N_9529);
and UO_1174 (O_1174,N_9722,N_9868);
and UO_1175 (O_1175,N_9823,N_9923);
and UO_1176 (O_1176,N_9784,N_9854);
and UO_1177 (O_1177,N_9540,N_9563);
nand UO_1178 (O_1178,N_9654,N_9828);
nor UO_1179 (O_1179,N_9570,N_9688);
or UO_1180 (O_1180,N_9774,N_9513);
nand UO_1181 (O_1181,N_9580,N_9639);
nand UO_1182 (O_1182,N_9740,N_9878);
nor UO_1183 (O_1183,N_9564,N_9894);
nor UO_1184 (O_1184,N_9715,N_9923);
and UO_1185 (O_1185,N_9706,N_9608);
nand UO_1186 (O_1186,N_9953,N_9836);
nand UO_1187 (O_1187,N_9506,N_9686);
nor UO_1188 (O_1188,N_9636,N_9934);
nor UO_1189 (O_1189,N_9508,N_9904);
or UO_1190 (O_1190,N_9925,N_9509);
nand UO_1191 (O_1191,N_9767,N_9731);
or UO_1192 (O_1192,N_9576,N_9500);
and UO_1193 (O_1193,N_9833,N_9961);
nor UO_1194 (O_1194,N_9947,N_9722);
or UO_1195 (O_1195,N_9647,N_9743);
and UO_1196 (O_1196,N_9964,N_9631);
or UO_1197 (O_1197,N_9913,N_9894);
or UO_1198 (O_1198,N_9659,N_9733);
or UO_1199 (O_1199,N_9606,N_9991);
and UO_1200 (O_1200,N_9911,N_9824);
or UO_1201 (O_1201,N_9846,N_9613);
nor UO_1202 (O_1202,N_9781,N_9766);
and UO_1203 (O_1203,N_9647,N_9679);
and UO_1204 (O_1204,N_9810,N_9899);
nor UO_1205 (O_1205,N_9528,N_9787);
and UO_1206 (O_1206,N_9795,N_9636);
nand UO_1207 (O_1207,N_9502,N_9674);
nor UO_1208 (O_1208,N_9879,N_9796);
xor UO_1209 (O_1209,N_9508,N_9782);
nand UO_1210 (O_1210,N_9982,N_9699);
or UO_1211 (O_1211,N_9976,N_9808);
and UO_1212 (O_1212,N_9815,N_9906);
xnor UO_1213 (O_1213,N_9803,N_9579);
or UO_1214 (O_1214,N_9716,N_9867);
nor UO_1215 (O_1215,N_9561,N_9984);
or UO_1216 (O_1216,N_9604,N_9853);
or UO_1217 (O_1217,N_9500,N_9671);
and UO_1218 (O_1218,N_9994,N_9705);
or UO_1219 (O_1219,N_9684,N_9884);
nand UO_1220 (O_1220,N_9526,N_9848);
or UO_1221 (O_1221,N_9744,N_9667);
nor UO_1222 (O_1222,N_9709,N_9642);
or UO_1223 (O_1223,N_9587,N_9844);
xor UO_1224 (O_1224,N_9968,N_9865);
or UO_1225 (O_1225,N_9995,N_9756);
and UO_1226 (O_1226,N_9631,N_9589);
and UO_1227 (O_1227,N_9770,N_9836);
and UO_1228 (O_1228,N_9561,N_9662);
nand UO_1229 (O_1229,N_9796,N_9706);
or UO_1230 (O_1230,N_9641,N_9709);
or UO_1231 (O_1231,N_9611,N_9995);
xnor UO_1232 (O_1232,N_9788,N_9667);
nand UO_1233 (O_1233,N_9638,N_9958);
and UO_1234 (O_1234,N_9828,N_9809);
nand UO_1235 (O_1235,N_9593,N_9994);
nor UO_1236 (O_1236,N_9992,N_9638);
and UO_1237 (O_1237,N_9602,N_9562);
nor UO_1238 (O_1238,N_9631,N_9537);
and UO_1239 (O_1239,N_9542,N_9781);
nor UO_1240 (O_1240,N_9727,N_9939);
nor UO_1241 (O_1241,N_9928,N_9761);
nor UO_1242 (O_1242,N_9873,N_9542);
nor UO_1243 (O_1243,N_9513,N_9963);
and UO_1244 (O_1244,N_9630,N_9653);
xnor UO_1245 (O_1245,N_9935,N_9835);
xor UO_1246 (O_1246,N_9920,N_9809);
nand UO_1247 (O_1247,N_9883,N_9581);
nor UO_1248 (O_1248,N_9815,N_9884);
nor UO_1249 (O_1249,N_9661,N_9576);
and UO_1250 (O_1250,N_9959,N_9690);
xnor UO_1251 (O_1251,N_9874,N_9852);
nand UO_1252 (O_1252,N_9761,N_9908);
nor UO_1253 (O_1253,N_9633,N_9725);
nand UO_1254 (O_1254,N_9917,N_9614);
nand UO_1255 (O_1255,N_9705,N_9788);
nor UO_1256 (O_1256,N_9784,N_9510);
nor UO_1257 (O_1257,N_9932,N_9929);
nor UO_1258 (O_1258,N_9571,N_9982);
nand UO_1259 (O_1259,N_9923,N_9813);
and UO_1260 (O_1260,N_9801,N_9541);
and UO_1261 (O_1261,N_9545,N_9963);
and UO_1262 (O_1262,N_9808,N_9758);
nand UO_1263 (O_1263,N_9868,N_9827);
and UO_1264 (O_1264,N_9649,N_9860);
or UO_1265 (O_1265,N_9560,N_9590);
xor UO_1266 (O_1266,N_9576,N_9508);
or UO_1267 (O_1267,N_9809,N_9843);
nand UO_1268 (O_1268,N_9651,N_9944);
and UO_1269 (O_1269,N_9562,N_9732);
and UO_1270 (O_1270,N_9684,N_9846);
nand UO_1271 (O_1271,N_9647,N_9889);
or UO_1272 (O_1272,N_9898,N_9723);
nand UO_1273 (O_1273,N_9662,N_9811);
or UO_1274 (O_1274,N_9996,N_9915);
nor UO_1275 (O_1275,N_9587,N_9775);
nand UO_1276 (O_1276,N_9747,N_9978);
or UO_1277 (O_1277,N_9933,N_9664);
xor UO_1278 (O_1278,N_9520,N_9604);
and UO_1279 (O_1279,N_9832,N_9558);
and UO_1280 (O_1280,N_9874,N_9659);
nand UO_1281 (O_1281,N_9912,N_9916);
or UO_1282 (O_1282,N_9634,N_9776);
nand UO_1283 (O_1283,N_9670,N_9510);
or UO_1284 (O_1284,N_9826,N_9685);
or UO_1285 (O_1285,N_9800,N_9828);
nand UO_1286 (O_1286,N_9641,N_9655);
xor UO_1287 (O_1287,N_9853,N_9548);
or UO_1288 (O_1288,N_9741,N_9947);
nor UO_1289 (O_1289,N_9518,N_9931);
nor UO_1290 (O_1290,N_9711,N_9804);
nand UO_1291 (O_1291,N_9912,N_9913);
or UO_1292 (O_1292,N_9636,N_9966);
xor UO_1293 (O_1293,N_9921,N_9752);
nand UO_1294 (O_1294,N_9764,N_9803);
nand UO_1295 (O_1295,N_9783,N_9587);
or UO_1296 (O_1296,N_9544,N_9953);
nor UO_1297 (O_1297,N_9502,N_9918);
xnor UO_1298 (O_1298,N_9689,N_9569);
or UO_1299 (O_1299,N_9794,N_9624);
xor UO_1300 (O_1300,N_9974,N_9530);
and UO_1301 (O_1301,N_9937,N_9954);
and UO_1302 (O_1302,N_9891,N_9721);
nor UO_1303 (O_1303,N_9808,N_9578);
or UO_1304 (O_1304,N_9838,N_9876);
and UO_1305 (O_1305,N_9913,N_9999);
and UO_1306 (O_1306,N_9707,N_9505);
xor UO_1307 (O_1307,N_9579,N_9553);
xnor UO_1308 (O_1308,N_9910,N_9680);
and UO_1309 (O_1309,N_9869,N_9981);
or UO_1310 (O_1310,N_9699,N_9895);
nand UO_1311 (O_1311,N_9625,N_9999);
and UO_1312 (O_1312,N_9518,N_9719);
nand UO_1313 (O_1313,N_9907,N_9654);
and UO_1314 (O_1314,N_9838,N_9887);
and UO_1315 (O_1315,N_9514,N_9851);
and UO_1316 (O_1316,N_9595,N_9888);
nor UO_1317 (O_1317,N_9987,N_9610);
or UO_1318 (O_1318,N_9784,N_9742);
and UO_1319 (O_1319,N_9862,N_9545);
nor UO_1320 (O_1320,N_9819,N_9724);
or UO_1321 (O_1321,N_9857,N_9543);
nand UO_1322 (O_1322,N_9860,N_9670);
nand UO_1323 (O_1323,N_9653,N_9715);
nor UO_1324 (O_1324,N_9962,N_9724);
and UO_1325 (O_1325,N_9898,N_9527);
nor UO_1326 (O_1326,N_9776,N_9690);
nor UO_1327 (O_1327,N_9844,N_9504);
or UO_1328 (O_1328,N_9540,N_9535);
xor UO_1329 (O_1329,N_9816,N_9748);
or UO_1330 (O_1330,N_9523,N_9873);
and UO_1331 (O_1331,N_9793,N_9578);
and UO_1332 (O_1332,N_9976,N_9737);
and UO_1333 (O_1333,N_9515,N_9603);
or UO_1334 (O_1334,N_9987,N_9917);
or UO_1335 (O_1335,N_9522,N_9741);
and UO_1336 (O_1336,N_9684,N_9578);
or UO_1337 (O_1337,N_9844,N_9808);
and UO_1338 (O_1338,N_9849,N_9807);
nand UO_1339 (O_1339,N_9655,N_9652);
and UO_1340 (O_1340,N_9853,N_9784);
nand UO_1341 (O_1341,N_9858,N_9622);
nand UO_1342 (O_1342,N_9704,N_9538);
xor UO_1343 (O_1343,N_9741,N_9560);
and UO_1344 (O_1344,N_9520,N_9646);
nand UO_1345 (O_1345,N_9531,N_9849);
nor UO_1346 (O_1346,N_9606,N_9961);
and UO_1347 (O_1347,N_9816,N_9828);
nand UO_1348 (O_1348,N_9841,N_9533);
xnor UO_1349 (O_1349,N_9543,N_9668);
nor UO_1350 (O_1350,N_9959,N_9857);
nor UO_1351 (O_1351,N_9996,N_9796);
nand UO_1352 (O_1352,N_9748,N_9549);
and UO_1353 (O_1353,N_9556,N_9866);
xor UO_1354 (O_1354,N_9667,N_9557);
and UO_1355 (O_1355,N_9604,N_9644);
and UO_1356 (O_1356,N_9769,N_9836);
and UO_1357 (O_1357,N_9775,N_9977);
and UO_1358 (O_1358,N_9814,N_9736);
nor UO_1359 (O_1359,N_9632,N_9924);
or UO_1360 (O_1360,N_9981,N_9776);
or UO_1361 (O_1361,N_9856,N_9776);
or UO_1362 (O_1362,N_9740,N_9715);
nor UO_1363 (O_1363,N_9753,N_9689);
or UO_1364 (O_1364,N_9839,N_9560);
xor UO_1365 (O_1365,N_9624,N_9790);
and UO_1366 (O_1366,N_9973,N_9831);
or UO_1367 (O_1367,N_9727,N_9635);
or UO_1368 (O_1368,N_9649,N_9533);
xnor UO_1369 (O_1369,N_9855,N_9681);
xnor UO_1370 (O_1370,N_9750,N_9514);
nor UO_1371 (O_1371,N_9889,N_9787);
nor UO_1372 (O_1372,N_9574,N_9718);
or UO_1373 (O_1373,N_9760,N_9906);
nand UO_1374 (O_1374,N_9935,N_9742);
nor UO_1375 (O_1375,N_9678,N_9983);
xnor UO_1376 (O_1376,N_9663,N_9768);
nand UO_1377 (O_1377,N_9931,N_9546);
or UO_1378 (O_1378,N_9716,N_9592);
and UO_1379 (O_1379,N_9724,N_9967);
xor UO_1380 (O_1380,N_9882,N_9785);
and UO_1381 (O_1381,N_9709,N_9501);
nand UO_1382 (O_1382,N_9511,N_9920);
and UO_1383 (O_1383,N_9650,N_9756);
and UO_1384 (O_1384,N_9584,N_9789);
and UO_1385 (O_1385,N_9901,N_9601);
nand UO_1386 (O_1386,N_9698,N_9753);
nand UO_1387 (O_1387,N_9987,N_9886);
and UO_1388 (O_1388,N_9699,N_9861);
nand UO_1389 (O_1389,N_9662,N_9744);
and UO_1390 (O_1390,N_9975,N_9806);
or UO_1391 (O_1391,N_9591,N_9709);
nor UO_1392 (O_1392,N_9701,N_9822);
and UO_1393 (O_1393,N_9859,N_9952);
xnor UO_1394 (O_1394,N_9651,N_9589);
and UO_1395 (O_1395,N_9915,N_9731);
and UO_1396 (O_1396,N_9781,N_9900);
and UO_1397 (O_1397,N_9943,N_9620);
or UO_1398 (O_1398,N_9819,N_9902);
and UO_1399 (O_1399,N_9960,N_9791);
nor UO_1400 (O_1400,N_9668,N_9872);
and UO_1401 (O_1401,N_9507,N_9616);
nor UO_1402 (O_1402,N_9655,N_9777);
nand UO_1403 (O_1403,N_9564,N_9905);
nor UO_1404 (O_1404,N_9779,N_9597);
and UO_1405 (O_1405,N_9746,N_9551);
and UO_1406 (O_1406,N_9894,N_9806);
nand UO_1407 (O_1407,N_9521,N_9774);
or UO_1408 (O_1408,N_9567,N_9504);
xor UO_1409 (O_1409,N_9559,N_9875);
xnor UO_1410 (O_1410,N_9542,N_9714);
nand UO_1411 (O_1411,N_9755,N_9726);
nand UO_1412 (O_1412,N_9548,N_9638);
nor UO_1413 (O_1413,N_9598,N_9809);
nand UO_1414 (O_1414,N_9729,N_9826);
nand UO_1415 (O_1415,N_9972,N_9927);
nor UO_1416 (O_1416,N_9605,N_9770);
and UO_1417 (O_1417,N_9888,N_9774);
nor UO_1418 (O_1418,N_9551,N_9943);
nor UO_1419 (O_1419,N_9679,N_9538);
nand UO_1420 (O_1420,N_9892,N_9811);
nor UO_1421 (O_1421,N_9993,N_9632);
nand UO_1422 (O_1422,N_9740,N_9884);
or UO_1423 (O_1423,N_9795,N_9747);
xor UO_1424 (O_1424,N_9509,N_9699);
and UO_1425 (O_1425,N_9782,N_9571);
nand UO_1426 (O_1426,N_9543,N_9787);
nand UO_1427 (O_1427,N_9835,N_9580);
nand UO_1428 (O_1428,N_9791,N_9605);
nand UO_1429 (O_1429,N_9796,N_9918);
nand UO_1430 (O_1430,N_9975,N_9592);
or UO_1431 (O_1431,N_9822,N_9527);
nand UO_1432 (O_1432,N_9874,N_9804);
nor UO_1433 (O_1433,N_9850,N_9539);
nand UO_1434 (O_1434,N_9790,N_9893);
nand UO_1435 (O_1435,N_9529,N_9757);
or UO_1436 (O_1436,N_9590,N_9798);
and UO_1437 (O_1437,N_9567,N_9631);
nand UO_1438 (O_1438,N_9820,N_9517);
and UO_1439 (O_1439,N_9948,N_9655);
nor UO_1440 (O_1440,N_9869,N_9506);
or UO_1441 (O_1441,N_9584,N_9667);
or UO_1442 (O_1442,N_9832,N_9823);
and UO_1443 (O_1443,N_9838,N_9985);
or UO_1444 (O_1444,N_9677,N_9894);
or UO_1445 (O_1445,N_9738,N_9921);
nand UO_1446 (O_1446,N_9801,N_9993);
or UO_1447 (O_1447,N_9513,N_9750);
nand UO_1448 (O_1448,N_9860,N_9595);
or UO_1449 (O_1449,N_9777,N_9788);
nand UO_1450 (O_1450,N_9912,N_9945);
nand UO_1451 (O_1451,N_9918,N_9999);
and UO_1452 (O_1452,N_9672,N_9688);
nand UO_1453 (O_1453,N_9921,N_9926);
and UO_1454 (O_1454,N_9729,N_9854);
or UO_1455 (O_1455,N_9650,N_9599);
and UO_1456 (O_1456,N_9714,N_9536);
xor UO_1457 (O_1457,N_9700,N_9668);
nand UO_1458 (O_1458,N_9832,N_9724);
nand UO_1459 (O_1459,N_9818,N_9700);
and UO_1460 (O_1460,N_9634,N_9937);
nand UO_1461 (O_1461,N_9560,N_9766);
nand UO_1462 (O_1462,N_9831,N_9930);
xnor UO_1463 (O_1463,N_9884,N_9658);
nand UO_1464 (O_1464,N_9715,N_9544);
or UO_1465 (O_1465,N_9714,N_9795);
nor UO_1466 (O_1466,N_9562,N_9712);
xor UO_1467 (O_1467,N_9823,N_9524);
nor UO_1468 (O_1468,N_9517,N_9661);
and UO_1469 (O_1469,N_9732,N_9704);
nand UO_1470 (O_1470,N_9667,N_9867);
or UO_1471 (O_1471,N_9933,N_9915);
nor UO_1472 (O_1472,N_9878,N_9767);
and UO_1473 (O_1473,N_9992,N_9776);
and UO_1474 (O_1474,N_9883,N_9943);
or UO_1475 (O_1475,N_9539,N_9953);
nand UO_1476 (O_1476,N_9856,N_9891);
nand UO_1477 (O_1477,N_9683,N_9500);
or UO_1478 (O_1478,N_9701,N_9823);
or UO_1479 (O_1479,N_9813,N_9583);
and UO_1480 (O_1480,N_9608,N_9880);
and UO_1481 (O_1481,N_9958,N_9507);
and UO_1482 (O_1482,N_9810,N_9690);
or UO_1483 (O_1483,N_9815,N_9655);
nor UO_1484 (O_1484,N_9652,N_9979);
or UO_1485 (O_1485,N_9732,N_9953);
or UO_1486 (O_1486,N_9791,N_9857);
nor UO_1487 (O_1487,N_9761,N_9634);
nand UO_1488 (O_1488,N_9518,N_9605);
nand UO_1489 (O_1489,N_9502,N_9607);
xnor UO_1490 (O_1490,N_9728,N_9677);
nor UO_1491 (O_1491,N_9848,N_9582);
and UO_1492 (O_1492,N_9680,N_9707);
xnor UO_1493 (O_1493,N_9689,N_9763);
nor UO_1494 (O_1494,N_9608,N_9939);
and UO_1495 (O_1495,N_9608,N_9978);
xor UO_1496 (O_1496,N_9827,N_9867);
and UO_1497 (O_1497,N_9714,N_9861);
nor UO_1498 (O_1498,N_9919,N_9974);
and UO_1499 (O_1499,N_9567,N_9901);
endmodule