module basic_1500_15000_2000_10_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_113,In_902);
and U1 (N_1,In_55,In_638);
or U2 (N_2,In_741,In_1451);
or U3 (N_3,In_691,In_947);
nor U4 (N_4,In_77,In_629);
xnor U5 (N_5,In_23,In_1);
nor U6 (N_6,In_361,In_402);
and U7 (N_7,In_129,In_447);
and U8 (N_8,In_207,In_1343);
or U9 (N_9,In_292,In_170);
nor U10 (N_10,In_556,In_1445);
nand U11 (N_11,In_1070,In_53);
nor U12 (N_12,In_731,In_824);
and U13 (N_13,In_637,In_1236);
and U14 (N_14,In_1361,In_503);
nor U15 (N_15,In_99,In_2);
and U16 (N_16,In_516,In_1217);
nand U17 (N_17,In_1219,In_359);
nand U18 (N_18,In_490,In_937);
xor U19 (N_19,In_1276,In_1313);
nand U20 (N_20,In_158,In_456);
and U21 (N_21,In_240,In_621);
xnor U22 (N_22,In_1179,In_1244);
and U23 (N_23,In_1087,In_1115);
nand U24 (N_24,In_585,In_1254);
nor U25 (N_25,In_524,In_1015);
nand U26 (N_26,In_1303,In_1443);
nand U27 (N_27,In_466,In_430);
xor U28 (N_28,In_438,In_460);
nor U29 (N_29,In_1129,In_215);
and U30 (N_30,In_1470,In_1337);
nor U31 (N_31,In_195,In_840);
and U32 (N_32,In_1142,In_242);
or U33 (N_33,In_308,In_174);
and U34 (N_34,In_198,In_1346);
nor U35 (N_35,In_718,In_832);
and U36 (N_36,In_111,In_1358);
or U37 (N_37,In_648,In_1101);
nor U38 (N_38,In_1274,In_385);
and U39 (N_39,In_1251,In_1357);
nor U40 (N_40,In_374,In_1355);
nand U41 (N_41,In_1237,In_462);
nand U42 (N_42,In_1222,In_1452);
nand U43 (N_43,In_1412,In_1292);
and U44 (N_44,In_507,In_1456);
or U45 (N_45,In_44,In_1260);
nand U46 (N_46,In_719,In_666);
and U47 (N_47,In_1160,In_246);
or U48 (N_48,In_1284,In_1110);
or U49 (N_49,In_802,In_543);
nand U50 (N_50,In_258,In_728);
nand U51 (N_51,In_310,In_189);
and U52 (N_52,In_1029,In_375);
and U53 (N_53,In_1293,In_508);
or U54 (N_54,In_997,In_378);
nand U55 (N_55,In_121,In_57);
nand U56 (N_56,In_150,In_674);
and U57 (N_57,In_1498,In_140);
or U58 (N_58,In_1130,In_283);
or U59 (N_59,In_297,In_326);
and U60 (N_60,In_572,In_67);
nor U61 (N_61,In_1095,In_749);
nand U62 (N_62,In_949,In_118);
and U63 (N_63,In_880,In_519);
or U64 (N_64,In_576,In_847);
nor U65 (N_65,In_311,In_155);
nand U66 (N_66,In_269,In_1282);
xor U67 (N_67,In_843,In_1050);
nor U68 (N_68,In_686,In_1479);
nand U69 (N_69,In_1442,In_1118);
and U70 (N_70,In_1281,In_38);
nor U71 (N_71,In_793,In_876);
nand U72 (N_72,In_397,In_1378);
and U73 (N_73,In_659,In_1288);
nand U74 (N_74,In_1255,In_1111);
nor U75 (N_75,In_608,In_935);
or U76 (N_76,In_9,In_914);
xnor U77 (N_77,In_325,In_722);
nand U78 (N_78,In_1128,In_881);
nor U79 (N_79,In_1194,In_603);
nand U80 (N_80,In_236,In_484);
nand U81 (N_81,In_336,In_681);
and U82 (N_82,In_833,In_328);
or U83 (N_83,In_882,In_509);
nand U84 (N_84,In_1472,In_231);
xnor U85 (N_85,In_1082,In_921);
nor U86 (N_86,In_227,In_829);
nor U87 (N_87,In_1403,In_281);
or U88 (N_88,In_262,In_748);
and U89 (N_89,In_126,In_967);
nor U90 (N_90,In_160,In_522);
or U91 (N_91,In_669,In_554);
nand U92 (N_92,In_293,In_321);
xnor U93 (N_93,In_106,In_1354);
nand U94 (N_94,In_134,In_1467);
and U95 (N_95,In_534,In_1259);
nor U96 (N_96,In_1060,In_774);
xnor U97 (N_97,In_738,In_151);
xor U98 (N_98,In_1027,In_750);
and U99 (N_99,In_1196,In_841);
nand U100 (N_100,In_785,In_1489);
nor U101 (N_101,In_998,In_428);
or U102 (N_102,In_379,In_1342);
nor U103 (N_103,In_1333,In_859);
xor U104 (N_104,In_354,In_517);
and U105 (N_105,In_600,In_999);
or U106 (N_106,In_414,In_973);
nor U107 (N_107,In_389,In_219);
and U108 (N_108,In_815,In_955);
nor U109 (N_109,In_795,In_499);
or U110 (N_110,In_756,In_1163);
nand U111 (N_111,In_1484,In_1113);
nand U112 (N_112,In_1409,In_980);
and U113 (N_113,In_651,In_1381);
and U114 (N_114,In_1065,In_768);
and U115 (N_115,In_1395,In_1102);
nor U116 (N_116,In_238,In_229);
or U117 (N_117,In_747,In_695);
nand U118 (N_118,In_527,In_458);
and U119 (N_119,In_510,In_230);
nand U120 (N_120,In_734,In_869);
nor U121 (N_121,In_333,In_1339);
or U122 (N_122,In_825,In_1450);
nor U123 (N_123,In_645,In_591);
and U124 (N_124,In_941,In_425);
xor U125 (N_125,In_1195,In_1324);
nor U126 (N_126,In_1422,In_184);
nor U127 (N_127,In_525,In_141);
xor U128 (N_128,In_604,In_1338);
nor U129 (N_129,In_237,In_888);
xor U130 (N_130,In_363,In_42);
xor U131 (N_131,In_294,In_1204);
and U132 (N_132,In_839,In_515);
nor U133 (N_133,In_1444,In_857);
and U134 (N_134,In_1143,In_1059);
xnor U135 (N_135,In_715,In_302);
and U136 (N_136,In_1134,In_551);
or U137 (N_137,In_900,In_1076);
and U138 (N_138,In_454,In_557);
nand U139 (N_139,In_301,In_1400);
nand U140 (N_140,In_1480,In_1038);
and U141 (N_141,In_1158,In_190);
or U142 (N_142,In_817,In_790);
and U143 (N_143,In_116,In_133);
nand U144 (N_144,In_1426,In_684);
and U145 (N_145,In_78,In_1225);
nand U146 (N_146,In_893,In_1345);
nand U147 (N_147,In_784,In_894);
nor U148 (N_148,In_1220,In_300);
nor U149 (N_149,In_1334,In_1249);
nand U150 (N_150,In_685,In_470);
nand U151 (N_151,In_982,In_1272);
and U152 (N_152,In_1265,In_1122);
nor U153 (N_153,In_930,In_214);
nor U154 (N_154,In_586,In_767);
nand U155 (N_155,In_612,In_675);
nor U156 (N_156,In_1298,In_271);
or U157 (N_157,In_419,In_306);
or U158 (N_158,In_1336,In_1148);
nor U159 (N_159,In_809,In_316);
and U160 (N_160,In_1019,In_1429);
nand U161 (N_161,In_210,In_948);
or U162 (N_162,In_1241,In_994);
nor U163 (N_163,In_779,In_26);
nor U164 (N_164,In_580,In_1018);
nor U165 (N_165,In_1235,In_979);
and U166 (N_166,In_1469,In_991);
nor U167 (N_167,In_186,In_746);
or U168 (N_168,In_459,In_1316);
or U169 (N_169,In_907,In_241);
nand U170 (N_170,In_878,In_777);
or U171 (N_171,In_1374,In_1407);
and U172 (N_172,In_661,In_593);
and U173 (N_173,In_1359,In_827);
or U174 (N_174,In_1210,In_69);
or U175 (N_175,In_495,In_916);
and U176 (N_176,In_1417,In_327);
or U177 (N_177,In_567,In_1205);
nor U178 (N_178,In_1414,In_1492);
and U179 (N_179,In_655,In_1040);
xnor U180 (N_180,In_698,In_1032);
or U181 (N_181,In_1197,In_234);
nor U182 (N_182,In_1155,In_701);
nor U183 (N_183,In_164,In_11);
nand U184 (N_184,In_1081,In_1003);
nand U185 (N_185,In_217,In_1362);
nand U186 (N_186,In_149,In_259);
nor U187 (N_187,In_745,In_71);
nand U188 (N_188,In_619,In_1151);
or U189 (N_189,In_533,In_114);
and U190 (N_190,In_1031,In_1493);
nor U191 (N_191,In_1043,In_555);
nand U192 (N_192,In_912,In_1476);
nor U193 (N_193,In_1468,In_200);
nor U194 (N_194,In_1089,In_176);
and U195 (N_195,In_920,In_399);
nor U196 (N_196,In_112,In_1256);
or U197 (N_197,In_532,In_1435);
or U198 (N_198,In_1030,In_319);
nand U199 (N_199,In_128,In_760);
or U200 (N_200,In_1137,In_971);
nor U201 (N_201,In_781,In_696);
or U202 (N_202,In_1080,In_432);
nor U203 (N_203,In_1014,In_423);
or U204 (N_204,In_906,In_1297);
nand U205 (N_205,In_773,In_1107);
nand U206 (N_206,In_547,In_1002);
nand U207 (N_207,In_1312,In_349);
nor U208 (N_208,In_1423,In_506);
and U209 (N_209,In_957,In_257);
or U210 (N_210,In_607,In_125);
and U211 (N_211,In_560,In_526);
or U212 (N_212,In_243,In_985);
nand U213 (N_213,In_1389,In_602);
nand U214 (N_214,In_411,In_1411);
nand U215 (N_215,In_183,In_1454);
nand U216 (N_216,In_1457,In_1329);
and U217 (N_217,In_1300,In_867);
and U218 (N_218,In_372,In_735);
nand U219 (N_219,In_280,In_1079);
nor U220 (N_220,In_435,In_1073);
nand U221 (N_221,In_27,In_305);
and U222 (N_222,In_1120,In_465);
nor U223 (N_223,In_928,In_729);
and U224 (N_224,In_670,In_248);
nand U225 (N_225,In_1286,In_52);
nand U226 (N_226,In_620,In_348);
nand U227 (N_227,In_1017,In_676);
nand U228 (N_228,In_384,In_537);
or U229 (N_229,In_961,In_1419);
and U230 (N_230,In_690,In_1275);
or U231 (N_231,In_886,In_418);
or U232 (N_232,In_171,In_1287);
nand U233 (N_233,In_513,In_594);
or U234 (N_234,In_1366,In_531);
nand U235 (N_235,In_889,In_1356);
and U236 (N_236,In_1352,In_960);
and U237 (N_237,In_1228,In_633);
and U238 (N_238,In_179,In_943);
and U239 (N_239,In_653,In_7);
xor U240 (N_240,In_1278,In_733);
or U241 (N_241,In_703,In_751);
xor U242 (N_242,In_613,In_1223);
nor U243 (N_243,In_660,In_765);
nor U244 (N_244,In_1415,In_107);
xor U245 (N_245,In_92,In_617);
and U246 (N_246,In_182,In_1152);
xnor U247 (N_247,In_650,In_426);
or U248 (N_248,In_964,In_75);
nand U249 (N_249,In_1104,In_1033);
and U250 (N_250,In_723,In_1035);
and U251 (N_251,In_954,In_712);
nand U252 (N_252,In_579,In_144);
nor U253 (N_253,In_628,In_1495);
and U254 (N_254,In_1238,In_481);
and U255 (N_255,In_656,In_521);
xor U256 (N_256,In_573,In_1126);
nand U257 (N_257,In_1091,In_958);
and U258 (N_258,In_1315,In_761);
nand U259 (N_259,In_119,In_331);
and U260 (N_260,In_1185,In_1135);
nand U261 (N_261,In_595,In_122);
xnor U262 (N_262,In_282,In_1174);
and U263 (N_263,In_202,In_687);
nand U264 (N_264,In_1474,In_1421);
nor U265 (N_265,In_1318,In_450);
and U266 (N_266,In_658,In_1264);
and U267 (N_267,In_1125,In_261);
or U268 (N_268,In_1216,In_911);
and U269 (N_269,In_1039,In_683);
nor U270 (N_270,In_1156,In_104);
and U271 (N_271,In_704,In_875);
nor U272 (N_272,In_714,In_463);
nor U273 (N_273,In_940,In_177);
or U274 (N_274,In_10,In_335);
or U275 (N_275,In_969,In_1436);
and U276 (N_276,In_1206,In_877);
or U277 (N_277,In_568,In_291);
nor U278 (N_278,In_864,In_1034);
and U279 (N_279,In_473,In_546);
or U280 (N_280,In_866,In_213);
or U281 (N_281,In_1092,In_918);
or U282 (N_282,In_870,In_1180);
nand U283 (N_283,In_887,In_853);
and U284 (N_284,In_216,In_501);
xnor U285 (N_285,In_1416,In_976);
or U286 (N_286,In_850,In_407);
xnor U287 (N_287,In_762,In_740);
and U288 (N_288,In_1392,In_1077);
nand U289 (N_289,In_1100,In_253);
nand U290 (N_290,In_1119,In_800);
or U291 (N_291,In_1046,In_461);
nand U292 (N_292,In_244,In_1116);
nand U293 (N_293,In_1384,In_1330);
nand U294 (N_294,In_845,In_185);
and U295 (N_295,In_791,In_1377);
or U296 (N_296,In_544,In_680);
nor U297 (N_297,In_1133,In_938);
nand U298 (N_298,In_946,In_156);
or U299 (N_299,In_1062,In_8);
xnor U300 (N_300,In_1103,In_1098);
or U301 (N_301,In_672,In_636);
and U302 (N_302,In_1273,In_159);
nand U303 (N_303,In_1383,In_341);
xnor U304 (N_304,In_285,In_356);
or U305 (N_305,In_373,In_288);
nor U306 (N_306,In_1042,In_480);
and U307 (N_307,In_1296,In_1289);
or U308 (N_308,In_175,In_491);
nand U309 (N_309,In_1227,In_381);
nand U310 (N_310,In_330,In_1351);
nand U311 (N_311,In_726,In_494);
nand U312 (N_312,In_347,In_564);
or U313 (N_313,In_449,In_1376);
nor U314 (N_314,In_266,In_1413);
nand U315 (N_315,In_102,In_706);
nor U316 (N_316,In_278,In_1008);
or U317 (N_317,In_816,In_996);
nor U318 (N_318,In_766,In_563);
nand U319 (N_319,In_96,In_1044);
or U320 (N_320,In_570,In_1386);
nor U321 (N_321,In_377,In_338);
nor U322 (N_322,In_1460,In_452);
nand U323 (N_323,In_1001,In_1475);
or U324 (N_324,In_689,In_1154);
and U325 (N_325,In_279,In_720);
and U326 (N_326,In_1406,In_788);
and U327 (N_327,In_60,In_694);
and U328 (N_328,In_1319,In_51);
or U329 (N_329,In_1370,In_1348);
or U330 (N_330,In_558,In_191);
or U331 (N_331,In_272,In_1487);
nand U332 (N_332,In_1139,In_298);
or U333 (N_333,In_181,In_624);
nand U334 (N_334,In_1149,In_172);
and U335 (N_335,In_623,In_32);
and U336 (N_336,In_754,In_865);
and U337 (N_337,In_482,In_844);
and U338 (N_338,In_1232,In_952);
and U339 (N_339,In_1314,In_0);
nor U340 (N_340,In_798,In_1153);
and U341 (N_341,In_422,In_108);
or U342 (N_342,In_1290,In_799);
or U343 (N_343,In_639,In_837);
and U344 (N_344,In_970,In_403);
or U345 (N_345,In_549,In_1162);
nor U346 (N_346,In_862,In_1307);
and U347 (N_347,In_367,In_1045);
and U348 (N_348,In_1064,In_1140);
or U349 (N_349,In_22,In_443);
and U350 (N_350,In_782,In_31);
nand U351 (N_351,In_1271,In_1369);
nor U352 (N_352,In_883,In_610);
nand U353 (N_353,In_1397,In_667);
or U354 (N_354,In_357,In_1323);
and U355 (N_355,In_1388,In_786);
or U356 (N_356,In_131,In_764);
or U357 (N_357,In_566,In_20);
and U358 (N_358,In_380,In_50);
nor U359 (N_359,In_1213,In_835);
or U360 (N_360,In_705,In_664);
and U361 (N_361,In_1047,In_487);
nand U362 (N_362,In_406,In_274);
nand U363 (N_363,In_1379,In_445);
nand U364 (N_364,In_950,In_673);
and U365 (N_365,In_700,In_1311);
or U366 (N_366,In_277,In_332);
nor U367 (N_367,In_863,In_153);
nor U368 (N_368,In_370,In_654);
or U369 (N_369,In_1215,In_929);
nor U370 (N_370,In_1071,In_1202);
nand U371 (N_371,In_437,In_1268);
xnor U372 (N_372,In_1173,In_197);
or U373 (N_373,In_1013,In_1067);
or U374 (N_374,In_1302,In_1327);
or U375 (N_375,In_529,In_255);
nand U376 (N_376,In_1418,In_1277);
nand U377 (N_377,In_632,In_987);
or U378 (N_378,In_471,In_169);
or U379 (N_379,In_74,In_369);
and U380 (N_380,In_1497,In_136);
and U381 (N_381,In_942,In_187);
nor U382 (N_382,In_431,In_590);
nand U383 (N_383,In_13,In_630);
and U384 (N_384,In_264,In_485);
nand U385 (N_385,In_646,In_662);
and U386 (N_386,In_404,In_993);
or U387 (N_387,In_858,In_1209);
and U388 (N_388,In_974,In_1446);
and U389 (N_389,In_100,In_1398);
nor U390 (N_390,In_605,In_752);
or U391 (N_391,In_1427,In_345);
nor U392 (N_392,In_1375,In_489);
or U393 (N_393,In_1471,In_1478);
or U394 (N_394,In_514,In_1437);
nand U395 (N_395,In_1431,In_1463);
nand U396 (N_396,In_220,In_5);
and U397 (N_397,In_80,In_296);
and U398 (N_398,In_45,In_1041);
and U399 (N_399,In_708,In_329);
xor U400 (N_400,In_1477,In_797);
and U401 (N_401,In_442,In_860);
nor U402 (N_402,In_1052,In_1161);
nand U403 (N_403,In_1069,In_73);
and U404 (N_404,In_351,In_364);
and U405 (N_405,In_625,In_1257);
nor U406 (N_406,In_205,In_956);
and U407 (N_407,In_127,In_193);
or U408 (N_408,In_771,In_981);
and U409 (N_409,In_1109,In_801);
nor U410 (N_410,In_1270,In_56);
xor U411 (N_411,In_309,In_39);
nor U412 (N_412,In_772,In_178);
xnor U413 (N_413,In_688,In_409);
and U414 (N_414,In_388,In_441);
and U415 (N_415,In_725,In_682);
nand U416 (N_416,In_416,In_753);
and U417 (N_417,In_317,In_523);
nand U418 (N_418,In_142,In_891);
or U419 (N_419,In_464,In_61);
nor U420 (N_420,In_87,In_1283);
and U421 (N_421,In_115,In_644);
nor U422 (N_422,In_469,In_989);
or U423 (N_423,In_842,In_834);
or U424 (N_424,In_545,In_201);
nand U425 (N_425,In_40,In_1121);
and U426 (N_426,In_1138,In_736);
and U427 (N_427,In_312,In_913);
and U428 (N_428,In_910,In_146);
xor U429 (N_429,In_717,In_939);
nor U430 (N_430,In_588,In_1198);
or U431 (N_431,In_4,In_826);
nand U432 (N_432,In_352,In_1306);
nand U433 (N_433,In_17,In_1368);
and U434 (N_434,In_440,In_211);
nor U435 (N_435,In_758,In_575);
nand U436 (N_436,In_631,In_1058);
xor U437 (N_437,In_247,In_713);
or U438 (N_438,In_854,In_344);
and U439 (N_439,In_16,In_355);
nor U440 (N_440,In_1165,In_538);
and U441 (N_441,In_1394,In_1176);
or U442 (N_442,In_1022,In_831);
or U443 (N_443,In_975,In_1072);
and U444 (N_444,In_697,In_420);
and U445 (N_445,In_1253,In_79);
and U446 (N_446,In_540,In_589);
nand U447 (N_447,In_615,In_1247);
nand U448 (N_448,In_830,In_43);
or U449 (N_449,In_596,In_41);
nand U450 (N_450,In_1186,In_35);
nor U451 (N_451,In_3,In_168);
or U452 (N_452,In_1168,In_1083);
and U453 (N_453,In_64,In_478);
and U454 (N_454,In_810,In_123);
nand U455 (N_455,In_1074,In_1150);
and U456 (N_456,In_770,In_1170);
nand U457 (N_457,In_1026,In_1230);
nand U458 (N_458,In_1136,In_143);
and U459 (N_459,In_897,In_265);
nand U460 (N_460,In_59,In_710);
nor U461 (N_461,In_977,In_535);
xnor U462 (N_462,In_1199,In_678);
and U463 (N_463,In_72,In_223);
and U464 (N_464,In_1234,In_665);
or U465 (N_465,In_1483,In_1499);
nand U466 (N_466,In_1169,In_598);
xnor U467 (N_467,In_86,In_587);
or U468 (N_468,In_36,In_1233);
and U469 (N_469,In_276,In_1016);
xnor U470 (N_470,In_1455,In_1240);
or U471 (N_471,In_390,In_368);
nor U472 (N_472,In_599,In_1491);
nand U473 (N_473,In_1433,In_899);
xnor U474 (N_474,In_256,In_304);
nor U475 (N_475,In_787,In_846);
nand U476 (N_476,In_1208,In_19);
nand U477 (N_477,In_157,In_789);
nand U478 (N_478,In_1490,In_1193);
and U479 (N_479,In_872,In_1299);
and U480 (N_480,In_836,In_1266);
nor U481 (N_481,In_14,In_28);
xor U482 (N_482,In_95,In_1360);
and U483 (N_483,In_393,In_320);
nor U484 (N_484,In_476,In_552);
nor U485 (N_485,In_933,In_1243);
and U486 (N_486,In_63,In_323);
nor U487 (N_487,In_417,In_192);
nor U488 (N_488,In_286,In_105);
nor U489 (N_489,In_83,In_1291);
nand U490 (N_490,In_926,In_1321);
or U491 (N_491,In_643,In_1239);
nand U492 (N_492,In_1305,In_1465);
nor U493 (N_493,In_315,In_353);
nand U494 (N_494,In_362,In_1448);
nor U495 (N_495,In_1211,In_565);
and U496 (N_496,In_421,In_1068);
nand U497 (N_497,In_1404,In_874);
nor U498 (N_498,In_436,In_467);
nand U499 (N_499,In_1063,In_1159);
or U500 (N_500,In_792,In_366);
nor U501 (N_501,In_709,In_763);
nor U502 (N_502,In_1353,In_931);
xnor U503 (N_503,In_135,In_1075);
or U504 (N_504,In_1494,In_822);
or U505 (N_505,In_744,In_635);
or U506 (N_506,In_995,In_1428);
nor U507 (N_507,In_505,In_601);
nor U508 (N_508,In_1410,In_1380);
nor U509 (N_509,In_249,In_821);
nor U510 (N_510,In_721,In_222);
or U511 (N_511,In_1112,In_562);
nand U512 (N_512,In_1310,In_1396);
xor U513 (N_513,In_1105,In_1117);
and U514 (N_514,In_1246,In_512);
xnor U515 (N_515,In_965,In_1371);
or U516 (N_516,In_455,In_502);
nand U517 (N_517,In_711,In_972);
or U518 (N_518,In_260,In_270);
xor U519 (N_519,In_70,In_818);
and U520 (N_520,In_945,In_702);
or U521 (N_521,In_21,In_1309);
nand U522 (N_522,In_959,In_885);
and U523 (N_523,In_475,In_1184);
nand U524 (N_524,In_769,In_203);
and U525 (N_525,In_371,In_427);
nand U526 (N_526,In_58,In_1004);
or U527 (N_527,In_1099,In_1365);
or U528 (N_528,In_84,In_923);
nor U529 (N_529,In_29,In_1261);
or U530 (N_530,In_439,In_559);
or U531 (N_531,In_34,In_103);
nand U532 (N_532,In_62,In_553);
or U533 (N_533,In_622,In_520);
nor U534 (N_534,In_268,In_641);
nor U535 (N_535,In_692,In_966);
nor U536 (N_536,In_152,In_1373);
nor U537 (N_537,In_88,In_429);
and U538 (N_538,In_915,In_1229);
nor U539 (N_539,In_1093,In_1024);
or U540 (N_540,In_1201,In_1326);
xnor U541 (N_541,In_1025,In_1191);
xor U542 (N_542,In_1363,In_1461);
or U543 (N_543,In_468,In_232);
xnor U544 (N_544,In_1123,In_879);
and U545 (N_545,In_303,In_161);
nor U546 (N_546,In_451,In_884);
xor U547 (N_547,In_1028,In_139);
and U548 (N_548,In_395,In_504);
or U549 (N_549,In_1399,In_343);
nor U550 (N_550,In_322,In_794);
and U551 (N_551,In_94,In_1057);
nand U552 (N_552,In_412,In_649);
xnor U553 (N_553,In_640,In_1007);
or U554 (N_554,In_97,In_1408);
or U555 (N_555,In_346,In_212);
or U556 (N_556,In_226,In_254);
nor U557 (N_557,In_1182,In_24);
and U558 (N_558,In_730,In_394);
nand U559 (N_559,In_273,In_896);
or U560 (N_560,In_851,In_805);
and U561 (N_561,In_365,In_1340);
or U562 (N_562,In_1012,In_609);
or U563 (N_563,In_627,In_909);
nand U564 (N_564,In_1245,In_1192);
nand U565 (N_565,In_614,In_196);
and U566 (N_566,In_1420,In_89);
or U567 (N_567,In_1382,In_235);
nor U568 (N_568,In_838,In_120);
nor U569 (N_569,In_1011,In_1224);
nand U570 (N_570,In_988,In_1485);
nor U571 (N_571,In_548,In_224);
and U572 (N_572,In_1294,In_1084);
or U573 (N_573,In_387,In_1486);
or U574 (N_574,In_814,In_511);
and U575 (N_575,In_1023,In_908);
nor U576 (N_576,In_1390,In_561);
nand U577 (N_577,In_1189,In_677);
xnor U578 (N_578,In_927,In_446);
nand U579 (N_579,In_1055,In_820);
nor U580 (N_580,In_1066,In_803);
xor U581 (N_581,In_811,In_386);
xor U582 (N_582,In_1335,In_204);
and U583 (N_583,In_1187,In_1258);
and U584 (N_584,In_1364,In_167);
nand U585 (N_585,In_616,In_1440);
and U586 (N_586,In_1488,In_1088);
or U587 (N_587,In_453,In_342);
nand U588 (N_588,In_1438,In_813);
and U589 (N_589,In_1037,In_457);
nand U590 (N_590,In_1464,In_1183);
and U591 (N_591,In_65,In_154);
or U592 (N_592,In_324,In_340);
xnor U593 (N_593,In_574,In_1021);
nand U594 (N_594,In_117,In_221);
nand U595 (N_595,In_1166,In_634);
nand U596 (N_596,In_334,In_1207);
nand U597 (N_597,In_924,In_990);
nor U598 (N_598,In_318,In_647);
xor U599 (N_599,In_919,In_162);
or U600 (N_600,In_147,In_433);
and U601 (N_601,In_1218,In_757);
or U602 (N_602,In_1226,In_1462);
nor U603 (N_603,In_932,In_1263);
or U604 (N_604,In_486,In_582);
nand U605 (N_605,In_1175,In_163);
and U606 (N_606,In_1006,In_299);
nand U607 (N_607,In_498,In_218);
nor U608 (N_608,In_1181,In_124);
or U609 (N_609,In_1020,In_1295);
or U610 (N_610,In_807,In_663);
nand U611 (N_611,In_951,In_37);
or U612 (N_612,In_295,In_1331);
or U613 (N_613,In_98,In_871);
nand U614 (N_614,In_925,In_500);
or U615 (N_615,In_1496,In_1106);
and U616 (N_616,In_1402,In_898);
nand U617 (N_617,In_1372,In_1350);
nand U618 (N_618,In_360,In_339);
or U619 (N_619,In_1203,In_6);
nor U620 (N_620,In_48,In_1393);
and U621 (N_621,In_1344,In_550);
nor U622 (N_622,In_1441,In_138);
nor U623 (N_623,In_109,In_652);
nor U624 (N_624,In_776,In_1332);
xor U625 (N_625,In_1061,In_1131);
or U626 (N_626,In_1177,In_1459);
xor U627 (N_627,In_759,In_1430);
or U628 (N_628,In_626,In_479);
nand U629 (N_629,In_1157,In_1434);
and U630 (N_630,In_130,In_1328);
and U631 (N_631,In_963,In_1250);
xnor U632 (N_632,In_1094,In_225);
nor U633 (N_633,In_166,In_448);
nand U634 (N_634,In_541,In_823);
nand U635 (N_635,In_33,In_496);
nand U636 (N_636,In_82,In_584);
xor U637 (N_637,In_1279,In_1096);
nand U638 (N_638,In_855,In_85);
or U639 (N_639,In_314,In_1048);
nor U640 (N_640,In_984,In_806);
nor U641 (N_641,In_693,In_1200);
nand U642 (N_642,In_542,In_780);
or U643 (N_643,In_424,In_778);
nor U644 (N_644,In_1304,In_890);
or U645 (N_645,In_400,In_434);
and U646 (N_646,In_410,In_1349);
nor U647 (N_647,In_1425,In_856);
and U648 (N_648,In_905,In_18);
nor U649 (N_649,In_868,In_199);
nand U650 (N_650,In_1301,In_1214);
nand U651 (N_651,In_1145,In_405);
or U652 (N_652,In_25,In_852);
and U653 (N_653,In_15,In_492);
xnor U654 (N_654,In_828,In_1171);
and U655 (N_655,In_992,In_383);
or U656 (N_656,In_1212,In_245);
and U657 (N_657,In_1449,In_1221);
nand U658 (N_658,In_250,In_1049);
or U659 (N_659,In_577,In_518);
nor U660 (N_660,In_583,In_101);
nand U661 (N_661,In_1391,In_284);
or U662 (N_662,In_901,In_148);
or U663 (N_663,In_986,In_699);
nor U664 (N_664,In_93,In_657);
or U665 (N_665,In_569,In_743);
nor U666 (N_666,In_861,In_1262);
xor U667 (N_667,In_1424,In_873);
or U668 (N_668,In_936,In_208);
nor U669 (N_669,In_1167,In_1124);
xnor U670 (N_670,In_707,In_90);
xor U671 (N_671,In_1188,In_165);
nor U672 (N_672,In_536,In_1447);
and U673 (N_673,In_739,In_1078);
nor U674 (N_674,In_1000,In_1252);
nand U675 (N_675,In_275,In_1127);
or U676 (N_676,In_1458,In_1347);
or U677 (N_677,In_1114,In_173);
and U678 (N_678,In_1325,In_1051);
nor U679 (N_679,In_983,In_727);
xor U680 (N_680,In_668,In_1320);
nor U681 (N_681,In_968,In_180);
or U682 (N_682,In_1308,In_1387);
or U683 (N_683,In_1280,In_1482);
and U684 (N_684,In_597,In_188);
and U685 (N_685,In_808,In_904);
and U686 (N_686,In_944,In_581);
nand U687 (N_687,In_953,In_1132);
or U688 (N_688,In_1036,In_194);
or U689 (N_689,In_1439,In_137);
nor U690 (N_690,In_396,In_290);
nand U691 (N_691,In_81,In_775);
xor U692 (N_692,In_978,In_1056);
nand U693 (N_693,In_472,In_350);
nand U694 (N_694,In_1146,In_724);
nor U695 (N_695,In_962,In_488);
or U696 (N_696,In_528,In_206);
nand U697 (N_697,In_1053,In_263);
and U698 (N_698,In_239,In_606);
nand U699 (N_699,In_642,In_1009);
nor U700 (N_700,In_1242,In_30);
or U701 (N_701,In_892,In_392);
or U702 (N_702,In_228,In_849);
nand U703 (N_703,In_1144,In_1269);
and U704 (N_704,In_1086,In_497);
and U705 (N_705,In_812,In_477);
or U706 (N_706,In_848,In_1401);
xnor U707 (N_707,In_1085,In_1466);
nor U708 (N_708,In_408,In_1097);
nand U709 (N_709,In_1147,In_66);
xnor U710 (N_710,In_12,In_267);
or U711 (N_711,In_611,In_917);
xnor U712 (N_712,In_1164,In_1010);
and U713 (N_713,In_1285,In_391);
nand U714 (N_714,In_755,In_307);
nor U715 (N_715,In_819,In_737);
xnor U716 (N_716,In_132,In_287);
or U717 (N_717,In_1172,In_618);
nand U718 (N_718,In_1453,In_91);
nor U719 (N_719,In_671,In_68);
or U720 (N_720,In_1108,In_679);
xnor U721 (N_721,In_1405,In_401);
nand U722 (N_722,In_804,In_251);
nand U723 (N_723,In_54,In_1317);
nand U724 (N_724,In_252,In_313);
nand U725 (N_725,In_233,In_145);
nor U726 (N_726,In_1322,In_796);
and U727 (N_727,In_49,In_1090);
nand U728 (N_728,In_415,In_1005);
and U729 (N_729,In_592,In_493);
nor U730 (N_730,In_1054,In_444);
or U731 (N_731,In_1367,In_732);
and U732 (N_732,In_1190,In_413);
and U733 (N_733,In_716,In_895);
and U734 (N_734,In_1481,In_110);
xor U735 (N_735,In_76,In_47);
or U736 (N_736,In_209,In_358);
nor U737 (N_737,In_1341,In_376);
or U738 (N_738,In_1385,In_474);
nor U739 (N_739,In_337,In_783);
nor U740 (N_740,In_1473,In_398);
nor U741 (N_741,In_1231,In_46);
nor U742 (N_742,In_530,In_539);
nand U743 (N_743,In_903,In_571);
or U744 (N_744,In_742,In_1248);
nor U745 (N_745,In_382,In_934);
xnor U746 (N_746,In_1267,In_1141);
nor U747 (N_747,In_578,In_1432);
nor U748 (N_748,In_483,In_922);
xor U749 (N_749,In_1178,In_289);
nor U750 (N_750,In_1476,In_538);
nand U751 (N_751,In_1087,In_1248);
nor U752 (N_752,In_1446,In_697);
nor U753 (N_753,In_193,In_666);
xor U754 (N_754,In_832,In_110);
or U755 (N_755,In_905,In_1353);
or U756 (N_756,In_974,In_1003);
nor U757 (N_757,In_535,In_164);
or U758 (N_758,In_341,In_1018);
xnor U759 (N_759,In_425,In_1377);
nand U760 (N_760,In_1073,In_860);
nand U761 (N_761,In_403,In_726);
and U762 (N_762,In_640,In_662);
nor U763 (N_763,In_1155,In_924);
nand U764 (N_764,In_1139,In_348);
and U765 (N_765,In_903,In_1466);
nand U766 (N_766,In_93,In_235);
nand U767 (N_767,In_566,In_450);
nor U768 (N_768,In_558,In_51);
xnor U769 (N_769,In_1184,In_1302);
nor U770 (N_770,In_1099,In_238);
or U771 (N_771,In_701,In_791);
or U772 (N_772,In_874,In_402);
or U773 (N_773,In_774,In_1096);
nand U774 (N_774,In_1267,In_1445);
nor U775 (N_775,In_1234,In_88);
nand U776 (N_776,In_1174,In_711);
nor U777 (N_777,In_783,In_407);
nor U778 (N_778,In_643,In_777);
nand U779 (N_779,In_125,In_366);
and U780 (N_780,In_79,In_169);
and U781 (N_781,In_1242,In_617);
nor U782 (N_782,In_190,In_338);
xnor U783 (N_783,In_404,In_925);
and U784 (N_784,In_509,In_1048);
xor U785 (N_785,In_674,In_1359);
nand U786 (N_786,In_1193,In_136);
nand U787 (N_787,In_1258,In_1246);
nor U788 (N_788,In_523,In_1002);
and U789 (N_789,In_264,In_602);
and U790 (N_790,In_1075,In_609);
nor U791 (N_791,In_1373,In_1005);
and U792 (N_792,In_399,In_370);
nor U793 (N_793,In_1419,In_657);
nor U794 (N_794,In_1208,In_188);
nor U795 (N_795,In_983,In_1318);
or U796 (N_796,In_212,In_799);
and U797 (N_797,In_1436,In_89);
and U798 (N_798,In_99,In_57);
nand U799 (N_799,In_724,In_1264);
or U800 (N_800,In_1471,In_736);
or U801 (N_801,In_1400,In_170);
nand U802 (N_802,In_6,In_933);
and U803 (N_803,In_297,In_1143);
nand U804 (N_804,In_1380,In_1450);
nor U805 (N_805,In_979,In_463);
nand U806 (N_806,In_1179,In_467);
nand U807 (N_807,In_1324,In_462);
nand U808 (N_808,In_1055,In_1415);
nor U809 (N_809,In_618,In_829);
and U810 (N_810,In_1457,In_1474);
or U811 (N_811,In_618,In_360);
nand U812 (N_812,In_622,In_465);
nor U813 (N_813,In_666,In_489);
and U814 (N_814,In_347,In_252);
or U815 (N_815,In_1254,In_1318);
nand U816 (N_816,In_342,In_329);
nand U817 (N_817,In_100,In_538);
xor U818 (N_818,In_1096,In_637);
or U819 (N_819,In_1302,In_110);
nand U820 (N_820,In_1407,In_579);
nand U821 (N_821,In_845,In_738);
xor U822 (N_822,In_959,In_1143);
or U823 (N_823,In_203,In_1389);
or U824 (N_824,In_621,In_1494);
and U825 (N_825,In_1252,In_513);
xnor U826 (N_826,In_726,In_1467);
or U827 (N_827,In_452,In_1413);
and U828 (N_828,In_284,In_1124);
nand U829 (N_829,In_1223,In_790);
nor U830 (N_830,In_1076,In_169);
or U831 (N_831,In_1268,In_115);
or U832 (N_832,In_680,In_317);
nor U833 (N_833,In_1080,In_263);
nand U834 (N_834,In_1382,In_1053);
or U835 (N_835,In_1492,In_701);
and U836 (N_836,In_262,In_792);
and U837 (N_837,In_937,In_1216);
and U838 (N_838,In_1294,In_484);
or U839 (N_839,In_287,In_1451);
xnor U840 (N_840,In_48,In_162);
xor U841 (N_841,In_1178,In_771);
or U842 (N_842,In_286,In_694);
nand U843 (N_843,In_473,In_572);
nand U844 (N_844,In_322,In_1405);
xor U845 (N_845,In_1170,In_1295);
xor U846 (N_846,In_235,In_1);
xor U847 (N_847,In_609,In_1280);
or U848 (N_848,In_143,In_738);
or U849 (N_849,In_1433,In_887);
nand U850 (N_850,In_264,In_171);
nor U851 (N_851,In_1349,In_816);
and U852 (N_852,In_1173,In_782);
or U853 (N_853,In_893,In_179);
or U854 (N_854,In_98,In_41);
nor U855 (N_855,In_1470,In_771);
or U856 (N_856,In_634,In_467);
nor U857 (N_857,In_1107,In_600);
nor U858 (N_858,In_1057,In_1238);
or U859 (N_859,In_1298,In_808);
and U860 (N_860,In_1219,In_1078);
xnor U861 (N_861,In_441,In_1234);
and U862 (N_862,In_1366,In_814);
and U863 (N_863,In_1119,In_261);
xnor U864 (N_864,In_533,In_585);
nand U865 (N_865,In_674,In_590);
and U866 (N_866,In_689,In_509);
or U867 (N_867,In_604,In_265);
nor U868 (N_868,In_1421,In_1312);
nor U869 (N_869,In_1281,In_1099);
nor U870 (N_870,In_1207,In_504);
nand U871 (N_871,In_1282,In_1284);
or U872 (N_872,In_1124,In_391);
and U873 (N_873,In_857,In_541);
nand U874 (N_874,In_1392,In_80);
xnor U875 (N_875,In_1173,In_837);
or U876 (N_876,In_1346,In_340);
nand U877 (N_877,In_1145,In_1371);
or U878 (N_878,In_1124,In_633);
nand U879 (N_879,In_527,In_1426);
xor U880 (N_880,In_1025,In_438);
nor U881 (N_881,In_1295,In_423);
or U882 (N_882,In_1454,In_925);
and U883 (N_883,In_1295,In_1002);
nand U884 (N_884,In_1012,In_1485);
or U885 (N_885,In_169,In_122);
nor U886 (N_886,In_577,In_586);
and U887 (N_887,In_415,In_815);
nand U888 (N_888,In_151,In_460);
and U889 (N_889,In_1359,In_1298);
and U890 (N_890,In_997,In_1121);
and U891 (N_891,In_113,In_532);
nor U892 (N_892,In_538,In_1271);
nor U893 (N_893,In_1226,In_479);
and U894 (N_894,In_976,In_896);
xnor U895 (N_895,In_524,In_1230);
nor U896 (N_896,In_770,In_674);
nor U897 (N_897,In_9,In_343);
and U898 (N_898,In_1075,In_1015);
nor U899 (N_899,In_1071,In_492);
nand U900 (N_900,In_1385,In_1223);
nand U901 (N_901,In_195,In_58);
or U902 (N_902,In_422,In_1273);
nand U903 (N_903,In_460,In_369);
nand U904 (N_904,In_1041,In_842);
or U905 (N_905,In_580,In_273);
and U906 (N_906,In_877,In_1084);
nand U907 (N_907,In_755,In_934);
and U908 (N_908,In_1318,In_1437);
xor U909 (N_909,In_714,In_1064);
nand U910 (N_910,In_1235,In_1387);
or U911 (N_911,In_102,In_882);
nor U912 (N_912,In_574,In_772);
and U913 (N_913,In_1284,In_1115);
and U914 (N_914,In_85,In_1469);
nor U915 (N_915,In_290,In_399);
nand U916 (N_916,In_616,In_153);
or U917 (N_917,In_967,In_1186);
nor U918 (N_918,In_1393,In_402);
and U919 (N_919,In_320,In_681);
nor U920 (N_920,In_905,In_1098);
nand U921 (N_921,In_427,In_134);
xor U922 (N_922,In_724,In_426);
xnor U923 (N_923,In_1080,In_492);
nor U924 (N_924,In_89,In_1460);
nor U925 (N_925,In_1143,In_1413);
nand U926 (N_926,In_1304,In_248);
nor U927 (N_927,In_1215,In_792);
nand U928 (N_928,In_88,In_230);
nand U929 (N_929,In_798,In_218);
nor U930 (N_930,In_55,In_77);
nand U931 (N_931,In_243,In_812);
nand U932 (N_932,In_35,In_895);
nand U933 (N_933,In_1021,In_582);
nor U934 (N_934,In_986,In_1099);
nand U935 (N_935,In_282,In_890);
nand U936 (N_936,In_634,In_946);
or U937 (N_937,In_223,In_608);
and U938 (N_938,In_336,In_718);
or U939 (N_939,In_358,In_1023);
nor U940 (N_940,In_1289,In_1273);
xor U941 (N_941,In_588,In_15);
or U942 (N_942,In_237,In_25);
xnor U943 (N_943,In_47,In_1046);
nor U944 (N_944,In_35,In_266);
and U945 (N_945,In_773,In_61);
and U946 (N_946,In_827,In_1043);
and U947 (N_947,In_1206,In_820);
and U948 (N_948,In_1211,In_893);
nor U949 (N_949,In_369,In_1018);
nor U950 (N_950,In_587,In_909);
and U951 (N_951,In_18,In_388);
or U952 (N_952,In_234,In_798);
or U953 (N_953,In_34,In_100);
nor U954 (N_954,In_521,In_122);
nor U955 (N_955,In_651,In_1288);
nor U956 (N_956,In_294,In_1279);
nand U957 (N_957,In_710,In_1026);
xor U958 (N_958,In_1468,In_88);
and U959 (N_959,In_173,In_1481);
nor U960 (N_960,In_230,In_453);
nand U961 (N_961,In_357,In_1078);
or U962 (N_962,In_306,In_695);
and U963 (N_963,In_1205,In_18);
xnor U964 (N_964,In_1315,In_773);
nand U965 (N_965,In_1062,In_1222);
nor U966 (N_966,In_555,In_147);
or U967 (N_967,In_507,In_372);
xnor U968 (N_968,In_1214,In_630);
and U969 (N_969,In_857,In_167);
or U970 (N_970,In_1018,In_560);
xor U971 (N_971,In_1089,In_801);
nor U972 (N_972,In_1123,In_592);
and U973 (N_973,In_1302,In_601);
nand U974 (N_974,In_764,In_189);
nand U975 (N_975,In_361,In_1410);
or U976 (N_976,In_983,In_745);
and U977 (N_977,In_1142,In_1023);
nand U978 (N_978,In_961,In_1375);
nor U979 (N_979,In_1338,In_323);
and U980 (N_980,In_931,In_309);
nor U981 (N_981,In_772,In_518);
and U982 (N_982,In_294,In_705);
nor U983 (N_983,In_1254,In_637);
and U984 (N_984,In_243,In_503);
nor U985 (N_985,In_160,In_1463);
nand U986 (N_986,In_243,In_1293);
and U987 (N_987,In_1229,In_416);
xor U988 (N_988,In_846,In_1363);
and U989 (N_989,In_781,In_1405);
xnor U990 (N_990,In_107,In_820);
nand U991 (N_991,In_426,In_33);
nor U992 (N_992,In_1302,In_1038);
xnor U993 (N_993,In_1202,In_605);
nor U994 (N_994,In_516,In_548);
or U995 (N_995,In_1337,In_67);
or U996 (N_996,In_769,In_693);
xnor U997 (N_997,In_514,In_1152);
nand U998 (N_998,In_168,In_1004);
nand U999 (N_999,In_1031,In_1477);
nor U1000 (N_1000,In_693,In_235);
nor U1001 (N_1001,In_0,In_1307);
nand U1002 (N_1002,In_390,In_146);
nor U1003 (N_1003,In_924,In_480);
and U1004 (N_1004,In_984,In_417);
or U1005 (N_1005,In_841,In_567);
nor U1006 (N_1006,In_1216,In_933);
nand U1007 (N_1007,In_763,In_224);
or U1008 (N_1008,In_848,In_1269);
and U1009 (N_1009,In_385,In_145);
nor U1010 (N_1010,In_631,In_890);
nor U1011 (N_1011,In_1472,In_678);
and U1012 (N_1012,In_301,In_537);
and U1013 (N_1013,In_892,In_1288);
or U1014 (N_1014,In_26,In_1327);
nor U1015 (N_1015,In_171,In_892);
and U1016 (N_1016,In_1464,In_431);
nor U1017 (N_1017,In_1040,In_316);
nor U1018 (N_1018,In_33,In_1444);
nand U1019 (N_1019,In_932,In_204);
xnor U1020 (N_1020,In_1099,In_989);
nor U1021 (N_1021,In_1371,In_1205);
nor U1022 (N_1022,In_1356,In_67);
and U1023 (N_1023,In_673,In_880);
nor U1024 (N_1024,In_778,In_399);
nor U1025 (N_1025,In_728,In_51);
nand U1026 (N_1026,In_956,In_1011);
nor U1027 (N_1027,In_335,In_1494);
or U1028 (N_1028,In_687,In_1112);
or U1029 (N_1029,In_639,In_1394);
and U1030 (N_1030,In_461,In_833);
nor U1031 (N_1031,In_1066,In_994);
or U1032 (N_1032,In_517,In_1399);
nand U1033 (N_1033,In_1383,In_1387);
nand U1034 (N_1034,In_314,In_363);
or U1035 (N_1035,In_1290,In_397);
nor U1036 (N_1036,In_473,In_1259);
nor U1037 (N_1037,In_1393,In_109);
nand U1038 (N_1038,In_1116,In_1239);
nand U1039 (N_1039,In_1111,In_446);
nand U1040 (N_1040,In_524,In_64);
nor U1041 (N_1041,In_302,In_99);
nor U1042 (N_1042,In_811,In_992);
xor U1043 (N_1043,In_518,In_1050);
nor U1044 (N_1044,In_557,In_1270);
and U1045 (N_1045,In_317,In_919);
nor U1046 (N_1046,In_491,In_257);
or U1047 (N_1047,In_499,In_636);
nand U1048 (N_1048,In_865,In_1492);
nand U1049 (N_1049,In_1384,In_1492);
and U1050 (N_1050,In_63,In_385);
xnor U1051 (N_1051,In_960,In_790);
nor U1052 (N_1052,In_552,In_1469);
xor U1053 (N_1053,In_1426,In_328);
nand U1054 (N_1054,In_212,In_1222);
nand U1055 (N_1055,In_560,In_235);
and U1056 (N_1056,In_269,In_498);
or U1057 (N_1057,In_560,In_144);
or U1058 (N_1058,In_719,In_876);
or U1059 (N_1059,In_273,In_76);
nand U1060 (N_1060,In_274,In_367);
nand U1061 (N_1061,In_1007,In_233);
xnor U1062 (N_1062,In_109,In_430);
nand U1063 (N_1063,In_1474,In_689);
and U1064 (N_1064,In_904,In_569);
and U1065 (N_1065,In_633,In_913);
or U1066 (N_1066,In_518,In_189);
nor U1067 (N_1067,In_1375,In_1489);
or U1068 (N_1068,In_835,In_30);
nor U1069 (N_1069,In_1454,In_1210);
xor U1070 (N_1070,In_252,In_75);
and U1071 (N_1071,In_306,In_685);
nand U1072 (N_1072,In_1388,In_503);
nor U1073 (N_1073,In_307,In_612);
and U1074 (N_1074,In_167,In_699);
nand U1075 (N_1075,In_873,In_789);
or U1076 (N_1076,In_936,In_981);
and U1077 (N_1077,In_360,In_281);
nand U1078 (N_1078,In_323,In_1013);
nand U1079 (N_1079,In_708,In_468);
or U1080 (N_1080,In_581,In_684);
and U1081 (N_1081,In_15,In_1018);
or U1082 (N_1082,In_593,In_12);
or U1083 (N_1083,In_181,In_197);
and U1084 (N_1084,In_179,In_711);
nor U1085 (N_1085,In_1143,In_1069);
xor U1086 (N_1086,In_1107,In_139);
nor U1087 (N_1087,In_982,In_1379);
and U1088 (N_1088,In_1110,In_1305);
nor U1089 (N_1089,In_595,In_36);
xor U1090 (N_1090,In_745,In_1096);
nand U1091 (N_1091,In_1203,In_1238);
or U1092 (N_1092,In_14,In_1221);
nand U1093 (N_1093,In_699,In_1029);
and U1094 (N_1094,In_896,In_817);
nor U1095 (N_1095,In_1275,In_266);
and U1096 (N_1096,In_1060,In_530);
nand U1097 (N_1097,In_539,In_625);
xor U1098 (N_1098,In_811,In_516);
or U1099 (N_1099,In_1026,In_1297);
xnor U1100 (N_1100,In_600,In_378);
and U1101 (N_1101,In_53,In_992);
and U1102 (N_1102,In_901,In_1378);
and U1103 (N_1103,In_580,In_1440);
and U1104 (N_1104,In_467,In_894);
xnor U1105 (N_1105,In_622,In_1033);
and U1106 (N_1106,In_877,In_1102);
or U1107 (N_1107,In_928,In_339);
or U1108 (N_1108,In_63,In_1291);
nor U1109 (N_1109,In_1276,In_216);
nand U1110 (N_1110,In_1216,In_120);
nor U1111 (N_1111,In_891,In_719);
xor U1112 (N_1112,In_1220,In_152);
or U1113 (N_1113,In_1144,In_1336);
and U1114 (N_1114,In_764,In_642);
nor U1115 (N_1115,In_333,In_888);
nand U1116 (N_1116,In_9,In_122);
nand U1117 (N_1117,In_412,In_602);
and U1118 (N_1118,In_1185,In_1207);
and U1119 (N_1119,In_163,In_421);
or U1120 (N_1120,In_315,In_152);
nand U1121 (N_1121,In_132,In_248);
nor U1122 (N_1122,In_1238,In_1230);
xor U1123 (N_1123,In_1462,In_69);
nor U1124 (N_1124,In_827,In_1006);
nor U1125 (N_1125,In_881,In_1472);
and U1126 (N_1126,In_1241,In_1168);
or U1127 (N_1127,In_147,In_136);
or U1128 (N_1128,In_644,In_256);
nor U1129 (N_1129,In_68,In_236);
xor U1130 (N_1130,In_1002,In_439);
nor U1131 (N_1131,In_1476,In_874);
and U1132 (N_1132,In_721,In_719);
and U1133 (N_1133,In_604,In_322);
nand U1134 (N_1134,In_472,In_1323);
or U1135 (N_1135,In_1239,In_1299);
or U1136 (N_1136,In_1397,In_22);
and U1137 (N_1137,In_998,In_169);
or U1138 (N_1138,In_1295,In_1407);
and U1139 (N_1139,In_824,In_1298);
and U1140 (N_1140,In_801,In_846);
nor U1141 (N_1141,In_538,In_859);
and U1142 (N_1142,In_1036,In_1097);
nor U1143 (N_1143,In_771,In_781);
and U1144 (N_1144,In_500,In_284);
or U1145 (N_1145,In_28,In_618);
xnor U1146 (N_1146,In_1476,In_1295);
nand U1147 (N_1147,In_212,In_1291);
nor U1148 (N_1148,In_205,In_681);
nand U1149 (N_1149,In_159,In_1424);
xor U1150 (N_1150,In_376,In_1072);
nand U1151 (N_1151,In_1059,In_1468);
nand U1152 (N_1152,In_1061,In_1221);
nor U1153 (N_1153,In_896,In_1171);
and U1154 (N_1154,In_1318,In_355);
nand U1155 (N_1155,In_72,In_444);
nand U1156 (N_1156,In_1039,In_79);
nor U1157 (N_1157,In_71,In_1127);
nand U1158 (N_1158,In_47,In_123);
and U1159 (N_1159,In_354,In_1213);
nand U1160 (N_1160,In_898,In_214);
nand U1161 (N_1161,In_22,In_699);
or U1162 (N_1162,In_804,In_779);
nor U1163 (N_1163,In_1411,In_254);
nor U1164 (N_1164,In_1171,In_995);
nor U1165 (N_1165,In_355,In_136);
xnor U1166 (N_1166,In_135,In_1041);
or U1167 (N_1167,In_171,In_519);
nand U1168 (N_1168,In_772,In_94);
or U1169 (N_1169,In_1397,In_234);
or U1170 (N_1170,In_341,In_930);
and U1171 (N_1171,In_603,In_227);
nand U1172 (N_1172,In_681,In_427);
nand U1173 (N_1173,In_1040,In_581);
nor U1174 (N_1174,In_21,In_1272);
and U1175 (N_1175,In_1308,In_1338);
nor U1176 (N_1176,In_50,In_1357);
and U1177 (N_1177,In_904,In_1120);
and U1178 (N_1178,In_606,In_657);
or U1179 (N_1179,In_775,In_518);
or U1180 (N_1180,In_712,In_470);
and U1181 (N_1181,In_1368,In_1251);
nand U1182 (N_1182,In_1421,In_1226);
nand U1183 (N_1183,In_385,In_1247);
nand U1184 (N_1184,In_148,In_1194);
nand U1185 (N_1185,In_465,In_1327);
nor U1186 (N_1186,In_967,In_537);
xor U1187 (N_1187,In_95,In_418);
or U1188 (N_1188,In_1357,In_1205);
nand U1189 (N_1189,In_1047,In_194);
xor U1190 (N_1190,In_217,In_1078);
and U1191 (N_1191,In_643,In_1224);
nor U1192 (N_1192,In_642,In_1467);
nand U1193 (N_1193,In_176,In_897);
xor U1194 (N_1194,In_421,In_261);
xor U1195 (N_1195,In_924,In_751);
nand U1196 (N_1196,In_928,In_1220);
nand U1197 (N_1197,In_845,In_439);
nor U1198 (N_1198,In_585,In_1074);
nand U1199 (N_1199,In_849,In_29);
or U1200 (N_1200,In_354,In_1282);
nor U1201 (N_1201,In_293,In_104);
nand U1202 (N_1202,In_90,In_10);
xor U1203 (N_1203,In_1122,In_634);
nor U1204 (N_1204,In_985,In_859);
nand U1205 (N_1205,In_362,In_708);
nor U1206 (N_1206,In_822,In_323);
and U1207 (N_1207,In_1024,In_1451);
or U1208 (N_1208,In_1342,In_406);
nor U1209 (N_1209,In_1093,In_628);
nand U1210 (N_1210,In_28,In_144);
nor U1211 (N_1211,In_922,In_995);
nand U1212 (N_1212,In_62,In_294);
nor U1213 (N_1213,In_410,In_367);
xor U1214 (N_1214,In_331,In_230);
and U1215 (N_1215,In_145,In_1075);
nand U1216 (N_1216,In_689,In_597);
nand U1217 (N_1217,In_449,In_1444);
or U1218 (N_1218,In_700,In_1286);
or U1219 (N_1219,In_1322,In_1032);
nor U1220 (N_1220,In_82,In_123);
or U1221 (N_1221,In_1463,In_838);
nand U1222 (N_1222,In_877,In_425);
or U1223 (N_1223,In_516,In_723);
nand U1224 (N_1224,In_269,In_788);
nor U1225 (N_1225,In_817,In_1189);
nand U1226 (N_1226,In_1051,In_936);
and U1227 (N_1227,In_1124,In_795);
xnor U1228 (N_1228,In_1410,In_417);
and U1229 (N_1229,In_163,In_664);
and U1230 (N_1230,In_478,In_367);
nand U1231 (N_1231,In_1095,In_488);
nor U1232 (N_1232,In_1448,In_1179);
or U1233 (N_1233,In_288,In_1092);
and U1234 (N_1234,In_1164,In_569);
or U1235 (N_1235,In_11,In_185);
nand U1236 (N_1236,In_327,In_864);
nand U1237 (N_1237,In_1378,In_1459);
nor U1238 (N_1238,In_723,In_107);
or U1239 (N_1239,In_132,In_233);
and U1240 (N_1240,In_750,In_929);
and U1241 (N_1241,In_1109,In_1069);
nand U1242 (N_1242,In_877,In_1009);
nand U1243 (N_1243,In_756,In_636);
nand U1244 (N_1244,In_271,In_1146);
or U1245 (N_1245,In_66,In_1173);
or U1246 (N_1246,In_335,In_921);
xnor U1247 (N_1247,In_647,In_153);
nand U1248 (N_1248,In_716,In_1155);
or U1249 (N_1249,In_1477,In_978);
and U1250 (N_1250,In_887,In_1435);
and U1251 (N_1251,In_767,In_376);
nand U1252 (N_1252,In_336,In_842);
nand U1253 (N_1253,In_270,In_1229);
nand U1254 (N_1254,In_1106,In_339);
and U1255 (N_1255,In_1357,In_92);
and U1256 (N_1256,In_1407,In_613);
nor U1257 (N_1257,In_1102,In_1290);
and U1258 (N_1258,In_324,In_971);
and U1259 (N_1259,In_236,In_797);
or U1260 (N_1260,In_1310,In_1267);
and U1261 (N_1261,In_923,In_1306);
nor U1262 (N_1262,In_95,In_635);
and U1263 (N_1263,In_813,In_442);
or U1264 (N_1264,In_916,In_966);
and U1265 (N_1265,In_7,In_1425);
nand U1266 (N_1266,In_155,In_267);
nor U1267 (N_1267,In_609,In_149);
or U1268 (N_1268,In_327,In_1248);
nor U1269 (N_1269,In_1130,In_353);
or U1270 (N_1270,In_95,In_1331);
and U1271 (N_1271,In_1436,In_589);
and U1272 (N_1272,In_591,In_1387);
and U1273 (N_1273,In_864,In_422);
and U1274 (N_1274,In_1307,In_94);
nor U1275 (N_1275,In_358,In_1468);
or U1276 (N_1276,In_182,In_245);
nor U1277 (N_1277,In_1091,In_780);
nand U1278 (N_1278,In_835,In_1240);
nand U1279 (N_1279,In_607,In_108);
or U1280 (N_1280,In_676,In_1290);
and U1281 (N_1281,In_1264,In_671);
nand U1282 (N_1282,In_141,In_918);
nor U1283 (N_1283,In_127,In_1368);
nand U1284 (N_1284,In_360,In_303);
nor U1285 (N_1285,In_664,In_537);
and U1286 (N_1286,In_528,In_389);
and U1287 (N_1287,In_988,In_867);
nand U1288 (N_1288,In_733,In_349);
nor U1289 (N_1289,In_305,In_223);
nor U1290 (N_1290,In_384,In_90);
and U1291 (N_1291,In_1320,In_89);
nand U1292 (N_1292,In_1,In_1145);
nor U1293 (N_1293,In_999,In_47);
and U1294 (N_1294,In_598,In_241);
or U1295 (N_1295,In_181,In_1136);
nor U1296 (N_1296,In_566,In_99);
or U1297 (N_1297,In_1102,In_1017);
or U1298 (N_1298,In_2,In_418);
nor U1299 (N_1299,In_1321,In_452);
or U1300 (N_1300,In_340,In_302);
nand U1301 (N_1301,In_1279,In_493);
nand U1302 (N_1302,In_625,In_1182);
or U1303 (N_1303,In_560,In_930);
and U1304 (N_1304,In_567,In_1372);
and U1305 (N_1305,In_1083,In_1472);
nor U1306 (N_1306,In_156,In_143);
or U1307 (N_1307,In_990,In_542);
nor U1308 (N_1308,In_934,In_112);
and U1309 (N_1309,In_719,In_1087);
and U1310 (N_1310,In_425,In_1189);
nand U1311 (N_1311,In_408,In_183);
nand U1312 (N_1312,In_711,In_455);
or U1313 (N_1313,In_1269,In_887);
or U1314 (N_1314,In_1449,In_301);
or U1315 (N_1315,In_275,In_661);
xnor U1316 (N_1316,In_1354,In_692);
nor U1317 (N_1317,In_1427,In_279);
nand U1318 (N_1318,In_438,In_795);
nand U1319 (N_1319,In_1465,In_1021);
or U1320 (N_1320,In_709,In_198);
nor U1321 (N_1321,In_779,In_1490);
nor U1322 (N_1322,In_1259,In_927);
and U1323 (N_1323,In_999,In_44);
nor U1324 (N_1324,In_1408,In_1319);
and U1325 (N_1325,In_638,In_40);
or U1326 (N_1326,In_309,In_982);
nand U1327 (N_1327,In_866,In_69);
and U1328 (N_1328,In_356,In_1132);
or U1329 (N_1329,In_791,In_536);
or U1330 (N_1330,In_946,In_868);
xnor U1331 (N_1331,In_1412,In_1442);
or U1332 (N_1332,In_1361,In_1405);
nand U1333 (N_1333,In_818,In_708);
and U1334 (N_1334,In_702,In_749);
or U1335 (N_1335,In_1340,In_933);
nor U1336 (N_1336,In_1357,In_870);
nor U1337 (N_1337,In_311,In_1396);
and U1338 (N_1338,In_1100,In_601);
xor U1339 (N_1339,In_337,In_257);
nor U1340 (N_1340,In_224,In_76);
or U1341 (N_1341,In_340,In_1347);
and U1342 (N_1342,In_1170,In_1016);
nand U1343 (N_1343,In_950,In_1450);
nand U1344 (N_1344,In_506,In_519);
or U1345 (N_1345,In_1152,In_104);
nor U1346 (N_1346,In_824,In_1250);
or U1347 (N_1347,In_1028,In_968);
nand U1348 (N_1348,In_1327,In_649);
nand U1349 (N_1349,In_50,In_1430);
or U1350 (N_1350,In_39,In_880);
nand U1351 (N_1351,In_1341,In_45);
nand U1352 (N_1352,In_1004,In_1222);
nor U1353 (N_1353,In_43,In_356);
and U1354 (N_1354,In_414,In_385);
or U1355 (N_1355,In_28,In_1472);
nand U1356 (N_1356,In_722,In_951);
nand U1357 (N_1357,In_1051,In_20);
or U1358 (N_1358,In_1334,In_652);
or U1359 (N_1359,In_522,In_312);
or U1360 (N_1360,In_795,In_1202);
nand U1361 (N_1361,In_433,In_59);
xor U1362 (N_1362,In_301,In_352);
nor U1363 (N_1363,In_1328,In_1412);
or U1364 (N_1364,In_993,In_307);
and U1365 (N_1365,In_441,In_862);
and U1366 (N_1366,In_1283,In_880);
nand U1367 (N_1367,In_1065,In_1158);
nand U1368 (N_1368,In_950,In_1193);
nor U1369 (N_1369,In_43,In_462);
nand U1370 (N_1370,In_1010,In_1221);
and U1371 (N_1371,In_392,In_363);
nand U1372 (N_1372,In_620,In_1143);
nor U1373 (N_1373,In_1404,In_206);
nor U1374 (N_1374,In_556,In_1396);
or U1375 (N_1375,In_9,In_608);
and U1376 (N_1376,In_919,In_332);
and U1377 (N_1377,In_972,In_618);
nand U1378 (N_1378,In_926,In_396);
or U1379 (N_1379,In_783,In_1488);
or U1380 (N_1380,In_260,In_891);
or U1381 (N_1381,In_639,In_636);
nand U1382 (N_1382,In_569,In_975);
nand U1383 (N_1383,In_1114,In_158);
nand U1384 (N_1384,In_144,In_48);
nor U1385 (N_1385,In_161,In_793);
xnor U1386 (N_1386,In_54,In_509);
nand U1387 (N_1387,In_1427,In_1082);
xor U1388 (N_1388,In_110,In_1012);
nor U1389 (N_1389,In_186,In_1062);
nor U1390 (N_1390,In_1245,In_130);
and U1391 (N_1391,In_800,In_64);
and U1392 (N_1392,In_673,In_1485);
and U1393 (N_1393,In_596,In_1328);
nand U1394 (N_1394,In_521,In_1419);
nor U1395 (N_1395,In_545,In_413);
or U1396 (N_1396,In_898,In_159);
nand U1397 (N_1397,In_1129,In_1255);
or U1398 (N_1398,In_148,In_1152);
nor U1399 (N_1399,In_692,In_1348);
and U1400 (N_1400,In_621,In_1251);
nor U1401 (N_1401,In_341,In_1411);
nand U1402 (N_1402,In_740,In_1221);
and U1403 (N_1403,In_809,In_353);
xnor U1404 (N_1404,In_303,In_1009);
and U1405 (N_1405,In_1439,In_685);
xor U1406 (N_1406,In_188,In_644);
and U1407 (N_1407,In_1165,In_67);
nand U1408 (N_1408,In_243,In_1012);
and U1409 (N_1409,In_548,In_71);
nor U1410 (N_1410,In_583,In_638);
nand U1411 (N_1411,In_256,In_1027);
and U1412 (N_1412,In_1154,In_306);
nor U1413 (N_1413,In_183,In_483);
or U1414 (N_1414,In_844,In_1385);
and U1415 (N_1415,In_73,In_989);
or U1416 (N_1416,In_1112,In_404);
or U1417 (N_1417,In_1310,In_1054);
nor U1418 (N_1418,In_728,In_548);
and U1419 (N_1419,In_1031,In_1307);
or U1420 (N_1420,In_80,In_1303);
nor U1421 (N_1421,In_48,In_730);
or U1422 (N_1422,In_572,In_1455);
or U1423 (N_1423,In_1467,In_677);
or U1424 (N_1424,In_443,In_1218);
or U1425 (N_1425,In_1146,In_566);
nand U1426 (N_1426,In_179,In_534);
nand U1427 (N_1427,In_673,In_1191);
nor U1428 (N_1428,In_903,In_522);
nand U1429 (N_1429,In_483,In_961);
or U1430 (N_1430,In_820,In_425);
xnor U1431 (N_1431,In_809,In_1276);
or U1432 (N_1432,In_533,In_304);
or U1433 (N_1433,In_6,In_12);
nand U1434 (N_1434,In_971,In_459);
or U1435 (N_1435,In_1175,In_230);
or U1436 (N_1436,In_151,In_1473);
nand U1437 (N_1437,In_812,In_143);
or U1438 (N_1438,In_1140,In_1294);
and U1439 (N_1439,In_1269,In_446);
nor U1440 (N_1440,In_454,In_1434);
or U1441 (N_1441,In_1116,In_317);
or U1442 (N_1442,In_1156,In_466);
or U1443 (N_1443,In_612,In_1216);
and U1444 (N_1444,In_567,In_1196);
or U1445 (N_1445,In_1372,In_1339);
nand U1446 (N_1446,In_572,In_190);
nand U1447 (N_1447,In_537,In_361);
nor U1448 (N_1448,In_1080,In_1041);
and U1449 (N_1449,In_1003,In_754);
and U1450 (N_1450,In_172,In_978);
nor U1451 (N_1451,In_1429,In_864);
nand U1452 (N_1452,In_1190,In_592);
xnor U1453 (N_1453,In_126,In_996);
and U1454 (N_1454,In_239,In_318);
and U1455 (N_1455,In_1244,In_654);
nor U1456 (N_1456,In_1310,In_242);
nor U1457 (N_1457,In_730,In_465);
and U1458 (N_1458,In_471,In_999);
and U1459 (N_1459,In_1256,In_804);
xor U1460 (N_1460,In_313,In_836);
nand U1461 (N_1461,In_746,In_874);
or U1462 (N_1462,In_123,In_1437);
nand U1463 (N_1463,In_91,In_216);
nand U1464 (N_1464,In_1105,In_13);
or U1465 (N_1465,In_449,In_1346);
nor U1466 (N_1466,In_187,In_503);
nor U1467 (N_1467,In_1408,In_1450);
nor U1468 (N_1468,In_1088,In_1458);
and U1469 (N_1469,In_158,In_463);
and U1470 (N_1470,In_997,In_197);
or U1471 (N_1471,In_749,In_255);
and U1472 (N_1472,In_568,In_1024);
and U1473 (N_1473,In_912,In_198);
or U1474 (N_1474,In_1315,In_1214);
nand U1475 (N_1475,In_307,In_625);
nor U1476 (N_1476,In_388,In_1440);
xor U1477 (N_1477,In_512,In_1479);
nor U1478 (N_1478,In_529,In_823);
and U1479 (N_1479,In_903,In_1065);
nor U1480 (N_1480,In_836,In_473);
and U1481 (N_1481,In_117,In_944);
nand U1482 (N_1482,In_118,In_94);
xor U1483 (N_1483,In_902,In_696);
nand U1484 (N_1484,In_92,In_946);
nand U1485 (N_1485,In_762,In_554);
nor U1486 (N_1486,In_1090,In_319);
or U1487 (N_1487,In_247,In_1277);
and U1488 (N_1488,In_1225,In_366);
and U1489 (N_1489,In_556,In_111);
or U1490 (N_1490,In_645,In_603);
xnor U1491 (N_1491,In_202,In_649);
nand U1492 (N_1492,In_1101,In_473);
and U1493 (N_1493,In_1146,In_226);
xnor U1494 (N_1494,In_1141,In_794);
and U1495 (N_1495,In_837,In_1267);
and U1496 (N_1496,In_816,In_1114);
or U1497 (N_1497,In_129,In_1307);
nor U1498 (N_1498,In_46,In_1393);
nor U1499 (N_1499,In_386,In_1211);
or U1500 (N_1500,N_478,N_147);
or U1501 (N_1501,N_208,N_506);
nor U1502 (N_1502,N_1323,N_581);
nor U1503 (N_1503,N_122,N_1024);
nand U1504 (N_1504,N_883,N_594);
or U1505 (N_1505,N_635,N_287);
nand U1506 (N_1506,N_177,N_1163);
xor U1507 (N_1507,N_0,N_788);
nor U1508 (N_1508,N_910,N_318);
nand U1509 (N_1509,N_653,N_659);
nor U1510 (N_1510,N_731,N_1231);
or U1511 (N_1511,N_1472,N_1460);
nand U1512 (N_1512,N_523,N_1100);
and U1513 (N_1513,N_1482,N_400);
and U1514 (N_1514,N_903,N_288);
or U1515 (N_1515,N_357,N_45);
or U1516 (N_1516,N_829,N_102);
xor U1517 (N_1517,N_819,N_1415);
or U1518 (N_1518,N_466,N_921);
and U1519 (N_1519,N_912,N_1421);
nand U1520 (N_1520,N_1063,N_764);
nor U1521 (N_1521,N_1322,N_338);
xnor U1522 (N_1522,N_94,N_1099);
nand U1523 (N_1523,N_1467,N_399);
nor U1524 (N_1524,N_951,N_176);
nor U1525 (N_1525,N_741,N_629);
and U1526 (N_1526,N_541,N_1009);
nand U1527 (N_1527,N_92,N_175);
nor U1528 (N_1528,N_354,N_620);
and U1529 (N_1529,N_114,N_336);
nor U1530 (N_1530,N_1027,N_1022);
or U1531 (N_1531,N_803,N_527);
nor U1532 (N_1532,N_518,N_929);
xor U1533 (N_1533,N_926,N_39);
nand U1534 (N_1534,N_121,N_98);
and U1535 (N_1535,N_369,N_1309);
or U1536 (N_1536,N_791,N_631);
or U1537 (N_1537,N_1021,N_187);
xnor U1538 (N_1538,N_210,N_285);
nand U1539 (N_1539,N_566,N_660);
nor U1540 (N_1540,N_289,N_55);
nand U1541 (N_1541,N_1432,N_645);
xnor U1542 (N_1542,N_93,N_1423);
nor U1543 (N_1543,N_1229,N_312);
and U1544 (N_1544,N_107,N_186);
nand U1545 (N_1545,N_1481,N_615);
and U1546 (N_1546,N_862,N_1439);
and U1547 (N_1547,N_251,N_936);
nor U1548 (N_1548,N_1417,N_668);
xor U1549 (N_1549,N_589,N_56);
nand U1550 (N_1550,N_901,N_1388);
nand U1551 (N_1551,N_815,N_691);
xnor U1552 (N_1552,N_712,N_36);
nor U1553 (N_1553,N_1375,N_663);
nand U1554 (N_1554,N_1320,N_1148);
or U1555 (N_1555,N_667,N_1137);
or U1556 (N_1556,N_1040,N_173);
xnor U1557 (N_1557,N_999,N_1488);
and U1558 (N_1558,N_447,N_676);
nor U1559 (N_1559,N_738,N_1332);
or U1560 (N_1560,N_586,N_1463);
nand U1561 (N_1561,N_627,N_345);
nand U1562 (N_1562,N_410,N_1136);
or U1563 (N_1563,N_1113,N_967);
or U1564 (N_1564,N_670,N_626);
nor U1565 (N_1565,N_1110,N_584);
and U1566 (N_1566,N_623,N_442);
nor U1567 (N_1567,N_1193,N_907);
nand U1568 (N_1568,N_1219,N_1311);
nor U1569 (N_1569,N_255,N_11);
or U1570 (N_1570,N_1365,N_892);
xnor U1571 (N_1571,N_1476,N_625);
nand U1572 (N_1572,N_979,N_1343);
nand U1573 (N_1573,N_1103,N_524);
nor U1574 (N_1574,N_278,N_1290);
and U1575 (N_1575,N_512,N_46);
and U1576 (N_1576,N_1215,N_1354);
and U1577 (N_1577,N_622,N_927);
nor U1578 (N_1578,N_178,N_314);
or U1579 (N_1579,N_476,N_1294);
and U1580 (N_1580,N_1392,N_840);
nand U1581 (N_1581,N_1457,N_82);
or U1582 (N_1582,N_1165,N_120);
xor U1583 (N_1583,N_600,N_1093);
and U1584 (N_1584,N_785,N_727);
and U1585 (N_1585,N_641,N_80);
and U1586 (N_1586,N_772,N_511);
xnor U1587 (N_1587,N_456,N_1259);
or U1588 (N_1588,N_1102,N_1014);
and U1589 (N_1589,N_215,N_1387);
nand U1590 (N_1590,N_1428,N_1123);
and U1591 (N_1591,N_202,N_1043);
nand U1592 (N_1592,N_726,N_1418);
and U1593 (N_1593,N_679,N_482);
or U1594 (N_1594,N_780,N_133);
nand U1595 (N_1595,N_1321,N_847);
or U1596 (N_1596,N_1207,N_262);
xnor U1597 (N_1597,N_925,N_274);
or U1598 (N_1598,N_953,N_284);
nor U1599 (N_1599,N_734,N_575);
nand U1600 (N_1600,N_869,N_1328);
or U1601 (N_1601,N_704,N_1389);
or U1602 (N_1602,N_1041,N_245);
nand U1603 (N_1603,N_219,N_1000);
or U1604 (N_1604,N_978,N_790);
and U1605 (N_1605,N_1443,N_1085);
and U1606 (N_1606,N_153,N_908);
nand U1607 (N_1607,N_918,N_1178);
nor U1608 (N_1608,N_307,N_1292);
nand U1609 (N_1609,N_1273,N_1245);
nor U1610 (N_1610,N_761,N_398);
xnor U1611 (N_1611,N_1285,N_1307);
and U1612 (N_1612,N_1445,N_1382);
nand U1613 (N_1613,N_64,N_954);
or U1614 (N_1614,N_583,N_181);
nor U1615 (N_1615,N_789,N_313);
xor U1616 (N_1616,N_864,N_1240);
nand U1617 (N_1617,N_1166,N_436);
or U1618 (N_1618,N_477,N_905);
nand U1619 (N_1619,N_207,N_188);
nor U1620 (N_1620,N_481,N_909);
nor U1621 (N_1621,N_1187,N_1055);
nor U1622 (N_1622,N_516,N_880);
or U1623 (N_1623,N_674,N_1045);
and U1624 (N_1624,N_1282,N_928);
nor U1625 (N_1625,N_27,N_1096);
nand U1626 (N_1626,N_1026,N_339);
or U1627 (N_1627,N_248,N_261);
or U1628 (N_1628,N_100,N_533);
and U1629 (N_1629,N_579,N_706);
nor U1630 (N_1630,N_787,N_1056);
nand U1631 (N_1631,N_1456,N_1304);
and U1632 (N_1632,N_460,N_856);
nor U1633 (N_1633,N_458,N_654);
or U1634 (N_1634,N_1475,N_1441);
nor U1635 (N_1635,N_375,N_521);
nand U1636 (N_1636,N_1190,N_662);
nand U1637 (N_1637,N_1331,N_1160);
and U1638 (N_1638,N_142,N_795);
and U1639 (N_1639,N_146,N_993);
xnor U1640 (N_1640,N_14,N_1153);
nand U1641 (N_1641,N_637,N_868);
and U1642 (N_1642,N_1217,N_271);
and U1643 (N_1643,N_746,N_413);
nor U1644 (N_1644,N_1084,N_537);
or U1645 (N_1645,N_280,N_1083);
nor U1646 (N_1646,N_1372,N_522);
and U1647 (N_1647,N_1402,N_947);
xor U1648 (N_1648,N_747,N_152);
xor U1649 (N_1649,N_801,N_802);
nor U1650 (N_1650,N_1279,N_1330);
or U1651 (N_1651,N_1408,N_557);
or U1652 (N_1652,N_902,N_63);
nand U1653 (N_1653,N_303,N_520);
nand U1654 (N_1654,N_291,N_1248);
nand U1655 (N_1655,N_54,N_783);
nand U1656 (N_1656,N_1012,N_180);
nand U1657 (N_1657,N_295,N_1204);
and U1658 (N_1658,N_965,N_1139);
or U1659 (N_1659,N_337,N_690);
nand U1660 (N_1660,N_1434,N_420);
and U1661 (N_1661,N_112,N_552);
nand U1662 (N_1662,N_1288,N_655);
nand U1663 (N_1663,N_531,N_652);
or U1664 (N_1664,N_479,N_150);
nor U1665 (N_1665,N_322,N_20);
and U1666 (N_1666,N_818,N_920);
xor U1667 (N_1667,N_1003,N_608);
nor U1668 (N_1668,N_24,N_1345);
nand U1669 (N_1669,N_1237,N_1244);
nor U1670 (N_1670,N_342,N_71);
nor U1671 (N_1671,N_415,N_561);
or U1672 (N_1672,N_1274,N_311);
and U1673 (N_1673,N_1334,N_1031);
or U1674 (N_1674,N_425,N_1379);
and U1675 (N_1675,N_651,N_1023);
xnor U1676 (N_1676,N_214,N_316);
and U1677 (N_1677,N_97,N_195);
or U1678 (N_1678,N_1002,N_159);
nand U1679 (N_1679,N_964,N_675);
nand U1680 (N_1680,N_841,N_1074);
nand U1681 (N_1681,N_444,N_1315);
xor U1682 (N_1682,N_1477,N_639);
and U1683 (N_1683,N_700,N_863);
nor U1684 (N_1684,N_301,N_365);
nor U1685 (N_1685,N_534,N_1414);
and U1686 (N_1686,N_833,N_143);
nand U1687 (N_1687,N_1422,N_244);
and U1688 (N_1688,N_1186,N_373);
nor U1689 (N_1689,N_148,N_1368);
nand U1690 (N_1690,N_1358,N_96);
or U1691 (N_1691,N_1342,N_474);
nand U1692 (N_1692,N_31,N_1132);
nor U1693 (N_1693,N_1130,N_406);
nor U1694 (N_1694,N_1234,N_1424);
and U1695 (N_1695,N_1069,N_385);
or U1696 (N_1696,N_1438,N_1452);
or U1697 (N_1697,N_347,N_179);
and U1698 (N_1698,N_720,N_644);
nor U1699 (N_1699,N_1453,N_315);
nor U1700 (N_1700,N_1386,N_235);
nor U1701 (N_1701,N_1196,N_12);
and U1702 (N_1702,N_366,N_368);
nor U1703 (N_1703,N_688,N_718);
nand U1704 (N_1704,N_1407,N_695);
and U1705 (N_1705,N_1177,N_328);
nand U1706 (N_1706,N_241,N_270);
nor U1707 (N_1707,N_762,N_1067);
nor U1708 (N_1708,N_633,N_199);
nand U1709 (N_1709,N_427,N_596);
nand U1710 (N_1710,N_1241,N_1369);
and U1711 (N_1711,N_254,N_1306);
nor U1712 (N_1712,N_1192,N_1433);
nand U1713 (N_1713,N_590,N_725);
or U1714 (N_1714,N_602,N_752);
or U1715 (N_1715,N_814,N_10);
and U1716 (N_1716,N_944,N_6);
nor U1717 (N_1717,N_543,N_1280);
nor U1718 (N_1718,N_1376,N_41);
and U1719 (N_1719,N_129,N_1222);
nand U1720 (N_1720,N_1066,N_1498);
nand U1721 (N_1721,N_414,N_4);
xnor U1722 (N_1722,N_983,N_1390);
nor U1723 (N_1723,N_835,N_1474);
nand U1724 (N_1724,N_528,N_1138);
nor U1725 (N_1725,N_732,N_703);
nor U1726 (N_1726,N_906,N_52);
nor U1727 (N_1727,N_713,N_457);
and U1728 (N_1728,N_904,N_1201);
nand U1729 (N_1729,N_1122,N_857);
nor U1730 (N_1730,N_751,N_111);
or U1731 (N_1731,N_238,N_1161);
or U1732 (N_1732,N_606,N_517);
or U1733 (N_1733,N_922,N_430);
or U1734 (N_1734,N_578,N_616);
and U1735 (N_1735,N_698,N_1269);
nor U1736 (N_1736,N_530,N_394);
nand U1737 (N_1737,N_246,N_431);
and U1738 (N_1738,N_418,N_302);
and U1739 (N_1739,N_432,N_1361);
or U1740 (N_1740,N_35,N_1194);
nand U1741 (N_1741,N_709,N_1220);
and U1742 (N_1742,N_630,N_405);
nand U1743 (N_1743,N_201,N_666);
nor U1744 (N_1744,N_189,N_996);
and U1745 (N_1745,N_108,N_1019);
nor U1746 (N_1746,N_230,N_292);
and U1747 (N_1747,N_1145,N_1454);
or U1748 (N_1748,N_433,N_475);
and U1749 (N_1749,N_1303,N_642);
and U1750 (N_1750,N_573,N_79);
nor U1751 (N_1751,N_831,N_1105);
nand U1752 (N_1752,N_1291,N_1370);
nor U1753 (N_1753,N_937,N_931);
nand U1754 (N_1754,N_1243,N_90);
nand U1755 (N_1755,N_1250,N_809);
nand U1756 (N_1756,N_1068,N_853);
nor U1757 (N_1757,N_1141,N_852);
nor U1758 (N_1758,N_872,N_44);
or U1759 (N_1759,N_551,N_154);
or U1760 (N_1760,N_1164,N_434);
and U1761 (N_1761,N_1227,N_823);
or U1762 (N_1762,N_1039,N_1104);
or U1763 (N_1763,N_721,N_1494);
and U1764 (N_1764,N_169,N_1347);
and U1765 (N_1765,N_1242,N_396);
nand U1766 (N_1766,N_735,N_770);
nand U1767 (N_1767,N_705,N_848);
xor U1768 (N_1768,N_825,N_372);
nand U1769 (N_1769,N_1173,N_23);
and U1770 (N_1770,N_69,N_268);
nor U1771 (N_1771,N_267,N_913);
or U1772 (N_1772,N_451,N_610);
nor U1773 (N_1773,N_885,N_66);
xor U1774 (N_1774,N_658,N_1111);
xor U1775 (N_1775,N_198,N_813);
nor U1776 (N_1776,N_513,N_439);
and U1777 (N_1777,N_149,N_497);
nand U1778 (N_1778,N_332,N_234);
or U1779 (N_1779,N_500,N_1072);
xnor U1780 (N_1780,N_1064,N_499);
or U1781 (N_1781,N_1403,N_404);
nand U1782 (N_1782,N_206,N_250);
nand U1783 (N_1783,N_697,N_165);
and U1784 (N_1784,N_992,N_13);
nor U1785 (N_1785,N_1366,N_1451);
or U1786 (N_1786,N_988,N_265);
and U1787 (N_1787,N_807,N_222);
and U1788 (N_1788,N_775,N_955);
xnor U1789 (N_1789,N_1124,N_1058);
nor U1790 (N_1790,N_845,N_156);
or U1791 (N_1791,N_1413,N_382);
nor U1792 (N_1792,N_827,N_836);
nand U1793 (N_1793,N_744,N_1289);
and U1794 (N_1794,N_1281,N_330);
nor U1795 (N_1795,N_225,N_317);
xor U1796 (N_1796,N_1268,N_1091);
nor U1797 (N_1797,N_72,N_304);
nand U1798 (N_1798,N_151,N_1140);
nor U1799 (N_1799,N_17,N_125);
nor U1800 (N_1800,N_1335,N_919);
or U1801 (N_1801,N_21,N_1429);
nor U1802 (N_1802,N_15,N_784);
nand U1803 (N_1803,N_1004,N_2);
xnor U1804 (N_1804,N_419,N_480);
or U1805 (N_1805,N_587,N_381);
xor U1806 (N_1806,N_1473,N_886);
xnor U1807 (N_1807,N_582,N_259);
or U1808 (N_1808,N_275,N_42);
nand U1809 (N_1809,N_76,N_1075);
nor U1810 (N_1810,N_281,N_383);
nand U1811 (N_1811,N_598,N_677);
nor U1812 (N_1812,N_29,N_341);
or U1813 (N_1813,N_397,N_1257);
xor U1814 (N_1814,N_650,N_503);
xor U1815 (N_1815,N_1065,N_877);
nand U1816 (N_1816,N_443,N_145);
and U1817 (N_1817,N_604,N_1125);
nand U1818 (N_1818,N_1131,N_1404);
or U1819 (N_1819,N_804,N_585);
xor U1820 (N_1820,N_438,N_1209);
and U1821 (N_1821,N_621,N_1094);
nor U1822 (N_1822,N_916,N_38);
nor U1823 (N_1823,N_981,N_221);
nor U1824 (N_1824,N_646,N_605);
nor U1825 (N_1825,N_47,N_170);
and U1826 (N_1826,N_1496,N_1081);
nor U1827 (N_1827,N_1020,N_1295);
and U1828 (N_1828,N_564,N_1049);
or U1829 (N_1829,N_1169,N_859);
nor U1830 (N_1830,N_970,N_1133);
nor U1831 (N_1831,N_297,N_7);
nand U1832 (N_1832,N_1296,N_1262);
or U1833 (N_1833,N_990,N_1470);
and U1834 (N_1834,N_811,N_32);
or U1835 (N_1835,N_948,N_555);
or U1836 (N_1836,N_334,N_138);
nand U1837 (N_1837,N_733,N_661);
nand U1838 (N_1838,N_493,N_286);
nand U1839 (N_1839,N_535,N_386);
nand U1840 (N_1840,N_1459,N_3);
nor U1841 (N_1841,N_1168,N_716);
xnor U1842 (N_1842,N_1329,N_1486);
or U1843 (N_1843,N_1060,N_200);
or U1844 (N_1844,N_1420,N_888);
or U1845 (N_1845,N_258,N_851);
nand U1846 (N_1846,N_973,N_782);
nor U1847 (N_1847,N_1126,N_532);
nand U1848 (N_1848,N_84,N_305);
nor U1849 (N_1849,N_437,N_1483);
and U1850 (N_1850,N_619,N_540);
nor U1851 (N_1851,N_1442,N_184);
nand U1852 (N_1852,N_486,N_865);
nor U1853 (N_1853,N_75,N_968);
nor U1854 (N_1854,N_1151,N_837);
and U1855 (N_1855,N_753,N_471);
and U1856 (N_1856,N_1208,N_371);
nor U1857 (N_1857,N_340,N_306);
or U1858 (N_1858,N_157,N_308);
and U1859 (N_1859,N_158,N_352);
nand U1860 (N_1860,N_239,N_448);
nor U1861 (N_1861,N_957,N_812);
and U1862 (N_1862,N_127,N_18);
nor U1863 (N_1863,N_1490,N_393);
and U1864 (N_1864,N_797,N_465);
nor U1865 (N_1865,N_1272,N_130);
nor U1866 (N_1866,N_509,N_424);
or U1867 (N_1867,N_1184,N_1362);
nand U1868 (N_1868,N_1359,N_1088);
xnor U1869 (N_1869,N_538,N_544);
or U1870 (N_1870,N_998,N_966);
nor U1871 (N_1871,N_1319,N_749);
and U1872 (N_1872,N_467,N_550);
or U1873 (N_1873,N_455,N_893);
nor U1874 (N_1874,N_839,N_980);
or U1875 (N_1875,N_1010,N_1032);
nor U1876 (N_1876,N_1212,N_1230);
nand U1877 (N_1877,N_1437,N_299);
or U1878 (N_1878,N_924,N_1175);
nor U1879 (N_1879,N_942,N_362);
nor U1880 (N_1880,N_329,N_53);
or U1881 (N_1881,N_501,N_1317);
nand U1882 (N_1882,N_1211,N_1198);
or U1883 (N_1883,N_1051,N_755);
nor U1884 (N_1884,N_1344,N_1393);
or U1885 (N_1885,N_640,N_231);
nor U1886 (N_1886,N_9,N_490);
nor U1887 (N_1887,N_298,N_1391);
nor U1888 (N_1888,N_1412,N_873);
nor U1889 (N_1889,N_923,N_331);
and U1890 (N_1890,N_717,N_1265);
nor U1891 (N_1891,N_462,N_1191);
nand U1892 (N_1892,N_678,N_441);
nor U1893 (N_1893,N_539,N_1478);
or U1894 (N_1894,N_1152,N_236);
and U1895 (N_1895,N_1238,N_612);
or U1896 (N_1896,N_634,N_894);
nand U1897 (N_1897,N_220,N_570);
nor U1898 (N_1898,N_350,N_226);
or U1899 (N_1899,N_1016,N_333);
nand U1900 (N_1900,N_229,N_242);
or U1901 (N_1901,N_624,N_693);
nand U1902 (N_1902,N_1214,N_1033);
nand U1903 (N_1903,N_89,N_25);
xor U1904 (N_1904,N_1117,N_118);
nor U1905 (N_1905,N_325,N_1346);
or U1906 (N_1906,N_1233,N_875);
xor U1907 (N_1907,N_1061,N_171);
nand U1908 (N_1908,N_1293,N_203);
xor U1909 (N_1909,N_935,N_806);
nand U1910 (N_1910,N_1223,N_822);
nand U1911 (N_1911,N_793,N_283);
nor U1912 (N_1912,N_1286,N_1070);
xor U1913 (N_1913,N_387,N_1384);
nor U1914 (N_1914,N_850,N_1373);
and U1915 (N_1915,N_769,N_5);
xor U1916 (N_1916,N_781,N_1254);
nand U1917 (N_1917,N_756,N_380);
or U1918 (N_1918,N_743,N_854);
nor U1919 (N_1919,N_1005,N_702);
or U1920 (N_1920,N_440,N_140);
or U1921 (N_1921,N_519,N_1299);
nor U1922 (N_1922,N_1006,N_1277);
nor U1923 (N_1923,N_1011,N_416);
or U1924 (N_1924,N_607,N_1394);
or U1925 (N_1925,N_1260,N_472);
and U1926 (N_1926,N_799,N_273);
and U1927 (N_1927,N_952,N_1087);
or U1928 (N_1928,N_294,N_423);
nand U1929 (N_1929,N_326,N_30);
nand U1930 (N_1930,N_574,N_636);
and U1931 (N_1931,N_67,N_1410);
nor U1932 (N_1932,N_861,N_1448);
nand U1933 (N_1933,N_1050,N_356);
nand U1934 (N_1934,N_737,N_946);
nand U1935 (N_1935,N_971,N_778);
nand U1936 (N_1936,N_1419,N_959);
xnor U1937 (N_1937,N_1251,N_997);
or U1938 (N_1938,N_277,N_989);
xnor U1939 (N_1939,N_1302,N_536);
nor U1940 (N_1940,N_483,N_542);
or U1941 (N_1941,N_632,N_421);
and U1942 (N_1942,N_963,N_665);
nand U1943 (N_1943,N_1340,N_1305);
xnor U1944 (N_1944,N_135,N_568);
nor U1945 (N_1945,N_264,N_742);
nor U1946 (N_1946,N_445,N_351);
and U1947 (N_1947,N_249,N_1409);
nand U1948 (N_1948,N_1179,N_263);
or U1949 (N_1949,N_685,N_1156);
or U1950 (N_1950,N_1200,N_849);
nand U1951 (N_1951,N_866,N_131);
nand U1952 (N_1952,N_450,N_593);
or U1953 (N_1953,N_617,N_323);
and U1954 (N_1954,N_740,N_1339);
or U1955 (N_1955,N_934,N_205);
nand U1956 (N_1956,N_601,N_353);
nand U1957 (N_1957,N_681,N_1035);
nand U1958 (N_1958,N_81,N_1092);
nor U1959 (N_1959,N_719,N_1158);
or U1960 (N_1960,N_16,N_1310);
xor U1961 (N_1961,N_300,N_977);
and U1962 (N_1962,N_969,N_1015);
or U1963 (N_1963,N_1495,N_57);
nor U1964 (N_1964,N_559,N_673);
nor U1965 (N_1965,N_166,N_1449);
and U1966 (N_1966,N_588,N_609);
and U1967 (N_1967,N_408,N_232);
and U1968 (N_1968,N_1425,N_1395);
or U1969 (N_1969,N_1155,N_190);
nand U1970 (N_1970,N_496,N_1492);
nor U1971 (N_1971,N_355,N_1098);
and U1972 (N_1972,N_1308,N_1400);
and U1973 (N_1973,N_560,N_464);
xnor U1974 (N_1974,N_321,N_119);
and U1975 (N_1975,N_85,N_580);
nand U1976 (N_1976,N_669,N_429);
xor U1977 (N_1977,N_1357,N_945);
and U1978 (N_1978,N_817,N_1116);
and U1979 (N_1979,N_510,N_105);
nand U1980 (N_1980,N_370,N_878);
nand U1981 (N_1981,N_1287,N_1313);
xor U1982 (N_1982,N_914,N_1034);
nor U1983 (N_1983,N_1399,N_943);
nor U1984 (N_1984,N_1082,N_377);
and U1985 (N_1985,N_599,N_253);
and U1986 (N_1986,N_1071,N_707);
nand U1987 (N_1987,N_1018,N_1183);
nor U1988 (N_1988,N_1465,N_358);
nand U1989 (N_1989,N_473,N_1297);
or U1990 (N_1990,N_830,N_1174);
and U1991 (N_1991,N_95,N_569);
nand U1992 (N_1992,N_1150,N_116);
nand U1993 (N_1993,N_1176,N_1489);
nand U1994 (N_1994,N_1225,N_1333);
and U1995 (N_1995,N_487,N_1485);
or U1996 (N_1996,N_765,N_364);
nor U1997 (N_1997,N_1188,N_1007);
xnor U1998 (N_1998,N_899,N_656);
and U1999 (N_1999,N_1106,N_1154);
nor U2000 (N_2000,N_768,N_269);
and U2001 (N_2001,N_881,N_858);
nor U2002 (N_2002,N_991,N_240);
nand U2003 (N_2003,N_113,N_1363);
nand U2004 (N_2004,N_834,N_74);
or U2005 (N_2005,N_1,N_389);
nor U2006 (N_2006,N_1162,N_1261);
or U2007 (N_2007,N_745,N_260);
nand U2008 (N_2008,N_213,N_545);
or U2009 (N_2009,N_879,N_1197);
xnor U2010 (N_2010,N_1159,N_452);
nor U2011 (N_2011,N_124,N_192);
and U2012 (N_2012,N_614,N_648);
nand U2013 (N_2013,N_193,N_359);
nand U2014 (N_2014,N_961,N_1129);
or U2015 (N_2015,N_1221,N_191);
xnor U2016 (N_2016,N_1406,N_26);
nand U2017 (N_2017,N_870,N_736);
and U2018 (N_2018,N_1440,N_547);
and U2019 (N_2019,N_276,N_218);
and U2020 (N_2020,N_1300,N_495);
and U2021 (N_2021,N_1271,N_1107);
and U2022 (N_2022,N_412,N_1351);
nand U2023 (N_2023,N_1458,N_563);
nand U2024 (N_2024,N_463,N_172);
nor U2025 (N_2025,N_91,N_77);
and U2026 (N_2026,N_1054,N_554);
xnor U2027 (N_2027,N_832,N_1089);
and U2028 (N_2028,N_1461,N_1398);
or U2029 (N_2029,N_710,N_417);
and U2030 (N_2030,N_671,N_760);
or U2031 (N_2031,N_882,N_1314);
or U2032 (N_2032,N_469,N_618);
nor U2033 (N_2033,N_1213,N_526);
or U2034 (N_2034,N_571,N_1120);
nor U2035 (N_2035,N_1336,N_1232);
or U2036 (N_2036,N_1147,N_344);
nor U2037 (N_2037,N_507,N_1446);
nand U2038 (N_2038,N_390,N_1205);
and U2039 (N_2039,N_1042,N_110);
and U2040 (N_2040,N_115,N_272);
nand U2041 (N_2041,N_887,N_958);
nor U2042 (N_2042,N_86,N_320);
nor U2043 (N_2043,N_686,N_1275);
nand U2044 (N_2044,N_1108,N_88);
xnor U2045 (N_2045,N_1350,N_139);
or U2046 (N_2046,N_1078,N_1252);
or U2047 (N_2047,N_391,N_1324);
nor U2048 (N_2048,N_376,N_613);
nand U2049 (N_2049,N_504,N_73);
nand U2050 (N_2050,N_895,N_794);
and U2051 (N_2051,N_319,N_577);
or U2052 (N_2052,N_682,N_78);
and U2053 (N_2053,N_722,N_1109);
or U2054 (N_2054,N_546,N_1127);
and U2055 (N_2055,N_962,N_132);
nand U2056 (N_2056,N_938,N_1086);
and U2057 (N_2057,N_1468,N_1037);
nor U2058 (N_2058,N_558,N_1218);
nand U2059 (N_2059,N_1008,N_638);
xnor U2060 (N_2060,N_374,N_174);
nor U2061 (N_2061,N_576,N_361);
xnor U2062 (N_2062,N_798,N_360);
nor U2063 (N_2063,N_247,N_1278);
and U2064 (N_2064,N_657,N_1101);
nand U2065 (N_2065,N_1325,N_821);
xnor U2066 (N_2066,N_1480,N_1142);
xnor U2067 (N_2067,N_1224,N_349);
nand U2068 (N_2068,N_379,N_1264);
nand U2069 (N_2069,N_1316,N_805);
nand U2070 (N_2070,N_956,N_134);
and U2071 (N_2071,N_844,N_327);
nor U2072 (N_2072,N_446,N_1499);
nand U2073 (N_2073,N_1469,N_1228);
and U2074 (N_2074,N_1170,N_941);
or U2075 (N_2075,N_233,N_796);
nand U2076 (N_2076,N_792,N_1327);
or U2077 (N_2077,N_426,N_960);
or U2078 (N_2078,N_1364,N_137);
and U2079 (N_2079,N_1435,N_194);
xnor U2080 (N_2080,N_1046,N_1466);
or U2081 (N_2081,N_1118,N_217);
nand U2082 (N_2082,N_826,N_128);
or U2083 (N_2083,N_1180,N_611);
and U2084 (N_2084,N_771,N_324);
and U2085 (N_2085,N_1097,N_724);
and U2086 (N_2086,N_891,N_1263);
nor U2087 (N_2087,N_939,N_409);
xor U2088 (N_2088,N_468,N_689);
nor U2089 (N_2089,N_1210,N_1276);
nand U2090 (N_2090,N_1203,N_407);
or U2091 (N_2091,N_33,N_243);
nor U2092 (N_2092,N_411,N_1057);
nand U2093 (N_2093,N_51,N_309);
xor U2094 (N_2094,N_1115,N_348);
xor U2095 (N_2095,N_99,N_1484);
nand U2096 (N_2096,N_592,N_22);
and U2097 (N_2097,N_1167,N_296);
nor U2098 (N_2098,N_196,N_182);
and U2099 (N_2099,N_223,N_562);
or U2100 (N_2100,N_141,N_68);
and U2101 (N_2101,N_28,N_683);
nor U2102 (N_2102,N_1149,N_1013);
and U2103 (N_2103,N_1146,N_846);
nand U2104 (N_2104,N_461,N_1121);
nor U2105 (N_2105,N_867,N_1444);
nand U2106 (N_2106,N_1326,N_933);
and U2107 (N_2107,N_1235,N_982);
nand U2108 (N_2108,N_986,N_708);
nand U2109 (N_2109,N_730,N_729);
nand U2110 (N_2110,N_714,N_1427);
nand U2111 (N_2111,N_59,N_728);
nor U2112 (N_2112,N_1236,N_485);
xnor U2113 (N_2113,N_1171,N_1255);
or U2114 (N_2114,N_1182,N_774);
or U2115 (N_2115,N_1464,N_949);
nand U2116 (N_2116,N_553,N_164);
xor U2117 (N_2117,N_828,N_876);
or U2118 (N_2118,N_106,N_197);
or U2119 (N_2119,N_1185,N_591);
and U2120 (N_2120,N_61,N_459);
or U2121 (N_2121,N_800,N_395);
and U2122 (N_2122,N_266,N_548);
nor U2123 (N_2123,N_1076,N_889);
and U2124 (N_2124,N_1436,N_628);
or U2125 (N_2125,N_1134,N_454);
or U2126 (N_2126,N_505,N_204);
or U2127 (N_2127,N_1079,N_1266);
or U2128 (N_2128,N_1044,N_723);
xnor U2129 (N_2129,N_256,N_1038);
or U2130 (N_2130,N_363,N_748);
nor U2131 (N_2131,N_525,N_101);
and U2132 (N_2132,N_972,N_779);
and U2133 (N_2133,N_838,N_1356);
or U2134 (N_2134,N_1431,N_1284);
nand U2135 (N_2135,N_975,N_1360);
nand U2136 (N_2136,N_162,N_209);
or U2137 (N_2137,N_759,N_1381);
and U2138 (N_2138,N_508,N_1001);
or U2139 (N_2139,N_168,N_647);
nand U2140 (N_2140,N_402,N_290);
nor U2141 (N_2141,N_672,N_987);
nand U2142 (N_2142,N_995,N_494);
or U2143 (N_2143,N_252,N_1030);
nand U2144 (N_2144,N_842,N_1430);
and U2145 (N_2145,N_1090,N_163);
nor U2146 (N_2146,N_565,N_367);
or U2147 (N_2147,N_1455,N_422);
or U2148 (N_2148,N_279,N_1114);
and U2149 (N_2149,N_1298,N_123);
nand U2150 (N_2150,N_871,N_766);
xor U2151 (N_2151,N_1247,N_1239);
xor U2152 (N_2152,N_860,N_515);
nor U2153 (N_2153,N_346,N_49);
nor U2154 (N_2154,N_1380,N_183);
and U2155 (N_2155,N_874,N_572);
xnor U2156 (N_2156,N_1073,N_758);
or U2157 (N_2157,N_776,N_824);
or U2158 (N_2158,N_1487,N_786);
or U2159 (N_2159,N_109,N_1348);
or U2160 (N_2160,N_388,N_915);
and U2161 (N_2161,N_43,N_597);
xor U2162 (N_2162,N_126,N_898);
and U2163 (N_2163,N_884,N_8);
or U2164 (N_2164,N_1337,N_1497);
and U2165 (N_2165,N_843,N_104);
or U2166 (N_2166,N_1416,N_711);
nor U2167 (N_2167,N_1256,N_696);
or U2168 (N_2168,N_715,N_750);
or U2169 (N_2169,N_167,N_1447);
or U2170 (N_2170,N_216,N_816);
nand U2171 (N_2171,N_687,N_985);
nor U2172 (N_2172,N_1258,N_1450);
and U2173 (N_2173,N_556,N_1189);
or U2174 (N_2174,N_1199,N_343);
xor U2175 (N_2175,N_1053,N_19);
and U2176 (N_2176,N_161,N_767);
nand U2177 (N_2177,N_1385,N_1355);
and U2178 (N_2178,N_808,N_1077);
and U2179 (N_2179,N_1397,N_37);
nand U2180 (N_2180,N_1491,N_60);
and U2181 (N_2181,N_1028,N_237);
or U2182 (N_2182,N_34,N_310);
nor U2183 (N_2183,N_1202,N_1206);
or U2184 (N_2184,N_917,N_664);
nor U2185 (N_2185,N_1048,N_70);
and U2186 (N_2186,N_224,N_595);
and U2187 (N_2187,N_87,N_1352);
nand U2188 (N_2188,N_228,N_136);
nor U2189 (N_2189,N_940,N_160);
or U2190 (N_2190,N_1267,N_1112);
or U2191 (N_2191,N_1025,N_83);
or U2192 (N_2192,N_820,N_684);
nand U2193 (N_2193,N_502,N_984);
or U2194 (N_2194,N_1181,N_1283);
or U2195 (N_2195,N_1062,N_1157);
nand U2196 (N_2196,N_403,N_470);
or U2197 (N_2197,N_549,N_810);
nor U2198 (N_2198,N_1426,N_1301);
xor U2199 (N_2199,N_1318,N_492);
or U2200 (N_2200,N_974,N_900);
or U2201 (N_2201,N_567,N_257);
nand U2202 (N_2202,N_976,N_392);
and U2203 (N_2203,N_1338,N_1396);
nand U2204 (N_2204,N_694,N_890);
xor U2205 (N_2205,N_932,N_1047);
and U2206 (N_2206,N_692,N_1216);
xor U2207 (N_2207,N_428,N_896);
or U2208 (N_2208,N_1341,N_1367);
and U2209 (N_2209,N_401,N_994);
xnor U2210 (N_2210,N_1059,N_930);
nor U2211 (N_2211,N_1052,N_144);
nor U2212 (N_2212,N_293,N_1119);
nand U2213 (N_2213,N_1128,N_1312);
or U2214 (N_2214,N_773,N_117);
nor U2215 (N_2215,N_103,N_211);
or U2216 (N_2216,N_1401,N_378);
nand U2217 (N_2217,N_491,N_603);
and U2218 (N_2218,N_484,N_1377);
or U2219 (N_2219,N_384,N_1144);
nand U2220 (N_2220,N_58,N_453);
or U2221 (N_2221,N_1036,N_1029);
and U2222 (N_2222,N_1253,N_514);
or U2223 (N_2223,N_855,N_48);
and U2224 (N_2224,N_435,N_699);
or U2225 (N_2225,N_1471,N_1349);
nor U2226 (N_2226,N_282,N_643);
or U2227 (N_2227,N_1371,N_1246);
xnor U2228 (N_2228,N_1172,N_62);
xor U2229 (N_2229,N_529,N_185);
nor U2230 (N_2230,N_489,N_911);
and U2231 (N_2231,N_777,N_50);
or U2232 (N_2232,N_1017,N_757);
xor U2233 (N_2233,N_1226,N_1195);
nand U2234 (N_2234,N_65,N_40);
xor U2235 (N_2235,N_335,N_212);
nand U2236 (N_2236,N_950,N_449);
and U2237 (N_2237,N_1493,N_1249);
nand U2238 (N_2238,N_763,N_701);
and U2239 (N_2239,N_1479,N_739);
nor U2240 (N_2240,N_1383,N_1374);
nor U2241 (N_2241,N_1270,N_1095);
xor U2242 (N_2242,N_1080,N_155);
or U2243 (N_2243,N_1411,N_754);
and U2244 (N_2244,N_1405,N_680);
and U2245 (N_2245,N_1378,N_1135);
nor U2246 (N_2246,N_649,N_1462);
nand U2247 (N_2247,N_897,N_1143);
nor U2248 (N_2248,N_498,N_227);
or U2249 (N_2249,N_1353,N_488);
and U2250 (N_2250,N_216,N_57);
or U2251 (N_2251,N_1202,N_681);
nand U2252 (N_2252,N_548,N_356);
and U2253 (N_2253,N_999,N_1286);
or U2254 (N_2254,N_231,N_1113);
nand U2255 (N_2255,N_166,N_684);
and U2256 (N_2256,N_294,N_28);
and U2257 (N_2257,N_502,N_948);
or U2258 (N_2258,N_687,N_330);
or U2259 (N_2259,N_1013,N_1087);
or U2260 (N_2260,N_470,N_948);
nor U2261 (N_2261,N_1219,N_321);
nor U2262 (N_2262,N_806,N_297);
or U2263 (N_2263,N_1063,N_1351);
and U2264 (N_2264,N_1130,N_337);
nand U2265 (N_2265,N_447,N_344);
and U2266 (N_2266,N_500,N_998);
nand U2267 (N_2267,N_793,N_374);
and U2268 (N_2268,N_561,N_130);
nor U2269 (N_2269,N_126,N_138);
or U2270 (N_2270,N_546,N_1169);
or U2271 (N_2271,N_936,N_1240);
and U2272 (N_2272,N_732,N_243);
nand U2273 (N_2273,N_1357,N_1201);
nand U2274 (N_2274,N_719,N_219);
nor U2275 (N_2275,N_298,N_231);
or U2276 (N_2276,N_1289,N_1258);
and U2277 (N_2277,N_816,N_1022);
or U2278 (N_2278,N_128,N_968);
and U2279 (N_2279,N_1425,N_971);
and U2280 (N_2280,N_126,N_337);
nor U2281 (N_2281,N_1302,N_66);
nor U2282 (N_2282,N_959,N_1278);
xor U2283 (N_2283,N_527,N_518);
nor U2284 (N_2284,N_178,N_584);
and U2285 (N_2285,N_510,N_530);
nand U2286 (N_2286,N_230,N_1471);
or U2287 (N_2287,N_498,N_910);
and U2288 (N_2288,N_741,N_469);
xnor U2289 (N_2289,N_275,N_992);
and U2290 (N_2290,N_885,N_446);
nand U2291 (N_2291,N_680,N_90);
nor U2292 (N_2292,N_601,N_115);
and U2293 (N_2293,N_1467,N_26);
nor U2294 (N_2294,N_1418,N_1440);
nand U2295 (N_2295,N_347,N_350);
nand U2296 (N_2296,N_833,N_814);
and U2297 (N_2297,N_1173,N_1457);
nor U2298 (N_2298,N_1230,N_1033);
xor U2299 (N_2299,N_302,N_1386);
and U2300 (N_2300,N_237,N_706);
nand U2301 (N_2301,N_1384,N_1499);
nand U2302 (N_2302,N_256,N_345);
or U2303 (N_2303,N_804,N_493);
and U2304 (N_2304,N_1035,N_646);
and U2305 (N_2305,N_481,N_877);
nand U2306 (N_2306,N_416,N_1351);
and U2307 (N_2307,N_1386,N_1200);
nand U2308 (N_2308,N_1353,N_1164);
and U2309 (N_2309,N_1060,N_413);
nand U2310 (N_2310,N_717,N_593);
or U2311 (N_2311,N_1410,N_674);
nand U2312 (N_2312,N_1418,N_1235);
or U2313 (N_2313,N_1116,N_837);
nand U2314 (N_2314,N_1249,N_1182);
nor U2315 (N_2315,N_1424,N_244);
nand U2316 (N_2316,N_1113,N_161);
nor U2317 (N_2317,N_1007,N_1101);
nor U2318 (N_2318,N_239,N_1456);
xnor U2319 (N_2319,N_842,N_871);
or U2320 (N_2320,N_897,N_383);
or U2321 (N_2321,N_1119,N_700);
or U2322 (N_2322,N_136,N_1469);
nand U2323 (N_2323,N_284,N_442);
xor U2324 (N_2324,N_65,N_756);
or U2325 (N_2325,N_1209,N_1213);
nor U2326 (N_2326,N_928,N_810);
nor U2327 (N_2327,N_883,N_617);
nand U2328 (N_2328,N_37,N_80);
and U2329 (N_2329,N_987,N_750);
nor U2330 (N_2330,N_356,N_1102);
or U2331 (N_2331,N_1033,N_1247);
xor U2332 (N_2332,N_1022,N_1246);
xor U2333 (N_2333,N_329,N_308);
nor U2334 (N_2334,N_612,N_1161);
nor U2335 (N_2335,N_520,N_9);
nor U2336 (N_2336,N_720,N_0);
nor U2337 (N_2337,N_1200,N_1170);
nor U2338 (N_2338,N_799,N_560);
and U2339 (N_2339,N_378,N_400);
nand U2340 (N_2340,N_1449,N_1293);
and U2341 (N_2341,N_860,N_1148);
and U2342 (N_2342,N_1477,N_256);
xor U2343 (N_2343,N_923,N_595);
nand U2344 (N_2344,N_814,N_1237);
xor U2345 (N_2345,N_967,N_190);
and U2346 (N_2346,N_1266,N_1201);
nand U2347 (N_2347,N_144,N_283);
and U2348 (N_2348,N_1232,N_764);
and U2349 (N_2349,N_854,N_509);
nand U2350 (N_2350,N_1129,N_1067);
nor U2351 (N_2351,N_990,N_764);
nand U2352 (N_2352,N_317,N_132);
or U2353 (N_2353,N_1201,N_6);
or U2354 (N_2354,N_438,N_1425);
or U2355 (N_2355,N_580,N_1009);
or U2356 (N_2356,N_691,N_1001);
and U2357 (N_2357,N_346,N_1139);
and U2358 (N_2358,N_57,N_1165);
or U2359 (N_2359,N_900,N_90);
nand U2360 (N_2360,N_327,N_1270);
or U2361 (N_2361,N_1451,N_263);
nand U2362 (N_2362,N_866,N_614);
nand U2363 (N_2363,N_874,N_1175);
nand U2364 (N_2364,N_45,N_66);
or U2365 (N_2365,N_1256,N_1052);
nor U2366 (N_2366,N_899,N_523);
xor U2367 (N_2367,N_1403,N_542);
and U2368 (N_2368,N_1347,N_995);
and U2369 (N_2369,N_1369,N_1393);
nand U2370 (N_2370,N_506,N_262);
nand U2371 (N_2371,N_1110,N_1429);
and U2372 (N_2372,N_1247,N_1103);
nor U2373 (N_2373,N_1409,N_873);
or U2374 (N_2374,N_239,N_1274);
or U2375 (N_2375,N_1059,N_100);
nor U2376 (N_2376,N_663,N_1249);
nand U2377 (N_2377,N_1497,N_984);
and U2378 (N_2378,N_1031,N_190);
xor U2379 (N_2379,N_735,N_1380);
and U2380 (N_2380,N_1185,N_296);
or U2381 (N_2381,N_241,N_338);
or U2382 (N_2382,N_1112,N_1476);
and U2383 (N_2383,N_825,N_83);
and U2384 (N_2384,N_462,N_1216);
nor U2385 (N_2385,N_413,N_346);
and U2386 (N_2386,N_1276,N_1401);
or U2387 (N_2387,N_141,N_800);
xnor U2388 (N_2388,N_397,N_344);
or U2389 (N_2389,N_1273,N_616);
or U2390 (N_2390,N_60,N_1136);
xnor U2391 (N_2391,N_939,N_541);
or U2392 (N_2392,N_1127,N_607);
or U2393 (N_2393,N_574,N_332);
nor U2394 (N_2394,N_600,N_546);
and U2395 (N_2395,N_530,N_527);
nand U2396 (N_2396,N_881,N_1467);
and U2397 (N_2397,N_1373,N_1432);
or U2398 (N_2398,N_1197,N_557);
xnor U2399 (N_2399,N_418,N_122);
nor U2400 (N_2400,N_1387,N_81);
nand U2401 (N_2401,N_623,N_867);
nor U2402 (N_2402,N_1362,N_872);
nand U2403 (N_2403,N_320,N_497);
nor U2404 (N_2404,N_823,N_1128);
nand U2405 (N_2405,N_457,N_1017);
nand U2406 (N_2406,N_1358,N_347);
or U2407 (N_2407,N_999,N_269);
or U2408 (N_2408,N_919,N_1146);
xor U2409 (N_2409,N_8,N_17);
and U2410 (N_2410,N_1493,N_1379);
or U2411 (N_2411,N_129,N_1205);
nand U2412 (N_2412,N_681,N_1085);
and U2413 (N_2413,N_753,N_704);
or U2414 (N_2414,N_1366,N_608);
nand U2415 (N_2415,N_46,N_105);
nor U2416 (N_2416,N_137,N_1454);
nor U2417 (N_2417,N_189,N_714);
xor U2418 (N_2418,N_1384,N_303);
nand U2419 (N_2419,N_245,N_504);
or U2420 (N_2420,N_638,N_1274);
nor U2421 (N_2421,N_274,N_437);
or U2422 (N_2422,N_482,N_7);
xnor U2423 (N_2423,N_326,N_1151);
xnor U2424 (N_2424,N_1104,N_964);
nand U2425 (N_2425,N_1276,N_719);
nor U2426 (N_2426,N_356,N_249);
and U2427 (N_2427,N_244,N_1264);
nor U2428 (N_2428,N_504,N_969);
xnor U2429 (N_2429,N_1477,N_108);
nand U2430 (N_2430,N_1346,N_997);
nor U2431 (N_2431,N_1119,N_387);
and U2432 (N_2432,N_1061,N_868);
xor U2433 (N_2433,N_852,N_71);
and U2434 (N_2434,N_693,N_1328);
nand U2435 (N_2435,N_451,N_539);
nand U2436 (N_2436,N_516,N_1309);
or U2437 (N_2437,N_545,N_276);
or U2438 (N_2438,N_440,N_460);
nor U2439 (N_2439,N_969,N_1312);
nor U2440 (N_2440,N_601,N_1467);
or U2441 (N_2441,N_1453,N_1013);
nor U2442 (N_2442,N_1102,N_849);
nor U2443 (N_2443,N_191,N_1108);
nand U2444 (N_2444,N_299,N_336);
nor U2445 (N_2445,N_181,N_425);
or U2446 (N_2446,N_1247,N_485);
xnor U2447 (N_2447,N_1401,N_631);
or U2448 (N_2448,N_451,N_702);
xor U2449 (N_2449,N_639,N_418);
or U2450 (N_2450,N_828,N_1056);
nand U2451 (N_2451,N_1478,N_1354);
and U2452 (N_2452,N_545,N_912);
or U2453 (N_2453,N_652,N_947);
and U2454 (N_2454,N_1474,N_463);
and U2455 (N_2455,N_1129,N_413);
or U2456 (N_2456,N_476,N_1063);
or U2457 (N_2457,N_617,N_1231);
xnor U2458 (N_2458,N_1459,N_1117);
nor U2459 (N_2459,N_229,N_588);
nand U2460 (N_2460,N_1244,N_1262);
nor U2461 (N_2461,N_150,N_369);
or U2462 (N_2462,N_761,N_432);
nor U2463 (N_2463,N_877,N_128);
or U2464 (N_2464,N_1100,N_286);
and U2465 (N_2465,N_506,N_49);
and U2466 (N_2466,N_159,N_151);
and U2467 (N_2467,N_452,N_1166);
nand U2468 (N_2468,N_1259,N_690);
nor U2469 (N_2469,N_1239,N_186);
and U2470 (N_2470,N_833,N_414);
nand U2471 (N_2471,N_394,N_1131);
nor U2472 (N_2472,N_1111,N_196);
xnor U2473 (N_2473,N_1195,N_1184);
and U2474 (N_2474,N_855,N_30);
and U2475 (N_2475,N_1216,N_1121);
and U2476 (N_2476,N_841,N_1144);
and U2477 (N_2477,N_51,N_1346);
and U2478 (N_2478,N_1381,N_1392);
or U2479 (N_2479,N_1260,N_855);
nor U2480 (N_2480,N_1336,N_923);
or U2481 (N_2481,N_442,N_673);
nor U2482 (N_2482,N_787,N_936);
or U2483 (N_2483,N_717,N_1002);
or U2484 (N_2484,N_712,N_413);
nand U2485 (N_2485,N_1162,N_151);
nor U2486 (N_2486,N_1462,N_759);
nor U2487 (N_2487,N_272,N_169);
and U2488 (N_2488,N_147,N_1209);
nor U2489 (N_2489,N_1313,N_93);
and U2490 (N_2490,N_943,N_320);
xor U2491 (N_2491,N_1470,N_613);
nor U2492 (N_2492,N_248,N_293);
or U2493 (N_2493,N_526,N_597);
nand U2494 (N_2494,N_1334,N_981);
xnor U2495 (N_2495,N_1414,N_397);
or U2496 (N_2496,N_1054,N_911);
nor U2497 (N_2497,N_619,N_995);
or U2498 (N_2498,N_515,N_539);
nand U2499 (N_2499,N_950,N_660);
nand U2500 (N_2500,N_1435,N_864);
nand U2501 (N_2501,N_490,N_796);
or U2502 (N_2502,N_452,N_1196);
or U2503 (N_2503,N_602,N_709);
nor U2504 (N_2504,N_1152,N_157);
nor U2505 (N_2505,N_604,N_190);
nor U2506 (N_2506,N_892,N_881);
xnor U2507 (N_2507,N_794,N_332);
nand U2508 (N_2508,N_638,N_175);
and U2509 (N_2509,N_864,N_576);
and U2510 (N_2510,N_702,N_613);
nand U2511 (N_2511,N_106,N_224);
or U2512 (N_2512,N_726,N_466);
and U2513 (N_2513,N_1479,N_297);
and U2514 (N_2514,N_1299,N_910);
nor U2515 (N_2515,N_161,N_622);
nand U2516 (N_2516,N_22,N_374);
nor U2517 (N_2517,N_486,N_1160);
or U2518 (N_2518,N_144,N_1439);
or U2519 (N_2519,N_1037,N_230);
nand U2520 (N_2520,N_985,N_1071);
or U2521 (N_2521,N_475,N_495);
and U2522 (N_2522,N_1368,N_953);
or U2523 (N_2523,N_1356,N_1394);
and U2524 (N_2524,N_457,N_682);
nand U2525 (N_2525,N_1320,N_707);
nor U2526 (N_2526,N_1150,N_37);
xor U2527 (N_2527,N_926,N_756);
nand U2528 (N_2528,N_1283,N_449);
and U2529 (N_2529,N_1453,N_133);
nand U2530 (N_2530,N_1292,N_693);
or U2531 (N_2531,N_488,N_793);
nor U2532 (N_2532,N_176,N_17);
nand U2533 (N_2533,N_43,N_980);
xnor U2534 (N_2534,N_131,N_538);
and U2535 (N_2535,N_734,N_425);
nor U2536 (N_2536,N_1116,N_157);
xor U2537 (N_2537,N_1281,N_900);
and U2538 (N_2538,N_1246,N_331);
or U2539 (N_2539,N_439,N_537);
and U2540 (N_2540,N_862,N_370);
nor U2541 (N_2541,N_204,N_1262);
nor U2542 (N_2542,N_1004,N_410);
nand U2543 (N_2543,N_1128,N_587);
nor U2544 (N_2544,N_547,N_8);
nor U2545 (N_2545,N_61,N_586);
nand U2546 (N_2546,N_89,N_615);
or U2547 (N_2547,N_1306,N_649);
nand U2548 (N_2548,N_130,N_257);
or U2549 (N_2549,N_453,N_265);
or U2550 (N_2550,N_962,N_277);
or U2551 (N_2551,N_934,N_1042);
nor U2552 (N_2552,N_1081,N_749);
or U2553 (N_2553,N_567,N_712);
nor U2554 (N_2554,N_903,N_594);
nand U2555 (N_2555,N_379,N_783);
nor U2556 (N_2556,N_489,N_1201);
nand U2557 (N_2557,N_1443,N_1289);
and U2558 (N_2558,N_1380,N_680);
xnor U2559 (N_2559,N_809,N_172);
nand U2560 (N_2560,N_977,N_337);
nand U2561 (N_2561,N_121,N_1049);
or U2562 (N_2562,N_1132,N_943);
and U2563 (N_2563,N_76,N_768);
or U2564 (N_2564,N_958,N_831);
and U2565 (N_2565,N_224,N_107);
or U2566 (N_2566,N_982,N_278);
and U2567 (N_2567,N_636,N_590);
and U2568 (N_2568,N_1243,N_803);
nor U2569 (N_2569,N_980,N_1167);
nand U2570 (N_2570,N_1456,N_1102);
nor U2571 (N_2571,N_737,N_862);
nor U2572 (N_2572,N_259,N_993);
nor U2573 (N_2573,N_846,N_1125);
or U2574 (N_2574,N_274,N_1479);
nor U2575 (N_2575,N_717,N_932);
nor U2576 (N_2576,N_972,N_964);
or U2577 (N_2577,N_1334,N_258);
and U2578 (N_2578,N_1465,N_376);
and U2579 (N_2579,N_1278,N_192);
nor U2580 (N_2580,N_1455,N_133);
nand U2581 (N_2581,N_1174,N_450);
nand U2582 (N_2582,N_634,N_48);
and U2583 (N_2583,N_95,N_887);
nand U2584 (N_2584,N_833,N_308);
nand U2585 (N_2585,N_900,N_215);
and U2586 (N_2586,N_468,N_1400);
nor U2587 (N_2587,N_826,N_821);
or U2588 (N_2588,N_354,N_1295);
or U2589 (N_2589,N_763,N_1153);
and U2590 (N_2590,N_1099,N_106);
and U2591 (N_2591,N_1450,N_1051);
nor U2592 (N_2592,N_833,N_16);
nand U2593 (N_2593,N_312,N_879);
or U2594 (N_2594,N_1315,N_756);
nand U2595 (N_2595,N_1071,N_1334);
nor U2596 (N_2596,N_470,N_345);
nand U2597 (N_2597,N_490,N_308);
nor U2598 (N_2598,N_513,N_842);
or U2599 (N_2599,N_306,N_784);
or U2600 (N_2600,N_899,N_464);
nor U2601 (N_2601,N_1493,N_1053);
or U2602 (N_2602,N_925,N_996);
and U2603 (N_2603,N_1441,N_736);
or U2604 (N_2604,N_1383,N_703);
nor U2605 (N_2605,N_1141,N_1015);
nand U2606 (N_2606,N_257,N_353);
or U2607 (N_2607,N_931,N_661);
xor U2608 (N_2608,N_1051,N_1027);
and U2609 (N_2609,N_1154,N_506);
or U2610 (N_2610,N_861,N_600);
nand U2611 (N_2611,N_46,N_936);
or U2612 (N_2612,N_1092,N_837);
or U2613 (N_2613,N_283,N_68);
xnor U2614 (N_2614,N_1478,N_1447);
xor U2615 (N_2615,N_664,N_768);
nand U2616 (N_2616,N_1250,N_1354);
and U2617 (N_2617,N_807,N_1416);
or U2618 (N_2618,N_1002,N_51);
nor U2619 (N_2619,N_84,N_1433);
nand U2620 (N_2620,N_59,N_1312);
xnor U2621 (N_2621,N_1338,N_178);
nor U2622 (N_2622,N_789,N_1072);
nor U2623 (N_2623,N_477,N_356);
or U2624 (N_2624,N_1385,N_427);
nand U2625 (N_2625,N_1386,N_444);
nand U2626 (N_2626,N_905,N_73);
or U2627 (N_2627,N_268,N_530);
or U2628 (N_2628,N_480,N_143);
or U2629 (N_2629,N_1447,N_258);
xnor U2630 (N_2630,N_992,N_972);
nand U2631 (N_2631,N_269,N_457);
nand U2632 (N_2632,N_1324,N_1274);
xnor U2633 (N_2633,N_227,N_119);
nor U2634 (N_2634,N_1128,N_1417);
and U2635 (N_2635,N_1050,N_1152);
nor U2636 (N_2636,N_189,N_1455);
or U2637 (N_2637,N_1424,N_721);
nor U2638 (N_2638,N_572,N_980);
xor U2639 (N_2639,N_1494,N_857);
nand U2640 (N_2640,N_1492,N_58);
xnor U2641 (N_2641,N_126,N_731);
or U2642 (N_2642,N_895,N_1001);
nand U2643 (N_2643,N_270,N_938);
nand U2644 (N_2644,N_1478,N_556);
or U2645 (N_2645,N_266,N_850);
and U2646 (N_2646,N_657,N_1232);
or U2647 (N_2647,N_1228,N_8);
nor U2648 (N_2648,N_1258,N_73);
and U2649 (N_2649,N_1425,N_12);
xor U2650 (N_2650,N_536,N_315);
and U2651 (N_2651,N_824,N_773);
nor U2652 (N_2652,N_1334,N_1107);
and U2653 (N_2653,N_327,N_59);
nand U2654 (N_2654,N_374,N_647);
or U2655 (N_2655,N_1423,N_309);
nand U2656 (N_2656,N_916,N_240);
nand U2657 (N_2657,N_1273,N_39);
nor U2658 (N_2658,N_1000,N_987);
nor U2659 (N_2659,N_677,N_1385);
nand U2660 (N_2660,N_270,N_1386);
and U2661 (N_2661,N_1344,N_1242);
or U2662 (N_2662,N_1393,N_1435);
xor U2663 (N_2663,N_738,N_764);
nor U2664 (N_2664,N_935,N_230);
and U2665 (N_2665,N_1203,N_906);
and U2666 (N_2666,N_670,N_619);
and U2667 (N_2667,N_912,N_708);
and U2668 (N_2668,N_210,N_553);
nand U2669 (N_2669,N_60,N_586);
and U2670 (N_2670,N_748,N_835);
or U2671 (N_2671,N_1489,N_1126);
xor U2672 (N_2672,N_844,N_707);
nor U2673 (N_2673,N_327,N_374);
nor U2674 (N_2674,N_1265,N_755);
nand U2675 (N_2675,N_410,N_0);
nor U2676 (N_2676,N_931,N_144);
nand U2677 (N_2677,N_1071,N_1411);
nand U2678 (N_2678,N_57,N_1244);
xnor U2679 (N_2679,N_265,N_92);
or U2680 (N_2680,N_197,N_630);
nor U2681 (N_2681,N_531,N_791);
or U2682 (N_2682,N_712,N_1257);
nor U2683 (N_2683,N_1329,N_755);
or U2684 (N_2684,N_602,N_1358);
and U2685 (N_2685,N_1403,N_698);
or U2686 (N_2686,N_60,N_115);
nand U2687 (N_2687,N_786,N_956);
nand U2688 (N_2688,N_1205,N_525);
and U2689 (N_2689,N_1062,N_529);
nand U2690 (N_2690,N_277,N_502);
and U2691 (N_2691,N_301,N_461);
or U2692 (N_2692,N_843,N_1410);
or U2693 (N_2693,N_1062,N_829);
and U2694 (N_2694,N_757,N_720);
and U2695 (N_2695,N_264,N_1417);
and U2696 (N_2696,N_1329,N_951);
xor U2697 (N_2697,N_1437,N_1215);
nand U2698 (N_2698,N_1079,N_1036);
nand U2699 (N_2699,N_527,N_2);
or U2700 (N_2700,N_960,N_659);
xor U2701 (N_2701,N_608,N_1077);
and U2702 (N_2702,N_202,N_1457);
or U2703 (N_2703,N_1059,N_651);
nand U2704 (N_2704,N_365,N_708);
or U2705 (N_2705,N_728,N_203);
and U2706 (N_2706,N_624,N_1149);
and U2707 (N_2707,N_1180,N_634);
nand U2708 (N_2708,N_911,N_494);
nand U2709 (N_2709,N_1110,N_901);
nor U2710 (N_2710,N_1144,N_703);
and U2711 (N_2711,N_1476,N_477);
nor U2712 (N_2712,N_943,N_726);
xnor U2713 (N_2713,N_223,N_354);
nand U2714 (N_2714,N_1336,N_161);
xnor U2715 (N_2715,N_1259,N_701);
xor U2716 (N_2716,N_904,N_16);
xor U2717 (N_2717,N_250,N_991);
or U2718 (N_2718,N_1326,N_24);
nor U2719 (N_2719,N_635,N_911);
and U2720 (N_2720,N_390,N_818);
and U2721 (N_2721,N_729,N_961);
and U2722 (N_2722,N_1334,N_1220);
and U2723 (N_2723,N_842,N_1480);
nor U2724 (N_2724,N_2,N_1228);
or U2725 (N_2725,N_55,N_452);
and U2726 (N_2726,N_1148,N_1030);
nor U2727 (N_2727,N_965,N_137);
nor U2728 (N_2728,N_887,N_1149);
or U2729 (N_2729,N_146,N_1478);
or U2730 (N_2730,N_1214,N_750);
and U2731 (N_2731,N_433,N_1414);
nor U2732 (N_2732,N_1444,N_1029);
and U2733 (N_2733,N_1307,N_506);
or U2734 (N_2734,N_706,N_91);
and U2735 (N_2735,N_381,N_729);
or U2736 (N_2736,N_540,N_1314);
or U2737 (N_2737,N_1024,N_696);
or U2738 (N_2738,N_984,N_1414);
nor U2739 (N_2739,N_555,N_18);
and U2740 (N_2740,N_690,N_1189);
nand U2741 (N_2741,N_1061,N_348);
and U2742 (N_2742,N_450,N_211);
nor U2743 (N_2743,N_1149,N_1483);
nor U2744 (N_2744,N_1083,N_741);
nor U2745 (N_2745,N_437,N_746);
nand U2746 (N_2746,N_576,N_1144);
nand U2747 (N_2747,N_218,N_1488);
and U2748 (N_2748,N_684,N_1220);
nand U2749 (N_2749,N_1435,N_1063);
nand U2750 (N_2750,N_208,N_126);
or U2751 (N_2751,N_1344,N_1311);
and U2752 (N_2752,N_791,N_394);
nor U2753 (N_2753,N_1406,N_969);
or U2754 (N_2754,N_574,N_598);
or U2755 (N_2755,N_1442,N_1091);
and U2756 (N_2756,N_1100,N_380);
nor U2757 (N_2757,N_43,N_695);
or U2758 (N_2758,N_1113,N_1189);
and U2759 (N_2759,N_1010,N_1210);
nand U2760 (N_2760,N_311,N_1095);
nand U2761 (N_2761,N_235,N_245);
nor U2762 (N_2762,N_1457,N_1390);
nor U2763 (N_2763,N_1362,N_808);
nor U2764 (N_2764,N_1194,N_547);
xnor U2765 (N_2765,N_423,N_882);
nand U2766 (N_2766,N_1293,N_1094);
nand U2767 (N_2767,N_185,N_1055);
xnor U2768 (N_2768,N_866,N_87);
xnor U2769 (N_2769,N_84,N_272);
nor U2770 (N_2770,N_660,N_974);
or U2771 (N_2771,N_796,N_286);
nand U2772 (N_2772,N_710,N_374);
nor U2773 (N_2773,N_876,N_1088);
and U2774 (N_2774,N_1228,N_924);
xor U2775 (N_2775,N_1375,N_1279);
nand U2776 (N_2776,N_1127,N_679);
nor U2777 (N_2777,N_235,N_907);
xnor U2778 (N_2778,N_109,N_552);
and U2779 (N_2779,N_800,N_348);
or U2780 (N_2780,N_1184,N_1381);
or U2781 (N_2781,N_392,N_964);
nor U2782 (N_2782,N_1157,N_1279);
or U2783 (N_2783,N_711,N_475);
nor U2784 (N_2784,N_12,N_1359);
nand U2785 (N_2785,N_1149,N_1331);
and U2786 (N_2786,N_1114,N_672);
xor U2787 (N_2787,N_970,N_766);
and U2788 (N_2788,N_995,N_1045);
or U2789 (N_2789,N_550,N_1386);
nand U2790 (N_2790,N_1322,N_714);
xor U2791 (N_2791,N_842,N_1477);
nand U2792 (N_2792,N_211,N_686);
nand U2793 (N_2793,N_1237,N_731);
or U2794 (N_2794,N_614,N_157);
nor U2795 (N_2795,N_1321,N_1149);
and U2796 (N_2796,N_463,N_811);
nor U2797 (N_2797,N_168,N_907);
nand U2798 (N_2798,N_417,N_1239);
and U2799 (N_2799,N_245,N_509);
or U2800 (N_2800,N_703,N_973);
nand U2801 (N_2801,N_858,N_1090);
or U2802 (N_2802,N_1313,N_636);
and U2803 (N_2803,N_382,N_426);
and U2804 (N_2804,N_1294,N_1115);
nor U2805 (N_2805,N_380,N_1395);
nand U2806 (N_2806,N_1221,N_109);
and U2807 (N_2807,N_25,N_237);
nand U2808 (N_2808,N_1406,N_1186);
or U2809 (N_2809,N_358,N_1410);
nor U2810 (N_2810,N_640,N_661);
and U2811 (N_2811,N_427,N_1414);
and U2812 (N_2812,N_1249,N_1209);
nor U2813 (N_2813,N_1377,N_397);
or U2814 (N_2814,N_1103,N_467);
or U2815 (N_2815,N_1106,N_753);
or U2816 (N_2816,N_430,N_1240);
nand U2817 (N_2817,N_460,N_683);
or U2818 (N_2818,N_1450,N_1058);
nor U2819 (N_2819,N_1370,N_179);
nor U2820 (N_2820,N_539,N_634);
nor U2821 (N_2821,N_261,N_449);
nor U2822 (N_2822,N_1241,N_1090);
nor U2823 (N_2823,N_455,N_1012);
nor U2824 (N_2824,N_649,N_497);
and U2825 (N_2825,N_143,N_157);
nand U2826 (N_2826,N_348,N_7);
and U2827 (N_2827,N_1015,N_1371);
nand U2828 (N_2828,N_138,N_256);
nor U2829 (N_2829,N_163,N_638);
and U2830 (N_2830,N_1155,N_1317);
nor U2831 (N_2831,N_1167,N_1196);
nand U2832 (N_2832,N_928,N_1134);
or U2833 (N_2833,N_673,N_567);
and U2834 (N_2834,N_419,N_1436);
xor U2835 (N_2835,N_293,N_787);
nand U2836 (N_2836,N_90,N_1062);
xor U2837 (N_2837,N_1190,N_1412);
or U2838 (N_2838,N_323,N_333);
nor U2839 (N_2839,N_450,N_1256);
nor U2840 (N_2840,N_456,N_1015);
nand U2841 (N_2841,N_699,N_1346);
or U2842 (N_2842,N_1478,N_1126);
nor U2843 (N_2843,N_1192,N_544);
nand U2844 (N_2844,N_72,N_1051);
xnor U2845 (N_2845,N_441,N_733);
and U2846 (N_2846,N_1146,N_1138);
and U2847 (N_2847,N_759,N_1362);
and U2848 (N_2848,N_742,N_1084);
or U2849 (N_2849,N_900,N_1161);
and U2850 (N_2850,N_1361,N_617);
or U2851 (N_2851,N_798,N_1134);
nor U2852 (N_2852,N_1416,N_1003);
nand U2853 (N_2853,N_747,N_1202);
or U2854 (N_2854,N_827,N_1374);
and U2855 (N_2855,N_208,N_295);
nor U2856 (N_2856,N_806,N_1083);
nor U2857 (N_2857,N_759,N_829);
or U2858 (N_2858,N_707,N_801);
or U2859 (N_2859,N_1337,N_440);
xor U2860 (N_2860,N_802,N_1337);
nor U2861 (N_2861,N_575,N_1190);
and U2862 (N_2862,N_235,N_906);
and U2863 (N_2863,N_945,N_1313);
nor U2864 (N_2864,N_833,N_1380);
nand U2865 (N_2865,N_1239,N_414);
nand U2866 (N_2866,N_462,N_93);
xor U2867 (N_2867,N_1063,N_810);
nor U2868 (N_2868,N_476,N_679);
nand U2869 (N_2869,N_224,N_947);
xor U2870 (N_2870,N_1439,N_262);
or U2871 (N_2871,N_1498,N_627);
nand U2872 (N_2872,N_109,N_1411);
nand U2873 (N_2873,N_271,N_234);
and U2874 (N_2874,N_293,N_629);
nor U2875 (N_2875,N_83,N_885);
and U2876 (N_2876,N_526,N_571);
nand U2877 (N_2877,N_88,N_492);
nor U2878 (N_2878,N_1279,N_1462);
nor U2879 (N_2879,N_1247,N_1145);
or U2880 (N_2880,N_1280,N_1407);
or U2881 (N_2881,N_1200,N_446);
nor U2882 (N_2882,N_794,N_29);
nand U2883 (N_2883,N_80,N_1478);
and U2884 (N_2884,N_125,N_1033);
nand U2885 (N_2885,N_705,N_1117);
nand U2886 (N_2886,N_161,N_1036);
or U2887 (N_2887,N_1023,N_339);
xor U2888 (N_2888,N_1139,N_966);
and U2889 (N_2889,N_247,N_253);
nor U2890 (N_2890,N_926,N_1296);
nand U2891 (N_2891,N_530,N_638);
or U2892 (N_2892,N_171,N_384);
and U2893 (N_2893,N_792,N_223);
or U2894 (N_2894,N_480,N_375);
nor U2895 (N_2895,N_406,N_508);
nor U2896 (N_2896,N_854,N_296);
nor U2897 (N_2897,N_312,N_1199);
xnor U2898 (N_2898,N_1040,N_1246);
and U2899 (N_2899,N_1324,N_1157);
and U2900 (N_2900,N_878,N_270);
and U2901 (N_2901,N_1303,N_573);
nor U2902 (N_2902,N_531,N_566);
nor U2903 (N_2903,N_700,N_981);
nand U2904 (N_2904,N_586,N_365);
nor U2905 (N_2905,N_381,N_999);
and U2906 (N_2906,N_494,N_489);
nand U2907 (N_2907,N_86,N_1409);
or U2908 (N_2908,N_1401,N_1399);
xor U2909 (N_2909,N_1325,N_240);
and U2910 (N_2910,N_1206,N_746);
or U2911 (N_2911,N_847,N_914);
or U2912 (N_2912,N_135,N_214);
nand U2913 (N_2913,N_1308,N_978);
and U2914 (N_2914,N_345,N_633);
and U2915 (N_2915,N_1347,N_406);
and U2916 (N_2916,N_356,N_1495);
or U2917 (N_2917,N_339,N_1213);
nor U2918 (N_2918,N_641,N_960);
nand U2919 (N_2919,N_936,N_1179);
or U2920 (N_2920,N_181,N_723);
or U2921 (N_2921,N_1484,N_0);
and U2922 (N_2922,N_1217,N_329);
nand U2923 (N_2923,N_272,N_24);
or U2924 (N_2924,N_743,N_1328);
nor U2925 (N_2925,N_624,N_15);
and U2926 (N_2926,N_291,N_433);
nand U2927 (N_2927,N_337,N_153);
nor U2928 (N_2928,N_66,N_901);
or U2929 (N_2929,N_917,N_982);
and U2930 (N_2930,N_1100,N_1204);
nand U2931 (N_2931,N_1497,N_380);
and U2932 (N_2932,N_1367,N_976);
nor U2933 (N_2933,N_1159,N_794);
nand U2934 (N_2934,N_1274,N_629);
nand U2935 (N_2935,N_1229,N_630);
or U2936 (N_2936,N_189,N_242);
nor U2937 (N_2937,N_138,N_841);
nand U2938 (N_2938,N_847,N_750);
and U2939 (N_2939,N_883,N_714);
and U2940 (N_2940,N_909,N_905);
and U2941 (N_2941,N_732,N_1172);
and U2942 (N_2942,N_645,N_1315);
or U2943 (N_2943,N_864,N_759);
nand U2944 (N_2944,N_1034,N_280);
and U2945 (N_2945,N_1132,N_468);
nand U2946 (N_2946,N_1333,N_1109);
nand U2947 (N_2947,N_1235,N_300);
or U2948 (N_2948,N_731,N_950);
and U2949 (N_2949,N_1173,N_355);
nor U2950 (N_2950,N_418,N_1314);
nand U2951 (N_2951,N_936,N_168);
xnor U2952 (N_2952,N_1246,N_1480);
nand U2953 (N_2953,N_610,N_1120);
nor U2954 (N_2954,N_1344,N_1391);
xor U2955 (N_2955,N_675,N_615);
nand U2956 (N_2956,N_744,N_509);
nand U2957 (N_2957,N_723,N_315);
xnor U2958 (N_2958,N_541,N_5);
xor U2959 (N_2959,N_1230,N_390);
xnor U2960 (N_2960,N_1441,N_723);
and U2961 (N_2961,N_1212,N_1143);
and U2962 (N_2962,N_1179,N_893);
or U2963 (N_2963,N_548,N_1141);
and U2964 (N_2964,N_789,N_492);
nor U2965 (N_2965,N_1196,N_754);
nand U2966 (N_2966,N_1054,N_357);
nand U2967 (N_2967,N_184,N_1473);
or U2968 (N_2968,N_362,N_1164);
or U2969 (N_2969,N_1264,N_1102);
nor U2970 (N_2970,N_962,N_63);
nor U2971 (N_2971,N_1140,N_1015);
or U2972 (N_2972,N_648,N_249);
and U2973 (N_2973,N_690,N_32);
nand U2974 (N_2974,N_522,N_1315);
nor U2975 (N_2975,N_383,N_1214);
nand U2976 (N_2976,N_261,N_205);
nand U2977 (N_2977,N_322,N_1347);
and U2978 (N_2978,N_1448,N_45);
nand U2979 (N_2979,N_312,N_279);
nor U2980 (N_2980,N_904,N_982);
nor U2981 (N_2981,N_1433,N_192);
and U2982 (N_2982,N_1081,N_626);
or U2983 (N_2983,N_158,N_187);
or U2984 (N_2984,N_539,N_709);
or U2985 (N_2985,N_113,N_1142);
nor U2986 (N_2986,N_594,N_1493);
and U2987 (N_2987,N_546,N_1242);
and U2988 (N_2988,N_141,N_582);
or U2989 (N_2989,N_803,N_1154);
nor U2990 (N_2990,N_600,N_1160);
xnor U2991 (N_2991,N_391,N_1167);
nand U2992 (N_2992,N_837,N_1105);
nor U2993 (N_2993,N_122,N_1261);
xnor U2994 (N_2994,N_768,N_355);
or U2995 (N_2995,N_1207,N_1350);
or U2996 (N_2996,N_837,N_416);
nand U2997 (N_2997,N_301,N_709);
nor U2998 (N_2998,N_679,N_1213);
nor U2999 (N_2999,N_1319,N_741);
nand U3000 (N_3000,N_2337,N_2375);
and U3001 (N_3001,N_2409,N_1881);
or U3002 (N_3002,N_2436,N_2043);
or U3003 (N_3003,N_1931,N_2153);
nor U3004 (N_3004,N_2201,N_2020);
and U3005 (N_3005,N_2804,N_2574);
and U3006 (N_3006,N_1521,N_2262);
or U3007 (N_3007,N_2114,N_1919);
or U3008 (N_3008,N_2341,N_1866);
and U3009 (N_3009,N_1758,N_2744);
xnor U3010 (N_3010,N_2584,N_2921);
or U3011 (N_3011,N_1777,N_2297);
nand U3012 (N_3012,N_2031,N_1786);
and U3013 (N_3013,N_2887,N_2922);
and U3014 (N_3014,N_1699,N_1560);
and U3015 (N_3015,N_2325,N_2671);
or U3016 (N_3016,N_1981,N_2159);
and U3017 (N_3017,N_2801,N_2179);
nand U3018 (N_3018,N_2276,N_2902);
nor U3019 (N_3019,N_2663,N_2395);
or U3020 (N_3020,N_2401,N_2965);
nand U3021 (N_3021,N_2040,N_1679);
or U3022 (N_3022,N_1853,N_1558);
and U3023 (N_3023,N_1501,N_2996);
nand U3024 (N_3024,N_2165,N_2094);
or U3025 (N_3025,N_2431,N_2726);
nand U3026 (N_3026,N_2309,N_2277);
nor U3027 (N_3027,N_2974,N_2414);
nand U3028 (N_3028,N_2110,N_1988);
and U3029 (N_3029,N_2970,N_1604);
or U3030 (N_3030,N_2731,N_2077);
nor U3031 (N_3031,N_2381,N_1960);
nor U3032 (N_3032,N_2232,N_2346);
nor U3033 (N_3033,N_1536,N_2241);
xor U3034 (N_3034,N_2966,N_2925);
nor U3035 (N_3035,N_2670,N_2315);
nand U3036 (N_3036,N_2610,N_1606);
nor U3037 (N_3037,N_2454,N_1894);
and U3038 (N_3038,N_2724,N_2957);
or U3039 (N_3039,N_2131,N_2271);
nor U3040 (N_3040,N_2076,N_1792);
and U3041 (N_3041,N_2597,N_2356);
and U3042 (N_3042,N_2907,N_2591);
or U3043 (N_3043,N_2764,N_1909);
nor U3044 (N_3044,N_2013,N_2142);
or U3045 (N_3045,N_2893,N_2373);
nand U3046 (N_3046,N_2362,N_1599);
or U3047 (N_3047,N_2543,N_1936);
and U3048 (N_3048,N_1872,N_2419);
and U3049 (N_3049,N_2427,N_2856);
and U3050 (N_3050,N_1592,N_2377);
nor U3051 (N_3051,N_2439,N_2066);
nor U3052 (N_3052,N_2392,N_2188);
nand U3053 (N_3053,N_1889,N_1959);
or U3054 (N_3054,N_1736,N_2620);
or U3055 (N_3055,N_2548,N_1746);
xnor U3056 (N_3056,N_2545,N_1913);
nor U3057 (N_3057,N_2184,N_2060);
and U3058 (N_3058,N_2983,N_1554);
xnor U3059 (N_3059,N_1682,N_1581);
xnor U3060 (N_3060,N_1869,N_2446);
or U3061 (N_3061,N_2552,N_2187);
nand U3062 (N_3062,N_1624,N_2499);
nor U3063 (N_3063,N_2012,N_1979);
or U3064 (N_3064,N_2960,N_2803);
nand U3065 (N_3065,N_2448,N_2068);
and U3066 (N_3066,N_1769,N_2929);
xnor U3067 (N_3067,N_2511,N_1993);
nand U3068 (N_3068,N_2604,N_1755);
nor U3069 (N_3069,N_1867,N_2927);
and U3070 (N_3070,N_2776,N_2593);
xnor U3071 (N_3071,N_2127,N_2169);
and U3072 (N_3072,N_2123,N_2898);
nor U3073 (N_3073,N_1731,N_2816);
and U3074 (N_3074,N_2483,N_2254);
nand U3075 (N_3075,N_2083,N_1799);
nor U3076 (N_3076,N_2949,N_2659);
or U3077 (N_3077,N_2716,N_2273);
and U3078 (N_3078,N_1659,N_2697);
nor U3079 (N_3079,N_1984,N_1669);
nor U3080 (N_3080,N_2458,N_2197);
nand U3081 (N_3081,N_2476,N_1636);
and U3082 (N_3082,N_2000,N_1626);
nor U3083 (N_3083,N_2494,N_2952);
xor U3084 (N_3084,N_1531,N_1875);
nand U3085 (N_3085,N_2363,N_2553);
and U3086 (N_3086,N_1857,N_1500);
nand U3087 (N_3087,N_1818,N_2866);
xor U3088 (N_3088,N_2986,N_1610);
or U3089 (N_3089,N_1963,N_1860);
nand U3090 (N_3090,N_1762,N_1822);
nor U3091 (N_3091,N_2836,N_2531);
nor U3092 (N_3092,N_1635,N_2332);
or U3093 (N_3093,N_2979,N_1790);
or U3094 (N_3094,N_2585,N_1888);
nor U3095 (N_3095,N_1874,N_1575);
nor U3096 (N_3096,N_2438,N_2738);
xor U3097 (N_3097,N_2781,N_2529);
and U3098 (N_3098,N_2871,N_2528);
nor U3099 (N_3099,N_1905,N_2581);
or U3100 (N_3100,N_1961,N_2735);
xnor U3101 (N_3101,N_2256,N_2968);
nor U3102 (N_3102,N_2813,N_1706);
nor U3103 (N_3103,N_1847,N_1844);
xor U3104 (N_3104,N_2366,N_2486);
or U3105 (N_3105,N_2025,N_1781);
or U3106 (N_3106,N_2238,N_1852);
nand U3107 (N_3107,N_2673,N_1780);
nor U3108 (N_3108,N_2630,N_2221);
nor U3109 (N_3109,N_1691,N_2089);
nor U3110 (N_3110,N_1672,N_2555);
nor U3111 (N_3111,N_2121,N_2030);
nand U3112 (N_3112,N_1942,N_1808);
or U3113 (N_3113,N_1851,N_2718);
or U3114 (N_3114,N_2074,N_2487);
and U3115 (N_3115,N_2041,N_2311);
nor U3116 (N_3116,N_1613,N_2765);
nor U3117 (N_3117,N_2888,N_2867);
nor U3118 (N_3118,N_2139,N_1548);
or U3119 (N_3119,N_2189,N_1897);
and U3120 (N_3120,N_2863,N_2705);
nor U3121 (N_3121,N_2666,N_1796);
or U3122 (N_3122,N_2444,N_1623);
or U3123 (N_3123,N_2513,N_2470);
and U3124 (N_3124,N_2795,N_1700);
nor U3125 (N_3125,N_2296,N_2194);
or U3126 (N_3126,N_1957,N_2044);
and U3127 (N_3127,N_2017,N_2371);
or U3128 (N_3128,N_1768,N_1764);
or U3129 (N_3129,N_1910,N_2707);
or U3130 (N_3130,N_2995,N_1681);
or U3131 (N_3131,N_2843,N_1650);
nor U3132 (N_3132,N_2293,N_2956);
nor U3133 (N_3133,N_2609,N_2643);
xor U3134 (N_3134,N_2834,N_1729);
nor U3135 (N_3135,N_2903,N_2980);
nor U3136 (N_3136,N_2561,N_2521);
or U3137 (N_3137,N_2096,N_2533);
nor U3138 (N_3138,N_2814,N_2632);
nor U3139 (N_3139,N_1696,N_1924);
nand U3140 (N_3140,N_2789,N_2938);
and U3141 (N_3141,N_1972,N_2291);
nand U3142 (N_3142,N_1564,N_2116);
nor U3143 (N_3143,N_2772,N_1773);
nand U3144 (N_3144,N_1983,N_1540);
or U3145 (N_3145,N_2876,N_2622);
or U3146 (N_3146,N_2474,N_2313);
and U3147 (N_3147,N_2991,N_1716);
or U3148 (N_3148,N_1666,N_1987);
nand U3149 (N_3149,N_2546,N_2879);
nand U3150 (N_3150,N_1520,N_2465);
nor U3151 (N_3151,N_2619,N_2092);
xnor U3152 (N_3152,N_1545,N_2605);
or U3153 (N_3153,N_2917,N_2481);
nor U3154 (N_3154,N_2695,N_2451);
nand U3155 (N_3155,N_2398,N_2248);
nand U3156 (N_3156,N_1783,N_1566);
and U3157 (N_3157,N_2336,N_1843);
xnor U3158 (N_3158,N_1589,N_2790);
nor U3159 (N_3159,N_1748,N_2421);
nand U3160 (N_3160,N_2088,N_1958);
nor U3161 (N_3161,N_1555,N_2576);
nand U3162 (N_3162,N_2894,N_1514);
or U3163 (N_3163,N_2640,N_2073);
nor U3164 (N_3164,N_2161,N_1649);
or U3165 (N_3165,N_2994,N_2785);
nor U3166 (N_3166,N_2100,N_2881);
nor U3167 (N_3167,N_1991,N_2330);
and U3168 (N_3168,N_2851,N_1864);
nor U3169 (N_3169,N_2450,N_2082);
nor U3170 (N_3170,N_1802,N_2459);
nand U3171 (N_3171,N_2386,N_2027);
nor U3172 (N_3172,N_2771,N_2149);
and U3173 (N_3173,N_1845,N_1761);
nor U3174 (N_3174,N_2655,N_2385);
and U3175 (N_3175,N_1590,N_1904);
nand U3176 (N_3176,N_2941,N_2207);
and U3177 (N_3177,N_1661,N_2146);
nand U3178 (N_3178,N_1718,N_1711);
nand U3179 (N_3179,N_2412,N_1891);
and U3180 (N_3180,N_2612,N_2274);
nand U3181 (N_3181,N_2407,N_2503);
nand U3182 (N_3182,N_2471,N_1600);
or U3183 (N_3183,N_2754,N_1738);
nor U3184 (N_3184,N_2777,N_2278);
nand U3185 (N_3185,N_1791,N_2302);
or U3186 (N_3186,N_1563,N_2572);
and U3187 (N_3187,N_1819,N_2455);
nand U3188 (N_3188,N_2406,N_2554);
nand U3189 (N_3189,N_2286,N_2259);
and U3190 (N_3190,N_2683,N_2512);
and U3191 (N_3191,N_2223,N_1879);
nor U3192 (N_3192,N_2239,N_2686);
nor U3193 (N_3193,N_2034,N_2825);
nand U3194 (N_3194,N_1788,N_1896);
xnor U3195 (N_3195,N_2024,N_1900);
nand U3196 (N_3196,N_2310,N_2509);
nor U3197 (N_3197,N_1982,N_1601);
nor U3198 (N_3198,N_2761,N_2099);
or U3199 (N_3199,N_2331,N_2987);
or U3200 (N_3200,N_2872,N_1974);
nand U3201 (N_3201,N_2323,N_2753);
xnor U3202 (N_3202,N_1975,N_2079);
or U3203 (N_3203,N_1719,N_2279);
nor U3204 (N_3204,N_1684,N_2954);
nor U3205 (N_3205,N_2452,N_2447);
and U3206 (N_3206,N_2711,N_2155);
or U3207 (N_3207,N_1577,N_1638);
and U3208 (N_3208,N_2069,N_2890);
nor U3209 (N_3209,N_1756,N_1932);
nor U3210 (N_3210,N_1651,N_1642);
and U3211 (N_3211,N_2918,N_2908);
nand U3212 (N_3212,N_1703,N_2618);
nand U3213 (N_3213,N_1929,N_1578);
or U3214 (N_3214,N_2992,N_1944);
nand U3215 (N_3215,N_2065,N_2281);
and U3216 (N_3216,N_2827,N_2896);
or U3217 (N_3217,N_2090,N_2958);
nor U3218 (N_3218,N_2226,N_2741);
or U3219 (N_3219,N_2947,N_2260);
nor U3220 (N_3220,N_1561,N_2018);
or U3221 (N_3221,N_1837,N_2607);
and U3222 (N_3222,N_1854,N_2157);
or U3223 (N_3223,N_2010,N_1992);
xnor U3224 (N_3224,N_2118,N_1953);
and U3225 (N_3225,N_2897,N_2886);
nor U3226 (N_3226,N_2299,N_2029);
or U3227 (N_3227,N_2147,N_2747);
and U3228 (N_3228,N_1705,N_2393);
or U3229 (N_3229,N_2294,N_1528);
nor U3230 (N_3230,N_1968,N_2782);
or U3231 (N_3231,N_1516,N_2959);
and U3232 (N_3232,N_2570,N_1625);
xor U3233 (N_3233,N_1620,N_2690);
nor U3234 (N_3234,N_2397,N_2849);
or U3235 (N_3235,N_1708,N_2931);
or U3236 (N_3236,N_1882,N_2773);
xor U3237 (N_3237,N_2823,N_2084);
nor U3238 (N_3238,N_1977,N_2878);
or U3239 (N_3239,N_2183,N_2768);
or U3240 (N_3240,N_2757,N_1573);
or U3241 (N_3241,N_1687,N_2687);
or U3242 (N_3242,N_2312,N_2339);
nor U3243 (N_3243,N_2300,N_2998);
and U3244 (N_3244,N_2535,N_1583);
nor U3245 (N_3245,N_2500,N_2936);
and U3246 (N_3246,N_2423,N_2829);
nor U3247 (N_3247,N_1933,N_1934);
and U3248 (N_3248,N_1701,N_2046);
and U3249 (N_3249,N_2517,N_2181);
and U3250 (N_3250,N_2045,N_1662);
or U3251 (N_3251,N_1774,N_1895);
nor U3252 (N_3252,N_1513,N_2853);
xnor U3253 (N_3253,N_1765,N_2490);
nor U3254 (N_3254,N_1943,N_1697);
nand U3255 (N_3255,N_2740,N_2178);
and U3256 (N_3256,N_2914,N_2091);
or U3257 (N_3257,N_2628,N_2793);
or U3258 (N_3258,N_1653,N_1937);
nor U3259 (N_3259,N_2399,N_2383);
nor U3260 (N_3260,N_2380,N_1996);
or U3261 (N_3261,N_2389,N_2348);
and U3262 (N_3262,N_2057,N_1926);
or U3263 (N_3263,N_2290,N_2767);
nand U3264 (N_3264,N_2345,N_2387);
nand U3265 (N_3265,N_1710,N_2606);
nand U3266 (N_3266,N_2493,N_2022);
and U3267 (N_3267,N_2463,N_2266);
nand U3268 (N_3268,N_2864,N_2963);
nor U3269 (N_3269,N_1525,N_2205);
nand U3270 (N_3270,N_1784,N_1743);
nor U3271 (N_3271,N_2847,N_2577);
nand U3272 (N_3272,N_2563,N_2441);
nand U3273 (N_3273,N_1886,N_1628);
and U3274 (N_3274,N_1643,N_1639);
or U3275 (N_3275,N_2435,N_1939);
xnor U3276 (N_3276,N_2404,N_1585);
nor U3277 (N_3277,N_2749,N_2520);
or U3278 (N_3278,N_2005,N_2176);
or U3279 (N_3279,N_2854,N_2275);
nor U3280 (N_3280,N_2304,N_2355);
xor U3281 (N_3281,N_1645,N_1817);
and U3282 (N_3282,N_2059,N_2478);
nand U3283 (N_3283,N_1771,N_2284);
nor U3284 (N_3284,N_2411,N_1546);
and U3285 (N_3285,N_1921,N_2138);
nor U3286 (N_3286,N_1749,N_2558);
xnor U3287 (N_3287,N_2006,N_1654);
nand U3288 (N_3288,N_2608,N_1720);
nor U3289 (N_3289,N_2562,N_2684);
and U3290 (N_3290,N_2725,N_2812);
nor U3291 (N_3291,N_2198,N_2261);
or U3292 (N_3292,N_2977,N_2722);
or U3293 (N_3293,N_2839,N_2353);
and U3294 (N_3294,N_2924,N_2811);
and U3295 (N_3295,N_2932,N_1778);
nand U3296 (N_3296,N_2358,N_1883);
or U3297 (N_3297,N_2955,N_2351);
xnor U3298 (N_3298,N_2728,N_2466);
nor U3299 (N_3299,N_2616,N_2685);
nor U3300 (N_3300,N_2115,N_2180);
and U3301 (N_3301,N_2243,N_2272);
or U3302 (N_3302,N_1805,N_2578);
or U3303 (N_3303,N_2085,N_1633);
nor U3304 (N_3304,N_2244,N_1734);
nand U3305 (N_3305,N_2942,N_1518);
nor U3306 (N_3306,N_2665,N_2587);
xnor U3307 (N_3307,N_2588,N_2301);
or U3308 (N_3308,N_2497,N_2442);
nand U3309 (N_3309,N_2703,N_2384);
xor U3310 (N_3310,N_1779,N_2743);
nand U3311 (N_3311,N_2733,N_1832);
or U3312 (N_3312,N_1775,N_2719);
or U3313 (N_3313,N_2349,N_1914);
and U3314 (N_3314,N_2095,N_2873);
xor U3315 (N_3315,N_1715,N_1925);
nor U3316 (N_3316,N_1787,N_2015);
nand U3317 (N_3317,N_2729,N_1693);
nand U3318 (N_3318,N_2850,N_2786);
and U3319 (N_3319,N_2694,N_2642);
xor U3320 (N_3320,N_2329,N_1807);
or U3321 (N_3321,N_1906,N_2857);
nand U3322 (N_3322,N_2717,N_2911);
nor U3323 (N_3323,N_2342,N_2318);
nor U3324 (N_3324,N_2920,N_1584);
xnor U3325 (N_3325,N_2571,N_2586);
and U3326 (N_3326,N_2210,N_1876);
xnor U3327 (N_3327,N_2048,N_1508);
nand U3328 (N_3328,N_1997,N_2388);
or U3329 (N_3329,N_2904,N_1688);
nor U3330 (N_3330,N_2805,N_2443);
nor U3331 (N_3331,N_2975,N_1967);
or U3332 (N_3332,N_2633,N_1709);
nor U3333 (N_3333,N_1795,N_2948);
and U3334 (N_3334,N_2997,N_2830);
nand U3335 (N_3335,N_2333,N_2255);
and U3336 (N_3336,N_2237,N_2328);
or U3337 (N_3337,N_2133,N_2564);
nand U3338 (N_3338,N_1782,N_2800);
nor U3339 (N_3339,N_2320,N_1752);
nor U3340 (N_3340,N_1702,N_1893);
nor U3341 (N_3341,N_1927,N_1800);
nand U3342 (N_3342,N_2762,N_2852);
or U3343 (N_3343,N_2219,N_1928);
xnor U3344 (N_3344,N_2658,N_2752);
xor U3345 (N_3345,N_2171,N_2602);
nand U3346 (N_3346,N_2540,N_1737);
and U3347 (N_3347,N_1814,N_2064);
nor U3348 (N_3348,N_2915,N_2787);
and U3349 (N_3349,N_2990,N_2295);
nor U3350 (N_3350,N_2837,N_1884);
and U3351 (N_3351,N_2425,N_1863);
and U3352 (N_3352,N_1732,N_2023);
nor U3353 (N_3353,N_2107,N_2322);
and U3354 (N_3354,N_2739,N_2208);
and U3355 (N_3355,N_1789,N_2168);
xor U3356 (N_3356,N_2748,N_2737);
and U3357 (N_3357,N_2527,N_1683);
nand U3358 (N_3358,N_1562,N_2242);
nor U3359 (N_3359,N_2473,N_1861);
xor U3360 (N_3360,N_2627,N_1603);
xor U3361 (N_3361,N_1949,N_1576);
or U3362 (N_3362,N_2750,N_2488);
nand U3363 (N_3363,N_1574,N_2334);
nor U3364 (N_3364,N_2360,N_2327);
nand U3365 (N_3365,N_2042,N_2506);
nor U3366 (N_3366,N_2660,N_2049);
and U3367 (N_3367,N_1511,N_2810);
nor U3368 (N_3368,N_2352,N_2287);
or U3369 (N_3369,N_2111,N_2113);
nand U3370 (N_3370,N_2840,N_2892);
xor U3371 (N_3371,N_2534,N_2831);
and U3372 (N_3372,N_2220,N_2723);
and U3373 (N_3373,N_2209,N_2379);
nor U3374 (N_3374,N_2859,N_2418);
and U3375 (N_3375,N_1689,N_2714);
and U3376 (N_3376,N_2001,N_2306);
nor U3377 (N_3377,N_2962,N_2826);
nor U3378 (N_3378,N_2820,N_2774);
nor U3379 (N_3379,N_1815,N_2403);
nor U3380 (N_3380,N_1630,N_1887);
xnor U3381 (N_3381,N_2449,N_2678);
nor U3382 (N_3382,N_2253,N_1579);
nand U3383 (N_3383,N_1674,N_2654);
nor U3384 (N_3384,N_2087,N_1803);
or U3385 (N_3385,N_2532,N_2211);
and U3386 (N_3386,N_2440,N_2647);
and U3387 (N_3387,N_2037,N_2639);
and U3388 (N_3388,N_1544,N_2542);
nand U3389 (N_3389,N_1713,N_2817);
and U3390 (N_3390,N_1885,N_2547);
xor U3391 (N_3391,N_1526,N_1652);
and U3392 (N_3392,N_1597,N_1903);
and U3393 (N_3393,N_1766,N_2889);
and U3394 (N_3394,N_1522,N_2568);
and U3395 (N_3395,N_2185,N_2215);
nand U3396 (N_3396,N_2652,N_1586);
or U3397 (N_3397,N_2706,N_2519);
nor U3398 (N_3398,N_2901,N_1549);
nor U3399 (N_3399,N_2390,N_1846);
nor U3400 (N_3400,N_2510,N_1835);
nand U3401 (N_3401,N_1725,N_2071);
or U3402 (N_3402,N_2758,N_2505);
or U3403 (N_3403,N_2961,N_2106);
nor U3404 (N_3404,N_2573,N_1945);
nor U3405 (N_3405,N_2682,N_2880);
and U3406 (N_3406,N_1940,N_2819);
nand U3407 (N_3407,N_1717,N_1823);
nand U3408 (N_3408,N_2422,N_2457);
xnor U3409 (N_3409,N_1918,N_2415);
nand U3410 (N_3410,N_1922,N_2788);
xnor U3411 (N_3411,N_2794,N_2496);
nand U3412 (N_3412,N_1670,N_1901);
and U3413 (N_3413,N_1858,N_2420);
nor U3414 (N_3414,N_2230,N_2245);
nand U3415 (N_3415,N_2050,N_2696);
xnor U3416 (N_3416,N_2233,N_2445);
and U3417 (N_3417,N_2154,N_1916);
xnor U3418 (N_3418,N_2596,N_2314);
or U3419 (N_3419,N_1728,N_1772);
or U3420 (N_3420,N_2550,N_1986);
nor U3421 (N_3421,N_2075,N_1878);
or U3422 (N_3422,N_2217,N_2526);
nor U3423 (N_3423,N_1950,N_2335);
xnor U3424 (N_3424,N_1730,N_1827);
and U3425 (N_3425,N_2844,N_2821);
nor U3426 (N_3426,N_2638,N_2280);
and U3427 (N_3427,N_2900,N_1831);
and U3428 (N_3428,N_1838,N_2636);
xor U3429 (N_3429,N_2967,N_1533);
and U3430 (N_3430,N_2978,N_2137);
xor U3431 (N_3431,N_2635,N_1735);
and U3432 (N_3432,N_1724,N_1641);
nand U3433 (N_3433,N_1547,N_1917);
nand U3434 (N_3434,N_1722,N_1995);
nor U3435 (N_3435,N_2783,N_2579);
nor U3436 (N_3436,N_1542,N_2134);
nand U3437 (N_3437,N_1631,N_2182);
nor U3438 (N_3438,N_2746,N_2734);
or U3439 (N_3439,N_2222,N_2489);
nor U3440 (N_3440,N_2689,N_1677);
nor U3441 (N_3441,N_2347,N_2730);
nand U3442 (N_3442,N_2592,N_1617);
or U3443 (N_3443,N_2634,N_2033);
xor U3444 (N_3444,N_2462,N_2148);
nor U3445 (N_3445,N_2288,N_2912);
and U3446 (N_3446,N_1744,N_2426);
and U3447 (N_3447,N_2408,N_2985);
nand U3448 (N_3448,N_2516,N_2021);
nor U3449 (N_3449,N_2943,N_2946);
and U3450 (N_3450,N_1841,N_1998);
and U3451 (N_3451,N_1629,N_1523);
or U3452 (N_3452,N_2240,N_2264);
or U3453 (N_3453,N_1763,N_2190);
nand U3454 (N_3454,N_2316,N_2796);
nand U3455 (N_3455,N_1816,N_2195);
nand U3456 (N_3456,N_2080,N_2594);
nor U3457 (N_3457,N_2374,N_1714);
xor U3458 (N_3458,N_2475,N_2598);
nand U3459 (N_3459,N_2675,N_2214);
and U3460 (N_3460,N_2935,N_2112);
or U3461 (N_3461,N_2565,N_1742);
or U3462 (N_3462,N_1873,N_2202);
xnor U3463 (N_3463,N_1656,N_2953);
nor U3464 (N_3464,N_2806,N_1612);
nor U3465 (N_3465,N_2808,N_1595);
or U3466 (N_3466,N_1541,N_2651);
nand U3467 (N_3467,N_1660,N_2104);
nor U3468 (N_3468,N_2950,N_2417);
or U3469 (N_3469,N_2203,N_2906);
and U3470 (N_3470,N_2231,N_2143);
and U3471 (N_3471,N_2715,N_2132);
nand U3472 (N_3472,N_2575,N_2861);
and U3473 (N_3473,N_1820,N_2101);
xor U3474 (N_3474,N_1582,N_2434);
nor U3475 (N_3475,N_2688,N_2919);
or U3476 (N_3476,N_1667,N_2538);
or U3477 (N_3477,N_2004,N_1767);
nand U3478 (N_3478,N_2484,N_2338);
and U3479 (N_3479,N_2899,N_1840);
nor U3480 (N_3480,N_2402,N_1834);
nand U3481 (N_3481,N_2964,N_2976);
nand U3482 (N_3482,N_1552,N_1990);
nand U3483 (N_3483,N_1707,N_2712);
or U3484 (N_3484,N_2833,N_2428);
and U3485 (N_3485,N_2160,N_2269);
nor U3486 (N_3486,N_2072,N_1676);
nand U3487 (N_3487,N_1892,N_1871);
nand U3488 (N_3488,N_2822,N_2775);
xor U3489 (N_3489,N_2815,N_2855);
nor U3490 (N_3490,N_1826,N_2560);
or U3491 (N_3491,N_1980,N_1648);
and U3492 (N_3492,N_2828,N_2615);
nor U3493 (N_3493,N_2218,N_2709);
nand U3494 (N_3494,N_2109,N_2472);
or U3495 (N_3495,N_1759,N_2626);
or U3496 (N_3496,N_2480,N_1754);
xnor U3497 (N_3497,N_1739,N_2600);
nand U3498 (N_3498,N_1740,N_1741);
and U3499 (N_3499,N_2097,N_2677);
and U3500 (N_3500,N_1726,N_1856);
nor U3501 (N_3501,N_2559,N_2525);
nand U3502 (N_3502,N_1568,N_1828);
xnor U3503 (N_3503,N_2206,N_1946);
or U3504 (N_3504,N_1964,N_2344);
nor U3505 (N_3505,N_2166,N_2755);
or U3506 (N_3506,N_2495,N_1868);
nor U3507 (N_3507,N_1534,N_2674);
or U3508 (N_3508,N_2557,N_2523);
and U3509 (N_3509,N_2910,N_2081);
or U3510 (N_3510,N_1570,N_2865);
and U3511 (N_3511,N_2934,N_2125);
or U3512 (N_3512,N_1948,N_2988);
nor U3513 (N_3513,N_2877,N_2732);
nor U3514 (N_3514,N_2135,N_2759);
nand U3515 (N_3515,N_1733,N_1890);
and U3516 (N_3516,N_1598,N_1673);
xnor U3517 (N_3517,N_1657,N_2350);
and U3518 (N_3518,N_2763,N_2047);
nor U3519 (N_3519,N_2213,N_2710);
or U3520 (N_3520,N_2152,N_2644);
and U3521 (N_3521,N_2544,N_2011);
and U3522 (N_3522,N_2376,N_1678);
or U3523 (N_3523,N_1647,N_1503);
nor U3524 (N_3524,N_2951,N_2939);
or U3525 (N_3525,N_1557,N_1804);
nand U3526 (N_3526,N_2163,N_1849);
and U3527 (N_3527,N_2780,N_2498);
or U3528 (N_3528,N_2186,N_2882);
nand U3529 (N_3529,N_2945,N_2926);
nand U3530 (N_3530,N_2172,N_2204);
nor U3531 (N_3531,N_2982,N_2928);
or U3532 (N_3532,N_2303,N_2649);
nand U3533 (N_3533,N_2039,N_2895);
nor U3534 (N_3534,N_2614,N_2541);
and U3535 (N_3535,N_1824,N_2225);
and U3536 (N_3536,N_1509,N_1971);
and U3537 (N_3537,N_2212,N_2019);
nor U3538 (N_3538,N_2832,N_2108);
or U3539 (N_3539,N_2003,N_1668);
and U3540 (N_3540,N_1809,N_1538);
and U3541 (N_3541,N_1750,N_2086);
nand U3542 (N_3542,N_2818,N_2129);
or U3543 (N_3543,N_2124,N_1915);
nand U3544 (N_3544,N_1539,N_1637);
or U3545 (N_3545,N_1596,N_1902);
and U3546 (N_3546,N_1760,N_2250);
and U3547 (N_3547,N_1859,N_1941);
xnor U3548 (N_3548,N_1751,N_2364);
nor U3549 (N_3549,N_2307,N_2664);
xnor U3550 (N_3550,N_1966,N_2770);
nor U3551 (N_3551,N_2656,N_1685);
nor U3552 (N_3552,N_1512,N_1850);
and U3553 (N_3553,N_2319,N_1543);
or U3554 (N_3554,N_2885,N_1952);
nand U3555 (N_3555,N_1615,N_1912);
or U3556 (N_3556,N_2549,N_1565);
and U3557 (N_3557,N_1692,N_2002);
xor U3558 (N_3558,N_1793,N_2224);
and U3559 (N_3559,N_2469,N_1594);
nor U3560 (N_3560,N_2756,N_2289);
nand U3561 (N_3561,N_1962,N_2067);
nor U3562 (N_3562,N_2354,N_1954);
nor U3563 (N_3563,N_2539,N_1947);
nor U3564 (N_3564,N_2692,N_2883);
nand U3565 (N_3565,N_2467,N_2582);
and U3566 (N_3566,N_2164,N_2760);
and U3567 (N_3567,N_2191,N_2285);
nand U3568 (N_3568,N_2802,N_2372);
and U3569 (N_3569,N_2007,N_1898);
xnor U3570 (N_3570,N_2824,N_1698);
nand U3571 (N_3571,N_2016,N_2631);
nor U3572 (N_3572,N_1619,N_2365);
and U3573 (N_3573,N_1999,N_2062);
nor U3574 (N_3574,N_2053,N_2916);
xnor U3575 (N_3575,N_2361,N_1556);
and U3576 (N_3576,N_2891,N_2324);
nor U3577 (N_3577,N_2601,N_1680);
xnor U3578 (N_3578,N_2841,N_1664);
xor U3579 (N_3579,N_2136,N_2669);
nand U3580 (N_3580,N_2321,N_2151);
nand U3581 (N_3581,N_2751,N_2784);
nor U3582 (N_3582,N_2282,N_1821);
and U3583 (N_3583,N_2357,N_1551);
nor U3584 (N_3584,N_2485,N_2246);
or U3585 (N_3585,N_1580,N_1797);
nor U3586 (N_3586,N_1644,N_1646);
or U3587 (N_3587,N_2869,N_1829);
xnor U3588 (N_3588,N_1640,N_1812);
nor U3589 (N_3589,N_1978,N_2681);
or U3590 (N_3590,N_2093,N_2263);
or U3591 (N_3591,N_1690,N_1955);
xnor U3592 (N_3592,N_2433,N_1723);
nand U3593 (N_3593,N_2477,N_2502);
and U3594 (N_3594,N_1727,N_2405);
and U3595 (N_3595,N_1839,N_2055);
or U3596 (N_3596,N_1504,N_2394);
xor U3597 (N_3597,N_2727,N_1524);
and U3598 (N_3598,N_2672,N_1602);
nand U3599 (N_3599,N_2258,N_2721);
or U3600 (N_3600,N_1627,N_2720);
or U3601 (N_3601,N_1865,N_2973);
xnor U3602 (N_3602,N_2884,N_2491);
nand U3603 (N_3603,N_1559,N_2989);
nand U3604 (N_3604,N_2369,N_2566);
nor U3605 (N_3605,N_2035,N_2993);
or U3606 (N_3606,N_2268,N_1956);
or U3607 (N_3607,N_2396,N_2120);
nor U3608 (N_3608,N_2700,N_2326);
nand U3609 (N_3609,N_2052,N_2779);
nor U3610 (N_3610,N_2699,N_2140);
or U3611 (N_3611,N_2858,N_2479);
or U3612 (N_3612,N_2972,N_2056);
nand U3613 (N_3613,N_1965,N_2391);
nor U3614 (N_3614,N_1569,N_2522);
and U3615 (N_3615,N_2536,N_2736);
nand U3616 (N_3616,N_2595,N_2105);
nor U3617 (N_3617,N_1899,N_1572);
nor U3618 (N_3618,N_1611,N_1911);
and U3619 (N_3619,N_2424,N_2175);
nand U3620 (N_3620,N_1794,N_2680);
or U3621 (N_3621,N_2556,N_2769);
or U3622 (N_3622,N_2032,N_1567);
or U3623 (N_3623,N_2842,N_2251);
and U3624 (N_3624,N_1530,N_2874);
nand U3625 (N_3625,N_2624,N_2645);
nor U3626 (N_3626,N_2937,N_1506);
and U3627 (N_3627,N_2378,N_1655);
and U3628 (N_3628,N_1607,N_1537);
nand U3629 (N_3629,N_1671,N_1632);
or U3630 (N_3630,N_1985,N_2589);
nor U3631 (N_3631,N_2036,N_2098);
and U3632 (N_3632,N_2359,N_2070);
nor U3633 (N_3633,N_2216,N_2058);
or U3634 (N_3634,N_2501,N_2646);
and U3635 (N_3635,N_2305,N_2228);
nand U3636 (N_3636,N_1813,N_1938);
or U3637 (N_3637,N_2192,N_2199);
or U3638 (N_3638,N_1989,N_2657);
nor U3639 (N_3639,N_2648,N_1622);
nand U3640 (N_3640,N_2835,N_2611);
and U3641 (N_3641,N_1608,N_2370);
xor U3642 (N_3642,N_2456,N_2613);
xor U3643 (N_3643,N_1973,N_1609);
xnor U3644 (N_3644,N_2766,N_2909);
and U3645 (N_3645,N_1994,N_2662);
xnor U3646 (N_3646,N_2530,N_2200);
and U3647 (N_3647,N_2368,N_2508);
nor U3648 (N_3648,N_1935,N_1686);
or U3649 (N_3649,N_2676,N_2809);
or U3650 (N_3650,N_1930,N_1502);
nand U3651 (N_3651,N_1836,N_2460);
nor U3652 (N_3652,N_1825,N_1862);
or U3653 (N_3653,N_1923,N_2868);
nand U3654 (N_3654,N_2940,N_2078);
nand U3655 (N_3655,N_1535,N_2061);
nand U3656 (N_3656,N_2126,N_2119);
or U3657 (N_3657,N_2846,N_2063);
or U3658 (N_3658,N_1877,N_2933);
xnor U3659 (N_3659,N_1753,N_2807);
nor U3660 (N_3660,N_1616,N_2461);
or U3661 (N_3661,N_2343,N_2905);
and U3662 (N_3662,N_2464,N_1920);
and U3663 (N_3663,N_2167,N_1785);
nand U3664 (N_3664,N_1675,N_2875);
or U3665 (N_3665,N_2117,N_2944);
nor U3666 (N_3666,N_2701,N_2416);
nand U3667 (N_3667,N_1842,N_2637);
nand U3668 (N_3668,N_1694,N_2298);
nand U3669 (N_3669,N_2569,N_2492);
nor U3670 (N_3670,N_2292,N_2122);
nor U3671 (N_3671,N_1798,N_2567);
xnor U3672 (N_3672,N_1907,N_2051);
nor U3673 (N_3673,N_2173,N_2130);
or U3674 (N_3674,N_2141,N_2382);
nor U3675 (N_3675,N_2797,N_2518);
or U3676 (N_3676,N_2507,N_1747);
and U3677 (N_3677,N_1969,N_2650);
or U3678 (N_3678,N_1745,N_2698);
and U3679 (N_3679,N_1591,N_2580);
nor U3680 (N_3680,N_1951,N_2504);
nor U3681 (N_3681,N_2340,N_2603);
and U3682 (N_3682,N_2679,N_1505);
or U3683 (N_3683,N_2145,N_2144);
nor U3684 (N_3684,N_2413,N_2468);
nand U3685 (N_3685,N_1532,N_1510);
nand U3686 (N_3686,N_2247,N_2778);
nor U3687 (N_3687,N_2014,N_2102);
xor U3688 (N_3688,N_2400,N_1529);
nand U3689 (N_3689,N_2667,N_2162);
nand U3690 (N_3690,N_2515,N_2170);
nor U3691 (N_3691,N_2482,N_1757);
and U3692 (N_3692,N_2969,N_1515);
nor U3693 (N_3693,N_1880,N_2283);
and U3694 (N_3694,N_2838,N_1811);
or U3695 (N_3695,N_1970,N_2583);
nand U3696 (N_3696,N_1848,N_2999);
and U3697 (N_3697,N_2930,N_2984);
and U3698 (N_3698,N_2229,N_2156);
nor U3699 (N_3699,N_1665,N_2196);
nand U3700 (N_3700,N_2177,N_2913);
or U3701 (N_3701,N_2267,N_1801);
nor U3702 (N_3702,N_1519,N_2693);
or U3703 (N_3703,N_1704,N_1587);
nor U3704 (N_3704,N_2799,N_1571);
nor U3705 (N_3705,N_2150,N_2798);
nor U3706 (N_3706,N_1527,N_2668);
or U3707 (N_3707,N_2236,N_2923);
or U3708 (N_3708,N_2971,N_2174);
nor U3709 (N_3709,N_2429,N_2453);
nor U3710 (N_3710,N_2026,N_2038);
nand U3711 (N_3711,N_2054,N_1976);
and U3712 (N_3712,N_1806,N_2234);
nor U3713 (N_3713,N_1658,N_2249);
nor U3714 (N_3714,N_2791,N_2028);
and U3715 (N_3715,N_1855,N_2410);
nand U3716 (N_3716,N_2708,N_2128);
nor U3717 (N_3717,N_1507,N_2870);
nand U3718 (N_3718,N_2713,N_2742);
nor U3719 (N_3719,N_2860,N_2265);
nand U3720 (N_3720,N_2653,N_2009);
or U3721 (N_3721,N_2625,N_2702);
and U3722 (N_3722,N_2524,N_2661);
xor U3723 (N_3723,N_1588,N_1695);
xnor U3724 (N_3724,N_2845,N_2252);
nand U3725 (N_3725,N_2641,N_1712);
nor U3726 (N_3726,N_2862,N_1621);
nor U3727 (N_3727,N_2227,N_1830);
or U3728 (N_3728,N_2704,N_2103);
and U3729 (N_3729,N_2629,N_1634);
nand U3730 (N_3730,N_1550,N_1553);
and U3731 (N_3731,N_2317,N_2590);
nand U3732 (N_3732,N_1770,N_2257);
or U3733 (N_3733,N_2270,N_2623);
or U3734 (N_3734,N_1593,N_1776);
or U3735 (N_3735,N_2691,N_1908);
nand U3736 (N_3736,N_2158,N_2551);
and U3737 (N_3737,N_2367,N_2981);
and U3738 (N_3738,N_1833,N_1517);
nand U3739 (N_3739,N_2235,N_2792);
and U3740 (N_3740,N_2514,N_1618);
and U3741 (N_3741,N_1614,N_1810);
or U3742 (N_3742,N_2621,N_1721);
and U3743 (N_3743,N_1663,N_2617);
and U3744 (N_3744,N_2432,N_2599);
and U3745 (N_3745,N_2308,N_2193);
nor U3746 (N_3746,N_2745,N_1605);
nor U3747 (N_3747,N_2437,N_2848);
and U3748 (N_3748,N_2008,N_2537);
nor U3749 (N_3749,N_2430,N_1870);
nand U3750 (N_3750,N_2918,N_1703);
nor U3751 (N_3751,N_2573,N_2741);
nand U3752 (N_3752,N_2190,N_2279);
xnor U3753 (N_3753,N_2506,N_2382);
nand U3754 (N_3754,N_1877,N_1689);
xor U3755 (N_3755,N_2347,N_2001);
or U3756 (N_3756,N_2415,N_2606);
nor U3757 (N_3757,N_2270,N_1537);
or U3758 (N_3758,N_1524,N_2463);
xor U3759 (N_3759,N_2340,N_1524);
or U3760 (N_3760,N_2517,N_1999);
nand U3761 (N_3761,N_2271,N_2317);
nor U3762 (N_3762,N_2886,N_2946);
nor U3763 (N_3763,N_2516,N_2175);
and U3764 (N_3764,N_1672,N_1660);
nand U3765 (N_3765,N_1694,N_2045);
nand U3766 (N_3766,N_2033,N_2149);
nand U3767 (N_3767,N_2224,N_2177);
nand U3768 (N_3768,N_1829,N_2972);
and U3769 (N_3769,N_1881,N_2402);
nand U3770 (N_3770,N_2655,N_2241);
xnor U3771 (N_3771,N_2171,N_2221);
and U3772 (N_3772,N_2810,N_1792);
nand U3773 (N_3773,N_2952,N_2700);
nor U3774 (N_3774,N_2800,N_1850);
nor U3775 (N_3775,N_1773,N_1720);
and U3776 (N_3776,N_1927,N_2265);
xor U3777 (N_3777,N_2112,N_2873);
nand U3778 (N_3778,N_1575,N_2581);
and U3779 (N_3779,N_2109,N_1936);
nand U3780 (N_3780,N_2670,N_1969);
nor U3781 (N_3781,N_1646,N_1539);
nor U3782 (N_3782,N_1824,N_2174);
nand U3783 (N_3783,N_2188,N_2216);
nand U3784 (N_3784,N_2828,N_2576);
nand U3785 (N_3785,N_1832,N_2572);
or U3786 (N_3786,N_1928,N_1976);
nor U3787 (N_3787,N_2263,N_1520);
nand U3788 (N_3788,N_2912,N_2299);
nand U3789 (N_3789,N_1634,N_2035);
and U3790 (N_3790,N_2838,N_1823);
or U3791 (N_3791,N_2438,N_1802);
nand U3792 (N_3792,N_2422,N_1646);
nand U3793 (N_3793,N_2231,N_1712);
nand U3794 (N_3794,N_1846,N_1978);
or U3795 (N_3795,N_1800,N_1582);
nor U3796 (N_3796,N_1957,N_1764);
or U3797 (N_3797,N_1875,N_2314);
nor U3798 (N_3798,N_1871,N_2927);
nor U3799 (N_3799,N_1886,N_2716);
nor U3800 (N_3800,N_2664,N_2365);
nor U3801 (N_3801,N_2774,N_2570);
or U3802 (N_3802,N_2527,N_2679);
xnor U3803 (N_3803,N_2046,N_2513);
nor U3804 (N_3804,N_2267,N_2377);
nor U3805 (N_3805,N_1730,N_2695);
nor U3806 (N_3806,N_1731,N_2237);
nor U3807 (N_3807,N_2167,N_2531);
and U3808 (N_3808,N_1735,N_2952);
and U3809 (N_3809,N_2090,N_2411);
nor U3810 (N_3810,N_1616,N_2453);
and U3811 (N_3811,N_2200,N_2784);
nand U3812 (N_3812,N_2873,N_2468);
nor U3813 (N_3813,N_1966,N_1767);
nor U3814 (N_3814,N_2707,N_2064);
and U3815 (N_3815,N_1800,N_2295);
xnor U3816 (N_3816,N_1759,N_1746);
nor U3817 (N_3817,N_2552,N_2846);
or U3818 (N_3818,N_1784,N_1558);
nand U3819 (N_3819,N_1746,N_2125);
and U3820 (N_3820,N_2296,N_2784);
and U3821 (N_3821,N_1975,N_2313);
or U3822 (N_3822,N_2987,N_2485);
xor U3823 (N_3823,N_1614,N_2050);
xor U3824 (N_3824,N_2460,N_2363);
nand U3825 (N_3825,N_2137,N_2106);
nand U3826 (N_3826,N_2323,N_1723);
and U3827 (N_3827,N_1878,N_2848);
nor U3828 (N_3828,N_1939,N_2036);
nor U3829 (N_3829,N_2745,N_2312);
nand U3830 (N_3830,N_1703,N_2084);
nand U3831 (N_3831,N_2104,N_2529);
nor U3832 (N_3832,N_1865,N_2209);
and U3833 (N_3833,N_2068,N_2967);
and U3834 (N_3834,N_2097,N_2584);
nor U3835 (N_3835,N_2259,N_2421);
or U3836 (N_3836,N_2013,N_1558);
xnor U3837 (N_3837,N_1858,N_2855);
nor U3838 (N_3838,N_2886,N_2263);
and U3839 (N_3839,N_1699,N_2574);
xor U3840 (N_3840,N_2309,N_2408);
and U3841 (N_3841,N_2449,N_1690);
nor U3842 (N_3842,N_2451,N_2229);
nand U3843 (N_3843,N_2445,N_1589);
or U3844 (N_3844,N_2443,N_1672);
nand U3845 (N_3845,N_1852,N_2656);
nand U3846 (N_3846,N_2652,N_1873);
nor U3847 (N_3847,N_2116,N_2470);
and U3848 (N_3848,N_2869,N_2090);
nand U3849 (N_3849,N_2998,N_1608);
or U3850 (N_3850,N_1871,N_2470);
or U3851 (N_3851,N_2135,N_2348);
nor U3852 (N_3852,N_2255,N_2643);
and U3853 (N_3853,N_2453,N_2430);
or U3854 (N_3854,N_2263,N_1952);
or U3855 (N_3855,N_1724,N_2966);
and U3856 (N_3856,N_2388,N_2663);
nand U3857 (N_3857,N_2579,N_1661);
or U3858 (N_3858,N_2645,N_1598);
or U3859 (N_3859,N_1570,N_1560);
or U3860 (N_3860,N_2846,N_2966);
and U3861 (N_3861,N_2611,N_2957);
nor U3862 (N_3862,N_2900,N_1799);
nor U3863 (N_3863,N_1877,N_1883);
and U3864 (N_3864,N_1957,N_2979);
and U3865 (N_3865,N_2630,N_2463);
nand U3866 (N_3866,N_1725,N_2134);
and U3867 (N_3867,N_2922,N_1512);
or U3868 (N_3868,N_2266,N_1891);
nor U3869 (N_3869,N_1966,N_2403);
nand U3870 (N_3870,N_2516,N_2433);
and U3871 (N_3871,N_2235,N_1794);
and U3872 (N_3872,N_1745,N_1666);
nor U3873 (N_3873,N_2897,N_2581);
or U3874 (N_3874,N_2117,N_2198);
nor U3875 (N_3875,N_2733,N_2540);
nand U3876 (N_3876,N_2608,N_1597);
xor U3877 (N_3877,N_2585,N_1961);
nand U3878 (N_3878,N_2177,N_2985);
or U3879 (N_3879,N_2065,N_2380);
xnor U3880 (N_3880,N_1958,N_2646);
xnor U3881 (N_3881,N_1718,N_2299);
nand U3882 (N_3882,N_1637,N_1960);
and U3883 (N_3883,N_2919,N_2193);
nand U3884 (N_3884,N_2144,N_2389);
nand U3885 (N_3885,N_2423,N_2808);
xnor U3886 (N_3886,N_2682,N_2265);
xnor U3887 (N_3887,N_2838,N_2686);
and U3888 (N_3888,N_1919,N_1855);
and U3889 (N_3889,N_1628,N_1990);
nor U3890 (N_3890,N_1597,N_2504);
or U3891 (N_3891,N_1545,N_2681);
or U3892 (N_3892,N_1507,N_2241);
and U3893 (N_3893,N_1890,N_2897);
and U3894 (N_3894,N_2139,N_1863);
and U3895 (N_3895,N_2667,N_2748);
or U3896 (N_3896,N_2677,N_2727);
or U3897 (N_3897,N_2016,N_1546);
nand U3898 (N_3898,N_2677,N_1894);
nor U3899 (N_3899,N_1809,N_2193);
or U3900 (N_3900,N_2279,N_2326);
or U3901 (N_3901,N_1554,N_2514);
or U3902 (N_3902,N_2621,N_2592);
and U3903 (N_3903,N_2107,N_1514);
nor U3904 (N_3904,N_1509,N_2809);
xnor U3905 (N_3905,N_1610,N_1622);
xnor U3906 (N_3906,N_2700,N_2402);
nor U3907 (N_3907,N_1716,N_1736);
nand U3908 (N_3908,N_2964,N_2403);
nand U3909 (N_3909,N_2075,N_1920);
xor U3910 (N_3910,N_2988,N_1911);
or U3911 (N_3911,N_2742,N_1833);
nand U3912 (N_3912,N_2674,N_2560);
or U3913 (N_3913,N_2798,N_1906);
or U3914 (N_3914,N_2756,N_2878);
nor U3915 (N_3915,N_1647,N_1740);
and U3916 (N_3916,N_1782,N_2240);
or U3917 (N_3917,N_2616,N_1710);
nor U3918 (N_3918,N_2801,N_1826);
xor U3919 (N_3919,N_1614,N_2015);
nand U3920 (N_3920,N_2149,N_2851);
or U3921 (N_3921,N_1690,N_1686);
or U3922 (N_3922,N_2087,N_2107);
or U3923 (N_3923,N_1820,N_1865);
or U3924 (N_3924,N_1538,N_2325);
nor U3925 (N_3925,N_2869,N_2542);
nand U3926 (N_3926,N_2598,N_1645);
xor U3927 (N_3927,N_1750,N_2095);
and U3928 (N_3928,N_2924,N_2221);
nand U3929 (N_3929,N_2187,N_2947);
nor U3930 (N_3930,N_1875,N_2258);
and U3931 (N_3931,N_1507,N_1624);
or U3932 (N_3932,N_2132,N_1607);
or U3933 (N_3933,N_2001,N_2040);
or U3934 (N_3934,N_2513,N_2140);
xor U3935 (N_3935,N_2419,N_1602);
nand U3936 (N_3936,N_1583,N_2416);
nor U3937 (N_3937,N_1803,N_1638);
nor U3938 (N_3938,N_2566,N_2172);
nand U3939 (N_3939,N_1601,N_2944);
nand U3940 (N_3940,N_2667,N_1952);
nand U3941 (N_3941,N_1578,N_1579);
nand U3942 (N_3942,N_1716,N_2334);
nor U3943 (N_3943,N_1526,N_1809);
and U3944 (N_3944,N_2740,N_2644);
xor U3945 (N_3945,N_1764,N_2370);
and U3946 (N_3946,N_2183,N_1970);
and U3947 (N_3947,N_2174,N_1914);
or U3948 (N_3948,N_2915,N_2805);
nor U3949 (N_3949,N_1794,N_1502);
or U3950 (N_3950,N_2540,N_1758);
nor U3951 (N_3951,N_1888,N_2761);
nand U3952 (N_3952,N_2833,N_2571);
nor U3953 (N_3953,N_2516,N_1980);
nor U3954 (N_3954,N_2394,N_2431);
nor U3955 (N_3955,N_2676,N_2366);
and U3956 (N_3956,N_2577,N_2324);
nor U3957 (N_3957,N_2272,N_2341);
or U3958 (N_3958,N_2601,N_2551);
and U3959 (N_3959,N_2613,N_2234);
or U3960 (N_3960,N_2917,N_1518);
and U3961 (N_3961,N_1885,N_1820);
nand U3962 (N_3962,N_2154,N_2874);
nor U3963 (N_3963,N_2805,N_2285);
and U3964 (N_3964,N_2806,N_2718);
or U3965 (N_3965,N_2350,N_1980);
or U3966 (N_3966,N_2919,N_1775);
nor U3967 (N_3967,N_1855,N_1531);
nor U3968 (N_3968,N_2447,N_2512);
nand U3969 (N_3969,N_1506,N_2110);
nand U3970 (N_3970,N_2169,N_1795);
or U3971 (N_3971,N_2212,N_2959);
and U3972 (N_3972,N_1715,N_2914);
or U3973 (N_3973,N_1625,N_1626);
nand U3974 (N_3974,N_2932,N_2335);
nor U3975 (N_3975,N_1561,N_1782);
nand U3976 (N_3976,N_1520,N_1727);
nand U3977 (N_3977,N_1883,N_2771);
nand U3978 (N_3978,N_2787,N_2069);
and U3979 (N_3979,N_2275,N_1505);
or U3980 (N_3980,N_2654,N_2554);
nand U3981 (N_3981,N_1742,N_2186);
xnor U3982 (N_3982,N_2849,N_2100);
nor U3983 (N_3983,N_1814,N_2206);
xnor U3984 (N_3984,N_1873,N_2790);
xnor U3985 (N_3985,N_1908,N_2611);
and U3986 (N_3986,N_2475,N_1656);
nand U3987 (N_3987,N_2332,N_2619);
and U3988 (N_3988,N_1861,N_2623);
nand U3989 (N_3989,N_1512,N_1542);
nor U3990 (N_3990,N_2367,N_2190);
or U3991 (N_3991,N_1864,N_2751);
and U3992 (N_3992,N_2123,N_2529);
nand U3993 (N_3993,N_1795,N_2865);
xnor U3994 (N_3994,N_2868,N_2224);
or U3995 (N_3995,N_1989,N_2334);
and U3996 (N_3996,N_1940,N_2035);
or U3997 (N_3997,N_1994,N_1587);
or U3998 (N_3998,N_2501,N_2250);
nor U3999 (N_3999,N_1551,N_2735);
nor U4000 (N_4000,N_2175,N_2758);
nor U4001 (N_4001,N_1546,N_1717);
and U4002 (N_4002,N_1678,N_2989);
nand U4003 (N_4003,N_2007,N_2369);
xor U4004 (N_4004,N_1542,N_2780);
and U4005 (N_4005,N_1882,N_1881);
and U4006 (N_4006,N_1837,N_2714);
xnor U4007 (N_4007,N_2347,N_2711);
nor U4008 (N_4008,N_2832,N_1982);
xor U4009 (N_4009,N_2576,N_2280);
nor U4010 (N_4010,N_2602,N_2806);
or U4011 (N_4011,N_1786,N_2135);
or U4012 (N_4012,N_2536,N_1792);
nor U4013 (N_4013,N_1874,N_2783);
nor U4014 (N_4014,N_2608,N_2338);
or U4015 (N_4015,N_2928,N_2783);
or U4016 (N_4016,N_1601,N_2156);
nand U4017 (N_4017,N_2594,N_1750);
or U4018 (N_4018,N_1739,N_1625);
xor U4019 (N_4019,N_2753,N_2869);
nor U4020 (N_4020,N_2766,N_2341);
or U4021 (N_4021,N_2956,N_2770);
nand U4022 (N_4022,N_1510,N_1890);
or U4023 (N_4023,N_2198,N_2694);
nand U4024 (N_4024,N_2358,N_2402);
or U4025 (N_4025,N_2511,N_2497);
nand U4026 (N_4026,N_1899,N_2498);
or U4027 (N_4027,N_2330,N_2245);
or U4028 (N_4028,N_1533,N_2427);
nand U4029 (N_4029,N_2320,N_2539);
nand U4030 (N_4030,N_2395,N_2492);
nor U4031 (N_4031,N_1910,N_2937);
nor U4032 (N_4032,N_2448,N_2720);
nor U4033 (N_4033,N_1934,N_1958);
or U4034 (N_4034,N_2348,N_2701);
or U4035 (N_4035,N_1897,N_2329);
or U4036 (N_4036,N_2469,N_2804);
and U4037 (N_4037,N_2292,N_2343);
or U4038 (N_4038,N_1762,N_2812);
nand U4039 (N_4039,N_1961,N_2033);
nand U4040 (N_4040,N_2959,N_1714);
nand U4041 (N_4041,N_2598,N_2078);
nor U4042 (N_4042,N_2682,N_2551);
or U4043 (N_4043,N_2342,N_2145);
or U4044 (N_4044,N_2744,N_1926);
nand U4045 (N_4045,N_1881,N_2704);
xnor U4046 (N_4046,N_1716,N_2321);
or U4047 (N_4047,N_2910,N_2327);
or U4048 (N_4048,N_2635,N_2301);
and U4049 (N_4049,N_2964,N_2624);
nand U4050 (N_4050,N_1505,N_1724);
nand U4051 (N_4051,N_2736,N_2374);
nand U4052 (N_4052,N_2210,N_1706);
nand U4053 (N_4053,N_2171,N_2520);
xnor U4054 (N_4054,N_2392,N_2261);
nand U4055 (N_4055,N_2331,N_2186);
or U4056 (N_4056,N_2599,N_2122);
and U4057 (N_4057,N_1726,N_2539);
and U4058 (N_4058,N_2634,N_1723);
and U4059 (N_4059,N_2216,N_2804);
nor U4060 (N_4060,N_1767,N_2451);
and U4061 (N_4061,N_2694,N_2789);
or U4062 (N_4062,N_2765,N_2017);
nand U4063 (N_4063,N_1790,N_2824);
nor U4064 (N_4064,N_2306,N_1940);
nor U4065 (N_4065,N_2487,N_1919);
nand U4066 (N_4066,N_2064,N_1665);
nand U4067 (N_4067,N_2548,N_1648);
nor U4068 (N_4068,N_1703,N_2755);
and U4069 (N_4069,N_1754,N_2848);
and U4070 (N_4070,N_2331,N_1541);
nand U4071 (N_4071,N_2254,N_2545);
nor U4072 (N_4072,N_1716,N_2945);
and U4073 (N_4073,N_2990,N_1855);
xor U4074 (N_4074,N_2004,N_2354);
or U4075 (N_4075,N_2260,N_1786);
and U4076 (N_4076,N_2293,N_2928);
nand U4077 (N_4077,N_2020,N_2163);
nand U4078 (N_4078,N_2821,N_1600);
nor U4079 (N_4079,N_2900,N_1880);
and U4080 (N_4080,N_2808,N_2137);
and U4081 (N_4081,N_1969,N_2173);
and U4082 (N_4082,N_2767,N_1928);
and U4083 (N_4083,N_2856,N_2900);
nor U4084 (N_4084,N_2301,N_2947);
nor U4085 (N_4085,N_2755,N_2883);
or U4086 (N_4086,N_1855,N_2568);
nor U4087 (N_4087,N_1735,N_2954);
nor U4088 (N_4088,N_2731,N_1626);
nor U4089 (N_4089,N_1708,N_2777);
nor U4090 (N_4090,N_1787,N_2057);
and U4091 (N_4091,N_2153,N_1598);
xnor U4092 (N_4092,N_2907,N_2642);
nand U4093 (N_4093,N_2546,N_2265);
xor U4094 (N_4094,N_2964,N_1737);
or U4095 (N_4095,N_2645,N_1881);
nand U4096 (N_4096,N_2451,N_2256);
and U4097 (N_4097,N_2643,N_2390);
or U4098 (N_4098,N_2213,N_1907);
xor U4099 (N_4099,N_2128,N_2646);
or U4100 (N_4100,N_2337,N_1842);
and U4101 (N_4101,N_1699,N_2186);
and U4102 (N_4102,N_2063,N_2295);
nand U4103 (N_4103,N_2521,N_1588);
nand U4104 (N_4104,N_2075,N_2496);
nor U4105 (N_4105,N_1972,N_1622);
nand U4106 (N_4106,N_2188,N_2680);
and U4107 (N_4107,N_2827,N_1865);
nor U4108 (N_4108,N_2977,N_2388);
or U4109 (N_4109,N_2048,N_2200);
nor U4110 (N_4110,N_2725,N_1601);
nand U4111 (N_4111,N_2234,N_2354);
and U4112 (N_4112,N_2590,N_1710);
nor U4113 (N_4113,N_2037,N_2083);
nor U4114 (N_4114,N_2694,N_2041);
nand U4115 (N_4115,N_2149,N_2132);
and U4116 (N_4116,N_2043,N_2434);
nor U4117 (N_4117,N_2361,N_2418);
nand U4118 (N_4118,N_1582,N_2215);
nor U4119 (N_4119,N_2473,N_2238);
and U4120 (N_4120,N_2377,N_2120);
or U4121 (N_4121,N_1901,N_2422);
nor U4122 (N_4122,N_1829,N_2935);
or U4123 (N_4123,N_2309,N_2878);
nor U4124 (N_4124,N_2061,N_1581);
nor U4125 (N_4125,N_1628,N_2212);
nand U4126 (N_4126,N_2633,N_2481);
or U4127 (N_4127,N_1654,N_2451);
or U4128 (N_4128,N_1701,N_1829);
and U4129 (N_4129,N_2913,N_2594);
or U4130 (N_4130,N_1806,N_1501);
and U4131 (N_4131,N_2950,N_2221);
and U4132 (N_4132,N_2346,N_2630);
xnor U4133 (N_4133,N_1657,N_2167);
or U4134 (N_4134,N_2940,N_2938);
nor U4135 (N_4135,N_1985,N_2848);
or U4136 (N_4136,N_1775,N_1980);
nor U4137 (N_4137,N_2829,N_2164);
nand U4138 (N_4138,N_1562,N_2720);
nand U4139 (N_4139,N_2637,N_1927);
nand U4140 (N_4140,N_2411,N_2426);
nor U4141 (N_4141,N_2904,N_1510);
and U4142 (N_4142,N_2276,N_2178);
or U4143 (N_4143,N_2616,N_2931);
and U4144 (N_4144,N_2970,N_1793);
xor U4145 (N_4145,N_2022,N_2354);
nand U4146 (N_4146,N_1573,N_1953);
nand U4147 (N_4147,N_2605,N_2590);
and U4148 (N_4148,N_2025,N_2547);
nor U4149 (N_4149,N_2340,N_2991);
and U4150 (N_4150,N_1981,N_2788);
and U4151 (N_4151,N_2191,N_2634);
or U4152 (N_4152,N_2187,N_2339);
or U4153 (N_4153,N_2400,N_1740);
nand U4154 (N_4154,N_2962,N_2152);
nor U4155 (N_4155,N_2892,N_2059);
and U4156 (N_4156,N_1880,N_1739);
and U4157 (N_4157,N_1936,N_1927);
and U4158 (N_4158,N_2663,N_2059);
or U4159 (N_4159,N_1812,N_2120);
or U4160 (N_4160,N_2229,N_1754);
and U4161 (N_4161,N_2395,N_2586);
and U4162 (N_4162,N_1901,N_2425);
nor U4163 (N_4163,N_1732,N_2919);
nand U4164 (N_4164,N_2663,N_2056);
and U4165 (N_4165,N_1902,N_1969);
nor U4166 (N_4166,N_2887,N_1814);
and U4167 (N_4167,N_1827,N_2402);
or U4168 (N_4168,N_2024,N_2338);
and U4169 (N_4169,N_1741,N_2631);
and U4170 (N_4170,N_2277,N_2658);
nand U4171 (N_4171,N_2155,N_2989);
or U4172 (N_4172,N_1971,N_2102);
or U4173 (N_4173,N_1931,N_1792);
nor U4174 (N_4174,N_1778,N_2959);
or U4175 (N_4175,N_1933,N_2109);
and U4176 (N_4176,N_2767,N_1861);
nand U4177 (N_4177,N_1853,N_2420);
nor U4178 (N_4178,N_1664,N_2858);
nand U4179 (N_4179,N_2633,N_2863);
or U4180 (N_4180,N_2790,N_1959);
or U4181 (N_4181,N_2759,N_1700);
nor U4182 (N_4182,N_2216,N_2277);
and U4183 (N_4183,N_2065,N_2885);
and U4184 (N_4184,N_1818,N_2252);
and U4185 (N_4185,N_2134,N_1853);
nor U4186 (N_4186,N_2525,N_1942);
nand U4187 (N_4187,N_1635,N_2194);
and U4188 (N_4188,N_2327,N_2255);
or U4189 (N_4189,N_1730,N_2296);
nor U4190 (N_4190,N_2480,N_2472);
and U4191 (N_4191,N_2478,N_2871);
xnor U4192 (N_4192,N_2755,N_2164);
and U4193 (N_4193,N_2638,N_2045);
and U4194 (N_4194,N_1972,N_2653);
and U4195 (N_4195,N_2470,N_2986);
nand U4196 (N_4196,N_1532,N_2218);
nor U4197 (N_4197,N_2650,N_1984);
nor U4198 (N_4198,N_2453,N_2985);
nand U4199 (N_4199,N_1926,N_1720);
or U4200 (N_4200,N_2829,N_2717);
nand U4201 (N_4201,N_2885,N_2211);
xor U4202 (N_4202,N_1628,N_2317);
nand U4203 (N_4203,N_2068,N_1825);
xnor U4204 (N_4204,N_2411,N_2239);
nor U4205 (N_4205,N_2559,N_2269);
nor U4206 (N_4206,N_2926,N_2814);
and U4207 (N_4207,N_2055,N_2828);
nand U4208 (N_4208,N_1904,N_1561);
and U4209 (N_4209,N_2573,N_2371);
and U4210 (N_4210,N_2597,N_2539);
nand U4211 (N_4211,N_1684,N_1598);
nor U4212 (N_4212,N_2500,N_1919);
nand U4213 (N_4213,N_1796,N_1720);
or U4214 (N_4214,N_2019,N_2636);
or U4215 (N_4215,N_2011,N_2522);
or U4216 (N_4216,N_2757,N_2588);
nor U4217 (N_4217,N_2092,N_1573);
and U4218 (N_4218,N_2151,N_2254);
or U4219 (N_4219,N_2565,N_2878);
and U4220 (N_4220,N_1690,N_2596);
nor U4221 (N_4221,N_1569,N_1829);
nand U4222 (N_4222,N_2176,N_2275);
or U4223 (N_4223,N_2668,N_2387);
and U4224 (N_4224,N_1962,N_2200);
nor U4225 (N_4225,N_2718,N_2000);
and U4226 (N_4226,N_2864,N_2081);
nand U4227 (N_4227,N_2381,N_2207);
nor U4228 (N_4228,N_1776,N_2699);
nand U4229 (N_4229,N_2408,N_2085);
or U4230 (N_4230,N_2699,N_2597);
or U4231 (N_4231,N_2062,N_2260);
and U4232 (N_4232,N_2714,N_1936);
and U4233 (N_4233,N_1696,N_1616);
nand U4234 (N_4234,N_1676,N_1564);
xor U4235 (N_4235,N_2511,N_2309);
and U4236 (N_4236,N_2237,N_1948);
nand U4237 (N_4237,N_1701,N_1699);
nor U4238 (N_4238,N_2579,N_2217);
or U4239 (N_4239,N_2327,N_2490);
nand U4240 (N_4240,N_1742,N_1891);
nor U4241 (N_4241,N_2127,N_1774);
or U4242 (N_4242,N_2836,N_2898);
and U4243 (N_4243,N_2603,N_2491);
nor U4244 (N_4244,N_1718,N_2014);
nand U4245 (N_4245,N_2664,N_2780);
nor U4246 (N_4246,N_2300,N_2428);
xnor U4247 (N_4247,N_1573,N_2557);
nor U4248 (N_4248,N_1938,N_1772);
or U4249 (N_4249,N_2126,N_2772);
nor U4250 (N_4250,N_2182,N_2960);
nand U4251 (N_4251,N_2261,N_2921);
nor U4252 (N_4252,N_2829,N_2948);
and U4253 (N_4253,N_2639,N_1878);
nand U4254 (N_4254,N_2632,N_2053);
and U4255 (N_4255,N_2597,N_2358);
and U4256 (N_4256,N_2005,N_2184);
nor U4257 (N_4257,N_2827,N_2394);
nand U4258 (N_4258,N_1994,N_2511);
nor U4259 (N_4259,N_2192,N_2366);
nand U4260 (N_4260,N_1570,N_2138);
or U4261 (N_4261,N_2951,N_2186);
and U4262 (N_4262,N_2090,N_2934);
nor U4263 (N_4263,N_1543,N_2575);
nor U4264 (N_4264,N_2717,N_1887);
or U4265 (N_4265,N_1835,N_1688);
nand U4266 (N_4266,N_2601,N_2969);
or U4267 (N_4267,N_2678,N_2205);
xor U4268 (N_4268,N_2580,N_1852);
nor U4269 (N_4269,N_2452,N_2821);
xnor U4270 (N_4270,N_2147,N_2746);
and U4271 (N_4271,N_1827,N_2649);
nand U4272 (N_4272,N_2386,N_2146);
nand U4273 (N_4273,N_2063,N_2670);
and U4274 (N_4274,N_2906,N_2351);
or U4275 (N_4275,N_2453,N_1813);
or U4276 (N_4276,N_2242,N_2695);
or U4277 (N_4277,N_1676,N_1662);
or U4278 (N_4278,N_2553,N_2905);
nor U4279 (N_4279,N_2857,N_2361);
or U4280 (N_4280,N_1777,N_2902);
and U4281 (N_4281,N_1566,N_2765);
and U4282 (N_4282,N_2284,N_2962);
or U4283 (N_4283,N_2974,N_2183);
and U4284 (N_4284,N_2463,N_1918);
xnor U4285 (N_4285,N_1607,N_1946);
nand U4286 (N_4286,N_2523,N_1618);
xor U4287 (N_4287,N_2698,N_2645);
nor U4288 (N_4288,N_2924,N_2306);
xnor U4289 (N_4289,N_1984,N_2900);
or U4290 (N_4290,N_2641,N_2370);
or U4291 (N_4291,N_1732,N_2027);
nor U4292 (N_4292,N_2089,N_2094);
or U4293 (N_4293,N_2882,N_2256);
nand U4294 (N_4294,N_1634,N_2520);
nor U4295 (N_4295,N_1854,N_2970);
nand U4296 (N_4296,N_2562,N_2175);
and U4297 (N_4297,N_2193,N_2738);
nor U4298 (N_4298,N_2478,N_2792);
and U4299 (N_4299,N_2077,N_2180);
nor U4300 (N_4300,N_2302,N_2561);
nor U4301 (N_4301,N_2073,N_2882);
nand U4302 (N_4302,N_2334,N_2805);
or U4303 (N_4303,N_1590,N_1878);
xor U4304 (N_4304,N_2425,N_1833);
nand U4305 (N_4305,N_2776,N_2319);
nor U4306 (N_4306,N_1847,N_1835);
or U4307 (N_4307,N_2901,N_2383);
or U4308 (N_4308,N_1699,N_1577);
nor U4309 (N_4309,N_1633,N_1685);
nor U4310 (N_4310,N_2337,N_1591);
nand U4311 (N_4311,N_2309,N_2724);
and U4312 (N_4312,N_2938,N_2533);
nand U4313 (N_4313,N_2332,N_2361);
and U4314 (N_4314,N_2848,N_1803);
nor U4315 (N_4315,N_1565,N_1766);
nor U4316 (N_4316,N_1652,N_2471);
or U4317 (N_4317,N_2370,N_1652);
or U4318 (N_4318,N_2890,N_2552);
or U4319 (N_4319,N_1597,N_2197);
and U4320 (N_4320,N_2211,N_2089);
nor U4321 (N_4321,N_1615,N_1889);
and U4322 (N_4322,N_2739,N_1537);
xor U4323 (N_4323,N_1654,N_2530);
and U4324 (N_4324,N_2387,N_2940);
nor U4325 (N_4325,N_2469,N_1948);
and U4326 (N_4326,N_2029,N_1565);
nand U4327 (N_4327,N_2778,N_2430);
nand U4328 (N_4328,N_1588,N_2656);
nor U4329 (N_4329,N_2127,N_2842);
or U4330 (N_4330,N_2005,N_1799);
and U4331 (N_4331,N_2523,N_2001);
nor U4332 (N_4332,N_2528,N_1545);
and U4333 (N_4333,N_2731,N_2175);
nor U4334 (N_4334,N_2978,N_2818);
nor U4335 (N_4335,N_2443,N_1546);
nand U4336 (N_4336,N_2526,N_2718);
nand U4337 (N_4337,N_2025,N_2734);
nand U4338 (N_4338,N_2475,N_1833);
xor U4339 (N_4339,N_1938,N_2987);
or U4340 (N_4340,N_2620,N_1513);
or U4341 (N_4341,N_2071,N_2850);
nor U4342 (N_4342,N_2500,N_1654);
and U4343 (N_4343,N_1945,N_2376);
or U4344 (N_4344,N_1599,N_1764);
nor U4345 (N_4345,N_2010,N_2000);
nand U4346 (N_4346,N_2591,N_1828);
nor U4347 (N_4347,N_1511,N_2165);
and U4348 (N_4348,N_1674,N_2502);
nor U4349 (N_4349,N_1544,N_2743);
and U4350 (N_4350,N_2908,N_2282);
or U4351 (N_4351,N_2396,N_1977);
or U4352 (N_4352,N_2171,N_2315);
nand U4353 (N_4353,N_1742,N_2665);
and U4354 (N_4354,N_2494,N_1931);
nor U4355 (N_4355,N_2248,N_2018);
nor U4356 (N_4356,N_2503,N_2654);
and U4357 (N_4357,N_2873,N_2297);
and U4358 (N_4358,N_1951,N_2943);
and U4359 (N_4359,N_2205,N_2617);
or U4360 (N_4360,N_1980,N_2826);
nor U4361 (N_4361,N_1573,N_2540);
and U4362 (N_4362,N_2115,N_2474);
and U4363 (N_4363,N_1820,N_2106);
nand U4364 (N_4364,N_2446,N_2393);
nand U4365 (N_4365,N_2556,N_1833);
nor U4366 (N_4366,N_2688,N_1779);
and U4367 (N_4367,N_2554,N_2076);
or U4368 (N_4368,N_1687,N_2083);
nand U4369 (N_4369,N_2475,N_2463);
and U4370 (N_4370,N_1588,N_2860);
and U4371 (N_4371,N_2580,N_1869);
xnor U4372 (N_4372,N_2963,N_1626);
xor U4373 (N_4373,N_2065,N_1608);
and U4374 (N_4374,N_2260,N_1680);
or U4375 (N_4375,N_2557,N_2953);
and U4376 (N_4376,N_2364,N_2395);
and U4377 (N_4377,N_1779,N_2976);
nand U4378 (N_4378,N_2309,N_2018);
nand U4379 (N_4379,N_2776,N_2946);
nor U4380 (N_4380,N_1936,N_2786);
xor U4381 (N_4381,N_1816,N_2910);
and U4382 (N_4382,N_2349,N_1879);
and U4383 (N_4383,N_1660,N_2839);
or U4384 (N_4384,N_2805,N_2289);
nand U4385 (N_4385,N_2680,N_1955);
or U4386 (N_4386,N_2055,N_2570);
xnor U4387 (N_4387,N_2450,N_2032);
or U4388 (N_4388,N_2195,N_2876);
or U4389 (N_4389,N_2197,N_2633);
nor U4390 (N_4390,N_2220,N_2537);
nor U4391 (N_4391,N_1805,N_2265);
or U4392 (N_4392,N_2235,N_1590);
nand U4393 (N_4393,N_1516,N_2306);
nor U4394 (N_4394,N_2260,N_1726);
nand U4395 (N_4395,N_1600,N_2874);
and U4396 (N_4396,N_2053,N_1784);
xnor U4397 (N_4397,N_2155,N_2464);
or U4398 (N_4398,N_2747,N_1504);
nor U4399 (N_4399,N_2588,N_2494);
or U4400 (N_4400,N_2194,N_1864);
and U4401 (N_4401,N_2990,N_1504);
nand U4402 (N_4402,N_2750,N_2235);
xnor U4403 (N_4403,N_1700,N_2592);
or U4404 (N_4404,N_2170,N_2575);
nor U4405 (N_4405,N_2224,N_2594);
nand U4406 (N_4406,N_2945,N_2206);
nor U4407 (N_4407,N_2460,N_1889);
and U4408 (N_4408,N_1788,N_1771);
nand U4409 (N_4409,N_2961,N_1686);
or U4410 (N_4410,N_2124,N_1944);
nor U4411 (N_4411,N_1831,N_2517);
nand U4412 (N_4412,N_2356,N_1852);
or U4413 (N_4413,N_2360,N_2349);
or U4414 (N_4414,N_2390,N_2727);
nor U4415 (N_4415,N_2824,N_2857);
xnor U4416 (N_4416,N_2398,N_1911);
or U4417 (N_4417,N_2002,N_1800);
or U4418 (N_4418,N_1719,N_2299);
nand U4419 (N_4419,N_2590,N_1850);
nor U4420 (N_4420,N_2439,N_1801);
and U4421 (N_4421,N_1503,N_1825);
nand U4422 (N_4422,N_1549,N_2772);
or U4423 (N_4423,N_2592,N_2084);
nand U4424 (N_4424,N_2750,N_1729);
or U4425 (N_4425,N_2266,N_2881);
or U4426 (N_4426,N_2870,N_2582);
nor U4427 (N_4427,N_1742,N_2095);
nor U4428 (N_4428,N_2878,N_1958);
and U4429 (N_4429,N_2174,N_2022);
nand U4430 (N_4430,N_2790,N_2849);
nor U4431 (N_4431,N_1791,N_2153);
nand U4432 (N_4432,N_2547,N_2933);
and U4433 (N_4433,N_2955,N_2354);
or U4434 (N_4434,N_2446,N_1823);
or U4435 (N_4435,N_2192,N_1738);
nor U4436 (N_4436,N_1884,N_1967);
nand U4437 (N_4437,N_2008,N_2377);
nand U4438 (N_4438,N_2706,N_2185);
and U4439 (N_4439,N_2320,N_1948);
and U4440 (N_4440,N_2733,N_1554);
or U4441 (N_4441,N_2844,N_2930);
or U4442 (N_4442,N_1887,N_2880);
or U4443 (N_4443,N_1918,N_1902);
nor U4444 (N_4444,N_2217,N_2382);
nor U4445 (N_4445,N_2194,N_1831);
or U4446 (N_4446,N_2874,N_2029);
xnor U4447 (N_4447,N_2213,N_2141);
and U4448 (N_4448,N_2718,N_2204);
nand U4449 (N_4449,N_2860,N_1877);
xnor U4450 (N_4450,N_2763,N_2067);
nand U4451 (N_4451,N_2585,N_2405);
or U4452 (N_4452,N_2535,N_1904);
xnor U4453 (N_4453,N_2919,N_2120);
xor U4454 (N_4454,N_2758,N_2121);
nor U4455 (N_4455,N_1739,N_2771);
xor U4456 (N_4456,N_2937,N_2180);
and U4457 (N_4457,N_2584,N_1906);
and U4458 (N_4458,N_2050,N_2232);
xor U4459 (N_4459,N_2928,N_2057);
and U4460 (N_4460,N_1878,N_2047);
and U4461 (N_4461,N_2293,N_2306);
nor U4462 (N_4462,N_2303,N_2850);
and U4463 (N_4463,N_2749,N_2169);
xnor U4464 (N_4464,N_2225,N_2629);
xor U4465 (N_4465,N_2170,N_1998);
nor U4466 (N_4466,N_2262,N_2313);
and U4467 (N_4467,N_2109,N_1752);
nand U4468 (N_4468,N_1847,N_1944);
or U4469 (N_4469,N_2360,N_1534);
or U4470 (N_4470,N_2401,N_1798);
nor U4471 (N_4471,N_1834,N_2737);
and U4472 (N_4472,N_2858,N_1722);
nor U4473 (N_4473,N_1851,N_2676);
nor U4474 (N_4474,N_2715,N_2879);
nor U4475 (N_4475,N_2345,N_2818);
or U4476 (N_4476,N_2364,N_1831);
nor U4477 (N_4477,N_2545,N_2859);
nand U4478 (N_4478,N_1746,N_1564);
xor U4479 (N_4479,N_2508,N_1929);
nand U4480 (N_4480,N_1600,N_2966);
nor U4481 (N_4481,N_2771,N_2569);
and U4482 (N_4482,N_2210,N_1942);
nand U4483 (N_4483,N_2295,N_2168);
nand U4484 (N_4484,N_2085,N_1988);
nor U4485 (N_4485,N_1798,N_1534);
and U4486 (N_4486,N_2738,N_2083);
nor U4487 (N_4487,N_1789,N_2590);
xor U4488 (N_4488,N_2888,N_1785);
xnor U4489 (N_4489,N_2198,N_2638);
nand U4490 (N_4490,N_2910,N_2707);
xor U4491 (N_4491,N_2500,N_2778);
nor U4492 (N_4492,N_2127,N_1851);
nand U4493 (N_4493,N_2030,N_2741);
or U4494 (N_4494,N_2711,N_2480);
nand U4495 (N_4495,N_2639,N_1681);
nor U4496 (N_4496,N_1868,N_2134);
or U4497 (N_4497,N_1905,N_2606);
or U4498 (N_4498,N_1904,N_1525);
nand U4499 (N_4499,N_2781,N_2619);
nor U4500 (N_4500,N_3435,N_3942);
and U4501 (N_4501,N_3106,N_4037);
and U4502 (N_4502,N_3980,N_3406);
and U4503 (N_4503,N_3950,N_4430);
nor U4504 (N_4504,N_3121,N_3838);
nor U4505 (N_4505,N_3241,N_3753);
nor U4506 (N_4506,N_3040,N_3978);
or U4507 (N_4507,N_3342,N_3655);
nor U4508 (N_4508,N_3494,N_3005);
or U4509 (N_4509,N_3683,N_3642);
and U4510 (N_4510,N_3270,N_3763);
nor U4511 (N_4511,N_3557,N_4347);
xor U4512 (N_4512,N_4401,N_3824);
xnor U4513 (N_4513,N_3138,N_3203);
nor U4514 (N_4514,N_3955,N_4487);
and U4515 (N_4515,N_3455,N_3305);
or U4516 (N_4516,N_3501,N_3625);
nor U4517 (N_4517,N_3880,N_4084);
xor U4518 (N_4518,N_3427,N_4197);
nand U4519 (N_4519,N_3362,N_3048);
nor U4520 (N_4520,N_3611,N_3000);
or U4521 (N_4521,N_3179,N_4396);
or U4522 (N_4522,N_3459,N_3626);
and U4523 (N_4523,N_3968,N_3224);
nand U4524 (N_4524,N_3214,N_3223);
and U4525 (N_4525,N_3065,N_4170);
nand U4526 (N_4526,N_3031,N_4132);
nand U4527 (N_4527,N_3189,N_4230);
nor U4528 (N_4528,N_3654,N_4425);
nor U4529 (N_4529,N_3096,N_3628);
and U4530 (N_4530,N_3656,N_3149);
nand U4531 (N_4531,N_4423,N_3566);
or U4532 (N_4532,N_3762,N_4195);
and U4533 (N_4533,N_4448,N_4204);
nand U4534 (N_4534,N_3727,N_3559);
nand U4535 (N_4535,N_3580,N_4360);
or U4536 (N_4536,N_4044,N_4367);
nand U4537 (N_4537,N_4129,N_4182);
or U4538 (N_4538,N_4461,N_3385);
nor U4539 (N_4539,N_4322,N_4394);
nor U4540 (N_4540,N_4474,N_3396);
nand U4541 (N_4541,N_3154,N_4026);
nand U4542 (N_4542,N_4240,N_3855);
nand U4543 (N_4543,N_3146,N_3939);
nor U4544 (N_4544,N_3132,N_4428);
nand U4545 (N_4545,N_3809,N_4496);
xor U4546 (N_4546,N_4450,N_3018);
and U4547 (N_4547,N_3380,N_3541);
or U4548 (N_4548,N_4316,N_3114);
nor U4549 (N_4549,N_3488,N_4387);
nand U4550 (N_4550,N_4146,N_3002);
or U4551 (N_4551,N_3721,N_4305);
and U4552 (N_4552,N_3877,N_3732);
or U4553 (N_4553,N_3907,N_3049);
nand U4554 (N_4554,N_3868,N_4335);
nor U4555 (N_4555,N_3982,N_4490);
or U4556 (N_4556,N_3785,N_4073);
nor U4557 (N_4557,N_3848,N_4268);
and U4558 (N_4558,N_3169,N_3116);
and U4559 (N_4559,N_4028,N_3148);
xnor U4560 (N_4560,N_4295,N_3467);
or U4561 (N_4561,N_4097,N_4093);
and U4562 (N_4562,N_3531,N_3818);
nand U4563 (N_4563,N_4482,N_3996);
nor U4564 (N_4564,N_3060,N_3830);
nand U4565 (N_4565,N_3572,N_3885);
xor U4566 (N_4566,N_4294,N_3082);
nor U4567 (N_4567,N_4143,N_4223);
or U4568 (N_4568,N_3402,N_3783);
xor U4569 (N_4569,N_3956,N_3073);
and U4570 (N_4570,N_4460,N_3252);
or U4571 (N_4571,N_3685,N_4329);
nand U4572 (N_4572,N_4087,N_3024);
nand U4573 (N_4573,N_3123,N_3847);
and U4574 (N_4574,N_3011,N_3101);
nand U4575 (N_4575,N_3480,N_4039);
or U4576 (N_4576,N_3367,N_3587);
nand U4577 (N_4577,N_3664,N_3786);
or U4578 (N_4578,N_3858,N_3299);
nand U4579 (N_4579,N_3886,N_3959);
or U4580 (N_4580,N_3567,N_3781);
nand U4581 (N_4581,N_3784,N_4236);
nor U4582 (N_4582,N_3411,N_3545);
xnor U4583 (N_4583,N_3248,N_4242);
nand U4584 (N_4584,N_3334,N_3921);
nor U4585 (N_4585,N_4331,N_3846);
or U4586 (N_4586,N_4019,N_3666);
nor U4587 (N_4587,N_4493,N_3387);
or U4588 (N_4588,N_3012,N_3193);
or U4589 (N_4589,N_3679,N_3449);
nand U4590 (N_4590,N_3794,N_3039);
nor U4591 (N_4591,N_3481,N_3926);
or U4592 (N_4592,N_3124,N_3941);
and U4593 (N_4593,N_3057,N_3551);
or U4594 (N_4594,N_4250,N_3987);
or U4595 (N_4595,N_3760,N_3358);
nor U4596 (N_4596,N_4036,N_3902);
and U4597 (N_4597,N_3303,N_4272);
or U4598 (N_4598,N_3033,N_3069);
and U4599 (N_4599,N_3554,N_4210);
and U4600 (N_4600,N_4465,N_4131);
nor U4601 (N_4601,N_3620,N_3401);
or U4602 (N_4602,N_4116,N_3227);
nor U4603 (N_4603,N_3979,N_4366);
nand U4604 (N_4604,N_3696,N_3776);
and U4605 (N_4605,N_3053,N_3875);
and U4606 (N_4606,N_3294,N_3135);
and U4607 (N_4607,N_3475,N_3465);
and U4608 (N_4608,N_3974,N_3930);
and U4609 (N_4609,N_3341,N_4311);
or U4610 (N_4610,N_3232,N_3474);
and U4611 (N_4611,N_4441,N_3969);
or U4612 (N_4612,N_4163,N_3262);
nand U4613 (N_4613,N_3859,N_3328);
nor U4614 (N_4614,N_3756,N_3623);
nor U4615 (N_4615,N_4162,N_3307);
and U4616 (N_4616,N_3920,N_3616);
and U4617 (N_4617,N_3092,N_3340);
xor U4618 (N_4618,N_4386,N_4446);
nand U4619 (N_4619,N_3729,N_3218);
xnor U4620 (N_4620,N_3538,N_4255);
and U4621 (N_4621,N_3374,N_3471);
nand U4622 (N_4622,N_3400,N_3463);
nand U4623 (N_4623,N_3842,N_3194);
and U4624 (N_4624,N_4390,N_4058);
nand U4625 (N_4625,N_4383,N_3278);
and U4626 (N_4626,N_3993,N_3243);
nand U4627 (N_4627,N_3726,N_4222);
nand U4628 (N_4628,N_4439,N_4300);
nand U4629 (N_4629,N_3681,N_3422);
nand U4630 (N_4630,N_3010,N_3535);
or U4631 (N_4631,N_3713,N_3035);
nand U4632 (N_4632,N_4385,N_4106);
and U4633 (N_4633,N_3433,N_3196);
or U4634 (N_4634,N_3759,N_3686);
nor U4635 (N_4635,N_3394,N_4147);
nor U4636 (N_4636,N_3235,N_3582);
and U4637 (N_4637,N_4302,N_4171);
and U4638 (N_4638,N_3943,N_4371);
nor U4639 (N_4639,N_4160,N_3302);
nor U4640 (N_4640,N_4091,N_3122);
nor U4641 (N_4641,N_3928,N_3962);
nand U4642 (N_4642,N_3780,N_3349);
nor U4643 (N_4643,N_3316,N_3970);
xor U4644 (N_4644,N_4090,N_3163);
or U4645 (N_4645,N_3238,N_3524);
nand U4646 (N_4646,N_3404,N_3895);
nand U4647 (N_4647,N_4382,N_3280);
nand U4648 (N_4648,N_3577,N_3403);
and U4649 (N_4649,N_3491,N_3355);
and U4650 (N_4650,N_4225,N_4442);
nand U4651 (N_4651,N_3100,N_3198);
or U4652 (N_4652,N_3306,N_4488);
nand U4653 (N_4653,N_3339,N_3560);
nand U4654 (N_4654,N_3782,N_3151);
xor U4655 (N_4655,N_3703,N_4440);
and U4656 (N_4656,N_3917,N_3910);
nand U4657 (N_4657,N_4486,N_3127);
nand U4658 (N_4658,N_4475,N_3896);
or U4659 (N_4659,N_4320,N_3201);
nand U4660 (N_4660,N_4009,N_4117);
xor U4661 (N_4661,N_3790,N_4031);
nor U4662 (N_4662,N_3849,N_3253);
nor U4663 (N_4663,N_3225,N_4103);
and U4664 (N_4664,N_4296,N_4115);
or U4665 (N_4665,N_4457,N_4310);
nor U4666 (N_4666,N_3515,N_3212);
nand U4667 (N_4667,N_3213,N_3343);
nand U4668 (N_4668,N_3923,N_3884);
and U4669 (N_4669,N_3722,N_3388);
nand U4670 (N_4670,N_3797,N_3323);
xor U4671 (N_4671,N_3561,N_4027);
nand U4672 (N_4672,N_4484,N_3022);
nand U4673 (N_4673,N_4071,N_3694);
nor U4674 (N_4674,N_4054,N_4246);
and U4675 (N_4675,N_4104,N_4133);
xor U4676 (N_4676,N_4410,N_3317);
and U4677 (N_4677,N_3177,N_3505);
nand U4678 (N_4678,N_4224,N_4001);
nand U4679 (N_4679,N_3431,N_4232);
or U4680 (N_4680,N_3321,N_3511);
and U4681 (N_4681,N_3382,N_3245);
or U4682 (N_4682,N_4243,N_4291);
or U4683 (N_4683,N_3803,N_4041);
nor U4684 (N_4684,N_4288,N_3417);
nor U4685 (N_4685,N_4489,N_4023);
and U4686 (N_4686,N_3140,N_4076);
or U4687 (N_4687,N_3940,N_3992);
nor U4688 (N_4688,N_3166,N_3688);
or U4689 (N_4689,N_3247,N_3016);
nor U4690 (N_4690,N_4277,N_4048);
nand U4691 (N_4691,N_3586,N_3264);
nand U4692 (N_4692,N_3630,N_3874);
or U4693 (N_4693,N_4168,N_3439);
and U4694 (N_4694,N_4145,N_3768);
nand U4695 (N_4695,N_3596,N_4180);
nor U4696 (N_4696,N_3640,N_3742);
xnor U4697 (N_4697,N_3322,N_3775);
and U4698 (N_4698,N_4262,N_3426);
or U4699 (N_4699,N_3102,N_4079);
and U4700 (N_4700,N_3960,N_3584);
nor U4701 (N_4701,N_3038,N_4021);
or U4702 (N_4702,N_3025,N_3935);
and U4703 (N_4703,N_4464,N_3222);
xnor U4704 (N_4704,N_3200,N_4343);
nor U4705 (N_4705,N_3936,N_4453);
nand U4706 (N_4706,N_4424,N_3922);
and U4707 (N_4707,N_4338,N_3347);
and U4708 (N_4708,N_3826,N_3714);
nor U4709 (N_4709,N_3424,N_3746);
and U4710 (N_4710,N_3291,N_3823);
nor U4711 (N_4711,N_3649,N_3613);
nand U4712 (N_4712,N_4319,N_4196);
and U4713 (N_4713,N_3639,N_3951);
nor U4714 (N_4714,N_3412,N_3054);
nor U4715 (N_4715,N_3453,N_4051);
nor U4716 (N_4716,N_4042,N_3164);
nand U4717 (N_4717,N_3160,N_4015);
nand U4718 (N_4718,N_3338,N_3576);
nand U4719 (N_4719,N_3953,N_4161);
nor U4720 (N_4720,N_3712,N_4426);
xnor U4721 (N_4721,N_4176,N_3525);
xor U4722 (N_4722,N_3393,N_3904);
and U4723 (N_4723,N_4353,N_4267);
nand U4724 (N_4724,N_4467,N_3704);
or U4725 (N_4725,N_4415,N_3632);
nand U4726 (N_4726,N_3828,N_3444);
and U4727 (N_4727,N_3643,N_3041);
nand U4728 (N_4728,N_3606,N_3813);
or U4729 (N_4729,N_3944,N_3076);
xnor U4730 (N_4730,N_4238,N_3256);
and U4731 (N_4731,N_3258,N_4211);
nand U4732 (N_4732,N_3948,N_4315);
xor U4733 (N_4733,N_3677,N_3492);
nand U4734 (N_4734,N_3423,N_3389);
or U4735 (N_4735,N_3432,N_4417);
nand U4736 (N_4736,N_3635,N_3171);
xnor U4737 (N_4737,N_3029,N_3529);
nor U4738 (N_4738,N_4152,N_4138);
and U4739 (N_4739,N_4228,N_3711);
or U4740 (N_4740,N_3692,N_3812);
nand U4741 (N_4741,N_3691,N_3973);
nor U4742 (N_4742,N_4149,N_3274);
nand U4743 (N_4743,N_3251,N_4392);
nor U4744 (N_4744,N_3315,N_3185);
nor U4745 (N_4745,N_3326,N_3815);
or U4746 (N_4746,N_4378,N_4047);
nor U4747 (N_4747,N_3972,N_3330);
nor U4748 (N_4748,N_3377,N_3420);
nand U4749 (N_4749,N_4188,N_3633);
and U4750 (N_4750,N_4194,N_3070);
or U4751 (N_4751,N_3118,N_3650);
and U4752 (N_4752,N_3636,N_3373);
nor U4753 (N_4753,N_3622,N_3142);
or U4754 (N_4754,N_4234,N_3084);
nand U4755 (N_4755,N_4485,N_3878);
nand U4756 (N_4756,N_3836,N_3591);
and U4757 (N_4757,N_3631,N_3221);
xor U4758 (N_4758,N_4095,N_4017);
nand U4759 (N_4759,N_3188,N_3310);
or U4760 (N_4760,N_4127,N_3817);
and U4761 (N_4761,N_3129,N_3344);
xor U4762 (N_4762,N_3839,N_4256);
nor U4763 (N_4763,N_4356,N_4123);
and U4764 (N_4764,N_4139,N_3210);
nand U4765 (N_4765,N_3747,N_3473);
nor U4766 (N_4766,N_3787,N_3808);
nand U4767 (N_4767,N_3697,N_3006);
or U4768 (N_4768,N_3573,N_3105);
and U4769 (N_4769,N_3653,N_3044);
and U4770 (N_4770,N_3219,N_3231);
nand U4771 (N_4771,N_3067,N_4248);
and U4772 (N_4772,N_3663,N_4308);
nor U4773 (N_4773,N_4283,N_3043);
or U4774 (N_4774,N_3986,N_4444);
or U4775 (N_4775,N_4261,N_4433);
nand U4776 (N_4776,N_3670,N_3440);
nor U4777 (N_4777,N_3372,N_3725);
or U4778 (N_4778,N_4284,N_3181);
nor U4779 (N_4779,N_4056,N_4362);
or U4780 (N_4780,N_3020,N_4339);
nor U4781 (N_4781,N_4350,N_3599);
xnor U4782 (N_4782,N_4345,N_3564);
nor U4783 (N_4783,N_3736,N_4406);
nand U4784 (N_4784,N_3500,N_3845);
xor U4785 (N_4785,N_3365,N_4063);
xor U4786 (N_4786,N_3479,N_3995);
or U4787 (N_4787,N_3055,N_3282);
nor U4788 (N_4788,N_3695,N_4334);
and U4789 (N_4789,N_3856,N_4221);
and U4790 (N_4790,N_3876,N_3791);
nand U4791 (N_4791,N_4274,N_3614);
or U4792 (N_4792,N_3352,N_3673);
nor U4793 (N_4793,N_4030,N_3337);
xor U4794 (N_4794,N_3502,N_3217);
nand U4795 (N_4795,N_3047,N_3693);
and U4796 (N_4796,N_4134,N_3066);
or U4797 (N_4797,N_3383,N_3168);
or U4798 (N_4798,N_3216,N_4150);
nand U4799 (N_4799,N_3883,N_3175);
nand U4800 (N_4800,N_3007,N_4411);
nand U4801 (N_4801,N_3857,N_3289);
or U4802 (N_4802,N_4404,N_3764);
or U4803 (N_4803,N_3139,N_3802);
or U4804 (N_4804,N_3528,N_4323);
or U4805 (N_4805,N_4178,N_4456);
nor U4806 (N_4806,N_3772,N_3835);
nand U4807 (N_4807,N_3061,N_3254);
nand U4808 (N_4808,N_4218,N_3346);
or U4809 (N_4809,N_3965,N_4239);
and U4810 (N_4810,N_3165,N_3745);
xnor U4811 (N_4811,N_3843,N_3792);
or U4812 (N_4812,N_3126,N_3507);
nor U4813 (N_4813,N_3205,N_3113);
and U4814 (N_4814,N_3381,N_3119);
xnor U4815 (N_4815,N_3134,N_3230);
and U4816 (N_4816,N_4269,N_3071);
nand U4817 (N_4817,N_3450,N_3228);
nor U4818 (N_4818,N_3448,N_4402);
nand U4819 (N_4819,N_4109,N_3441);
nand U4820 (N_4820,N_3281,N_3668);
nor U4821 (N_4821,N_3510,N_3867);
nor U4822 (N_4822,N_3689,N_4033);
nor U4823 (N_4823,N_3313,N_4077);
nand U4824 (N_4824,N_3821,N_4083);
nand U4825 (N_4825,N_3752,N_3646);
nor U4826 (N_4826,N_3309,N_3675);
or U4827 (N_4827,N_3568,N_3648);
nor U4828 (N_4828,N_3028,N_3518);
xnor U4829 (N_4829,N_4096,N_4011);
or U4830 (N_4830,N_3509,N_3170);
and U4831 (N_4831,N_3615,N_4443);
nor U4832 (N_4832,N_3700,N_3085);
xnor U4833 (N_4833,N_4355,N_3701);
nand U4834 (N_4834,N_3008,N_4251);
nand U4835 (N_4835,N_4298,N_4463);
nor U4836 (N_4836,N_3530,N_3516);
and U4837 (N_4837,N_3136,N_4376);
xor U4838 (N_4838,N_3112,N_3279);
nand U4839 (N_4839,N_4122,N_4307);
nor U4840 (N_4840,N_3128,N_3325);
or U4841 (N_4841,N_4244,N_4328);
and U4842 (N_4842,N_4226,N_3853);
nand U4843 (N_4843,N_3137,N_3314);
or U4844 (N_4844,N_3522,N_3523);
nand U4845 (N_4845,N_3977,N_3651);
xor U4846 (N_4846,N_3915,N_3312);
or U4847 (N_4847,N_3671,N_4275);
and U4848 (N_4848,N_4372,N_3644);
nor U4849 (N_4849,N_4301,N_4304);
xnor U4850 (N_4850,N_3718,N_3399);
or U4851 (N_4851,N_4388,N_4181);
or U4852 (N_4852,N_4368,N_4113);
or U4853 (N_4853,N_3037,N_4157);
or U4854 (N_4854,N_4422,N_4053);
nand U4855 (N_4855,N_3945,N_4016);
or U4856 (N_4856,N_3618,N_3534);
xor U4857 (N_4857,N_4330,N_4451);
and U4858 (N_4858,N_3336,N_3133);
nor U4859 (N_4859,N_3348,N_3796);
nand U4860 (N_4860,N_3144,N_3089);
or U4861 (N_4861,N_3147,N_3271);
xnor U4862 (N_4862,N_4190,N_3865);
nor U4863 (N_4863,N_4341,N_4193);
nor U4864 (N_4864,N_3997,N_4156);
nor U4865 (N_4865,N_3699,N_4429);
or U4866 (N_4866,N_3998,N_4481);
and U4867 (N_4867,N_3097,N_4081);
nor U4868 (N_4868,N_3023,N_3478);
or U4869 (N_4869,N_4070,N_3735);
nand U4870 (N_4870,N_4124,N_4389);
and U4871 (N_4871,N_3825,N_4349);
nand U4872 (N_4872,N_3659,N_4061);
nand U4873 (N_4873,N_4260,N_3539);
nor U4874 (N_4874,N_3709,N_4292);
xor U4875 (N_4875,N_3589,N_3609);
and U4876 (N_4876,N_4142,N_3706);
nor U4877 (N_4877,N_4006,N_3487);
or U4878 (N_4878,N_4324,N_3298);
nand U4879 (N_4879,N_4498,N_3369);
nor U4880 (N_4880,N_4059,N_3192);
or U4881 (N_4881,N_4471,N_3800);
or U4882 (N_4882,N_3680,N_3414);
or U4883 (N_4883,N_3612,N_4420);
nand U4884 (N_4884,N_4379,N_4400);
and U4885 (N_4885,N_3707,N_4370);
and U4886 (N_4886,N_3255,N_3384);
or U4887 (N_4887,N_3434,N_3829);
and U4888 (N_4888,N_3822,N_3485);
or U4889 (N_4889,N_3887,N_4468);
or U4890 (N_4890,N_3131,N_4029);
and U4891 (N_4891,N_3543,N_4094);
or U4892 (N_4892,N_3015,N_3575);
nand U4893 (N_4893,N_4495,N_3226);
nor U4894 (N_4894,N_3864,N_3619);
and U4895 (N_4895,N_4049,N_3311);
nor U4896 (N_4896,N_4233,N_4351);
or U4897 (N_4897,N_3811,N_4192);
xnor U4898 (N_4898,N_3484,N_4003);
nand U4899 (N_4899,N_3779,N_3368);
nand U4900 (N_4900,N_3913,N_4212);
nor U4901 (N_4901,N_4395,N_3470);
or U4902 (N_4902,N_4235,N_4494);
or U4903 (N_4903,N_3929,N_4340);
nor U4904 (N_4904,N_4273,N_3111);
nor U4905 (N_4905,N_3483,N_3585);
nor U4906 (N_4906,N_4214,N_4231);
nand U4907 (N_4907,N_4068,N_4447);
or U4908 (N_4908,N_4069,N_4012);
nor U4909 (N_4909,N_3242,N_3269);
and U4910 (N_4910,N_3296,N_3087);
or U4911 (N_4911,N_3045,N_4144);
nor U4912 (N_4912,N_4259,N_3167);
nand U4913 (N_4913,N_3908,N_3728);
or U4914 (N_4914,N_3287,N_3295);
nor U4915 (N_4915,N_3056,N_3017);
nand U4916 (N_4916,N_4175,N_4459);
or U4917 (N_4917,N_4111,N_3571);
nand U4918 (N_4918,N_4452,N_3851);
nor U4919 (N_4919,N_4492,N_4164);
nand U4920 (N_4920,N_3579,N_3263);
nand U4921 (N_4921,N_3027,N_3852);
nor U4922 (N_4922,N_3985,N_3761);
xor U4923 (N_4923,N_4409,N_4241);
nand U4924 (N_4924,N_4432,N_3120);
nand U4925 (N_4925,N_4120,N_4419);
or U4926 (N_4926,N_3621,N_3984);
nand U4927 (N_4927,N_4365,N_3195);
nor U4928 (N_4928,N_4314,N_3766);
nor U4929 (N_4929,N_3174,N_3319);
and U4930 (N_4930,N_3418,N_4247);
nor U4931 (N_4931,N_3009,N_3098);
or U4932 (N_4932,N_3145,N_4128);
nand U4933 (N_4933,N_3257,N_3155);
and U4934 (N_4934,N_4408,N_3837);
xor U4935 (N_4935,N_3861,N_4369);
nor U4936 (N_4936,N_4306,N_3240);
xnor U4937 (N_4937,N_3103,N_4321);
nor U4938 (N_4938,N_4121,N_3486);
and U4939 (N_4939,N_3593,N_3873);
or U4940 (N_4940,N_3079,N_3359);
nor U4941 (N_4941,N_4289,N_4318);
or U4942 (N_4942,N_3215,N_3769);
nor U4943 (N_4943,N_3891,N_3597);
and U4944 (N_4944,N_3261,N_3905);
nor U4945 (N_4945,N_4013,N_3464);
nand U4946 (N_4946,N_3909,N_4470);
nor U4947 (N_4947,N_3652,N_3831);
and U4948 (N_4948,N_3392,N_3526);
or U4949 (N_4949,N_3117,N_4159);
nand U4950 (N_4950,N_3157,N_4297);
and U4951 (N_4951,N_3419,N_3335);
nor U4952 (N_4952,N_4000,N_4332);
or U4953 (N_4953,N_4346,N_3806);
or U4954 (N_4954,N_3860,N_4399);
and U4955 (N_4955,N_3207,N_3078);
xor U4956 (N_4956,N_4279,N_4022);
nor U4957 (N_4957,N_4333,N_3496);
nor U4958 (N_4958,N_4397,N_4045);
or U4959 (N_4959,N_3237,N_3378);
or U4960 (N_4960,N_3260,N_3125);
or U4961 (N_4961,N_3684,N_3546);
xor U4962 (N_4962,N_3436,N_4174);
nor U4963 (N_4963,N_3919,N_3916);
nand U4964 (N_4964,N_3042,N_3517);
or U4965 (N_4965,N_3641,N_3717);
xor U4966 (N_4966,N_4435,N_3594);
nor U4967 (N_4967,N_3413,N_4062);
nand U4968 (N_4968,N_3946,N_3866);
nor U4969 (N_4969,N_3482,N_3647);
or U4970 (N_4970,N_3397,N_4398);
nor U4971 (N_4971,N_3454,N_3442);
and U4972 (N_4972,N_3019,N_4359);
nand U4973 (N_4973,N_4427,N_3268);
and U4974 (N_4974,N_4472,N_3988);
or U4975 (N_4975,N_3527,N_3156);
and U4976 (N_4976,N_4177,N_3892);
or U4977 (N_4977,N_4454,N_3428);
or U4978 (N_4978,N_3050,N_3981);
nand U4979 (N_4979,N_3932,N_3143);
nand U4980 (N_4980,N_3710,N_3190);
and U4981 (N_4981,N_4187,N_3519);
and U4982 (N_4982,N_3911,N_4098);
nand U4983 (N_4983,N_4374,N_4153);
and U4984 (N_4984,N_4449,N_3608);
nand U4985 (N_4985,N_4086,N_4245);
nor U4986 (N_4986,N_3461,N_3451);
nand U4987 (N_4987,N_4140,N_3975);
nand U4988 (N_4988,N_3533,N_4391);
xnor U4989 (N_4989,N_3810,N_3588);
nor U4990 (N_4990,N_3958,N_4491);
nor U4991 (N_4991,N_3964,N_3889);
or U4992 (N_4992,N_3208,N_4034);
nand U4993 (N_4993,N_3906,N_4309);
nand U4994 (N_4994,N_3390,N_3331);
nor U4995 (N_4995,N_4055,N_3765);
nor U4996 (N_4996,N_3046,N_4183);
or U4997 (N_4997,N_4141,N_3108);
nand U4998 (N_4998,N_4201,N_4198);
and U4999 (N_4999,N_3773,N_3356);
and U5000 (N_5000,N_3366,N_4110);
nand U5001 (N_5001,N_3493,N_3293);
nand U5002 (N_5002,N_4108,N_3900);
and U5003 (N_5003,N_3150,N_3605);
and U5004 (N_5004,N_3793,N_3267);
or U5005 (N_5005,N_4271,N_4455);
nor U5006 (N_5006,N_3276,N_3462);
or U5007 (N_5007,N_4361,N_3739);
or U5008 (N_5008,N_4155,N_4130);
or U5009 (N_5009,N_3804,N_4018);
or U5010 (N_5010,N_3583,N_3233);
nor U5011 (N_5011,N_3537,N_3778);
xor U5012 (N_5012,N_4167,N_3871);
or U5013 (N_5013,N_4278,N_4137);
nor U5014 (N_5014,N_3409,N_4072);
nand U5015 (N_5015,N_3197,N_3607);
or U5016 (N_5016,N_3246,N_4281);
nand U5017 (N_5017,N_4327,N_3807);
nand U5018 (N_5018,N_4148,N_3199);
or U5019 (N_5019,N_3840,N_3407);
nor U5020 (N_5020,N_3898,N_3063);
and U5021 (N_5021,N_3602,N_3272);
and U5022 (N_5022,N_4413,N_4065);
or U5023 (N_5023,N_4480,N_3445);
nor U5024 (N_5024,N_4462,N_3059);
nor U5025 (N_5025,N_4219,N_4357);
or U5026 (N_5026,N_4265,N_3574);
or U5027 (N_5027,N_3211,N_3976);
nand U5028 (N_5028,N_3104,N_3410);
and U5029 (N_5029,N_4299,N_3771);
or U5030 (N_5030,N_4266,N_4080);
nor U5031 (N_5031,N_4217,N_4497);
nor U5032 (N_5032,N_4344,N_3026);
nand U5033 (N_5033,N_3890,N_3881);
or U5034 (N_5034,N_3495,N_4125);
and U5035 (N_5035,N_4412,N_3301);
nand U5036 (N_5036,N_3661,N_3521);
nand U5037 (N_5037,N_3805,N_4057);
nor U5038 (N_5038,N_4276,N_4282);
or U5039 (N_5039,N_3477,N_3540);
nor U5040 (N_5040,N_4100,N_3755);
or U5041 (N_5041,N_3547,N_3967);
nor U5042 (N_5042,N_4290,N_4473);
nand U5043 (N_5043,N_4336,N_4184);
and U5044 (N_5044,N_4257,N_3304);
and U5045 (N_5045,N_3719,N_4254);
nand U5046 (N_5046,N_4135,N_3052);
and U5047 (N_5047,N_4200,N_4136);
nand U5048 (N_5048,N_3130,N_3083);
and U5049 (N_5049,N_3952,N_4375);
or U5050 (N_5050,N_3429,N_3705);
xor U5051 (N_5051,N_3357,N_3110);
nor U5052 (N_5052,N_4434,N_3991);
nor U5053 (N_5053,N_3370,N_4354);
or U5054 (N_5054,N_4263,N_3658);
nand U5055 (N_5055,N_4431,N_3239);
nor U5056 (N_5056,N_3749,N_3080);
or U5057 (N_5057,N_4215,N_3629);
or U5058 (N_5058,N_3032,N_3767);
nand U5059 (N_5059,N_4038,N_4206);
or U5060 (N_5060,N_3452,N_3789);
and U5061 (N_5061,N_3416,N_3520);
nand U5062 (N_5062,N_3933,N_3924);
and U5063 (N_5063,N_4438,N_3879);
xor U5064 (N_5064,N_3740,N_3250);
and U5065 (N_5065,N_3513,N_3814);
or U5066 (N_5066,N_3265,N_3318);
and U5067 (N_5067,N_3954,N_3634);
or U5068 (N_5068,N_3363,N_3731);
xor U5069 (N_5069,N_3425,N_3744);
or U5070 (N_5070,N_4202,N_3284);
nand U5071 (N_5071,N_3415,N_3178);
or U5072 (N_5072,N_3820,N_3447);
and U5073 (N_5073,N_3074,N_3499);
nand U5074 (N_5074,N_3176,N_3329);
or U5075 (N_5075,N_3562,N_4220);
nor U5076 (N_5076,N_3667,N_3598);
xnor U5077 (N_5077,N_3446,N_4205);
nor U5078 (N_5078,N_3172,N_3672);
or U5079 (N_5079,N_4052,N_3162);
or U5080 (N_5080,N_3801,N_3081);
xnor U5081 (N_5081,N_4293,N_3665);
nand U5082 (N_5082,N_3581,N_3698);
nor U5083 (N_5083,N_3182,N_4092);
or U5084 (N_5084,N_3555,N_3099);
and U5085 (N_5085,N_3075,N_3361);
and U5086 (N_5086,N_4066,N_3934);
and U5087 (N_5087,N_3738,N_3220);
nand U5088 (N_5088,N_4107,N_3443);
nand U5089 (N_5089,N_4007,N_3183);
or U5090 (N_5090,N_3234,N_3669);
nor U5091 (N_5091,N_4249,N_3186);
nor U5092 (N_5092,N_3300,N_4179);
nand U5093 (N_5093,N_3720,N_3570);
xor U5094 (N_5094,N_4458,N_3963);
nor U5095 (N_5095,N_4252,N_4024);
nor U5096 (N_5096,N_4032,N_4207);
nand U5097 (N_5097,N_3003,N_3292);
nor U5098 (N_5098,N_4384,N_3437);
nor U5099 (N_5099,N_3350,N_3638);
nor U5100 (N_5100,N_3754,N_4208);
or U5101 (N_5101,N_4337,N_3737);
xor U5102 (N_5102,N_3748,N_3503);
nand U5103 (N_5103,N_4040,N_3184);
nand U5104 (N_5104,N_3914,N_3645);
and U5105 (N_5105,N_3062,N_4209);
nor U5106 (N_5106,N_3662,N_3592);
nor U5107 (N_5107,N_3508,N_3816);
nand U5108 (N_5108,N_3229,N_3903);
nor U5109 (N_5109,N_4381,N_3925);
and U5110 (N_5110,N_4203,N_3989);
and U5111 (N_5111,N_3068,N_3285);
nor U5112 (N_5112,N_3244,N_3209);
and U5113 (N_5113,N_3458,N_3690);
and U5114 (N_5114,N_4199,N_3273);
or U5115 (N_5115,N_3819,N_3354);
xor U5116 (N_5116,N_3109,N_4105);
xor U5117 (N_5117,N_3536,N_3795);
and U5118 (N_5118,N_3173,N_4005);
nor U5119 (N_5119,N_3637,N_3072);
nand U5120 (N_5120,N_3107,N_4172);
nor U5121 (N_5121,N_3833,N_3093);
nand U5122 (N_5122,N_3894,N_3832);
nand U5123 (N_5123,N_3553,N_3506);
nand U5124 (N_5124,N_3489,N_3724);
or U5125 (N_5125,N_3532,N_3565);
nor U5126 (N_5126,N_3206,N_3715);
and U5127 (N_5127,N_3798,N_4380);
nand U5128 (N_5128,N_3617,N_3834);
nand U5129 (N_5129,N_4165,N_4166);
or U5130 (N_5130,N_4437,N_4060);
nand U5131 (N_5131,N_4102,N_3090);
nand U5132 (N_5132,N_3777,N_3799);
xnor U5133 (N_5133,N_3332,N_3590);
and U5134 (N_5134,N_3734,N_3512);
nand U5135 (N_5135,N_3949,N_3141);
nor U5136 (N_5136,N_3757,N_3774);
and U5137 (N_5137,N_3869,N_3058);
or U5138 (N_5138,N_3994,N_3204);
nand U5139 (N_5139,N_4285,N_3468);
and U5140 (N_5140,N_3386,N_4436);
nor U5141 (N_5141,N_3901,N_3034);
and U5142 (N_5142,N_3862,N_4088);
or U5143 (N_5143,N_3014,N_3660);
or U5144 (N_5144,N_3674,N_3333);
nand U5145 (N_5145,N_3723,N_3405);
xnor U5146 (N_5146,N_3202,N_3320);
and U5147 (N_5147,N_4342,N_3957);
xor U5148 (N_5148,N_4280,N_3277);
nor U5149 (N_5149,N_3391,N_4326);
nor U5150 (N_5150,N_3983,N_4020);
or U5151 (N_5151,N_3161,N_3091);
or U5152 (N_5152,N_3460,N_3086);
nand U5153 (N_5153,N_3364,N_4189);
nor U5154 (N_5154,N_4078,N_4010);
or U5155 (N_5155,N_3498,N_3918);
or U5156 (N_5156,N_4258,N_4004);
nand U5157 (N_5157,N_3021,N_3395);
or U5158 (N_5158,N_3872,N_3999);
nor U5159 (N_5159,N_3870,N_3476);
nor U5160 (N_5160,N_3259,N_4303);
and U5161 (N_5161,N_4227,N_4477);
and U5162 (N_5162,N_4476,N_3236);
or U5163 (N_5163,N_3376,N_3882);
xnor U5164 (N_5164,N_3550,N_4317);
nor U5165 (N_5165,N_4445,N_4479);
xnor U5166 (N_5166,N_3353,N_4416);
and U5167 (N_5167,N_3490,N_3327);
and U5168 (N_5168,N_3610,N_3360);
nor U5169 (N_5169,N_3603,N_4075);
and U5170 (N_5170,N_3730,N_4119);
nand U5171 (N_5171,N_4064,N_4126);
and U5172 (N_5172,N_4185,N_3379);
or U5173 (N_5173,N_3678,N_4067);
and U5174 (N_5174,N_3159,N_3472);
or U5175 (N_5175,N_3931,N_4008);
xnor U5176 (N_5176,N_4421,N_4253);
nand U5177 (N_5177,N_4085,N_4101);
and U5178 (N_5178,N_3716,N_4405);
nand U5179 (N_5179,N_4414,N_4466);
and U5180 (N_5180,N_3051,N_3758);
or U5181 (N_5181,N_3095,N_3863);
and U5182 (N_5182,N_4112,N_3421);
nand U5183 (N_5183,N_4186,N_3375);
nand U5184 (N_5184,N_4312,N_4325);
nand U5185 (N_5185,N_3595,N_4270);
nand U5186 (N_5186,N_3888,N_3297);
nor U5187 (N_5187,N_3308,N_3854);
or U5188 (N_5188,N_3249,N_3153);
nor U5189 (N_5189,N_3013,N_4118);
and U5190 (N_5190,N_4407,N_3733);
xnor U5191 (N_5191,N_3682,N_4264);
nand U5192 (N_5192,N_3947,N_4151);
xnor U5193 (N_5193,N_3457,N_4352);
nor U5194 (N_5194,N_3004,N_3841);
or U5195 (N_5195,N_3558,N_3899);
or U5196 (N_5196,N_3578,N_4154);
nor U5197 (N_5197,N_3514,N_3030);
or U5198 (N_5198,N_3544,N_3912);
and U5199 (N_5199,N_3556,N_4173);
nand U5200 (N_5200,N_4191,N_4237);
nand U5201 (N_5201,N_3094,N_3743);
nand U5202 (N_5202,N_3469,N_4035);
or U5203 (N_5203,N_3275,N_3938);
and U5204 (N_5204,N_4393,N_4469);
and U5205 (N_5205,N_3563,N_3750);
and U5206 (N_5206,N_3708,N_3497);
nand U5207 (N_5207,N_4099,N_3036);
or U5208 (N_5208,N_4043,N_4364);
or U5209 (N_5209,N_4046,N_3158);
or U5210 (N_5210,N_3600,N_3398);
nand U5211 (N_5211,N_4363,N_3937);
or U5212 (N_5212,N_3180,N_3286);
and U5213 (N_5213,N_3408,N_3676);
nand U5214 (N_5214,N_4050,N_4014);
nor U5215 (N_5215,N_3971,N_4403);
or U5216 (N_5216,N_3702,N_4158);
nand U5217 (N_5217,N_3351,N_4358);
and U5218 (N_5218,N_3604,N_3751);
and U5219 (N_5219,N_3345,N_4229);
nor U5220 (N_5220,N_3504,N_4418);
or U5221 (N_5221,N_3788,N_3077);
or U5222 (N_5222,N_3266,N_4169);
nand U5223 (N_5223,N_4082,N_3961);
xnor U5224 (N_5224,N_3844,N_4483);
nor U5225 (N_5225,N_3187,N_3601);
or U5226 (N_5226,N_3548,N_4286);
and U5227 (N_5227,N_3624,N_4114);
and U5228 (N_5228,N_3552,N_3324);
or U5229 (N_5229,N_4089,N_3088);
nor U5230 (N_5230,N_3001,N_3897);
nand U5231 (N_5231,N_4499,N_3430);
nand U5232 (N_5232,N_3115,N_3893);
and U5233 (N_5233,N_3152,N_3966);
nor U5234 (N_5234,N_3371,N_3283);
or U5235 (N_5235,N_3827,N_4216);
or U5236 (N_5236,N_3290,N_3687);
nand U5237 (N_5237,N_3288,N_3657);
and U5238 (N_5238,N_3466,N_4002);
or U5239 (N_5239,N_4313,N_3927);
nor U5240 (N_5240,N_3569,N_3741);
nor U5241 (N_5241,N_3064,N_4213);
and U5242 (N_5242,N_4478,N_4348);
or U5243 (N_5243,N_4287,N_3770);
nor U5244 (N_5244,N_3850,N_3542);
and U5245 (N_5245,N_4373,N_4377);
and U5246 (N_5246,N_4025,N_3990);
and U5247 (N_5247,N_3456,N_3627);
or U5248 (N_5248,N_4074,N_3191);
and U5249 (N_5249,N_3549,N_3438);
nor U5250 (N_5250,N_3597,N_3060);
and U5251 (N_5251,N_3833,N_3162);
xor U5252 (N_5252,N_4493,N_4055);
nand U5253 (N_5253,N_3809,N_3754);
or U5254 (N_5254,N_4326,N_3718);
nor U5255 (N_5255,N_3214,N_3117);
or U5256 (N_5256,N_3198,N_4414);
and U5257 (N_5257,N_4188,N_4448);
nand U5258 (N_5258,N_3835,N_3766);
and U5259 (N_5259,N_4313,N_3556);
nand U5260 (N_5260,N_3938,N_3092);
nor U5261 (N_5261,N_3979,N_3641);
xnor U5262 (N_5262,N_4159,N_4271);
nand U5263 (N_5263,N_3291,N_3012);
xnor U5264 (N_5264,N_3668,N_4080);
or U5265 (N_5265,N_4137,N_4353);
nand U5266 (N_5266,N_3453,N_3224);
and U5267 (N_5267,N_3241,N_3629);
or U5268 (N_5268,N_4239,N_4412);
nor U5269 (N_5269,N_3274,N_4097);
and U5270 (N_5270,N_3225,N_3018);
nor U5271 (N_5271,N_3695,N_4126);
or U5272 (N_5272,N_4327,N_3865);
xnor U5273 (N_5273,N_3879,N_3398);
nor U5274 (N_5274,N_3165,N_3975);
xor U5275 (N_5275,N_3266,N_3056);
and U5276 (N_5276,N_3895,N_4222);
xnor U5277 (N_5277,N_3542,N_3564);
and U5278 (N_5278,N_3712,N_3926);
nand U5279 (N_5279,N_4138,N_3890);
and U5280 (N_5280,N_4029,N_4214);
or U5281 (N_5281,N_3083,N_4442);
nor U5282 (N_5282,N_3462,N_4498);
and U5283 (N_5283,N_4016,N_3003);
nand U5284 (N_5284,N_3915,N_3895);
or U5285 (N_5285,N_4486,N_4198);
nand U5286 (N_5286,N_3096,N_3058);
nor U5287 (N_5287,N_4252,N_3574);
xor U5288 (N_5288,N_4028,N_4436);
and U5289 (N_5289,N_3018,N_3058);
xor U5290 (N_5290,N_3691,N_3303);
xor U5291 (N_5291,N_3149,N_4176);
nor U5292 (N_5292,N_3410,N_3896);
or U5293 (N_5293,N_3437,N_4357);
or U5294 (N_5294,N_3191,N_4044);
nand U5295 (N_5295,N_4168,N_4017);
or U5296 (N_5296,N_3226,N_3575);
nor U5297 (N_5297,N_4079,N_3084);
or U5298 (N_5298,N_4112,N_4404);
or U5299 (N_5299,N_4100,N_4231);
nor U5300 (N_5300,N_4337,N_4194);
nor U5301 (N_5301,N_4112,N_3257);
nand U5302 (N_5302,N_4319,N_4086);
nand U5303 (N_5303,N_3292,N_3994);
or U5304 (N_5304,N_3195,N_3129);
and U5305 (N_5305,N_3086,N_3345);
or U5306 (N_5306,N_3358,N_3168);
nor U5307 (N_5307,N_3763,N_3180);
and U5308 (N_5308,N_3679,N_3860);
or U5309 (N_5309,N_3159,N_4229);
nor U5310 (N_5310,N_3403,N_4197);
and U5311 (N_5311,N_3381,N_3787);
nor U5312 (N_5312,N_4194,N_3790);
or U5313 (N_5313,N_3350,N_4073);
nor U5314 (N_5314,N_3790,N_3585);
nand U5315 (N_5315,N_3986,N_3601);
nand U5316 (N_5316,N_4013,N_3356);
nor U5317 (N_5317,N_3062,N_3581);
and U5318 (N_5318,N_3881,N_4229);
nor U5319 (N_5319,N_4376,N_3446);
nor U5320 (N_5320,N_3194,N_3075);
xor U5321 (N_5321,N_3493,N_3247);
xnor U5322 (N_5322,N_4351,N_3118);
nor U5323 (N_5323,N_3045,N_3433);
or U5324 (N_5324,N_3207,N_4273);
xor U5325 (N_5325,N_3871,N_4141);
and U5326 (N_5326,N_3012,N_4062);
nand U5327 (N_5327,N_3238,N_3127);
nor U5328 (N_5328,N_3881,N_4130);
or U5329 (N_5329,N_3528,N_3703);
and U5330 (N_5330,N_3222,N_4332);
xor U5331 (N_5331,N_3998,N_3686);
nor U5332 (N_5332,N_3095,N_3987);
and U5333 (N_5333,N_4237,N_3491);
or U5334 (N_5334,N_4377,N_3752);
nand U5335 (N_5335,N_3502,N_3988);
nor U5336 (N_5336,N_3554,N_3314);
or U5337 (N_5337,N_4073,N_3526);
xnor U5338 (N_5338,N_4210,N_3060);
or U5339 (N_5339,N_3153,N_4304);
nor U5340 (N_5340,N_3335,N_3295);
nor U5341 (N_5341,N_3580,N_3319);
or U5342 (N_5342,N_3570,N_4041);
xnor U5343 (N_5343,N_3167,N_4459);
and U5344 (N_5344,N_3140,N_3987);
nor U5345 (N_5345,N_3550,N_3674);
or U5346 (N_5346,N_4324,N_3428);
or U5347 (N_5347,N_3438,N_3759);
nor U5348 (N_5348,N_3880,N_4307);
nand U5349 (N_5349,N_3917,N_3626);
or U5350 (N_5350,N_3801,N_3762);
nor U5351 (N_5351,N_3865,N_3921);
nor U5352 (N_5352,N_3984,N_3587);
nand U5353 (N_5353,N_3479,N_3040);
nor U5354 (N_5354,N_3782,N_4125);
nor U5355 (N_5355,N_4135,N_4215);
nor U5356 (N_5356,N_3668,N_3284);
nand U5357 (N_5357,N_3707,N_3023);
and U5358 (N_5358,N_3763,N_4138);
nand U5359 (N_5359,N_4348,N_3865);
nand U5360 (N_5360,N_3555,N_3488);
nand U5361 (N_5361,N_3255,N_3326);
or U5362 (N_5362,N_3329,N_3638);
xor U5363 (N_5363,N_4291,N_3849);
or U5364 (N_5364,N_3998,N_3250);
xnor U5365 (N_5365,N_3794,N_4411);
nor U5366 (N_5366,N_3084,N_3190);
xor U5367 (N_5367,N_3174,N_3073);
xnor U5368 (N_5368,N_4483,N_3134);
nand U5369 (N_5369,N_3588,N_3434);
xor U5370 (N_5370,N_3375,N_4038);
nand U5371 (N_5371,N_3074,N_3510);
nor U5372 (N_5372,N_4067,N_3064);
and U5373 (N_5373,N_4478,N_4055);
and U5374 (N_5374,N_3385,N_3169);
nor U5375 (N_5375,N_4208,N_4454);
or U5376 (N_5376,N_4127,N_3978);
and U5377 (N_5377,N_3595,N_3509);
or U5378 (N_5378,N_3202,N_4234);
nor U5379 (N_5379,N_3536,N_3735);
and U5380 (N_5380,N_4369,N_3334);
and U5381 (N_5381,N_4177,N_4158);
nor U5382 (N_5382,N_4438,N_3557);
nor U5383 (N_5383,N_3617,N_3330);
xor U5384 (N_5384,N_4291,N_3652);
and U5385 (N_5385,N_4052,N_3292);
nor U5386 (N_5386,N_3079,N_4034);
nor U5387 (N_5387,N_4490,N_3317);
nor U5388 (N_5388,N_4354,N_3303);
or U5389 (N_5389,N_3917,N_3869);
and U5390 (N_5390,N_3446,N_3983);
nand U5391 (N_5391,N_3972,N_3906);
nand U5392 (N_5392,N_3752,N_3538);
nand U5393 (N_5393,N_3578,N_3911);
or U5394 (N_5394,N_3726,N_3960);
nor U5395 (N_5395,N_3540,N_4079);
or U5396 (N_5396,N_3489,N_3408);
nand U5397 (N_5397,N_3012,N_3549);
nor U5398 (N_5398,N_3334,N_4039);
or U5399 (N_5399,N_3227,N_4442);
nand U5400 (N_5400,N_3191,N_4234);
nor U5401 (N_5401,N_4144,N_3605);
nor U5402 (N_5402,N_3168,N_4438);
and U5403 (N_5403,N_3397,N_4096);
nand U5404 (N_5404,N_3775,N_3915);
nor U5405 (N_5405,N_3512,N_4379);
nand U5406 (N_5406,N_4396,N_3797);
or U5407 (N_5407,N_3121,N_3038);
nand U5408 (N_5408,N_3728,N_3202);
nand U5409 (N_5409,N_4348,N_4273);
and U5410 (N_5410,N_3026,N_4019);
or U5411 (N_5411,N_3657,N_3357);
and U5412 (N_5412,N_3523,N_3902);
or U5413 (N_5413,N_3372,N_4201);
or U5414 (N_5414,N_4415,N_3144);
nor U5415 (N_5415,N_3417,N_3729);
nor U5416 (N_5416,N_3285,N_4102);
xnor U5417 (N_5417,N_3049,N_4499);
nand U5418 (N_5418,N_3153,N_3402);
or U5419 (N_5419,N_4320,N_3026);
and U5420 (N_5420,N_3166,N_3722);
or U5421 (N_5421,N_4270,N_3468);
nor U5422 (N_5422,N_3868,N_3493);
nand U5423 (N_5423,N_3631,N_3536);
nor U5424 (N_5424,N_3028,N_3766);
nor U5425 (N_5425,N_4438,N_3905);
xor U5426 (N_5426,N_3129,N_3114);
or U5427 (N_5427,N_3425,N_3375);
xnor U5428 (N_5428,N_3032,N_3153);
nand U5429 (N_5429,N_3316,N_3838);
and U5430 (N_5430,N_4143,N_3629);
xnor U5431 (N_5431,N_4041,N_3317);
nor U5432 (N_5432,N_3954,N_4270);
nor U5433 (N_5433,N_3564,N_4312);
nand U5434 (N_5434,N_3650,N_3505);
and U5435 (N_5435,N_3394,N_3908);
nor U5436 (N_5436,N_3666,N_3978);
nor U5437 (N_5437,N_3089,N_3735);
xor U5438 (N_5438,N_3532,N_3633);
nor U5439 (N_5439,N_4122,N_4155);
nor U5440 (N_5440,N_3281,N_3129);
xor U5441 (N_5441,N_3924,N_4488);
nor U5442 (N_5442,N_3576,N_4167);
xnor U5443 (N_5443,N_4336,N_3548);
or U5444 (N_5444,N_3220,N_3929);
and U5445 (N_5445,N_4219,N_3856);
and U5446 (N_5446,N_4333,N_4058);
or U5447 (N_5447,N_4006,N_3127);
xnor U5448 (N_5448,N_3839,N_3796);
and U5449 (N_5449,N_4395,N_4011);
and U5450 (N_5450,N_4067,N_3221);
or U5451 (N_5451,N_3298,N_3362);
or U5452 (N_5452,N_4248,N_4332);
and U5453 (N_5453,N_4131,N_3547);
nor U5454 (N_5454,N_3569,N_3677);
nor U5455 (N_5455,N_4017,N_3225);
nand U5456 (N_5456,N_3902,N_4322);
nor U5457 (N_5457,N_4089,N_3655);
or U5458 (N_5458,N_3988,N_4050);
nand U5459 (N_5459,N_3959,N_3899);
nand U5460 (N_5460,N_3156,N_3725);
and U5461 (N_5461,N_3126,N_4462);
nor U5462 (N_5462,N_3145,N_4396);
and U5463 (N_5463,N_4148,N_3948);
nor U5464 (N_5464,N_3271,N_3816);
and U5465 (N_5465,N_3223,N_3560);
nand U5466 (N_5466,N_4393,N_3340);
nor U5467 (N_5467,N_3797,N_3826);
and U5468 (N_5468,N_3755,N_4130);
and U5469 (N_5469,N_3610,N_3779);
or U5470 (N_5470,N_3722,N_3441);
nand U5471 (N_5471,N_3512,N_3784);
or U5472 (N_5472,N_3215,N_3498);
and U5473 (N_5473,N_4479,N_3212);
or U5474 (N_5474,N_3719,N_4495);
or U5475 (N_5475,N_3366,N_4045);
nand U5476 (N_5476,N_3747,N_3199);
nor U5477 (N_5477,N_3655,N_3458);
or U5478 (N_5478,N_3526,N_3159);
xnor U5479 (N_5479,N_3052,N_3693);
nor U5480 (N_5480,N_4003,N_4076);
nand U5481 (N_5481,N_3579,N_4151);
and U5482 (N_5482,N_4179,N_4269);
xor U5483 (N_5483,N_4032,N_4241);
or U5484 (N_5484,N_3367,N_4454);
nor U5485 (N_5485,N_3094,N_4413);
nand U5486 (N_5486,N_4474,N_3638);
nor U5487 (N_5487,N_3669,N_3366);
or U5488 (N_5488,N_4115,N_3113);
nand U5489 (N_5489,N_4028,N_4432);
or U5490 (N_5490,N_3517,N_4402);
or U5491 (N_5491,N_3798,N_3103);
or U5492 (N_5492,N_4311,N_3318);
and U5493 (N_5493,N_4257,N_3314);
or U5494 (N_5494,N_3570,N_4498);
or U5495 (N_5495,N_4077,N_3788);
nand U5496 (N_5496,N_3688,N_3319);
nand U5497 (N_5497,N_4232,N_3010);
or U5498 (N_5498,N_4439,N_3806);
xnor U5499 (N_5499,N_3363,N_3347);
nand U5500 (N_5500,N_4476,N_4178);
nor U5501 (N_5501,N_3536,N_3434);
and U5502 (N_5502,N_3504,N_3017);
or U5503 (N_5503,N_4204,N_4168);
nor U5504 (N_5504,N_4289,N_3328);
xor U5505 (N_5505,N_3575,N_4426);
and U5506 (N_5506,N_4142,N_4033);
or U5507 (N_5507,N_4222,N_4190);
nand U5508 (N_5508,N_4232,N_3695);
or U5509 (N_5509,N_3551,N_4198);
and U5510 (N_5510,N_3868,N_3762);
nand U5511 (N_5511,N_3180,N_4330);
or U5512 (N_5512,N_4093,N_3036);
nand U5513 (N_5513,N_3093,N_3331);
nand U5514 (N_5514,N_4424,N_3849);
nand U5515 (N_5515,N_3546,N_4225);
or U5516 (N_5516,N_3657,N_3835);
xor U5517 (N_5517,N_3502,N_4380);
xnor U5518 (N_5518,N_3998,N_3838);
nor U5519 (N_5519,N_4325,N_3585);
nor U5520 (N_5520,N_3551,N_3301);
xnor U5521 (N_5521,N_3547,N_4362);
and U5522 (N_5522,N_3437,N_3243);
nor U5523 (N_5523,N_3488,N_3561);
and U5524 (N_5524,N_4319,N_3989);
or U5525 (N_5525,N_3845,N_3168);
or U5526 (N_5526,N_3000,N_3211);
and U5527 (N_5527,N_4018,N_4193);
nand U5528 (N_5528,N_4203,N_3722);
nor U5529 (N_5529,N_3866,N_4233);
xnor U5530 (N_5530,N_3880,N_4279);
or U5531 (N_5531,N_3028,N_3824);
nor U5532 (N_5532,N_3085,N_3234);
xor U5533 (N_5533,N_4265,N_3257);
or U5534 (N_5534,N_4177,N_4009);
or U5535 (N_5535,N_3580,N_3558);
nor U5536 (N_5536,N_3121,N_3703);
nor U5537 (N_5537,N_3560,N_3117);
and U5538 (N_5538,N_3612,N_3868);
or U5539 (N_5539,N_4239,N_4056);
and U5540 (N_5540,N_3886,N_4411);
nand U5541 (N_5541,N_3135,N_3686);
and U5542 (N_5542,N_3779,N_3407);
or U5543 (N_5543,N_3827,N_3922);
or U5544 (N_5544,N_3493,N_3590);
or U5545 (N_5545,N_4196,N_3337);
nor U5546 (N_5546,N_3480,N_4048);
nand U5547 (N_5547,N_3817,N_3175);
or U5548 (N_5548,N_3267,N_3683);
nor U5549 (N_5549,N_3277,N_3470);
nor U5550 (N_5550,N_3077,N_3681);
nand U5551 (N_5551,N_3544,N_3257);
and U5552 (N_5552,N_3779,N_4284);
nand U5553 (N_5553,N_3082,N_3563);
nor U5554 (N_5554,N_4404,N_3475);
nand U5555 (N_5555,N_3270,N_4169);
xor U5556 (N_5556,N_3898,N_4055);
or U5557 (N_5557,N_3714,N_3682);
xnor U5558 (N_5558,N_4359,N_3316);
nand U5559 (N_5559,N_3330,N_3202);
nand U5560 (N_5560,N_3365,N_4260);
nor U5561 (N_5561,N_4063,N_3975);
nor U5562 (N_5562,N_3133,N_3508);
and U5563 (N_5563,N_3816,N_3182);
nor U5564 (N_5564,N_4039,N_4155);
nor U5565 (N_5565,N_3441,N_3970);
nand U5566 (N_5566,N_3355,N_4159);
and U5567 (N_5567,N_4434,N_3295);
or U5568 (N_5568,N_3467,N_3521);
or U5569 (N_5569,N_3789,N_3355);
and U5570 (N_5570,N_3406,N_4294);
and U5571 (N_5571,N_3173,N_3837);
nor U5572 (N_5572,N_4222,N_3071);
or U5573 (N_5573,N_4174,N_3808);
or U5574 (N_5574,N_3148,N_4132);
or U5575 (N_5575,N_4080,N_3380);
and U5576 (N_5576,N_3968,N_3067);
nand U5577 (N_5577,N_3614,N_3101);
nand U5578 (N_5578,N_3206,N_3848);
nand U5579 (N_5579,N_4364,N_3380);
xnor U5580 (N_5580,N_3623,N_4312);
nand U5581 (N_5581,N_3261,N_3746);
and U5582 (N_5582,N_3847,N_3572);
or U5583 (N_5583,N_3964,N_3480);
xnor U5584 (N_5584,N_3925,N_4103);
and U5585 (N_5585,N_4167,N_4239);
nor U5586 (N_5586,N_3837,N_3867);
nand U5587 (N_5587,N_3675,N_3773);
nand U5588 (N_5588,N_3067,N_4312);
nand U5589 (N_5589,N_3641,N_3695);
and U5590 (N_5590,N_4105,N_3399);
or U5591 (N_5591,N_3179,N_3483);
nor U5592 (N_5592,N_4047,N_4212);
xnor U5593 (N_5593,N_3868,N_4089);
and U5594 (N_5594,N_3788,N_4001);
and U5595 (N_5595,N_4298,N_4084);
nand U5596 (N_5596,N_3057,N_4052);
nand U5597 (N_5597,N_4431,N_4043);
nand U5598 (N_5598,N_3471,N_3279);
and U5599 (N_5599,N_3729,N_4195);
xnor U5600 (N_5600,N_3773,N_3419);
or U5601 (N_5601,N_3230,N_4097);
xnor U5602 (N_5602,N_3414,N_3432);
or U5603 (N_5603,N_4077,N_3166);
or U5604 (N_5604,N_4178,N_3311);
and U5605 (N_5605,N_3424,N_4248);
and U5606 (N_5606,N_3401,N_3828);
xnor U5607 (N_5607,N_4172,N_3757);
nand U5608 (N_5608,N_4324,N_3036);
and U5609 (N_5609,N_3252,N_3266);
xnor U5610 (N_5610,N_3668,N_3244);
or U5611 (N_5611,N_3697,N_4328);
and U5612 (N_5612,N_4063,N_4234);
or U5613 (N_5613,N_3354,N_4174);
nand U5614 (N_5614,N_3207,N_3608);
or U5615 (N_5615,N_3675,N_3210);
nand U5616 (N_5616,N_4281,N_3723);
and U5617 (N_5617,N_3245,N_4034);
nor U5618 (N_5618,N_3342,N_4302);
nand U5619 (N_5619,N_4016,N_4452);
nand U5620 (N_5620,N_3787,N_4239);
nand U5621 (N_5621,N_3839,N_3591);
nand U5622 (N_5622,N_4430,N_3754);
nand U5623 (N_5623,N_4304,N_3335);
xnor U5624 (N_5624,N_3912,N_3287);
or U5625 (N_5625,N_3830,N_3261);
and U5626 (N_5626,N_4113,N_3263);
and U5627 (N_5627,N_3455,N_3804);
and U5628 (N_5628,N_3098,N_3255);
nand U5629 (N_5629,N_3203,N_3453);
and U5630 (N_5630,N_3613,N_3517);
and U5631 (N_5631,N_3246,N_3414);
xor U5632 (N_5632,N_3374,N_3858);
nor U5633 (N_5633,N_4306,N_3875);
nand U5634 (N_5634,N_3025,N_3246);
or U5635 (N_5635,N_3122,N_3246);
or U5636 (N_5636,N_3457,N_4305);
nand U5637 (N_5637,N_4364,N_4427);
nand U5638 (N_5638,N_4182,N_3908);
and U5639 (N_5639,N_4387,N_4187);
and U5640 (N_5640,N_4484,N_4416);
xnor U5641 (N_5641,N_3582,N_3539);
nand U5642 (N_5642,N_4487,N_4043);
nor U5643 (N_5643,N_4401,N_3683);
and U5644 (N_5644,N_3583,N_4232);
or U5645 (N_5645,N_4399,N_4088);
nor U5646 (N_5646,N_4428,N_4132);
and U5647 (N_5647,N_3106,N_3379);
xor U5648 (N_5648,N_3563,N_3544);
or U5649 (N_5649,N_3371,N_4477);
nand U5650 (N_5650,N_3472,N_3422);
nor U5651 (N_5651,N_3921,N_3460);
nor U5652 (N_5652,N_3227,N_4053);
nand U5653 (N_5653,N_3713,N_4385);
xor U5654 (N_5654,N_3861,N_4057);
nand U5655 (N_5655,N_3555,N_4201);
nand U5656 (N_5656,N_4350,N_3330);
or U5657 (N_5657,N_4075,N_4255);
xnor U5658 (N_5658,N_3549,N_4351);
and U5659 (N_5659,N_3299,N_3938);
nor U5660 (N_5660,N_3594,N_3980);
and U5661 (N_5661,N_3041,N_3574);
nor U5662 (N_5662,N_4323,N_3347);
and U5663 (N_5663,N_3612,N_3145);
or U5664 (N_5664,N_3535,N_3481);
nand U5665 (N_5665,N_4132,N_3050);
nor U5666 (N_5666,N_3404,N_3477);
nand U5667 (N_5667,N_4476,N_4085);
nor U5668 (N_5668,N_4258,N_3678);
and U5669 (N_5669,N_3921,N_3186);
xor U5670 (N_5670,N_4107,N_4067);
and U5671 (N_5671,N_3373,N_3801);
nand U5672 (N_5672,N_3037,N_4464);
nor U5673 (N_5673,N_3743,N_3335);
nand U5674 (N_5674,N_4415,N_4196);
or U5675 (N_5675,N_4253,N_3031);
and U5676 (N_5676,N_3600,N_3793);
or U5677 (N_5677,N_3695,N_3541);
or U5678 (N_5678,N_4438,N_3824);
nand U5679 (N_5679,N_3532,N_3678);
nor U5680 (N_5680,N_3397,N_3149);
nand U5681 (N_5681,N_3116,N_3135);
or U5682 (N_5682,N_3954,N_3527);
and U5683 (N_5683,N_4298,N_3321);
or U5684 (N_5684,N_3045,N_3126);
xor U5685 (N_5685,N_3555,N_3945);
nand U5686 (N_5686,N_4073,N_4248);
nor U5687 (N_5687,N_3607,N_3491);
or U5688 (N_5688,N_4252,N_4235);
nand U5689 (N_5689,N_3071,N_4191);
xor U5690 (N_5690,N_4270,N_3507);
nor U5691 (N_5691,N_3068,N_4434);
nand U5692 (N_5692,N_3019,N_3201);
or U5693 (N_5693,N_3336,N_3142);
and U5694 (N_5694,N_4243,N_4401);
nand U5695 (N_5695,N_3542,N_4041);
xor U5696 (N_5696,N_4095,N_4423);
nand U5697 (N_5697,N_4049,N_4264);
or U5698 (N_5698,N_3866,N_4250);
nor U5699 (N_5699,N_3517,N_3578);
or U5700 (N_5700,N_3191,N_3980);
xnor U5701 (N_5701,N_3947,N_3712);
and U5702 (N_5702,N_3987,N_4226);
or U5703 (N_5703,N_4169,N_4040);
nand U5704 (N_5704,N_4339,N_3028);
xnor U5705 (N_5705,N_4336,N_3106);
nand U5706 (N_5706,N_3847,N_4250);
nor U5707 (N_5707,N_3703,N_4314);
nor U5708 (N_5708,N_4180,N_4088);
and U5709 (N_5709,N_3454,N_3255);
nand U5710 (N_5710,N_3271,N_3714);
nor U5711 (N_5711,N_4381,N_3784);
nand U5712 (N_5712,N_4397,N_4141);
and U5713 (N_5713,N_3014,N_3510);
nor U5714 (N_5714,N_4384,N_4048);
xnor U5715 (N_5715,N_3089,N_3771);
xnor U5716 (N_5716,N_4418,N_3594);
and U5717 (N_5717,N_3427,N_3405);
nor U5718 (N_5718,N_3882,N_3160);
nor U5719 (N_5719,N_3898,N_3161);
or U5720 (N_5720,N_3366,N_3854);
and U5721 (N_5721,N_4069,N_3320);
and U5722 (N_5722,N_3425,N_3094);
nand U5723 (N_5723,N_3902,N_3427);
nor U5724 (N_5724,N_3511,N_4106);
or U5725 (N_5725,N_4498,N_3421);
or U5726 (N_5726,N_4071,N_3456);
or U5727 (N_5727,N_3290,N_3977);
nand U5728 (N_5728,N_3781,N_4275);
or U5729 (N_5729,N_4392,N_3245);
nor U5730 (N_5730,N_4238,N_4002);
and U5731 (N_5731,N_3379,N_3476);
or U5732 (N_5732,N_3809,N_3923);
nor U5733 (N_5733,N_3981,N_3592);
nor U5734 (N_5734,N_3606,N_4289);
nor U5735 (N_5735,N_3539,N_3590);
nand U5736 (N_5736,N_4455,N_3241);
or U5737 (N_5737,N_4422,N_4269);
or U5738 (N_5738,N_3916,N_3798);
nand U5739 (N_5739,N_3730,N_3591);
nand U5740 (N_5740,N_4296,N_3453);
nor U5741 (N_5741,N_3933,N_4018);
or U5742 (N_5742,N_3213,N_3605);
nand U5743 (N_5743,N_3152,N_3727);
and U5744 (N_5744,N_3542,N_3870);
nor U5745 (N_5745,N_4185,N_4121);
nand U5746 (N_5746,N_4197,N_4172);
or U5747 (N_5747,N_3723,N_4031);
or U5748 (N_5748,N_3522,N_3357);
nor U5749 (N_5749,N_3592,N_3073);
or U5750 (N_5750,N_3502,N_4470);
or U5751 (N_5751,N_4049,N_3646);
xor U5752 (N_5752,N_4407,N_3922);
and U5753 (N_5753,N_4332,N_3792);
or U5754 (N_5754,N_3824,N_4215);
nor U5755 (N_5755,N_4336,N_3165);
nor U5756 (N_5756,N_4189,N_3757);
xnor U5757 (N_5757,N_3654,N_3787);
nand U5758 (N_5758,N_3555,N_3140);
and U5759 (N_5759,N_4258,N_3216);
nand U5760 (N_5760,N_3336,N_3180);
nor U5761 (N_5761,N_4140,N_3040);
and U5762 (N_5762,N_3215,N_3043);
xor U5763 (N_5763,N_3835,N_3878);
or U5764 (N_5764,N_4425,N_3827);
nand U5765 (N_5765,N_3337,N_4088);
or U5766 (N_5766,N_4019,N_3961);
or U5767 (N_5767,N_3682,N_4150);
and U5768 (N_5768,N_3966,N_4394);
or U5769 (N_5769,N_4439,N_3183);
nand U5770 (N_5770,N_4372,N_3920);
and U5771 (N_5771,N_4388,N_4079);
nor U5772 (N_5772,N_3335,N_4293);
nand U5773 (N_5773,N_3795,N_3190);
nor U5774 (N_5774,N_3176,N_3634);
or U5775 (N_5775,N_4108,N_3122);
and U5776 (N_5776,N_3333,N_3063);
nor U5777 (N_5777,N_4413,N_3985);
nand U5778 (N_5778,N_4062,N_4210);
and U5779 (N_5779,N_3753,N_3074);
or U5780 (N_5780,N_4038,N_3937);
or U5781 (N_5781,N_4277,N_3856);
or U5782 (N_5782,N_4093,N_4406);
nand U5783 (N_5783,N_4173,N_3552);
and U5784 (N_5784,N_3709,N_3740);
nand U5785 (N_5785,N_3176,N_3594);
nand U5786 (N_5786,N_3441,N_4043);
or U5787 (N_5787,N_3055,N_3424);
nand U5788 (N_5788,N_4063,N_3311);
or U5789 (N_5789,N_4060,N_3529);
nor U5790 (N_5790,N_4491,N_3024);
or U5791 (N_5791,N_3006,N_4076);
nand U5792 (N_5792,N_3905,N_3780);
xnor U5793 (N_5793,N_3646,N_4293);
or U5794 (N_5794,N_3557,N_3342);
nor U5795 (N_5795,N_3017,N_3473);
or U5796 (N_5796,N_3941,N_4011);
or U5797 (N_5797,N_3617,N_3118);
or U5798 (N_5798,N_3141,N_3667);
or U5799 (N_5799,N_3822,N_4280);
and U5800 (N_5800,N_3258,N_4198);
or U5801 (N_5801,N_3352,N_3237);
nor U5802 (N_5802,N_3431,N_4203);
or U5803 (N_5803,N_3897,N_3821);
nand U5804 (N_5804,N_4102,N_4383);
xor U5805 (N_5805,N_4494,N_4155);
nand U5806 (N_5806,N_3056,N_4137);
or U5807 (N_5807,N_3641,N_3063);
and U5808 (N_5808,N_3369,N_3713);
xnor U5809 (N_5809,N_3593,N_4493);
or U5810 (N_5810,N_4199,N_4403);
or U5811 (N_5811,N_4017,N_4146);
nor U5812 (N_5812,N_3552,N_3918);
nand U5813 (N_5813,N_3436,N_3301);
nand U5814 (N_5814,N_3698,N_4315);
and U5815 (N_5815,N_4481,N_3052);
nor U5816 (N_5816,N_4038,N_4021);
or U5817 (N_5817,N_3090,N_4477);
or U5818 (N_5818,N_4356,N_3505);
xor U5819 (N_5819,N_3301,N_3994);
and U5820 (N_5820,N_4120,N_3732);
and U5821 (N_5821,N_3901,N_3196);
or U5822 (N_5822,N_3676,N_4222);
nor U5823 (N_5823,N_3721,N_3917);
nor U5824 (N_5824,N_3062,N_3037);
nor U5825 (N_5825,N_3549,N_3837);
nand U5826 (N_5826,N_3821,N_3079);
or U5827 (N_5827,N_3631,N_4017);
and U5828 (N_5828,N_4455,N_4303);
and U5829 (N_5829,N_3266,N_4115);
nand U5830 (N_5830,N_4352,N_4156);
and U5831 (N_5831,N_3742,N_3856);
xnor U5832 (N_5832,N_3759,N_3313);
or U5833 (N_5833,N_4260,N_3102);
and U5834 (N_5834,N_3836,N_3578);
and U5835 (N_5835,N_3978,N_3604);
nand U5836 (N_5836,N_4451,N_3956);
nor U5837 (N_5837,N_3819,N_3890);
and U5838 (N_5838,N_3950,N_3005);
nand U5839 (N_5839,N_4055,N_3475);
and U5840 (N_5840,N_3898,N_4413);
and U5841 (N_5841,N_3548,N_3447);
or U5842 (N_5842,N_3742,N_3941);
nor U5843 (N_5843,N_3761,N_3404);
xor U5844 (N_5844,N_3021,N_3273);
nand U5845 (N_5845,N_3408,N_3202);
nand U5846 (N_5846,N_3589,N_3368);
nor U5847 (N_5847,N_4258,N_4463);
nand U5848 (N_5848,N_3189,N_4467);
and U5849 (N_5849,N_3690,N_4149);
nand U5850 (N_5850,N_3813,N_4474);
and U5851 (N_5851,N_3961,N_3413);
xor U5852 (N_5852,N_3515,N_4112);
and U5853 (N_5853,N_4230,N_3955);
nor U5854 (N_5854,N_3549,N_3701);
and U5855 (N_5855,N_3546,N_3176);
and U5856 (N_5856,N_4092,N_3090);
nor U5857 (N_5857,N_3086,N_4362);
and U5858 (N_5858,N_3852,N_3666);
and U5859 (N_5859,N_3821,N_4437);
and U5860 (N_5860,N_4175,N_3474);
nor U5861 (N_5861,N_3393,N_3407);
nand U5862 (N_5862,N_3588,N_3104);
nor U5863 (N_5863,N_4414,N_4340);
nand U5864 (N_5864,N_3508,N_3883);
nand U5865 (N_5865,N_3595,N_3738);
or U5866 (N_5866,N_4191,N_4103);
nand U5867 (N_5867,N_4193,N_3171);
xnor U5868 (N_5868,N_3467,N_3374);
nand U5869 (N_5869,N_4111,N_3192);
nand U5870 (N_5870,N_4210,N_3458);
or U5871 (N_5871,N_3864,N_4022);
and U5872 (N_5872,N_3363,N_3413);
or U5873 (N_5873,N_4150,N_4416);
or U5874 (N_5874,N_3070,N_3238);
xor U5875 (N_5875,N_3942,N_3236);
nand U5876 (N_5876,N_3783,N_3577);
or U5877 (N_5877,N_3329,N_3273);
nand U5878 (N_5878,N_3824,N_4388);
and U5879 (N_5879,N_3457,N_3222);
nor U5880 (N_5880,N_4064,N_3821);
and U5881 (N_5881,N_3275,N_3478);
or U5882 (N_5882,N_3988,N_3333);
xor U5883 (N_5883,N_3539,N_4373);
xnor U5884 (N_5884,N_3855,N_3427);
or U5885 (N_5885,N_3646,N_3973);
nor U5886 (N_5886,N_3794,N_3564);
and U5887 (N_5887,N_3638,N_3574);
nand U5888 (N_5888,N_3419,N_3733);
nand U5889 (N_5889,N_3610,N_4421);
or U5890 (N_5890,N_3264,N_4459);
nand U5891 (N_5891,N_3127,N_3073);
nand U5892 (N_5892,N_3868,N_3792);
nor U5893 (N_5893,N_3859,N_4232);
and U5894 (N_5894,N_4306,N_3220);
nand U5895 (N_5895,N_3631,N_4421);
or U5896 (N_5896,N_3115,N_3000);
or U5897 (N_5897,N_3852,N_4025);
xnor U5898 (N_5898,N_4013,N_4232);
and U5899 (N_5899,N_4181,N_4408);
nor U5900 (N_5900,N_3664,N_4217);
nor U5901 (N_5901,N_3824,N_4081);
nor U5902 (N_5902,N_3648,N_4345);
nor U5903 (N_5903,N_3217,N_3823);
nor U5904 (N_5904,N_3183,N_3608);
and U5905 (N_5905,N_4325,N_4335);
xnor U5906 (N_5906,N_3049,N_4342);
nand U5907 (N_5907,N_3706,N_3035);
nor U5908 (N_5908,N_4283,N_4270);
nor U5909 (N_5909,N_3777,N_3288);
xnor U5910 (N_5910,N_3491,N_3811);
or U5911 (N_5911,N_4184,N_3765);
nand U5912 (N_5912,N_4113,N_4482);
nand U5913 (N_5913,N_4458,N_4011);
and U5914 (N_5914,N_3551,N_3952);
nand U5915 (N_5915,N_4405,N_4073);
nand U5916 (N_5916,N_3335,N_4445);
and U5917 (N_5917,N_4419,N_4016);
and U5918 (N_5918,N_3055,N_4453);
or U5919 (N_5919,N_4365,N_3880);
xor U5920 (N_5920,N_3245,N_4263);
and U5921 (N_5921,N_3971,N_3669);
and U5922 (N_5922,N_3923,N_4179);
or U5923 (N_5923,N_4018,N_3536);
nor U5924 (N_5924,N_4245,N_3689);
or U5925 (N_5925,N_3312,N_4349);
and U5926 (N_5926,N_3478,N_3274);
xnor U5927 (N_5927,N_3600,N_4057);
and U5928 (N_5928,N_3734,N_4477);
or U5929 (N_5929,N_4131,N_3454);
and U5930 (N_5930,N_4084,N_4434);
or U5931 (N_5931,N_3521,N_4441);
nor U5932 (N_5932,N_3732,N_4182);
or U5933 (N_5933,N_3055,N_4021);
nor U5934 (N_5934,N_3269,N_3602);
or U5935 (N_5935,N_3709,N_4253);
nand U5936 (N_5936,N_3504,N_3662);
nand U5937 (N_5937,N_3903,N_3024);
xnor U5938 (N_5938,N_3563,N_3137);
or U5939 (N_5939,N_3097,N_4357);
nor U5940 (N_5940,N_3374,N_3320);
nor U5941 (N_5941,N_3654,N_3461);
nand U5942 (N_5942,N_3291,N_4123);
nand U5943 (N_5943,N_3228,N_3954);
nor U5944 (N_5944,N_3230,N_3242);
and U5945 (N_5945,N_3462,N_3318);
xnor U5946 (N_5946,N_3074,N_3739);
and U5947 (N_5947,N_3557,N_4131);
nor U5948 (N_5948,N_3595,N_3990);
nor U5949 (N_5949,N_3962,N_4427);
and U5950 (N_5950,N_4019,N_3249);
nand U5951 (N_5951,N_4117,N_3813);
nor U5952 (N_5952,N_3140,N_4418);
nor U5953 (N_5953,N_3821,N_4113);
nor U5954 (N_5954,N_3447,N_3618);
xor U5955 (N_5955,N_3604,N_3989);
and U5956 (N_5956,N_3815,N_3306);
nand U5957 (N_5957,N_3022,N_3719);
nand U5958 (N_5958,N_4131,N_3841);
nor U5959 (N_5959,N_3744,N_3329);
nand U5960 (N_5960,N_4069,N_3778);
nand U5961 (N_5961,N_3595,N_3793);
and U5962 (N_5962,N_3200,N_3835);
nand U5963 (N_5963,N_4351,N_3027);
xnor U5964 (N_5964,N_4087,N_3227);
and U5965 (N_5965,N_3863,N_3774);
and U5966 (N_5966,N_4260,N_3779);
nand U5967 (N_5967,N_3679,N_3133);
nand U5968 (N_5968,N_3782,N_4340);
and U5969 (N_5969,N_3850,N_3666);
nor U5970 (N_5970,N_4261,N_3756);
or U5971 (N_5971,N_3344,N_3841);
or U5972 (N_5972,N_3732,N_3274);
nand U5973 (N_5973,N_3470,N_4438);
and U5974 (N_5974,N_3090,N_4016);
xor U5975 (N_5975,N_3697,N_4446);
or U5976 (N_5976,N_3628,N_3456);
nor U5977 (N_5977,N_3188,N_4117);
nor U5978 (N_5978,N_3271,N_3583);
or U5979 (N_5979,N_3886,N_4102);
xnor U5980 (N_5980,N_3022,N_3826);
nand U5981 (N_5981,N_4077,N_3285);
nor U5982 (N_5982,N_3718,N_4309);
nor U5983 (N_5983,N_3204,N_4494);
xnor U5984 (N_5984,N_3212,N_3350);
nand U5985 (N_5985,N_3541,N_3582);
and U5986 (N_5986,N_3280,N_3986);
nor U5987 (N_5987,N_4154,N_3599);
and U5988 (N_5988,N_3760,N_3987);
nor U5989 (N_5989,N_4295,N_3374);
or U5990 (N_5990,N_3025,N_3220);
nand U5991 (N_5991,N_3859,N_3703);
or U5992 (N_5992,N_3933,N_3237);
nand U5993 (N_5993,N_3184,N_3607);
nor U5994 (N_5994,N_3542,N_4226);
xnor U5995 (N_5995,N_4091,N_3667);
nand U5996 (N_5996,N_3788,N_4063);
nor U5997 (N_5997,N_4128,N_3310);
or U5998 (N_5998,N_4347,N_3219);
nor U5999 (N_5999,N_3261,N_3345);
nor U6000 (N_6000,N_5793,N_4527);
or U6001 (N_6001,N_5926,N_5181);
and U6002 (N_6002,N_5459,N_5760);
nor U6003 (N_6003,N_4892,N_5269);
nor U6004 (N_6004,N_5057,N_5894);
nor U6005 (N_6005,N_5489,N_4961);
nand U6006 (N_6006,N_4612,N_5464);
nor U6007 (N_6007,N_5511,N_5712);
nor U6008 (N_6008,N_4954,N_5123);
nor U6009 (N_6009,N_5102,N_4721);
nand U6010 (N_6010,N_4918,N_5780);
or U6011 (N_6011,N_4907,N_5940);
and U6012 (N_6012,N_5659,N_5525);
nand U6013 (N_6013,N_4898,N_5412);
and U6014 (N_6014,N_4606,N_5627);
and U6015 (N_6015,N_5128,N_5152);
and U6016 (N_6016,N_5858,N_5770);
or U6017 (N_6017,N_4849,N_5556);
or U6018 (N_6018,N_4819,N_5893);
or U6019 (N_6019,N_5968,N_4882);
nor U6020 (N_6020,N_4590,N_5538);
or U6021 (N_6021,N_5141,N_4838);
nand U6022 (N_6022,N_5772,N_4618);
nand U6023 (N_6023,N_5837,N_5228);
nand U6024 (N_6024,N_4733,N_4862);
nand U6025 (N_6025,N_5138,N_5160);
and U6026 (N_6026,N_5104,N_5891);
nand U6027 (N_6027,N_5040,N_5761);
and U6028 (N_6028,N_4801,N_5775);
and U6029 (N_6029,N_4637,N_5618);
or U6030 (N_6030,N_4916,N_4641);
xnor U6031 (N_6031,N_5355,N_4750);
or U6032 (N_6032,N_5059,N_5285);
nand U6033 (N_6033,N_5653,N_5447);
nand U6034 (N_6034,N_5062,N_5897);
nand U6035 (N_6035,N_5192,N_4589);
or U6036 (N_6036,N_5290,N_5589);
nand U6037 (N_6037,N_5796,N_4682);
or U6038 (N_6038,N_4561,N_5453);
nor U6039 (N_6039,N_4663,N_4989);
and U6040 (N_6040,N_5949,N_5432);
or U6041 (N_6041,N_5963,N_5016);
nor U6042 (N_6042,N_5762,N_4760);
and U6043 (N_6043,N_5452,N_5711);
nor U6044 (N_6044,N_5764,N_4509);
and U6045 (N_6045,N_5222,N_5946);
and U6046 (N_6046,N_5261,N_4611);
and U6047 (N_6047,N_5737,N_4963);
nand U6048 (N_6048,N_4741,N_4924);
nor U6049 (N_6049,N_4577,N_4762);
or U6050 (N_6050,N_5882,N_4787);
nand U6051 (N_6051,N_4514,N_5942);
and U6052 (N_6052,N_4708,N_5503);
xor U6053 (N_6053,N_4523,N_4854);
xor U6054 (N_6054,N_5929,N_5568);
or U6055 (N_6055,N_5258,N_5672);
nand U6056 (N_6056,N_4973,N_4666);
nand U6057 (N_6057,N_5203,N_5451);
or U6058 (N_6058,N_4588,N_5133);
xor U6059 (N_6059,N_4568,N_5270);
xnor U6060 (N_6060,N_5778,N_5878);
and U6061 (N_6061,N_4883,N_4504);
nor U6062 (N_6062,N_5064,N_5082);
and U6063 (N_6063,N_4692,N_5231);
or U6064 (N_6064,N_5210,N_5395);
nand U6065 (N_6065,N_5925,N_5422);
nor U6066 (N_6066,N_4863,N_4518);
nand U6067 (N_6067,N_5041,N_5500);
xnor U6068 (N_6068,N_4915,N_5528);
xnor U6069 (N_6069,N_5721,N_5534);
and U6070 (N_6070,N_5508,N_5311);
nor U6071 (N_6071,N_5811,N_5972);
and U6072 (N_6072,N_4811,N_5300);
or U6073 (N_6073,N_5429,N_5874);
nand U6074 (N_6074,N_5235,N_4749);
or U6075 (N_6075,N_5971,N_5936);
and U6076 (N_6076,N_4695,N_5822);
and U6077 (N_6077,N_4541,N_5901);
or U6078 (N_6078,N_5092,N_4667);
nand U6079 (N_6079,N_5410,N_4809);
nand U6080 (N_6080,N_5933,N_4713);
xor U6081 (N_6081,N_5714,N_5176);
and U6082 (N_6082,N_5177,N_5973);
nor U6083 (N_6083,N_4903,N_5073);
or U6084 (N_6084,N_5388,N_5582);
or U6085 (N_6085,N_5099,N_5666);
nor U6086 (N_6086,N_5595,N_4922);
nand U6087 (N_6087,N_5403,N_5875);
nor U6088 (N_6088,N_4554,N_4745);
and U6089 (N_6089,N_5912,N_4634);
nand U6090 (N_6090,N_5649,N_5739);
nand U6091 (N_6091,N_5325,N_5785);
nor U6092 (N_6092,N_5143,N_5517);
nor U6093 (N_6093,N_4813,N_5080);
or U6094 (N_6094,N_5724,N_4572);
nor U6095 (N_6095,N_5472,N_5363);
nor U6096 (N_6096,N_5314,N_5637);
nand U6097 (N_6097,N_5864,N_5977);
or U6098 (N_6098,N_5431,N_4619);
nor U6099 (N_6099,N_5510,N_4607);
nor U6100 (N_6100,N_4912,N_4670);
nor U6101 (N_6101,N_4624,N_5928);
xnor U6102 (N_6102,N_4983,N_4727);
nor U6103 (N_6103,N_5624,N_4691);
and U6104 (N_6104,N_5906,N_4786);
nor U6105 (N_6105,N_4650,N_4818);
nand U6106 (N_6106,N_4761,N_5107);
or U6107 (N_6107,N_4816,N_5809);
and U6108 (N_6108,N_5899,N_4753);
and U6109 (N_6109,N_4859,N_5297);
xnor U6110 (N_6110,N_5254,N_5846);
nand U6111 (N_6111,N_4742,N_5163);
nor U6112 (N_6112,N_5246,N_5162);
nor U6113 (N_6113,N_4976,N_5602);
nand U6114 (N_6114,N_5634,N_5910);
nor U6115 (N_6115,N_4709,N_4850);
nand U6116 (N_6116,N_5576,N_5540);
and U6117 (N_6117,N_5257,N_5207);
nand U6118 (N_6118,N_5543,N_4779);
or U6119 (N_6119,N_5260,N_5629);
nor U6120 (N_6120,N_4841,N_5838);
and U6121 (N_6121,N_5515,N_4793);
nand U6122 (N_6122,N_5371,N_5156);
and U6123 (N_6123,N_5449,N_5026);
and U6124 (N_6124,N_4759,N_4946);
nor U6125 (N_6125,N_5049,N_5168);
or U6126 (N_6126,N_4703,N_5698);
and U6127 (N_6127,N_4757,N_5684);
xnor U6128 (N_6128,N_5750,N_4716);
nor U6129 (N_6129,N_5075,N_5250);
nor U6130 (N_6130,N_4808,N_5524);
nor U6131 (N_6131,N_5930,N_4605);
nor U6132 (N_6132,N_5504,N_5896);
or U6133 (N_6133,N_5658,N_5333);
nor U6134 (N_6134,N_5433,N_4675);
xor U6135 (N_6135,N_4914,N_5571);
nor U6136 (N_6136,N_5272,N_4890);
nor U6137 (N_6137,N_5743,N_5917);
or U6138 (N_6138,N_4913,N_5173);
nand U6139 (N_6139,N_5436,N_4604);
xnor U6140 (N_6140,N_5052,N_4580);
or U6141 (N_6141,N_5200,N_5286);
nand U6142 (N_6142,N_5498,N_5547);
nand U6143 (N_6143,N_4584,N_4955);
nand U6144 (N_6144,N_5889,N_4705);
and U6145 (N_6145,N_5587,N_5063);
nor U6146 (N_6146,N_5601,N_5979);
nand U6147 (N_6147,N_4598,N_5639);
or U6148 (N_6148,N_5310,N_5387);
or U6149 (N_6149,N_5526,N_4535);
and U6150 (N_6150,N_4943,N_5321);
or U6151 (N_6151,N_5004,N_4851);
xor U6152 (N_6152,N_5264,N_5347);
nand U6153 (N_6153,N_5651,N_5931);
or U6154 (N_6154,N_5379,N_4647);
nand U6155 (N_6155,N_5784,N_4755);
nand U6156 (N_6156,N_5315,N_5130);
nand U6157 (N_6157,N_4586,N_5189);
and U6158 (N_6158,N_5172,N_5011);
nand U6159 (N_6159,N_5742,N_5167);
nor U6160 (N_6160,N_5663,N_4774);
or U6161 (N_6161,N_5442,N_5271);
and U6162 (N_6162,N_4627,N_5749);
or U6163 (N_6163,N_5677,N_5370);
or U6164 (N_6164,N_4575,N_5990);
or U6165 (N_6165,N_5487,N_4904);
nand U6166 (N_6166,N_5343,N_4860);
nor U6167 (N_6167,N_5044,N_5094);
and U6168 (N_6168,N_5396,N_5213);
nor U6169 (N_6169,N_5497,N_5032);
nor U6170 (N_6170,N_5390,N_5118);
nand U6171 (N_6171,N_5126,N_5042);
nor U6172 (N_6172,N_5230,N_5887);
or U6173 (N_6173,N_5787,N_4764);
nor U6174 (N_6174,N_5090,N_5050);
nand U6175 (N_6175,N_4694,N_4763);
or U6176 (N_6176,N_4521,N_4872);
nand U6177 (N_6177,N_5056,N_5017);
and U6178 (N_6178,N_5252,N_5998);
nand U6179 (N_6179,N_5021,N_5707);
and U6180 (N_6180,N_4526,N_4971);
xnor U6181 (N_6181,N_5117,N_4563);
nand U6182 (N_6182,N_4965,N_5259);
or U6183 (N_6183,N_5071,N_4843);
and U6184 (N_6184,N_4696,N_5440);
or U6185 (N_6185,N_5648,N_5765);
nand U6186 (N_6186,N_5546,N_5733);
nand U6187 (N_6187,N_4977,N_5855);
nor U6188 (N_6188,N_5923,N_4567);
and U6189 (N_6189,N_5754,N_5608);
xor U6190 (N_6190,N_5895,N_5706);
nor U6191 (N_6191,N_5959,N_5611);
or U6192 (N_6192,N_5372,N_4926);
nand U6193 (N_6193,N_5996,N_5782);
nor U6194 (N_6194,N_4969,N_5091);
or U6195 (N_6195,N_5043,N_5243);
or U6196 (N_6196,N_5598,N_5329);
or U6197 (N_6197,N_5575,N_5614);
or U6198 (N_6198,N_4592,N_5225);
nor U6199 (N_6199,N_5084,N_4622);
or U6200 (N_6200,N_5872,N_5559);
nor U6201 (N_6201,N_5305,N_5730);
and U6202 (N_6202,N_5288,N_4780);
xnor U6203 (N_6203,N_5475,N_5430);
nor U6204 (N_6204,N_4923,N_4729);
or U6205 (N_6205,N_5353,N_4669);
xor U6206 (N_6206,N_5951,N_5450);
or U6207 (N_6207,N_5691,N_4942);
and U6208 (N_6208,N_4751,N_5514);
or U6209 (N_6209,N_4783,N_5037);
nor U6210 (N_6210,N_5384,N_4905);
or U6211 (N_6211,N_4778,N_4972);
nand U6212 (N_6212,N_4505,N_5253);
and U6213 (N_6213,N_5954,N_5217);
xnor U6214 (N_6214,N_5078,N_5952);
nand U6215 (N_6215,N_5086,N_5561);
xnor U6216 (N_6216,N_4995,N_5284);
nor U6217 (N_6217,N_4502,N_4875);
xnor U6218 (N_6218,N_5718,N_5600);
nand U6219 (N_6219,N_4700,N_4834);
or U6220 (N_6220,N_5402,N_5628);
nor U6221 (N_6221,N_5696,N_4658);
or U6222 (N_6222,N_5960,N_5014);
or U6223 (N_6223,N_5890,N_5345);
or U6224 (N_6224,N_4654,N_4925);
nor U6225 (N_6225,N_5067,N_5365);
nor U6226 (N_6226,N_5581,N_4992);
or U6227 (N_6227,N_4948,N_5974);
nor U6228 (N_6228,N_5808,N_5194);
nand U6229 (N_6229,N_4996,N_4840);
or U6230 (N_6230,N_4827,N_4744);
nand U6231 (N_6231,N_5299,N_5638);
xor U6232 (N_6232,N_5792,N_5913);
nand U6233 (N_6233,N_4579,N_5407);
or U6234 (N_6234,N_5401,N_4506);
nand U6235 (N_6235,N_5630,N_5939);
and U6236 (N_6236,N_5751,N_4656);
or U6237 (N_6237,N_5334,N_5380);
nor U6238 (N_6238,N_4994,N_4551);
or U6239 (N_6239,N_4833,N_5135);
and U6240 (N_6240,N_5512,N_5723);
or U6241 (N_6241,N_5220,N_5495);
nand U6242 (N_6242,N_4799,N_4565);
nand U6243 (N_6243,N_4917,N_5171);
nor U6244 (N_6244,N_5385,N_5287);
nor U6245 (N_6245,N_5485,N_5069);
xor U6246 (N_6246,N_5492,N_5175);
nand U6247 (N_6247,N_4908,N_5665);
and U6248 (N_6248,N_5873,N_5027);
nor U6249 (N_6249,N_4929,N_5854);
nor U6250 (N_6250,N_4517,N_5655);
nor U6251 (N_6251,N_4776,N_4934);
nand U6252 (N_6252,N_4548,N_4546);
nand U6253 (N_6253,N_5573,N_5716);
nor U6254 (N_6254,N_4661,N_5834);
or U6255 (N_6255,N_5159,N_5776);
nor U6256 (N_6256,N_5660,N_5522);
nand U6257 (N_6257,N_5359,N_4609);
and U6258 (N_6258,N_5745,N_5298);
and U6259 (N_6259,N_5885,N_4951);
nor U6260 (N_6260,N_5095,N_5763);
nand U6261 (N_6261,N_5802,N_4507);
or U6262 (N_6262,N_4555,N_5439);
xnor U6263 (N_6263,N_5381,N_5606);
nor U6264 (N_6264,N_5198,N_4769);
nor U6265 (N_6265,N_5356,N_4594);
nor U6266 (N_6266,N_5641,N_4714);
and U6267 (N_6267,N_5268,N_5640);
xnor U6268 (N_6268,N_5603,N_5362);
and U6269 (N_6269,N_5881,N_4981);
or U6270 (N_6270,N_5109,N_4931);
or U6271 (N_6271,N_5866,N_4897);
nand U6272 (N_6272,N_5132,N_5383);
nor U6273 (N_6273,N_4886,N_4765);
nand U6274 (N_6274,N_5552,N_5456);
nand U6275 (N_6275,N_5470,N_4777);
xor U6276 (N_6276,N_5705,N_4638);
or U6277 (N_6277,N_5943,N_5612);
nand U6278 (N_6278,N_5077,N_5239);
nor U6279 (N_6279,N_5294,N_5860);
nor U6280 (N_6280,N_5404,N_5605);
or U6281 (N_6281,N_5070,N_4562);
xor U6282 (N_6282,N_5377,N_4718);
nand U6283 (N_6283,N_5216,N_5694);
nand U6284 (N_6284,N_5348,N_5320);
and U6285 (N_6285,N_4911,N_5636);
and U6286 (N_6286,N_5088,N_4593);
nand U6287 (N_6287,N_5237,N_5756);
nand U6288 (N_6288,N_5266,N_4735);
and U6289 (N_6289,N_5165,N_4791);
nand U6290 (N_6290,N_5335,N_5732);
and U6291 (N_6291,N_5744,N_5700);
and U6292 (N_6292,N_5850,N_5527);
and U6293 (N_6293,N_5024,N_5862);
and U6294 (N_6294,N_5994,N_5114);
nor U6295 (N_6295,N_4693,N_5557);
or U6296 (N_6296,N_5566,N_5318);
and U6297 (N_6297,N_5830,N_4528);
nor U6298 (N_6298,N_5389,N_4775);
nor U6299 (N_6299,N_4869,N_5188);
and U6300 (N_6300,N_5617,N_4940);
xor U6301 (N_6301,N_4649,N_5970);
nor U6302 (N_6302,N_5437,N_5678);
nor U6303 (N_6303,N_5360,N_5789);
and U6304 (N_6304,N_4864,N_5865);
or U6305 (N_6305,N_5471,N_4902);
nor U6306 (N_6306,N_5704,N_4599);
and U6307 (N_6307,N_5484,N_5186);
nor U6308 (N_6308,N_4553,N_4895);
and U6309 (N_6309,N_5153,N_5393);
or U6310 (N_6310,N_4617,N_5767);
xnor U6311 (N_6311,N_5616,N_5755);
or U6312 (N_6312,N_5273,N_5670);
or U6313 (N_6313,N_4960,N_4974);
or U6314 (N_6314,N_4970,N_4831);
and U6315 (N_6315,N_5255,N_5183);
nor U6316 (N_6316,N_5542,N_5047);
and U6317 (N_6317,N_4631,N_4725);
xnor U6318 (N_6318,N_4957,N_5903);
or U6319 (N_6319,N_5976,N_5840);
nor U6320 (N_6320,N_5029,N_5620);
nor U6321 (N_6321,N_4560,N_4797);
and U6322 (N_6322,N_5740,N_5746);
xnor U6323 (N_6323,N_5131,N_5445);
nand U6324 (N_6324,N_5425,N_5920);
nand U6325 (N_6325,N_4671,N_4547);
and U6326 (N_6326,N_4800,N_4773);
nand U6327 (N_6327,N_5209,N_4737);
or U6328 (N_6328,N_4986,N_4645);
nor U6329 (N_6329,N_4510,N_4532);
or U6330 (N_6330,N_4959,N_5134);
and U6331 (N_6331,N_5145,N_5251);
nand U6332 (N_6332,N_4569,N_5274);
nor U6333 (N_6333,N_4500,N_4712);
nand U6334 (N_6334,N_4719,N_5342);
nand U6335 (N_6335,N_5679,N_4564);
or U6336 (N_6336,N_5908,N_4978);
and U6337 (N_6337,N_5814,N_5580);
or U6338 (N_6338,N_5491,N_5911);
nand U6339 (N_6339,N_5097,N_5991);
or U6340 (N_6340,N_5597,N_5753);
and U6341 (N_6341,N_5720,N_5693);
nor U6342 (N_6342,N_5108,N_5010);
nor U6343 (N_6343,N_4866,N_4602);
and U6344 (N_6344,N_5205,N_5702);
or U6345 (N_6345,N_5867,N_5178);
or U6346 (N_6346,N_4544,N_5242);
or U6347 (N_6347,N_5909,N_5719);
nor U6348 (N_6348,N_5275,N_5844);
and U6349 (N_6349,N_5826,N_4756);
or U6350 (N_6350,N_5588,N_5791);
nand U6351 (N_6351,N_4533,N_5279);
and U6352 (N_6352,N_5309,N_5632);
or U6353 (N_6353,N_5871,N_4530);
nor U6354 (N_6354,N_5956,N_5002);
xor U6355 (N_6355,N_4676,N_5572);
or U6356 (N_6356,N_4571,N_5563);
xor U6357 (N_6357,N_5842,N_4858);
nor U6358 (N_6358,N_4928,N_4825);
and U6359 (N_6359,N_5212,N_5236);
and U6360 (N_6360,N_5594,N_5339);
and U6361 (N_6361,N_5758,N_5351);
or U6362 (N_6362,N_5523,N_5697);
or U6363 (N_6363,N_4807,N_4614);
nor U6364 (N_6364,N_5009,N_5562);
xnor U6365 (N_6365,N_5140,N_5149);
or U6366 (N_6366,N_4880,N_5932);
nor U6367 (N_6367,N_5825,N_5992);
nand U6368 (N_6368,N_5280,N_4648);
nor U6369 (N_6369,N_5898,N_4615);
or U6370 (N_6370,N_4520,N_5934);
or U6371 (N_6371,N_4683,N_4956);
or U6372 (N_6372,N_5817,N_5812);
nand U6373 (N_6373,N_5306,N_4806);
nand U6374 (N_6374,N_5619,N_5675);
nand U6375 (N_6375,N_5344,N_5068);
and U6376 (N_6376,N_4870,N_4595);
or U6377 (N_6377,N_5918,N_4830);
xor U6378 (N_6378,N_5046,N_4842);
and U6379 (N_6379,N_4921,N_5708);
and U6380 (N_6380,N_5686,N_4852);
xor U6381 (N_6381,N_4576,N_5661);
or U6382 (N_6382,N_5101,N_5643);
nand U6383 (N_6383,N_5144,N_4620);
or U6384 (N_6384,N_4689,N_4516);
or U6385 (N_6385,N_5227,N_5599);
nand U6386 (N_6386,N_4893,N_4865);
nand U6387 (N_6387,N_5397,N_5000);
xor U6388 (N_6388,N_5529,N_4853);
or U6389 (N_6389,N_4785,N_5013);
or U6390 (N_6390,N_5736,N_5741);
xor U6391 (N_6391,N_4794,N_4540);
nand U6392 (N_6392,N_5997,N_5626);
or U6393 (N_6393,N_5113,N_5766);
nand U6394 (N_6394,N_4796,N_4947);
nand U6395 (N_6395,N_5710,N_4873);
and U6396 (N_6396,N_5234,N_4587);
and U6397 (N_6397,N_5382,N_5590);
nor U6398 (N_6398,N_5341,N_5414);
or U6399 (N_6399,N_4884,N_5821);
nor U6400 (N_6400,N_5465,N_5501);
or U6401 (N_6401,N_5861,N_4881);
nand U6402 (N_6402,N_4900,N_5211);
nor U6403 (N_6403,N_5486,N_5457);
or U6404 (N_6404,N_5950,N_5116);
or U6405 (N_6405,N_5074,N_5989);
or U6406 (N_6406,N_4896,N_5291);
or U6407 (N_6407,N_5419,N_5870);
nand U6408 (N_6408,N_4672,N_4508);
nor U6409 (N_6409,N_5759,N_5622);
nand U6410 (N_6410,N_5033,N_4720);
and U6411 (N_6411,N_5957,N_5405);
nor U6412 (N_6412,N_5975,N_5922);
or U6413 (N_6413,N_5448,N_5961);
nand U6414 (N_6414,N_4674,N_5435);
xor U6415 (N_6415,N_5803,N_5229);
nor U6416 (N_6416,N_5336,N_5174);
or U6417 (N_6417,N_5646,N_5916);
or U6418 (N_6418,N_4767,N_5927);
and U6419 (N_6419,N_5295,N_5610);
and U6420 (N_6420,N_5948,N_5847);
or U6421 (N_6421,N_4747,N_4628);
or U6422 (N_6422,N_5035,N_5146);
xor U6423 (N_6423,N_5852,N_5191);
nor U6424 (N_6424,N_5490,N_4621);
and U6425 (N_6425,N_4710,N_5549);
or U6426 (N_6426,N_5302,N_4855);
nor U6427 (N_6427,N_5006,N_4732);
or U6428 (N_6428,N_5967,N_5584);
nand U6429 (N_6429,N_4552,N_5105);
nor U6430 (N_6430,N_4529,N_5039);
and U6431 (N_6431,N_4821,N_5642);
nand U6432 (N_6432,N_5729,N_5654);
nand U6433 (N_6433,N_5625,N_5502);
nor U6434 (N_6434,N_5900,N_5819);
nor U6435 (N_6435,N_5478,N_5003);
or U6436 (N_6436,N_4937,N_5394);
and U6437 (N_6437,N_5966,N_4846);
nand U6438 (N_6438,N_4804,N_5446);
nand U6439 (N_6439,N_4524,N_5988);
nor U6440 (N_6440,N_5127,N_5408);
or U6441 (N_6441,N_5028,N_4874);
and U6442 (N_6442,N_4781,N_5187);
nor U6443 (N_6443,N_5221,N_5119);
nor U6444 (N_6444,N_5944,N_5079);
nand U6445 (N_6445,N_5418,N_4687);
xor U6446 (N_6446,N_5965,N_5829);
and U6447 (N_6447,N_5218,N_5777);
nand U6448 (N_6448,N_4975,N_4616);
or U6449 (N_6449,N_4788,N_5815);
xor U6450 (N_6450,N_5262,N_4679);
nand U6451 (N_6451,N_5958,N_5735);
nor U6452 (N_6452,N_5748,N_5537);
nor U6453 (N_6453,N_5180,N_5185);
nor U6454 (N_6454,N_5757,N_4574);
nand U6455 (N_6455,N_4906,N_4899);
nand U6456 (N_6456,N_4690,N_5773);
or U6457 (N_6457,N_5352,N_5247);
xnor U6458 (N_6458,N_5505,N_4662);
nand U6459 (N_6459,N_5564,N_5674);
and U6460 (N_6460,N_5322,N_4731);
nand U6461 (N_6461,N_5462,N_5494);
or U6462 (N_6462,N_5001,N_5361);
and U6463 (N_6463,N_4789,N_4944);
and U6464 (N_6464,N_5657,N_4608);
or U6465 (N_6465,N_5621,N_4715);
and U6466 (N_6466,N_4888,N_5434);
or U6467 (N_6467,N_5921,N_4771);
or U6468 (N_6468,N_4702,N_5689);
nor U6469 (N_6469,N_5150,N_4784);
and U6470 (N_6470,N_4536,N_5645);
or U6471 (N_6471,N_4982,N_4738);
or U6472 (N_6472,N_4857,N_4817);
nor U6473 (N_6473,N_5307,N_5303);
and U6474 (N_6474,N_4939,N_4740);
and U6475 (N_6475,N_4558,N_4739);
xnor U6476 (N_6476,N_5463,N_5350);
nor U6477 (N_6477,N_5652,N_5807);
and U6478 (N_6478,N_5087,N_5518);
or U6479 (N_6479,N_5148,N_4967);
xnor U6480 (N_6480,N_4832,N_5053);
and U6481 (N_6481,N_5367,N_5289);
xor U6482 (N_6482,N_5859,N_5593);
nor U6483 (N_6483,N_4877,N_5985);
nor U6484 (N_6484,N_4688,N_5623);
nor U6485 (N_6485,N_4748,N_5281);
xor U6486 (N_6486,N_5206,N_4630);
nand U6487 (N_6487,N_5788,N_5986);
nor U6488 (N_6488,N_5015,N_5938);
or U6489 (N_6489,N_5398,N_5100);
xnor U6490 (N_6490,N_5806,N_5884);
nand U6491 (N_6491,N_5240,N_5995);
nor U6492 (N_6492,N_5019,N_5530);
nand U6493 (N_6493,N_4644,N_5386);
nand U6494 (N_6494,N_5012,N_5747);
or U6495 (N_6495,N_5110,N_4889);
nand U6496 (N_6496,N_4894,N_4626);
nor U6497 (N_6497,N_5790,N_5249);
nor U6498 (N_6498,N_4887,N_5399);
and U6499 (N_6499,N_5699,N_4550);
and U6500 (N_6500,N_5513,N_4629);
and U6501 (N_6501,N_4531,N_5179);
nand U6502 (N_6502,N_4752,N_5214);
or U6503 (N_6503,N_5476,N_5828);
or U6504 (N_6504,N_4585,N_4582);
or U6505 (N_6505,N_5282,N_5798);
nand U6506 (N_6506,N_5553,N_5725);
nand U6507 (N_6507,N_5539,N_5466);
nor U6508 (N_6508,N_5833,N_5378);
nor U6509 (N_6509,N_5208,N_5544);
and U6510 (N_6510,N_5136,N_4603);
nor U6511 (N_6511,N_4820,N_5953);
nor U6512 (N_6512,N_5795,N_5703);
and U6513 (N_6513,N_5233,N_5054);
nand U6514 (N_6514,N_4511,N_5337);
and U6515 (N_6515,N_5112,N_4930);
or U6516 (N_6516,N_5241,N_5554);
and U6517 (N_6517,N_5982,N_4920);
or U6518 (N_6518,N_4938,N_4932);
or U6519 (N_6519,N_5184,N_5454);
or U6520 (N_6520,N_4839,N_4962);
nand U6521 (N_6521,N_4643,N_4723);
or U6522 (N_6522,N_5536,N_4927);
and U6523 (N_6523,N_5935,N_5415);
nand U6524 (N_6524,N_4968,N_5987);
and U6525 (N_6525,N_4591,N_4772);
xnor U6526 (N_6526,N_5324,N_4697);
or U6527 (N_6527,N_5416,N_5786);
nand U6528 (N_6528,N_5734,N_5820);
nand U6529 (N_6529,N_5499,N_5283);
nand U6530 (N_6530,N_5905,N_5197);
nand U6531 (N_6531,N_4726,N_4919);
nor U6532 (N_6532,N_5644,N_5779);
and U6533 (N_6533,N_4993,N_4990);
or U6534 (N_6534,N_4699,N_5596);
or U6535 (N_6535,N_4542,N_4657);
nand U6536 (N_6536,N_5877,N_5781);
or U6537 (N_6537,N_4871,N_4945);
nand U6538 (N_6538,N_5521,N_5330);
or U6539 (N_6539,N_5089,N_5421);
nand U6540 (N_6540,N_5904,N_5031);
nand U6541 (N_6541,N_4522,N_5892);
and U6542 (N_6542,N_5574,N_5420);
and U6543 (N_6543,N_5045,N_4724);
or U6544 (N_6544,N_4991,N_5196);
nor U6545 (N_6545,N_5915,N_5941);
nand U6546 (N_6546,N_5164,N_5577);
xnor U6547 (N_6547,N_4861,N_4891);
nand U6548 (N_6548,N_5550,N_5244);
nand U6549 (N_6549,N_5469,N_4513);
or U6550 (N_6550,N_5879,N_4653);
nor U6551 (N_6551,N_5633,N_5848);
or U6552 (N_6552,N_4868,N_4635);
and U6553 (N_6553,N_5106,N_4698);
nor U6554 (N_6554,N_5650,N_5955);
and U6555 (N_6555,N_5248,N_5692);
and U6556 (N_6556,N_5937,N_5317);
and U6557 (N_6557,N_4573,N_5332);
nand U6558 (N_6558,N_4988,N_4766);
or U6559 (N_6559,N_4678,N_4549);
nor U6560 (N_6560,N_5276,N_5083);
or U6561 (N_6561,N_5924,N_5662);
xor U6562 (N_6562,N_4736,N_5664);
nand U6563 (N_6563,N_5667,N_4501);
nand U6564 (N_6564,N_5836,N_5313);
nor U6565 (N_6565,N_4684,N_5292);
nor U6566 (N_6566,N_4984,N_4566);
and U6567 (N_6567,N_4885,N_4734);
nand U6568 (N_6568,N_4826,N_4835);
xor U6569 (N_6569,N_5687,N_5701);
and U6570 (N_6570,N_5034,N_5585);
and U6571 (N_6571,N_4997,N_4673);
and U6572 (N_6572,N_5157,N_5731);
nor U6573 (N_6573,N_4557,N_5983);
and U6574 (N_6574,N_5535,N_4534);
nor U6575 (N_6575,N_5728,N_5631);
and U6576 (N_6576,N_5768,N_5558);
or U6577 (N_6577,N_4642,N_5869);
and U6578 (N_6578,N_4770,N_5683);
or U6579 (N_6579,N_5125,N_5800);
or U6580 (N_6580,N_4876,N_5441);
and U6581 (N_6581,N_4704,N_5374);
nand U6582 (N_6582,N_5366,N_4792);
and U6583 (N_6583,N_5443,N_5509);
and U6584 (N_6584,N_4559,N_5520);
and U6585 (N_6585,N_4601,N_4525);
nor U6586 (N_6586,N_5098,N_5999);
and U6587 (N_6587,N_5481,N_4822);
xnor U6588 (N_6588,N_5409,N_5005);
nor U6589 (N_6589,N_5567,N_4660);
and U6590 (N_6590,N_5265,N_4707);
nand U6591 (N_6591,N_5048,N_5219);
or U6592 (N_6592,N_5835,N_5831);
nand U6593 (N_6593,N_4909,N_5426);
nand U6594 (N_6594,N_5147,N_4706);
nand U6595 (N_6595,N_5308,N_4768);
nand U6596 (N_6596,N_5738,N_5424);
nor U6597 (N_6597,N_4844,N_5458);
or U6598 (N_6598,N_5727,N_5555);
and U6599 (N_6599,N_5215,N_5055);
and U6600 (N_6600,N_5488,N_5801);
nor U6601 (N_6601,N_5592,N_5316);
and U6602 (N_6602,N_5886,N_5226);
nor U6603 (N_6603,N_4632,N_5224);
or U6604 (N_6604,N_5851,N_4659);
nand U6605 (N_6605,N_4685,N_5473);
nand U6606 (N_6606,N_5919,N_5072);
or U6607 (N_6607,N_5061,N_4999);
xnor U6608 (N_6608,N_5195,N_4795);
nand U6609 (N_6609,N_5085,N_5139);
xnor U6610 (N_6610,N_4754,N_5907);
and U6611 (N_6611,N_5392,N_5682);
nor U6612 (N_6612,N_4953,N_5477);
or U6613 (N_6613,N_5673,N_5081);
xor U6614 (N_6614,N_5681,N_4823);
nand U6615 (N_6615,N_4987,N_5124);
nor U6616 (N_6616,N_4878,N_5161);
nor U6617 (N_6617,N_4570,N_4515);
nor U6618 (N_6618,N_5984,N_5096);
and U6619 (N_6619,N_4538,N_4802);
and U6620 (N_6620,N_5841,N_5375);
and U6621 (N_6621,N_4503,N_5615);
and U6622 (N_6622,N_5981,N_5717);
nor U6623 (N_6623,N_5853,N_5843);
or U6624 (N_6624,N_4837,N_5076);
and U6625 (N_6625,N_5223,N_5506);
or U6626 (N_6626,N_5122,N_4728);
nor U6627 (N_6627,N_5368,N_4782);
nor U6628 (N_6628,N_5376,N_5340);
or U6629 (N_6629,N_5121,N_5155);
and U6630 (N_6630,N_5369,N_5025);
or U6631 (N_6631,N_4543,N_5560);
nand U6632 (N_6632,N_5613,N_5312);
nand U6633 (N_6633,N_4651,N_4758);
nor U6634 (N_6634,N_5455,N_5319);
nand U6635 (N_6635,N_4985,N_5794);
or U6636 (N_6636,N_4815,N_5713);
or U6637 (N_6637,N_4836,N_5474);
nand U6638 (N_6638,N_5516,N_5066);
nor U6639 (N_6639,N_4901,N_4798);
and U6640 (N_6640,N_5823,N_5263);
and U6641 (N_6641,N_5293,N_4646);
nand U6642 (N_6642,N_4600,N_5480);
and U6643 (N_6643,N_5635,N_5296);
nor U6644 (N_6644,N_4636,N_4597);
and U6645 (N_6645,N_4941,N_5813);
or U6646 (N_6646,N_5199,N_5170);
nor U6647 (N_6647,N_5533,N_4803);
xnor U6648 (N_6648,N_5357,N_5111);
and U6649 (N_6649,N_5676,N_5945);
nand U6650 (N_6650,N_5695,N_5115);
xnor U6651 (N_6651,N_4583,N_4805);
or U6652 (N_6652,N_5680,N_4701);
and U6653 (N_6653,N_5151,N_4640);
or U6654 (N_6654,N_4730,N_5810);
and U6655 (N_6655,N_5301,N_5888);
or U6656 (N_6656,N_4958,N_5586);
nor U6657 (N_6657,N_5668,N_5137);
nor U6658 (N_6658,N_5548,N_5444);
nand U6659 (N_6659,N_5771,N_5058);
or U6660 (N_6660,N_5579,N_4639);
nand U6661 (N_6661,N_5816,N_5120);
xnor U6662 (N_6662,N_4681,N_5964);
or U6663 (N_6663,N_4519,N_5245);
and U6664 (N_6664,N_5364,N_5774);
nor U6665 (N_6665,N_5715,N_5093);
and U6666 (N_6666,N_5008,N_5583);
and U6667 (N_6667,N_5578,N_4686);
or U6668 (N_6668,N_5204,N_4665);
or U6669 (N_6669,N_5129,N_5818);
nor U6670 (N_6670,N_5978,N_4545);
nand U6671 (N_6671,N_5947,N_5354);
nor U6672 (N_6672,N_5876,N_5827);
or U6673 (N_6673,N_5065,N_5685);
and U6674 (N_6674,N_4812,N_5752);
or U6675 (N_6675,N_5182,N_5839);
or U6676 (N_6676,N_4814,N_5256);
nor U6677 (N_6677,N_5804,N_4578);
and U6678 (N_6678,N_5902,N_5400);
nor U6679 (N_6679,N_5604,N_5202);
nand U6680 (N_6680,N_5326,N_4828);
or U6681 (N_6681,N_5007,N_4829);
and U6682 (N_6682,N_4512,N_5482);
nand U6683 (N_6683,N_5483,N_5327);
and U6684 (N_6684,N_4910,N_5158);
nand U6685 (N_6685,N_4625,N_5722);
or U6686 (N_6686,N_5709,N_5036);
and U6687 (N_6687,N_5980,N_5391);
nor U6688 (N_6688,N_5856,N_4847);
or U6689 (N_6689,N_5358,N_5030);
and U6690 (N_6690,N_5849,N_5154);
and U6691 (N_6691,N_5461,N_4743);
nor U6692 (N_6692,N_4845,N_5413);
and U6693 (N_6693,N_5428,N_4539);
xnor U6694 (N_6694,N_5824,N_4680);
or U6695 (N_6695,N_5438,N_5962);
and U6696 (N_6696,N_4655,N_5323);
nand U6697 (N_6697,N_4664,N_5845);
nor U6698 (N_6698,N_5166,N_5277);
and U6699 (N_6699,N_4623,N_5669);
or U6700 (N_6700,N_5060,N_4790);
nand U6701 (N_6701,N_5338,N_5018);
or U6702 (N_6702,N_5783,N_4952);
or U6703 (N_6703,N_5569,N_5328);
xor U6704 (N_6704,N_5671,N_5278);
nand U6705 (N_6705,N_5993,N_5656);
xnor U6706 (N_6706,N_5201,N_5799);
or U6707 (N_6707,N_5880,N_4824);
nor U6708 (N_6708,N_5690,N_4633);
xor U6709 (N_6709,N_4722,N_5411);
nor U6710 (N_6710,N_4867,N_4613);
and U6711 (N_6711,N_4556,N_5467);
and U6712 (N_6712,N_5331,N_4610);
xnor U6713 (N_6713,N_5423,N_5193);
and U6714 (N_6714,N_5427,N_5883);
or U6715 (N_6715,N_5609,N_5531);
and U6716 (N_6716,N_5726,N_5914);
or U6717 (N_6717,N_4677,N_5022);
or U6718 (N_6718,N_5541,N_5805);
nand U6719 (N_6719,N_5190,N_4933);
xnor U6720 (N_6720,N_5647,N_4980);
or U6721 (N_6721,N_5349,N_5863);
nand U6722 (N_6722,N_4936,N_5051);
nor U6723 (N_6723,N_5688,N_4998);
or U6724 (N_6724,N_4935,N_5607);
and U6725 (N_6725,N_4856,N_5532);
nor U6726 (N_6726,N_5493,N_4581);
xor U6727 (N_6727,N_5267,N_5232);
xnor U6728 (N_6728,N_5496,N_5460);
and U6729 (N_6729,N_4810,N_5797);
or U6730 (N_6730,N_4879,N_5969);
nand U6731 (N_6731,N_5142,N_4964);
nor U6732 (N_6732,N_5023,N_4979);
or U6733 (N_6733,N_5769,N_5468);
nand U6734 (N_6734,N_5868,N_5406);
xnor U6735 (N_6735,N_5551,N_5020);
or U6736 (N_6736,N_4966,N_4717);
nand U6737 (N_6737,N_5238,N_5417);
nand U6738 (N_6738,N_5857,N_4652);
or U6739 (N_6739,N_5832,N_5346);
nand U6740 (N_6740,N_4668,N_5373);
nor U6741 (N_6741,N_4596,N_5519);
nand U6742 (N_6742,N_4950,N_5545);
nand U6743 (N_6743,N_4848,N_5507);
or U6744 (N_6744,N_5038,N_5565);
nor U6745 (N_6745,N_4746,N_4949);
nand U6746 (N_6746,N_5103,N_5304);
or U6747 (N_6747,N_5169,N_5591);
and U6748 (N_6748,N_4711,N_4537);
nand U6749 (N_6749,N_5479,N_5570);
nand U6750 (N_6750,N_5565,N_5723);
nor U6751 (N_6751,N_5278,N_4906);
nor U6752 (N_6752,N_4829,N_5945);
or U6753 (N_6753,N_4515,N_5942);
nor U6754 (N_6754,N_4513,N_5369);
nand U6755 (N_6755,N_4688,N_5102);
and U6756 (N_6756,N_5943,N_4838);
xnor U6757 (N_6757,N_5664,N_5134);
or U6758 (N_6758,N_5995,N_4740);
and U6759 (N_6759,N_4556,N_4667);
nand U6760 (N_6760,N_5118,N_5580);
and U6761 (N_6761,N_4834,N_4797);
and U6762 (N_6762,N_5982,N_4934);
or U6763 (N_6763,N_4576,N_5111);
nand U6764 (N_6764,N_4735,N_5496);
and U6765 (N_6765,N_4821,N_5906);
and U6766 (N_6766,N_4706,N_5992);
nand U6767 (N_6767,N_4632,N_5023);
nor U6768 (N_6768,N_4615,N_4821);
and U6769 (N_6769,N_5991,N_5496);
and U6770 (N_6770,N_4775,N_5906);
nor U6771 (N_6771,N_5240,N_4833);
nand U6772 (N_6772,N_4776,N_4522);
and U6773 (N_6773,N_5302,N_4949);
or U6774 (N_6774,N_5018,N_5850);
or U6775 (N_6775,N_4529,N_5199);
and U6776 (N_6776,N_5764,N_4662);
nor U6777 (N_6777,N_4892,N_4637);
or U6778 (N_6778,N_4883,N_5666);
nand U6779 (N_6779,N_5743,N_4749);
and U6780 (N_6780,N_5330,N_4909);
nor U6781 (N_6781,N_5923,N_4634);
nand U6782 (N_6782,N_4842,N_5177);
and U6783 (N_6783,N_5004,N_5307);
or U6784 (N_6784,N_5107,N_5484);
or U6785 (N_6785,N_5790,N_5193);
and U6786 (N_6786,N_4540,N_4806);
xnor U6787 (N_6787,N_5387,N_5256);
and U6788 (N_6788,N_5881,N_5297);
nor U6789 (N_6789,N_5598,N_5862);
or U6790 (N_6790,N_5068,N_5411);
nor U6791 (N_6791,N_5452,N_5617);
and U6792 (N_6792,N_5509,N_4774);
or U6793 (N_6793,N_4561,N_5642);
nor U6794 (N_6794,N_4600,N_4899);
nor U6795 (N_6795,N_5413,N_4562);
xnor U6796 (N_6796,N_4761,N_5090);
xor U6797 (N_6797,N_5581,N_4804);
nor U6798 (N_6798,N_5744,N_5174);
or U6799 (N_6799,N_5378,N_5463);
nand U6800 (N_6800,N_5605,N_5222);
or U6801 (N_6801,N_5985,N_4982);
nand U6802 (N_6802,N_5877,N_5072);
nor U6803 (N_6803,N_4520,N_5029);
nor U6804 (N_6804,N_4725,N_5940);
and U6805 (N_6805,N_4670,N_4819);
nand U6806 (N_6806,N_5206,N_5561);
or U6807 (N_6807,N_4640,N_5250);
and U6808 (N_6808,N_5709,N_5064);
nor U6809 (N_6809,N_5888,N_5948);
or U6810 (N_6810,N_4825,N_4740);
or U6811 (N_6811,N_5211,N_5577);
nor U6812 (N_6812,N_4625,N_5016);
xnor U6813 (N_6813,N_4520,N_5852);
nor U6814 (N_6814,N_5102,N_4896);
nand U6815 (N_6815,N_4947,N_4720);
nor U6816 (N_6816,N_4980,N_4667);
nor U6817 (N_6817,N_5593,N_5928);
or U6818 (N_6818,N_5836,N_5327);
or U6819 (N_6819,N_4777,N_4698);
nand U6820 (N_6820,N_5592,N_5359);
nand U6821 (N_6821,N_5315,N_5781);
or U6822 (N_6822,N_4663,N_5601);
nor U6823 (N_6823,N_5392,N_4768);
nand U6824 (N_6824,N_4859,N_4506);
nor U6825 (N_6825,N_4846,N_4546);
and U6826 (N_6826,N_5551,N_4840);
nor U6827 (N_6827,N_4968,N_5123);
nor U6828 (N_6828,N_4695,N_4507);
nand U6829 (N_6829,N_4516,N_4948);
nand U6830 (N_6830,N_5234,N_5490);
and U6831 (N_6831,N_4911,N_4791);
nor U6832 (N_6832,N_5651,N_5447);
nor U6833 (N_6833,N_5633,N_5414);
or U6834 (N_6834,N_5570,N_5328);
nand U6835 (N_6835,N_5601,N_4932);
nand U6836 (N_6836,N_5067,N_5769);
nand U6837 (N_6837,N_4944,N_5712);
nor U6838 (N_6838,N_5739,N_5223);
nor U6839 (N_6839,N_5327,N_5933);
and U6840 (N_6840,N_5190,N_4840);
nor U6841 (N_6841,N_5187,N_5115);
nand U6842 (N_6842,N_4778,N_5646);
or U6843 (N_6843,N_5079,N_5593);
nand U6844 (N_6844,N_5127,N_5325);
and U6845 (N_6845,N_5008,N_4797);
nor U6846 (N_6846,N_5965,N_5498);
nor U6847 (N_6847,N_5607,N_4599);
nand U6848 (N_6848,N_5217,N_4982);
or U6849 (N_6849,N_4884,N_5607);
nand U6850 (N_6850,N_4615,N_5491);
nor U6851 (N_6851,N_5507,N_5918);
or U6852 (N_6852,N_4640,N_5234);
or U6853 (N_6853,N_4887,N_5317);
nor U6854 (N_6854,N_5956,N_4920);
or U6855 (N_6855,N_5288,N_5518);
or U6856 (N_6856,N_4830,N_4971);
nand U6857 (N_6857,N_4912,N_5746);
or U6858 (N_6858,N_5890,N_5432);
nor U6859 (N_6859,N_5710,N_5867);
or U6860 (N_6860,N_5887,N_4822);
or U6861 (N_6861,N_5888,N_5413);
nor U6862 (N_6862,N_5604,N_4523);
nor U6863 (N_6863,N_5445,N_5894);
or U6864 (N_6864,N_4839,N_4809);
nor U6865 (N_6865,N_5581,N_5959);
xor U6866 (N_6866,N_5886,N_5093);
nor U6867 (N_6867,N_5718,N_4762);
and U6868 (N_6868,N_5165,N_5386);
nand U6869 (N_6869,N_5035,N_5132);
and U6870 (N_6870,N_5302,N_4713);
nor U6871 (N_6871,N_4778,N_4585);
or U6872 (N_6872,N_5863,N_5325);
nand U6873 (N_6873,N_5021,N_4552);
and U6874 (N_6874,N_5736,N_5723);
nor U6875 (N_6875,N_5777,N_5829);
nor U6876 (N_6876,N_5613,N_5412);
nor U6877 (N_6877,N_5280,N_4766);
and U6878 (N_6878,N_5561,N_5630);
nor U6879 (N_6879,N_5210,N_5676);
and U6880 (N_6880,N_4772,N_4502);
or U6881 (N_6881,N_4512,N_5344);
and U6882 (N_6882,N_5823,N_5802);
xnor U6883 (N_6883,N_5972,N_5626);
nor U6884 (N_6884,N_5446,N_4719);
xnor U6885 (N_6885,N_5163,N_4602);
or U6886 (N_6886,N_4798,N_5020);
and U6887 (N_6887,N_5142,N_5635);
nand U6888 (N_6888,N_5049,N_4639);
and U6889 (N_6889,N_5535,N_5240);
or U6890 (N_6890,N_4712,N_5303);
and U6891 (N_6891,N_5950,N_5752);
and U6892 (N_6892,N_5063,N_5823);
and U6893 (N_6893,N_4558,N_5727);
or U6894 (N_6894,N_4923,N_4712);
xor U6895 (N_6895,N_4923,N_5622);
nor U6896 (N_6896,N_5573,N_4807);
and U6897 (N_6897,N_4830,N_5126);
xnor U6898 (N_6898,N_5771,N_5208);
or U6899 (N_6899,N_5286,N_4780);
nand U6900 (N_6900,N_5615,N_5366);
nand U6901 (N_6901,N_5315,N_4859);
nor U6902 (N_6902,N_5057,N_4662);
and U6903 (N_6903,N_5811,N_5436);
or U6904 (N_6904,N_4760,N_4931);
or U6905 (N_6905,N_5194,N_4570);
nand U6906 (N_6906,N_5025,N_4567);
and U6907 (N_6907,N_5664,N_4843);
or U6908 (N_6908,N_5069,N_4939);
nand U6909 (N_6909,N_5320,N_5220);
nand U6910 (N_6910,N_5449,N_4530);
or U6911 (N_6911,N_4919,N_5592);
nand U6912 (N_6912,N_5792,N_4939);
nand U6913 (N_6913,N_4763,N_5196);
and U6914 (N_6914,N_5395,N_5876);
xor U6915 (N_6915,N_4569,N_5910);
nor U6916 (N_6916,N_4884,N_5030);
nand U6917 (N_6917,N_4860,N_5092);
and U6918 (N_6918,N_5628,N_5635);
nor U6919 (N_6919,N_5196,N_5720);
nor U6920 (N_6920,N_5631,N_5961);
xor U6921 (N_6921,N_5001,N_5309);
or U6922 (N_6922,N_5727,N_5627);
or U6923 (N_6923,N_5334,N_5640);
nor U6924 (N_6924,N_4763,N_4569);
nand U6925 (N_6925,N_5466,N_5715);
nor U6926 (N_6926,N_5323,N_5593);
or U6927 (N_6927,N_5152,N_4995);
and U6928 (N_6928,N_4690,N_5926);
or U6929 (N_6929,N_5125,N_4858);
or U6930 (N_6930,N_5453,N_5932);
nor U6931 (N_6931,N_5260,N_5533);
nor U6932 (N_6932,N_5628,N_5100);
nand U6933 (N_6933,N_5772,N_4840);
nand U6934 (N_6934,N_4823,N_5906);
nand U6935 (N_6935,N_5747,N_5883);
xor U6936 (N_6936,N_5227,N_4582);
nand U6937 (N_6937,N_5159,N_4674);
nand U6938 (N_6938,N_4765,N_5489);
or U6939 (N_6939,N_5454,N_4658);
nor U6940 (N_6940,N_4873,N_5233);
nor U6941 (N_6941,N_5627,N_5411);
and U6942 (N_6942,N_5993,N_4713);
or U6943 (N_6943,N_5070,N_5947);
or U6944 (N_6944,N_5429,N_5161);
or U6945 (N_6945,N_5698,N_4639);
and U6946 (N_6946,N_5418,N_5018);
nor U6947 (N_6947,N_4941,N_5328);
and U6948 (N_6948,N_5325,N_5220);
nor U6949 (N_6949,N_4561,N_5457);
nand U6950 (N_6950,N_5475,N_4844);
xnor U6951 (N_6951,N_5295,N_5478);
nor U6952 (N_6952,N_4726,N_5160);
and U6953 (N_6953,N_5571,N_5755);
nand U6954 (N_6954,N_5809,N_5181);
or U6955 (N_6955,N_5367,N_5657);
nand U6956 (N_6956,N_5709,N_5533);
nand U6957 (N_6957,N_5242,N_5516);
nor U6958 (N_6958,N_4696,N_5638);
xnor U6959 (N_6959,N_5040,N_5053);
xor U6960 (N_6960,N_5463,N_4731);
and U6961 (N_6961,N_4894,N_4873);
nand U6962 (N_6962,N_5248,N_4642);
nand U6963 (N_6963,N_5318,N_4732);
or U6964 (N_6964,N_4846,N_5552);
and U6965 (N_6965,N_5015,N_5153);
or U6966 (N_6966,N_5600,N_5019);
and U6967 (N_6967,N_4863,N_5335);
and U6968 (N_6968,N_4738,N_5087);
xnor U6969 (N_6969,N_5326,N_4825);
and U6970 (N_6970,N_4652,N_4536);
and U6971 (N_6971,N_5112,N_4619);
or U6972 (N_6972,N_5863,N_5973);
nand U6973 (N_6973,N_4952,N_4543);
xnor U6974 (N_6974,N_5691,N_4757);
nor U6975 (N_6975,N_5982,N_4865);
or U6976 (N_6976,N_5954,N_4725);
nand U6977 (N_6977,N_5151,N_4871);
nand U6978 (N_6978,N_5179,N_4732);
or U6979 (N_6979,N_4824,N_5487);
nand U6980 (N_6980,N_5802,N_5327);
nand U6981 (N_6981,N_5208,N_5648);
and U6982 (N_6982,N_4954,N_4542);
or U6983 (N_6983,N_4898,N_5901);
nand U6984 (N_6984,N_4644,N_5523);
nor U6985 (N_6985,N_5371,N_5687);
and U6986 (N_6986,N_4898,N_5744);
xor U6987 (N_6987,N_5725,N_5472);
nand U6988 (N_6988,N_4651,N_5754);
or U6989 (N_6989,N_5746,N_4663);
nor U6990 (N_6990,N_5180,N_4998);
nor U6991 (N_6991,N_5226,N_5215);
nand U6992 (N_6992,N_4973,N_5507);
nor U6993 (N_6993,N_5599,N_5405);
and U6994 (N_6994,N_5988,N_4804);
xor U6995 (N_6995,N_4988,N_5822);
or U6996 (N_6996,N_5007,N_5161);
nor U6997 (N_6997,N_4536,N_4706);
and U6998 (N_6998,N_4624,N_4691);
or U6999 (N_6999,N_5500,N_4530);
or U7000 (N_7000,N_4766,N_4906);
and U7001 (N_7001,N_4794,N_4977);
nor U7002 (N_7002,N_5556,N_4687);
nor U7003 (N_7003,N_4866,N_5770);
nand U7004 (N_7004,N_5862,N_5990);
nand U7005 (N_7005,N_5268,N_4769);
nand U7006 (N_7006,N_5280,N_5661);
nand U7007 (N_7007,N_5516,N_5221);
and U7008 (N_7008,N_5395,N_5119);
nor U7009 (N_7009,N_4872,N_5346);
and U7010 (N_7010,N_4687,N_5858);
nor U7011 (N_7011,N_5933,N_4591);
and U7012 (N_7012,N_4672,N_5565);
and U7013 (N_7013,N_5752,N_5646);
or U7014 (N_7014,N_5687,N_5137);
nor U7015 (N_7015,N_4967,N_5141);
or U7016 (N_7016,N_5126,N_4746);
or U7017 (N_7017,N_4706,N_4606);
or U7018 (N_7018,N_5319,N_4581);
or U7019 (N_7019,N_5656,N_5096);
nor U7020 (N_7020,N_5316,N_5533);
nor U7021 (N_7021,N_5795,N_5163);
nand U7022 (N_7022,N_5479,N_5156);
and U7023 (N_7023,N_5486,N_5153);
and U7024 (N_7024,N_4923,N_5304);
nor U7025 (N_7025,N_5491,N_4617);
xnor U7026 (N_7026,N_4722,N_5078);
or U7027 (N_7027,N_5905,N_5061);
nor U7028 (N_7028,N_5128,N_4551);
nand U7029 (N_7029,N_5280,N_4919);
or U7030 (N_7030,N_5964,N_4987);
nand U7031 (N_7031,N_4595,N_5903);
or U7032 (N_7032,N_5033,N_5170);
nand U7033 (N_7033,N_4594,N_5344);
or U7034 (N_7034,N_5066,N_5098);
and U7035 (N_7035,N_4551,N_5241);
and U7036 (N_7036,N_5175,N_5771);
and U7037 (N_7037,N_5826,N_4709);
xnor U7038 (N_7038,N_4764,N_5816);
and U7039 (N_7039,N_4844,N_5157);
or U7040 (N_7040,N_5789,N_5558);
nand U7041 (N_7041,N_4508,N_5191);
and U7042 (N_7042,N_5103,N_4578);
and U7043 (N_7043,N_5933,N_5896);
nand U7044 (N_7044,N_5144,N_5691);
xor U7045 (N_7045,N_4548,N_5709);
nor U7046 (N_7046,N_5591,N_4836);
and U7047 (N_7047,N_5230,N_4934);
nand U7048 (N_7048,N_4793,N_4931);
or U7049 (N_7049,N_5240,N_4640);
or U7050 (N_7050,N_5465,N_4776);
and U7051 (N_7051,N_5211,N_4529);
or U7052 (N_7052,N_5520,N_5715);
nand U7053 (N_7053,N_5852,N_4927);
and U7054 (N_7054,N_5557,N_4881);
nand U7055 (N_7055,N_5605,N_5031);
or U7056 (N_7056,N_4965,N_4630);
nand U7057 (N_7057,N_5631,N_5030);
nor U7058 (N_7058,N_4983,N_5564);
xor U7059 (N_7059,N_4924,N_5095);
and U7060 (N_7060,N_4589,N_5593);
or U7061 (N_7061,N_5823,N_4588);
xnor U7062 (N_7062,N_5770,N_5482);
or U7063 (N_7063,N_5966,N_4871);
nand U7064 (N_7064,N_5457,N_4696);
and U7065 (N_7065,N_5669,N_5101);
nand U7066 (N_7066,N_5334,N_4648);
nor U7067 (N_7067,N_5020,N_5077);
nor U7068 (N_7068,N_5807,N_5837);
nor U7069 (N_7069,N_5799,N_5831);
nor U7070 (N_7070,N_4521,N_4856);
nand U7071 (N_7071,N_5414,N_5068);
xor U7072 (N_7072,N_4754,N_4826);
or U7073 (N_7073,N_5227,N_5238);
nor U7074 (N_7074,N_4935,N_5139);
xor U7075 (N_7075,N_5413,N_5540);
or U7076 (N_7076,N_4690,N_5436);
nand U7077 (N_7077,N_5480,N_5345);
nand U7078 (N_7078,N_5683,N_4622);
and U7079 (N_7079,N_5338,N_4908);
nand U7080 (N_7080,N_4611,N_5859);
xnor U7081 (N_7081,N_5564,N_5844);
nand U7082 (N_7082,N_4918,N_5624);
or U7083 (N_7083,N_5512,N_5194);
nor U7084 (N_7084,N_5464,N_4537);
and U7085 (N_7085,N_5496,N_5874);
or U7086 (N_7086,N_4873,N_5334);
or U7087 (N_7087,N_5722,N_5152);
nand U7088 (N_7088,N_4965,N_5690);
nand U7089 (N_7089,N_4636,N_5300);
nand U7090 (N_7090,N_5585,N_5607);
and U7091 (N_7091,N_4671,N_5448);
or U7092 (N_7092,N_5406,N_5127);
xor U7093 (N_7093,N_4921,N_4584);
and U7094 (N_7094,N_4533,N_4572);
nand U7095 (N_7095,N_4630,N_4883);
nor U7096 (N_7096,N_5600,N_4947);
nor U7097 (N_7097,N_5044,N_4910);
or U7098 (N_7098,N_5528,N_5739);
nand U7099 (N_7099,N_5805,N_5930);
nand U7100 (N_7100,N_4751,N_5193);
or U7101 (N_7101,N_5888,N_4675);
and U7102 (N_7102,N_5393,N_4633);
nand U7103 (N_7103,N_5934,N_5808);
and U7104 (N_7104,N_4877,N_5953);
and U7105 (N_7105,N_4581,N_4853);
nor U7106 (N_7106,N_4843,N_5287);
nor U7107 (N_7107,N_4518,N_5219);
xnor U7108 (N_7108,N_5293,N_5115);
nor U7109 (N_7109,N_5382,N_4974);
or U7110 (N_7110,N_4597,N_5614);
or U7111 (N_7111,N_5272,N_5172);
and U7112 (N_7112,N_4646,N_5703);
nand U7113 (N_7113,N_5658,N_5794);
nand U7114 (N_7114,N_5976,N_4735);
nor U7115 (N_7115,N_4782,N_5192);
nand U7116 (N_7116,N_4751,N_5521);
nand U7117 (N_7117,N_5351,N_5017);
nor U7118 (N_7118,N_4894,N_5000);
or U7119 (N_7119,N_5696,N_4768);
and U7120 (N_7120,N_5207,N_4863);
nor U7121 (N_7121,N_5473,N_5752);
or U7122 (N_7122,N_5696,N_5856);
nor U7123 (N_7123,N_4709,N_5824);
nand U7124 (N_7124,N_5269,N_4790);
nand U7125 (N_7125,N_5091,N_4726);
nor U7126 (N_7126,N_5074,N_5888);
nor U7127 (N_7127,N_4862,N_5883);
and U7128 (N_7128,N_5662,N_5550);
and U7129 (N_7129,N_4939,N_5067);
nand U7130 (N_7130,N_5207,N_4597);
or U7131 (N_7131,N_4593,N_4848);
nor U7132 (N_7132,N_4784,N_5490);
or U7133 (N_7133,N_4698,N_4852);
or U7134 (N_7134,N_5302,N_5001);
or U7135 (N_7135,N_4502,N_4607);
nor U7136 (N_7136,N_5791,N_5964);
nor U7137 (N_7137,N_5279,N_4747);
or U7138 (N_7138,N_5149,N_5581);
xnor U7139 (N_7139,N_5759,N_5659);
or U7140 (N_7140,N_4985,N_5270);
or U7141 (N_7141,N_5055,N_4981);
nand U7142 (N_7142,N_5339,N_5274);
xor U7143 (N_7143,N_4544,N_5144);
nand U7144 (N_7144,N_4675,N_5745);
xor U7145 (N_7145,N_4644,N_4846);
and U7146 (N_7146,N_5954,N_5766);
xnor U7147 (N_7147,N_5870,N_4922);
nor U7148 (N_7148,N_5868,N_5210);
nor U7149 (N_7149,N_4738,N_5986);
nand U7150 (N_7150,N_4703,N_4678);
and U7151 (N_7151,N_5983,N_5479);
nand U7152 (N_7152,N_5528,N_5297);
xnor U7153 (N_7153,N_4648,N_4865);
or U7154 (N_7154,N_5398,N_4983);
nand U7155 (N_7155,N_5550,N_5509);
nand U7156 (N_7156,N_5482,N_5528);
and U7157 (N_7157,N_5989,N_4877);
xnor U7158 (N_7158,N_5648,N_5699);
and U7159 (N_7159,N_4686,N_5310);
nor U7160 (N_7160,N_5116,N_5905);
xnor U7161 (N_7161,N_5522,N_4683);
or U7162 (N_7162,N_5531,N_5183);
xor U7163 (N_7163,N_5575,N_5893);
or U7164 (N_7164,N_5619,N_5199);
nand U7165 (N_7165,N_4567,N_5677);
xor U7166 (N_7166,N_4967,N_4739);
and U7167 (N_7167,N_4876,N_4994);
nand U7168 (N_7168,N_5414,N_5392);
nor U7169 (N_7169,N_5656,N_4973);
xnor U7170 (N_7170,N_5331,N_5801);
nand U7171 (N_7171,N_4885,N_5149);
nand U7172 (N_7172,N_5764,N_4770);
or U7173 (N_7173,N_5113,N_5849);
nand U7174 (N_7174,N_5456,N_4655);
and U7175 (N_7175,N_5523,N_5758);
xnor U7176 (N_7176,N_4867,N_5671);
nand U7177 (N_7177,N_4982,N_4620);
or U7178 (N_7178,N_5622,N_5562);
or U7179 (N_7179,N_5060,N_5420);
nor U7180 (N_7180,N_5013,N_5581);
or U7181 (N_7181,N_4640,N_5034);
nand U7182 (N_7182,N_4993,N_5616);
nand U7183 (N_7183,N_4847,N_5307);
nor U7184 (N_7184,N_5139,N_5956);
or U7185 (N_7185,N_5409,N_4712);
nand U7186 (N_7186,N_4611,N_4600);
and U7187 (N_7187,N_4648,N_4806);
nor U7188 (N_7188,N_5523,N_5996);
nand U7189 (N_7189,N_5262,N_4997);
and U7190 (N_7190,N_5173,N_5305);
and U7191 (N_7191,N_5155,N_5906);
xor U7192 (N_7192,N_5832,N_5304);
or U7193 (N_7193,N_5923,N_5315);
nand U7194 (N_7194,N_5385,N_5199);
or U7195 (N_7195,N_5364,N_5512);
and U7196 (N_7196,N_5691,N_5595);
nor U7197 (N_7197,N_5392,N_5678);
and U7198 (N_7198,N_5914,N_4776);
or U7199 (N_7199,N_4843,N_4663);
xor U7200 (N_7200,N_5454,N_5130);
or U7201 (N_7201,N_5175,N_4944);
or U7202 (N_7202,N_5571,N_4891);
xor U7203 (N_7203,N_5037,N_4565);
nor U7204 (N_7204,N_4798,N_5315);
and U7205 (N_7205,N_5517,N_5676);
or U7206 (N_7206,N_5418,N_5231);
and U7207 (N_7207,N_5789,N_4986);
or U7208 (N_7208,N_5138,N_5681);
or U7209 (N_7209,N_4939,N_4978);
xnor U7210 (N_7210,N_5956,N_5369);
nand U7211 (N_7211,N_5414,N_5307);
nand U7212 (N_7212,N_5542,N_5075);
nand U7213 (N_7213,N_4824,N_5627);
xor U7214 (N_7214,N_4513,N_5185);
nor U7215 (N_7215,N_5986,N_5103);
nor U7216 (N_7216,N_5498,N_4514);
or U7217 (N_7217,N_4712,N_5508);
and U7218 (N_7218,N_4652,N_5915);
nor U7219 (N_7219,N_5367,N_5209);
or U7220 (N_7220,N_5306,N_5824);
or U7221 (N_7221,N_4634,N_5268);
or U7222 (N_7222,N_5434,N_5564);
and U7223 (N_7223,N_4971,N_4691);
nand U7224 (N_7224,N_5306,N_4607);
nor U7225 (N_7225,N_4502,N_4881);
nor U7226 (N_7226,N_5874,N_4555);
and U7227 (N_7227,N_4577,N_4939);
nand U7228 (N_7228,N_5015,N_5728);
nand U7229 (N_7229,N_4724,N_4617);
nand U7230 (N_7230,N_5347,N_5847);
and U7231 (N_7231,N_5290,N_4915);
nand U7232 (N_7232,N_5592,N_4704);
and U7233 (N_7233,N_5050,N_5584);
nand U7234 (N_7234,N_5559,N_5150);
nand U7235 (N_7235,N_5996,N_4669);
nand U7236 (N_7236,N_5505,N_5534);
and U7237 (N_7237,N_5397,N_4727);
nor U7238 (N_7238,N_4867,N_4803);
and U7239 (N_7239,N_5716,N_5238);
or U7240 (N_7240,N_5389,N_5034);
or U7241 (N_7241,N_5530,N_5748);
and U7242 (N_7242,N_5989,N_5577);
and U7243 (N_7243,N_5489,N_5988);
and U7244 (N_7244,N_4833,N_5092);
and U7245 (N_7245,N_5984,N_5936);
or U7246 (N_7246,N_5820,N_5852);
nand U7247 (N_7247,N_4674,N_5554);
nor U7248 (N_7248,N_5643,N_5641);
and U7249 (N_7249,N_5126,N_5171);
or U7250 (N_7250,N_4673,N_4948);
nor U7251 (N_7251,N_5528,N_5421);
nor U7252 (N_7252,N_4931,N_5226);
and U7253 (N_7253,N_5391,N_5486);
nand U7254 (N_7254,N_5737,N_4648);
nor U7255 (N_7255,N_5056,N_5946);
nor U7256 (N_7256,N_5350,N_5014);
nand U7257 (N_7257,N_4894,N_5090);
and U7258 (N_7258,N_4597,N_5724);
or U7259 (N_7259,N_5754,N_5923);
and U7260 (N_7260,N_4616,N_4505);
or U7261 (N_7261,N_5103,N_5015);
nand U7262 (N_7262,N_5820,N_5528);
nor U7263 (N_7263,N_5726,N_4741);
or U7264 (N_7264,N_4718,N_4530);
or U7265 (N_7265,N_4841,N_5637);
and U7266 (N_7266,N_5658,N_4750);
and U7267 (N_7267,N_5679,N_5172);
nor U7268 (N_7268,N_5605,N_5432);
or U7269 (N_7269,N_4708,N_5443);
nor U7270 (N_7270,N_4945,N_5561);
and U7271 (N_7271,N_4901,N_4521);
and U7272 (N_7272,N_5575,N_5211);
and U7273 (N_7273,N_4825,N_5745);
and U7274 (N_7274,N_5294,N_5859);
and U7275 (N_7275,N_4556,N_5105);
xnor U7276 (N_7276,N_5286,N_5720);
or U7277 (N_7277,N_5012,N_4785);
or U7278 (N_7278,N_4628,N_5713);
nor U7279 (N_7279,N_4541,N_5032);
nor U7280 (N_7280,N_4529,N_5674);
nor U7281 (N_7281,N_5117,N_5683);
nor U7282 (N_7282,N_5150,N_5083);
xnor U7283 (N_7283,N_4953,N_5533);
xnor U7284 (N_7284,N_5569,N_4858);
and U7285 (N_7285,N_5689,N_5727);
or U7286 (N_7286,N_4972,N_5938);
nor U7287 (N_7287,N_5682,N_4991);
nor U7288 (N_7288,N_5759,N_4949);
and U7289 (N_7289,N_4709,N_5844);
xor U7290 (N_7290,N_5784,N_4794);
nand U7291 (N_7291,N_5985,N_5997);
and U7292 (N_7292,N_5784,N_5677);
nor U7293 (N_7293,N_4795,N_4947);
nor U7294 (N_7294,N_5594,N_4532);
nor U7295 (N_7295,N_5955,N_5463);
and U7296 (N_7296,N_5936,N_5377);
and U7297 (N_7297,N_4643,N_5508);
xor U7298 (N_7298,N_4943,N_4511);
and U7299 (N_7299,N_5705,N_5998);
and U7300 (N_7300,N_5484,N_5521);
nand U7301 (N_7301,N_4949,N_5047);
and U7302 (N_7302,N_5623,N_5617);
and U7303 (N_7303,N_5104,N_5961);
nor U7304 (N_7304,N_5520,N_5668);
nor U7305 (N_7305,N_5811,N_5257);
and U7306 (N_7306,N_5700,N_5360);
nand U7307 (N_7307,N_5938,N_5098);
nor U7308 (N_7308,N_5431,N_4529);
or U7309 (N_7309,N_4514,N_5312);
nand U7310 (N_7310,N_4830,N_5938);
nor U7311 (N_7311,N_5542,N_5674);
and U7312 (N_7312,N_5608,N_5532);
or U7313 (N_7313,N_5361,N_4719);
and U7314 (N_7314,N_5945,N_5536);
and U7315 (N_7315,N_5073,N_5508);
and U7316 (N_7316,N_5647,N_4653);
nand U7317 (N_7317,N_5726,N_4586);
nand U7318 (N_7318,N_5380,N_5357);
nor U7319 (N_7319,N_5476,N_5717);
nor U7320 (N_7320,N_5673,N_5473);
or U7321 (N_7321,N_5766,N_5631);
nand U7322 (N_7322,N_5298,N_4938);
or U7323 (N_7323,N_5582,N_5314);
or U7324 (N_7324,N_5084,N_5408);
nand U7325 (N_7325,N_4507,N_5148);
xnor U7326 (N_7326,N_5934,N_4513);
nor U7327 (N_7327,N_5810,N_4522);
nor U7328 (N_7328,N_5681,N_5474);
nand U7329 (N_7329,N_4533,N_5930);
and U7330 (N_7330,N_5469,N_5427);
nand U7331 (N_7331,N_5206,N_5068);
and U7332 (N_7332,N_4553,N_5573);
and U7333 (N_7333,N_5093,N_5589);
or U7334 (N_7334,N_5906,N_4971);
nor U7335 (N_7335,N_5934,N_5682);
nor U7336 (N_7336,N_5025,N_4974);
and U7337 (N_7337,N_5446,N_4885);
nand U7338 (N_7338,N_5785,N_4759);
or U7339 (N_7339,N_5521,N_5526);
nor U7340 (N_7340,N_5062,N_5476);
xnor U7341 (N_7341,N_5741,N_5609);
nor U7342 (N_7342,N_5724,N_4549);
xnor U7343 (N_7343,N_4985,N_4666);
xnor U7344 (N_7344,N_5285,N_4783);
and U7345 (N_7345,N_5218,N_4819);
or U7346 (N_7346,N_5030,N_5199);
or U7347 (N_7347,N_5243,N_5851);
or U7348 (N_7348,N_5513,N_5559);
nand U7349 (N_7349,N_5497,N_4609);
nand U7350 (N_7350,N_5314,N_4669);
and U7351 (N_7351,N_5022,N_4977);
nor U7352 (N_7352,N_4722,N_5599);
nor U7353 (N_7353,N_5874,N_4563);
xnor U7354 (N_7354,N_5195,N_4664);
xnor U7355 (N_7355,N_4837,N_4807);
nor U7356 (N_7356,N_5779,N_5568);
nand U7357 (N_7357,N_5118,N_4543);
nor U7358 (N_7358,N_5217,N_4609);
nand U7359 (N_7359,N_5093,N_4646);
xor U7360 (N_7360,N_5279,N_4682);
or U7361 (N_7361,N_5423,N_5642);
or U7362 (N_7362,N_5706,N_5998);
or U7363 (N_7363,N_5686,N_5806);
nand U7364 (N_7364,N_4992,N_4842);
xnor U7365 (N_7365,N_5540,N_5721);
nor U7366 (N_7366,N_5155,N_4861);
and U7367 (N_7367,N_5790,N_4964);
xnor U7368 (N_7368,N_4968,N_5419);
nand U7369 (N_7369,N_5025,N_4599);
or U7370 (N_7370,N_5331,N_5539);
nand U7371 (N_7371,N_5113,N_5210);
nor U7372 (N_7372,N_4831,N_4531);
or U7373 (N_7373,N_4740,N_4693);
nor U7374 (N_7374,N_5603,N_5882);
or U7375 (N_7375,N_5478,N_5441);
nor U7376 (N_7376,N_4970,N_5379);
xor U7377 (N_7377,N_5117,N_5721);
and U7378 (N_7378,N_5593,N_5508);
and U7379 (N_7379,N_5144,N_5540);
or U7380 (N_7380,N_5321,N_5391);
nor U7381 (N_7381,N_4752,N_5646);
xnor U7382 (N_7382,N_4958,N_5136);
or U7383 (N_7383,N_4565,N_4619);
nand U7384 (N_7384,N_5363,N_4753);
or U7385 (N_7385,N_4500,N_5530);
nor U7386 (N_7386,N_5926,N_4575);
or U7387 (N_7387,N_5301,N_4760);
or U7388 (N_7388,N_5003,N_4763);
or U7389 (N_7389,N_5190,N_4510);
and U7390 (N_7390,N_5342,N_5482);
or U7391 (N_7391,N_4919,N_5932);
nor U7392 (N_7392,N_5740,N_5611);
and U7393 (N_7393,N_5163,N_5352);
and U7394 (N_7394,N_5194,N_5836);
nor U7395 (N_7395,N_4581,N_4501);
and U7396 (N_7396,N_4862,N_5777);
nor U7397 (N_7397,N_4808,N_4708);
or U7398 (N_7398,N_5763,N_5032);
or U7399 (N_7399,N_4992,N_4789);
nor U7400 (N_7400,N_4591,N_4526);
or U7401 (N_7401,N_4825,N_5653);
and U7402 (N_7402,N_5259,N_4634);
nand U7403 (N_7403,N_5926,N_5664);
nor U7404 (N_7404,N_5967,N_5740);
xnor U7405 (N_7405,N_4716,N_5288);
or U7406 (N_7406,N_5682,N_5471);
xnor U7407 (N_7407,N_4869,N_4809);
or U7408 (N_7408,N_5517,N_5879);
xor U7409 (N_7409,N_4579,N_4804);
or U7410 (N_7410,N_5194,N_4511);
or U7411 (N_7411,N_4569,N_5542);
or U7412 (N_7412,N_4886,N_4743);
xnor U7413 (N_7413,N_4940,N_4542);
and U7414 (N_7414,N_5933,N_4643);
or U7415 (N_7415,N_5130,N_5927);
nor U7416 (N_7416,N_5819,N_4713);
xor U7417 (N_7417,N_5020,N_4778);
nand U7418 (N_7418,N_5816,N_5973);
nand U7419 (N_7419,N_5419,N_5175);
nor U7420 (N_7420,N_4597,N_5469);
nand U7421 (N_7421,N_5391,N_5346);
and U7422 (N_7422,N_5640,N_4678);
nor U7423 (N_7423,N_5828,N_5853);
or U7424 (N_7424,N_5557,N_5526);
and U7425 (N_7425,N_4818,N_4635);
or U7426 (N_7426,N_4960,N_5121);
or U7427 (N_7427,N_5718,N_5374);
or U7428 (N_7428,N_5508,N_4682);
nand U7429 (N_7429,N_5315,N_5809);
nand U7430 (N_7430,N_4522,N_5195);
nor U7431 (N_7431,N_4978,N_4508);
xnor U7432 (N_7432,N_5726,N_4645);
xnor U7433 (N_7433,N_5386,N_5034);
and U7434 (N_7434,N_5847,N_5805);
or U7435 (N_7435,N_4501,N_5556);
nor U7436 (N_7436,N_4727,N_4933);
or U7437 (N_7437,N_4951,N_5458);
and U7438 (N_7438,N_5099,N_5727);
nor U7439 (N_7439,N_5986,N_4868);
nand U7440 (N_7440,N_5739,N_5196);
xnor U7441 (N_7441,N_5981,N_4821);
and U7442 (N_7442,N_5882,N_4532);
and U7443 (N_7443,N_5694,N_5703);
nand U7444 (N_7444,N_5027,N_5848);
and U7445 (N_7445,N_4914,N_5155);
nand U7446 (N_7446,N_4610,N_5386);
xnor U7447 (N_7447,N_4926,N_4989);
and U7448 (N_7448,N_5451,N_5349);
nand U7449 (N_7449,N_4756,N_5092);
or U7450 (N_7450,N_5230,N_5666);
nand U7451 (N_7451,N_5666,N_4619);
and U7452 (N_7452,N_5475,N_5850);
and U7453 (N_7453,N_4772,N_5151);
nand U7454 (N_7454,N_5685,N_4884);
or U7455 (N_7455,N_5279,N_5298);
and U7456 (N_7456,N_5571,N_4655);
nor U7457 (N_7457,N_5405,N_5169);
nand U7458 (N_7458,N_4522,N_4736);
nand U7459 (N_7459,N_5815,N_5493);
and U7460 (N_7460,N_5117,N_4892);
xnor U7461 (N_7461,N_5022,N_4759);
nor U7462 (N_7462,N_4889,N_5864);
nand U7463 (N_7463,N_4680,N_5387);
or U7464 (N_7464,N_5637,N_5561);
nor U7465 (N_7465,N_4808,N_5976);
xor U7466 (N_7466,N_5999,N_5614);
nand U7467 (N_7467,N_5407,N_5138);
or U7468 (N_7468,N_5265,N_5145);
xnor U7469 (N_7469,N_4911,N_5730);
xnor U7470 (N_7470,N_5684,N_5557);
or U7471 (N_7471,N_5429,N_4782);
and U7472 (N_7472,N_4707,N_4646);
nor U7473 (N_7473,N_5535,N_4567);
nand U7474 (N_7474,N_5962,N_5817);
and U7475 (N_7475,N_4809,N_4836);
nor U7476 (N_7476,N_5359,N_5288);
xor U7477 (N_7477,N_4940,N_5679);
nand U7478 (N_7478,N_4670,N_5927);
nor U7479 (N_7479,N_4827,N_5409);
or U7480 (N_7480,N_5094,N_5381);
nand U7481 (N_7481,N_4500,N_5119);
or U7482 (N_7482,N_5552,N_5272);
nor U7483 (N_7483,N_4749,N_5398);
nand U7484 (N_7484,N_5081,N_5413);
and U7485 (N_7485,N_5063,N_5372);
nand U7486 (N_7486,N_4767,N_4734);
nand U7487 (N_7487,N_4808,N_4950);
xor U7488 (N_7488,N_5718,N_5745);
or U7489 (N_7489,N_5576,N_5268);
nor U7490 (N_7490,N_4820,N_4610);
or U7491 (N_7491,N_5640,N_5002);
nand U7492 (N_7492,N_4992,N_4939);
nor U7493 (N_7493,N_4794,N_5836);
or U7494 (N_7494,N_4800,N_4901);
nor U7495 (N_7495,N_5647,N_4798);
and U7496 (N_7496,N_5475,N_4662);
or U7497 (N_7497,N_5575,N_4891);
nor U7498 (N_7498,N_5683,N_5568);
and U7499 (N_7499,N_5215,N_5362);
and U7500 (N_7500,N_7151,N_6911);
nand U7501 (N_7501,N_7331,N_6881);
xor U7502 (N_7502,N_7213,N_6790);
and U7503 (N_7503,N_7434,N_6666);
or U7504 (N_7504,N_6299,N_6157);
nand U7505 (N_7505,N_6990,N_7405);
and U7506 (N_7506,N_6768,N_7013);
nand U7507 (N_7507,N_6365,N_7252);
nor U7508 (N_7508,N_6786,N_6198);
nor U7509 (N_7509,N_6691,N_6648);
and U7510 (N_7510,N_6285,N_7322);
nor U7511 (N_7511,N_6282,N_7253);
nor U7512 (N_7512,N_6129,N_6572);
xor U7513 (N_7513,N_6701,N_7049);
and U7514 (N_7514,N_6669,N_6578);
and U7515 (N_7515,N_6793,N_6695);
or U7516 (N_7516,N_6671,N_6750);
or U7517 (N_7517,N_6583,N_7468);
nand U7518 (N_7518,N_6661,N_6754);
or U7519 (N_7519,N_6723,N_6022);
and U7520 (N_7520,N_6378,N_7382);
or U7521 (N_7521,N_6110,N_6771);
nor U7522 (N_7522,N_6882,N_7303);
nor U7523 (N_7523,N_7307,N_6773);
or U7524 (N_7524,N_6760,N_6289);
nor U7525 (N_7525,N_7248,N_6354);
nor U7526 (N_7526,N_7163,N_6505);
nand U7527 (N_7527,N_6512,N_6419);
nand U7528 (N_7528,N_6552,N_6788);
nor U7529 (N_7529,N_6872,N_7438);
and U7530 (N_7530,N_7246,N_6561);
xor U7531 (N_7531,N_6761,N_7366);
and U7532 (N_7532,N_7218,N_6167);
and U7533 (N_7533,N_7437,N_7183);
or U7534 (N_7534,N_7420,N_7235);
and U7535 (N_7535,N_6713,N_7141);
nor U7536 (N_7536,N_6966,N_7491);
or U7537 (N_7537,N_6772,N_6919);
nand U7538 (N_7538,N_7068,N_6000);
nand U7539 (N_7539,N_6868,N_6495);
or U7540 (N_7540,N_7374,N_6014);
nor U7541 (N_7541,N_6125,N_7326);
and U7542 (N_7542,N_6465,N_7257);
and U7543 (N_7543,N_7477,N_6392);
nor U7544 (N_7544,N_6267,N_6855);
xor U7545 (N_7545,N_7306,N_7067);
nand U7546 (N_7546,N_7269,N_7217);
nor U7547 (N_7547,N_6448,N_6159);
or U7548 (N_7548,N_7201,N_7011);
and U7549 (N_7549,N_6341,N_6844);
nand U7550 (N_7550,N_6399,N_7277);
or U7551 (N_7551,N_7283,N_6811);
or U7552 (N_7552,N_7056,N_7480);
or U7553 (N_7553,N_6853,N_7138);
xnor U7554 (N_7554,N_6890,N_6080);
or U7555 (N_7555,N_6309,N_6739);
nor U7556 (N_7556,N_6897,N_6953);
nor U7557 (N_7557,N_7202,N_7037);
nand U7558 (N_7558,N_6827,N_6117);
nor U7559 (N_7559,N_6931,N_6209);
and U7560 (N_7560,N_6182,N_6349);
nor U7561 (N_7561,N_6385,N_6049);
and U7562 (N_7562,N_7376,N_6092);
or U7563 (N_7563,N_7146,N_7465);
or U7564 (N_7564,N_6964,N_6412);
or U7565 (N_7565,N_6676,N_6456);
and U7566 (N_7566,N_6837,N_6703);
nand U7567 (N_7567,N_7294,N_6958);
or U7568 (N_7568,N_7057,N_6387);
nand U7569 (N_7569,N_6091,N_6556);
and U7570 (N_7570,N_6704,N_6176);
xor U7571 (N_7571,N_6292,N_6339);
nor U7572 (N_7572,N_7203,N_6943);
xor U7573 (N_7573,N_6698,N_6048);
nor U7574 (N_7574,N_6543,N_6065);
or U7575 (N_7575,N_7044,N_6652);
nor U7576 (N_7576,N_6846,N_6581);
nor U7577 (N_7577,N_6217,N_6122);
and U7578 (N_7578,N_7153,N_6781);
nor U7579 (N_7579,N_6431,N_7476);
nand U7580 (N_7580,N_7221,N_6161);
nor U7581 (N_7581,N_6832,N_6265);
nand U7582 (N_7582,N_6614,N_7096);
nor U7583 (N_7583,N_6900,N_7121);
or U7584 (N_7584,N_6395,N_6276);
or U7585 (N_7585,N_6974,N_6696);
or U7586 (N_7586,N_6109,N_7199);
nor U7587 (N_7587,N_6196,N_7375);
nor U7588 (N_7588,N_6679,N_6765);
nor U7589 (N_7589,N_7337,N_7082);
and U7590 (N_7590,N_7053,N_6440);
nand U7591 (N_7591,N_6263,N_6138);
nor U7592 (N_7592,N_6345,N_6893);
nand U7593 (N_7593,N_6449,N_7267);
or U7594 (N_7594,N_6386,N_6527);
or U7595 (N_7595,N_7394,N_7488);
nor U7596 (N_7596,N_6053,N_7352);
nand U7597 (N_7597,N_6088,N_7159);
and U7598 (N_7598,N_6571,N_6009);
xnor U7599 (N_7599,N_6993,N_6374);
and U7600 (N_7600,N_6221,N_6227);
nand U7601 (N_7601,N_7062,N_6314);
nor U7602 (N_7602,N_6537,N_6938);
and U7603 (N_7603,N_6650,N_7014);
and U7604 (N_7604,N_6797,N_6817);
xnor U7605 (N_7605,N_7169,N_6186);
nand U7606 (N_7606,N_7208,N_7008);
nand U7607 (N_7607,N_7481,N_7220);
or U7608 (N_7608,N_7412,N_7197);
nor U7609 (N_7609,N_6325,N_7418);
and U7610 (N_7610,N_7143,N_6865);
nor U7611 (N_7611,N_6226,N_6123);
nor U7612 (N_7612,N_7441,N_6023);
or U7613 (N_7613,N_7043,N_6904);
or U7614 (N_7614,N_6621,N_6778);
nand U7615 (N_7615,N_6442,N_6158);
nor U7616 (N_7616,N_6540,N_6864);
nor U7617 (N_7617,N_6375,N_7165);
nand U7618 (N_7618,N_6564,N_7264);
nor U7619 (N_7619,N_6798,N_7310);
xor U7620 (N_7620,N_7416,N_6275);
and U7621 (N_7621,N_6028,N_7462);
or U7622 (N_7622,N_7370,N_6601);
nor U7623 (N_7623,N_7009,N_7372);
or U7624 (N_7624,N_7320,N_7410);
or U7625 (N_7625,N_6424,N_7178);
nand U7626 (N_7626,N_6825,N_6428);
nor U7627 (N_7627,N_6469,N_6426);
nor U7628 (N_7628,N_7443,N_6526);
xor U7629 (N_7629,N_6409,N_7098);
nand U7630 (N_7630,N_7212,N_6845);
or U7631 (N_7631,N_6686,N_6052);
nor U7632 (N_7632,N_6178,N_6602);
nor U7633 (N_7633,N_6632,N_7135);
or U7634 (N_7634,N_6434,N_6201);
nor U7635 (N_7635,N_6318,N_6224);
or U7636 (N_7636,N_6905,N_6662);
xnor U7637 (N_7637,N_6004,N_6539);
xnor U7638 (N_7638,N_6241,N_6735);
nor U7639 (N_7639,N_6826,N_7429);
or U7640 (N_7640,N_7432,N_7260);
or U7641 (N_7641,N_7489,N_7229);
nand U7642 (N_7642,N_6690,N_6763);
or U7643 (N_7643,N_6220,N_7373);
nor U7644 (N_7644,N_6383,N_6188);
nand U7645 (N_7645,N_6368,N_6016);
or U7646 (N_7646,N_7099,N_7182);
or U7647 (N_7647,N_7139,N_6940);
nand U7648 (N_7648,N_6749,N_6821);
nor U7649 (N_7649,N_6351,N_6712);
xnor U7650 (N_7650,N_6187,N_7455);
nand U7651 (N_7651,N_6423,N_7118);
or U7652 (N_7652,N_6779,N_7285);
or U7653 (N_7653,N_6233,N_6699);
nor U7654 (N_7654,N_6847,N_6169);
or U7655 (N_7655,N_6170,N_7389);
nand U7656 (N_7656,N_6559,N_6095);
and U7657 (N_7657,N_6906,N_6711);
nand U7658 (N_7658,N_6764,N_6848);
nand U7659 (N_7659,N_6818,N_6271);
nor U7660 (N_7660,N_6758,N_6160);
and U7661 (N_7661,N_6199,N_6590);
nor U7662 (N_7662,N_6421,N_6251);
nand U7663 (N_7663,N_6420,N_6684);
and U7664 (N_7664,N_6076,N_6829);
xor U7665 (N_7665,N_6545,N_6727);
and U7666 (N_7666,N_6631,N_6664);
xor U7667 (N_7667,N_6393,N_6474);
and U7668 (N_7668,N_7150,N_7251);
and U7669 (N_7669,N_6903,N_6099);
nand U7670 (N_7670,N_6247,N_7494);
or U7671 (N_7671,N_7181,N_6618);
nor U7672 (N_7672,N_6101,N_6896);
xnor U7673 (N_7673,N_6784,N_6127);
and U7674 (N_7674,N_7095,N_7238);
nand U7675 (N_7675,N_7194,N_7027);
nor U7676 (N_7676,N_6935,N_6461);
nor U7677 (N_7677,N_6061,N_6946);
nand U7678 (N_7678,N_7454,N_6145);
nand U7679 (N_7679,N_6360,N_6907);
nand U7680 (N_7680,N_6577,N_6926);
and U7681 (N_7681,N_6398,N_7004);
nor U7682 (N_7682,N_7089,N_6432);
nor U7683 (N_7683,N_6370,N_7365);
nand U7684 (N_7684,N_7347,N_6492);
or U7685 (N_7685,N_7002,N_6834);
nor U7686 (N_7686,N_6789,N_7116);
and U7687 (N_7687,N_6457,N_7325);
nand U7688 (N_7688,N_6005,N_7070);
or U7689 (N_7689,N_7256,N_6215);
or U7690 (N_7690,N_7487,N_6291);
nor U7691 (N_7691,N_7423,N_6534);
nor U7692 (N_7692,N_6642,N_6113);
and U7693 (N_7693,N_6525,N_7433);
nand U7694 (N_7694,N_7332,N_6706);
nand U7695 (N_7695,N_7395,N_6249);
xnor U7696 (N_7696,N_6082,N_7399);
nand U7697 (N_7697,N_6154,N_6523);
or U7698 (N_7698,N_7299,N_7396);
or U7699 (N_7699,N_7342,N_6193);
nand U7700 (N_7700,N_6796,N_6979);
nand U7701 (N_7701,N_7234,N_7363);
nor U7702 (N_7702,N_6720,N_6142);
nor U7703 (N_7703,N_6274,N_6530);
and U7704 (N_7704,N_6073,N_6102);
nor U7705 (N_7705,N_6787,N_6453);
nand U7706 (N_7706,N_7362,N_6927);
or U7707 (N_7707,N_7329,N_6210);
nor U7708 (N_7708,N_6433,N_6932);
and U7709 (N_7709,N_7452,N_7401);
nand U7710 (N_7710,N_6565,N_7411);
or U7711 (N_7711,N_7016,N_7078);
and U7712 (N_7712,N_7207,N_7469);
nand U7713 (N_7713,N_6719,N_6260);
xor U7714 (N_7714,N_6230,N_6836);
or U7715 (N_7715,N_6253,N_6619);
nand U7716 (N_7716,N_6327,N_7149);
xnor U7717 (N_7717,N_6783,N_6121);
and U7718 (N_7718,N_7266,N_6767);
and U7719 (N_7719,N_6232,N_6418);
nor U7720 (N_7720,N_6737,N_6438);
and U7721 (N_7721,N_7304,N_7398);
or U7722 (N_7722,N_6566,N_6718);
nand U7723 (N_7723,N_6891,N_7451);
nor U7724 (N_7724,N_6860,N_7247);
and U7725 (N_7725,N_6447,N_6443);
and U7726 (N_7726,N_6298,N_6924);
and U7727 (N_7727,N_6623,N_6155);
and U7728 (N_7728,N_7313,N_7431);
xnor U7729 (N_7729,N_6839,N_7227);
or U7730 (N_7730,N_6002,N_6770);
nand U7731 (N_7731,N_6400,N_6925);
and U7732 (N_7732,N_6501,N_6902);
or U7733 (N_7733,N_6476,N_7426);
or U7734 (N_7734,N_7085,N_6863);
or U7735 (N_7735,N_6639,N_6658);
nand U7736 (N_7736,N_6532,N_7196);
or U7737 (N_7737,N_6672,N_6626);
nand U7738 (N_7738,N_7075,N_7239);
nand U7739 (N_7739,N_7028,N_6963);
nor U7740 (N_7740,N_6394,N_7359);
or U7741 (N_7741,N_7175,N_6384);
and U7742 (N_7742,N_7076,N_7093);
and U7743 (N_7743,N_7367,N_6637);
nand U7744 (N_7744,N_6143,N_6558);
and U7745 (N_7745,N_6549,N_6219);
or U7746 (N_7746,N_6223,N_6777);
and U7747 (N_7747,N_7003,N_7392);
nor U7748 (N_7748,N_6038,N_7161);
and U7749 (N_7749,N_6236,N_6280);
nand U7750 (N_7750,N_6295,N_7343);
nor U7751 (N_7751,N_6544,N_7292);
nor U7752 (N_7752,N_6550,N_6850);
or U7753 (N_7753,N_7327,N_6975);
and U7754 (N_7754,N_6801,N_7258);
and U7755 (N_7755,N_6814,N_6586);
nor U7756 (N_7756,N_7479,N_7496);
nor U7757 (N_7757,N_6522,N_7134);
nand U7758 (N_7758,N_6269,N_7275);
or U7759 (N_7759,N_7409,N_6389);
nand U7760 (N_7760,N_6934,N_7038);
and U7761 (N_7761,N_6311,N_7176);
and U7762 (N_7762,N_6162,N_6111);
and U7763 (N_7763,N_6611,N_6753);
and U7764 (N_7764,N_6063,N_6516);
nand U7765 (N_7765,N_6830,N_6894);
nor U7766 (N_7766,N_7152,N_6415);
nor U7767 (N_7767,N_7147,N_7115);
and U7768 (N_7768,N_7458,N_6876);
nand U7769 (N_7769,N_6008,N_7336);
nor U7770 (N_7770,N_6823,N_7103);
nor U7771 (N_7771,N_7460,N_6211);
or U7772 (N_7772,N_6301,N_7127);
nor U7773 (N_7773,N_7059,N_7400);
or U7774 (N_7774,N_6488,N_7249);
and U7775 (N_7775,N_6659,N_7015);
and U7776 (N_7776,N_6518,N_7309);
nor U7777 (N_7777,N_7225,N_7171);
nand U7778 (N_7778,N_6514,N_7377);
nand U7779 (N_7779,N_6467,N_7271);
nor U7780 (N_7780,N_7066,N_6908);
or U7781 (N_7781,N_6213,N_6264);
or U7782 (N_7782,N_7279,N_6151);
and U7783 (N_7783,N_6745,N_6195);
or U7784 (N_7784,N_6388,N_6283);
xnor U7785 (N_7785,N_6315,N_6910);
xnor U7786 (N_7786,N_6235,N_6948);
nand U7787 (N_7787,N_6597,N_6607);
nor U7788 (N_7788,N_6120,N_7424);
and U7789 (N_7789,N_7334,N_6569);
and U7790 (N_7790,N_6367,N_6744);
nand U7791 (N_7791,N_7284,N_7061);
and U7792 (N_7792,N_6715,N_6736);
or U7793 (N_7793,N_6272,N_6802);
or U7794 (N_7794,N_7348,N_6965);
nor U7795 (N_7795,N_6087,N_6324);
or U7796 (N_7796,N_6281,N_7301);
and U7797 (N_7797,N_6058,N_6775);
and U7798 (N_7798,N_6460,N_7107);
or U7799 (N_7799,N_6104,N_7032);
nand U7800 (N_7800,N_6390,N_6163);
and U7801 (N_7801,N_6687,N_6653);
nor U7802 (N_7802,N_6451,N_6268);
nand U7803 (N_7803,N_6310,N_7200);
or U7804 (N_7804,N_6513,N_6689);
and U7805 (N_7805,N_6654,N_7007);
and U7806 (N_7806,N_6562,N_6870);
and U7807 (N_7807,N_6681,N_7091);
xnor U7808 (N_7808,N_6225,N_6446);
and U7809 (N_7809,N_6321,N_6404);
or U7810 (N_7810,N_6939,N_6057);
xnor U7811 (N_7811,N_6989,N_6616);
xor U7812 (N_7812,N_7064,N_6273);
nand U7813 (N_7813,N_6929,N_6702);
nor U7814 (N_7814,N_6807,N_6084);
nand U7815 (N_7815,N_7498,N_6144);
or U7816 (N_7816,N_7231,N_7210);
nor U7817 (N_7817,N_7162,N_6915);
or U7818 (N_7818,N_7472,N_6857);
nand U7819 (N_7819,N_6785,N_6075);
or U7820 (N_7820,N_7383,N_7020);
and U7821 (N_7821,N_7358,N_6140);
and U7822 (N_7822,N_7485,N_7270);
xor U7823 (N_7823,N_7074,N_6692);
nand U7824 (N_7824,N_6636,N_6175);
or U7825 (N_7825,N_7019,N_7077);
xor U7826 (N_7826,N_7486,N_6520);
or U7827 (N_7827,N_6984,N_6100);
nor U7828 (N_7828,N_6331,N_7110);
xnor U7829 (N_7829,N_6498,N_7447);
and U7830 (N_7830,N_7223,N_6725);
and U7831 (N_7831,N_6304,N_6229);
nor U7832 (N_7832,N_6670,N_6620);
nand U7833 (N_7833,N_7295,N_7349);
nor U7834 (N_7834,N_6531,N_7421);
nand U7835 (N_7835,N_6806,N_7205);
and U7836 (N_7836,N_6307,N_6835);
nand U7837 (N_7837,N_6851,N_6396);
nor U7838 (N_7838,N_6794,N_7224);
nand U7839 (N_7839,N_7189,N_6766);
nand U7840 (N_7840,N_6657,N_6849);
nand U7841 (N_7841,N_6957,N_7330);
and U7842 (N_7842,N_7250,N_7047);
and U7843 (N_7843,N_7177,N_6804);
nand U7844 (N_7844,N_6403,N_7105);
or U7845 (N_7845,N_7195,N_7168);
nor U7846 (N_7846,N_6981,N_7191);
or U7847 (N_7847,N_6665,N_6936);
nand U7848 (N_7848,N_6810,N_7495);
nand U7849 (N_7849,N_6340,N_6694);
xor U7850 (N_7850,N_6485,N_6972);
and U7851 (N_7851,N_6883,N_7404);
or U7852 (N_7852,N_6027,N_6051);
and U7853 (N_7853,N_6463,N_7346);
or U7854 (N_7854,N_6444,N_6098);
nor U7855 (N_7855,N_7351,N_6067);
and U7856 (N_7856,N_7371,N_6730);
nand U7857 (N_7857,N_6494,N_7033);
or U7858 (N_7858,N_6647,N_6477);
and U7859 (N_7859,N_6332,N_6371);
and U7860 (N_7860,N_7393,N_6553);
and U7861 (N_7861,N_6430,N_6576);
or U7862 (N_7862,N_7435,N_6089);
nor U7863 (N_7863,N_6867,N_6279);
nand U7864 (N_7864,N_6490,N_6108);
and U7865 (N_7865,N_7018,N_6288);
and U7866 (N_7866,N_7123,N_6997);
nand U7867 (N_7867,N_6792,N_6046);
nand U7868 (N_7868,N_6885,N_7034);
and U7869 (N_7869,N_6316,N_7474);
and U7870 (N_7870,N_6567,N_6733);
or U7871 (N_7871,N_7272,N_7436);
and U7872 (N_7872,N_6372,N_7132);
nand U7873 (N_7873,N_6959,N_6800);
or U7874 (N_7874,N_6916,N_7364);
and U7875 (N_7875,N_6001,N_6740);
nor U7876 (N_7876,N_7198,N_6093);
nand U7877 (N_7877,N_6776,N_7117);
or U7878 (N_7878,N_7104,N_6563);
nand U7879 (N_7879,N_7324,N_6714);
or U7880 (N_7880,N_6344,N_6751);
and U7881 (N_7881,N_6605,N_7293);
or U7882 (N_7882,N_7108,N_6491);
nor U7883 (N_7883,N_6064,N_6356);
or U7884 (N_7884,N_6017,N_6475);
xnor U7885 (N_7885,N_7154,N_6380);
nor U7886 (N_7886,N_6180,N_7245);
nor U7887 (N_7887,N_6551,N_6560);
nand U7888 (N_7888,N_6007,N_6177);
and U7889 (N_7889,N_7041,N_7164);
and U7890 (N_7890,N_7125,N_7440);
nor U7891 (N_7891,N_6174,N_6697);
xor U7892 (N_7892,N_6606,N_6536);
nand U7893 (N_7893,N_6330,N_7222);
and U7894 (N_7894,N_6252,N_6248);
nor U7895 (N_7895,N_6668,N_6866);
and U7896 (N_7896,N_7386,N_6074);
or U7897 (N_7897,N_6146,N_6244);
xnor U7898 (N_7898,N_6270,N_7054);
nand U7899 (N_7899,N_7006,N_6933);
nand U7900 (N_7900,N_6542,N_6308);
and U7901 (N_7901,N_6838,N_7214);
xnor U7902 (N_7902,N_6573,N_6141);
and U7903 (N_7903,N_6808,N_7471);
nand U7904 (N_7904,N_6585,N_7024);
xor U7905 (N_7905,N_7063,N_6489);
nand U7906 (N_7906,N_6819,N_6326);
or U7907 (N_7907,N_7417,N_6410);
nand U7908 (N_7908,N_6342,N_6886);
nand U7909 (N_7909,N_7022,N_7291);
nor U7910 (N_7910,N_6242,N_7470);
and U7911 (N_7911,N_6171,N_7237);
and U7912 (N_7912,N_7084,N_6239);
xor U7913 (N_7913,N_6427,N_6954);
or U7914 (N_7914,N_7317,N_6930);
or U7915 (N_7915,N_7130,N_6364);
or U7916 (N_7916,N_6651,N_6921);
or U7917 (N_7917,N_6548,N_6094);
nand U7918 (N_7918,N_7157,N_7300);
and U7919 (N_7919,N_7339,N_6312);
nand U7920 (N_7920,N_6589,N_6214);
nand U7921 (N_7921,N_7360,N_6296);
nor U7922 (N_7922,N_7280,N_7296);
and U7923 (N_7923,N_7137,N_6917);
or U7924 (N_7924,N_7287,N_7273);
or U7925 (N_7925,N_6119,N_7345);
nand U7926 (N_7926,N_6204,N_6033);
nor U7927 (N_7927,N_6630,N_6164);
nor U7928 (N_7928,N_6854,N_6624);
nand U7929 (N_7929,N_6976,N_7145);
and U7930 (N_7930,N_7422,N_6960);
or U7931 (N_7931,N_6859,N_6320);
or U7932 (N_7932,N_6509,N_6436);
or U7933 (N_7933,N_6136,N_6728);
or U7934 (N_7934,N_6039,N_6570);
nor U7935 (N_7935,N_7106,N_7158);
and U7936 (N_7936,N_6056,N_6824);
or U7937 (N_7937,N_6638,N_6898);
xor U7938 (N_7938,N_6401,N_6507);
nand U7939 (N_7939,N_6083,N_6153);
nand U7940 (N_7940,N_6502,N_6613);
nand U7941 (N_7941,N_7144,N_6521);
and U7942 (N_7942,N_6391,N_7428);
or U7943 (N_7943,N_6709,N_6300);
and U7944 (N_7944,N_7459,N_7338);
nor U7945 (N_7945,N_6405,N_6337);
xor U7946 (N_7946,N_7188,N_6131);
nor U7947 (N_7947,N_6126,N_6015);
nand U7948 (N_7948,N_6173,N_6708);
nor U7949 (N_7949,N_6366,N_6035);
and U7950 (N_7950,N_6294,N_7023);
nand U7951 (N_7951,N_6018,N_7414);
and U7952 (N_7952,N_6259,N_7088);
xnor U7953 (N_7953,N_6774,N_6203);
nor U7954 (N_7954,N_6257,N_6888);
or U7955 (N_7955,N_6071,N_6899);
nor U7956 (N_7956,N_7219,N_6200);
nor U7957 (N_7957,N_7243,N_6478);
nand U7958 (N_7958,N_7045,N_7478);
and U7959 (N_7959,N_6962,N_6479);
and U7960 (N_7960,N_6471,N_6184);
or U7961 (N_7961,N_6517,N_6435);
nor U7962 (N_7962,N_7354,N_6036);
and U7963 (N_7963,N_6425,N_7052);
xor U7964 (N_7964,N_7397,N_6085);
nor U7965 (N_7965,N_7323,N_6496);
or U7966 (N_7966,N_6944,N_6942);
nor U7967 (N_7967,N_6752,N_6081);
xor U7968 (N_7968,N_6700,N_6947);
or U7969 (N_7969,N_7340,N_6608);
xor U7970 (N_7970,N_7381,N_7005);
and U7971 (N_7971,N_7430,N_6856);
nand U7972 (N_7972,N_6815,N_6041);
nand U7973 (N_7973,N_7119,N_6194);
and U7974 (N_7974,N_6805,N_6166);
nor U7975 (N_7975,N_6013,N_7259);
nor U7976 (N_7976,N_6499,N_7180);
nor U7977 (N_7977,N_6987,N_7456);
nor U7978 (N_7978,N_6887,N_6707);
nand U7979 (N_7979,N_6066,N_6968);
nor U7980 (N_7980,N_6584,N_6493);
and U7981 (N_7981,N_6951,N_7156);
nand U7982 (N_7982,N_6831,N_6515);
or U7983 (N_7983,N_7419,N_6317);
or U7984 (N_7984,N_6667,N_6472);
nand U7985 (N_7985,N_6680,N_7142);
xnor U7986 (N_7986,N_7079,N_6688);
nor U7987 (N_7987,N_6945,N_7000);
nor U7988 (N_7988,N_6216,N_6950);
and U7989 (N_7989,N_6503,N_6413);
and U7990 (N_7990,N_6323,N_6743);
or U7991 (N_7991,N_6192,N_6470);
and U7992 (N_7992,N_7446,N_7262);
or U7993 (N_7993,N_6003,N_7297);
xor U7994 (N_7994,N_6302,N_7328);
and U7995 (N_7995,N_6133,N_7042);
nand U7996 (N_7996,N_6181,N_6971);
nand U7997 (N_7997,N_7211,N_6612);
nor U7998 (N_7998,N_6032,N_6504);
nand U7999 (N_7999,N_6165,N_6646);
or U8000 (N_8000,N_7148,N_6258);
and U8001 (N_8001,N_7333,N_7321);
nor U8002 (N_8002,N_6168,N_6977);
or U8003 (N_8003,N_6486,N_6852);
nand U8004 (N_8004,N_6031,N_7112);
nor U8005 (N_8005,N_6625,N_7390);
nand U8006 (N_8006,N_6742,N_7101);
nand U8007 (N_8007,N_7133,N_6437);
and U8008 (N_8008,N_6574,N_7100);
and U8009 (N_8009,N_6982,N_6114);
and U8010 (N_8010,N_7233,N_6363);
and U8011 (N_8011,N_6190,N_6685);
nor U8012 (N_8012,N_6909,N_6043);
nor U8013 (N_8013,N_6633,N_6617);
and U8014 (N_8014,N_6012,N_7483);
nor U8015 (N_8015,N_6519,N_6615);
nor U8016 (N_8016,N_6290,N_7242);
and U8017 (N_8017,N_6068,N_7318);
nand U8018 (N_8018,N_7427,N_6459);
and U8019 (N_8019,N_7350,N_6955);
nor U8020 (N_8020,N_6635,N_6030);
nor U8021 (N_8021,N_6062,N_6130);
nor U8022 (N_8022,N_6045,N_6988);
and U8023 (N_8023,N_6884,N_7314);
nand U8024 (N_8024,N_6649,N_6949);
or U8025 (N_8025,N_6724,N_6487);
nor U8026 (N_8026,N_7425,N_6928);
and U8027 (N_8027,N_6991,N_6115);
xor U8028 (N_8028,N_6579,N_6877);
and U8029 (N_8029,N_6889,N_7475);
nor U8030 (N_8030,N_6006,N_6970);
and U8031 (N_8031,N_6350,N_7030);
nor U8032 (N_8032,N_6149,N_7206);
or U8033 (N_8033,N_6078,N_6506);
nor U8034 (N_8034,N_7312,N_6529);
xnor U8035 (N_8035,N_6054,N_7391);
or U8036 (N_8036,N_6462,N_6336);
nor U8037 (N_8037,N_7092,N_7001);
and U8038 (N_8038,N_6923,N_6809);
or U8039 (N_8039,N_7261,N_7081);
xnor U8040 (N_8040,N_7450,N_6640);
nand U8041 (N_8041,N_7241,N_6059);
or U8042 (N_8042,N_7129,N_7087);
nand U8043 (N_8043,N_6880,N_6060);
nand U8044 (N_8044,N_7276,N_6622);
nand U8045 (N_8045,N_6246,N_6042);
or U8046 (N_8046,N_6599,N_7492);
xor U8047 (N_8047,N_7356,N_7385);
or U8048 (N_8048,N_6998,N_7482);
nor U8049 (N_8049,N_7069,N_7073);
and U8050 (N_8050,N_6132,N_7228);
xnor U8051 (N_8051,N_7173,N_7124);
nand U8052 (N_8052,N_6875,N_6079);
nor U8053 (N_8053,N_7406,N_7379);
nand U8054 (N_8054,N_7319,N_6254);
and U8055 (N_8055,N_6795,N_7185);
nand U8056 (N_8056,N_6228,N_7473);
nand U8057 (N_8057,N_6357,N_6629);
or U8058 (N_8058,N_6952,N_7466);
and U8059 (N_8059,N_6734,N_6037);
nor U8060 (N_8060,N_6358,N_6705);
xor U8061 (N_8061,N_7216,N_6961);
nand U8062 (N_8062,N_6025,N_6441);
nand U8063 (N_8063,N_6941,N_7344);
nand U8064 (N_8064,N_7449,N_6722);
nor U8065 (N_8065,N_6995,N_7353);
xor U8066 (N_8066,N_6759,N_6450);
nand U8067 (N_8067,N_7120,N_6748);
or U8068 (N_8068,N_6782,N_6841);
nor U8069 (N_8069,N_7268,N_6628);
nor U8070 (N_8070,N_7128,N_6297);
nand U8071 (N_8071,N_6179,N_7413);
or U8072 (N_8072,N_7186,N_7072);
or U8073 (N_8073,N_6197,N_6107);
or U8074 (N_8074,N_6352,N_7226);
nor U8075 (N_8075,N_6417,N_6994);
or U8076 (N_8076,N_6644,N_6677);
and U8077 (N_8077,N_6147,N_7126);
or U8078 (N_8078,N_6746,N_7035);
nand U8079 (N_8079,N_6603,N_7278);
and U8080 (N_8080,N_6922,N_7387);
or U8081 (N_8081,N_7311,N_6338);
nor U8082 (N_8082,N_6077,N_7050);
nand U8083 (N_8083,N_7457,N_6097);
nand U8084 (N_8084,N_6407,N_6124);
nand U8085 (N_8085,N_6445,N_6675);
or U8086 (N_8086,N_7021,N_7467);
and U8087 (N_8087,N_6726,N_6137);
nor U8088 (N_8088,N_6334,N_7240);
nand U8089 (N_8089,N_6710,N_6992);
and U8090 (N_8090,N_7369,N_6020);
or U8091 (N_8091,N_7170,N_7493);
and U8092 (N_8092,N_6547,N_7286);
and U8093 (N_8093,N_7039,N_6816);
or U8094 (N_8094,N_7017,N_6355);
xor U8095 (N_8095,N_6822,N_6050);
and U8096 (N_8096,N_7355,N_6070);
and U8097 (N_8097,N_6918,N_6287);
nor U8098 (N_8098,N_6069,N_6484);
and U8099 (N_8099,N_6382,N_6879);
nand U8100 (N_8100,N_6587,N_7453);
and U8101 (N_8101,N_7179,N_6591);
or U8102 (N_8102,N_7290,N_6483);
and U8103 (N_8103,N_7232,N_6376);
or U8104 (N_8104,N_6634,N_6592);
or U8105 (N_8105,N_7236,N_6105);
nand U8106 (N_8106,N_7281,N_6874);
nor U8107 (N_8107,N_7357,N_6112);
and U8108 (N_8108,N_7302,N_6842);
nand U8109 (N_8109,N_7255,N_6021);
or U8110 (N_8110,N_7408,N_6422);
nor U8111 (N_8111,N_6029,N_6999);
and U8112 (N_8112,N_7361,N_6191);
and U8113 (N_8113,N_6218,N_6118);
nor U8114 (N_8114,N_7174,N_7190);
and U8115 (N_8115,N_6208,N_7097);
nand U8116 (N_8116,N_6359,N_7263);
and U8117 (N_8117,N_6328,N_6156);
nor U8118 (N_8118,N_7113,N_6305);
or U8119 (N_8119,N_6335,N_7060);
nand U8120 (N_8120,N_7071,N_6454);
or U8121 (N_8121,N_7065,N_7445);
nor U8122 (N_8122,N_6497,N_6901);
or U8123 (N_8123,N_7368,N_7388);
and U8124 (N_8124,N_6343,N_6799);
nor U8125 (N_8125,N_6262,N_7442);
and U8126 (N_8126,N_6861,N_6996);
nor U8127 (N_8127,N_6693,N_6980);
or U8128 (N_8128,N_7341,N_7499);
and U8129 (N_8129,N_6481,N_6116);
xnor U8130 (N_8130,N_6044,N_6843);
nor U8131 (N_8131,N_7316,N_7415);
and U8132 (N_8132,N_7090,N_7187);
or U8133 (N_8133,N_7114,N_6261);
and U8134 (N_8134,N_6452,N_6055);
and U8135 (N_8135,N_7254,N_6464);
nor U8136 (N_8136,N_6986,N_6466);
nor U8137 (N_8137,N_6206,N_6813);
xor U8138 (N_8138,N_6245,N_6222);
nor U8139 (N_8139,N_6862,N_7274);
nand U8140 (N_8140,N_7131,N_6554);
and U8141 (N_8141,N_6757,N_6237);
xnor U8142 (N_8142,N_6381,N_6150);
or U8143 (N_8143,N_7497,N_6373);
or U8144 (N_8144,N_6871,N_6369);
or U8145 (N_8145,N_6627,N_6508);
nand U8146 (N_8146,N_6172,N_6546);
nor U8147 (N_8147,N_7192,N_7102);
nand U8148 (N_8148,N_6780,N_6956);
nand U8149 (N_8149,N_6306,N_6303);
and U8150 (N_8150,N_6538,N_6011);
nor U8151 (N_8151,N_6185,N_6973);
nand U8152 (N_8152,N_6482,N_6240);
nand U8153 (N_8153,N_6873,N_6717);
nand U8154 (N_8154,N_6582,N_6912);
or U8155 (N_8155,N_6610,N_6580);
and U8156 (N_8156,N_6769,N_6568);
nand U8157 (N_8157,N_6148,N_6869);
nand U8158 (N_8158,N_6878,N_7166);
nand U8159 (N_8159,N_7380,N_7403);
xor U8160 (N_8160,N_7155,N_6411);
nand U8161 (N_8161,N_6596,N_6402);
or U8162 (N_8162,N_6812,N_6673);
and U8163 (N_8163,N_7378,N_6913);
nand U8164 (N_8164,N_6732,N_6010);
nor U8165 (N_8165,N_6293,N_6683);
nand U8166 (N_8166,N_7461,N_6983);
nor U8167 (N_8167,N_6716,N_6641);
nor U8168 (N_8168,N_6828,N_6019);
nor U8169 (N_8169,N_6346,N_7036);
or U8170 (N_8170,N_7230,N_6643);
nand U8171 (N_8171,N_6655,N_7167);
nor U8172 (N_8172,N_6286,N_6555);
nand U8173 (N_8173,N_7083,N_6152);
nor U8174 (N_8174,N_6353,N_7402);
nor U8175 (N_8175,N_6238,N_6250);
or U8176 (N_8176,N_6920,N_6588);
nor U8177 (N_8177,N_6072,N_6858);
and U8178 (N_8178,N_6212,N_6791);
or U8179 (N_8179,N_7282,N_6439);
xnor U8180 (N_8180,N_6377,N_6598);
and U8181 (N_8181,N_7335,N_6738);
xnor U8182 (N_8182,N_7298,N_6510);
nor U8183 (N_8183,N_6535,N_6595);
nor U8184 (N_8184,N_6895,N_6663);
nor U8185 (N_8185,N_7215,N_6397);
xnor U8186 (N_8186,N_7046,N_7029);
and U8187 (N_8187,N_7010,N_7407);
or U8188 (N_8188,N_7244,N_6284);
or U8189 (N_8189,N_7305,N_6333);
nor U8190 (N_8190,N_6937,N_6034);
and U8191 (N_8191,N_6762,N_6040);
or U8192 (N_8192,N_6967,N_6674);
and U8193 (N_8193,N_6329,N_6557);
nand U8194 (N_8194,N_7055,N_6408);
nor U8195 (N_8195,N_6347,N_6255);
nand U8196 (N_8196,N_6480,N_6406);
nor U8197 (N_8197,N_6645,N_6096);
or U8198 (N_8198,N_7439,N_6820);
nand U8199 (N_8199,N_6234,N_7315);
and U8200 (N_8200,N_6414,N_6277);
and U8201 (N_8201,N_7484,N_6106);
and U8202 (N_8202,N_6090,N_6183);
nor U8203 (N_8203,N_6756,N_6205);
nand U8204 (N_8204,N_6047,N_6243);
or U8205 (N_8205,N_7040,N_6985);
or U8206 (N_8206,N_6207,N_6429);
or U8207 (N_8207,N_6833,N_6511);
nor U8208 (N_8208,N_6528,N_6348);
nor U8209 (N_8209,N_6729,N_6892);
nand U8210 (N_8210,N_7184,N_6473);
and U8211 (N_8211,N_7012,N_7288);
or U8212 (N_8212,N_6202,N_7048);
nor U8213 (N_8213,N_7109,N_7265);
nand U8214 (N_8214,N_6741,N_6914);
nand U8215 (N_8215,N_6604,N_7025);
nand U8216 (N_8216,N_7026,N_6266);
and U8217 (N_8217,N_7051,N_7289);
xor U8218 (N_8218,N_7140,N_7464);
nand U8219 (N_8219,N_7308,N_7111);
xor U8220 (N_8220,N_6575,N_6319);
xnor U8221 (N_8221,N_6416,N_6609);
nand U8222 (N_8222,N_7490,N_6747);
nor U8223 (N_8223,N_6660,N_6455);
and U8224 (N_8224,N_7094,N_6379);
xor U8225 (N_8225,N_6969,N_6458);
nand U8226 (N_8226,N_6231,N_7209);
nor U8227 (N_8227,N_7058,N_6103);
xor U8228 (N_8228,N_7463,N_6682);
nor U8229 (N_8229,N_7204,N_6600);
xnor U8230 (N_8230,N_6755,N_6313);
nand U8231 (N_8231,N_7080,N_6803);
or U8232 (N_8232,N_6468,N_6256);
or U8233 (N_8233,N_6026,N_6541);
and U8234 (N_8234,N_7160,N_6656);
nand U8235 (N_8235,N_6134,N_7172);
and U8236 (N_8236,N_7031,N_6524);
and U8237 (N_8237,N_6678,N_7086);
and U8238 (N_8238,N_6086,N_7193);
or U8239 (N_8239,N_6731,N_7448);
nand U8240 (N_8240,N_6128,N_6533);
or U8241 (N_8241,N_6322,N_6593);
nand U8242 (N_8242,N_6500,N_7122);
xnor U8243 (N_8243,N_7384,N_6721);
xnor U8244 (N_8244,N_6024,N_6189);
nor U8245 (N_8245,N_6840,N_6278);
xnor U8246 (N_8246,N_6978,N_6139);
and U8247 (N_8247,N_6362,N_7136);
and U8248 (N_8248,N_6135,N_7444);
nand U8249 (N_8249,N_6594,N_6361);
and U8250 (N_8250,N_6721,N_6763);
and U8251 (N_8251,N_7131,N_7154);
or U8252 (N_8252,N_7373,N_7413);
and U8253 (N_8253,N_6123,N_6937);
or U8254 (N_8254,N_6062,N_6662);
and U8255 (N_8255,N_7067,N_6902);
and U8256 (N_8256,N_6616,N_6143);
xnor U8257 (N_8257,N_6028,N_6532);
nor U8258 (N_8258,N_7293,N_6530);
nand U8259 (N_8259,N_6558,N_6557);
or U8260 (N_8260,N_6404,N_6136);
and U8261 (N_8261,N_6746,N_7259);
or U8262 (N_8262,N_6764,N_7159);
xor U8263 (N_8263,N_6559,N_6670);
xnor U8264 (N_8264,N_6295,N_7324);
or U8265 (N_8265,N_6609,N_6725);
nand U8266 (N_8266,N_7411,N_7173);
nand U8267 (N_8267,N_7022,N_6192);
nor U8268 (N_8268,N_7416,N_6652);
nor U8269 (N_8269,N_6236,N_6886);
nand U8270 (N_8270,N_7176,N_6329);
nand U8271 (N_8271,N_6760,N_7306);
and U8272 (N_8272,N_6262,N_6898);
nand U8273 (N_8273,N_6398,N_6884);
and U8274 (N_8274,N_6158,N_6315);
and U8275 (N_8275,N_7134,N_6697);
or U8276 (N_8276,N_7489,N_6474);
nand U8277 (N_8277,N_6130,N_6323);
and U8278 (N_8278,N_6722,N_6040);
nand U8279 (N_8279,N_7229,N_6999);
nor U8280 (N_8280,N_7155,N_6077);
and U8281 (N_8281,N_6190,N_6298);
and U8282 (N_8282,N_6744,N_7014);
and U8283 (N_8283,N_6644,N_6519);
or U8284 (N_8284,N_6626,N_7277);
or U8285 (N_8285,N_7480,N_6223);
or U8286 (N_8286,N_6773,N_6657);
nand U8287 (N_8287,N_6428,N_7225);
or U8288 (N_8288,N_6805,N_7413);
or U8289 (N_8289,N_6807,N_6244);
nand U8290 (N_8290,N_7032,N_6620);
nand U8291 (N_8291,N_6321,N_6510);
or U8292 (N_8292,N_7292,N_7148);
or U8293 (N_8293,N_6742,N_7499);
and U8294 (N_8294,N_6356,N_6919);
nor U8295 (N_8295,N_6288,N_7229);
and U8296 (N_8296,N_6957,N_6080);
nor U8297 (N_8297,N_6360,N_6314);
or U8298 (N_8298,N_6312,N_7481);
nor U8299 (N_8299,N_6553,N_6867);
nand U8300 (N_8300,N_7057,N_7095);
and U8301 (N_8301,N_6587,N_7427);
xor U8302 (N_8302,N_7185,N_6129);
xor U8303 (N_8303,N_6094,N_6434);
and U8304 (N_8304,N_6652,N_6049);
and U8305 (N_8305,N_6143,N_6305);
and U8306 (N_8306,N_6731,N_6322);
or U8307 (N_8307,N_6927,N_6647);
and U8308 (N_8308,N_6479,N_7391);
xnor U8309 (N_8309,N_6888,N_6492);
nor U8310 (N_8310,N_6500,N_6277);
nand U8311 (N_8311,N_7208,N_6412);
nor U8312 (N_8312,N_7286,N_6184);
nand U8313 (N_8313,N_6071,N_6827);
and U8314 (N_8314,N_6608,N_7039);
and U8315 (N_8315,N_6972,N_6326);
or U8316 (N_8316,N_7012,N_6093);
nand U8317 (N_8317,N_6247,N_7100);
and U8318 (N_8318,N_6893,N_6054);
or U8319 (N_8319,N_7374,N_6083);
or U8320 (N_8320,N_6736,N_6788);
nor U8321 (N_8321,N_7261,N_7097);
nor U8322 (N_8322,N_6375,N_6847);
nor U8323 (N_8323,N_7430,N_6849);
xor U8324 (N_8324,N_7380,N_7274);
and U8325 (N_8325,N_6290,N_6651);
xor U8326 (N_8326,N_6305,N_6469);
xnor U8327 (N_8327,N_6708,N_6273);
nand U8328 (N_8328,N_6454,N_7300);
xor U8329 (N_8329,N_7219,N_6950);
and U8330 (N_8330,N_6543,N_6457);
nand U8331 (N_8331,N_6546,N_6918);
nand U8332 (N_8332,N_6594,N_6401);
and U8333 (N_8333,N_7418,N_7337);
nor U8334 (N_8334,N_6202,N_7463);
xor U8335 (N_8335,N_7303,N_6288);
nor U8336 (N_8336,N_6182,N_6808);
and U8337 (N_8337,N_6448,N_6249);
and U8338 (N_8338,N_6753,N_6965);
nor U8339 (N_8339,N_7367,N_7229);
and U8340 (N_8340,N_6119,N_6092);
or U8341 (N_8341,N_6053,N_7200);
xor U8342 (N_8342,N_6563,N_6624);
and U8343 (N_8343,N_7407,N_7025);
or U8344 (N_8344,N_6692,N_6061);
and U8345 (N_8345,N_6358,N_7456);
nand U8346 (N_8346,N_6249,N_6142);
and U8347 (N_8347,N_6566,N_6342);
xnor U8348 (N_8348,N_7444,N_6281);
and U8349 (N_8349,N_6187,N_6683);
and U8350 (N_8350,N_7221,N_6592);
nor U8351 (N_8351,N_6613,N_6639);
and U8352 (N_8352,N_6352,N_6683);
nand U8353 (N_8353,N_6460,N_6388);
nor U8354 (N_8354,N_6289,N_6003);
or U8355 (N_8355,N_6716,N_6762);
or U8356 (N_8356,N_6510,N_6434);
or U8357 (N_8357,N_7297,N_6442);
or U8358 (N_8358,N_6056,N_7384);
nand U8359 (N_8359,N_6749,N_7187);
nand U8360 (N_8360,N_6486,N_7426);
nand U8361 (N_8361,N_6005,N_7087);
or U8362 (N_8362,N_6198,N_6408);
or U8363 (N_8363,N_6858,N_6588);
or U8364 (N_8364,N_6490,N_6299);
nor U8365 (N_8365,N_7291,N_7212);
xnor U8366 (N_8366,N_6372,N_6264);
xor U8367 (N_8367,N_6028,N_6603);
xor U8368 (N_8368,N_6060,N_6542);
nor U8369 (N_8369,N_7019,N_7400);
nor U8370 (N_8370,N_7266,N_6090);
and U8371 (N_8371,N_6093,N_6507);
xor U8372 (N_8372,N_6030,N_6252);
nor U8373 (N_8373,N_6021,N_7129);
nand U8374 (N_8374,N_6146,N_7255);
and U8375 (N_8375,N_6079,N_6762);
nand U8376 (N_8376,N_7384,N_6638);
xnor U8377 (N_8377,N_7341,N_6298);
nand U8378 (N_8378,N_6588,N_7478);
and U8379 (N_8379,N_7142,N_6459);
or U8380 (N_8380,N_6266,N_7108);
and U8381 (N_8381,N_7180,N_6205);
or U8382 (N_8382,N_6469,N_6329);
nand U8383 (N_8383,N_7294,N_7459);
and U8384 (N_8384,N_7112,N_6083);
or U8385 (N_8385,N_6642,N_6771);
or U8386 (N_8386,N_6246,N_7164);
nor U8387 (N_8387,N_7473,N_7070);
and U8388 (N_8388,N_6543,N_6763);
xnor U8389 (N_8389,N_6709,N_6560);
xnor U8390 (N_8390,N_6845,N_6809);
and U8391 (N_8391,N_6755,N_6100);
and U8392 (N_8392,N_6697,N_6813);
nand U8393 (N_8393,N_6392,N_6856);
nand U8394 (N_8394,N_6688,N_6449);
xnor U8395 (N_8395,N_6553,N_6140);
nor U8396 (N_8396,N_6639,N_6628);
nor U8397 (N_8397,N_7131,N_7188);
nor U8398 (N_8398,N_6427,N_6650);
nand U8399 (N_8399,N_6787,N_6605);
nor U8400 (N_8400,N_6019,N_7027);
nor U8401 (N_8401,N_7455,N_6858);
and U8402 (N_8402,N_6995,N_6786);
xor U8403 (N_8403,N_6789,N_6721);
and U8404 (N_8404,N_6922,N_7261);
nor U8405 (N_8405,N_6759,N_6483);
nor U8406 (N_8406,N_7232,N_6548);
nor U8407 (N_8407,N_6073,N_6274);
nor U8408 (N_8408,N_7342,N_6284);
or U8409 (N_8409,N_7180,N_6376);
nand U8410 (N_8410,N_6454,N_6966);
or U8411 (N_8411,N_6538,N_6153);
nor U8412 (N_8412,N_7280,N_6595);
nor U8413 (N_8413,N_7042,N_6594);
xor U8414 (N_8414,N_7257,N_6121);
nand U8415 (N_8415,N_7278,N_6567);
nor U8416 (N_8416,N_6750,N_6754);
or U8417 (N_8417,N_6239,N_6377);
nand U8418 (N_8418,N_7168,N_6552);
nor U8419 (N_8419,N_6223,N_6040);
or U8420 (N_8420,N_7158,N_7351);
nor U8421 (N_8421,N_6136,N_6712);
nor U8422 (N_8422,N_7409,N_6103);
and U8423 (N_8423,N_6956,N_7238);
nand U8424 (N_8424,N_6543,N_6675);
or U8425 (N_8425,N_6713,N_6513);
or U8426 (N_8426,N_7443,N_6034);
nand U8427 (N_8427,N_6406,N_6795);
xnor U8428 (N_8428,N_7131,N_6546);
nor U8429 (N_8429,N_6927,N_6905);
nor U8430 (N_8430,N_7207,N_6919);
nor U8431 (N_8431,N_6002,N_6371);
or U8432 (N_8432,N_6490,N_6156);
nor U8433 (N_8433,N_6085,N_6327);
or U8434 (N_8434,N_6123,N_6101);
nand U8435 (N_8435,N_7172,N_7193);
and U8436 (N_8436,N_6874,N_6658);
and U8437 (N_8437,N_6058,N_6042);
nand U8438 (N_8438,N_6387,N_7282);
nand U8439 (N_8439,N_6708,N_7323);
nand U8440 (N_8440,N_7146,N_6094);
or U8441 (N_8441,N_7295,N_6420);
nor U8442 (N_8442,N_6260,N_7269);
nand U8443 (N_8443,N_6727,N_7191);
nand U8444 (N_8444,N_7249,N_6550);
or U8445 (N_8445,N_7295,N_6436);
and U8446 (N_8446,N_6232,N_6576);
nor U8447 (N_8447,N_6715,N_6766);
nand U8448 (N_8448,N_6803,N_6625);
or U8449 (N_8449,N_6373,N_6120);
or U8450 (N_8450,N_6739,N_6332);
nor U8451 (N_8451,N_7192,N_6310);
nor U8452 (N_8452,N_6635,N_7238);
nor U8453 (N_8453,N_7093,N_6862);
xor U8454 (N_8454,N_6164,N_6421);
nor U8455 (N_8455,N_6177,N_7349);
nand U8456 (N_8456,N_6870,N_6551);
or U8457 (N_8457,N_6965,N_7240);
nand U8458 (N_8458,N_7129,N_7231);
nor U8459 (N_8459,N_6057,N_7493);
or U8460 (N_8460,N_6456,N_6793);
nand U8461 (N_8461,N_7248,N_6818);
nor U8462 (N_8462,N_6758,N_6429);
xnor U8463 (N_8463,N_6504,N_6477);
xnor U8464 (N_8464,N_6671,N_6037);
or U8465 (N_8465,N_7169,N_6602);
and U8466 (N_8466,N_6808,N_6924);
nor U8467 (N_8467,N_7276,N_6821);
nand U8468 (N_8468,N_6130,N_6366);
xnor U8469 (N_8469,N_6790,N_6603);
and U8470 (N_8470,N_6283,N_6088);
xor U8471 (N_8471,N_7177,N_6460);
or U8472 (N_8472,N_6593,N_6960);
nand U8473 (N_8473,N_6450,N_7377);
or U8474 (N_8474,N_6839,N_7019);
or U8475 (N_8475,N_6218,N_6772);
or U8476 (N_8476,N_6988,N_6513);
or U8477 (N_8477,N_6917,N_6571);
nor U8478 (N_8478,N_6186,N_6651);
or U8479 (N_8479,N_7027,N_6037);
or U8480 (N_8480,N_6786,N_7364);
nand U8481 (N_8481,N_6899,N_6296);
nor U8482 (N_8482,N_6258,N_6642);
nand U8483 (N_8483,N_7091,N_6312);
nor U8484 (N_8484,N_6709,N_7414);
nand U8485 (N_8485,N_6040,N_7170);
and U8486 (N_8486,N_7341,N_6508);
nand U8487 (N_8487,N_6598,N_6574);
nand U8488 (N_8488,N_6366,N_7382);
nand U8489 (N_8489,N_7255,N_7352);
nor U8490 (N_8490,N_6621,N_6117);
and U8491 (N_8491,N_6922,N_6826);
or U8492 (N_8492,N_6031,N_6375);
nand U8493 (N_8493,N_7134,N_6020);
nor U8494 (N_8494,N_6042,N_6932);
or U8495 (N_8495,N_7485,N_6431);
nor U8496 (N_8496,N_7010,N_6697);
and U8497 (N_8497,N_6822,N_6135);
and U8498 (N_8498,N_6663,N_6244);
nor U8499 (N_8499,N_6526,N_6919);
or U8500 (N_8500,N_6730,N_7314);
nor U8501 (N_8501,N_6830,N_6680);
and U8502 (N_8502,N_6851,N_6437);
nor U8503 (N_8503,N_6135,N_6677);
and U8504 (N_8504,N_7104,N_6482);
nor U8505 (N_8505,N_7124,N_6377);
nand U8506 (N_8506,N_6830,N_7276);
and U8507 (N_8507,N_7202,N_7419);
nor U8508 (N_8508,N_7060,N_7140);
and U8509 (N_8509,N_7138,N_7465);
and U8510 (N_8510,N_6462,N_6712);
and U8511 (N_8511,N_6465,N_7275);
nand U8512 (N_8512,N_7079,N_6457);
or U8513 (N_8513,N_6929,N_6707);
nand U8514 (N_8514,N_6862,N_6129);
xnor U8515 (N_8515,N_7414,N_7128);
nor U8516 (N_8516,N_6614,N_7495);
or U8517 (N_8517,N_7171,N_6699);
or U8518 (N_8518,N_6407,N_6942);
or U8519 (N_8519,N_7322,N_7111);
or U8520 (N_8520,N_6404,N_6332);
or U8521 (N_8521,N_6285,N_6598);
nand U8522 (N_8522,N_6522,N_6197);
nand U8523 (N_8523,N_7478,N_6728);
or U8524 (N_8524,N_6456,N_6472);
nor U8525 (N_8525,N_6406,N_6947);
and U8526 (N_8526,N_6151,N_6970);
or U8527 (N_8527,N_6901,N_7451);
or U8528 (N_8528,N_6070,N_6379);
and U8529 (N_8529,N_6396,N_7227);
or U8530 (N_8530,N_7421,N_6444);
or U8531 (N_8531,N_6671,N_6393);
nand U8532 (N_8532,N_6913,N_6800);
nand U8533 (N_8533,N_7354,N_7487);
or U8534 (N_8534,N_6917,N_6606);
and U8535 (N_8535,N_6262,N_6999);
nand U8536 (N_8536,N_7065,N_6175);
xnor U8537 (N_8537,N_6648,N_7107);
or U8538 (N_8538,N_6554,N_6369);
nand U8539 (N_8539,N_7329,N_7336);
nor U8540 (N_8540,N_7354,N_6558);
nor U8541 (N_8541,N_6756,N_7474);
nand U8542 (N_8542,N_6571,N_6370);
nand U8543 (N_8543,N_7497,N_6657);
xnor U8544 (N_8544,N_6481,N_6431);
nand U8545 (N_8545,N_6327,N_6507);
nor U8546 (N_8546,N_6450,N_6356);
nor U8547 (N_8547,N_6168,N_6149);
or U8548 (N_8548,N_6555,N_6208);
nor U8549 (N_8549,N_7358,N_6787);
or U8550 (N_8550,N_7197,N_6725);
nor U8551 (N_8551,N_6054,N_6204);
nand U8552 (N_8552,N_6631,N_6795);
and U8553 (N_8553,N_6942,N_7057);
nor U8554 (N_8554,N_6901,N_6728);
and U8555 (N_8555,N_6562,N_6760);
nand U8556 (N_8556,N_6341,N_6949);
nor U8557 (N_8557,N_6412,N_7151);
or U8558 (N_8558,N_6334,N_6096);
or U8559 (N_8559,N_6423,N_6178);
nor U8560 (N_8560,N_7350,N_6032);
or U8561 (N_8561,N_7029,N_6681);
nor U8562 (N_8562,N_6191,N_7091);
nor U8563 (N_8563,N_6423,N_6847);
and U8564 (N_8564,N_7089,N_6438);
and U8565 (N_8565,N_6586,N_7348);
nand U8566 (N_8566,N_6333,N_6318);
or U8567 (N_8567,N_6852,N_6533);
or U8568 (N_8568,N_6507,N_6508);
and U8569 (N_8569,N_6147,N_6296);
or U8570 (N_8570,N_6046,N_6339);
nor U8571 (N_8571,N_6157,N_6824);
and U8572 (N_8572,N_6150,N_6667);
nor U8573 (N_8573,N_6501,N_6058);
and U8574 (N_8574,N_7339,N_6894);
nand U8575 (N_8575,N_6846,N_7452);
and U8576 (N_8576,N_6259,N_6544);
and U8577 (N_8577,N_6158,N_6445);
xor U8578 (N_8578,N_7159,N_7115);
or U8579 (N_8579,N_7049,N_6037);
nand U8580 (N_8580,N_6744,N_7126);
nand U8581 (N_8581,N_6954,N_7454);
nand U8582 (N_8582,N_6331,N_7056);
nor U8583 (N_8583,N_7331,N_7445);
nand U8584 (N_8584,N_7206,N_7236);
nor U8585 (N_8585,N_6907,N_7105);
or U8586 (N_8586,N_6470,N_6207);
nand U8587 (N_8587,N_6346,N_6507);
and U8588 (N_8588,N_6310,N_6687);
xor U8589 (N_8589,N_7357,N_6100);
nor U8590 (N_8590,N_6020,N_7381);
nor U8591 (N_8591,N_7293,N_6355);
and U8592 (N_8592,N_6882,N_6544);
xnor U8593 (N_8593,N_6703,N_6150);
nand U8594 (N_8594,N_6131,N_7339);
nand U8595 (N_8595,N_6975,N_7145);
nand U8596 (N_8596,N_6357,N_6254);
nor U8597 (N_8597,N_6334,N_6202);
xnor U8598 (N_8598,N_7070,N_6369);
or U8599 (N_8599,N_7340,N_7215);
or U8600 (N_8600,N_6322,N_6455);
and U8601 (N_8601,N_7275,N_6259);
and U8602 (N_8602,N_7465,N_6090);
and U8603 (N_8603,N_7369,N_7491);
or U8604 (N_8604,N_6829,N_6625);
nand U8605 (N_8605,N_6647,N_6021);
xor U8606 (N_8606,N_6331,N_6319);
or U8607 (N_8607,N_6247,N_7409);
nand U8608 (N_8608,N_7269,N_7161);
nand U8609 (N_8609,N_6778,N_7376);
and U8610 (N_8610,N_7255,N_6064);
nor U8611 (N_8611,N_6379,N_7340);
nand U8612 (N_8612,N_7020,N_7260);
nor U8613 (N_8613,N_6087,N_6952);
or U8614 (N_8614,N_7342,N_6111);
nand U8615 (N_8615,N_6426,N_6937);
nand U8616 (N_8616,N_6580,N_6699);
nand U8617 (N_8617,N_6621,N_7019);
xnor U8618 (N_8618,N_6902,N_7405);
nand U8619 (N_8619,N_6574,N_7449);
xnor U8620 (N_8620,N_6886,N_7364);
and U8621 (N_8621,N_7380,N_7493);
or U8622 (N_8622,N_7299,N_7140);
or U8623 (N_8623,N_6285,N_6874);
nand U8624 (N_8624,N_6083,N_6934);
nand U8625 (N_8625,N_6800,N_6433);
and U8626 (N_8626,N_7287,N_6575);
or U8627 (N_8627,N_6939,N_6924);
nand U8628 (N_8628,N_7280,N_7438);
or U8629 (N_8629,N_6151,N_6443);
and U8630 (N_8630,N_7061,N_7286);
and U8631 (N_8631,N_7316,N_6496);
or U8632 (N_8632,N_7074,N_7358);
nor U8633 (N_8633,N_6863,N_7186);
nand U8634 (N_8634,N_6742,N_6930);
or U8635 (N_8635,N_6422,N_7164);
or U8636 (N_8636,N_6265,N_6054);
xnor U8637 (N_8637,N_7416,N_6332);
nor U8638 (N_8638,N_7439,N_7199);
or U8639 (N_8639,N_6661,N_6371);
nand U8640 (N_8640,N_6402,N_6103);
nor U8641 (N_8641,N_7422,N_6678);
and U8642 (N_8642,N_7072,N_6170);
and U8643 (N_8643,N_7105,N_6669);
nand U8644 (N_8644,N_6369,N_7094);
or U8645 (N_8645,N_7406,N_7059);
or U8646 (N_8646,N_7281,N_6651);
nor U8647 (N_8647,N_6418,N_6904);
nor U8648 (N_8648,N_6695,N_7204);
nor U8649 (N_8649,N_6406,N_6660);
nor U8650 (N_8650,N_6958,N_6753);
or U8651 (N_8651,N_6165,N_6900);
nor U8652 (N_8652,N_6467,N_6607);
nor U8653 (N_8653,N_6263,N_6513);
nor U8654 (N_8654,N_6785,N_7364);
nor U8655 (N_8655,N_6307,N_6230);
nor U8656 (N_8656,N_7304,N_7107);
nor U8657 (N_8657,N_6344,N_6716);
and U8658 (N_8658,N_6855,N_6960);
nor U8659 (N_8659,N_7400,N_7341);
and U8660 (N_8660,N_6910,N_7439);
nand U8661 (N_8661,N_6084,N_7037);
nand U8662 (N_8662,N_6911,N_6535);
nor U8663 (N_8663,N_7424,N_7409);
and U8664 (N_8664,N_6493,N_7042);
nand U8665 (N_8665,N_7063,N_7005);
nand U8666 (N_8666,N_6286,N_7161);
or U8667 (N_8667,N_7473,N_7007);
nand U8668 (N_8668,N_6733,N_6933);
nand U8669 (N_8669,N_6820,N_7193);
and U8670 (N_8670,N_7417,N_6379);
and U8671 (N_8671,N_6675,N_6115);
and U8672 (N_8672,N_6597,N_6975);
xnor U8673 (N_8673,N_6356,N_7016);
and U8674 (N_8674,N_7443,N_7262);
nand U8675 (N_8675,N_6100,N_6749);
nand U8676 (N_8676,N_6443,N_6992);
and U8677 (N_8677,N_6135,N_6371);
nor U8678 (N_8678,N_7465,N_7441);
and U8679 (N_8679,N_7160,N_6566);
nand U8680 (N_8680,N_6644,N_6498);
and U8681 (N_8681,N_6174,N_6004);
nand U8682 (N_8682,N_7073,N_6076);
nor U8683 (N_8683,N_6747,N_6446);
nand U8684 (N_8684,N_7381,N_7015);
nand U8685 (N_8685,N_7030,N_6010);
and U8686 (N_8686,N_7269,N_6969);
or U8687 (N_8687,N_6417,N_7096);
and U8688 (N_8688,N_6868,N_6847);
nand U8689 (N_8689,N_7267,N_7105);
nand U8690 (N_8690,N_6857,N_6207);
nor U8691 (N_8691,N_6642,N_6427);
nor U8692 (N_8692,N_6311,N_6384);
or U8693 (N_8693,N_6670,N_6654);
and U8694 (N_8694,N_6929,N_6118);
and U8695 (N_8695,N_7390,N_6165);
nand U8696 (N_8696,N_6319,N_6896);
nor U8697 (N_8697,N_6729,N_6947);
nor U8698 (N_8698,N_6015,N_7032);
or U8699 (N_8699,N_7020,N_6884);
and U8700 (N_8700,N_6111,N_6662);
xnor U8701 (N_8701,N_6517,N_7116);
or U8702 (N_8702,N_6480,N_7266);
or U8703 (N_8703,N_6208,N_6394);
nand U8704 (N_8704,N_6392,N_7177);
nor U8705 (N_8705,N_6021,N_6166);
nand U8706 (N_8706,N_7488,N_7170);
and U8707 (N_8707,N_6362,N_6198);
and U8708 (N_8708,N_6184,N_7086);
and U8709 (N_8709,N_6883,N_7065);
nor U8710 (N_8710,N_6797,N_7083);
nor U8711 (N_8711,N_7220,N_7260);
nor U8712 (N_8712,N_6645,N_6489);
xor U8713 (N_8713,N_6292,N_6456);
nor U8714 (N_8714,N_6760,N_7238);
nand U8715 (N_8715,N_6145,N_6674);
and U8716 (N_8716,N_6527,N_6651);
nor U8717 (N_8717,N_7004,N_6934);
and U8718 (N_8718,N_7149,N_7460);
nand U8719 (N_8719,N_6668,N_7254);
nand U8720 (N_8720,N_6040,N_6891);
or U8721 (N_8721,N_6644,N_7009);
xor U8722 (N_8722,N_7316,N_6176);
xnor U8723 (N_8723,N_7449,N_6891);
and U8724 (N_8724,N_7260,N_6805);
nor U8725 (N_8725,N_6154,N_7388);
and U8726 (N_8726,N_6795,N_7063);
and U8727 (N_8727,N_6927,N_6708);
or U8728 (N_8728,N_6261,N_7349);
nand U8729 (N_8729,N_6170,N_7033);
or U8730 (N_8730,N_6259,N_7238);
nand U8731 (N_8731,N_6636,N_6836);
nor U8732 (N_8732,N_6442,N_6426);
nand U8733 (N_8733,N_6444,N_6831);
or U8734 (N_8734,N_6953,N_6116);
nor U8735 (N_8735,N_6630,N_6824);
nand U8736 (N_8736,N_6469,N_6975);
nand U8737 (N_8737,N_6246,N_6229);
nand U8738 (N_8738,N_6216,N_6263);
and U8739 (N_8739,N_6059,N_6325);
and U8740 (N_8740,N_6037,N_7362);
nand U8741 (N_8741,N_6248,N_6124);
nor U8742 (N_8742,N_7397,N_6998);
or U8743 (N_8743,N_6351,N_6349);
nand U8744 (N_8744,N_6304,N_7002);
or U8745 (N_8745,N_7455,N_6476);
nand U8746 (N_8746,N_7434,N_6427);
xor U8747 (N_8747,N_6377,N_7383);
nor U8748 (N_8748,N_6114,N_7498);
nor U8749 (N_8749,N_7386,N_6452);
or U8750 (N_8750,N_7249,N_7095);
and U8751 (N_8751,N_7373,N_6453);
xnor U8752 (N_8752,N_7091,N_6136);
nand U8753 (N_8753,N_6486,N_6487);
and U8754 (N_8754,N_6718,N_7281);
nor U8755 (N_8755,N_6210,N_6018);
nor U8756 (N_8756,N_6842,N_6020);
nand U8757 (N_8757,N_7289,N_6053);
and U8758 (N_8758,N_7354,N_7311);
or U8759 (N_8759,N_7391,N_6648);
nand U8760 (N_8760,N_7051,N_7307);
nor U8761 (N_8761,N_6815,N_7176);
xnor U8762 (N_8762,N_6112,N_6360);
and U8763 (N_8763,N_6338,N_6573);
or U8764 (N_8764,N_6000,N_7005);
nand U8765 (N_8765,N_6848,N_6183);
and U8766 (N_8766,N_6019,N_6484);
nor U8767 (N_8767,N_7173,N_7061);
or U8768 (N_8768,N_7046,N_6704);
and U8769 (N_8769,N_6664,N_7443);
xor U8770 (N_8770,N_7270,N_6171);
and U8771 (N_8771,N_7044,N_6078);
nand U8772 (N_8772,N_6644,N_6521);
and U8773 (N_8773,N_6402,N_7233);
and U8774 (N_8774,N_6532,N_6301);
nor U8775 (N_8775,N_7331,N_7148);
nand U8776 (N_8776,N_6396,N_6199);
nand U8777 (N_8777,N_6280,N_6935);
xnor U8778 (N_8778,N_6619,N_6564);
and U8779 (N_8779,N_6746,N_6410);
or U8780 (N_8780,N_6805,N_6929);
nand U8781 (N_8781,N_6685,N_6035);
nand U8782 (N_8782,N_6063,N_6687);
nor U8783 (N_8783,N_6281,N_6104);
nand U8784 (N_8784,N_6331,N_6901);
nand U8785 (N_8785,N_6397,N_6962);
and U8786 (N_8786,N_6692,N_7223);
xnor U8787 (N_8787,N_7446,N_6677);
nor U8788 (N_8788,N_6554,N_7411);
and U8789 (N_8789,N_6987,N_6274);
nor U8790 (N_8790,N_6037,N_7377);
nor U8791 (N_8791,N_6078,N_6375);
and U8792 (N_8792,N_6877,N_6285);
nor U8793 (N_8793,N_7490,N_6084);
xnor U8794 (N_8794,N_6410,N_7270);
nand U8795 (N_8795,N_6607,N_6097);
nand U8796 (N_8796,N_6000,N_7056);
nor U8797 (N_8797,N_7046,N_7097);
nor U8798 (N_8798,N_6793,N_6067);
nand U8799 (N_8799,N_6704,N_7056);
nand U8800 (N_8800,N_6861,N_6485);
xnor U8801 (N_8801,N_6286,N_6199);
nor U8802 (N_8802,N_6564,N_6271);
xor U8803 (N_8803,N_7470,N_6906);
nor U8804 (N_8804,N_7328,N_7096);
nand U8805 (N_8805,N_6447,N_7128);
nor U8806 (N_8806,N_6865,N_7305);
and U8807 (N_8807,N_7286,N_7250);
or U8808 (N_8808,N_6709,N_6175);
nor U8809 (N_8809,N_6102,N_6561);
nor U8810 (N_8810,N_6087,N_7098);
or U8811 (N_8811,N_7190,N_6532);
or U8812 (N_8812,N_6431,N_7002);
nor U8813 (N_8813,N_7026,N_6569);
nor U8814 (N_8814,N_6984,N_7094);
nand U8815 (N_8815,N_6135,N_6465);
nor U8816 (N_8816,N_7497,N_6691);
nand U8817 (N_8817,N_6887,N_6525);
nand U8818 (N_8818,N_6564,N_6536);
or U8819 (N_8819,N_6306,N_6256);
nor U8820 (N_8820,N_7111,N_6522);
and U8821 (N_8821,N_6093,N_7098);
nand U8822 (N_8822,N_6741,N_7179);
and U8823 (N_8823,N_6087,N_7029);
nand U8824 (N_8824,N_7452,N_6462);
or U8825 (N_8825,N_6620,N_6183);
nor U8826 (N_8826,N_6192,N_6351);
nand U8827 (N_8827,N_7268,N_6705);
nand U8828 (N_8828,N_6783,N_6419);
nor U8829 (N_8829,N_6935,N_6326);
xor U8830 (N_8830,N_7177,N_6082);
xor U8831 (N_8831,N_7353,N_6797);
and U8832 (N_8832,N_6184,N_6655);
nand U8833 (N_8833,N_6123,N_6846);
and U8834 (N_8834,N_7047,N_7256);
nor U8835 (N_8835,N_7042,N_6942);
and U8836 (N_8836,N_6791,N_6668);
and U8837 (N_8837,N_7243,N_7180);
or U8838 (N_8838,N_6928,N_7487);
and U8839 (N_8839,N_6301,N_7376);
nand U8840 (N_8840,N_6810,N_7397);
xor U8841 (N_8841,N_6485,N_6199);
nand U8842 (N_8842,N_6869,N_7043);
or U8843 (N_8843,N_6484,N_6597);
nor U8844 (N_8844,N_6492,N_6608);
or U8845 (N_8845,N_7489,N_7396);
nand U8846 (N_8846,N_6262,N_7482);
xor U8847 (N_8847,N_7414,N_7280);
or U8848 (N_8848,N_6995,N_6506);
or U8849 (N_8849,N_7316,N_7210);
xnor U8850 (N_8850,N_6506,N_6226);
or U8851 (N_8851,N_6334,N_6652);
or U8852 (N_8852,N_6366,N_7209);
nand U8853 (N_8853,N_6370,N_6553);
nand U8854 (N_8854,N_6950,N_7246);
nor U8855 (N_8855,N_7287,N_7007);
nor U8856 (N_8856,N_6691,N_7005);
or U8857 (N_8857,N_6145,N_6825);
nand U8858 (N_8858,N_6488,N_6105);
nand U8859 (N_8859,N_7352,N_6969);
nand U8860 (N_8860,N_6711,N_6816);
xnor U8861 (N_8861,N_6625,N_6950);
and U8862 (N_8862,N_6008,N_6703);
and U8863 (N_8863,N_6564,N_6360);
xor U8864 (N_8864,N_7202,N_6720);
nor U8865 (N_8865,N_6306,N_6723);
and U8866 (N_8866,N_7140,N_7213);
xnor U8867 (N_8867,N_7448,N_6269);
nand U8868 (N_8868,N_6824,N_7288);
or U8869 (N_8869,N_6466,N_7432);
nand U8870 (N_8870,N_6945,N_6454);
nand U8871 (N_8871,N_6539,N_6492);
nand U8872 (N_8872,N_6563,N_6981);
and U8873 (N_8873,N_7253,N_6720);
or U8874 (N_8874,N_6733,N_7245);
nor U8875 (N_8875,N_6087,N_6145);
xnor U8876 (N_8876,N_7006,N_6898);
nor U8877 (N_8877,N_6902,N_7476);
nor U8878 (N_8878,N_6488,N_6780);
nand U8879 (N_8879,N_6943,N_6373);
nand U8880 (N_8880,N_6956,N_6816);
nand U8881 (N_8881,N_7075,N_6482);
nand U8882 (N_8882,N_6561,N_7275);
nor U8883 (N_8883,N_6859,N_6075);
nor U8884 (N_8884,N_7468,N_6202);
nand U8885 (N_8885,N_7248,N_6742);
or U8886 (N_8886,N_6362,N_6858);
or U8887 (N_8887,N_6226,N_6899);
nor U8888 (N_8888,N_6211,N_6278);
nand U8889 (N_8889,N_6247,N_7264);
and U8890 (N_8890,N_6350,N_6660);
nand U8891 (N_8891,N_6985,N_6101);
nor U8892 (N_8892,N_6785,N_6431);
xnor U8893 (N_8893,N_6237,N_6441);
or U8894 (N_8894,N_7413,N_6004);
and U8895 (N_8895,N_6403,N_6370);
and U8896 (N_8896,N_6142,N_7331);
and U8897 (N_8897,N_6147,N_7278);
nand U8898 (N_8898,N_6589,N_6269);
nand U8899 (N_8899,N_6799,N_7001);
nor U8900 (N_8900,N_6570,N_6809);
nand U8901 (N_8901,N_6539,N_6858);
nor U8902 (N_8902,N_6341,N_6007);
nand U8903 (N_8903,N_6694,N_6271);
and U8904 (N_8904,N_6873,N_6613);
or U8905 (N_8905,N_7201,N_6236);
nand U8906 (N_8906,N_6287,N_6225);
nand U8907 (N_8907,N_6113,N_6643);
or U8908 (N_8908,N_6416,N_7027);
and U8909 (N_8909,N_6031,N_6277);
xor U8910 (N_8910,N_6481,N_7343);
nand U8911 (N_8911,N_6086,N_7183);
nand U8912 (N_8912,N_7025,N_6753);
xnor U8913 (N_8913,N_6139,N_6584);
and U8914 (N_8914,N_6253,N_6079);
and U8915 (N_8915,N_6723,N_6864);
nor U8916 (N_8916,N_6284,N_6646);
or U8917 (N_8917,N_6579,N_6146);
nand U8918 (N_8918,N_6072,N_7248);
or U8919 (N_8919,N_6282,N_7185);
or U8920 (N_8920,N_6744,N_6325);
and U8921 (N_8921,N_6522,N_7477);
and U8922 (N_8922,N_6146,N_7045);
or U8923 (N_8923,N_7138,N_6902);
and U8924 (N_8924,N_6603,N_6438);
xor U8925 (N_8925,N_6090,N_6259);
nor U8926 (N_8926,N_7357,N_6350);
and U8927 (N_8927,N_6100,N_7028);
xnor U8928 (N_8928,N_7169,N_6017);
xor U8929 (N_8929,N_6215,N_7483);
nand U8930 (N_8930,N_6352,N_6210);
nand U8931 (N_8931,N_6151,N_6653);
nor U8932 (N_8932,N_6155,N_7064);
xnor U8933 (N_8933,N_6319,N_6723);
or U8934 (N_8934,N_6765,N_6808);
and U8935 (N_8935,N_7263,N_7402);
or U8936 (N_8936,N_7384,N_6028);
and U8937 (N_8937,N_7477,N_6396);
nand U8938 (N_8938,N_6919,N_6296);
and U8939 (N_8939,N_6552,N_7169);
or U8940 (N_8940,N_6221,N_6984);
nand U8941 (N_8941,N_6101,N_7326);
nor U8942 (N_8942,N_6138,N_7369);
and U8943 (N_8943,N_6644,N_6985);
xnor U8944 (N_8944,N_6275,N_7455);
nor U8945 (N_8945,N_7442,N_7107);
nor U8946 (N_8946,N_6725,N_6693);
and U8947 (N_8947,N_6343,N_7148);
nand U8948 (N_8948,N_6504,N_7485);
nor U8949 (N_8949,N_6316,N_6021);
or U8950 (N_8950,N_7424,N_6772);
or U8951 (N_8951,N_6984,N_6502);
and U8952 (N_8952,N_6604,N_6484);
and U8953 (N_8953,N_7019,N_7405);
nand U8954 (N_8954,N_6662,N_6151);
nor U8955 (N_8955,N_6205,N_6718);
or U8956 (N_8956,N_6425,N_6441);
nor U8957 (N_8957,N_6299,N_6815);
nand U8958 (N_8958,N_6235,N_6393);
nor U8959 (N_8959,N_6313,N_7222);
nand U8960 (N_8960,N_6816,N_6748);
nor U8961 (N_8961,N_6356,N_7028);
nor U8962 (N_8962,N_7219,N_6318);
nand U8963 (N_8963,N_6097,N_7262);
or U8964 (N_8964,N_6872,N_7230);
nor U8965 (N_8965,N_6636,N_7389);
or U8966 (N_8966,N_6394,N_6577);
and U8967 (N_8967,N_7260,N_6798);
and U8968 (N_8968,N_7413,N_6057);
or U8969 (N_8969,N_6616,N_6337);
xor U8970 (N_8970,N_6268,N_6058);
nor U8971 (N_8971,N_6124,N_6743);
and U8972 (N_8972,N_6241,N_7297);
nor U8973 (N_8973,N_7385,N_6686);
nor U8974 (N_8974,N_7121,N_6222);
or U8975 (N_8975,N_6026,N_6947);
nor U8976 (N_8976,N_6364,N_7447);
and U8977 (N_8977,N_6787,N_6651);
nand U8978 (N_8978,N_6603,N_6407);
nor U8979 (N_8979,N_6144,N_6133);
or U8980 (N_8980,N_6468,N_6235);
xnor U8981 (N_8981,N_6876,N_6463);
nor U8982 (N_8982,N_6942,N_6255);
nor U8983 (N_8983,N_7465,N_6739);
nor U8984 (N_8984,N_7440,N_6354);
nand U8985 (N_8985,N_6491,N_6385);
and U8986 (N_8986,N_7346,N_6631);
xor U8987 (N_8987,N_7444,N_6232);
nor U8988 (N_8988,N_7050,N_6162);
nand U8989 (N_8989,N_7421,N_6303);
and U8990 (N_8990,N_7483,N_6423);
nor U8991 (N_8991,N_6331,N_7201);
and U8992 (N_8992,N_6154,N_7063);
or U8993 (N_8993,N_6221,N_7113);
or U8994 (N_8994,N_6932,N_7103);
nor U8995 (N_8995,N_6472,N_6311);
nor U8996 (N_8996,N_6265,N_6392);
and U8997 (N_8997,N_6236,N_6248);
xor U8998 (N_8998,N_6909,N_6320);
nand U8999 (N_8999,N_6709,N_6923);
nor U9000 (N_9000,N_8410,N_8106);
and U9001 (N_9001,N_8067,N_8637);
and U9002 (N_9002,N_7925,N_7694);
xnor U9003 (N_9003,N_8408,N_8248);
or U9004 (N_9004,N_7834,N_8472);
or U9005 (N_9005,N_7936,N_8386);
xnor U9006 (N_9006,N_8990,N_7707);
nor U9007 (N_9007,N_8891,N_8275);
nor U9008 (N_9008,N_7656,N_8355);
or U9009 (N_9009,N_8166,N_8543);
or U9010 (N_9010,N_8489,N_8692);
nor U9011 (N_9011,N_8033,N_8391);
nand U9012 (N_9012,N_7818,N_8219);
and U9013 (N_9013,N_8149,N_8256);
nor U9014 (N_9014,N_8153,N_8208);
and U9015 (N_9015,N_8384,N_8231);
and U9016 (N_9016,N_7685,N_8631);
xnor U9017 (N_9017,N_8460,N_8794);
and U9018 (N_9018,N_7551,N_8700);
and U9019 (N_9019,N_8999,N_7941);
or U9020 (N_9020,N_8047,N_8838);
nor U9021 (N_9021,N_8674,N_8158);
and U9022 (N_9022,N_7655,N_8381);
nand U9023 (N_9023,N_8235,N_7533);
or U9024 (N_9024,N_8485,N_8445);
xor U9025 (N_9025,N_8301,N_7939);
nand U9026 (N_9026,N_8128,N_7602);
or U9027 (N_9027,N_7733,N_8252);
and U9028 (N_9028,N_7703,N_8026);
xnor U9029 (N_9029,N_8500,N_7552);
and U9030 (N_9030,N_8726,N_8441);
nor U9031 (N_9031,N_8874,N_8012);
nor U9032 (N_9032,N_8182,N_7704);
or U9033 (N_9033,N_8684,N_8463);
or U9034 (N_9034,N_7529,N_8348);
and U9035 (N_9035,N_8091,N_8627);
or U9036 (N_9036,N_7579,N_8200);
or U9037 (N_9037,N_8747,N_7962);
nor U9038 (N_9038,N_8191,N_7929);
nor U9039 (N_9039,N_8496,N_8306);
nand U9040 (N_9040,N_8713,N_8734);
and U9041 (N_9041,N_8373,N_8326);
nor U9042 (N_9042,N_8881,N_8172);
or U9043 (N_9043,N_8201,N_7930);
nor U9044 (N_9044,N_7937,N_8746);
or U9045 (N_9045,N_8540,N_8056);
nand U9046 (N_9046,N_8458,N_7938);
and U9047 (N_9047,N_8982,N_8666);
and U9048 (N_9048,N_8216,N_8588);
nand U9049 (N_9049,N_7840,N_8819);
and U9050 (N_9050,N_8926,N_8553);
nor U9051 (N_9051,N_7799,N_8076);
nand U9052 (N_9052,N_7627,N_8327);
or U9053 (N_9053,N_8097,N_7565);
nor U9054 (N_9054,N_8488,N_8101);
or U9055 (N_9055,N_7928,N_8476);
or U9056 (N_9056,N_8749,N_8592);
nand U9057 (N_9057,N_8967,N_8593);
nor U9058 (N_9058,N_7861,N_8577);
or U9059 (N_9059,N_8133,N_7924);
nand U9060 (N_9060,N_8725,N_8646);
nand U9061 (N_9061,N_8896,N_8731);
nor U9062 (N_9062,N_7695,N_8486);
and U9063 (N_9063,N_8234,N_8919);
or U9064 (N_9064,N_8676,N_8045);
xor U9065 (N_9065,N_8126,N_8352);
and U9066 (N_9066,N_7511,N_8143);
and U9067 (N_9067,N_8261,N_8343);
nor U9068 (N_9068,N_8279,N_7893);
nor U9069 (N_9069,N_8758,N_7761);
nand U9070 (N_9070,N_7868,N_8171);
and U9071 (N_9071,N_7915,N_8576);
nand U9072 (N_9072,N_7754,N_8648);
and U9073 (N_9073,N_7796,N_8541);
or U9074 (N_9074,N_8781,N_8040);
nand U9075 (N_9075,N_8462,N_7859);
nand U9076 (N_9076,N_8548,N_7735);
nand U9077 (N_9077,N_8183,N_7981);
nand U9078 (N_9078,N_7586,N_8764);
nand U9079 (N_9079,N_8699,N_7527);
xor U9080 (N_9080,N_7611,N_7774);
or U9081 (N_9081,N_8428,N_8945);
xor U9082 (N_9082,N_8491,N_7633);
or U9083 (N_9083,N_7901,N_8229);
nor U9084 (N_9084,N_7839,N_7566);
nand U9085 (N_9085,N_7699,N_7767);
and U9086 (N_9086,N_8319,N_7688);
or U9087 (N_9087,N_8804,N_8230);
nor U9088 (N_9088,N_8148,N_8759);
xnor U9089 (N_9089,N_8020,N_8581);
nor U9090 (N_9090,N_7987,N_8887);
and U9091 (N_9091,N_8910,N_7709);
and U9092 (N_9092,N_7885,N_7526);
nor U9093 (N_9093,N_8903,N_8413);
or U9094 (N_9094,N_7944,N_7788);
xnor U9095 (N_9095,N_7714,N_8087);
xor U9096 (N_9096,N_8653,N_7741);
and U9097 (N_9097,N_8711,N_8382);
and U9098 (N_9098,N_8293,N_7605);
nor U9099 (N_9099,N_8089,N_7785);
nand U9100 (N_9100,N_8082,N_7524);
nand U9101 (N_9101,N_8647,N_8170);
and U9102 (N_9102,N_8003,N_7532);
nand U9103 (N_9103,N_8835,N_7597);
or U9104 (N_9104,N_8342,N_7876);
and U9105 (N_9105,N_7860,N_7554);
nor U9106 (N_9106,N_8797,N_7781);
nor U9107 (N_9107,N_8771,N_8251);
and U9108 (N_9108,N_7592,N_8288);
xor U9109 (N_9109,N_8103,N_7968);
xnor U9110 (N_9110,N_7793,N_7825);
nand U9111 (N_9111,N_8132,N_8241);
nand U9112 (N_9112,N_8972,N_8029);
nor U9113 (N_9113,N_8770,N_7813);
nor U9114 (N_9114,N_8691,N_7803);
and U9115 (N_9115,N_8439,N_8115);
nand U9116 (N_9116,N_8741,N_8004);
and U9117 (N_9117,N_8015,N_8430);
and U9118 (N_9118,N_7920,N_8389);
nand U9119 (N_9119,N_7686,N_7510);
nand U9120 (N_9120,N_8016,N_7652);
nor U9121 (N_9121,N_8437,N_8120);
nor U9122 (N_9122,N_8336,N_8791);
and U9123 (N_9123,N_7878,N_8858);
and U9124 (N_9124,N_7895,N_7724);
and U9125 (N_9125,N_7623,N_8471);
and U9126 (N_9126,N_8308,N_8583);
nor U9127 (N_9127,N_8071,N_8058);
nand U9128 (N_9128,N_8287,N_8524);
and U9129 (N_9129,N_8936,N_8333);
nand U9130 (N_9130,N_8187,N_7872);
and U9131 (N_9131,N_8265,N_8986);
and U9132 (N_9132,N_7864,N_8147);
and U9133 (N_9133,N_8065,N_8694);
nor U9134 (N_9134,N_7805,N_8636);
nor U9135 (N_9135,N_7519,N_7585);
xnor U9136 (N_9136,N_8899,N_7549);
and U9137 (N_9137,N_8715,N_7535);
and U9138 (N_9138,N_8947,N_7628);
and U9139 (N_9139,N_8597,N_8754);
or U9140 (N_9140,N_8924,N_8433);
nand U9141 (N_9141,N_8240,N_8236);
and U9142 (N_9142,N_8189,N_7687);
nand U9143 (N_9143,N_8314,N_8497);
and U9144 (N_9144,N_7959,N_8824);
and U9145 (N_9145,N_8761,N_8412);
and U9146 (N_9146,N_8285,N_8821);
or U9147 (N_9147,N_8523,N_7556);
and U9148 (N_9148,N_8867,N_7951);
or U9149 (N_9149,N_8803,N_8415);
nor U9150 (N_9150,N_8787,N_7521);
nand U9151 (N_9151,N_7618,N_8173);
or U9152 (N_9152,N_7934,N_8845);
nand U9153 (N_9153,N_8397,N_8121);
xor U9154 (N_9154,N_8568,N_8928);
nand U9155 (N_9155,N_7518,N_8532);
xnor U9156 (N_9156,N_8547,N_8102);
nor U9157 (N_9157,N_7772,N_7643);
or U9158 (N_9158,N_8923,N_7997);
nor U9159 (N_9159,N_7783,N_8518);
or U9160 (N_9160,N_8813,N_7693);
and U9161 (N_9161,N_7789,N_8228);
nand U9162 (N_9162,N_8425,N_8066);
and U9163 (N_9163,N_8882,N_7850);
or U9164 (N_9164,N_8828,N_8331);
nor U9165 (N_9165,N_8639,N_8169);
nor U9166 (N_9166,N_8602,N_8565);
nand U9167 (N_9167,N_8657,N_7851);
and U9168 (N_9168,N_8502,N_8808);
nor U9169 (N_9169,N_8802,N_8013);
or U9170 (N_9170,N_7515,N_8450);
xnor U9171 (N_9171,N_8546,N_8575);
nor U9172 (N_9172,N_8728,N_7844);
xnor U9173 (N_9173,N_8633,N_8107);
nand U9174 (N_9174,N_7620,N_7911);
and U9175 (N_9175,N_8374,N_8805);
nand U9176 (N_9176,N_8468,N_7675);
and U9177 (N_9177,N_8626,N_8084);
nand U9178 (N_9178,N_7988,N_8669);
nor U9179 (N_9179,N_8151,N_8008);
nand U9180 (N_9180,N_7947,N_7570);
nor U9181 (N_9181,N_8253,N_7809);
or U9182 (N_9182,N_8861,N_8160);
nor U9183 (N_9183,N_8337,N_7976);
and U9184 (N_9184,N_8063,N_8806);
or U9185 (N_9185,N_8017,N_8205);
and U9186 (N_9186,N_8185,N_8522);
nor U9187 (N_9187,N_7562,N_8226);
nor U9188 (N_9188,N_8589,N_7677);
nand U9189 (N_9189,N_8359,N_8975);
and U9190 (N_9190,N_8510,N_7942);
or U9191 (N_9191,N_8300,N_8283);
or U9192 (N_9192,N_8753,N_8704);
or U9193 (N_9193,N_8979,N_7642);
or U9194 (N_9194,N_8705,N_8459);
nor U9195 (N_9195,N_8150,N_7952);
nand U9196 (N_9196,N_8053,N_8788);
xnor U9197 (N_9197,N_8048,N_7517);
nor U9198 (N_9198,N_8856,N_8188);
nand U9199 (N_9199,N_7973,N_8981);
nand U9200 (N_9200,N_7810,N_8949);
nor U9201 (N_9201,N_7587,N_8827);
and U9202 (N_9202,N_8709,N_8651);
nand U9203 (N_9203,N_8334,N_8843);
or U9204 (N_9204,N_8390,N_7525);
and U9205 (N_9205,N_8745,N_8141);
or U9206 (N_9206,N_7739,N_7923);
and U9207 (N_9207,N_7949,N_8362);
nand U9208 (N_9208,N_8364,N_8707);
or U9209 (N_9209,N_8034,N_8095);
or U9210 (N_9210,N_8378,N_8712);
nand U9211 (N_9211,N_8629,N_7553);
nor U9212 (N_9212,N_7720,N_8880);
nor U9213 (N_9213,N_8181,N_8831);
nor U9214 (N_9214,N_8552,N_7683);
and U9215 (N_9215,N_7994,N_7974);
nand U9216 (N_9216,N_8365,N_8206);
and U9217 (N_9217,N_8885,N_8001);
xnor U9218 (N_9218,N_8587,N_8558);
xnor U9219 (N_9219,N_8325,N_8706);
nand U9220 (N_9220,N_8022,N_8640);
xnor U9221 (N_9221,N_8904,N_8339);
or U9222 (N_9222,N_8075,N_7730);
nor U9223 (N_9223,N_8179,N_8869);
xor U9224 (N_9224,N_7865,N_7603);
and U9225 (N_9225,N_8601,N_8162);
nand U9226 (N_9226,N_8035,N_8872);
and U9227 (N_9227,N_7582,N_7610);
nor U9228 (N_9228,N_8784,N_7630);
or U9229 (N_9229,N_8567,N_7978);
and U9230 (N_9230,N_7742,N_7622);
nand U9231 (N_9231,N_7800,N_8438);
and U9232 (N_9232,N_8934,N_7877);
nand U9233 (N_9233,N_8796,N_8623);
xnor U9234 (N_9234,N_7564,N_7691);
or U9235 (N_9235,N_7722,N_7500);
and U9236 (N_9236,N_8387,N_8105);
nor U9237 (N_9237,N_8564,N_8744);
or U9238 (N_9238,N_8608,N_8743);
nand U9239 (N_9239,N_7975,N_8135);
nand U9240 (N_9240,N_7747,N_8578);
nor U9241 (N_9241,N_8911,N_8670);
nor U9242 (N_9242,N_7966,N_8139);
nand U9243 (N_9243,N_8638,N_8790);
nand U9244 (N_9244,N_8984,N_7650);
or U9245 (N_9245,N_8370,N_8544);
nand U9246 (N_9246,N_8596,N_8224);
nand U9247 (N_9247,N_8534,N_8730);
nand U9248 (N_9248,N_8144,N_7982);
nor U9249 (N_9249,N_8156,N_7894);
or U9250 (N_9250,N_7670,N_7571);
nor U9251 (N_9251,N_8958,N_8406);
and U9252 (N_9252,N_8930,N_8559);
or U9253 (N_9253,N_8393,N_8511);
and U9254 (N_9254,N_8878,N_8571);
nor U9255 (N_9255,N_8944,N_7639);
xnor U9256 (N_9256,N_8921,N_8695);
and U9257 (N_9257,N_8442,N_8624);
and U9258 (N_9258,N_8424,N_8816);
or U9259 (N_9259,N_7880,N_8255);
and U9260 (N_9260,N_7824,N_8655);
nor U9261 (N_9261,N_7738,N_7624);
nor U9262 (N_9262,N_8165,N_8570);
nand U9263 (N_9263,N_8850,N_7869);
xnor U9264 (N_9264,N_8516,N_7673);
nand U9265 (N_9265,N_7651,N_7829);
or U9266 (N_9266,N_8582,N_8603);
nand U9267 (N_9267,N_8551,N_8893);
nor U9268 (N_9268,N_8330,N_8697);
nand U9269 (N_9269,N_8723,N_7736);
and U9270 (N_9270,N_8338,N_8680);
and U9271 (N_9271,N_7692,N_8863);
and U9272 (N_9272,N_8215,N_8690);
nor U9273 (N_9273,N_8154,N_7879);
and U9274 (N_9274,N_8988,N_7757);
nand U9275 (N_9275,N_7819,N_8873);
nand U9276 (N_9276,N_8773,N_8487);
or U9277 (N_9277,N_8533,N_7862);
and U9278 (N_9278,N_7581,N_8937);
nor U9279 (N_9279,N_7794,N_7608);
nor U9280 (N_9280,N_8772,N_8092);
and U9281 (N_9281,N_7625,N_8940);
and U9282 (N_9282,N_8913,N_8898);
nor U9283 (N_9283,N_8482,N_8607);
nand U9284 (N_9284,N_8599,N_7890);
nand U9285 (N_9285,N_8826,N_8072);
or U9286 (N_9286,N_8006,N_7575);
xnor U9287 (N_9287,N_8585,N_8473);
xnor U9288 (N_9288,N_8069,N_8563);
or U9289 (N_9289,N_7826,N_8118);
and U9290 (N_9290,N_8780,N_8536);
xnor U9291 (N_9291,N_8902,N_7909);
nor U9292 (N_9292,N_8799,N_8227);
and U9293 (N_9293,N_7873,N_8852);
or U9294 (N_9294,N_8019,N_8595);
or U9295 (N_9295,N_7857,N_7782);
nor U9296 (N_9296,N_7726,N_8825);
nor U9297 (N_9297,N_8014,N_8615);
nor U9298 (N_9298,N_8420,N_7737);
and U9299 (N_9299,N_8517,N_8290);
or U9300 (N_9300,N_7927,N_8380);
or U9301 (N_9301,N_7647,N_8096);
nand U9302 (N_9302,N_7886,N_7584);
or U9303 (N_9303,N_8262,N_8545);
nor U9304 (N_9304,N_7537,N_7616);
xor U9305 (N_9305,N_8399,N_7559);
nand U9306 (N_9306,N_8854,N_8762);
nor U9307 (N_9307,N_7921,N_7821);
xnor U9308 (N_9308,N_7768,N_8405);
and U9309 (N_9309,N_7672,N_8064);
nor U9310 (N_9310,N_7971,N_8480);
or U9311 (N_9311,N_7943,N_8807);
and U9312 (N_9312,N_8748,N_7995);
nand U9313 (N_9313,N_7904,N_7980);
and U9314 (N_9314,N_8630,N_8613);
and U9315 (N_9315,N_7658,N_7907);
nor U9316 (N_9316,N_8515,N_8011);
or U9317 (N_9317,N_8783,N_8436);
xor U9318 (N_9318,N_8675,N_8619);
nand U9319 (N_9319,N_8137,N_8466);
and U9320 (N_9320,N_8009,N_8829);
nor U9321 (N_9321,N_7956,N_8451);
and U9322 (N_9322,N_8628,N_7832);
nand U9323 (N_9323,N_8973,N_8789);
nand U9324 (N_9324,N_8233,N_7931);
or U9325 (N_9325,N_8481,N_7506);
nor U9326 (N_9326,N_7591,N_7577);
nand U9327 (N_9327,N_7888,N_7769);
nor U9328 (N_9328,N_8916,N_8579);
or U9329 (N_9329,N_7569,N_8038);
nand U9330 (N_9330,N_8719,N_8611);
or U9331 (N_9331,N_8952,N_8682);
nand U9332 (N_9332,N_8080,N_8266);
nor U9333 (N_9333,N_7791,N_8217);
nor U9334 (N_9334,N_7644,N_7899);
nand U9335 (N_9335,N_7682,N_8186);
xor U9336 (N_9336,N_8573,N_8278);
nor U9337 (N_9337,N_7706,N_8204);
and U9338 (N_9338,N_8010,N_7626);
or U9339 (N_9339,N_8260,N_7653);
nand U9340 (N_9340,N_7634,N_7640);
xnor U9341 (N_9341,N_8740,N_8814);
nor U9342 (N_9342,N_7866,N_8422);
nor U9343 (N_9343,N_8586,N_7985);
nor U9344 (N_9344,N_8722,N_8388);
nor U9345 (N_9345,N_8088,N_7705);
nor U9346 (N_9346,N_8376,N_8310);
nor U9347 (N_9347,N_7775,N_8469);
nor U9348 (N_9348,N_8119,N_8131);
xnor U9349 (N_9349,N_8635,N_8043);
nand U9350 (N_9350,N_8621,N_8164);
nand U9351 (N_9351,N_8935,N_7891);
or U9352 (N_9352,N_7563,N_8906);
and U9353 (N_9353,N_8693,N_8363);
and U9354 (N_9354,N_8556,N_8786);
and U9355 (N_9355,N_7836,N_8823);
nor U9356 (N_9356,N_8777,N_8672);
nand U9357 (N_9357,N_8023,N_8429);
or U9358 (N_9358,N_8978,N_7522);
and U9359 (N_9359,N_8353,N_7977);
or U9360 (N_9360,N_8566,N_7967);
and U9361 (N_9361,N_8963,N_7950);
or U9362 (N_9362,N_8032,N_7910);
nor U9363 (N_9363,N_8848,N_7897);
nand U9364 (N_9364,N_8316,N_8375);
or U9365 (N_9365,N_7842,N_8645);
or U9366 (N_9366,N_8477,N_8605);
nand U9367 (N_9367,N_8720,N_7933);
xnor U9368 (N_9368,N_8098,N_8474);
and U9369 (N_9369,N_7654,N_8404);
xor U9370 (N_9370,N_7752,N_8432);
nand U9371 (N_9371,N_7711,N_7725);
or U9372 (N_9372,N_8968,N_8938);
nor U9373 (N_9373,N_7712,N_8453);
or U9374 (N_9374,N_8851,N_8073);
nor U9375 (N_9375,N_8769,N_7847);
xor U9376 (N_9376,N_8870,N_8604);
nand U9377 (N_9377,N_8245,N_8509);
nand U9378 (N_9378,N_7595,N_8562);
and U9379 (N_9379,N_8057,N_8259);
xor U9380 (N_9380,N_8110,N_7776);
nor U9381 (N_9381,N_7749,N_7721);
xor U9382 (N_9382,N_8915,N_8136);
or U9383 (N_9383,N_8493,N_7993);
or U9384 (N_9384,N_8941,N_8443);
nor U9385 (N_9385,N_7790,N_8320);
nor U9386 (N_9386,N_8195,N_7723);
xor U9387 (N_9387,N_8535,N_7960);
nand U9388 (N_9388,N_7513,N_7753);
nor U9389 (N_9389,N_8421,N_7986);
nand U9390 (N_9390,N_7935,N_8724);
nand U9391 (N_9391,N_8737,N_7567);
and U9392 (N_9392,N_8736,N_7708);
xor U9393 (N_9393,N_8554,N_8254);
nand U9394 (N_9394,N_7674,N_8876);
nand U9395 (N_9395,N_7786,N_7883);
nand U9396 (N_9396,N_7727,N_7913);
nand U9397 (N_9397,N_8667,N_8396);
and U9398 (N_9398,N_8247,N_7520);
nand U9399 (N_9399,N_8037,N_7679);
or U9400 (N_9400,N_8907,N_8484);
nand U9401 (N_9401,N_8305,N_8964);
nand U9402 (N_9402,N_8176,N_8347);
and U9403 (N_9403,N_8322,N_8357);
nand U9404 (N_9404,N_8529,N_7574);
or U9405 (N_9405,N_8041,N_7867);
nor U9406 (N_9406,N_8093,N_8857);
and U9407 (N_9407,N_8917,N_7681);
or U9408 (N_9408,N_8218,N_8785);
nor U9409 (N_9409,N_8108,N_8202);
xnor U9410 (N_9410,N_7702,N_8811);
or U9411 (N_9411,N_8385,N_7743);
and U9412 (N_9412,N_8822,N_8526);
xnor U9413 (N_9413,N_8159,N_7534);
or U9414 (N_9414,N_7680,N_8892);
nor U9415 (N_9415,N_7875,N_8992);
or U9416 (N_9416,N_8994,N_8312);
nor U9417 (N_9417,N_8129,N_8503);
and U9418 (N_9418,N_8817,N_7755);
nand U9419 (N_9419,N_8263,N_7612);
or U9420 (N_9420,N_8905,N_8212);
and U9421 (N_9421,N_8324,N_7760);
xnor U9422 (N_9422,N_8409,N_8197);
nand U9423 (N_9423,N_8448,N_8211);
nand U9424 (N_9424,N_8427,N_8847);
nand U9425 (N_9425,N_7838,N_7599);
and U9426 (N_9426,N_8888,N_8561);
or U9427 (N_9427,N_7871,N_8049);
and U9428 (N_9428,N_8900,N_7700);
nor U9429 (N_9429,N_7889,N_7667);
nand U9430 (N_9430,N_8721,N_8100);
or U9431 (N_9431,N_7874,N_8302);
nor U9432 (N_9432,N_7505,N_8400);
nor U9433 (N_9433,N_8329,N_8061);
nand U9434 (N_9434,N_8617,N_8000);
nor U9435 (N_9435,N_7848,N_8414);
or U9436 (N_9436,N_7771,N_7698);
xnor U9437 (N_9437,N_8508,N_8871);
or U9438 (N_9438,N_7719,N_8598);
nand U9439 (N_9439,N_7713,N_8304);
nor U9440 (N_9440,N_7996,N_8750);
xnor U9441 (N_9441,N_8190,N_8083);
xor U9442 (N_9442,N_8113,N_7716);
and U9443 (N_9443,N_8527,N_7822);
nor U9444 (N_9444,N_8099,N_8834);
and U9445 (N_9445,N_8452,N_8678);
or U9446 (N_9446,N_7765,N_8738);
and U9447 (N_9447,N_7762,N_8710);
and U9448 (N_9448,N_7573,N_8225);
and U9449 (N_9449,N_8161,N_8766);
nand U9450 (N_9450,N_8125,N_8757);
nor U9451 (N_9451,N_8078,N_8213);
nand U9452 (N_9452,N_7807,N_7831);
nor U9453 (N_9453,N_7906,N_8142);
nor U9454 (N_9454,N_7665,N_8618);
or U9455 (N_9455,N_8818,N_7945);
and U9456 (N_9456,N_7501,N_8920);
nand U9457 (N_9457,N_7792,N_8660);
nand U9458 (N_9458,N_8795,N_8701);
and U9459 (N_9459,N_8687,N_8402);
or U9460 (N_9460,N_7657,N_7827);
and U9461 (N_9461,N_8447,N_8280);
nor U9462 (N_9462,N_8323,N_7764);
nor U9463 (N_9463,N_8270,N_8643);
xor U9464 (N_9464,N_8395,N_8950);
or U9465 (N_9465,N_8501,N_7528);
xor U9466 (N_9466,N_7841,N_7999);
nand U9467 (N_9467,N_8192,N_7815);
xnor U9468 (N_9468,N_8932,N_7902);
nand U9469 (N_9469,N_8074,N_8238);
and U9470 (N_9470,N_7898,N_8686);
and U9471 (N_9471,N_7835,N_7863);
or U9472 (N_9472,N_8054,N_7811);
nor U9473 (N_9473,N_7852,N_8239);
or U9474 (N_9474,N_7645,N_7663);
or U9475 (N_9475,N_7560,N_7732);
and U9476 (N_9476,N_7979,N_7837);
nor U9477 (N_9477,N_7887,N_7849);
or U9478 (N_9478,N_8664,N_8506);
and U9479 (N_9479,N_8908,N_8514);
nor U9480 (N_9480,N_8318,N_8993);
or U9481 (N_9481,N_7882,N_7545);
nor U9482 (N_9482,N_8220,N_7598);
or U9483 (N_9483,N_7823,N_8090);
nand U9484 (N_9484,N_7555,N_7636);
nor U9485 (N_9485,N_8394,N_7690);
and U9486 (N_9486,N_8594,N_8531);
nand U9487 (N_9487,N_8830,N_8328);
or U9488 (N_9488,N_7621,N_8127);
or U9489 (N_9489,N_8232,N_8112);
xnor U9490 (N_9490,N_8860,N_8776);
and U9491 (N_9491,N_8809,N_8475);
nand U9492 (N_9492,N_8525,N_8221);
or U9493 (N_9493,N_8959,N_8361);
nand U9494 (N_9494,N_7940,N_8068);
and U9495 (N_9495,N_8309,N_8953);
and U9496 (N_9496,N_8842,N_8449);
nor U9497 (N_9497,N_8292,N_7814);
nand U9498 (N_9498,N_8349,N_7607);
or U9499 (N_9499,N_8606,N_8864);
and U9500 (N_9500,N_8733,N_7972);
xnor U9501 (N_9501,N_8966,N_7661);
nand U9502 (N_9502,N_7905,N_8401);
or U9503 (N_9503,N_8340,N_7870);
or U9504 (N_9504,N_8435,N_8895);
and U9505 (N_9505,N_8955,N_8271);
nor U9506 (N_9506,N_7932,N_7744);
nand U9507 (N_9507,N_8574,N_8977);
xor U9508 (N_9508,N_8550,N_7740);
nor U9509 (N_9509,N_8492,N_8398);
nand U9510 (N_9510,N_7641,N_8942);
and U9511 (N_9511,N_8194,N_7779);
nor U9512 (N_9512,N_8498,N_8649);
and U9513 (N_9513,N_7502,N_8350);
or U9514 (N_9514,N_7746,N_8138);
nor U9515 (N_9515,N_8483,N_7715);
or U9516 (N_9516,N_8590,N_7992);
nor U9517 (N_9517,N_8600,N_7853);
and U9518 (N_9518,N_7766,N_8273);
nor U9519 (N_9519,N_8859,N_8294);
and U9520 (N_9520,N_7717,N_8461);
or U9521 (N_9521,N_8507,N_8767);
or U9522 (N_9522,N_8059,N_8122);
nor U9523 (N_9523,N_8094,N_8157);
or U9524 (N_9524,N_7922,N_7648);
xnor U9525 (N_9525,N_7504,N_8021);
and U9526 (N_9526,N_8372,N_8086);
nor U9527 (N_9527,N_8951,N_7900);
or U9528 (N_9528,N_8849,N_8569);
and U9529 (N_9529,N_8203,N_8104);
xnor U9530 (N_9530,N_8210,N_7614);
or U9531 (N_9531,N_8267,N_8250);
nor U9532 (N_9532,N_8855,N_7916);
nand U9533 (N_9533,N_8321,N_8846);
or U9534 (N_9534,N_8584,N_8987);
nand U9535 (N_9535,N_8454,N_7548);
nor U9536 (N_9536,N_8954,N_8335);
and U9537 (N_9537,N_8444,N_8960);
nand U9538 (N_9538,N_7512,N_8840);
nor U9539 (N_9539,N_7632,N_7990);
and U9540 (N_9540,N_8081,N_8971);
and U9541 (N_9541,N_8717,N_8123);
nor U9542 (N_9542,N_7550,N_7926);
and U9543 (N_9543,N_8311,N_8175);
and U9544 (N_9544,N_7546,N_7806);
nor U9545 (N_9545,N_8264,N_7701);
nand U9546 (N_9546,N_7745,N_7804);
or U9547 (N_9547,N_8495,N_8996);
or U9548 (N_9548,N_7590,N_8222);
and U9549 (N_9549,N_8542,N_8756);
and U9550 (N_9550,N_8989,N_7958);
or U9551 (N_9551,N_8890,N_8555);
and U9552 (N_9552,N_8889,N_8193);
and U9553 (N_9553,N_8163,N_7763);
or U9554 (N_9554,N_8379,N_8196);
nor U9555 (N_9555,N_8499,N_8572);
or U9556 (N_9556,N_8752,N_8877);
nand U9557 (N_9557,N_8146,N_8052);
nor U9558 (N_9558,N_7953,N_8024);
and U9559 (N_9559,N_7812,N_7778);
or U9560 (N_9560,N_8354,N_7820);
nand U9561 (N_9561,N_8403,N_8612);
nor U9562 (N_9562,N_7808,N_8681);
and U9563 (N_9563,N_8276,N_7543);
nor U9564 (N_9564,N_8299,N_8411);
or U9565 (N_9565,N_8465,N_8114);
nor U9566 (N_9566,N_8303,N_8027);
and U9567 (N_9567,N_8152,N_7756);
and U9568 (N_9568,N_7547,N_8774);
nor U9569 (N_9569,N_7750,N_8416);
and U9570 (N_9570,N_7955,N_8866);
nand U9571 (N_9571,N_7649,N_7539);
or U9572 (N_9572,N_7678,N_8243);
nor U9573 (N_9573,N_7731,N_7646);
and U9574 (N_9574,N_8839,N_8519);
and U9575 (N_9575,N_8685,N_8298);
and U9576 (N_9576,N_8018,N_8168);
nand U9577 (N_9577,N_8418,N_8641);
and U9578 (N_9578,N_8281,N_7538);
and U9579 (N_9579,N_7671,N_7594);
nand U9580 (N_9580,N_8044,N_7748);
nor U9581 (N_9581,N_7881,N_8530);
nor U9582 (N_9582,N_8258,N_8644);
and U9583 (N_9583,N_7588,N_8696);
nand U9584 (N_9584,N_8661,N_8961);
xnor U9585 (N_9585,N_8755,N_8371);
and U9586 (N_9586,N_8549,N_8307);
or U9587 (N_9587,N_7583,N_8313);
nor U9588 (N_9588,N_8367,N_8933);
or U9589 (N_9589,N_8894,N_8622);
and U9590 (N_9590,N_8274,N_7964);
and U9591 (N_9591,N_8957,N_8853);
nand U9592 (N_9592,N_8199,N_7855);
or U9593 (N_9593,N_8286,N_8237);
nand U9594 (N_9594,N_8031,N_7845);
xnor U9595 (N_9595,N_8560,N_8948);
or U9596 (N_9596,N_8922,N_8538);
nor U9597 (N_9597,N_8868,N_8223);
and U9598 (N_9598,N_8257,N_8284);
nand U9599 (N_9599,N_8007,N_8242);
nand U9600 (N_9600,N_8030,N_7846);
xor U9601 (N_9601,N_8528,N_8844);
and U9602 (N_9602,N_8134,N_8616);
xnor U9603 (N_9603,N_8956,N_7858);
or U9604 (N_9604,N_8778,N_7773);
nand U9605 (N_9605,N_7798,N_8070);
nor U9606 (N_9606,N_8668,N_8426);
nor U9607 (N_9607,N_8614,N_8505);
nand U9608 (N_9608,N_8297,N_8025);
nor U9609 (N_9609,N_8085,N_7659);
xor U9610 (N_9610,N_7593,N_7637);
or U9611 (N_9611,N_8046,N_8407);
and U9612 (N_9612,N_8209,N_8291);
and U9613 (N_9613,N_8446,N_7801);
nand U9614 (N_9614,N_8650,N_8727);
nor U9615 (N_9615,N_8673,N_8351);
nor U9616 (N_9616,N_7884,N_7843);
or U9617 (N_9617,N_7896,N_8289);
or U9618 (N_9618,N_8155,N_8671);
and U9619 (N_9619,N_8077,N_8998);
and U9620 (N_9620,N_7770,N_7965);
or U9621 (N_9621,N_8580,N_7918);
nand U9622 (N_9622,N_7600,N_8479);
nor U9623 (N_9623,N_8419,N_7669);
and U9624 (N_9624,N_8116,N_7542);
nand U9625 (N_9625,N_7666,N_8177);
nor U9626 (N_9626,N_8768,N_8591);
nor U9627 (N_9627,N_7596,N_7514);
nand U9628 (N_9628,N_8782,N_8974);
nor U9629 (N_9629,N_7984,N_7631);
or U9630 (N_9630,N_8702,N_7544);
xor U9631 (N_9631,N_7751,N_8079);
and U9632 (N_9632,N_8272,N_8642);
nor U9633 (N_9633,N_7629,N_7963);
or U9634 (N_9634,N_7780,N_8356);
nand U9635 (N_9635,N_8698,N_8927);
nand U9636 (N_9636,N_8042,N_8662);
nor U9637 (N_9637,N_8760,N_7833);
nand U9638 (N_9638,N_7589,N_7817);
nand U9639 (N_9639,N_7948,N_8841);
nand U9640 (N_9640,N_8111,N_8884);
xnor U9641 (N_9641,N_7734,N_8659);
xnor U9642 (N_9642,N_7830,N_7684);
or U9643 (N_9643,N_8912,N_8812);
xnor U9644 (N_9644,N_8997,N_7970);
and U9645 (N_9645,N_8965,N_8679);
nand U9646 (N_9646,N_8801,N_7892);
nand U9647 (N_9647,N_8918,N_8180);
nor U9648 (N_9648,N_8832,N_8837);
and U9649 (N_9649,N_8943,N_8358);
nor U9650 (N_9650,N_7619,N_8714);
nor U9651 (N_9651,N_8929,N_8360);
or U9652 (N_9652,N_7509,N_7568);
nor U9653 (N_9653,N_7728,N_8490);
xor U9654 (N_9654,N_8464,N_8383);
nor U9655 (N_9655,N_8494,N_7635);
and U9656 (N_9656,N_8632,N_8268);
nand U9657 (N_9657,N_8703,N_8800);
or U9658 (N_9658,N_7961,N_7664);
xor U9659 (N_9659,N_8991,N_7604);
or U9660 (N_9660,N_8366,N_7710);
or U9661 (N_9661,N_8976,N_8886);
nor U9662 (N_9662,N_8062,N_8879);
nand U9663 (N_9663,N_8742,N_7578);
xnor U9664 (N_9664,N_8368,N_8875);
nand U9665 (N_9665,N_8815,N_7854);
nor U9666 (N_9666,N_8798,N_7523);
xnor U9667 (N_9667,N_8665,N_8392);
nand U9668 (N_9668,N_8793,N_7998);
nor U9669 (N_9669,N_7609,N_8520);
and U9670 (N_9670,N_8688,N_8269);
nand U9671 (N_9671,N_8434,N_8763);
and U9672 (N_9672,N_7729,N_7516);
nand U9673 (N_9673,N_8055,N_8652);
nand U9674 (N_9674,N_8663,N_8537);
nand U9675 (N_9675,N_8862,N_7601);
or U9676 (N_9676,N_8145,N_8295);
or U9677 (N_9677,N_8332,N_7662);
nand U9678 (N_9678,N_8246,N_8440);
xnor U9679 (N_9679,N_8346,N_8513);
nand U9680 (N_9680,N_8689,N_7689);
nand U9681 (N_9681,N_7969,N_7557);
or U9682 (N_9682,N_8620,N_8625);
and U9683 (N_9683,N_7507,N_7787);
or U9684 (N_9684,N_8369,N_7957);
and U9685 (N_9685,N_8775,N_7503);
nor U9686 (N_9686,N_8198,N_8249);
or U9687 (N_9687,N_8931,N_8683);
and U9688 (N_9688,N_8039,N_8431);
and U9689 (N_9689,N_8377,N_8467);
and U9690 (N_9690,N_7606,N_7983);
nand U9691 (N_9691,N_7914,N_7917);
or U9692 (N_9692,N_8512,N_8124);
and U9693 (N_9693,N_8282,N_7795);
nand U9694 (N_9694,N_7676,N_8716);
nand U9695 (N_9695,N_8658,N_7777);
or U9696 (N_9696,N_8417,N_7660);
or U9697 (N_9697,N_8244,N_7617);
and U9698 (N_9698,N_7668,N_8317);
nor U9699 (N_9699,N_8732,N_8735);
and U9700 (N_9700,N_8901,N_8909);
nor U9701 (N_9701,N_8656,N_8117);
nand U9702 (N_9702,N_8939,N_7508);
or U9703 (N_9703,N_8820,N_8609);
nor U9704 (N_9704,N_7536,N_8140);
or U9705 (N_9705,N_8833,N_8296);
or U9706 (N_9706,N_7828,N_8610);
and U9707 (N_9707,N_8946,N_8174);
or U9708 (N_9708,N_8130,N_7530);
nor U9709 (N_9709,N_7784,N_8792);
and U9710 (N_9710,N_8729,N_8883);
and U9711 (N_9711,N_8478,N_8810);
or U9712 (N_9712,N_8983,N_7580);
nand U9713 (N_9713,N_7615,N_8865);
or U9714 (N_9714,N_8969,N_8005);
nor U9715 (N_9715,N_8751,N_8634);
nand U9716 (N_9716,N_8167,N_8028);
nand U9717 (N_9717,N_7919,N_7576);
and U9718 (N_9718,N_8962,N_7912);
or U9719 (N_9719,N_7558,N_7638);
nor U9720 (N_9720,N_8345,N_8708);
or U9721 (N_9721,N_8504,N_8765);
nand U9722 (N_9722,N_8455,N_8995);
nor U9723 (N_9723,N_8341,N_8677);
and U9724 (N_9724,N_7531,N_8980);
nor U9725 (N_9725,N_8207,N_7561);
nor U9726 (N_9726,N_8925,N_8718);
nor U9727 (N_9727,N_7903,N_8539);
nand U9728 (N_9728,N_8178,N_8985);
or U9729 (N_9729,N_8109,N_7697);
and U9730 (N_9730,N_7802,N_7797);
or U9731 (N_9731,N_7989,N_7718);
or U9732 (N_9732,N_8456,N_8470);
or U9733 (N_9733,N_8739,N_8002);
and U9734 (N_9734,N_8036,N_8423);
nor U9735 (N_9735,N_7991,N_8060);
and U9736 (N_9736,N_7954,N_7856);
and U9737 (N_9737,N_8836,N_7540);
and U9738 (N_9738,N_8457,N_8970);
or U9739 (N_9739,N_8557,N_8277);
nand U9740 (N_9740,N_7908,N_7758);
nor U9741 (N_9741,N_7572,N_8779);
nor U9742 (N_9742,N_7541,N_8050);
nand U9743 (N_9743,N_7696,N_8184);
nand U9744 (N_9744,N_7613,N_8654);
and U9745 (N_9745,N_7946,N_8521);
xnor U9746 (N_9746,N_7816,N_8914);
or U9747 (N_9747,N_7759,N_8051);
and U9748 (N_9748,N_8897,N_8315);
xor U9749 (N_9749,N_8344,N_8214);
xnor U9750 (N_9750,N_8385,N_7757);
or U9751 (N_9751,N_8461,N_7544);
and U9752 (N_9752,N_8556,N_8673);
nor U9753 (N_9753,N_8437,N_8908);
and U9754 (N_9754,N_8697,N_7858);
or U9755 (N_9755,N_7917,N_7752);
nor U9756 (N_9756,N_8228,N_8638);
xnor U9757 (N_9757,N_7917,N_7580);
or U9758 (N_9758,N_8395,N_7753);
nand U9759 (N_9759,N_8783,N_7556);
nand U9760 (N_9760,N_8506,N_8648);
and U9761 (N_9761,N_8866,N_8747);
nor U9762 (N_9762,N_7824,N_7831);
nor U9763 (N_9763,N_8893,N_8647);
and U9764 (N_9764,N_7594,N_7521);
nor U9765 (N_9765,N_7855,N_7845);
or U9766 (N_9766,N_8061,N_8229);
nand U9767 (N_9767,N_8254,N_7954);
and U9768 (N_9768,N_8743,N_8800);
nor U9769 (N_9769,N_8248,N_7857);
nand U9770 (N_9770,N_8355,N_8221);
nand U9771 (N_9771,N_7956,N_8773);
nand U9772 (N_9772,N_8119,N_7520);
or U9773 (N_9773,N_8841,N_7588);
and U9774 (N_9774,N_8789,N_7886);
and U9775 (N_9775,N_7538,N_8123);
nor U9776 (N_9776,N_7583,N_7911);
nand U9777 (N_9777,N_7737,N_8876);
or U9778 (N_9778,N_7976,N_8367);
and U9779 (N_9779,N_8122,N_8917);
nand U9780 (N_9780,N_7681,N_8733);
nand U9781 (N_9781,N_8253,N_8116);
and U9782 (N_9782,N_7515,N_8649);
nor U9783 (N_9783,N_7594,N_8760);
or U9784 (N_9784,N_7502,N_8863);
nor U9785 (N_9785,N_8758,N_8231);
nor U9786 (N_9786,N_8951,N_8875);
nor U9787 (N_9787,N_8117,N_8084);
and U9788 (N_9788,N_8697,N_8183);
nor U9789 (N_9789,N_8145,N_7754);
nand U9790 (N_9790,N_8854,N_8895);
nand U9791 (N_9791,N_7812,N_8319);
nor U9792 (N_9792,N_7635,N_8396);
nor U9793 (N_9793,N_8854,N_8267);
nand U9794 (N_9794,N_8797,N_8676);
nand U9795 (N_9795,N_8213,N_8115);
nand U9796 (N_9796,N_7830,N_8543);
or U9797 (N_9797,N_8521,N_8522);
or U9798 (N_9798,N_8926,N_8795);
xor U9799 (N_9799,N_8889,N_8693);
and U9800 (N_9800,N_8013,N_8486);
nand U9801 (N_9801,N_8508,N_8765);
xor U9802 (N_9802,N_8826,N_7761);
and U9803 (N_9803,N_7863,N_8757);
xor U9804 (N_9804,N_7509,N_8914);
or U9805 (N_9805,N_8971,N_8109);
nor U9806 (N_9806,N_7830,N_7767);
xor U9807 (N_9807,N_7947,N_7603);
and U9808 (N_9808,N_8228,N_7816);
nor U9809 (N_9809,N_7668,N_8031);
and U9810 (N_9810,N_8782,N_7986);
nor U9811 (N_9811,N_7992,N_8954);
xor U9812 (N_9812,N_8293,N_7595);
or U9813 (N_9813,N_8604,N_7731);
and U9814 (N_9814,N_8985,N_7650);
or U9815 (N_9815,N_7515,N_8978);
nand U9816 (N_9816,N_8158,N_8733);
or U9817 (N_9817,N_8381,N_7747);
nand U9818 (N_9818,N_8547,N_8082);
and U9819 (N_9819,N_8808,N_8782);
nand U9820 (N_9820,N_7925,N_8119);
or U9821 (N_9821,N_8170,N_8034);
and U9822 (N_9822,N_7504,N_8989);
nand U9823 (N_9823,N_8052,N_8749);
nand U9824 (N_9824,N_7791,N_7846);
xor U9825 (N_9825,N_8464,N_8647);
xor U9826 (N_9826,N_7851,N_7745);
and U9827 (N_9827,N_7786,N_8123);
nand U9828 (N_9828,N_8752,N_7987);
or U9829 (N_9829,N_8595,N_8507);
or U9830 (N_9830,N_8894,N_7979);
nand U9831 (N_9831,N_7580,N_8999);
xor U9832 (N_9832,N_8525,N_7981);
nor U9833 (N_9833,N_8997,N_7971);
or U9834 (N_9834,N_8444,N_7991);
or U9835 (N_9835,N_8076,N_8149);
nor U9836 (N_9836,N_8874,N_7660);
or U9837 (N_9837,N_8744,N_8023);
xor U9838 (N_9838,N_7748,N_8354);
nor U9839 (N_9839,N_8771,N_7628);
nand U9840 (N_9840,N_8513,N_8631);
and U9841 (N_9841,N_8366,N_8841);
nor U9842 (N_9842,N_7925,N_7634);
nor U9843 (N_9843,N_7636,N_8642);
or U9844 (N_9844,N_8772,N_8449);
or U9845 (N_9845,N_8626,N_8121);
or U9846 (N_9846,N_8383,N_8518);
and U9847 (N_9847,N_8232,N_8881);
and U9848 (N_9848,N_8309,N_8151);
and U9849 (N_9849,N_7757,N_8096);
or U9850 (N_9850,N_8960,N_7535);
nor U9851 (N_9851,N_7959,N_8662);
and U9852 (N_9852,N_8532,N_8747);
nor U9853 (N_9853,N_8500,N_8929);
nand U9854 (N_9854,N_8133,N_8926);
and U9855 (N_9855,N_8369,N_8201);
and U9856 (N_9856,N_8227,N_8977);
and U9857 (N_9857,N_8394,N_7500);
and U9858 (N_9858,N_7724,N_7997);
nand U9859 (N_9859,N_8228,N_7943);
and U9860 (N_9860,N_8995,N_7560);
or U9861 (N_9861,N_8123,N_7506);
or U9862 (N_9862,N_8013,N_8833);
or U9863 (N_9863,N_8474,N_8815);
nor U9864 (N_9864,N_8256,N_8088);
nand U9865 (N_9865,N_8507,N_7820);
nor U9866 (N_9866,N_8183,N_8347);
or U9867 (N_9867,N_8505,N_8201);
or U9868 (N_9868,N_8003,N_8665);
and U9869 (N_9869,N_7953,N_8278);
nor U9870 (N_9870,N_8019,N_7748);
nor U9871 (N_9871,N_8825,N_8888);
and U9872 (N_9872,N_7945,N_8634);
nor U9873 (N_9873,N_8526,N_7782);
nand U9874 (N_9874,N_7777,N_7767);
or U9875 (N_9875,N_8714,N_8649);
and U9876 (N_9876,N_7569,N_8941);
xnor U9877 (N_9877,N_8398,N_8264);
or U9878 (N_9878,N_8195,N_8896);
or U9879 (N_9879,N_8689,N_8821);
nor U9880 (N_9880,N_8838,N_8993);
nand U9881 (N_9881,N_7815,N_8222);
nand U9882 (N_9882,N_8950,N_7800);
nor U9883 (N_9883,N_7761,N_8171);
nor U9884 (N_9884,N_8746,N_8804);
or U9885 (N_9885,N_8499,N_8732);
or U9886 (N_9886,N_7830,N_8680);
xnor U9887 (N_9887,N_8139,N_8929);
and U9888 (N_9888,N_8288,N_8421);
nand U9889 (N_9889,N_7766,N_8272);
or U9890 (N_9890,N_8712,N_7694);
or U9891 (N_9891,N_8116,N_8746);
nand U9892 (N_9892,N_8619,N_8980);
xor U9893 (N_9893,N_8577,N_8093);
nor U9894 (N_9894,N_8854,N_8825);
and U9895 (N_9895,N_8337,N_7863);
nand U9896 (N_9896,N_7941,N_7944);
nor U9897 (N_9897,N_8862,N_8811);
and U9898 (N_9898,N_8910,N_8474);
or U9899 (N_9899,N_8933,N_7955);
nand U9900 (N_9900,N_7549,N_7577);
or U9901 (N_9901,N_7559,N_8640);
and U9902 (N_9902,N_8982,N_8051);
nor U9903 (N_9903,N_7758,N_7832);
nand U9904 (N_9904,N_8605,N_7914);
nor U9905 (N_9905,N_7585,N_8714);
or U9906 (N_9906,N_7863,N_8934);
nor U9907 (N_9907,N_7766,N_8821);
nand U9908 (N_9908,N_8188,N_8140);
and U9909 (N_9909,N_8846,N_7745);
and U9910 (N_9910,N_8841,N_8695);
nor U9911 (N_9911,N_8171,N_7917);
xnor U9912 (N_9912,N_8214,N_8924);
or U9913 (N_9913,N_8765,N_7588);
nor U9914 (N_9914,N_8945,N_8964);
and U9915 (N_9915,N_7885,N_7834);
or U9916 (N_9916,N_7576,N_8824);
and U9917 (N_9917,N_7704,N_8255);
and U9918 (N_9918,N_7699,N_8831);
nor U9919 (N_9919,N_8417,N_8956);
nand U9920 (N_9920,N_8256,N_7915);
and U9921 (N_9921,N_8867,N_8596);
and U9922 (N_9922,N_8184,N_8789);
nand U9923 (N_9923,N_8632,N_8570);
and U9924 (N_9924,N_8105,N_8407);
xnor U9925 (N_9925,N_8810,N_8463);
nor U9926 (N_9926,N_8799,N_8204);
and U9927 (N_9927,N_7919,N_7550);
or U9928 (N_9928,N_8686,N_8542);
nor U9929 (N_9929,N_7822,N_8340);
nor U9930 (N_9930,N_8613,N_7574);
nor U9931 (N_9931,N_7792,N_8324);
nand U9932 (N_9932,N_8332,N_8738);
or U9933 (N_9933,N_8898,N_8583);
nand U9934 (N_9934,N_8800,N_8122);
and U9935 (N_9935,N_8492,N_7825);
nor U9936 (N_9936,N_8389,N_7759);
and U9937 (N_9937,N_8516,N_7591);
nand U9938 (N_9938,N_8452,N_8418);
and U9939 (N_9939,N_8477,N_7742);
or U9940 (N_9940,N_7539,N_8206);
xor U9941 (N_9941,N_7511,N_8015);
or U9942 (N_9942,N_8993,N_7591);
and U9943 (N_9943,N_8083,N_7771);
and U9944 (N_9944,N_8211,N_7536);
nor U9945 (N_9945,N_8905,N_8324);
nand U9946 (N_9946,N_7921,N_8864);
nand U9947 (N_9947,N_8258,N_7898);
nor U9948 (N_9948,N_8381,N_8959);
nor U9949 (N_9949,N_7899,N_8838);
and U9950 (N_9950,N_8440,N_7859);
or U9951 (N_9951,N_8214,N_8879);
or U9952 (N_9952,N_7909,N_8689);
or U9953 (N_9953,N_8197,N_7911);
and U9954 (N_9954,N_7625,N_7956);
and U9955 (N_9955,N_7619,N_7829);
or U9956 (N_9956,N_7559,N_7980);
and U9957 (N_9957,N_8782,N_8859);
xnor U9958 (N_9958,N_8292,N_8860);
and U9959 (N_9959,N_7638,N_7829);
and U9960 (N_9960,N_8788,N_7629);
nand U9961 (N_9961,N_7682,N_8037);
nor U9962 (N_9962,N_7836,N_7684);
nor U9963 (N_9963,N_7526,N_7740);
or U9964 (N_9964,N_8132,N_8027);
nand U9965 (N_9965,N_7625,N_8184);
nand U9966 (N_9966,N_7817,N_8386);
and U9967 (N_9967,N_8835,N_8393);
nor U9968 (N_9968,N_7860,N_8148);
and U9969 (N_9969,N_8879,N_7789);
nand U9970 (N_9970,N_7556,N_8206);
nand U9971 (N_9971,N_8776,N_7944);
and U9972 (N_9972,N_8414,N_7616);
nor U9973 (N_9973,N_7773,N_7533);
xnor U9974 (N_9974,N_7508,N_8050);
or U9975 (N_9975,N_8511,N_8621);
nand U9976 (N_9976,N_8110,N_8236);
xor U9977 (N_9977,N_8376,N_8644);
or U9978 (N_9978,N_8212,N_8794);
and U9979 (N_9979,N_7617,N_8199);
and U9980 (N_9980,N_8682,N_8728);
nand U9981 (N_9981,N_8914,N_8988);
and U9982 (N_9982,N_8550,N_7647);
and U9983 (N_9983,N_8392,N_8428);
and U9984 (N_9984,N_8069,N_8589);
and U9985 (N_9985,N_8251,N_7663);
xnor U9986 (N_9986,N_8844,N_7729);
or U9987 (N_9987,N_8108,N_8153);
nor U9988 (N_9988,N_8194,N_7803);
xor U9989 (N_9989,N_7815,N_8660);
nand U9990 (N_9990,N_8758,N_7701);
or U9991 (N_9991,N_7922,N_8241);
or U9992 (N_9992,N_8491,N_7780);
nor U9993 (N_9993,N_8985,N_8104);
and U9994 (N_9994,N_8677,N_7807);
and U9995 (N_9995,N_8745,N_8539);
nor U9996 (N_9996,N_7574,N_7624);
and U9997 (N_9997,N_7597,N_8057);
or U9998 (N_9998,N_8356,N_8748);
nor U9999 (N_9999,N_8632,N_8492);
nand U10000 (N_10000,N_8175,N_7678);
nor U10001 (N_10001,N_8399,N_8916);
nand U10002 (N_10002,N_8183,N_8928);
xnor U10003 (N_10003,N_8901,N_8757);
or U10004 (N_10004,N_8426,N_7632);
nand U10005 (N_10005,N_7552,N_7521);
or U10006 (N_10006,N_7730,N_8619);
nand U10007 (N_10007,N_7686,N_7572);
xnor U10008 (N_10008,N_8325,N_8960);
nor U10009 (N_10009,N_8193,N_7953);
nand U10010 (N_10010,N_8034,N_8689);
nand U10011 (N_10011,N_7934,N_8882);
nand U10012 (N_10012,N_7885,N_7884);
nand U10013 (N_10013,N_8727,N_8519);
or U10014 (N_10014,N_8042,N_7690);
and U10015 (N_10015,N_8993,N_8889);
xor U10016 (N_10016,N_8158,N_7622);
xnor U10017 (N_10017,N_8051,N_8181);
nor U10018 (N_10018,N_8255,N_7536);
xor U10019 (N_10019,N_7977,N_7520);
nand U10020 (N_10020,N_8563,N_8797);
or U10021 (N_10021,N_8981,N_8351);
nor U10022 (N_10022,N_7881,N_7874);
and U10023 (N_10023,N_8181,N_8554);
nor U10024 (N_10024,N_8740,N_7625);
nor U10025 (N_10025,N_8549,N_8535);
and U10026 (N_10026,N_8667,N_8444);
or U10027 (N_10027,N_8035,N_7783);
nand U10028 (N_10028,N_8030,N_8529);
nor U10029 (N_10029,N_8544,N_8674);
nor U10030 (N_10030,N_8536,N_8917);
or U10031 (N_10031,N_8991,N_7659);
xor U10032 (N_10032,N_8812,N_8743);
nand U10033 (N_10033,N_7522,N_8376);
and U10034 (N_10034,N_7768,N_8883);
nor U10035 (N_10035,N_8927,N_7802);
nand U10036 (N_10036,N_8627,N_8950);
xor U10037 (N_10037,N_8609,N_7545);
nor U10038 (N_10038,N_8266,N_8865);
or U10039 (N_10039,N_7599,N_8584);
nand U10040 (N_10040,N_8106,N_8091);
nand U10041 (N_10041,N_7507,N_8412);
nor U10042 (N_10042,N_7524,N_7953);
or U10043 (N_10043,N_8687,N_8046);
or U10044 (N_10044,N_7995,N_7521);
or U10045 (N_10045,N_8779,N_8675);
or U10046 (N_10046,N_8711,N_7634);
nor U10047 (N_10047,N_7553,N_7585);
nand U10048 (N_10048,N_8161,N_8791);
or U10049 (N_10049,N_8830,N_7910);
nor U10050 (N_10050,N_7989,N_8422);
nand U10051 (N_10051,N_7877,N_7996);
nand U10052 (N_10052,N_8107,N_8367);
nor U10053 (N_10053,N_8713,N_7911);
and U10054 (N_10054,N_8664,N_8583);
or U10055 (N_10055,N_8456,N_8208);
nand U10056 (N_10056,N_8719,N_8498);
or U10057 (N_10057,N_8780,N_8971);
nor U10058 (N_10058,N_8293,N_7903);
or U10059 (N_10059,N_8773,N_8858);
nand U10060 (N_10060,N_8013,N_8638);
nor U10061 (N_10061,N_7696,N_8644);
and U10062 (N_10062,N_8075,N_8874);
nor U10063 (N_10063,N_8405,N_8000);
nor U10064 (N_10064,N_7898,N_8803);
and U10065 (N_10065,N_8090,N_8557);
nor U10066 (N_10066,N_8205,N_8523);
or U10067 (N_10067,N_8406,N_8377);
or U10068 (N_10068,N_8453,N_8065);
and U10069 (N_10069,N_7695,N_8894);
and U10070 (N_10070,N_8405,N_7635);
and U10071 (N_10071,N_8217,N_8180);
and U10072 (N_10072,N_8810,N_8298);
or U10073 (N_10073,N_8999,N_7967);
or U10074 (N_10074,N_8796,N_8741);
nor U10075 (N_10075,N_8826,N_7905);
and U10076 (N_10076,N_7834,N_8826);
nand U10077 (N_10077,N_8746,N_8066);
nor U10078 (N_10078,N_8421,N_8300);
or U10079 (N_10079,N_8019,N_8831);
nand U10080 (N_10080,N_8037,N_8457);
nor U10081 (N_10081,N_8004,N_7699);
nor U10082 (N_10082,N_7971,N_8271);
and U10083 (N_10083,N_8862,N_7818);
xnor U10084 (N_10084,N_8915,N_7562);
nor U10085 (N_10085,N_8179,N_8243);
nand U10086 (N_10086,N_7755,N_8117);
nor U10087 (N_10087,N_7910,N_8277);
nor U10088 (N_10088,N_8112,N_8179);
or U10089 (N_10089,N_8763,N_8820);
and U10090 (N_10090,N_8847,N_8156);
nor U10091 (N_10091,N_8697,N_8768);
and U10092 (N_10092,N_7581,N_8501);
and U10093 (N_10093,N_8691,N_8715);
and U10094 (N_10094,N_8130,N_7908);
nor U10095 (N_10095,N_8772,N_8016);
nor U10096 (N_10096,N_8383,N_7581);
xor U10097 (N_10097,N_8794,N_8145);
nor U10098 (N_10098,N_8677,N_8811);
nand U10099 (N_10099,N_8564,N_7912);
or U10100 (N_10100,N_8266,N_7518);
nand U10101 (N_10101,N_8487,N_8962);
and U10102 (N_10102,N_8662,N_7850);
and U10103 (N_10103,N_8110,N_7516);
or U10104 (N_10104,N_7800,N_7536);
or U10105 (N_10105,N_7930,N_7817);
nor U10106 (N_10106,N_7594,N_7731);
xor U10107 (N_10107,N_8494,N_8130);
or U10108 (N_10108,N_8364,N_8343);
or U10109 (N_10109,N_8115,N_8905);
nor U10110 (N_10110,N_7704,N_8194);
and U10111 (N_10111,N_7902,N_7724);
or U10112 (N_10112,N_8225,N_7687);
nor U10113 (N_10113,N_8168,N_8815);
nor U10114 (N_10114,N_8943,N_8638);
nor U10115 (N_10115,N_8395,N_8364);
or U10116 (N_10116,N_7819,N_8457);
and U10117 (N_10117,N_8029,N_7617);
nor U10118 (N_10118,N_8795,N_8276);
nor U10119 (N_10119,N_8095,N_8317);
or U10120 (N_10120,N_7665,N_8627);
nor U10121 (N_10121,N_7627,N_8353);
or U10122 (N_10122,N_7721,N_8781);
and U10123 (N_10123,N_8137,N_8759);
nand U10124 (N_10124,N_8337,N_7517);
nand U10125 (N_10125,N_7600,N_8262);
or U10126 (N_10126,N_8234,N_8453);
xnor U10127 (N_10127,N_8885,N_8700);
nor U10128 (N_10128,N_8788,N_8740);
xnor U10129 (N_10129,N_7590,N_8630);
or U10130 (N_10130,N_8377,N_8114);
and U10131 (N_10131,N_8437,N_8400);
xnor U10132 (N_10132,N_7966,N_8426);
or U10133 (N_10133,N_8117,N_7516);
and U10134 (N_10134,N_7670,N_8227);
nand U10135 (N_10135,N_8699,N_8739);
or U10136 (N_10136,N_8711,N_8385);
and U10137 (N_10137,N_8783,N_7979);
or U10138 (N_10138,N_8737,N_7849);
nor U10139 (N_10139,N_7758,N_8412);
and U10140 (N_10140,N_7736,N_8425);
nor U10141 (N_10141,N_8011,N_8593);
or U10142 (N_10142,N_7893,N_7564);
nor U10143 (N_10143,N_7815,N_7553);
nor U10144 (N_10144,N_8525,N_7708);
or U10145 (N_10145,N_8141,N_8094);
nand U10146 (N_10146,N_8690,N_8969);
nor U10147 (N_10147,N_7693,N_7991);
and U10148 (N_10148,N_8522,N_8383);
or U10149 (N_10149,N_8906,N_7923);
nor U10150 (N_10150,N_8126,N_8135);
nor U10151 (N_10151,N_7658,N_8777);
or U10152 (N_10152,N_8502,N_8050);
and U10153 (N_10153,N_8833,N_8770);
or U10154 (N_10154,N_8276,N_8806);
nor U10155 (N_10155,N_8397,N_7683);
and U10156 (N_10156,N_8252,N_7789);
or U10157 (N_10157,N_8986,N_8251);
nor U10158 (N_10158,N_7798,N_8583);
and U10159 (N_10159,N_8027,N_8139);
xor U10160 (N_10160,N_8065,N_8766);
nand U10161 (N_10161,N_8106,N_7912);
or U10162 (N_10162,N_8983,N_8976);
or U10163 (N_10163,N_8135,N_8623);
xor U10164 (N_10164,N_7783,N_8125);
nor U10165 (N_10165,N_8347,N_7879);
nor U10166 (N_10166,N_7626,N_8719);
nor U10167 (N_10167,N_8534,N_8342);
nand U10168 (N_10168,N_8914,N_8461);
or U10169 (N_10169,N_8567,N_8730);
xor U10170 (N_10170,N_7759,N_8597);
nor U10171 (N_10171,N_8910,N_7863);
and U10172 (N_10172,N_7780,N_8671);
or U10173 (N_10173,N_8632,N_8317);
nor U10174 (N_10174,N_7982,N_8496);
or U10175 (N_10175,N_8707,N_8827);
and U10176 (N_10176,N_8855,N_8571);
or U10177 (N_10177,N_8816,N_8761);
nand U10178 (N_10178,N_8538,N_7667);
or U10179 (N_10179,N_8603,N_7965);
or U10180 (N_10180,N_8564,N_8928);
and U10181 (N_10181,N_7547,N_7913);
and U10182 (N_10182,N_8173,N_7784);
xnor U10183 (N_10183,N_8615,N_7551);
xnor U10184 (N_10184,N_8660,N_8720);
and U10185 (N_10185,N_7594,N_8766);
and U10186 (N_10186,N_7736,N_7989);
xnor U10187 (N_10187,N_7661,N_7903);
and U10188 (N_10188,N_8071,N_8230);
or U10189 (N_10189,N_8043,N_8650);
and U10190 (N_10190,N_8869,N_7532);
and U10191 (N_10191,N_8233,N_7935);
nor U10192 (N_10192,N_8507,N_7756);
or U10193 (N_10193,N_8496,N_7931);
nand U10194 (N_10194,N_7823,N_8132);
and U10195 (N_10195,N_8854,N_8562);
nand U10196 (N_10196,N_8207,N_8216);
nor U10197 (N_10197,N_7875,N_8916);
nor U10198 (N_10198,N_7856,N_8968);
and U10199 (N_10199,N_8392,N_7979);
or U10200 (N_10200,N_8558,N_7932);
and U10201 (N_10201,N_8758,N_8803);
nand U10202 (N_10202,N_8235,N_8213);
and U10203 (N_10203,N_8451,N_7637);
and U10204 (N_10204,N_8146,N_8554);
or U10205 (N_10205,N_8329,N_8973);
nor U10206 (N_10206,N_8927,N_8925);
nor U10207 (N_10207,N_7879,N_8405);
or U10208 (N_10208,N_7644,N_8989);
nand U10209 (N_10209,N_8562,N_8903);
or U10210 (N_10210,N_7792,N_7761);
and U10211 (N_10211,N_8357,N_7550);
or U10212 (N_10212,N_8907,N_8562);
nand U10213 (N_10213,N_8289,N_7937);
and U10214 (N_10214,N_8014,N_8169);
nor U10215 (N_10215,N_7513,N_8680);
nor U10216 (N_10216,N_8548,N_8483);
nand U10217 (N_10217,N_8941,N_8818);
nand U10218 (N_10218,N_8160,N_8529);
xor U10219 (N_10219,N_8329,N_7871);
nor U10220 (N_10220,N_8343,N_7795);
or U10221 (N_10221,N_8680,N_8031);
nand U10222 (N_10222,N_8253,N_8784);
and U10223 (N_10223,N_7599,N_7987);
nor U10224 (N_10224,N_7540,N_8441);
nor U10225 (N_10225,N_7903,N_7836);
nor U10226 (N_10226,N_8768,N_8342);
xor U10227 (N_10227,N_7631,N_8133);
and U10228 (N_10228,N_8065,N_7577);
nand U10229 (N_10229,N_7583,N_8839);
or U10230 (N_10230,N_7929,N_8336);
or U10231 (N_10231,N_8032,N_8176);
nor U10232 (N_10232,N_7513,N_8049);
nor U10233 (N_10233,N_8919,N_8789);
nand U10234 (N_10234,N_8434,N_8149);
and U10235 (N_10235,N_8357,N_8502);
or U10236 (N_10236,N_8084,N_8935);
and U10237 (N_10237,N_8506,N_8931);
nor U10238 (N_10238,N_7817,N_8272);
and U10239 (N_10239,N_8701,N_8860);
or U10240 (N_10240,N_8159,N_7550);
and U10241 (N_10241,N_8934,N_8060);
nand U10242 (N_10242,N_8752,N_8179);
nand U10243 (N_10243,N_7717,N_7715);
nor U10244 (N_10244,N_7756,N_7588);
nor U10245 (N_10245,N_8357,N_7780);
nor U10246 (N_10246,N_7670,N_7533);
nand U10247 (N_10247,N_8153,N_7728);
or U10248 (N_10248,N_7882,N_8177);
nand U10249 (N_10249,N_8457,N_8461);
or U10250 (N_10250,N_8574,N_7876);
nor U10251 (N_10251,N_8414,N_7656);
nand U10252 (N_10252,N_8805,N_7864);
or U10253 (N_10253,N_7885,N_8672);
xnor U10254 (N_10254,N_7540,N_8485);
nor U10255 (N_10255,N_8159,N_8857);
or U10256 (N_10256,N_8709,N_7787);
xor U10257 (N_10257,N_8117,N_8397);
xnor U10258 (N_10258,N_8857,N_8701);
nand U10259 (N_10259,N_8077,N_7875);
and U10260 (N_10260,N_7549,N_8425);
or U10261 (N_10261,N_7639,N_7500);
nand U10262 (N_10262,N_8807,N_8499);
and U10263 (N_10263,N_8765,N_7652);
or U10264 (N_10264,N_7841,N_7804);
xor U10265 (N_10265,N_8857,N_8919);
nor U10266 (N_10266,N_7764,N_8485);
or U10267 (N_10267,N_8977,N_8216);
or U10268 (N_10268,N_7676,N_8892);
nor U10269 (N_10269,N_8588,N_8625);
xnor U10270 (N_10270,N_8464,N_7624);
or U10271 (N_10271,N_7956,N_8808);
nor U10272 (N_10272,N_8130,N_8510);
xor U10273 (N_10273,N_8877,N_8211);
and U10274 (N_10274,N_7722,N_8303);
nor U10275 (N_10275,N_7613,N_7624);
nand U10276 (N_10276,N_7768,N_7789);
or U10277 (N_10277,N_7630,N_7976);
nand U10278 (N_10278,N_8785,N_8723);
or U10279 (N_10279,N_7759,N_8626);
or U10280 (N_10280,N_7964,N_8714);
or U10281 (N_10281,N_8169,N_7980);
xnor U10282 (N_10282,N_8925,N_7875);
and U10283 (N_10283,N_8172,N_8715);
or U10284 (N_10284,N_7654,N_8849);
and U10285 (N_10285,N_8872,N_8256);
and U10286 (N_10286,N_8327,N_8071);
or U10287 (N_10287,N_7798,N_7648);
nand U10288 (N_10288,N_8052,N_7917);
xor U10289 (N_10289,N_7639,N_7840);
xor U10290 (N_10290,N_7617,N_8529);
xnor U10291 (N_10291,N_8683,N_8340);
xnor U10292 (N_10292,N_8722,N_8321);
or U10293 (N_10293,N_8107,N_7890);
or U10294 (N_10294,N_7819,N_7685);
and U10295 (N_10295,N_7743,N_7718);
and U10296 (N_10296,N_8410,N_7888);
nand U10297 (N_10297,N_8482,N_8379);
nand U10298 (N_10298,N_8283,N_8184);
nand U10299 (N_10299,N_7764,N_8835);
nor U10300 (N_10300,N_8105,N_7892);
or U10301 (N_10301,N_8035,N_8123);
and U10302 (N_10302,N_8952,N_8705);
or U10303 (N_10303,N_8399,N_7764);
nand U10304 (N_10304,N_8874,N_8252);
nand U10305 (N_10305,N_8511,N_7594);
or U10306 (N_10306,N_8478,N_8903);
nand U10307 (N_10307,N_8696,N_8467);
and U10308 (N_10308,N_7609,N_8632);
nand U10309 (N_10309,N_7615,N_7753);
or U10310 (N_10310,N_8006,N_8607);
nand U10311 (N_10311,N_7789,N_8206);
xnor U10312 (N_10312,N_8518,N_8185);
xor U10313 (N_10313,N_7512,N_7899);
and U10314 (N_10314,N_7632,N_8640);
and U10315 (N_10315,N_8953,N_8434);
or U10316 (N_10316,N_8381,N_8979);
nor U10317 (N_10317,N_8901,N_8680);
nand U10318 (N_10318,N_8254,N_8392);
nor U10319 (N_10319,N_8232,N_8984);
nand U10320 (N_10320,N_8510,N_8053);
nand U10321 (N_10321,N_8961,N_8071);
nor U10322 (N_10322,N_7550,N_8075);
or U10323 (N_10323,N_7925,N_8768);
nor U10324 (N_10324,N_8333,N_8269);
and U10325 (N_10325,N_7863,N_8201);
nand U10326 (N_10326,N_7850,N_7519);
and U10327 (N_10327,N_8517,N_8255);
or U10328 (N_10328,N_7880,N_8846);
or U10329 (N_10329,N_7938,N_8921);
xor U10330 (N_10330,N_8437,N_8406);
or U10331 (N_10331,N_8954,N_7934);
nand U10332 (N_10332,N_8741,N_7517);
or U10333 (N_10333,N_8448,N_8003);
and U10334 (N_10334,N_7619,N_8228);
nand U10335 (N_10335,N_7980,N_8409);
or U10336 (N_10336,N_7860,N_8101);
nor U10337 (N_10337,N_8330,N_7622);
nor U10338 (N_10338,N_8203,N_8728);
nand U10339 (N_10339,N_8412,N_7718);
or U10340 (N_10340,N_8953,N_8603);
or U10341 (N_10341,N_7919,N_7581);
nand U10342 (N_10342,N_8999,N_7675);
xnor U10343 (N_10343,N_8077,N_8237);
nor U10344 (N_10344,N_8292,N_8477);
nor U10345 (N_10345,N_8316,N_8031);
and U10346 (N_10346,N_8636,N_8317);
nor U10347 (N_10347,N_8108,N_8178);
or U10348 (N_10348,N_8974,N_8570);
or U10349 (N_10349,N_8352,N_7794);
nor U10350 (N_10350,N_8673,N_8657);
nand U10351 (N_10351,N_8708,N_8534);
xnor U10352 (N_10352,N_8312,N_7674);
or U10353 (N_10353,N_8923,N_8204);
xor U10354 (N_10354,N_8718,N_8116);
nand U10355 (N_10355,N_7603,N_7651);
or U10356 (N_10356,N_8631,N_7880);
and U10357 (N_10357,N_8383,N_8088);
or U10358 (N_10358,N_8028,N_8153);
nand U10359 (N_10359,N_7711,N_8020);
nor U10360 (N_10360,N_8204,N_8771);
and U10361 (N_10361,N_8354,N_8870);
nor U10362 (N_10362,N_7919,N_8420);
and U10363 (N_10363,N_7805,N_8329);
nand U10364 (N_10364,N_8407,N_8158);
or U10365 (N_10365,N_8654,N_8562);
and U10366 (N_10366,N_8982,N_7587);
and U10367 (N_10367,N_8173,N_8955);
or U10368 (N_10368,N_7556,N_8505);
xor U10369 (N_10369,N_7685,N_8806);
and U10370 (N_10370,N_8906,N_8157);
nand U10371 (N_10371,N_8265,N_8395);
or U10372 (N_10372,N_8464,N_8889);
and U10373 (N_10373,N_8928,N_8969);
nand U10374 (N_10374,N_8304,N_8624);
nor U10375 (N_10375,N_7981,N_7883);
or U10376 (N_10376,N_7915,N_7663);
or U10377 (N_10377,N_8077,N_8682);
or U10378 (N_10378,N_7696,N_8035);
or U10379 (N_10379,N_7542,N_8730);
and U10380 (N_10380,N_8751,N_8420);
nor U10381 (N_10381,N_8159,N_7640);
or U10382 (N_10382,N_7929,N_7581);
xnor U10383 (N_10383,N_8328,N_8003);
nor U10384 (N_10384,N_8914,N_7884);
nor U10385 (N_10385,N_7534,N_8245);
and U10386 (N_10386,N_8841,N_8170);
and U10387 (N_10387,N_8317,N_8634);
and U10388 (N_10388,N_7829,N_8551);
nand U10389 (N_10389,N_7873,N_8377);
xnor U10390 (N_10390,N_8878,N_8225);
and U10391 (N_10391,N_7551,N_8062);
or U10392 (N_10392,N_8318,N_8381);
and U10393 (N_10393,N_8164,N_7857);
or U10394 (N_10394,N_8193,N_7792);
and U10395 (N_10395,N_8613,N_8196);
and U10396 (N_10396,N_8356,N_7736);
nor U10397 (N_10397,N_8356,N_8754);
and U10398 (N_10398,N_8022,N_8463);
nor U10399 (N_10399,N_8854,N_8435);
xor U10400 (N_10400,N_8250,N_8624);
nand U10401 (N_10401,N_8332,N_8649);
nand U10402 (N_10402,N_8897,N_8114);
and U10403 (N_10403,N_7985,N_8463);
xor U10404 (N_10404,N_7533,N_8228);
nand U10405 (N_10405,N_8156,N_8270);
nor U10406 (N_10406,N_8725,N_8983);
nand U10407 (N_10407,N_8703,N_8696);
or U10408 (N_10408,N_7874,N_7941);
nor U10409 (N_10409,N_8893,N_7746);
and U10410 (N_10410,N_7877,N_7899);
and U10411 (N_10411,N_8999,N_7681);
xnor U10412 (N_10412,N_7879,N_8451);
and U10413 (N_10413,N_7604,N_8221);
and U10414 (N_10414,N_8199,N_8261);
xor U10415 (N_10415,N_7690,N_8786);
xnor U10416 (N_10416,N_7914,N_7588);
nand U10417 (N_10417,N_8727,N_8945);
nand U10418 (N_10418,N_8879,N_7888);
nor U10419 (N_10419,N_7808,N_7842);
or U10420 (N_10420,N_8737,N_7517);
and U10421 (N_10421,N_8919,N_8521);
and U10422 (N_10422,N_8020,N_7934);
nor U10423 (N_10423,N_8095,N_8323);
nor U10424 (N_10424,N_8810,N_8058);
nor U10425 (N_10425,N_8734,N_7592);
nor U10426 (N_10426,N_7554,N_8553);
or U10427 (N_10427,N_7576,N_8963);
nand U10428 (N_10428,N_8185,N_7530);
nand U10429 (N_10429,N_8325,N_8804);
xor U10430 (N_10430,N_8937,N_8208);
nand U10431 (N_10431,N_8613,N_7523);
nand U10432 (N_10432,N_8009,N_8967);
nor U10433 (N_10433,N_8886,N_7524);
nand U10434 (N_10434,N_8854,N_8456);
nor U10435 (N_10435,N_8952,N_7554);
or U10436 (N_10436,N_8787,N_8561);
and U10437 (N_10437,N_8954,N_8642);
nand U10438 (N_10438,N_8912,N_8806);
nor U10439 (N_10439,N_8244,N_8800);
and U10440 (N_10440,N_7507,N_8299);
or U10441 (N_10441,N_8311,N_8742);
xnor U10442 (N_10442,N_7790,N_8876);
nor U10443 (N_10443,N_7782,N_8181);
or U10444 (N_10444,N_8551,N_8914);
nor U10445 (N_10445,N_8672,N_8034);
and U10446 (N_10446,N_8002,N_7631);
nor U10447 (N_10447,N_8858,N_7767);
nand U10448 (N_10448,N_7651,N_7690);
and U10449 (N_10449,N_8247,N_7631);
nand U10450 (N_10450,N_8007,N_7584);
or U10451 (N_10451,N_8621,N_8916);
and U10452 (N_10452,N_7996,N_8457);
nor U10453 (N_10453,N_8596,N_8471);
xnor U10454 (N_10454,N_8625,N_7706);
nor U10455 (N_10455,N_7949,N_8835);
or U10456 (N_10456,N_7911,N_8340);
nand U10457 (N_10457,N_8134,N_7673);
or U10458 (N_10458,N_8091,N_8656);
xnor U10459 (N_10459,N_7812,N_8948);
or U10460 (N_10460,N_7750,N_7951);
xor U10461 (N_10461,N_8477,N_8407);
and U10462 (N_10462,N_7616,N_8749);
and U10463 (N_10463,N_7755,N_8684);
nand U10464 (N_10464,N_7915,N_8179);
nand U10465 (N_10465,N_8807,N_7800);
and U10466 (N_10466,N_7869,N_8068);
nor U10467 (N_10467,N_8073,N_7940);
xnor U10468 (N_10468,N_8363,N_7623);
or U10469 (N_10469,N_7509,N_8260);
or U10470 (N_10470,N_7994,N_7527);
nor U10471 (N_10471,N_8992,N_8064);
nor U10472 (N_10472,N_8528,N_8321);
nor U10473 (N_10473,N_8099,N_7701);
nand U10474 (N_10474,N_7695,N_7924);
nand U10475 (N_10475,N_8286,N_8517);
nor U10476 (N_10476,N_8727,N_8217);
or U10477 (N_10477,N_8991,N_7715);
and U10478 (N_10478,N_8953,N_7784);
and U10479 (N_10479,N_8418,N_7545);
or U10480 (N_10480,N_8847,N_7546);
and U10481 (N_10481,N_7710,N_7934);
nand U10482 (N_10482,N_7548,N_7913);
nor U10483 (N_10483,N_8271,N_8820);
nor U10484 (N_10484,N_8240,N_8247);
and U10485 (N_10485,N_7911,N_8686);
xor U10486 (N_10486,N_7954,N_8775);
or U10487 (N_10487,N_8438,N_7874);
and U10488 (N_10488,N_8552,N_8655);
xnor U10489 (N_10489,N_8854,N_7571);
or U10490 (N_10490,N_8174,N_8452);
nand U10491 (N_10491,N_8393,N_7698);
or U10492 (N_10492,N_7876,N_8373);
nand U10493 (N_10493,N_8807,N_8038);
or U10494 (N_10494,N_8635,N_8537);
nor U10495 (N_10495,N_7910,N_8924);
and U10496 (N_10496,N_8588,N_8047);
nor U10497 (N_10497,N_7615,N_8822);
nand U10498 (N_10498,N_7528,N_7614);
and U10499 (N_10499,N_8126,N_8992);
nand U10500 (N_10500,N_9555,N_10322);
or U10501 (N_10501,N_9028,N_10270);
nand U10502 (N_10502,N_10389,N_9043);
and U10503 (N_10503,N_9053,N_10498);
nor U10504 (N_10504,N_10196,N_9470);
or U10505 (N_10505,N_9133,N_9885);
and U10506 (N_10506,N_9360,N_10220);
and U10507 (N_10507,N_9515,N_9982);
and U10508 (N_10508,N_9729,N_10070);
nand U10509 (N_10509,N_9710,N_9206);
nand U10510 (N_10510,N_9665,N_10231);
nand U10511 (N_10511,N_10462,N_9613);
nor U10512 (N_10512,N_9277,N_9317);
nor U10513 (N_10513,N_9714,N_9839);
nor U10514 (N_10514,N_10272,N_10374);
nand U10515 (N_10515,N_10135,N_10364);
nand U10516 (N_10516,N_9962,N_9105);
or U10517 (N_10517,N_9732,N_9850);
nor U10518 (N_10518,N_10383,N_9436);
xor U10519 (N_10519,N_10012,N_9057);
or U10520 (N_10520,N_10044,N_9670);
xnor U10521 (N_10521,N_9611,N_10067);
nor U10522 (N_10522,N_9215,N_9622);
or U10523 (N_10523,N_9237,N_9516);
xnor U10524 (N_10524,N_9055,N_9848);
or U10525 (N_10525,N_9017,N_10485);
and U10526 (N_10526,N_9701,N_9987);
xor U10527 (N_10527,N_9617,N_9154);
or U10528 (N_10528,N_9468,N_10129);
nor U10529 (N_10529,N_10106,N_9199);
and U10530 (N_10530,N_10061,N_9740);
nor U10531 (N_10531,N_10042,N_10359);
nand U10532 (N_10532,N_10390,N_9928);
nor U10533 (N_10533,N_9148,N_9265);
nand U10534 (N_10534,N_9275,N_10217);
nand U10535 (N_10535,N_9218,N_10334);
nand U10536 (N_10536,N_10494,N_9464);
nand U10537 (N_10537,N_9172,N_9642);
or U10538 (N_10538,N_9669,N_9680);
and U10539 (N_10539,N_10266,N_9807);
nor U10540 (N_10540,N_9612,N_10232);
nand U10541 (N_10541,N_9441,N_9035);
and U10542 (N_10542,N_10090,N_9815);
or U10543 (N_10543,N_9245,N_10489);
nand U10544 (N_10544,N_10405,N_9200);
and U10545 (N_10545,N_9227,N_9633);
nor U10546 (N_10546,N_9262,N_9486);
and U10547 (N_10547,N_10013,N_9204);
or U10548 (N_10548,N_9306,N_9899);
or U10549 (N_10549,N_9523,N_9004);
nor U10550 (N_10550,N_9097,N_9968);
nand U10551 (N_10551,N_10078,N_10213);
nand U10552 (N_10552,N_9892,N_10077);
nor U10553 (N_10553,N_9062,N_10168);
nand U10554 (N_10554,N_10050,N_10165);
nor U10555 (N_10555,N_10252,N_9957);
xor U10556 (N_10556,N_10098,N_9726);
nor U10557 (N_10557,N_9514,N_9510);
nor U10558 (N_10558,N_9186,N_10195);
and U10559 (N_10559,N_9886,N_9312);
and U10560 (N_10560,N_10022,N_9346);
or U10561 (N_10561,N_10229,N_9361);
nand U10562 (N_10562,N_9111,N_10190);
or U10563 (N_10563,N_9537,N_9313);
nand U10564 (N_10564,N_9263,N_9679);
or U10565 (N_10565,N_9452,N_9945);
or U10566 (N_10566,N_9817,N_10162);
nand U10567 (N_10567,N_10166,N_10136);
nor U10568 (N_10568,N_10075,N_9616);
and U10569 (N_10569,N_9345,N_9458);
nor U10570 (N_10570,N_9884,N_9662);
nand U10571 (N_10571,N_9478,N_9251);
nand U10572 (N_10572,N_9634,N_9240);
nor U10573 (N_10573,N_9502,N_9503);
nor U10574 (N_10574,N_9750,N_10153);
nand U10575 (N_10575,N_10212,N_9309);
or U10576 (N_10576,N_9870,N_9337);
and U10577 (N_10577,N_9623,N_10149);
nand U10578 (N_10578,N_9910,N_10486);
nand U10579 (N_10579,N_9681,N_10309);
nor U10580 (N_10580,N_9585,N_9020);
nand U10581 (N_10581,N_9214,N_10036);
or U10582 (N_10582,N_10331,N_9042);
and U10583 (N_10583,N_10010,N_9751);
and U10584 (N_10584,N_9031,N_9040);
nor U10585 (N_10585,N_9619,N_9863);
nand U10586 (N_10586,N_9448,N_10219);
and U10587 (N_10587,N_10255,N_9404);
nor U10588 (N_10588,N_10385,N_10271);
xor U10589 (N_10589,N_9600,N_9134);
and U10590 (N_10590,N_9289,N_9354);
or U10591 (N_10591,N_10431,N_9904);
nand U10592 (N_10592,N_9326,N_10002);
xor U10593 (N_10593,N_9226,N_10296);
and U10594 (N_10594,N_9430,N_10436);
or U10595 (N_10595,N_10346,N_10257);
nand U10596 (N_10596,N_10282,N_9927);
nand U10597 (N_10597,N_9291,N_9121);
nand U10598 (N_10598,N_9953,N_9019);
or U10599 (N_10599,N_9718,N_9347);
or U10600 (N_10600,N_9694,N_9009);
nand U10601 (N_10601,N_9540,N_9217);
and U10602 (N_10602,N_9827,N_10244);
nor U10603 (N_10603,N_9089,N_9144);
and U10604 (N_10604,N_10267,N_10226);
or U10605 (N_10605,N_9706,N_10451);
nand U10606 (N_10606,N_10254,N_9435);
and U10607 (N_10607,N_9864,N_10315);
nor U10608 (N_10608,N_9270,N_9507);
nand U10609 (N_10609,N_10493,N_9985);
nand U10610 (N_10610,N_9654,N_10357);
nand U10611 (N_10611,N_9422,N_10068);
and U10612 (N_10612,N_9170,N_9488);
nor U10613 (N_10613,N_10102,N_9294);
nand U10614 (N_10614,N_9184,N_9806);
xor U10615 (N_10615,N_10201,N_9855);
nor U10616 (N_10616,N_9179,N_10120);
and U10617 (N_10617,N_10387,N_9010);
xnor U10618 (N_10618,N_10059,N_9846);
nor U10619 (N_10619,N_9090,N_9286);
and U10620 (N_10620,N_9770,N_10308);
xnor U10621 (N_10621,N_9152,N_10417);
nand U10622 (N_10622,N_9259,N_9618);
and U10623 (N_10623,N_10223,N_9842);
nand U10624 (N_10624,N_9446,N_9242);
xor U10625 (N_10625,N_9529,N_10432);
and U10626 (N_10626,N_10015,N_9857);
xor U10627 (N_10627,N_9194,N_9860);
and U10628 (N_10628,N_9657,N_10192);
nand U10629 (N_10629,N_10482,N_10341);
xnor U10630 (N_10630,N_9407,N_10142);
nor U10631 (N_10631,N_9224,N_9304);
xor U10632 (N_10632,N_10449,N_9691);
and U10633 (N_10633,N_10439,N_9584);
nor U10634 (N_10634,N_9508,N_9088);
or U10635 (N_10635,N_10178,N_9542);
or U10636 (N_10636,N_9548,N_9833);
or U10637 (N_10637,N_9971,N_9046);
nor U10638 (N_10638,N_10020,N_9742);
and U10639 (N_10639,N_10476,N_9673);
nor U10640 (N_10640,N_9812,N_10367);
and U10641 (N_10641,N_9069,N_9338);
nor U10642 (N_10642,N_10351,N_10285);
or U10643 (N_10643,N_10228,N_10128);
nand U10644 (N_10644,N_9257,N_10453);
nand U10645 (N_10645,N_10481,N_10048);
and U10646 (N_10646,N_9007,N_9798);
and U10647 (N_10647,N_10419,N_10450);
nor U10648 (N_10648,N_9961,N_10054);
nand U10649 (N_10649,N_10401,N_9038);
nand U10650 (N_10650,N_10366,N_9937);
nor U10651 (N_10651,N_9804,N_9450);
nor U10652 (N_10652,N_9522,N_9621);
and U10653 (N_10653,N_10009,N_9264);
nor U10654 (N_10654,N_9519,N_10193);
or U10655 (N_10655,N_10395,N_9014);
or U10656 (N_10656,N_10378,N_9072);
nor U10657 (N_10657,N_10248,N_9854);
and U10658 (N_10658,N_10421,N_10150);
nor U10659 (N_10659,N_9995,N_9965);
nand U10660 (N_10660,N_9279,N_9467);
or U10661 (N_10661,N_9760,N_9255);
and U10662 (N_10662,N_10053,N_10086);
nor U10663 (N_10663,N_10307,N_10400);
nand U10664 (N_10664,N_9856,N_10430);
or U10665 (N_10665,N_9387,N_9929);
and U10666 (N_10666,N_9689,N_10211);
nor U10667 (N_10667,N_9303,N_10454);
nor U10668 (N_10668,N_9849,N_9873);
nand U10669 (N_10669,N_9580,N_10353);
and U10670 (N_10670,N_10093,N_9058);
and U10671 (N_10671,N_10117,N_9820);
xor U10672 (N_10672,N_9177,N_9922);
nand U10673 (N_10673,N_9076,N_10208);
and U10674 (N_10674,N_9495,N_9274);
and U10675 (N_10675,N_9744,N_9250);
nand U10676 (N_10676,N_9321,N_10246);
or U10677 (N_10677,N_9518,N_9029);
nand U10678 (N_10678,N_10291,N_10202);
and U10679 (N_10679,N_9229,N_9119);
or U10680 (N_10680,N_9647,N_9541);
xnor U10681 (N_10681,N_10031,N_10371);
and U10682 (N_10682,N_10021,N_9244);
xor U10683 (N_10683,N_9801,N_9280);
or U10684 (N_10684,N_10377,N_9786);
nand U10685 (N_10685,N_9444,N_10392);
xor U10686 (N_10686,N_9759,N_10474);
nand U10687 (N_10687,N_9207,N_10260);
nand U10688 (N_10688,N_9233,N_10301);
xnor U10689 (N_10689,N_9341,N_9421);
nand U10690 (N_10690,N_9609,N_9941);
and U10691 (N_10691,N_9911,N_9986);
and U10692 (N_10692,N_10063,N_9512);
or U10693 (N_10693,N_9462,N_9728);
nand U10694 (N_10694,N_9324,N_9545);
and U10695 (N_10695,N_9693,N_10278);
or U10696 (N_10696,N_10235,N_10394);
and U10697 (N_10697,N_9165,N_9047);
or U10698 (N_10698,N_10163,N_9620);
nand U10699 (N_10699,N_9185,N_9389);
nand U10700 (N_10700,N_10052,N_10311);
nand U10701 (N_10701,N_10284,N_10115);
nand U10702 (N_10702,N_9946,N_10438);
or U10703 (N_10703,N_9091,N_10289);
nor U10704 (N_10704,N_9626,N_9077);
nand U10705 (N_10705,N_9586,N_9821);
nand U10706 (N_10706,N_9909,N_10473);
and U10707 (N_10707,N_10200,N_9339);
and U10708 (N_10708,N_9284,N_9330);
or U10709 (N_10709,N_10327,N_9060);
nor U10710 (N_10710,N_9591,N_9116);
nor U10711 (N_10711,N_9016,N_10380);
nor U10712 (N_10712,N_10411,N_9776);
xor U10713 (N_10713,N_10428,N_9638);
xnor U10714 (N_10714,N_9993,N_9045);
nor U10715 (N_10715,N_9103,N_10258);
or U10716 (N_10716,N_9107,N_9044);
nor U10717 (N_10717,N_10101,N_9766);
or U10718 (N_10718,N_9763,N_10001);
nor U10719 (N_10719,N_9325,N_9667);
or U10720 (N_10720,N_9805,N_10046);
nor U10721 (N_10721,N_9037,N_9906);
and U10722 (N_10722,N_9822,N_9695);
or U10723 (N_10723,N_10304,N_9323);
nand U10724 (N_10724,N_9533,N_9285);
and U10725 (N_10725,N_9506,N_9830);
and U10726 (N_10726,N_9717,N_9293);
nor U10727 (N_10727,N_9376,N_9219);
nand U10728 (N_10728,N_10256,N_10143);
or U10729 (N_10729,N_9923,N_9378);
nand U10730 (N_10730,N_9648,N_10137);
or U10731 (N_10731,N_10029,N_10424);
and U10732 (N_10732,N_9980,N_9383);
or U10733 (N_10733,N_9209,N_10250);
or U10734 (N_10734,N_9499,N_9705);
nor U10735 (N_10735,N_9132,N_10205);
nor U10736 (N_10736,N_9139,N_9003);
nor U10737 (N_10737,N_9746,N_9278);
nand U10738 (N_10738,N_9228,N_10434);
and U10739 (N_10739,N_9025,N_10003);
nand U10740 (N_10740,N_9108,N_10017);
and U10741 (N_10741,N_9774,N_9563);
nand U10742 (N_10742,N_9032,N_9001);
nand U10743 (N_10743,N_10122,N_9831);
xnor U10744 (N_10744,N_9550,N_9366);
nand U10745 (N_10745,N_10139,N_9949);
or U10746 (N_10746,N_9553,N_9015);
or U10747 (N_10747,N_9869,N_9160);
xor U10748 (N_10748,N_9178,N_10492);
or U10749 (N_10749,N_10455,N_9935);
nor U10750 (N_10750,N_10083,N_9725);
nor U10751 (N_10751,N_9465,N_10247);
xor U10752 (N_10752,N_10072,N_10466);
nand U10753 (N_10753,N_10373,N_9102);
nor U10754 (N_10754,N_9587,N_9865);
nand U10755 (N_10755,N_9656,N_10349);
nor U10756 (N_10756,N_9466,N_10119);
or U10757 (N_10757,N_9958,N_9417);
nand U10758 (N_10758,N_10147,N_10008);
nand U10759 (N_10759,N_9769,N_10241);
nand U10760 (N_10760,N_9546,N_9205);
and U10761 (N_10761,N_10306,N_9022);
nand U10762 (N_10762,N_10126,N_9943);
nand U10763 (N_10763,N_9399,N_9118);
and U10764 (N_10764,N_10495,N_9707);
nor U10765 (N_10765,N_9483,N_9527);
xnor U10766 (N_10766,N_9041,N_10207);
and U10767 (N_10767,N_9692,N_9790);
nor U10768 (N_10768,N_9268,N_9490);
nand U10769 (N_10769,N_9794,N_9329);
or U10770 (N_10770,N_9730,N_10032);
xnor U10771 (N_10771,N_9720,N_10300);
nor U10772 (N_10772,N_9898,N_9881);
or U10773 (N_10773,N_10314,N_10469);
or U10774 (N_10774,N_10375,N_9997);
nand U10775 (N_10775,N_9574,N_9445);
or U10776 (N_10776,N_9351,N_9409);
nor U10777 (N_10777,N_9595,N_10104);
nand U10778 (N_10778,N_10138,N_10082);
nand U10779 (N_10779,N_9547,N_9723);
nand U10780 (N_10780,N_10037,N_10172);
and U10781 (N_10781,N_9593,N_9627);
nand U10782 (N_10782,N_10110,N_10487);
and U10783 (N_10783,N_9646,N_10237);
and U10784 (N_10784,N_10189,N_9697);
or U10785 (N_10785,N_9597,N_10402);
nand U10786 (N_10786,N_9994,N_10006);
nand U10787 (N_10787,N_9168,N_10343);
nand U10788 (N_10788,N_9704,N_9114);
or U10789 (N_10789,N_10214,N_9355);
or U10790 (N_10790,N_10324,N_10362);
or U10791 (N_10791,N_10043,N_9400);
nand U10792 (N_10792,N_10016,N_10379);
or U10793 (N_10793,N_10345,N_9390);
and U10794 (N_10794,N_10496,N_9782);
and U10795 (N_10795,N_9123,N_9431);
or U10796 (N_10796,N_9933,N_10412);
nand U10797 (N_10797,N_9225,N_9727);
or U10798 (N_10798,N_9261,N_9938);
xor U10799 (N_10799,N_10161,N_9392);
or U10800 (N_10800,N_10151,N_10125);
and U10801 (N_10801,N_10121,N_9414);
nand U10802 (N_10802,N_9562,N_10381);
nor U10803 (N_10803,N_9582,N_9248);
or U10804 (N_10804,N_10339,N_9485);
or U10805 (N_10805,N_9979,N_10159);
or U10806 (N_10806,N_10164,N_10259);
nor U10807 (N_10807,N_9440,N_10415);
nand U10808 (N_10808,N_9298,N_9146);
nand U10809 (N_10809,N_10347,N_9137);
or U10810 (N_10810,N_9663,N_10410);
or U10811 (N_10811,N_9487,N_10361);
and U10812 (N_10812,N_9590,N_10234);
nand U10813 (N_10813,N_9283,N_9385);
or U10814 (N_10814,N_9579,N_9780);
or U10815 (N_10815,N_10095,N_10132);
or U10816 (N_10816,N_9398,N_9887);
nand U10817 (N_10817,N_9377,N_10169);
nand U10818 (N_10818,N_10464,N_10085);
nand U10819 (N_10819,N_9984,N_10127);
nor U10820 (N_10820,N_10092,N_9249);
nor U10821 (N_10821,N_9688,N_9074);
or U10822 (N_10822,N_9528,N_10338);
or U10823 (N_10823,N_10318,N_9629);
or U10824 (N_10824,N_9535,N_9916);
nand U10825 (N_10825,N_10414,N_9891);
nor U10826 (N_10826,N_9719,N_9188);
and U10827 (N_10827,N_10064,N_10108);
or U10828 (N_10828,N_10470,N_10317);
nand U10829 (N_10829,N_9424,N_9724);
xor U10830 (N_10830,N_10024,N_9155);
nor U10831 (N_10831,N_9388,N_9722);
or U10832 (N_10832,N_9405,N_9948);
and U10833 (N_10833,N_9491,N_10321);
and U10834 (N_10834,N_10174,N_9936);
nand U10835 (N_10835,N_10458,N_10388);
and U10836 (N_10836,N_10124,N_10484);
or U10837 (N_10837,N_9882,N_9308);
nor U10838 (N_10838,N_10177,N_9835);
or U10839 (N_10839,N_9628,N_9752);
or U10840 (N_10840,N_9824,N_9811);
or U10841 (N_10841,N_9650,N_9511);
or U10842 (N_10842,N_9415,N_9521);
xor U10843 (N_10843,N_10403,N_10263);
and U10844 (N_10844,N_9526,N_9189);
or U10845 (N_10845,N_9469,N_9454);
and U10846 (N_10846,N_9551,N_10183);
nand U10847 (N_10847,N_10471,N_9287);
nand U10848 (N_10848,N_10497,N_9051);
nor U10849 (N_10849,N_10134,N_9149);
nor U10850 (N_10850,N_9418,N_10397);
and U10851 (N_10851,N_9762,N_10283);
nor U10852 (N_10852,N_9826,N_9859);
or U10853 (N_10853,N_9434,N_9018);
nor U10854 (N_10854,N_9991,N_10055);
and U10855 (N_10855,N_9080,N_9307);
and U10856 (N_10856,N_10081,N_9645);
xnor U10857 (N_10857,N_9837,N_9156);
nor U10858 (N_10858,N_9034,N_9702);
or U10859 (N_10859,N_9344,N_9671);
or U10860 (N_10860,N_9903,N_9079);
and U10861 (N_10861,N_9216,N_9315);
and U10862 (N_10862,N_9158,N_9779);
and U10863 (N_10863,N_10176,N_9455);
nand U10864 (N_10864,N_9461,N_10230);
or U10865 (N_10865,N_9568,N_10198);
nand U10866 (N_10866,N_9247,N_10279);
nand U10867 (N_10867,N_10034,N_9482);
nor U10868 (N_10868,N_9592,N_9981);
and U10869 (N_10869,N_9808,N_9191);
or U10870 (N_10870,N_10365,N_10112);
or U10871 (N_10871,N_9397,N_9544);
or U10872 (N_10872,N_10038,N_9599);
xor U10873 (N_10873,N_10216,N_9713);
nor U10874 (N_10874,N_10039,N_9084);
and U10875 (N_10875,N_10281,N_9872);
nor U10876 (N_10876,N_9601,N_10144);
nor U10877 (N_10877,N_9411,N_10483);
and U10878 (N_10878,N_10107,N_10372);
and U10879 (N_10879,N_9637,N_9150);
and U10880 (N_10880,N_9739,N_9463);
or U10881 (N_10881,N_9099,N_9889);
nand U10882 (N_10882,N_10369,N_9425);
nand U10883 (N_10883,N_9024,N_10408);
or U10884 (N_10884,N_9708,N_9230);
or U10885 (N_10885,N_10264,N_9589);
xnor U10886 (N_10886,N_9311,N_10158);
nand U10887 (N_10887,N_9731,N_9061);
or U10888 (N_10888,N_9352,N_10344);
nor U10889 (N_10889,N_10005,N_9745);
and U10890 (N_10890,N_9552,N_10445);
and U10891 (N_10891,N_9788,N_9447);
nand U10892 (N_10892,N_9558,N_9484);
xnor U10893 (N_10893,N_9394,N_10251);
or U10894 (N_10894,N_9187,N_9554);
xnor U10895 (N_10895,N_10275,N_9819);
nor U10896 (N_10896,N_9059,N_10376);
nand U10897 (N_10897,N_9162,N_9078);
nand U10898 (N_10898,N_9813,N_10312);
or U10899 (N_10899,N_9145,N_9944);
nand U10900 (N_10900,N_10011,N_9687);
and U10901 (N_10901,N_9127,N_10167);
nor U10902 (N_10902,N_9380,N_9768);
and U10903 (N_10903,N_9333,N_10468);
and U10904 (N_10904,N_9988,N_10088);
xnor U10905 (N_10905,N_9320,N_10328);
xor U10906 (N_10906,N_9534,N_9142);
or U10907 (N_10907,N_10040,N_10243);
xnor U10908 (N_10908,N_10175,N_9932);
nand U10909 (N_10909,N_9234,N_10018);
or U10910 (N_10910,N_9532,N_9489);
and U10911 (N_10911,N_9026,N_9071);
or U10912 (N_10912,N_10459,N_10180);
and U10913 (N_10913,N_9070,N_10330);
or U10914 (N_10914,N_9963,N_9202);
and U10915 (N_10915,N_9841,N_9894);
nand U10916 (N_10916,N_9147,N_9565);
nor U10917 (N_10917,N_10360,N_9539);
and U10918 (N_10918,N_9931,N_10370);
nor U10919 (N_10919,N_9666,N_9777);
and U10920 (N_10920,N_9907,N_10416);
nor U10921 (N_10921,N_9747,N_9153);
nand U10922 (N_10922,N_9836,N_9169);
or U10923 (N_10923,N_9373,N_9743);
and U10924 (N_10924,N_9180,N_9793);
or U10925 (N_10925,N_10294,N_9810);
or U10926 (N_10926,N_9433,N_10096);
nand U10927 (N_10927,N_9260,N_10145);
or U10928 (N_10928,N_9136,N_10276);
or U10929 (N_10929,N_9082,N_9011);
xor U10930 (N_10930,N_10393,N_9143);
nor U10931 (N_10931,N_9192,N_9371);
and U10932 (N_10932,N_9379,N_9644);
nor U10933 (N_10933,N_10435,N_9602);
and U10934 (N_10934,N_9221,N_10225);
or U10935 (N_10935,N_9651,N_9951);
or U10936 (N_10936,N_10157,N_10221);
and U10937 (N_10937,N_10100,N_9068);
and U10938 (N_10938,N_9564,N_9998);
nand U10939 (N_10939,N_10491,N_9457);
nand U10940 (N_10940,N_10447,N_9640);
and U10941 (N_10941,N_9386,N_9176);
xor U10942 (N_10942,N_10184,N_10033);
and U10943 (N_10943,N_10027,N_9677);
and U10944 (N_10944,N_9791,N_9560);
nor U10945 (N_10945,N_9439,N_10350);
and U10946 (N_10946,N_10382,N_10472);
and U10947 (N_10947,N_9784,N_9749);
and U10948 (N_10948,N_9632,N_9851);
nand U10949 (N_10949,N_9874,N_9408);
nor U10950 (N_10950,N_9596,N_10261);
and U10951 (N_10951,N_9288,N_9615);
nor U10952 (N_10952,N_10280,N_9900);
and U10953 (N_10953,N_9427,N_10056);
and U10954 (N_10954,N_10062,N_9429);
or U10955 (N_10955,N_9924,N_9437);
or U10956 (N_10956,N_9631,N_9783);
xnor U10957 (N_10957,N_9258,N_9151);
nor U10958 (N_10958,N_9741,N_9343);
nand U10959 (N_10959,N_9847,N_9238);
or U10960 (N_10960,N_9736,N_9737);
and U10961 (N_10961,N_9109,N_10342);
xnor U10962 (N_10962,N_9348,N_9328);
or U10963 (N_10963,N_9124,N_9588);
nor U10964 (N_10964,N_10025,N_10477);
nor U10965 (N_10965,N_10118,N_10384);
nor U10966 (N_10966,N_9764,N_9253);
nand U10967 (N_10967,N_9456,N_10084);
or U10968 (N_10968,N_9384,N_10293);
or U10969 (N_10969,N_10303,N_9299);
and U10970 (N_10970,N_10467,N_9269);
nor U10971 (N_10971,N_9684,N_9748);
nor U10972 (N_10972,N_9138,N_9977);
nand U10973 (N_10973,N_9524,N_9173);
and U10974 (N_10974,N_9497,N_9403);
nand U10975 (N_10975,N_10295,N_9340);
nand U10976 (N_10976,N_9113,N_10049);
nand U10977 (N_10977,N_9712,N_9443);
nor U10978 (N_10978,N_9969,N_10335);
xor U10979 (N_10979,N_9525,N_10210);
nor U10980 (N_10980,N_9183,N_9252);
nand U10981 (N_10981,N_9879,N_9816);
nand U10982 (N_10982,N_9659,N_9067);
and U10983 (N_10983,N_9832,N_10404);
nor U10984 (N_10984,N_9370,N_9161);
nor U10985 (N_10985,N_9787,N_10222);
nor U10986 (N_10986,N_9083,N_9603);
and U10987 (N_10987,N_10181,N_9449);
or U10988 (N_10988,N_9543,N_10130);
nand U10989 (N_10989,N_9223,N_9190);
nor U10990 (N_10990,N_9419,N_9867);
or U10991 (N_10991,N_9319,N_9367);
and U10992 (N_10992,N_9033,N_9093);
nor U10993 (N_10993,N_10326,N_10057);
or U10994 (N_10994,N_9845,N_10490);
and U10995 (N_10995,N_9608,N_9880);
and U10996 (N_10996,N_9683,N_9063);
and U10997 (N_10997,N_9336,N_9085);
or U10998 (N_10998,N_9125,N_9301);
nand U10999 (N_10999,N_10045,N_9653);
nor U11000 (N_11000,N_9195,N_10074);
nand U11001 (N_11001,N_9501,N_9420);
or U11002 (N_11002,N_9364,N_9120);
and U11003 (N_11003,N_9048,N_9002);
or U11004 (N_11004,N_10305,N_9610);
nand U11005 (N_11005,N_10441,N_9362);
or U11006 (N_11006,N_9950,N_9175);
or U11007 (N_11007,N_9802,N_9871);
xor U11008 (N_11008,N_9754,N_10188);
nor U11009 (N_11009,N_9652,N_9635);
and U11010 (N_11010,N_9716,N_9901);
nand U11011 (N_11011,N_9682,N_10116);
nand U11012 (N_11012,N_9363,N_10480);
nor U11013 (N_11013,N_9734,N_9416);
and U11014 (N_11014,N_9598,N_10273);
or U11015 (N_11015,N_9231,N_10268);
or U11016 (N_11016,N_9013,N_10386);
or U11017 (N_11017,N_10197,N_10245);
nand U11018 (N_11018,N_9914,N_9800);
nand U11019 (N_11019,N_9919,N_9709);
nor U11020 (N_11020,N_9272,N_9171);
nor U11021 (N_11021,N_9908,N_10155);
or U11022 (N_11022,N_9104,N_10329);
or U11023 (N_11023,N_9735,N_9331);
nor U11024 (N_11024,N_9008,N_9853);
nor U11025 (N_11025,N_10433,N_9092);
or U11026 (N_11026,N_9239,N_10060);
nand U11027 (N_11027,N_9686,N_9428);
and U11028 (N_11028,N_9630,N_10313);
and U11029 (N_11029,N_9027,N_10409);
nand U11030 (N_11030,N_9825,N_9267);
xnor U11031 (N_11031,N_9604,N_9757);
and U11032 (N_11032,N_9246,N_9624);
and U11033 (N_11033,N_9607,N_9471);
nand U11034 (N_11034,N_9792,N_10156);
and U11035 (N_11035,N_9711,N_10336);
nor U11036 (N_11036,N_9594,N_9054);
xor U11037 (N_11037,N_9915,N_9005);
or U11038 (N_11038,N_9868,N_9858);
and U11039 (N_11039,N_10004,N_9122);
xor U11040 (N_11040,N_10087,N_9517);
nor U11041 (N_11041,N_10058,N_10499);
nand U11042 (N_11042,N_9942,N_10422);
and U11043 (N_11043,N_10356,N_10091);
nand U11044 (N_11044,N_10363,N_9789);
or U11045 (N_11045,N_9295,N_9636);
nor U11046 (N_11046,N_9834,N_9327);
nor U11047 (N_11047,N_9006,N_9476);
nand U11048 (N_11048,N_9081,N_9030);
nor U11049 (N_11049,N_9844,N_9256);
nand U11050 (N_11050,N_10028,N_10269);
and U11051 (N_11051,N_9576,N_9130);
xnor U11052 (N_11052,N_9381,N_10277);
nor U11053 (N_11053,N_9890,N_9065);
nand U11054 (N_11054,N_9128,N_9012);
and U11055 (N_11055,N_9966,N_9575);
nand U11056 (N_11056,N_9096,N_9531);
or U11057 (N_11057,N_9561,N_10302);
and U11058 (N_11058,N_9573,N_9322);
or U11059 (N_11059,N_9164,N_9318);
nor U11060 (N_11060,N_10286,N_10456);
or U11061 (N_11061,N_10240,N_9947);
nand U11062 (N_11062,N_9755,N_10133);
or U11063 (N_11063,N_10103,N_9182);
nand U11064 (N_11064,N_10080,N_9992);
nor U11065 (N_11065,N_10368,N_10154);
xor U11066 (N_11066,N_10348,N_9395);
nand U11067 (N_11067,N_9955,N_9472);
nand U11068 (N_11068,N_9773,N_9438);
nand U11069 (N_11069,N_9368,N_9193);
or U11070 (N_11070,N_9583,N_10000);
or U11071 (N_11071,N_9129,N_9674);
nor U11072 (N_11072,N_9316,N_9110);
and U11073 (N_11073,N_9174,N_10236);
nand U11074 (N_11074,N_9453,N_10292);
nor U11075 (N_11075,N_10463,N_9852);
nor U11076 (N_11076,N_10274,N_10413);
or U11077 (N_11077,N_9412,N_9357);
or U11078 (N_11078,N_10007,N_10140);
or U11079 (N_11079,N_9897,N_10023);
and U11080 (N_11080,N_9964,N_10239);
nor U11081 (N_11081,N_10340,N_9668);
or U11082 (N_11082,N_9799,N_9649);
nor U11083 (N_11083,N_9690,N_9396);
xnor U11084 (N_11084,N_9232,N_9862);
or U11085 (N_11085,N_10465,N_10051);
nor U11086 (N_11086,N_9557,N_10242);
or U11087 (N_11087,N_10191,N_9115);
nor U11088 (N_11088,N_9960,N_9999);
and U11089 (N_11089,N_9996,N_9775);
and U11090 (N_11090,N_9895,N_10396);
or U11091 (N_11091,N_9342,N_9235);
or U11092 (N_11092,N_10475,N_10203);
and U11093 (N_11093,N_9814,N_10109);
or U11094 (N_11094,N_9661,N_9492);
nor U11095 (N_11095,N_9967,N_9877);
or U11096 (N_11096,N_9520,N_9167);
or U11097 (N_11097,N_9201,N_9513);
and U11098 (N_11098,N_9369,N_9181);
or U11099 (N_11099,N_9254,N_9460);
nor U11100 (N_11100,N_9073,N_9410);
and U11101 (N_11101,N_9530,N_10337);
and U11102 (N_11102,N_10186,N_10290);
nand U11103 (N_11103,N_10148,N_10448);
nor U11104 (N_11104,N_9570,N_9210);
nand U11105 (N_11105,N_10047,N_9442);
nor U11106 (N_11106,N_10488,N_10094);
or U11107 (N_11107,N_9930,N_10206);
nor U11108 (N_11108,N_10238,N_10079);
nor U11109 (N_11109,N_9625,N_9296);
nor U11110 (N_11110,N_9578,N_9567);
and U11111 (N_11111,N_9393,N_9926);
and U11112 (N_11112,N_10209,N_9796);
nor U11113 (N_11113,N_9606,N_9538);
nor U11114 (N_11114,N_9353,N_9477);
or U11115 (N_11115,N_10297,N_9498);
nand U11116 (N_11116,N_9785,N_9356);
nand U11117 (N_11117,N_9056,N_10073);
nand U11118 (N_11118,N_10333,N_10406);
nor U11119 (N_11119,N_9838,N_10407);
xnor U11120 (N_11120,N_9925,N_9413);
nand U11121 (N_11121,N_9402,N_10187);
and U11122 (N_11122,N_9459,N_9496);
or U11123 (N_11123,N_9241,N_9700);
or U11124 (N_11124,N_9039,N_10316);
or U11125 (N_11125,N_9696,N_9141);
nand U11126 (N_11126,N_9305,N_10041);
and U11127 (N_11127,N_10170,N_9577);
nand U11128 (N_11128,N_9672,N_9699);
or U11129 (N_11129,N_9423,N_9212);
nor U11130 (N_11130,N_10099,N_9050);
xor U11131 (N_11131,N_10440,N_9896);
nor U11132 (N_11132,N_10425,N_9198);
nand U11133 (N_11133,N_9698,N_9920);
or U11134 (N_11134,N_9883,N_9509);
and U11135 (N_11135,N_9271,N_9350);
or U11136 (N_11136,N_10452,N_9117);
nand U11137 (N_11137,N_9952,N_9823);
nand U11138 (N_11138,N_9983,N_9281);
nor U11139 (N_11139,N_10423,N_9131);
and U11140 (N_11140,N_9536,N_9222);
and U11141 (N_11141,N_9297,N_9818);
nor U11142 (N_11142,N_10227,N_9314);
or U11143 (N_11143,N_9087,N_9614);
nand U11144 (N_11144,N_9781,N_9655);
or U11145 (N_11145,N_9213,N_9106);
xor U11146 (N_11146,N_9976,N_9276);
xor U11147 (N_11147,N_9211,N_9100);
or U11148 (N_11148,N_9203,N_10426);
nor U11149 (N_11149,N_10026,N_10019);
and U11150 (N_11150,N_9473,N_9166);
nor U11151 (N_11151,N_10089,N_9721);
and U11152 (N_11152,N_9391,N_9126);
xor U11153 (N_11153,N_10182,N_9359);
and U11154 (N_11154,N_9112,N_9406);
nor U11155 (N_11155,N_9989,N_9480);
nand U11156 (N_11156,N_10332,N_9843);
nor U11157 (N_11157,N_9266,N_9157);
xor U11158 (N_11158,N_9021,N_10310);
xor U11159 (N_11159,N_9715,N_9738);
nand U11160 (N_11160,N_9220,N_9335);
and U11161 (N_11161,N_10131,N_9052);
and U11162 (N_11162,N_9098,N_9678);
or U11163 (N_11163,N_10444,N_9605);
or U11164 (N_11164,N_10354,N_9196);
nor U11165 (N_11165,N_9236,N_9956);
and U11166 (N_11166,N_10194,N_9475);
or U11167 (N_11167,N_10418,N_9197);
xnor U11168 (N_11168,N_9829,N_10160);
xor U11169 (N_11169,N_9703,N_10179);
nand U11170 (N_11170,N_10113,N_9135);
or U11171 (N_11171,N_9401,N_9893);
or U11172 (N_11172,N_10443,N_10262);
and U11173 (N_11173,N_9494,N_10218);
nor U11174 (N_11174,N_9876,N_10111);
or U11175 (N_11175,N_9685,N_10429);
nand U11176 (N_11176,N_10420,N_9332);
nand U11177 (N_11177,N_10358,N_9761);
nor U11178 (N_11178,N_10355,N_9481);
or U11179 (N_11179,N_9140,N_10442);
and U11180 (N_11180,N_10287,N_9767);
nand U11181 (N_11181,N_9095,N_9959);
nand U11182 (N_11182,N_10427,N_9066);
nand U11183 (N_11183,N_10265,N_10457);
and U11184 (N_11184,N_9572,N_9372);
nand U11185 (N_11185,N_9972,N_9375);
nor U11186 (N_11186,N_9094,N_9493);
and U11187 (N_11187,N_9795,N_10065);
and U11188 (N_11188,N_9905,N_10391);
and U11189 (N_11189,N_10097,N_9809);
nand U11190 (N_11190,N_10105,N_9840);
nand U11191 (N_11191,N_10398,N_9451);
and U11192 (N_11192,N_9075,N_10224);
xnor U11193 (N_11193,N_9374,N_9049);
nand U11194 (N_11194,N_9753,N_9676);
nand U11195 (N_11195,N_9292,N_9349);
nand U11196 (N_11196,N_9756,N_10399);
nand U11197 (N_11197,N_10298,N_9549);
and U11198 (N_11198,N_10076,N_10071);
nand U11199 (N_11199,N_9771,N_9365);
or U11200 (N_11200,N_10066,N_9866);
and U11201 (N_11201,N_10199,N_9973);
nand U11202 (N_11202,N_9086,N_9975);
or U11203 (N_11203,N_9675,N_9664);
and U11204 (N_11204,N_9300,N_9559);
or U11205 (N_11205,N_10253,N_9643);
or U11206 (N_11206,N_9282,N_9159);
nand U11207 (N_11207,N_9569,N_9334);
nor U11208 (N_11208,N_9064,N_10030);
or U11209 (N_11209,N_9970,N_9036);
nor U11210 (N_11210,N_9913,N_9556);
and U11211 (N_11211,N_10233,N_10460);
and U11212 (N_11212,N_9978,N_9243);
xor U11213 (N_11213,N_9581,N_9934);
nand U11214 (N_11214,N_10035,N_10299);
nand U11215 (N_11215,N_9912,N_9290);
or U11216 (N_11216,N_10437,N_9504);
or U11217 (N_11217,N_10173,N_9733);
xnor U11218 (N_11218,N_9302,N_10461);
nand U11219 (N_11219,N_9658,N_9639);
or U11220 (N_11220,N_9875,N_10215);
nor U11221 (N_11221,N_9000,N_10288);
or U11222 (N_11222,N_9163,N_9990);
nand U11223 (N_11223,N_9902,N_9772);
and U11224 (N_11224,N_9566,N_10141);
nand U11225 (N_11225,N_10446,N_9101);
xnor U11226 (N_11226,N_9939,N_10352);
nand U11227 (N_11227,N_9954,N_10123);
and U11228 (N_11228,N_9432,N_10478);
nand U11229 (N_11229,N_9474,N_9940);
xor U11230 (N_11230,N_9310,N_9917);
or U11231 (N_11231,N_9778,N_9505);
xor U11232 (N_11232,N_10114,N_9758);
and U11233 (N_11233,N_9921,N_10320);
nor U11234 (N_11234,N_9479,N_10479);
nor U11235 (N_11235,N_10069,N_9273);
nand U11236 (N_11236,N_10146,N_9974);
nor U11237 (N_11237,N_10014,N_9571);
or U11238 (N_11238,N_9918,N_9500);
or U11239 (N_11239,N_9023,N_9765);
or U11240 (N_11240,N_10325,N_9382);
nand U11241 (N_11241,N_9878,N_10249);
and U11242 (N_11242,N_9426,N_9861);
nor U11243 (N_11243,N_10204,N_9828);
nor U11244 (N_11244,N_10319,N_9797);
xnor U11245 (N_11245,N_9888,N_10185);
nand U11246 (N_11246,N_10171,N_9641);
nand U11247 (N_11247,N_10323,N_9358);
xnor U11248 (N_11248,N_9803,N_9660);
nand U11249 (N_11249,N_9208,N_10152);
or U11250 (N_11250,N_9696,N_9700);
nand U11251 (N_11251,N_10264,N_10413);
nor U11252 (N_11252,N_9152,N_9998);
xnor U11253 (N_11253,N_10308,N_10387);
and U11254 (N_11254,N_10497,N_9262);
xor U11255 (N_11255,N_9787,N_9952);
nand U11256 (N_11256,N_9098,N_9394);
xnor U11257 (N_11257,N_9778,N_9682);
or U11258 (N_11258,N_9184,N_10432);
and U11259 (N_11259,N_9074,N_10244);
or U11260 (N_11260,N_9575,N_10083);
nand U11261 (N_11261,N_10037,N_9906);
nand U11262 (N_11262,N_9462,N_9937);
nand U11263 (N_11263,N_10329,N_9827);
and U11264 (N_11264,N_9251,N_9973);
and U11265 (N_11265,N_9950,N_10471);
or U11266 (N_11266,N_9176,N_9654);
xor U11267 (N_11267,N_10429,N_10492);
and U11268 (N_11268,N_9967,N_9617);
and U11269 (N_11269,N_9954,N_10065);
xnor U11270 (N_11270,N_9444,N_10332);
or U11271 (N_11271,N_9270,N_9774);
nor U11272 (N_11272,N_10081,N_9580);
nor U11273 (N_11273,N_9809,N_9856);
or U11274 (N_11274,N_9477,N_9724);
or U11275 (N_11275,N_10179,N_9418);
nand U11276 (N_11276,N_10220,N_9601);
and U11277 (N_11277,N_9528,N_9510);
or U11278 (N_11278,N_9695,N_9737);
nor U11279 (N_11279,N_9097,N_9522);
or U11280 (N_11280,N_10035,N_9483);
nor U11281 (N_11281,N_9074,N_10124);
and U11282 (N_11282,N_9226,N_9362);
nand U11283 (N_11283,N_9447,N_9085);
and U11284 (N_11284,N_9119,N_10065);
nor U11285 (N_11285,N_9553,N_10374);
and U11286 (N_11286,N_9306,N_9412);
xnor U11287 (N_11287,N_9643,N_9964);
or U11288 (N_11288,N_9874,N_9370);
nor U11289 (N_11289,N_10262,N_10033);
or U11290 (N_11290,N_10070,N_9298);
nand U11291 (N_11291,N_9711,N_9395);
nand U11292 (N_11292,N_10336,N_9761);
and U11293 (N_11293,N_9335,N_9217);
nor U11294 (N_11294,N_9439,N_9461);
and U11295 (N_11295,N_9747,N_9913);
nand U11296 (N_11296,N_9888,N_9771);
nand U11297 (N_11297,N_9370,N_10250);
and U11298 (N_11298,N_9634,N_9988);
and U11299 (N_11299,N_9345,N_9892);
and U11300 (N_11300,N_10248,N_10457);
or U11301 (N_11301,N_9989,N_9795);
and U11302 (N_11302,N_9249,N_9455);
or U11303 (N_11303,N_9611,N_10399);
and U11304 (N_11304,N_9237,N_10058);
nand U11305 (N_11305,N_9682,N_9848);
or U11306 (N_11306,N_9540,N_9866);
xnor U11307 (N_11307,N_9227,N_9290);
nand U11308 (N_11308,N_10455,N_9288);
xnor U11309 (N_11309,N_10026,N_9874);
xnor U11310 (N_11310,N_9327,N_9310);
nand U11311 (N_11311,N_10242,N_9113);
nor U11312 (N_11312,N_10209,N_9567);
nand U11313 (N_11313,N_9187,N_10462);
or U11314 (N_11314,N_9423,N_9523);
or U11315 (N_11315,N_9939,N_10487);
and U11316 (N_11316,N_9525,N_9266);
and U11317 (N_11317,N_9598,N_10270);
nor U11318 (N_11318,N_9894,N_9281);
nor U11319 (N_11319,N_10450,N_10300);
and U11320 (N_11320,N_10069,N_10009);
xnor U11321 (N_11321,N_9110,N_10048);
or U11322 (N_11322,N_10464,N_9290);
and U11323 (N_11323,N_9776,N_9831);
xnor U11324 (N_11324,N_9093,N_10294);
or U11325 (N_11325,N_10341,N_9005);
nand U11326 (N_11326,N_9471,N_9051);
xnor U11327 (N_11327,N_9496,N_10413);
nand U11328 (N_11328,N_10074,N_10219);
nand U11329 (N_11329,N_9299,N_9772);
nor U11330 (N_11330,N_9241,N_9163);
nand U11331 (N_11331,N_10358,N_10015);
and U11332 (N_11332,N_10142,N_10021);
nand U11333 (N_11333,N_9617,N_9321);
nand U11334 (N_11334,N_10215,N_9513);
nor U11335 (N_11335,N_10240,N_9744);
xor U11336 (N_11336,N_10438,N_9657);
nor U11337 (N_11337,N_9541,N_10437);
nor U11338 (N_11338,N_9435,N_9432);
nand U11339 (N_11339,N_9240,N_10175);
xor U11340 (N_11340,N_9420,N_10162);
nand U11341 (N_11341,N_10307,N_9613);
and U11342 (N_11342,N_10123,N_9906);
or U11343 (N_11343,N_9348,N_9018);
or U11344 (N_11344,N_9077,N_9578);
and U11345 (N_11345,N_9114,N_9974);
nand U11346 (N_11346,N_9191,N_9294);
xor U11347 (N_11347,N_10040,N_9666);
or U11348 (N_11348,N_10092,N_9086);
nor U11349 (N_11349,N_9901,N_9404);
nor U11350 (N_11350,N_9619,N_10148);
and U11351 (N_11351,N_9968,N_9004);
or U11352 (N_11352,N_9804,N_10034);
or U11353 (N_11353,N_9212,N_9262);
and U11354 (N_11354,N_9169,N_9042);
nor U11355 (N_11355,N_9859,N_9035);
nand U11356 (N_11356,N_9625,N_9979);
nor U11357 (N_11357,N_10401,N_9344);
and U11358 (N_11358,N_9357,N_10126);
and U11359 (N_11359,N_10043,N_9249);
or U11360 (N_11360,N_9119,N_9592);
or U11361 (N_11361,N_9055,N_10353);
or U11362 (N_11362,N_10495,N_9660);
nand U11363 (N_11363,N_10233,N_9820);
nor U11364 (N_11364,N_9245,N_9581);
nor U11365 (N_11365,N_9293,N_10422);
xor U11366 (N_11366,N_9508,N_9912);
or U11367 (N_11367,N_9930,N_10226);
or U11368 (N_11368,N_10421,N_9536);
and U11369 (N_11369,N_10221,N_10340);
xor U11370 (N_11370,N_10369,N_9887);
nor U11371 (N_11371,N_9901,N_10011);
and U11372 (N_11372,N_10311,N_9796);
and U11373 (N_11373,N_9212,N_9062);
nor U11374 (N_11374,N_9582,N_9054);
and U11375 (N_11375,N_9242,N_10437);
nand U11376 (N_11376,N_9604,N_9814);
nor U11377 (N_11377,N_9171,N_10120);
xnor U11378 (N_11378,N_9114,N_10190);
and U11379 (N_11379,N_9097,N_9137);
or U11380 (N_11380,N_9479,N_9033);
or U11381 (N_11381,N_9478,N_10216);
or U11382 (N_11382,N_9678,N_9739);
or U11383 (N_11383,N_9133,N_10344);
nand U11384 (N_11384,N_9740,N_9763);
nor U11385 (N_11385,N_10270,N_10334);
and U11386 (N_11386,N_10269,N_9104);
and U11387 (N_11387,N_10499,N_9791);
nand U11388 (N_11388,N_10296,N_9334);
xnor U11389 (N_11389,N_9894,N_9914);
and U11390 (N_11390,N_10440,N_9543);
xnor U11391 (N_11391,N_10405,N_10184);
and U11392 (N_11392,N_10073,N_10210);
or U11393 (N_11393,N_9186,N_9494);
nand U11394 (N_11394,N_9373,N_9961);
or U11395 (N_11395,N_9800,N_9709);
and U11396 (N_11396,N_9470,N_9069);
nand U11397 (N_11397,N_9071,N_9542);
and U11398 (N_11398,N_9359,N_10427);
xnor U11399 (N_11399,N_9670,N_9087);
nand U11400 (N_11400,N_9302,N_10197);
or U11401 (N_11401,N_9284,N_9797);
or U11402 (N_11402,N_9130,N_10471);
and U11403 (N_11403,N_9544,N_10318);
and U11404 (N_11404,N_9660,N_9048);
nand U11405 (N_11405,N_10470,N_10264);
and U11406 (N_11406,N_9149,N_10384);
or U11407 (N_11407,N_9167,N_10353);
and U11408 (N_11408,N_9591,N_10317);
or U11409 (N_11409,N_9313,N_10215);
or U11410 (N_11410,N_9801,N_9365);
nor U11411 (N_11411,N_9215,N_10287);
xor U11412 (N_11412,N_10030,N_9781);
or U11413 (N_11413,N_9623,N_10283);
nand U11414 (N_11414,N_9934,N_9535);
and U11415 (N_11415,N_9172,N_10164);
nor U11416 (N_11416,N_9520,N_10408);
nand U11417 (N_11417,N_9928,N_10181);
and U11418 (N_11418,N_9422,N_9158);
or U11419 (N_11419,N_9235,N_9781);
nor U11420 (N_11420,N_10195,N_9459);
and U11421 (N_11421,N_10185,N_9266);
nand U11422 (N_11422,N_10200,N_9184);
nor U11423 (N_11423,N_10117,N_9660);
nor U11424 (N_11424,N_9748,N_10157);
nor U11425 (N_11425,N_10370,N_10215);
and U11426 (N_11426,N_9595,N_10053);
xor U11427 (N_11427,N_10347,N_10149);
nand U11428 (N_11428,N_9449,N_9980);
nor U11429 (N_11429,N_9226,N_10428);
nand U11430 (N_11430,N_9202,N_9324);
nor U11431 (N_11431,N_9901,N_9727);
xnor U11432 (N_11432,N_10182,N_9083);
or U11433 (N_11433,N_9604,N_9748);
nand U11434 (N_11434,N_9069,N_9974);
xor U11435 (N_11435,N_10454,N_10374);
and U11436 (N_11436,N_10075,N_9527);
nor U11437 (N_11437,N_10436,N_9844);
nand U11438 (N_11438,N_9664,N_10464);
xor U11439 (N_11439,N_9863,N_10027);
and U11440 (N_11440,N_10201,N_9861);
or U11441 (N_11441,N_9462,N_10160);
or U11442 (N_11442,N_9450,N_10072);
and U11443 (N_11443,N_9577,N_9358);
and U11444 (N_11444,N_9239,N_9945);
or U11445 (N_11445,N_9461,N_9660);
nand U11446 (N_11446,N_10091,N_9268);
or U11447 (N_11447,N_10070,N_9804);
or U11448 (N_11448,N_9491,N_9380);
nor U11449 (N_11449,N_9641,N_9209);
nand U11450 (N_11450,N_9294,N_9747);
xnor U11451 (N_11451,N_10391,N_9865);
nor U11452 (N_11452,N_9853,N_9047);
or U11453 (N_11453,N_10039,N_9103);
nand U11454 (N_11454,N_10285,N_9044);
nand U11455 (N_11455,N_9128,N_9685);
nand U11456 (N_11456,N_10391,N_9670);
and U11457 (N_11457,N_9186,N_9888);
or U11458 (N_11458,N_9216,N_10214);
nand U11459 (N_11459,N_10043,N_10243);
and U11460 (N_11460,N_10042,N_9251);
and U11461 (N_11461,N_10492,N_9235);
nand U11462 (N_11462,N_10254,N_9038);
nand U11463 (N_11463,N_9711,N_10386);
or U11464 (N_11464,N_9511,N_9743);
and U11465 (N_11465,N_9567,N_9334);
and U11466 (N_11466,N_9789,N_9163);
nand U11467 (N_11467,N_9327,N_9666);
nand U11468 (N_11468,N_9513,N_10258);
or U11469 (N_11469,N_9091,N_9403);
and U11470 (N_11470,N_9620,N_9630);
nand U11471 (N_11471,N_9804,N_9420);
nor U11472 (N_11472,N_10444,N_10228);
or U11473 (N_11473,N_10442,N_10245);
nand U11474 (N_11474,N_9809,N_9263);
and U11475 (N_11475,N_9907,N_9827);
nand U11476 (N_11476,N_10051,N_9686);
nor U11477 (N_11477,N_9415,N_9405);
or U11478 (N_11478,N_10348,N_9228);
nand U11479 (N_11479,N_9224,N_10108);
and U11480 (N_11480,N_9857,N_9007);
nand U11481 (N_11481,N_9151,N_9648);
or U11482 (N_11482,N_9233,N_10030);
or U11483 (N_11483,N_9794,N_9889);
nor U11484 (N_11484,N_10295,N_9202);
nand U11485 (N_11485,N_9968,N_9624);
and U11486 (N_11486,N_9116,N_9080);
nor U11487 (N_11487,N_10234,N_9500);
or U11488 (N_11488,N_9051,N_9440);
xnor U11489 (N_11489,N_9603,N_9545);
or U11490 (N_11490,N_9545,N_9119);
or U11491 (N_11491,N_10092,N_9553);
nor U11492 (N_11492,N_10376,N_9896);
or U11493 (N_11493,N_9247,N_10123);
and U11494 (N_11494,N_10415,N_10342);
nor U11495 (N_11495,N_9864,N_9195);
and U11496 (N_11496,N_9307,N_10250);
nor U11497 (N_11497,N_10136,N_9543);
or U11498 (N_11498,N_10273,N_10320);
or U11499 (N_11499,N_9476,N_10345);
nand U11500 (N_11500,N_10274,N_10026);
nor U11501 (N_11501,N_10047,N_10098);
nand U11502 (N_11502,N_10095,N_9295);
nand U11503 (N_11503,N_9298,N_9481);
or U11504 (N_11504,N_9846,N_9860);
or U11505 (N_11505,N_9617,N_9258);
nor U11506 (N_11506,N_9232,N_9790);
or U11507 (N_11507,N_9662,N_10250);
or U11508 (N_11508,N_10025,N_9481);
or U11509 (N_11509,N_9483,N_9769);
xnor U11510 (N_11510,N_10069,N_9661);
nor U11511 (N_11511,N_9990,N_9034);
nand U11512 (N_11512,N_9687,N_9613);
nor U11513 (N_11513,N_9119,N_9944);
and U11514 (N_11514,N_10454,N_9181);
nand U11515 (N_11515,N_9127,N_9769);
nand U11516 (N_11516,N_9904,N_9108);
or U11517 (N_11517,N_10092,N_9021);
nand U11518 (N_11518,N_9669,N_10461);
nand U11519 (N_11519,N_10312,N_10322);
nand U11520 (N_11520,N_10207,N_10275);
and U11521 (N_11521,N_9301,N_9094);
and U11522 (N_11522,N_9941,N_10081);
and U11523 (N_11523,N_9957,N_9759);
nand U11524 (N_11524,N_9925,N_9933);
or U11525 (N_11525,N_9005,N_9702);
and U11526 (N_11526,N_9100,N_9931);
or U11527 (N_11527,N_10448,N_10283);
and U11528 (N_11528,N_9041,N_9834);
or U11529 (N_11529,N_9537,N_10191);
nor U11530 (N_11530,N_10447,N_10419);
nor U11531 (N_11531,N_9314,N_9525);
nand U11532 (N_11532,N_10099,N_9911);
nor U11533 (N_11533,N_10204,N_10324);
or U11534 (N_11534,N_9451,N_9271);
or U11535 (N_11535,N_9871,N_9134);
or U11536 (N_11536,N_9151,N_10229);
nand U11537 (N_11537,N_9421,N_10401);
nor U11538 (N_11538,N_9966,N_9115);
xnor U11539 (N_11539,N_9416,N_9731);
nor U11540 (N_11540,N_9598,N_9993);
and U11541 (N_11541,N_10194,N_9227);
or U11542 (N_11542,N_9816,N_10360);
or U11543 (N_11543,N_9531,N_9169);
xor U11544 (N_11544,N_9686,N_9021);
nor U11545 (N_11545,N_10383,N_9883);
nand U11546 (N_11546,N_9863,N_9937);
or U11547 (N_11547,N_9718,N_9160);
xnor U11548 (N_11548,N_9956,N_9142);
xnor U11549 (N_11549,N_9483,N_9134);
nor U11550 (N_11550,N_10123,N_9085);
nand U11551 (N_11551,N_9417,N_9182);
nand U11552 (N_11552,N_10019,N_10200);
and U11553 (N_11553,N_9347,N_9698);
and U11554 (N_11554,N_9793,N_9757);
or U11555 (N_11555,N_9033,N_9615);
or U11556 (N_11556,N_10224,N_10396);
and U11557 (N_11557,N_9985,N_9528);
or U11558 (N_11558,N_9323,N_10027);
nor U11559 (N_11559,N_9549,N_9450);
or U11560 (N_11560,N_9575,N_9708);
xor U11561 (N_11561,N_10123,N_9517);
and U11562 (N_11562,N_9407,N_10396);
or U11563 (N_11563,N_9137,N_10410);
nor U11564 (N_11564,N_10015,N_9370);
nor U11565 (N_11565,N_10098,N_10454);
or U11566 (N_11566,N_9883,N_9125);
nand U11567 (N_11567,N_10363,N_9439);
and U11568 (N_11568,N_9359,N_10057);
or U11569 (N_11569,N_9399,N_9854);
nand U11570 (N_11570,N_9293,N_9817);
and U11571 (N_11571,N_9004,N_9532);
and U11572 (N_11572,N_9066,N_9822);
and U11573 (N_11573,N_9741,N_10318);
and U11574 (N_11574,N_9142,N_9939);
and U11575 (N_11575,N_9485,N_10052);
and U11576 (N_11576,N_9833,N_9954);
and U11577 (N_11577,N_9051,N_9031);
and U11578 (N_11578,N_9996,N_9713);
nor U11579 (N_11579,N_10003,N_9003);
nor U11580 (N_11580,N_10152,N_10459);
or U11581 (N_11581,N_9587,N_9943);
nand U11582 (N_11582,N_10488,N_9233);
or U11583 (N_11583,N_9514,N_9914);
or U11584 (N_11584,N_10173,N_9709);
nor U11585 (N_11585,N_10458,N_9676);
xnor U11586 (N_11586,N_10255,N_9794);
nor U11587 (N_11587,N_9354,N_9277);
and U11588 (N_11588,N_10209,N_10432);
or U11589 (N_11589,N_9483,N_9452);
and U11590 (N_11590,N_9329,N_10342);
and U11591 (N_11591,N_9095,N_10482);
xnor U11592 (N_11592,N_10313,N_10111);
or U11593 (N_11593,N_10424,N_9614);
or U11594 (N_11594,N_10489,N_9888);
and U11595 (N_11595,N_9836,N_9967);
xor U11596 (N_11596,N_9262,N_10358);
nand U11597 (N_11597,N_10420,N_9460);
xor U11598 (N_11598,N_10223,N_10342);
nor U11599 (N_11599,N_9302,N_9726);
and U11600 (N_11600,N_9103,N_9708);
and U11601 (N_11601,N_10340,N_10115);
nand U11602 (N_11602,N_9360,N_9411);
nor U11603 (N_11603,N_9102,N_9392);
xor U11604 (N_11604,N_9297,N_9502);
nand U11605 (N_11605,N_9545,N_9807);
or U11606 (N_11606,N_9530,N_10251);
and U11607 (N_11607,N_9392,N_9446);
nand U11608 (N_11608,N_10283,N_10423);
and U11609 (N_11609,N_10338,N_9601);
or U11610 (N_11610,N_9763,N_9508);
or U11611 (N_11611,N_9891,N_9746);
or U11612 (N_11612,N_9327,N_10002);
nor U11613 (N_11613,N_9278,N_9051);
nor U11614 (N_11614,N_9977,N_9300);
or U11615 (N_11615,N_9282,N_10136);
or U11616 (N_11616,N_9723,N_10233);
and U11617 (N_11617,N_9430,N_9775);
or U11618 (N_11618,N_10462,N_9655);
nor U11619 (N_11619,N_9179,N_9664);
nand U11620 (N_11620,N_9837,N_10411);
or U11621 (N_11621,N_10295,N_9958);
and U11622 (N_11622,N_9663,N_9125);
nor U11623 (N_11623,N_10118,N_10007);
nor U11624 (N_11624,N_9255,N_10166);
xnor U11625 (N_11625,N_9353,N_10389);
nand U11626 (N_11626,N_10344,N_10053);
nor U11627 (N_11627,N_9246,N_10290);
or U11628 (N_11628,N_9230,N_9107);
nor U11629 (N_11629,N_10463,N_9582);
nand U11630 (N_11630,N_10405,N_9911);
nor U11631 (N_11631,N_9283,N_9064);
nand U11632 (N_11632,N_9958,N_10142);
nand U11633 (N_11633,N_10216,N_9459);
nand U11634 (N_11634,N_10354,N_10289);
and U11635 (N_11635,N_9329,N_9042);
or U11636 (N_11636,N_9569,N_9086);
nor U11637 (N_11637,N_9773,N_9895);
and U11638 (N_11638,N_9639,N_9748);
and U11639 (N_11639,N_10129,N_9368);
nor U11640 (N_11640,N_9598,N_10091);
and U11641 (N_11641,N_9204,N_9614);
and U11642 (N_11642,N_9869,N_9292);
or U11643 (N_11643,N_9294,N_9662);
nor U11644 (N_11644,N_10000,N_9818);
nor U11645 (N_11645,N_9009,N_9966);
xor U11646 (N_11646,N_9140,N_10421);
nand U11647 (N_11647,N_9575,N_9046);
nor U11648 (N_11648,N_10402,N_10375);
and U11649 (N_11649,N_9276,N_10299);
or U11650 (N_11650,N_9794,N_10212);
nand U11651 (N_11651,N_9183,N_9364);
and U11652 (N_11652,N_10237,N_10289);
or U11653 (N_11653,N_10166,N_10174);
nor U11654 (N_11654,N_9522,N_10379);
nand U11655 (N_11655,N_9818,N_10396);
or U11656 (N_11656,N_9492,N_9476);
and U11657 (N_11657,N_9234,N_9925);
or U11658 (N_11658,N_9908,N_9451);
or U11659 (N_11659,N_10472,N_9434);
or U11660 (N_11660,N_9557,N_9921);
or U11661 (N_11661,N_9191,N_10360);
xor U11662 (N_11662,N_9339,N_9948);
or U11663 (N_11663,N_9246,N_9932);
nor U11664 (N_11664,N_9746,N_9892);
and U11665 (N_11665,N_10374,N_9232);
and U11666 (N_11666,N_9620,N_10472);
xnor U11667 (N_11667,N_9579,N_10190);
or U11668 (N_11668,N_9727,N_9171);
nand U11669 (N_11669,N_9572,N_9939);
nor U11670 (N_11670,N_9804,N_10083);
nor U11671 (N_11671,N_10231,N_9900);
xnor U11672 (N_11672,N_10112,N_9332);
and U11673 (N_11673,N_10258,N_9199);
nor U11674 (N_11674,N_9948,N_9572);
nor U11675 (N_11675,N_9818,N_9107);
or U11676 (N_11676,N_9252,N_9941);
nor U11677 (N_11677,N_9034,N_9448);
or U11678 (N_11678,N_10177,N_10264);
xor U11679 (N_11679,N_9953,N_9249);
nand U11680 (N_11680,N_10322,N_10333);
nand U11681 (N_11681,N_9234,N_10341);
nand U11682 (N_11682,N_9914,N_10212);
nor U11683 (N_11683,N_9577,N_10497);
and U11684 (N_11684,N_9857,N_9126);
nor U11685 (N_11685,N_9051,N_10469);
xnor U11686 (N_11686,N_9468,N_9863);
and U11687 (N_11687,N_9833,N_9140);
nand U11688 (N_11688,N_10093,N_9703);
and U11689 (N_11689,N_10203,N_9902);
and U11690 (N_11690,N_9075,N_9372);
xor U11691 (N_11691,N_10140,N_10486);
nand U11692 (N_11692,N_9984,N_9460);
nand U11693 (N_11693,N_10305,N_9046);
or U11694 (N_11694,N_9350,N_9338);
nor U11695 (N_11695,N_9774,N_9622);
nand U11696 (N_11696,N_9423,N_9064);
nor U11697 (N_11697,N_9707,N_9086);
or U11698 (N_11698,N_9215,N_9777);
or U11699 (N_11699,N_9211,N_9274);
and U11700 (N_11700,N_9692,N_9473);
and U11701 (N_11701,N_9580,N_9292);
nand U11702 (N_11702,N_10261,N_9774);
nor U11703 (N_11703,N_9508,N_9945);
nor U11704 (N_11704,N_10464,N_10480);
nand U11705 (N_11705,N_9044,N_9454);
or U11706 (N_11706,N_9324,N_10045);
nand U11707 (N_11707,N_9399,N_9323);
nor U11708 (N_11708,N_10318,N_9538);
nand U11709 (N_11709,N_10470,N_9854);
nand U11710 (N_11710,N_9615,N_9788);
nand U11711 (N_11711,N_9968,N_9850);
or U11712 (N_11712,N_9260,N_10425);
and U11713 (N_11713,N_10100,N_9601);
nand U11714 (N_11714,N_10490,N_10214);
and U11715 (N_11715,N_10326,N_9610);
and U11716 (N_11716,N_9250,N_9645);
nand U11717 (N_11717,N_10355,N_10480);
and U11718 (N_11718,N_9010,N_9161);
nand U11719 (N_11719,N_10242,N_10160);
nand U11720 (N_11720,N_10385,N_9127);
and U11721 (N_11721,N_10246,N_9462);
nand U11722 (N_11722,N_9762,N_9289);
and U11723 (N_11723,N_9266,N_9306);
nand U11724 (N_11724,N_9792,N_10411);
or U11725 (N_11725,N_9760,N_9484);
xor U11726 (N_11726,N_9388,N_9421);
and U11727 (N_11727,N_9261,N_9280);
or U11728 (N_11728,N_10359,N_9488);
nand U11729 (N_11729,N_9317,N_10384);
nor U11730 (N_11730,N_10363,N_10337);
and U11731 (N_11731,N_9903,N_9917);
xnor U11732 (N_11732,N_9952,N_9046);
nand U11733 (N_11733,N_9879,N_9046);
or U11734 (N_11734,N_10069,N_10378);
or U11735 (N_11735,N_9733,N_9384);
xnor U11736 (N_11736,N_10218,N_10191);
nand U11737 (N_11737,N_9213,N_9523);
nor U11738 (N_11738,N_10115,N_9170);
or U11739 (N_11739,N_10411,N_9662);
or U11740 (N_11740,N_10091,N_10436);
nand U11741 (N_11741,N_9647,N_9877);
or U11742 (N_11742,N_9099,N_9319);
nand U11743 (N_11743,N_9828,N_10217);
or U11744 (N_11744,N_9538,N_9699);
nor U11745 (N_11745,N_9341,N_9702);
or U11746 (N_11746,N_9223,N_9626);
nand U11747 (N_11747,N_10307,N_9939);
or U11748 (N_11748,N_9076,N_10198);
nor U11749 (N_11749,N_10431,N_10124);
nor U11750 (N_11750,N_10133,N_10100);
or U11751 (N_11751,N_9015,N_10031);
nor U11752 (N_11752,N_9393,N_9475);
and U11753 (N_11753,N_9188,N_10037);
xor U11754 (N_11754,N_10183,N_9484);
or U11755 (N_11755,N_9942,N_9268);
nand U11756 (N_11756,N_10132,N_9249);
xor U11757 (N_11757,N_9784,N_9581);
and U11758 (N_11758,N_9995,N_10052);
or U11759 (N_11759,N_10033,N_10190);
nand U11760 (N_11760,N_9057,N_9532);
or U11761 (N_11761,N_10031,N_10300);
nand U11762 (N_11762,N_9878,N_9816);
or U11763 (N_11763,N_9748,N_10467);
nor U11764 (N_11764,N_10455,N_10499);
or U11765 (N_11765,N_10108,N_9845);
nand U11766 (N_11766,N_10388,N_10042);
nand U11767 (N_11767,N_9889,N_10312);
nor U11768 (N_11768,N_9273,N_9228);
and U11769 (N_11769,N_10132,N_9435);
xor U11770 (N_11770,N_9411,N_9609);
or U11771 (N_11771,N_9640,N_10046);
nor U11772 (N_11772,N_10474,N_9835);
or U11773 (N_11773,N_9669,N_9181);
and U11774 (N_11774,N_9271,N_10416);
and U11775 (N_11775,N_9957,N_9043);
xnor U11776 (N_11776,N_9382,N_9367);
nor U11777 (N_11777,N_9121,N_10147);
nor U11778 (N_11778,N_9595,N_10402);
nor U11779 (N_11779,N_9099,N_9357);
or U11780 (N_11780,N_9834,N_9737);
xnor U11781 (N_11781,N_9582,N_9780);
nand U11782 (N_11782,N_9574,N_10165);
or U11783 (N_11783,N_9193,N_10407);
or U11784 (N_11784,N_9496,N_9771);
and U11785 (N_11785,N_10241,N_9693);
or U11786 (N_11786,N_9329,N_9774);
nand U11787 (N_11787,N_9708,N_10112);
nor U11788 (N_11788,N_10308,N_9620);
nor U11789 (N_11789,N_9000,N_9303);
xnor U11790 (N_11790,N_9039,N_10273);
or U11791 (N_11791,N_9244,N_9252);
or U11792 (N_11792,N_9271,N_10118);
nor U11793 (N_11793,N_9350,N_10494);
nand U11794 (N_11794,N_10180,N_9339);
nor U11795 (N_11795,N_10347,N_10012);
nand U11796 (N_11796,N_9138,N_10193);
or U11797 (N_11797,N_9783,N_9625);
and U11798 (N_11798,N_9040,N_9791);
nand U11799 (N_11799,N_9396,N_9419);
xnor U11800 (N_11800,N_10390,N_9666);
and U11801 (N_11801,N_10092,N_10148);
xor U11802 (N_11802,N_10040,N_10297);
or U11803 (N_11803,N_9668,N_10481);
nand U11804 (N_11804,N_9058,N_9109);
nor U11805 (N_11805,N_9414,N_9901);
or U11806 (N_11806,N_10006,N_9559);
or U11807 (N_11807,N_9012,N_9660);
xnor U11808 (N_11808,N_10282,N_9329);
nand U11809 (N_11809,N_9701,N_10351);
nor U11810 (N_11810,N_9222,N_10184);
and U11811 (N_11811,N_9180,N_9525);
or U11812 (N_11812,N_10125,N_9723);
xor U11813 (N_11813,N_9350,N_9383);
xnor U11814 (N_11814,N_9153,N_10401);
xnor U11815 (N_11815,N_9816,N_9530);
nor U11816 (N_11816,N_9874,N_9172);
nor U11817 (N_11817,N_9007,N_9880);
or U11818 (N_11818,N_10137,N_9733);
or U11819 (N_11819,N_9121,N_9036);
or U11820 (N_11820,N_10072,N_10428);
nand U11821 (N_11821,N_9619,N_9600);
or U11822 (N_11822,N_10034,N_9600);
nand U11823 (N_11823,N_9828,N_9905);
nor U11824 (N_11824,N_10070,N_9097);
nor U11825 (N_11825,N_9094,N_9748);
nand U11826 (N_11826,N_9046,N_9740);
and U11827 (N_11827,N_9334,N_9944);
nand U11828 (N_11828,N_10068,N_9533);
nand U11829 (N_11829,N_9291,N_9171);
nor U11830 (N_11830,N_9473,N_9733);
or U11831 (N_11831,N_9420,N_9417);
xnor U11832 (N_11832,N_9704,N_10137);
and U11833 (N_11833,N_9529,N_10070);
and U11834 (N_11834,N_9644,N_10254);
nand U11835 (N_11835,N_10451,N_10079);
nand U11836 (N_11836,N_9568,N_9771);
xnor U11837 (N_11837,N_10281,N_9909);
nor U11838 (N_11838,N_10477,N_10081);
and U11839 (N_11839,N_9251,N_9672);
and U11840 (N_11840,N_10360,N_9421);
and U11841 (N_11841,N_9724,N_9337);
or U11842 (N_11842,N_9727,N_9434);
nand U11843 (N_11843,N_9579,N_9493);
and U11844 (N_11844,N_9448,N_10001);
nand U11845 (N_11845,N_9429,N_10260);
or U11846 (N_11846,N_9076,N_9658);
nand U11847 (N_11847,N_10208,N_9802);
or U11848 (N_11848,N_9465,N_9768);
nor U11849 (N_11849,N_9390,N_9616);
xor U11850 (N_11850,N_9404,N_9814);
nand U11851 (N_11851,N_9908,N_9383);
xor U11852 (N_11852,N_9484,N_10467);
nand U11853 (N_11853,N_9668,N_9817);
nand U11854 (N_11854,N_10197,N_10303);
xnor U11855 (N_11855,N_10076,N_9833);
nor U11856 (N_11856,N_9139,N_9848);
or U11857 (N_11857,N_9897,N_9845);
and U11858 (N_11858,N_10118,N_10013);
nand U11859 (N_11859,N_9835,N_10467);
or U11860 (N_11860,N_9900,N_10180);
xor U11861 (N_11861,N_9567,N_10005);
nand U11862 (N_11862,N_9939,N_9426);
or U11863 (N_11863,N_9097,N_9496);
nor U11864 (N_11864,N_9955,N_9572);
or U11865 (N_11865,N_9546,N_9579);
xor U11866 (N_11866,N_9183,N_10370);
xor U11867 (N_11867,N_9099,N_10183);
xor U11868 (N_11868,N_9021,N_9277);
and U11869 (N_11869,N_10286,N_10050);
nand U11870 (N_11870,N_9760,N_9990);
or U11871 (N_11871,N_9592,N_9128);
nand U11872 (N_11872,N_9620,N_10352);
xor U11873 (N_11873,N_10296,N_9040);
xnor U11874 (N_11874,N_9816,N_9188);
nor U11875 (N_11875,N_10375,N_9239);
nand U11876 (N_11876,N_10284,N_10433);
nor U11877 (N_11877,N_9447,N_9462);
nor U11878 (N_11878,N_9923,N_10066);
nor U11879 (N_11879,N_9895,N_10297);
and U11880 (N_11880,N_9103,N_9044);
nor U11881 (N_11881,N_10082,N_10013);
xnor U11882 (N_11882,N_9450,N_10375);
nor U11883 (N_11883,N_10258,N_10481);
nor U11884 (N_11884,N_9300,N_10374);
nor U11885 (N_11885,N_9846,N_9254);
nor U11886 (N_11886,N_9769,N_9972);
or U11887 (N_11887,N_9945,N_9565);
or U11888 (N_11888,N_9794,N_9985);
or U11889 (N_11889,N_10459,N_9239);
or U11890 (N_11890,N_9172,N_9480);
nand U11891 (N_11891,N_9794,N_9703);
nor U11892 (N_11892,N_9322,N_10455);
nor U11893 (N_11893,N_9942,N_10363);
nand U11894 (N_11894,N_9385,N_10142);
or U11895 (N_11895,N_9901,N_9214);
nor U11896 (N_11896,N_10113,N_9197);
nor U11897 (N_11897,N_9418,N_9581);
nand U11898 (N_11898,N_9324,N_9961);
or U11899 (N_11899,N_9302,N_9328);
or U11900 (N_11900,N_9285,N_9408);
xnor U11901 (N_11901,N_10079,N_9412);
xnor U11902 (N_11902,N_9339,N_9120);
or U11903 (N_11903,N_9857,N_9584);
or U11904 (N_11904,N_10198,N_9655);
nor U11905 (N_11905,N_9637,N_10444);
nand U11906 (N_11906,N_9731,N_10392);
nand U11907 (N_11907,N_9623,N_9297);
or U11908 (N_11908,N_9141,N_10433);
nor U11909 (N_11909,N_9591,N_10337);
or U11910 (N_11910,N_10353,N_9843);
and U11911 (N_11911,N_9784,N_9344);
xor U11912 (N_11912,N_10211,N_10296);
nand U11913 (N_11913,N_10023,N_9465);
nand U11914 (N_11914,N_10193,N_9176);
nand U11915 (N_11915,N_9409,N_9642);
or U11916 (N_11916,N_10485,N_9528);
and U11917 (N_11917,N_10388,N_10231);
and U11918 (N_11918,N_9891,N_9025);
nand U11919 (N_11919,N_10108,N_9748);
nor U11920 (N_11920,N_10037,N_9017);
nand U11921 (N_11921,N_10034,N_9094);
or U11922 (N_11922,N_10232,N_9428);
nand U11923 (N_11923,N_10083,N_9383);
nand U11924 (N_11924,N_9981,N_9786);
nor U11925 (N_11925,N_10014,N_9358);
nand U11926 (N_11926,N_10117,N_10136);
nor U11927 (N_11927,N_9496,N_10320);
nand U11928 (N_11928,N_9020,N_9050);
and U11929 (N_11929,N_10271,N_9481);
nor U11930 (N_11930,N_9351,N_9783);
and U11931 (N_11931,N_9887,N_9733);
nand U11932 (N_11932,N_9255,N_9028);
or U11933 (N_11933,N_10354,N_10004);
and U11934 (N_11934,N_9545,N_9654);
nor U11935 (N_11935,N_9301,N_10293);
nor U11936 (N_11936,N_10172,N_9523);
nor U11937 (N_11937,N_9071,N_9391);
and U11938 (N_11938,N_10084,N_10039);
nor U11939 (N_11939,N_9272,N_10159);
or U11940 (N_11940,N_9727,N_9910);
and U11941 (N_11941,N_9323,N_10093);
nand U11942 (N_11942,N_10376,N_10319);
xor U11943 (N_11943,N_10252,N_9927);
or U11944 (N_11944,N_9150,N_9039);
nand U11945 (N_11945,N_9801,N_9308);
nor U11946 (N_11946,N_10023,N_9236);
nor U11947 (N_11947,N_9254,N_9653);
or U11948 (N_11948,N_9913,N_10424);
nor U11949 (N_11949,N_9476,N_9232);
or U11950 (N_11950,N_9054,N_9081);
or U11951 (N_11951,N_9227,N_10486);
nand U11952 (N_11952,N_9998,N_10184);
nand U11953 (N_11953,N_9019,N_9675);
xor U11954 (N_11954,N_10323,N_10129);
xor U11955 (N_11955,N_9163,N_9676);
nand U11956 (N_11956,N_9170,N_9881);
or U11957 (N_11957,N_9224,N_9221);
nand U11958 (N_11958,N_9055,N_10384);
and U11959 (N_11959,N_9081,N_10340);
nand U11960 (N_11960,N_9514,N_10117);
xor U11961 (N_11961,N_9133,N_10094);
xor U11962 (N_11962,N_10264,N_9294);
or U11963 (N_11963,N_10294,N_10277);
nor U11964 (N_11964,N_9842,N_9869);
nor U11965 (N_11965,N_9991,N_9997);
or U11966 (N_11966,N_10100,N_9715);
nor U11967 (N_11967,N_9149,N_9543);
xor U11968 (N_11968,N_9223,N_10094);
and U11969 (N_11969,N_9762,N_9870);
nor U11970 (N_11970,N_9148,N_9039);
or U11971 (N_11971,N_10279,N_9045);
nand U11972 (N_11972,N_9837,N_10104);
nand U11973 (N_11973,N_10357,N_9966);
nor U11974 (N_11974,N_9491,N_9388);
xnor U11975 (N_11975,N_10002,N_9740);
nand U11976 (N_11976,N_10372,N_10479);
or U11977 (N_11977,N_10147,N_9198);
nand U11978 (N_11978,N_9284,N_9288);
or U11979 (N_11979,N_9220,N_9547);
or U11980 (N_11980,N_10074,N_9656);
xor U11981 (N_11981,N_9639,N_10276);
or U11982 (N_11982,N_9300,N_9421);
nor U11983 (N_11983,N_9992,N_10434);
nor U11984 (N_11984,N_9386,N_9275);
nand U11985 (N_11985,N_9945,N_9119);
or U11986 (N_11986,N_9834,N_9129);
nor U11987 (N_11987,N_9464,N_9918);
and U11988 (N_11988,N_10496,N_9066);
nand U11989 (N_11989,N_9136,N_9706);
or U11990 (N_11990,N_9038,N_10175);
and U11991 (N_11991,N_9634,N_10210);
nor U11992 (N_11992,N_9368,N_10404);
nor U11993 (N_11993,N_9829,N_9047);
and U11994 (N_11994,N_9045,N_9206);
and U11995 (N_11995,N_9504,N_9304);
or U11996 (N_11996,N_9544,N_10350);
nand U11997 (N_11997,N_10376,N_9630);
nand U11998 (N_11998,N_10376,N_10457);
nand U11999 (N_11999,N_9769,N_10465);
nor U12000 (N_12000,N_11943,N_11301);
and U12001 (N_12001,N_11510,N_10814);
and U12002 (N_12002,N_10753,N_11090);
xnor U12003 (N_12003,N_10661,N_11092);
nand U12004 (N_12004,N_10938,N_10971);
nor U12005 (N_12005,N_11010,N_10839);
nor U12006 (N_12006,N_10685,N_11720);
or U12007 (N_12007,N_10723,N_11332);
and U12008 (N_12008,N_10763,N_11341);
or U12009 (N_12009,N_11956,N_11819);
xor U12010 (N_12010,N_11232,N_10698);
and U12011 (N_12011,N_11096,N_11048);
nand U12012 (N_12012,N_11363,N_11877);
nor U12013 (N_12013,N_10801,N_11480);
nor U12014 (N_12014,N_10773,N_11704);
nand U12015 (N_12015,N_11831,N_11841);
nand U12016 (N_12016,N_11388,N_10770);
or U12017 (N_12017,N_11974,N_11658);
nand U12018 (N_12018,N_11492,N_11037);
nor U12019 (N_12019,N_10933,N_10541);
xor U12020 (N_12020,N_11427,N_10691);
xor U12021 (N_12021,N_11271,N_10833);
nor U12022 (N_12022,N_11715,N_11752);
and U12023 (N_12023,N_10767,N_11270);
and U12024 (N_12024,N_10690,N_10975);
xor U12025 (N_12025,N_11791,N_11944);
or U12026 (N_12026,N_10624,N_10582);
or U12027 (N_12027,N_10623,N_11891);
nand U12028 (N_12028,N_10654,N_10913);
and U12029 (N_12029,N_11884,N_10512);
nor U12030 (N_12030,N_10641,N_10703);
or U12031 (N_12031,N_10995,N_11909);
and U12032 (N_12032,N_11825,N_10630);
nor U12033 (N_12033,N_11848,N_11539);
or U12034 (N_12034,N_10579,N_11274);
nand U12035 (N_12035,N_10779,N_11112);
nor U12036 (N_12036,N_11662,N_11766);
nand U12037 (N_12037,N_11700,N_10550);
or U12038 (N_12038,N_11229,N_11666);
nor U12039 (N_12039,N_11078,N_11685);
nand U12040 (N_12040,N_11686,N_10872);
nor U12041 (N_12041,N_10710,N_11143);
nor U12042 (N_12042,N_11763,N_10859);
xor U12043 (N_12043,N_10775,N_11678);
nand U12044 (N_12044,N_11774,N_11489);
nor U12045 (N_12045,N_11642,N_11648);
xor U12046 (N_12046,N_11923,N_11703);
nor U12047 (N_12047,N_11213,N_11546);
nor U12048 (N_12048,N_11101,N_11870);
nand U12049 (N_12049,N_10789,N_10882);
xnor U12050 (N_12050,N_11983,N_11952);
nor U12051 (N_12051,N_11395,N_10840);
and U12052 (N_12052,N_11150,N_11739);
or U12053 (N_12053,N_11850,N_11479);
and U12054 (N_12054,N_10970,N_11838);
and U12055 (N_12055,N_10846,N_11279);
nor U12056 (N_12056,N_11194,N_11504);
or U12057 (N_12057,N_11623,N_10953);
nor U12058 (N_12058,N_11136,N_11840);
xnor U12059 (N_12059,N_11018,N_11424);
xor U12060 (N_12060,N_10988,N_11097);
and U12061 (N_12061,N_10602,N_11033);
or U12062 (N_12062,N_11968,N_11562);
nand U12063 (N_12063,N_11311,N_11744);
nor U12064 (N_12064,N_11303,N_11688);
nand U12065 (N_12065,N_10904,N_11231);
and U12066 (N_12066,N_11401,N_11799);
or U12067 (N_12067,N_11809,N_10722);
nand U12068 (N_12068,N_11812,N_11133);
nor U12069 (N_12069,N_10824,N_11059);
nor U12070 (N_12070,N_11695,N_11066);
nor U12071 (N_12071,N_10919,N_11663);
nand U12072 (N_12072,N_10662,N_10860);
nand U12073 (N_12073,N_10927,N_10709);
xnor U12074 (N_12074,N_11595,N_11660);
or U12075 (N_12075,N_11652,N_11501);
nand U12076 (N_12076,N_11972,N_11040);
and U12077 (N_12077,N_11965,N_11371);
nand U12078 (N_12078,N_10660,N_11731);
nand U12079 (N_12079,N_11076,N_11200);
or U12080 (N_12080,N_11467,N_11938);
or U12081 (N_12081,N_10517,N_10883);
xnor U12082 (N_12082,N_11331,N_11743);
and U12083 (N_12083,N_11179,N_11935);
nand U12084 (N_12084,N_11151,N_11188);
nor U12085 (N_12085,N_10819,N_10858);
nand U12086 (N_12086,N_11728,N_11434);
or U12087 (N_12087,N_10593,N_11975);
nand U12088 (N_12088,N_11951,N_10750);
or U12089 (N_12089,N_11497,N_10877);
nor U12090 (N_12090,N_11665,N_11697);
nand U12091 (N_12091,N_10989,N_11071);
nand U12092 (N_12092,N_11042,N_10893);
and U12093 (N_12093,N_11505,N_11741);
or U12094 (N_12094,N_10791,N_11913);
nor U12095 (N_12095,N_11586,N_11485);
or U12096 (N_12096,N_11158,N_11596);
xnor U12097 (N_12097,N_11340,N_11214);
or U12098 (N_12098,N_11468,N_11988);
xnor U12099 (N_12099,N_10962,N_10817);
nor U12100 (N_12100,N_11383,N_11577);
and U12101 (N_12101,N_11190,N_11751);
nor U12102 (N_12102,N_10577,N_10911);
and U12103 (N_12103,N_11220,N_11611);
nand U12104 (N_12104,N_11465,N_11374);
nand U12105 (N_12105,N_11954,N_11835);
or U12106 (N_12106,N_11769,N_11615);
or U12107 (N_12107,N_10669,N_11297);
or U12108 (N_12108,N_11117,N_10968);
nor U12109 (N_12109,N_11287,N_11285);
and U12110 (N_12110,N_10831,N_10559);
nor U12111 (N_12111,N_10925,N_11152);
or U12112 (N_12112,N_11367,N_10769);
nor U12113 (N_12113,N_11613,N_11277);
nor U12114 (N_12114,N_11472,N_11453);
nor U12115 (N_12115,N_10874,N_11708);
or U12116 (N_12116,N_10665,N_10578);
nor U12117 (N_12117,N_11722,N_10887);
nand U12118 (N_12118,N_10842,N_10596);
nand U12119 (N_12119,N_10552,N_11959);
or U12120 (N_12120,N_10570,N_11630);
and U12121 (N_12121,N_10542,N_11603);
xor U12122 (N_12122,N_11607,N_11717);
or U12123 (N_12123,N_10803,N_11425);
nor U12124 (N_12124,N_11254,N_10657);
and U12125 (N_12125,N_10896,N_10562);
nand U12126 (N_12126,N_11113,N_11627);
or U12127 (N_12127,N_10617,N_10906);
or U12128 (N_12128,N_11661,N_10986);
nor U12129 (N_12129,N_11500,N_11691);
nor U12130 (N_12130,N_11049,N_11647);
and U12131 (N_12131,N_10847,N_10683);
and U12132 (N_12132,N_10798,N_11865);
and U12133 (N_12133,N_10591,N_11084);
nand U12134 (N_12134,N_11571,N_10594);
and U12135 (N_12135,N_11324,N_11091);
or U12136 (N_12136,N_11377,N_11813);
nor U12137 (N_12137,N_11366,N_11197);
and U12138 (N_12138,N_11327,N_11714);
or U12139 (N_12139,N_11372,N_11278);
nor U12140 (N_12140,N_11748,N_11183);
nor U12141 (N_12141,N_11261,N_11885);
and U12142 (N_12142,N_11706,N_10734);
and U12143 (N_12143,N_11716,N_10565);
nor U12144 (N_12144,N_11430,N_10568);
and U12145 (N_12145,N_11138,N_11206);
nor U12146 (N_12146,N_11140,N_11128);
or U12147 (N_12147,N_11517,N_11106);
nand U12148 (N_12148,N_11435,N_11369);
nor U12149 (N_12149,N_11193,N_10950);
nand U12150 (N_12150,N_11432,N_11458);
and U12151 (N_12151,N_10885,N_10576);
nand U12152 (N_12152,N_10609,N_10870);
nand U12153 (N_12153,N_10606,N_11633);
or U12154 (N_12154,N_11142,N_10735);
and U12155 (N_12155,N_11878,N_10748);
nor U12156 (N_12156,N_10828,N_10561);
or U12157 (N_12157,N_11013,N_11629);
nor U12158 (N_12158,N_11225,N_11549);
nand U12159 (N_12159,N_11767,N_11275);
xor U12160 (N_12160,N_11223,N_10957);
nand U12161 (N_12161,N_10668,N_11309);
nor U12162 (N_12162,N_11664,N_11019);
nand U12163 (N_12163,N_11826,N_11025);
nand U12164 (N_12164,N_11569,N_11792);
xor U12165 (N_12165,N_11325,N_11990);
and U12166 (N_12166,N_11062,N_11413);
and U12167 (N_12167,N_11955,N_10777);
nor U12168 (N_12168,N_10905,N_10838);
xor U12169 (N_12169,N_10615,N_11568);
or U12170 (N_12170,N_10652,N_11359);
nor U12171 (N_12171,N_11796,N_10604);
xnor U12172 (N_12172,N_11585,N_10644);
nor U12173 (N_12173,N_11855,N_10642);
and U12174 (N_12174,N_11534,N_11864);
and U12175 (N_12175,N_11289,N_10535);
or U12176 (N_12176,N_11355,N_10943);
and U12177 (N_12177,N_11007,N_10857);
nand U12178 (N_12178,N_11851,N_10781);
nand U12179 (N_12179,N_11281,N_10731);
or U12180 (N_12180,N_10677,N_10929);
nand U12181 (N_12181,N_11445,N_11072);
or U12182 (N_12182,N_10848,N_11541);
nand U12183 (N_12183,N_11027,N_11391);
nor U12184 (N_12184,N_11230,N_11807);
and U12185 (N_12185,N_11455,N_11318);
and U12186 (N_12186,N_11985,N_11109);
or U12187 (N_12187,N_11482,N_11003);
or U12188 (N_12188,N_10634,N_11879);
or U12189 (N_12189,N_10794,N_11755);
nand U12190 (N_12190,N_11645,N_11429);
or U12191 (N_12191,N_11949,N_10705);
nand U12192 (N_12192,N_11637,N_11542);
xnor U12193 (N_12193,N_11119,N_11221);
nor U12194 (N_12194,N_11578,N_10761);
nand U12195 (N_12195,N_11973,N_10500);
nand U12196 (N_12196,N_11387,N_10524);
nor U12197 (N_12197,N_11868,N_11093);
nand U12198 (N_12198,N_11046,N_11937);
and U12199 (N_12199,N_11902,N_11525);
and U12200 (N_12200,N_11522,N_10707);
and U12201 (N_12201,N_11824,N_10759);
and U12202 (N_12202,N_11265,N_10649);
and U12203 (N_12203,N_11683,N_11020);
or U12204 (N_12204,N_11762,N_11654);
and U12205 (N_12205,N_10765,N_10627);
nor U12206 (N_12206,N_11358,N_10718);
or U12207 (N_12207,N_11996,N_11872);
or U12208 (N_12208,N_11618,N_11583);
or U12209 (N_12209,N_11460,N_11834);
and U12210 (N_12210,N_11643,N_11993);
or U12211 (N_12211,N_10937,N_11380);
xor U12212 (N_12212,N_10888,N_11895);
or U12213 (N_12213,N_11156,N_11908);
and U12214 (N_12214,N_11313,N_11530);
nor U12215 (N_12215,N_11047,N_11635);
or U12216 (N_12216,N_11998,N_10534);
or U12217 (N_12217,N_10967,N_11357);
xnor U12218 (N_12218,N_11181,N_11061);
nor U12219 (N_12219,N_10928,N_11684);
and U12220 (N_12220,N_11528,N_11853);
or U12221 (N_12221,N_10704,N_10567);
or U12222 (N_12222,N_11565,N_11982);
nor U12223 (N_12223,N_11070,N_11857);
nor U12224 (N_12224,N_10978,N_11368);
and U12225 (N_12225,N_11103,N_11911);
and U12226 (N_12226,N_10912,N_10645);
or U12227 (N_12227,N_10864,N_11130);
nor U12228 (N_12228,N_11619,N_11822);
or U12229 (N_12229,N_11417,N_11000);
or U12230 (N_12230,N_11723,N_10613);
nor U12231 (N_12231,N_11713,N_11579);
nand U12232 (N_12232,N_11828,N_10800);
or U12233 (N_12233,N_11334,N_11994);
and U12234 (N_12234,N_10876,N_11378);
and U12235 (N_12235,N_11349,N_11167);
nand U12236 (N_12236,N_10643,N_11947);
nor U12237 (N_12237,N_10572,N_11719);
nor U12238 (N_12238,N_11861,N_11449);
xor U12239 (N_12239,N_11195,N_11679);
and U12240 (N_12240,N_11800,N_10708);
xnor U12241 (N_12241,N_10889,N_10740);
xor U12242 (N_12242,N_11298,N_11111);
and U12243 (N_12243,N_11342,N_11602);
and U12244 (N_12244,N_11921,N_11893);
xor U12245 (N_12245,N_11085,N_11116);
nand U12246 (N_12246,N_11137,N_11593);
or U12247 (N_12247,N_11147,N_11503);
xnor U12248 (N_12248,N_11210,N_10597);
or U12249 (N_12249,N_11862,N_11980);
or U12250 (N_12250,N_11051,N_11651);
nand U12251 (N_12251,N_11330,N_10523);
nor U12252 (N_12252,N_10880,N_11842);
nor U12253 (N_12253,N_11749,N_11088);
and U12254 (N_12254,N_11304,N_10994);
and U12255 (N_12255,N_10891,N_11962);
xnor U12256 (N_12256,N_11738,N_11346);
and U12257 (N_12257,N_11361,N_11474);
nor U12258 (N_12258,N_10536,N_10670);
and U12259 (N_12259,N_10745,N_11022);
and U12260 (N_12260,N_11428,N_11919);
nor U12261 (N_12261,N_10659,N_11004);
nor U12262 (N_12262,N_11375,N_11702);
nand U12263 (N_12263,N_10974,N_11617);
xnor U12264 (N_12264,N_11162,N_11918);
or U12265 (N_12265,N_11668,N_11405);
nor U12266 (N_12266,N_11439,N_11269);
or U12267 (N_12267,N_11782,N_11258);
nor U12268 (N_12268,N_10672,N_10598);
and U12269 (N_12269,N_11543,N_10861);
or U12270 (N_12270,N_10895,N_10780);
and U12271 (N_12271,N_10530,N_10622);
nor U12272 (N_12272,N_10966,N_11552);
and U12273 (N_12273,N_10618,N_10676);
nor U12274 (N_12274,N_11291,N_11450);
and U12275 (N_12275,N_10981,N_10571);
nand U12276 (N_12276,N_10539,N_10818);
or U12277 (N_12277,N_11053,N_10737);
nor U12278 (N_12278,N_10506,N_10656);
xor U12279 (N_12279,N_11146,N_11100);
and U12280 (N_12280,N_11174,N_10648);
nor U12281 (N_12281,N_11575,N_11524);
or U12282 (N_12282,N_11581,N_10684);
nand U12283 (N_12283,N_11126,N_11017);
nand U12284 (N_12284,N_10589,N_11856);
and U12285 (N_12285,N_10793,N_10849);
xnor U12286 (N_12286,N_11745,N_10772);
or U12287 (N_12287,N_11634,N_11481);
nor U12288 (N_12288,N_11570,N_11867);
and U12289 (N_12289,N_11612,N_10525);
and U12290 (N_12290,N_11608,N_11789);
nor U12291 (N_12291,N_11094,N_10903);
or U12292 (N_12292,N_11351,N_11939);
and U12293 (N_12293,N_11888,N_11900);
nor U12294 (N_12294,N_10948,N_11243);
nor U12295 (N_12295,N_11015,N_11689);
or U12296 (N_12296,N_11166,N_11513);
nor U12297 (N_12297,N_11248,N_11566);
or U12298 (N_12298,N_11082,N_11680);
or U12299 (N_12299,N_11362,N_11710);
or U12300 (N_12300,N_10717,N_10547);
xnor U12301 (N_12301,N_11609,N_11564);
nor U12302 (N_12302,N_10931,N_11127);
nor U12303 (N_12303,N_11646,N_10558);
and U12304 (N_12304,N_11044,N_10741);
xor U12305 (N_12305,N_11961,N_10743);
or U12306 (N_12306,N_11916,N_11163);
xnor U12307 (N_12307,N_10946,N_10771);
nand U12308 (N_12308,N_11729,N_11933);
nor U12309 (N_12309,N_11423,N_10712);
nand U12310 (N_12310,N_10600,N_11063);
or U12311 (N_12311,N_11823,N_11526);
nor U12312 (N_12312,N_11029,N_11705);
xnor U12313 (N_12313,N_10746,N_11997);
nand U12314 (N_12314,N_11461,N_11589);
and U12315 (N_12315,N_11411,N_11941);
and U12316 (N_12316,N_10543,N_11173);
nand U12317 (N_12317,N_11196,N_11105);
nand U12318 (N_12318,N_11625,N_10738);
nand U12319 (N_12319,N_11892,N_11447);
xor U12320 (N_12320,N_11121,N_11312);
or U12321 (N_12321,N_10899,N_11153);
and U12322 (N_12322,N_11820,N_11337);
nor U12323 (N_12323,N_11457,N_10633);
or U12324 (N_12324,N_11536,N_11544);
and U12325 (N_12325,N_11175,N_11262);
nand U12326 (N_12326,N_10812,N_11400);
or U12327 (N_12327,N_11014,N_11470);
nor U12328 (N_12328,N_11315,N_10915);
or U12329 (N_12329,N_11307,N_10673);
or U12330 (N_12330,N_11986,N_11169);
nand U12331 (N_12331,N_11945,N_10663);
or U12332 (N_12332,N_10505,N_11914);
nand U12333 (N_12333,N_11365,N_11889);
or U12334 (N_12334,N_10605,N_11393);
nand U12335 (N_12335,N_10939,N_11960);
nor U12336 (N_12336,N_11592,N_10894);
and U12337 (N_12337,N_10727,N_10916);
or U12338 (N_12338,N_10788,N_10553);
nor U12339 (N_12339,N_11771,N_11164);
nor U12340 (N_12340,N_11416,N_10640);
or U12341 (N_12341,N_10914,N_11079);
xor U12342 (N_12342,N_11765,N_11494);
nor U12343 (N_12343,N_11860,N_11509);
and U12344 (N_12344,N_10575,N_11299);
or U12345 (N_12345,N_11976,N_11984);
or U12346 (N_12346,N_11977,N_11839);
and U12347 (N_12347,N_11557,N_11219);
nand U12348 (N_12348,N_11971,N_11317);
nor U12349 (N_12349,N_11008,N_10681);
nand U12350 (N_12350,N_10721,N_10776);
xor U12351 (N_12351,N_11038,N_10528);
nor U12352 (N_12352,N_11446,N_10688);
and U12353 (N_12353,N_11006,N_11732);
and U12354 (N_12354,N_11157,N_10960);
or U12355 (N_12355,N_11540,N_10884);
or U12356 (N_12356,N_11899,N_11348);
or U12357 (N_12357,N_11614,N_11120);
nand U12358 (N_12358,N_11292,N_11832);
nand U12359 (N_12359,N_11477,N_11328);
nand U12360 (N_12360,N_11060,N_11236);
xnor U12361 (N_12361,N_11740,N_11780);
and U12362 (N_12362,N_11054,N_11203);
or U12363 (N_12363,N_10647,N_11772);
nand U12364 (N_12364,N_11211,N_10521);
or U12365 (N_12365,N_11852,N_11198);
and U12366 (N_12366,N_10725,N_10736);
and U12367 (N_12367,N_10991,N_10785);
nand U12368 (N_12368,N_10823,N_10611);
and U12369 (N_12369,N_11701,N_11698);
or U12370 (N_12370,N_11376,N_10583);
or U12371 (N_12371,N_11582,N_11527);
or U12372 (N_12372,N_10782,N_11154);
or U12373 (N_12373,N_11573,N_10830);
nand U12374 (N_12374,N_10629,N_11360);
or U12375 (N_12375,N_10930,N_10898);
nand U12376 (N_12376,N_11632,N_11535);
nand U12377 (N_12377,N_11511,N_11883);
and U12378 (N_12378,N_10509,N_10573);
or U12379 (N_12379,N_11673,N_11123);
xor U12380 (N_12380,N_10832,N_10549);
or U12381 (N_12381,N_10856,N_10922);
nand U12382 (N_12382,N_10566,N_10632);
nor U12383 (N_12383,N_11830,N_11483);
nand U12384 (N_12384,N_11894,N_11216);
nand U12385 (N_12385,N_11160,N_11768);
nand U12386 (N_12386,N_11209,N_11779);
and U12387 (N_12387,N_11052,N_10796);
nor U12388 (N_12388,N_11110,N_11747);
or U12389 (N_12389,N_11240,N_11390);
nand U12390 (N_12390,N_11141,N_10826);
xor U12391 (N_12391,N_11026,N_10869);
nand U12392 (N_12392,N_11448,N_11606);
nand U12393 (N_12393,N_10892,N_11469);
and U12394 (N_12394,N_11370,N_10924);
and U12395 (N_12395,N_11260,N_11081);
or U12396 (N_12396,N_11727,N_11399);
xnor U12397 (N_12397,N_11810,N_10804);
nand U12398 (N_12398,N_11095,N_11381);
nor U12399 (N_12399,N_11537,N_11653);
and U12400 (N_12400,N_10822,N_10900);
nor U12401 (N_12401,N_11493,N_11350);
nor U12402 (N_12402,N_11069,N_11182);
nor U12403 (N_12403,N_11674,N_11516);
or U12404 (N_12404,N_11043,N_11237);
nor U12405 (N_12405,N_11616,N_11031);
or U12406 (N_12406,N_11897,N_11186);
nor U12407 (N_12407,N_11699,N_11672);
nor U12408 (N_12408,N_11556,N_10520);
nor U12409 (N_12409,N_10557,N_11929);
or U12410 (N_12410,N_10867,N_11605);
and U12411 (N_12411,N_10835,N_11131);
nor U12412 (N_12412,N_10638,N_11869);
and U12413 (N_12413,N_11979,N_10813);
nand U12414 (N_12414,N_10590,N_11969);
xor U12415 (N_12415,N_11319,N_11487);
nor U12416 (N_12416,N_11451,N_11065);
or U12417 (N_12417,N_11139,N_10733);
or U12418 (N_12418,N_11259,N_11594);
or U12419 (N_12419,N_11681,N_11035);
nor U12420 (N_12420,N_10809,N_10979);
or U12421 (N_12421,N_10799,N_10686);
nor U12422 (N_12422,N_11734,N_10514);
nand U12423 (N_12423,N_10650,N_11412);
and U12424 (N_12424,N_11067,N_10921);
nand U12425 (N_12425,N_11934,N_11574);
nand U12426 (N_12426,N_11242,N_11563);
or U12427 (N_12427,N_10532,N_10855);
or U12428 (N_12428,N_11966,N_11584);
nand U12429 (N_12429,N_11846,N_11843);
nor U12430 (N_12430,N_10901,N_11604);
or U12431 (N_12431,N_11981,N_11538);
and U12432 (N_12432,N_11178,N_10726);
nor U12433 (N_12433,N_11189,N_10502);
nand U12434 (N_12434,N_10845,N_10619);
and U12435 (N_12435,N_11518,N_11191);
xnor U12436 (N_12436,N_10701,N_10511);
nor U12437 (N_12437,N_11032,N_11402);
or U12438 (N_12438,N_11709,N_11129);
and U12439 (N_12439,N_11554,N_11978);
nand U12440 (N_12440,N_10908,N_10797);
xnor U12441 (N_12441,N_11415,N_11567);
and U12442 (N_12442,N_11250,N_10612);
nand U12443 (N_12443,N_11233,N_11904);
nand U12444 (N_12444,N_11322,N_10588);
nand U12445 (N_12445,N_11520,N_11125);
and U12446 (N_12446,N_11172,N_11758);
nor U12447 (N_12447,N_11249,N_10961);
or U12448 (N_12448,N_10653,N_11385);
and U12449 (N_12449,N_11431,N_11600);
xor U12450 (N_12450,N_11548,N_11283);
nor U12451 (N_12451,N_11045,N_10515);
xor U12452 (N_12452,N_10897,N_10729);
or U12453 (N_12453,N_11963,N_10976);
nand U12454 (N_12454,N_10866,N_10720);
or U12455 (N_12455,N_11290,N_11756);
nor U12456 (N_12456,N_11514,N_11009);
nor U12457 (N_12457,N_10516,N_11580);
or U12458 (N_12458,N_11987,N_10784);
or U12459 (N_12459,N_11737,N_11176);
or U12460 (N_12460,N_11601,N_11558);
xnor U12461 (N_12461,N_10836,N_10965);
nand U12462 (N_12462,N_11433,N_11906);
xnor U12463 (N_12463,N_11104,N_10992);
nor U12464 (N_12464,N_10503,N_11268);
and U12465 (N_12465,N_11389,N_10757);
nand U12466 (N_12466,N_11227,N_11426);
or U12467 (N_12467,N_11757,N_11296);
or U12468 (N_12468,N_10719,N_11827);
nand U12469 (N_12469,N_10693,N_11657);
and U12470 (N_12470,N_10658,N_11086);
nand U12471 (N_12471,N_11118,N_11742);
and U12472 (N_12472,N_11495,N_10694);
nand U12473 (N_12473,N_11712,N_10982);
or U12474 (N_12474,N_11055,N_11310);
nand U12475 (N_12475,N_11392,N_10716);
nor U12476 (N_12476,N_11488,N_10513);
and U12477 (N_12477,N_10910,N_10507);
nand U12478 (N_12478,N_11836,N_11553);
nor U12479 (N_12479,N_11108,N_10569);
nor U12480 (N_12480,N_10527,N_11475);
or U12481 (N_12481,N_11896,N_11898);
or U12482 (N_12482,N_11058,N_10764);
and U12483 (N_12483,N_11442,N_11675);
and U12484 (N_12484,N_11875,N_11671);
xor U12485 (N_12485,N_10918,N_10714);
or U12486 (N_12486,N_11329,N_11550);
nor U12487 (N_12487,N_10689,N_11034);
or U12488 (N_12488,N_10628,N_11199);
nand U12489 (N_12489,N_10651,N_11440);
nand U12490 (N_12490,N_10574,N_11547);
or U12491 (N_12491,N_10607,N_10853);
or U12492 (N_12492,N_11266,N_10696);
nand U12493 (N_12493,N_11354,N_11364);
nor U12494 (N_12494,N_11320,N_10581);
nand U12495 (N_12495,N_10526,N_11638);
nand U12496 (N_12496,N_11598,N_11948);
nor U12497 (N_12497,N_11486,N_11829);
or U12498 (N_12498,N_11316,N_11403);
nand U12499 (N_12499,N_11187,N_10890);
nor U12500 (N_12500,N_11523,N_11352);
or U12501 (N_12501,N_11644,N_10749);
or U12502 (N_12502,N_10625,N_11308);
or U12503 (N_12503,N_11967,N_10923);
nand U12504 (N_12504,N_11218,N_11050);
xor U12505 (N_12505,N_11833,N_10941);
nand U12506 (N_12506,N_11217,N_11491);
nor U12507 (N_12507,N_11039,N_11132);
and U12508 (N_12508,N_11011,N_10977);
nor U12509 (N_12509,N_10997,N_11247);
or U12510 (N_12510,N_11499,N_11761);
nor U12511 (N_12511,N_10533,N_10586);
nor U12512 (N_12512,N_11215,N_11905);
or U12513 (N_12513,N_11726,N_11591);
nand U12514 (N_12514,N_10755,N_11023);
nand U12515 (N_12515,N_11168,N_11273);
nor U12516 (N_12516,N_11437,N_10902);
or U12517 (N_12517,N_11655,N_11452);
or U12518 (N_12518,N_11572,N_11145);
nand U12519 (N_12519,N_10807,N_11272);
nand U12520 (N_12520,N_10584,N_10730);
or U12521 (N_12521,N_11456,N_11590);
nor U12522 (N_12522,N_11012,N_11932);
xor U12523 (N_12523,N_10675,N_11305);
nor U12524 (N_12524,N_10954,N_10806);
and U12525 (N_12525,N_11473,N_10816);
nand U12526 (N_12526,N_11854,N_10616);
xnor U12527 (N_12527,N_10646,N_11267);
and U12528 (N_12528,N_11610,N_11677);
nor U12529 (N_12529,N_11394,N_11928);
xnor U12530 (N_12530,N_11454,N_11866);
and U12531 (N_12531,N_11946,N_10504);
nor U12532 (N_12532,N_11759,N_11970);
xor U12533 (N_12533,N_11588,N_10821);
nand U12534 (N_12534,N_11667,N_11326);
nand U12535 (N_12535,N_11773,N_11597);
nand U12536 (N_12536,N_11676,N_11102);
and U12537 (N_12537,N_11811,N_11251);
nand U12538 (N_12538,N_11476,N_10601);
nor U12539 (N_12539,N_11404,N_10926);
and U12540 (N_12540,N_11794,N_10987);
xnor U12541 (N_12541,N_11323,N_11057);
nor U12542 (N_12542,N_11746,N_11353);
and U12543 (N_12543,N_11814,N_10851);
nand U12544 (N_12544,N_11235,N_11670);
or U12545 (N_12545,N_10614,N_10580);
or U12546 (N_12546,N_10537,N_10671);
or U12547 (N_12547,N_10635,N_10850);
or U12548 (N_12548,N_10501,N_10973);
nor U12549 (N_12549,N_10700,N_10706);
or U12550 (N_12550,N_11478,N_11649);
nor U12551 (N_12551,N_11001,N_11498);
or U12552 (N_12552,N_10990,N_11490);
and U12553 (N_12553,N_10998,N_11314);
nor U12554 (N_12554,N_10949,N_10554);
xnor U12555 (N_12555,N_10621,N_11177);
or U12556 (N_12556,N_10728,N_11622);
and U12557 (N_12557,N_11788,N_10969);
nor U12558 (N_12558,N_10620,N_11135);
or U12559 (N_12559,N_11074,N_11754);
or U12560 (N_12560,N_10942,N_11255);
or U12561 (N_12561,N_11419,N_11244);
and U12562 (N_12562,N_11784,N_11777);
xor U12563 (N_12563,N_10666,N_11238);
and U12564 (N_12564,N_11576,N_11922);
or U12565 (N_12565,N_11005,N_10983);
and U12566 (N_12566,N_11512,N_11409);
and U12567 (N_12567,N_11641,N_10964);
and U12568 (N_12568,N_10752,N_10873);
nor U12569 (N_12569,N_11245,N_10713);
nand U12570 (N_12570,N_10508,N_10993);
or U12571 (N_12571,N_10810,N_10760);
xor U12572 (N_12572,N_11443,N_11669);
xnor U12573 (N_12573,N_11422,N_11931);
or U12574 (N_12574,N_11859,N_11620);
and U12575 (N_12575,N_10636,N_10560);
xnor U12576 (N_12576,N_11282,N_11821);
and U12577 (N_12577,N_10868,N_11847);
and U12578 (N_12578,N_11502,N_11721);
and U12579 (N_12579,N_11725,N_11781);
xnor U12580 (N_12580,N_10599,N_10608);
and U12581 (N_12581,N_10699,N_11464);
or U12582 (N_12582,N_11874,N_10564);
nand U12583 (N_12583,N_11087,N_10711);
nand U12584 (N_12584,N_11384,N_10724);
or U12585 (N_12585,N_11992,N_10834);
nor U12586 (N_12586,N_10820,N_11212);
and U12587 (N_12587,N_11356,N_11692);
nor U12588 (N_12588,N_11626,N_11753);
and U12589 (N_12589,N_10692,N_11942);
nand U12590 (N_12590,N_11694,N_10790);
or U12591 (N_12591,N_10592,N_11075);
and U12592 (N_12592,N_10747,N_10585);
and U12593 (N_12593,N_11926,N_11264);
nor U12594 (N_12594,N_11907,N_11707);
or U12595 (N_12595,N_10952,N_11016);
nor U12596 (N_12596,N_11639,N_11024);
and U12597 (N_12597,N_11837,N_11295);
and U12598 (N_12598,N_11887,N_11815);
nand U12599 (N_12599,N_10531,N_11845);
nor U12600 (N_12600,N_11226,N_10959);
nor U12601 (N_12601,N_10756,N_11463);
nand U12602 (N_12602,N_10972,N_11336);
or U12603 (N_12603,N_10639,N_11155);
and U12604 (N_12604,N_11302,N_11321);
and U12605 (N_12605,N_11396,N_11335);
nor U12606 (N_12606,N_10951,N_11787);
nand U12607 (N_12607,N_11080,N_10637);
xor U12608 (N_12608,N_11805,N_10556);
nand U12609 (N_12609,N_11134,N_11345);
nor U12610 (N_12610,N_10844,N_11338);
nand U12611 (N_12611,N_11650,N_10827);
nor U12612 (N_12612,N_11201,N_11798);
nand U12613 (N_12613,N_11306,N_11041);
or U12614 (N_12614,N_11036,N_10674);
and U12615 (N_12615,N_11165,N_11690);
and U12616 (N_12616,N_10751,N_10510);
nand U12617 (N_12617,N_10679,N_11441);
nand U12618 (N_12618,N_11873,N_11280);
or U12619 (N_12619,N_10742,N_10862);
nor U12620 (N_12620,N_11161,N_11021);
nor U12621 (N_12621,N_10778,N_11687);
nor U12622 (N_12622,N_11184,N_11386);
nor U12623 (N_12623,N_11252,N_11115);
or U12624 (N_12624,N_11802,N_10825);
and U12625 (N_12625,N_11382,N_11999);
or U12626 (N_12626,N_11912,N_11628);
or U12627 (N_12627,N_10854,N_10678);
and U12628 (N_12628,N_10909,N_11185);
xor U12629 (N_12629,N_10664,N_10945);
or U12630 (N_12630,N_10680,N_11444);
or U12631 (N_12631,N_11293,N_11817);
and U12632 (N_12632,N_11631,N_10852);
nor U12633 (N_12633,N_10519,N_11030);
and U12634 (N_12634,N_11506,N_11682);
nand U12635 (N_12635,N_10795,N_10766);
nand U12636 (N_12636,N_11816,N_10829);
and U12637 (N_12637,N_11333,N_10595);
nand U12638 (N_12638,N_11901,N_10702);
nor U12639 (N_12639,N_10932,N_10548);
and U12640 (N_12640,N_11148,N_10802);
or U12641 (N_12641,N_11529,N_11953);
xor U12642 (N_12642,N_10522,N_11760);
nand U12643 (N_12643,N_11207,N_10631);
nand U12644 (N_12644,N_11733,N_10739);
or U12645 (N_12645,N_11533,N_10695);
nand U12646 (N_12646,N_11693,N_11122);
or U12647 (N_12647,N_11545,N_11804);
and U12648 (N_12648,N_10875,N_11640);
or U12649 (N_12649,N_11599,N_11964);
nand U12650 (N_12650,N_11950,N_11561);
nand U12651 (N_12651,N_11801,N_11144);
and U12652 (N_12652,N_10732,N_11844);
nor U12653 (N_12653,N_10955,N_11508);
or U12654 (N_12654,N_10603,N_10886);
nor U12655 (N_12655,N_11256,N_11924);
or U12656 (N_12656,N_10546,N_11718);
and U12657 (N_12657,N_10540,N_11228);
and U12658 (N_12658,N_11930,N_11344);
and U12659 (N_12659,N_11406,N_11736);
nor U12660 (N_12660,N_11343,N_10958);
or U12661 (N_12661,N_11797,N_11886);
nor U12662 (N_12662,N_10815,N_11056);
or U12663 (N_12663,N_10984,N_11462);
and U12664 (N_12664,N_11420,N_11786);
nand U12665 (N_12665,N_11636,N_11890);
nor U12666 (N_12666,N_11995,N_11515);
or U12667 (N_12667,N_11192,N_11903);
nor U12668 (N_12668,N_10879,N_10907);
nand U12669 (N_12669,N_10863,N_11849);
xor U12670 (N_12670,N_11496,N_11808);
nand U12671 (N_12671,N_11099,N_11149);
or U12672 (N_12672,N_11339,N_11276);
and U12673 (N_12673,N_11711,N_10837);
nand U12674 (N_12674,N_10538,N_11373);
or U12675 (N_12675,N_11205,N_11659);
nor U12676 (N_12676,N_10841,N_11484);
or U12677 (N_12677,N_11286,N_11559);
or U12678 (N_12678,N_11521,N_11253);
or U12679 (N_12679,N_11940,N_10865);
xnor U12680 (N_12680,N_11410,N_10774);
nor U12681 (N_12681,N_11284,N_11587);
or U12682 (N_12682,N_10811,N_11991);
xor U12683 (N_12683,N_10944,N_11560);
xnor U12684 (N_12684,N_10792,N_11871);
or U12685 (N_12685,N_11436,N_11818);
and U12686 (N_12686,N_11519,N_11783);
nor U12687 (N_12687,N_10529,N_10544);
nand U12688 (N_12688,N_10881,N_10940);
nor U12689 (N_12689,N_11750,N_11239);
or U12690 (N_12690,N_11863,N_10783);
nor U12691 (N_12691,N_11778,N_10768);
or U12692 (N_12692,N_11397,N_11858);
xnor U12693 (N_12693,N_10805,N_10551);
nand U12694 (N_12694,N_11414,N_11881);
and U12695 (N_12695,N_11882,N_11263);
or U12696 (N_12696,N_10917,N_11234);
or U12697 (N_12697,N_11204,N_11507);
or U12698 (N_12698,N_11957,N_11208);
nor U12699 (N_12699,N_10878,N_11927);
and U12700 (N_12700,N_10715,N_10787);
or U12701 (N_12701,N_10963,N_11257);
and U12702 (N_12702,N_11300,N_11925);
nand U12703 (N_12703,N_10999,N_11555);
and U12704 (N_12704,N_11114,N_11876);
or U12705 (N_12705,N_11246,N_11459);
or U12706 (N_12706,N_11730,N_11696);
nor U12707 (N_12707,N_10920,N_10754);
or U12708 (N_12708,N_11408,N_11531);
or U12709 (N_12709,N_11764,N_10626);
nor U12710 (N_12710,N_11222,N_10996);
or U12711 (N_12711,N_11180,N_11806);
xnor U12712 (N_12712,N_10786,N_10555);
or U12713 (N_12713,N_11958,N_11077);
nor U12714 (N_12714,N_10843,N_11466);
or U12715 (N_12715,N_10697,N_11159);
xor U12716 (N_12716,N_11551,N_10545);
xor U12717 (N_12717,N_10985,N_10655);
nor U12718 (N_12718,N_11785,N_11418);
nor U12719 (N_12719,N_11803,N_11910);
nand U12720 (N_12720,N_11735,N_11083);
or U12721 (N_12721,N_10934,N_11471);
or U12722 (N_12722,N_10563,N_11624);
and U12723 (N_12723,N_11790,N_11347);
and U12724 (N_12724,N_11920,N_11068);
xor U12725 (N_12725,N_10744,N_11124);
nand U12726 (N_12726,N_10667,N_11064);
nand U12727 (N_12727,N_10935,N_11098);
nand U12728 (N_12728,N_11089,N_10610);
or U12729 (N_12729,N_11936,N_11107);
nand U12730 (N_12730,N_11002,N_11407);
nor U12731 (N_12731,N_11438,N_10758);
xor U12732 (N_12732,N_11294,N_10980);
nor U12733 (N_12733,N_11880,N_11989);
or U12734 (N_12734,N_10762,N_11171);
and U12735 (N_12735,N_11776,N_11724);
and U12736 (N_12736,N_11917,N_10682);
and U12737 (N_12737,N_11028,N_10956);
nor U12738 (N_12738,N_10518,N_10687);
nor U12739 (N_12739,N_11073,N_11621);
xor U12740 (N_12740,N_10587,N_10936);
nand U12741 (N_12741,N_11775,N_11915);
nand U12742 (N_12742,N_11241,N_11224);
or U12743 (N_12743,N_11795,N_11656);
or U12744 (N_12744,N_10947,N_11170);
and U12745 (N_12745,N_11379,N_10808);
or U12746 (N_12746,N_11288,N_11532);
and U12747 (N_12747,N_10871,N_11770);
and U12748 (N_12748,N_11793,N_11421);
nand U12749 (N_12749,N_11398,N_11202);
and U12750 (N_12750,N_11913,N_11168);
and U12751 (N_12751,N_10557,N_11599);
nor U12752 (N_12752,N_11440,N_11394);
nand U12753 (N_12753,N_11856,N_11484);
nor U12754 (N_12754,N_10763,N_11468);
and U12755 (N_12755,N_11193,N_11483);
or U12756 (N_12756,N_11491,N_11570);
or U12757 (N_12757,N_11875,N_11658);
nor U12758 (N_12758,N_11692,N_11562);
xnor U12759 (N_12759,N_11966,N_11801);
or U12760 (N_12760,N_11285,N_11509);
or U12761 (N_12761,N_11322,N_11514);
or U12762 (N_12762,N_11481,N_11865);
nand U12763 (N_12763,N_11396,N_11519);
or U12764 (N_12764,N_11474,N_11573);
and U12765 (N_12765,N_11044,N_11995);
nor U12766 (N_12766,N_11235,N_10824);
xnor U12767 (N_12767,N_10640,N_10592);
nand U12768 (N_12768,N_10850,N_10736);
nor U12769 (N_12769,N_11185,N_11356);
nor U12770 (N_12770,N_11480,N_11937);
or U12771 (N_12771,N_10946,N_11948);
nor U12772 (N_12772,N_11865,N_11808);
nand U12773 (N_12773,N_10669,N_10971);
or U12774 (N_12774,N_10840,N_11154);
and U12775 (N_12775,N_11198,N_10965);
or U12776 (N_12776,N_10959,N_11257);
xor U12777 (N_12777,N_11867,N_10511);
and U12778 (N_12778,N_10758,N_11540);
nand U12779 (N_12779,N_11348,N_11626);
nor U12780 (N_12780,N_11579,N_11282);
nand U12781 (N_12781,N_11684,N_11129);
or U12782 (N_12782,N_11454,N_11096);
and U12783 (N_12783,N_10545,N_11804);
or U12784 (N_12784,N_11412,N_11494);
nand U12785 (N_12785,N_11051,N_11781);
nor U12786 (N_12786,N_11601,N_11917);
nand U12787 (N_12787,N_11088,N_10646);
nand U12788 (N_12788,N_10962,N_10527);
nor U12789 (N_12789,N_11749,N_11400);
or U12790 (N_12790,N_11870,N_11619);
nand U12791 (N_12791,N_11076,N_11887);
nand U12792 (N_12792,N_10535,N_11286);
and U12793 (N_12793,N_11731,N_11432);
or U12794 (N_12794,N_10769,N_10774);
and U12795 (N_12795,N_11997,N_11968);
and U12796 (N_12796,N_10540,N_11377);
nor U12797 (N_12797,N_10648,N_10520);
and U12798 (N_12798,N_11675,N_10544);
nand U12799 (N_12799,N_11369,N_11661);
xnor U12800 (N_12800,N_11323,N_11316);
and U12801 (N_12801,N_11551,N_11901);
or U12802 (N_12802,N_11650,N_10908);
or U12803 (N_12803,N_11031,N_11366);
and U12804 (N_12804,N_11705,N_10733);
xor U12805 (N_12805,N_10695,N_10965);
nand U12806 (N_12806,N_11584,N_11662);
or U12807 (N_12807,N_10835,N_11790);
and U12808 (N_12808,N_11889,N_11556);
or U12809 (N_12809,N_11680,N_11931);
and U12810 (N_12810,N_10595,N_11348);
or U12811 (N_12811,N_11890,N_11477);
nor U12812 (N_12812,N_10734,N_11608);
nor U12813 (N_12813,N_10641,N_10754);
or U12814 (N_12814,N_11060,N_11861);
nand U12815 (N_12815,N_10832,N_11271);
nand U12816 (N_12816,N_11428,N_11342);
and U12817 (N_12817,N_11352,N_10873);
nor U12818 (N_12818,N_11088,N_11639);
nor U12819 (N_12819,N_10710,N_10906);
and U12820 (N_12820,N_11429,N_11295);
or U12821 (N_12821,N_10828,N_10610);
or U12822 (N_12822,N_11695,N_11776);
xnor U12823 (N_12823,N_11405,N_10736);
or U12824 (N_12824,N_11642,N_10604);
nor U12825 (N_12825,N_11862,N_11743);
or U12826 (N_12826,N_11440,N_11166);
or U12827 (N_12827,N_11999,N_11885);
nor U12828 (N_12828,N_11557,N_10929);
nand U12829 (N_12829,N_10974,N_10616);
and U12830 (N_12830,N_10757,N_11298);
nor U12831 (N_12831,N_11776,N_11915);
and U12832 (N_12832,N_10718,N_11264);
nor U12833 (N_12833,N_10922,N_10849);
nand U12834 (N_12834,N_11190,N_11247);
or U12835 (N_12835,N_11286,N_11652);
or U12836 (N_12836,N_10674,N_11906);
and U12837 (N_12837,N_11982,N_11160);
or U12838 (N_12838,N_10778,N_10807);
and U12839 (N_12839,N_11697,N_11518);
nand U12840 (N_12840,N_10621,N_11968);
nand U12841 (N_12841,N_10653,N_10909);
nand U12842 (N_12842,N_11665,N_11479);
or U12843 (N_12843,N_11419,N_11627);
xnor U12844 (N_12844,N_10857,N_11086);
xor U12845 (N_12845,N_11950,N_11027);
and U12846 (N_12846,N_11883,N_10693);
xor U12847 (N_12847,N_10634,N_11797);
and U12848 (N_12848,N_11626,N_11244);
nor U12849 (N_12849,N_10649,N_10738);
and U12850 (N_12850,N_11829,N_11714);
nand U12851 (N_12851,N_11749,N_11705);
nor U12852 (N_12852,N_10777,N_11688);
and U12853 (N_12853,N_11358,N_11698);
nor U12854 (N_12854,N_11111,N_10873);
nand U12855 (N_12855,N_10586,N_11693);
or U12856 (N_12856,N_11234,N_11946);
or U12857 (N_12857,N_10702,N_11648);
or U12858 (N_12858,N_11737,N_11589);
and U12859 (N_12859,N_11257,N_11961);
or U12860 (N_12860,N_10638,N_10881);
xor U12861 (N_12861,N_11317,N_10697);
and U12862 (N_12862,N_10886,N_11365);
and U12863 (N_12863,N_11003,N_11292);
nand U12864 (N_12864,N_11798,N_10844);
and U12865 (N_12865,N_10718,N_11956);
nand U12866 (N_12866,N_10590,N_11132);
nor U12867 (N_12867,N_11638,N_11251);
nand U12868 (N_12868,N_10725,N_11531);
nand U12869 (N_12869,N_10510,N_11004);
or U12870 (N_12870,N_11749,N_10551);
nand U12871 (N_12871,N_11887,N_11712);
and U12872 (N_12872,N_10707,N_10516);
nand U12873 (N_12873,N_11806,N_11054);
and U12874 (N_12874,N_11319,N_11188);
nand U12875 (N_12875,N_11939,N_10957);
nor U12876 (N_12876,N_11989,N_11423);
and U12877 (N_12877,N_10813,N_11444);
nor U12878 (N_12878,N_11839,N_10971);
nor U12879 (N_12879,N_11576,N_10514);
and U12880 (N_12880,N_11540,N_11510);
nor U12881 (N_12881,N_11918,N_10674);
and U12882 (N_12882,N_11080,N_11022);
xnor U12883 (N_12883,N_11024,N_11266);
or U12884 (N_12884,N_10805,N_11854);
nand U12885 (N_12885,N_11309,N_10727);
or U12886 (N_12886,N_10725,N_10576);
nand U12887 (N_12887,N_11037,N_11689);
nand U12888 (N_12888,N_10863,N_10981);
or U12889 (N_12889,N_11393,N_11994);
and U12890 (N_12890,N_11849,N_10895);
and U12891 (N_12891,N_10645,N_11581);
xnor U12892 (N_12892,N_11910,N_10585);
or U12893 (N_12893,N_11958,N_11428);
or U12894 (N_12894,N_11380,N_11684);
nor U12895 (N_12895,N_10869,N_11890);
and U12896 (N_12896,N_11269,N_10709);
nor U12897 (N_12897,N_10603,N_11195);
nand U12898 (N_12898,N_10886,N_11631);
nand U12899 (N_12899,N_11130,N_11159);
nand U12900 (N_12900,N_11942,N_11605);
nor U12901 (N_12901,N_11019,N_11264);
nand U12902 (N_12902,N_10503,N_10663);
nand U12903 (N_12903,N_10851,N_11170);
nand U12904 (N_12904,N_10542,N_11233);
nand U12905 (N_12905,N_11369,N_11061);
or U12906 (N_12906,N_11945,N_11079);
and U12907 (N_12907,N_11049,N_11404);
or U12908 (N_12908,N_11633,N_11058);
and U12909 (N_12909,N_11418,N_11359);
and U12910 (N_12910,N_11471,N_11428);
nor U12911 (N_12911,N_11206,N_10796);
or U12912 (N_12912,N_11357,N_11314);
nor U12913 (N_12913,N_11267,N_11630);
nand U12914 (N_12914,N_11728,N_10967);
or U12915 (N_12915,N_11299,N_10539);
nor U12916 (N_12916,N_10838,N_11890);
and U12917 (N_12917,N_11013,N_11143);
or U12918 (N_12918,N_11373,N_11284);
or U12919 (N_12919,N_11365,N_10737);
nand U12920 (N_12920,N_11455,N_10575);
and U12921 (N_12921,N_11830,N_11227);
or U12922 (N_12922,N_11914,N_11800);
or U12923 (N_12923,N_11043,N_10921);
and U12924 (N_12924,N_10612,N_11600);
xnor U12925 (N_12925,N_11084,N_10732);
nor U12926 (N_12926,N_11903,N_11105);
or U12927 (N_12927,N_11352,N_11555);
nand U12928 (N_12928,N_11335,N_11167);
or U12929 (N_12929,N_11973,N_11385);
nor U12930 (N_12930,N_11200,N_11348);
xnor U12931 (N_12931,N_11018,N_11714);
nor U12932 (N_12932,N_10641,N_11254);
nand U12933 (N_12933,N_11800,N_10579);
nor U12934 (N_12934,N_11403,N_11001);
nand U12935 (N_12935,N_10643,N_11383);
xor U12936 (N_12936,N_10627,N_10517);
nand U12937 (N_12937,N_11453,N_11214);
or U12938 (N_12938,N_10914,N_10597);
or U12939 (N_12939,N_11973,N_10858);
nor U12940 (N_12940,N_11833,N_10562);
nor U12941 (N_12941,N_11404,N_11734);
and U12942 (N_12942,N_10843,N_11333);
and U12943 (N_12943,N_11941,N_10955);
nor U12944 (N_12944,N_10929,N_10993);
or U12945 (N_12945,N_11276,N_11347);
xnor U12946 (N_12946,N_10718,N_11703);
or U12947 (N_12947,N_10693,N_11518);
xor U12948 (N_12948,N_11629,N_10999);
nor U12949 (N_12949,N_11775,N_10844);
or U12950 (N_12950,N_11309,N_11644);
nor U12951 (N_12951,N_11044,N_11329);
or U12952 (N_12952,N_11113,N_11400);
nand U12953 (N_12953,N_11159,N_11858);
nand U12954 (N_12954,N_11664,N_11547);
nor U12955 (N_12955,N_10633,N_11957);
xnor U12956 (N_12956,N_11020,N_10811);
nor U12957 (N_12957,N_11541,N_11618);
nor U12958 (N_12958,N_11289,N_11442);
or U12959 (N_12959,N_11655,N_11225);
nor U12960 (N_12960,N_10821,N_11142);
or U12961 (N_12961,N_11341,N_11703);
and U12962 (N_12962,N_11664,N_10578);
or U12963 (N_12963,N_11513,N_11276);
nor U12964 (N_12964,N_10734,N_11534);
and U12965 (N_12965,N_11266,N_11740);
or U12966 (N_12966,N_10956,N_11950);
nor U12967 (N_12967,N_10702,N_11295);
nand U12968 (N_12968,N_11735,N_11252);
or U12969 (N_12969,N_10849,N_10929);
or U12970 (N_12970,N_10979,N_11407);
and U12971 (N_12971,N_11145,N_11781);
and U12972 (N_12972,N_10672,N_11675);
or U12973 (N_12973,N_11127,N_10565);
and U12974 (N_12974,N_11168,N_10927);
nand U12975 (N_12975,N_10815,N_10748);
nand U12976 (N_12976,N_10806,N_10585);
nor U12977 (N_12977,N_11528,N_11763);
nor U12978 (N_12978,N_11482,N_10775);
nor U12979 (N_12979,N_11169,N_10775);
and U12980 (N_12980,N_10902,N_10735);
and U12981 (N_12981,N_10620,N_11890);
nand U12982 (N_12982,N_11255,N_11158);
nand U12983 (N_12983,N_10709,N_11857);
nand U12984 (N_12984,N_10943,N_11450);
nand U12985 (N_12985,N_10729,N_11844);
nor U12986 (N_12986,N_11921,N_11529);
or U12987 (N_12987,N_11880,N_10995);
and U12988 (N_12988,N_11490,N_11279);
nor U12989 (N_12989,N_10796,N_11078);
and U12990 (N_12990,N_10562,N_11831);
xor U12991 (N_12991,N_11265,N_11379);
or U12992 (N_12992,N_11987,N_10827);
and U12993 (N_12993,N_11150,N_11791);
nor U12994 (N_12994,N_11276,N_10678);
and U12995 (N_12995,N_11056,N_11551);
nand U12996 (N_12996,N_11879,N_11050);
nand U12997 (N_12997,N_11690,N_11994);
and U12998 (N_12998,N_11476,N_11114);
or U12999 (N_12999,N_10660,N_10787);
nand U13000 (N_13000,N_11314,N_11887);
nor U13001 (N_13001,N_10788,N_11469);
or U13002 (N_13002,N_11992,N_11896);
xnor U13003 (N_13003,N_11563,N_10929);
or U13004 (N_13004,N_11882,N_10840);
and U13005 (N_13005,N_11079,N_10952);
and U13006 (N_13006,N_11931,N_10625);
nand U13007 (N_13007,N_10595,N_11435);
or U13008 (N_13008,N_11347,N_11079);
nand U13009 (N_13009,N_10929,N_10732);
or U13010 (N_13010,N_11768,N_11366);
nand U13011 (N_13011,N_10665,N_10747);
nor U13012 (N_13012,N_11711,N_10683);
and U13013 (N_13013,N_11705,N_11217);
and U13014 (N_13014,N_10534,N_11624);
or U13015 (N_13015,N_11126,N_11427);
and U13016 (N_13016,N_10845,N_11442);
or U13017 (N_13017,N_11682,N_10667);
and U13018 (N_13018,N_11066,N_11815);
and U13019 (N_13019,N_10595,N_10790);
nor U13020 (N_13020,N_11783,N_10975);
or U13021 (N_13021,N_11611,N_11722);
nand U13022 (N_13022,N_11162,N_11925);
and U13023 (N_13023,N_11795,N_10555);
nand U13024 (N_13024,N_11170,N_11005);
nor U13025 (N_13025,N_11699,N_10705);
or U13026 (N_13026,N_10550,N_10597);
or U13027 (N_13027,N_11802,N_11748);
and U13028 (N_13028,N_11239,N_11944);
or U13029 (N_13029,N_11207,N_11097);
and U13030 (N_13030,N_10734,N_11731);
nand U13031 (N_13031,N_10752,N_11077);
xnor U13032 (N_13032,N_11008,N_11636);
or U13033 (N_13033,N_10614,N_10746);
xor U13034 (N_13034,N_11523,N_10766);
or U13035 (N_13035,N_11001,N_10526);
nor U13036 (N_13036,N_11019,N_10836);
or U13037 (N_13037,N_11020,N_10814);
xor U13038 (N_13038,N_11793,N_11935);
and U13039 (N_13039,N_11260,N_10899);
and U13040 (N_13040,N_10985,N_10956);
and U13041 (N_13041,N_11872,N_11797);
or U13042 (N_13042,N_10757,N_10865);
and U13043 (N_13043,N_10744,N_11886);
or U13044 (N_13044,N_11229,N_11950);
or U13045 (N_13045,N_10756,N_10802);
or U13046 (N_13046,N_10507,N_11187);
nor U13047 (N_13047,N_11708,N_11220);
nor U13048 (N_13048,N_11287,N_11142);
nand U13049 (N_13049,N_11178,N_10602);
nor U13050 (N_13050,N_11083,N_11464);
nand U13051 (N_13051,N_11951,N_11295);
nor U13052 (N_13052,N_10502,N_11044);
nand U13053 (N_13053,N_10694,N_10568);
nand U13054 (N_13054,N_10759,N_11330);
nand U13055 (N_13055,N_10561,N_11479);
nor U13056 (N_13056,N_11575,N_11091);
nor U13057 (N_13057,N_11700,N_11114);
nor U13058 (N_13058,N_11462,N_10786);
nor U13059 (N_13059,N_11565,N_11937);
or U13060 (N_13060,N_11533,N_11360);
or U13061 (N_13061,N_10568,N_11880);
nand U13062 (N_13062,N_11923,N_11048);
or U13063 (N_13063,N_10934,N_11410);
xor U13064 (N_13064,N_11865,N_11314);
or U13065 (N_13065,N_10570,N_11882);
and U13066 (N_13066,N_11287,N_10904);
nand U13067 (N_13067,N_11390,N_11706);
nand U13068 (N_13068,N_11801,N_11794);
nor U13069 (N_13069,N_11784,N_11432);
and U13070 (N_13070,N_11874,N_11291);
or U13071 (N_13071,N_10712,N_10603);
nor U13072 (N_13072,N_11289,N_11261);
nand U13073 (N_13073,N_11046,N_10669);
or U13074 (N_13074,N_11589,N_10874);
and U13075 (N_13075,N_11768,N_11846);
nand U13076 (N_13076,N_11028,N_11209);
nor U13077 (N_13077,N_10929,N_10580);
and U13078 (N_13078,N_11535,N_11968);
nand U13079 (N_13079,N_11617,N_10586);
nor U13080 (N_13080,N_11828,N_11644);
or U13081 (N_13081,N_10864,N_11580);
or U13082 (N_13082,N_11988,N_11728);
nor U13083 (N_13083,N_10961,N_11866);
and U13084 (N_13084,N_10942,N_11669);
nor U13085 (N_13085,N_10791,N_11816);
nand U13086 (N_13086,N_10526,N_10518);
or U13087 (N_13087,N_11368,N_10714);
and U13088 (N_13088,N_10851,N_10661);
nor U13089 (N_13089,N_10885,N_11359);
nor U13090 (N_13090,N_11321,N_10544);
or U13091 (N_13091,N_11069,N_11553);
and U13092 (N_13092,N_11328,N_10565);
and U13093 (N_13093,N_10739,N_10779);
or U13094 (N_13094,N_11374,N_10804);
nand U13095 (N_13095,N_11838,N_11406);
and U13096 (N_13096,N_11084,N_11496);
nor U13097 (N_13097,N_11829,N_11701);
nand U13098 (N_13098,N_11408,N_11313);
and U13099 (N_13099,N_10908,N_10538);
and U13100 (N_13100,N_11303,N_11776);
and U13101 (N_13101,N_10566,N_10533);
nand U13102 (N_13102,N_11864,N_10805);
xor U13103 (N_13103,N_11159,N_11751);
or U13104 (N_13104,N_10735,N_11428);
or U13105 (N_13105,N_11027,N_10854);
xnor U13106 (N_13106,N_11070,N_10547);
xnor U13107 (N_13107,N_11518,N_11747);
nor U13108 (N_13108,N_10579,N_11618);
nor U13109 (N_13109,N_10578,N_10702);
nor U13110 (N_13110,N_10970,N_11023);
nand U13111 (N_13111,N_10815,N_11117);
xor U13112 (N_13112,N_11360,N_11576);
and U13113 (N_13113,N_10878,N_11956);
nor U13114 (N_13114,N_10637,N_10558);
xnor U13115 (N_13115,N_11144,N_11106);
xor U13116 (N_13116,N_11080,N_11608);
xnor U13117 (N_13117,N_11234,N_10627);
nand U13118 (N_13118,N_11172,N_11461);
or U13119 (N_13119,N_11536,N_11223);
nand U13120 (N_13120,N_10951,N_10993);
and U13121 (N_13121,N_11301,N_11492);
nor U13122 (N_13122,N_11268,N_10772);
or U13123 (N_13123,N_11096,N_11127);
nand U13124 (N_13124,N_10625,N_11101);
nand U13125 (N_13125,N_10638,N_11146);
xnor U13126 (N_13126,N_11339,N_11966);
and U13127 (N_13127,N_11116,N_11185);
nand U13128 (N_13128,N_10831,N_11760);
and U13129 (N_13129,N_10654,N_10851);
xnor U13130 (N_13130,N_11334,N_11723);
or U13131 (N_13131,N_11457,N_11757);
xnor U13132 (N_13132,N_11459,N_11913);
nand U13133 (N_13133,N_11589,N_11793);
nand U13134 (N_13134,N_11188,N_11550);
or U13135 (N_13135,N_11749,N_11238);
or U13136 (N_13136,N_11427,N_10607);
xor U13137 (N_13137,N_11699,N_10698);
xnor U13138 (N_13138,N_11099,N_11506);
or U13139 (N_13139,N_11004,N_11806);
nand U13140 (N_13140,N_11115,N_11988);
xor U13141 (N_13141,N_10652,N_10537);
or U13142 (N_13142,N_10616,N_11550);
and U13143 (N_13143,N_11562,N_11248);
nor U13144 (N_13144,N_11958,N_11424);
and U13145 (N_13145,N_11150,N_11417);
xnor U13146 (N_13146,N_11614,N_10509);
and U13147 (N_13147,N_10633,N_10722);
or U13148 (N_13148,N_10732,N_10919);
xnor U13149 (N_13149,N_11493,N_10533);
nor U13150 (N_13150,N_11857,N_11676);
or U13151 (N_13151,N_11842,N_11483);
and U13152 (N_13152,N_11010,N_11792);
or U13153 (N_13153,N_11713,N_11769);
nand U13154 (N_13154,N_10765,N_10794);
or U13155 (N_13155,N_11336,N_11589);
or U13156 (N_13156,N_11785,N_11043);
nand U13157 (N_13157,N_11663,N_10718);
nor U13158 (N_13158,N_11555,N_11149);
nand U13159 (N_13159,N_11956,N_11351);
or U13160 (N_13160,N_11078,N_10826);
nor U13161 (N_13161,N_11361,N_10580);
or U13162 (N_13162,N_11047,N_11494);
xnor U13163 (N_13163,N_11298,N_10992);
and U13164 (N_13164,N_11718,N_11778);
nor U13165 (N_13165,N_11382,N_10845);
and U13166 (N_13166,N_11550,N_11065);
and U13167 (N_13167,N_10675,N_11868);
nor U13168 (N_13168,N_11264,N_10927);
nand U13169 (N_13169,N_11106,N_11786);
nor U13170 (N_13170,N_11688,N_10749);
nand U13171 (N_13171,N_11178,N_10694);
or U13172 (N_13172,N_10864,N_10515);
nor U13173 (N_13173,N_10621,N_10556);
nand U13174 (N_13174,N_10634,N_11973);
xnor U13175 (N_13175,N_11249,N_10965);
nand U13176 (N_13176,N_11049,N_11843);
and U13177 (N_13177,N_11230,N_10583);
xor U13178 (N_13178,N_11543,N_10648);
or U13179 (N_13179,N_11706,N_11157);
or U13180 (N_13180,N_11298,N_10950);
nor U13181 (N_13181,N_11557,N_11642);
or U13182 (N_13182,N_11442,N_10697);
xor U13183 (N_13183,N_11987,N_11038);
nor U13184 (N_13184,N_10614,N_11395);
or U13185 (N_13185,N_10986,N_10786);
nor U13186 (N_13186,N_11862,N_11258);
and U13187 (N_13187,N_10637,N_10583);
and U13188 (N_13188,N_11678,N_10520);
nand U13189 (N_13189,N_11402,N_11349);
nand U13190 (N_13190,N_11869,N_11523);
nor U13191 (N_13191,N_11132,N_10698);
and U13192 (N_13192,N_10831,N_10974);
or U13193 (N_13193,N_10988,N_10965);
or U13194 (N_13194,N_11649,N_11791);
nor U13195 (N_13195,N_11096,N_11695);
or U13196 (N_13196,N_11590,N_11547);
nand U13197 (N_13197,N_11821,N_11285);
or U13198 (N_13198,N_11902,N_11401);
nor U13199 (N_13199,N_11664,N_10865);
and U13200 (N_13200,N_11689,N_11437);
and U13201 (N_13201,N_10720,N_11305);
and U13202 (N_13202,N_11997,N_10561);
nand U13203 (N_13203,N_11588,N_11389);
nor U13204 (N_13204,N_11993,N_11330);
nand U13205 (N_13205,N_11362,N_11370);
nor U13206 (N_13206,N_11199,N_11398);
nand U13207 (N_13207,N_11331,N_11795);
nor U13208 (N_13208,N_11391,N_11442);
and U13209 (N_13209,N_11581,N_10699);
nand U13210 (N_13210,N_11395,N_11800);
nor U13211 (N_13211,N_11160,N_10523);
xnor U13212 (N_13212,N_11944,N_10620);
xor U13213 (N_13213,N_10836,N_11222);
nor U13214 (N_13214,N_11482,N_11204);
nand U13215 (N_13215,N_10742,N_10794);
nor U13216 (N_13216,N_11807,N_10759);
nand U13217 (N_13217,N_10982,N_11736);
nor U13218 (N_13218,N_11556,N_11241);
nand U13219 (N_13219,N_10873,N_11842);
nor U13220 (N_13220,N_10708,N_11948);
nand U13221 (N_13221,N_10934,N_10704);
nor U13222 (N_13222,N_11784,N_10931);
nor U13223 (N_13223,N_11210,N_11858);
nand U13224 (N_13224,N_11158,N_11047);
nor U13225 (N_13225,N_11562,N_11600);
xor U13226 (N_13226,N_10804,N_10890);
and U13227 (N_13227,N_10747,N_11657);
nand U13228 (N_13228,N_10811,N_11087);
and U13229 (N_13229,N_10670,N_10562);
nor U13230 (N_13230,N_11498,N_11461);
and U13231 (N_13231,N_11702,N_10646);
or U13232 (N_13232,N_11145,N_10661);
and U13233 (N_13233,N_11312,N_11644);
nand U13234 (N_13234,N_11485,N_11376);
nor U13235 (N_13235,N_10882,N_10533);
and U13236 (N_13236,N_11408,N_11660);
nand U13237 (N_13237,N_10719,N_11605);
nand U13238 (N_13238,N_11333,N_11234);
nand U13239 (N_13239,N_11601,N_10688);
nor U13240 (N_13240,N_10823,N_11008);
and U13241 (N_13241,N_11087,N_10874);
or U13242 (N_13242,N_10879,N_10911);
and U13243 (N_13243,N_11125,N_10909);
nand U13244 (N_13244,N_11078,N_11992);
or U13245 (N_13245,N_10537,N_11026);
nor U13246 (N_13246,N_11652,N_11154);
or U13247 (N_13247,N_10695,N_11633);
or U13248 (N_13248,N_10919,N_11236);
or U13249 (N_13249,N_11025,N_10744);
and U13250 (N_13250,N_11272,N_11002);
nand U13251 (N_13251,N_11442,N_11350);
and U13252 (N_13252,N_10582,N_11010);
xor U13253 (N_13253,N_11852,N_11954);
nor U13254 (N_13254,N_11733,N_11976);
nor U13255 (N_13255,N_11249,N_10845);
or U13256 (N_13256,N_11795,N_11647);
or U13257 (N_13257,N_11236,N_11524);
nand U13258 (N_13258,N_11666,N_11149);
and U13259 (N_13259,N_10853,N_11729);
and U13260 (N_13260,N_10737,N_10608);
or U13261 (N_13261,N_11736,N_10727);
nor U13262 (N_13262,N_11493,N_10826);
nand U13263 (N_13263,N_11995,N_10710);
nor U13264 (N_13264,N_11072,N_11628);
nor U13265 (N_13265,N_11017,N_10770);
and U13266 (N_13266,N_11206,N_11513);
nand U13267 (N_13267,N_11467,N_11119);
nand U13268 (N_13268,N_10904,N_10868);
or U13269 (N_13269,N_10813,N_10901);
nand U13270 (N_13270,N_11275,N_11882);
or U13271 (N_13271,N_11604,N_11448);
xor U13272 (N_13272,N_11089,N_10738);
or U13273 (N_13273,N_11592,N_11816);
nor U13274 (N_13274,N_11360,N_10798);
xnor U13275 (N_13275,N_11683,N_11209);
nor U13276 (N_13276,N_10714,N_10632);
nor U13277 (N_13277,N_11087,N_11502);
nor U13278 (N_13278,N_11899,N_11767);
nor U13279 (N_13279,N_10549,N_11531);
and U13280 (N_13280,N_11676,N_11443);
nor U13281 (N_13281,N_10815,N_11781);
nand U13282 (N_13282,N_11866,N_11003);
or U13283 (N_13283,N_10627,N_11645);
and U13284 (N_13284,N_11773,N_11706);
nor U13285 (N_13285,N_11953,N_11308);
nor U13286 (N_13286,N_11833,N_10869);
and U13287 (N_13287,N_11901,N_11479);
or U13288 (N_13288,N_11352,N_11584);
and U13289 (N_13289,N_11184,N_10867);
nor U13290 (N_13290,N_11046,N_11929);
nand U13291 (N_13291,N_10500,N_10945);
and U13292 (N_13292,N_11750,N_10696);
and U13293 (N_13293,N_11086,N_11642);
or U13294 (N_13294,N_11804,N_11908);
nand U13295 (N_13295,N_11319,N_11246);
nor U13296 (N_13296,N_11923,N_11848);
and U13297 (N_13297,N_11525,N_11498);
nand U13298 (N_13298,N_11396,N_11656);
or U13299 (N_13299,N_10944,N_11045);
nor U13300 (N_13300,N_10652,N_11143);
or U13301 (N_13301,N_11150,N_10952);
or U13302 (N_13302,N_11449,N_11214);
nor U13303 (N_13303,N_11452,N_11352);
nor U13304 (N_13304,N_10695,N_11553);
and U13305 (N_13305,N_10759,N_11462);
and U13306 (N_13306,N_10939,N_11443);
and U13307 (N_13307,N_10711,N_10870);
nand U13308 (N_13308,N_10819,N_11286);
nand U13309 (N_13309,N_11223,N_10842);
and U13310 (N_13310,N_11435,N_10899);
nand U13311 (N_13311,N_11948,N_11190);
or U13312 (N_13312,N_10660,N_10555);
nor U13313 (N_13313,N_11565,N_11274);
or U13314 (N_13314,N_11763,N_10634);
xor U13315 (N_13315,N_11020,N_11778);
or U13316 (N_13316,N_11536,N_11711);
and U13317 (N_13317,N_11250,N_10673);
nor U13318 (N_13318,N_11340,N_11125);
nor U13319 (N_13319,N_11784,N_11337);
and U13320 (N_13320,N_11217,N_11354);
and U13321 (N_13321,N_10716,N_10695);
nand U13322 (N_13322,N_11780,N_11351);
or U13323 (N_13323,N_10569,N_11458);
and U13324 (N_13324,N_10685,N_11369);
nor U13325 (N_13325,N_10534,N_11104);
xnor U13326 (N_13326,N_11910,N_11222);
nor U13327 (N_13327,N_11364,N_11592);
nor U13328 (N_13328,N_10691,N_11634);
xnor U13329 (N_13329,N_11354,N_11022);
or U13330 (N_13330,N_11024,N_11569);
or U13331 (N_13331,N_10600,N_10584);
and U13332 (N_13332,N_10826,N_10650);
xnor U13333 (N_13333,N_11784,N_10922);
or U13334 (N_13334,N_10955,N_11090);
nor U13335 (N_13335,N_10829,N_11972);
nor U13336 (N_13336,N_11082,N_10950);
and U13337 (N_13337,N_10688,N_11567);
nand U13338 (N_13338,N_10565,N_10829);
nand U13339 (N_13339,N_11157,N_11469);
and U13340 (N_13340,N_11237,N_10917);
nand U13341 (N_13341,N_11756,N_10981);
and U13342 (N_13342,N_10706,N_11306);
nand U13343 (N_13343,N_11330,N_11389);
or U13344 (N_13344,N_11942,N_10501);
or U13345 (N_13345,N_11782,N_11037);
nand U13346 (N_13346,N_11543,N_11169);
nor U13347 (N_13347,N_10979,N_10816);
or U13348 (N_13348,N_11446,N_11005);
or U13349 (N_13349,N_11212,N_10784);
xnor U13350 (N_13350,N_10820,N_10706);
and U13351 (N_13351,N_10913,N_10567);
and U13352 (N_13352,N_11150,N_11178);
nor U13353 (N_13353,N_11850,N_11014);
and U13354 (N_13354,N_11821,N_11928);
and U13355 (N_13355,N_11606,N_11477);
nor U13356 (N_13356,N_11165,N_11063);
nand U13357 (N_13357,N_11237,N_11543);
nand U13358 (N_13358,N_11301,N_11733);
and U13359 (N_13359,N_10965,N_11974);
nand U13360 (N_13360,N_11526,N_11578);
or U13361 (N_13361,N_11983,N_11745);
nor U13362 (N_13362,N_11690,N_11535);
nor U13363 (N_13363,N_10925,N_10577);
or U13364 (N_13364,N_10845,N_10611);
nand U13365 (N_13365,N_11203,N_11137);
or U13366 (N_13366,N_11172,N_11274);
and U13367 (N_13367,N_11220,N_11307);
nand U13368 (N_13368,N_11090,N_10902);
or U13369 (N_13369,N_10561,N_10942);
nor U13370 (N_13370,N_10611,N_11400);
and U13371 (N_13371,N_11343,N_11546);
nand U13372 (N_13372,N_11917,N_10947);
nor U13373 (N_13373,N_11569,N_11129);
nand U13374 (N_13374,N_11493,N_11220);
and U13375 (N_13375,N_10546,N_10529);
nand U13376 (N_13376,N_11516,N_10806);
nand U13377 (N_13377,N_11824,N_10545);
xor U13378 (N_13378,N_11075,N_10604);
and U13379 (N_13379,N_11760,N_11333);
or U13380 (N_13380,N_10917,N_11183);
and U13381 (N_13381,N_10873,N_11695);
nor U13382 (N_13382,N_11534,N_10945);
or U13383 (N_13383,N_10800,N_11298);
nand U13384 (N_13384,N_10646,N_10634);
nor U13385 (N_13385,N_11817,N_10657);
nand U13386 (N_13386,N_10533,N_11819);
nand U13387 (N_13387,N_11459,N_10608);
or U13388 (N_13388,N_11090,N_11212);
and U13389 (N_13389,N_11213,N_11704);
nor U13390 (N_13390,N_10540,N_10500);
or U13391 (N_13391,N_10987,N_11347);
or U13392 (N_13392,N_11878,N_11595);
or U13393 (N_13393,N_10909,N_10652);
nand U13394 (N_13394,N_10643,N_10691);
and U13395 (N_13395,N_10791,N_11646);
xor U13396 (N_13396,N_11270,N_11196);
and U13397 (N_13397,N_11132,N_11696);
nor U13398 (N_13398,N_10523,N_11995);
and U13399 (N_13399,N_11828,N_11307);
nand U13400 (N_13400,N_11081,N_11236);
nand U13401 (N_13401,N_10920,N_10815);
and U13402 (N_13402,N_11764,N_11990);
nand U13403 (N_13403,N_11483,N_10652);
and U13404 (N_13404,N_10703,N_11824);
or U13405 (N_13405,N_10827,N_10924);
and U13406 (N_13406,N_11828,N_11663);
nor U13407 (N_13407,N_11148,N_10666);
nor U13408 (N_13408,N_10922,N_11977);
nor U13409 (N_13409,N_11901,N_11162);
and U13410 (N_13410,N_11515,N_10570);
nor U13411 (N_13411,N_11456,N_11051);
nor U13412 (N_13412,N_11517,N_11232);
or U13413 (N_13413,N_10750,N_11251);
or U13414 (N_13414,N_10841,N_10897);
nor U13415 (N_13415,N_10572,N_10520);
and U13416 (N_13416,N_11155,N_10606);
nor U13417 (N_13417,N_11893,N_10951);
and U13418 (N_13418,N_11178,N_11890);
nor U13419 (N_13419,N_10573,N_10740);
nand U13420 (N_13420,N_10672,N_11432);
and U13421 (N_13421,N_11247,N_11458);
nand U13422 (N_13422,N_11294,N_10895);
and U13423 (N_13423,N_10756,N_11269);
or U13424 (N_13424,N_11116,N_11141);
and U13425 (N_13425,N_11559,N_10679);
or U13426 (N_13426,N_11587,N_10627);
nor U13427 (N_13427,N_10631,N_10822);
and U13428 (N_13428,N_11694,N_11301);
xnor U13429 (N_13429,N_11457,N_10616);
nand U13430 (N_13430,N_11069,N_10746);
and U13431 (N_13431,N_10816,N_10732);
nand U13432 (N_13432,N_11027,N_11091);
nor U13433 (N_13433,N_11966,N_10611);
and U13434 (N_13434,N_11212,N_11271);
or U13435 (N_13435,N_11143,N_11582);
nand U13436 (N_13436,N_10987,N_11826);
nand U13437 (N_13437,N_11258,N_11729);
nor U13438 (N_13438,N_10566,N_10929);
nand U13439 (N_13439,N_11129,N_11015);
nand U13440 (N_13440,N_10616,N_11675);
nor U13441 (N_13441,N_11046,N_11719);
xnor U13442 (N_13442,N_10538,N_11527);
nand U13443 (N_13443,N_11454,N_10986);
or U13444 (N_13444,N_11075,N_11717);
nor U13445 (N_13445,N_11465,N_11529);
or U13446 (N_13446,N_11388,N_11634);
nand U13447 (N_13447,N_10649,N_11766);
and U13448 (N_13448,N_10954,N_11618);
nor U13449 (N_13449,N_11016,N_11490);
xor U13450 (N_13450,N_11488,N_10973);
nor U13451 (N_13451,N_10501,N_10781);
nand U13452 (N_13452,N_11119,N_11209);
or U13453 (N_13453,N_11005,N_11884);
nand U13454 (N_13454,N_11163,N_11139);
or U13455 (N_13455,N_11168,N_10553);
nor U13456 (N_13456,N_11905,N_10942);
nand U13457 (N_13457,N_10833,N_11217);
or U13458 (N_13458,N_10846,N_11074);
nor U13459 (N_13459,N_11371,N_10974);
nor U13460 (N_13460,N_11718,N_11044);
nor U13461 (N_13461,N_11357,N_10533);
nand U13462 (N_13462,N_11319,N_10779);
nor U13463 (N_13463,N_11190,N_11208);
and U13464 (N_13464,N_11377,N_11086);
nor U13465 (N_13465,N_11122,N_11379);
or U13466 (N_13466,N_11462,N_10596);
nor U13467 (N_13467,N_10945,N_11624);
nand U13468 (N_13468,N_11909,N_10577);
nand U13469 (N_13469,N_10635,N_11759);
or U13470 (N_13470,N_11440,N_11352);
nand U13471 (N_13471,N_11427,N_11367);
xor U13472 (N_13472,N_11881,N_11196);
nor U13473 (N_13473,N_10666,N_11567);
nor U13474 (N_13474,N_11922,N_11804);
or U13475 (N_13475,N_11177,N_10578);
and U13476 (N_13476,N_11933,N_10880);
nor U13477 (N_13477,N_11551,N_10611);
and U13478 (N_13478,N_10537,N_11973);
nor U13479 (N_13479,N_11248,N_10732);
xor U13480 (N_13480,N_11931,N_11128);
nor U13481 (N_13481,N_11039,N_11959);
or U13482 (N_13482,N_11134,N_10812);
and U13483 (N_13483,N_10754,N_11284);
nand U13484 (N_13484,N_11799,N_10744);
or U13485 (N_13485,N_11859,N_11697);
or U13486 (N_13486,N_10770,N_10999);
nor U13487 (N_13487,N_11954,N_11810);
nand U13488 (N_13488,N_11974,N_10651);
or U13489 (N_13489,N_11904,N_11506);
nor U13490 (N_13490,N_11851,N_11279);
and U13491 (N_13491,N_10923,N_11024);
xnor U13492 (N_13492,N_11363,N_11654);
or U13493 (N_13493,N_10581,N_11707);
xor U13494 (N_13494,N_11480,N_11347);
nand U13495 (N_13495,N_11340,N_11643);
and U13496 (N_13496,N_11412,N_11510);
xnor U13497 (N_13497,N_10778,N_11592);
xor U13498 (N_13498,N_10773,N_10832);
nor U13499 (N_13499,N_11974,N_11117);
and U13500 (N_13500,N_13159,N_12511);
or U13501 (N_13501,N_12243,N_12110);
nand U13502 (N_13502,N_12076,N_12093);
nand U13503 (N_13503,N_13298,N_13343);
or U13504 (N_13504,N_12703,N_12995);
and U13505 (N_13505,N_13193,N_12289);
nor U13506 (N_13506,N_13339,N_12860);
and U13507 (N_13507,N_13313,N_12250);
nand U13508 (N_13508,N_13172,N_12214);
and U13509 (N_13509,N_12652,N_12442);
and U13510 (N_13510,N_12936,N_12976);
nor U13511 (N_13511,N_12241,N_12213);
and U13512 (N_13512,N_12272,N_13405);
xnor U13513 (N_13513,N_12819,N_12406);
nand U13514 (N_13514,N_13088,N_12147);
xnor U13515 (N_13515,N_12799,N_12464);
or U13516 (N_13516,N_13336,N_12552);
nor U13517 (N_13517,N_13455,N_12154);
nand U13518 (N_13518,N_12744,N_13457);
xnor U13519 (N_13519,N_12704,N_12440);
or U13520 (N_13520,N_13074,N_12475);
nor U13521 (N_13521,N_12596,N_12750);
nor U13522 (N_13522,N_13224,N_12606);
or U13523 (N_13523,N_12179,N_12875);
nor U13524 (N_13524,N_12638,N_12074);
nor U13525 (N_13525,N_13425,N_12623);
nor U13526 (N_13526,N_12062,N_12259);
nand U13527 (N_13527,N_12070,N_12222);
nor U13528 (N_13528,N_13129,N_12726);
nand U13529 (N_13529,N_12317,N_13024);
nand U13530 (N_13530,N_12348,N_13247);
nand U13531 (N_13531,N_12314,N_12457);
or U13532 (N_13532,N_12201,N_12480);
and U13533 (N_13533,N_12956,N_13165);
and U13534 (N_13534,N_12021,N_13104);
and U13535 (N_13535,N_13188,N_12275);
or U13536 (N_13536,N_12391,N_13005);
and U13537 (N_13537,N_12692,N_13107);
nand U13538 (N_13538,N_12741,N_12673);
nand U13539 (N_13539,N_12544,N_12683);
xnor U13540 (N_13540,N_12519,N_12612);
nor U13541 (N_13541,N_12411,N_12530);
nor U13542 (N_13542,N_13393,N_12418);
nand U13543 (N_13543,N_13387,N_13401);
and U13544 (N_13544,N_12835,N_13306);
or U13545 (N_13545,N_12791,N_13227);
or U13546 (N_13546,N_12928,N_12727);
and U13547 (N_13547,N_13178,N_12965);
xnor U13548 (N_13548,N_13469,N_13491);
or U13549 (N_13549,N_12907,N_12264);
nor U13550 (N_13550,N_13284,N_13004);
or U13551 (N_13551,N_12472,N_13158);
or U13552 (N_13552,N_13181,N_12378);
or U13553 (N_13553,N_13060,N_12576);
nor U13554 (N_13554,N_13324,N_12695);
and U13555 (N_13555,N_13090,N_13430);
or U13556 (N_13556,N_12631,N_13108);
nor U13557 (N_13557,N_12112,N_13226);
nand U13558 (N_13558,N_13128,N_12587);
or U13559 (N_13559,N_12651,N_13127);
or U13560 (N_13560,N_12253,N_12583);
and U13561 (N_13561,N_12063,N_12495);
and U13562 (N_13562,N_12034,N_12790);
or U13563 (N_13563,N_12292,N_12582);
nand U13564 (N_13564,N_13382,N_12877);
nor U13565 (N_13565,N_12142,N_12352);
and U13566 (N_13566,N_12882,N_12124);
nor U13567 (N_13567,N_13283,N_13293);
nand U13568 (N_13568,N_12466,N_12251);
nor U13569 (N_13569,N_12434,N_12861);
nor U13570 (N_13570,N_12917,N_13134);
nand U13571 (N_13571,N_12771,N_13021);
xnor U13572 (N_13572,N_13275,N_13039);
or U13573 (N_13573,N_13274,N_12891);
nand U13574 (N_13574,N_13453,N_12156);
nor U13575 (N_13575,N_12979,N_13404);
or U13576 (N_13576,N_13092,N_13011);
and U13577 (N_13577,N_13078,N_12349);
nor U13578 (N_13578,N_12007,N_12820);
and U13579 (N_13579,N_12479,N_12113);
or U13580 (N_13580,N_12534,N_12992);
and U13581 (N_13581,N_12354,N_12551);
nand U13582 (N_13582,N_12166,N_12721);
and U13583 (N_13583,N_12211,N_12117);
nand U13584 (N_13584,N_12944,N_13244);
nor U13585 (N_13585,N_12102,N_12746);
nor U13586 (N_13586,N_13157,N_13144);
or U13587 (N_13587,N_12485,N_12061);
or U13588 (N_13588,N_12850,N_12796);
or U13589 (N_13589,N_12384,N_12344);
and U13590 (N_13590,N_13229,N_13136);
or U13591 (N_13591,N_13034,N_12417);
xor U13592 (N_13592,N_12058,N_12219);
xor U13593 (N_13593,N_13190,N_13235);
or U13594 (N_13594,N_13103,N_12924);
nor U13595 (N_13595,N_12316,N_13186);
and U13596 (N_13596,N_12290,N_12018);
nand U13597 (N_13597,N_12421,N_12772);
nand U13598 (N_13598,N_12679,N_12180);
and U13599 (N_13599,N_12300,N_12035);
or U13600 (N_13600,N_12953,N_13036);
nor U13601 (N_13601,N_12604,N_12634);
or U13602 (N_13602,N_12616,N_13305);
or U13603 (N_13603,N_12257,N_12223);
nor U13604 (N_13604,N_12911,N_12724);
or U13605 (N_13605,N_13413,N_13041);
nand U13606 (N_13606,N_13345,N_12240);
nand U13607 (N_13607,N_13361,N_12000);
nor U13608 (N_13608,N_12015,N_12937);
nor U13609 (N_13609,N_12846,N_12165);
or U13610 (N_13610,N_12635,N_13485);
nor U13611 (N_13611,N_13400,N_12561);
xor U13612 (N_13612,N_12342,N_12330);
and U13613 (N_13613,N_12297,N_12146);
and U13614 (N_13614,N_12786,N_12873);
nand U13615 (N_13615,N_13403,N_12952);
xnor U13616 (N_13616,N_13046,N_12644);
and U13617 (N_13617,N_13091,N_13206);
nand U13618 (N_13618,N_13102,N_12218);
nand U13619 (N_13619,N_12263,N_12256);
and U13620 (N_13620,N_12362,N_13061);
or U13621 (N_13621,N_13198,N_13000);
nand U13622 (N_13622,N_12014,N_12525);
xnor U13623 (N_13623,N_12068,N_13473);
and U13624 (N_13624,N_12700,N_13341);
and U13625 (N_13625,N_12915,N_12232);
nor U13626 (N_13626,N_13049,N_13105);
or U13627 (N_13627,N_12709,N_12153);
xnor U13628 (N_13628,N_12131,N_12887);
nor U13629 (N_13629,N_13292,N_12880);
nand U13630 (N_13630,N_12826,N_12688);
nor U13631 (N_13631,N_13213,N_13205);
and U13632 (N_13632,N_12513,N_13223);
or U13633 (N_13633,N_13474,N_13208);
and U13634 (N_13634,N_12105,N_12867);
xnor U13635 (N_13635,N_12611,N_12728);
or U13636 (N_13636,N_12900,N_13154);
xor U13637 (N_13637,N_12716,N_12801);
and U13638 (N_13638,N_12975,N_12041);
nor U13639 (N_13639,N_13335,N_12702);
nand U13640 (N_13640,N_12234,N_12533);
nand U13641 (N_13641,N_12027,N_13201);
or U13642 (N_13642,N_12636,N_13492);
and U13643 (N_13643,N_12556,N_13360);
nor U13644 (N_13644,N_12617,N_12026);
and U13645 (N_13645,N_13266,N_13267);
or U13646 (N_13646,N_12224,N_13347);
nand U13647 (N_13647,N_12627,N_12849);
or U13648 (N_13648,N_12870,N_12394);
nor U13649 (N_13649,N_12422,N_12987);
and U13650 (N_13650,N_12336,N_12357);
or U13651 (N_13651,N_12591,N_13412);
and U13652 (N_13652,N_13318,N_13254);
and U13653 (N_13653,N_13315,N_13338);
nand U13654 (N_13654,N_12005,N_13153);
nor U13655 (N_13655,N_12751,N_13307);
and U13656 (N_13656,N_13197,N_13427);
nand U13657 (N_13657,N_12568,N_13019);
nor U13658 (N_13658,N_13076,N_13101);
nand U13659 (N_13659,N_12456,N_12413);
nand U13660 (N_13660,N_12549,N_12307);
nor U13661 (N_13661,N_12514,N_12176);
nor U13662 (N_13662,N_12712,N_12523);
nor U13663 (N_13663,N_12925,N_13013);
or U13664 (N_13664,N_12660,N_13278);
nand U13665 (N_13665,N_13351,N_12152);
nand U13666 (N_13666,N_13189,N_12943);
and U13667 (N_13667,N_13332,N_12960);
nand U13668 (N_13668,N_12686,N_12444);
nor U13669 (N_13669,N_12756,N_13058);
and U13670 (N_13670,N_13482,N_12586);
nor U13671 (N_13671,N_12040,N_13467);
or U13672 (N_13672,N_12198,N_13383);
or U13673 (N_13673,N_12051,N_13409);
nand U13674 (N_13674,N_13431,N_12524);
nand U13675 (N_13675,N_12844,N_12809);
or U13676 (N_13676,N_12607,N_13433);
nand U13677 (N_13677,N_12705,N_12518);
and U13678 (N_13678,N_12023,N_12984);
or U13679 (N_13679,N_13449,N_12885);
and U13680 (N_13680,N_12642,N_12004);
nor U13681 (N_13681,N_12465,N_13045);
and U13682 (N_13682,N_12935,N_13321);
nand U13683 (N_13683,N_12811,N_13269);
xnor U13684 (N_13684,N_13029,N_13312);
nand U13685 (N_13685,N_12983,N_12516);
or U13686 (N_13686,N_13211,N_12424);
xor U13687 (N_13687,N_13248,N_12496);
and U13688 (N_13688,N_12575,N_13150);
nand U13689 (N_13689,N_13459,N_13073);
nand U13690 (N_13690,N_12939,N_13083);
nand U13691 (N_13691,N_13466,N_12914);
and U13692 (N_13692,N_12333,N_12589);
nand U13693 (N_13693,N_12077,N_12087);
and U13694 (N_13694,N_12547,N_13255);
or U13695 (N_13695,N_13263,N_12399);
nand U13696 (N_13696,N_12507,N_13456);
or U13697 (N_13697,N_12904,N_12294);
and U13698 (N_13698,N_13007,N_12206);
nand U13699 (N_13699,N_12581,N_12610);
and U13700 (N_13700,N_12505,N_13098);
and U13701 (N_13701,N_13030,N_13216);
nor U13702 (N_13702,N_13418,N_13426);
nor U13703 (N_13703,N_13288,N_12557);
or U13704 (N_13704,N_12743,N_12654);
nor U13705 (N_13705,N_12940,N_13286);
nand U13706 (N_13706,N_12609,N_12392);
nor U13707 (N_13707,N_12386,N_12404);
or U13708 (N_13708,N_13033,N_13017);
and U13709 (N_13709,N_12816,N_12228);
or U13710 (N_13710,N_12193,N_13122);
or U13711 (N_13711,N_13093,N_12010);
nand U13712 (N_13712,N_12186,N_12590);
nand U13713 (N_13713,N_12753,N_12655);
nor U13714 (N_13714,N_12141,N_12571);
nor U13715 (N_13715,N_12455,N_13233);
and U13716 (N_13716,N_12210,N_12452);
nand U13717 (N_13717,N_12615,N_12208);
nor U13718 (N_13718,N_13204,N_12050);
or U13719 (N_13719,N_12020,N_13446);
nand U13720 (N_13720,N_13421,N_12526);
and U13721 (N_13721,N_13348,N_13450);
or U13722 (N_13722,N_12433,N_12269);
or U13723 (N_13723,N_13243,N_13121);
xor U13724 (N_13724,N_12787,N_12379);
and U13725 (N_13725,N_12215,N_12510);
or U13726 (N_13726,N_13476,N_12310);
nor U13727 (N_13727,N_13297,N_12934);
xnor U13728 (N_13728,N_13225,N_12578);
nand U13729 (N_13729,N_12874,N_12028);
xnor U13730 (N_13730,N_13494,N_12429);
nand U13731 (N_13731,N_12947,N_13008);
and U13732 (N_13732,N_13327,N_12948);
nand U13733 (N_13733,N_13068,N_13316);
nor U13734 (N_13734,N_12056,N_12871);
or U13735 (N_13735,N_12980,N_12012);
or U13736 (N_13736,N_13215,N_13020);
and U13737 (N_13737,N_13023,N_12780);
nor U13738 (N_13738,N_13042,N_13027);
nor U13739 (N_13739,N_12868,N_12419);
and U13740 (N_13740,N_12149,N_12381);
and U13741 (N_13741,N_12200,N_12287);
and U13742 (N_13742,N_12319,N_12897);
and U13743 (N_13743,N_12374,N_12098);
nand U13744 (N_13744,N_12912,N_12489);
and U13745 (N_13745,N_12121,N_12360);
and U13746 (N_13746,N_12343,N_12527);
or U13747 (N_13747,N_12955,N_12395);
and U13748 (N_13748,N_12420,N_12710);
and U13749 (N_13749,N_12967,N_12311);
nand U13750 (N_13750,N_12921,N_12991);
or U13751 (N_13751,N_12950,N_12192);
xnor U13752 (N_13752,N_13424,N_12650);
xnor U13753 (N_13753,N_12260,N_12331);
or U13754 (N_13754,N_12656,N_13370);
or U13755 (N_13755,N_13423,N_12235);
and U13756 (N_13756,N_12091,N_12385);
nor U13757 (N_13757,N_12299,N_12559);
nor U13758 (N_13758,N_12630,N_12126);
or U13759 (N_13759,N_12713,N_13463);
or U13760 (N_13760,N_12601,N_12225);
nor U13761 (N_13761,N_12963,N_13142);
nand U13762 (N_13762,N_13419,N_12069);
or U13763 (N_13763,N_12347,N_12680);
or U13764 (N_13764,N_12388,N_13493);
or U13765 (N_13765,N_12337,N_13460);
and U13766 (N_13766,N_12593,N_12238);
xnor U13767 (N_13767,N_12371,N_12261);
and U13768 (N_13768,N_13143,N_12500);
nor U13769 (N_13769,N_12375,N_13200);
nand U13770 (N_13770,N_13296,N_12504);
and U13771 (N_13771,N_12558,N_12775);
or U13772 (N_13772,N_12645,N_12770);
nor U13773 (N_13773,N_12339,N_12689);
nor U13774 (N_13774,N_12351,N_12229);
or U13775 (N_13775,N_12542,N_12158);
and U13776 (N_13776,N_12431,N_12376);
nor U13777 (N_13777,N_13119,N_12461);
xor U13778 (N_13778,N_12338,N_13116);
xnor U13779 (N_13779,N_12067,N_12132);
nor U13780 (N_13780,N_12084,N_13125);
nor U13781 (N_13781,N_12566,N_12451);
and U13782 (N_13782,N_12435,N_12691);
nor U13783 (N_13783,N_12818,N_13210);
or U13784 (N_13784,N_12535,N_12807);
nand U13785 (N_13785,N_13272,N_12450);
or U13786 (N_13786,N_13228,N_12964);
nand U13787 (N_13787,N_12862,N_12671);
or U13788 (N_13788,N_13322,N_12033);
or U13789 (N_13789,N_13395,N_13112);
nor U13790 (N_13790,N_13171,N_12237);
nand U13791 (N_13791,N_13349,N_12090);
and U13792 (N_13792,N_13477,N_12739);
or U13793 (N_13793,N_12555,N_13065);
nor U13794 (N_13794,N_12531,N_12829);
and U13795 (N_13795,N_13289,N_12390);
or U13796 (N_13796,N_12782,N_12170);
nand U13797 (N_13797,N_12988,N_13451);
or U13798 (N_13798,N_12373,N_12893);
nand U13799 (N_13799,N_12094,N_12400);
nand U13800 (N_13800,N_12150,N_13319);
xnor U13801 (N_13801,N_12055,N_13059);
and U13802 (N_13802,N_12764,N_12478);
nor U13803 (N_13803,N_13429,N_12682);
or U13804 (N_13804,N_12426,N_13110);
nand U13805 (N_13805,N_13145,N_12993);
nand U13806 (N_13806,N_12412,N_12878);
nor U13807 (N_13807,N_12060,N_12143);
nor U13808 (N_13808,N_12151,N_12605);
and U13809 (N_13809,N_12048,N_12570);
nor U13810 (N_13810,N_12959,N_12493);
and U13811 (N_13811,N_12127,N_12247);
nor U13812 (N_13812,N_12827,N_12720);
nor U13813 (N_13813,N_12546,N_12291);
and U13814 (N_13814,N_12301,N_13337);
nand U13815 (N_13815,N_13089,N_12437);
and U13816 (N_13816,N_13245,N_12477);
and U13817 (N_13817,N_12066,N_13135);
nor U13818 (N_13818,N_12296,N_12639);
and U13819 (N_13819,N_12101,N_13040);
nand U13820 (N_13820,N_12997,N_13246);
nor U13821 (N_13821,N_13120,N_12580);
nor U13822 (N_13822,N_12252,N_12288);
and U13823 (N_13823,N_12509,N_12996);
or U13824 (N_13824,N_13070,N_12136);
or U13825 (N_13825,N_13238,N_12830);
or U13826 (N_13826,N_12646,N_12502);
nand U13827 (N_13827,N_13362,N_12793);
or U13828 (N_13828,N_12031,N_12614);
or U13829 (N_13829,N_13115,N_13375);
or U13830 (N_13830,N_12981,N_13014);
and U13831 (N_13831,N_12968,N_12841);
and U13832 (N_13832,N_13420,N_13131);
nor U13833 (N_13833,N_13356,N_12777);
nand U13834 (N_13834,N_12476,N_12163);
or U13835 (N_13835,N_12664,N_13050);
or U13836 (N_13836,N_12410,N_12930);
or U13837 (N_13837,N_12595,N_13432);
or U13838 (N_13838,N_13468,N_13086);
and U13839 (N_13839,N_12189,N_12608);
nand U13840 (N_13840,N_12554,N_12160);
or U13841 (N_13841,N_13117,N_13152);
nor U13842 (N_13842,N_12115,N_12054);
and U13843 (N_13843,N_13273,N_12487);
or U13844 (N_13844,N_12017,N_12254);
xnor U13845 (N_13845,N_12078,N_13082);
nand U13846 (N_13846,N_12961,N_12765);
and U13847 (N_13847,N_12541,N_12231);
or U13848 (N_13848,N_13176,N_13488);
nor U13849 (N_13849,N_12266,N_12107);
nand U13850 (N_13850,N_12798,N_12926);
nand U13851 (N_13851,N_13410,N_12008);
and U13852 (N_13852,N_12239,N_12072);
and U13853 (N_13853,N_13416,N_12405);
xnor U13854 (N_13854,N_12800,N_12633);
and U13855 (N_13855,N_12574,N_13350);
and U13856 (N_13856,N_13422,N_12207);
xor U13857 (N_13857,N_13138,N_12203);
nor U13858 (N_13858,N_12693,N_12738);
and U13859 (N_13859,N_12687,N_12506);
and U13860 (N_13860,N_12220,N_12903);
nand U13861 (N_13861,N_12209,N_13282);
nand U13862 (N_13862,N_13130,N_13016);
and U13863 (N_13863,N_12825,N_12503);
nand U13864 (N_13864,N_13397,N_12856);
xnor U13865 (N_13865,N_13028,N_13271);
and U13866 (N_13866,N_12366,N_12803);
or U13867 (N_13867,N_12842,N_12889);
nor U13868 (N_13868,N_13114,N_12640);
nor U13869 (N_13869,N_12082,N_12064);
nand U13870 (N_13870,N_12677,N_12363);
xor U13871 (N_13871,N_13195,N_13085);
or U13872 (N_13872,N_13399,N_13465);
nor U13873 (N_13873,N_12145,N_13192);
nor U13874 (N_13874,N_12895,N_12923);
or U13875 (N_13875,N_12119,N_12901);
nand U13876 (N_13876,N_13163,N_13378);
nor U13877 (N_13877,N_12872,N_13231);
nor U13878 (N_13878,N_13380,N_13148);
or U13879 (N_13879,N_13003,N_12626);
nor U13880 (N_13880,N_12372,N_12382);
nand U13881 (N_13881,N_13290,N_12494);
xnor U13882 (N_13882,N_13408,N_12676);
or U13883 (N_13883,N_13471,N_12407);
nand U13884 (N_13884,N_13406,N_13072);
or U13885 (N_13885,N_12763,N_12217);
xnor U13886 (N_13886,N_12467,N_12364);
and U13887 (N_13887,N_13389,N_13268);
and U13888 (N_13888,N_12898,N_12075);
or U13889 (N_13889,N_13281,N_12945);
nand U13890 (N_13890,N_12236,N_12327);
and U13891 (N_13891,N_13483,N_13147);
or U13892 (N_13892,N_13212,N_12029);
or U13893 (N_13893,N_12579,N_12109);
or U13894 (N_13894,N_12760,N_12902);
nor U13895 (N_13895,N_13214,N_13140);
and U13896 (N_13896,N_12852,N_12757);
nand U13897 (N_13897,N_12468,N_13258);
nand U13898 (N_13898,N_12755,N_12804);
nand U13899 (N_13899,N_13084,N_13377);
or U13900 (N_13900,N_12168,N_13259);
or U13901 (N_13901,N_13006,N_12346);
nor U13902 (N_13902,N_12859,N_12335);
nor U13903 (N_13903,N_12309,N_12045);
xnor U13904 (N_13904,N_12318,N_13415);
nor U13905 (N_13905,N_12491,N_13295);
nand U13906 (N_13906,N_13166,N_12585);
and U13907 (N_13907,N_12255,N_12543);
nand U13908 (N_13908,N_12245,N_12740);
nor U13909 (N_13909,N_12308,N_12325);
nand U13910 (N_13910,N_12359,N_13484);
nor U13911 (N_13911,N_12563,N_13094);
and U13912 (N_13912,N_12032,N_12762);
nand U13913 (N_13913,N_13047,N_13454);
nand U13914 (N_13914,N_12661,N_12187);
nand U13915 (N_13915,N_12532,N_12624);
nor U13916 (N_13916,N_12280,N_12685);
or U13917 (N_13917,N_12813,N_13314);
nand U13918 (N_13918,N_12719,N_12792);
nor U13919 (N_13919,N_12037,N_12742);
nor U13920 (N_13920,N_12302,N_12171);
nor U13921 (N_13921,N_12324,N_12845);
nor U13922 (N_13922,N_12737,N_13390);
nand U13923 (N_13923,N_12182,N_12648);
nand U13924 (N_13924,N_12794,N_13280);
and U13925 (N_13925,N_12708,N_12512);
or U13926 (N_13926,N_13302,N_13264);
and U13927 (N_13927,N_12249,N_12175);
and U13928 (N_13928,N_12977,N_12003);
or U13929 (N_13929,N_12619,N_12722);
nand U13930 (N_13930,N_13179,N_12447);
and U13931 (N_13931,N_12528,N_13155);
nand U13932 (N_13932,N_12858,N_12905);
xnor U13933 (N_13933,N_12282,N_13048);
nand U13934 (N_13934,N_13022,N_13291);
nor U13935 (N_13935,N_12672,N_13261);
nand U13936 (N_13936,N_13062,N_12423);
and U13937 (N_13937,N_12922,N_12443);
nand U13938 (N_13938,N_12459,N_12886);
and U13939 (N_13939,N_13480,N_12377);
nor U13940 (N_13940,N_12401,N_12341);
and U13941 (N_13941,N_12736,N_13301);
nor U13942 (N_13942,N_13170,N_13097);
nor U13943 (N_13943,N_12322,N_12197);
or U13944 (N_13944,N_13294,N_13194);
nor U13945 (N_13945,N_12625,N_12184);
and U13946 (N_13946,N_12653,N_12515);
nor U13947 (N_13947,N_12498,N_13167);
nor U13948 (N_13948,N_12864,N_12320);
nand U13949 (N_13949,N_12957,N_13156);
and U13950 (N_13950,N_13417,N_13411);
nor U13951 (N_13951,N_12933,N_12321);
nand U13952 (N_13952,N_13187,N_13026);
nor U13953 (N_13953,N_12725,N_12083);
and U13954 (N_13954,N_12122,N_13160);
nand U13955 (N_13955,N_13219,N_12954);
xnor U13956 (N_13956,N_13442,N_13328);
nand U13957 (N_13957,N_13053,N_12353);
nand U13958 (N_13958,N_13240,N_12814);
nand U13959 (N_13959,N_12499,N_13262);
and U13960 (N_13960,N_12662,N_12567);
xnor U13961 (N_13961,N_13260,N_12537);
nor U13962 (N_13962,N_12538,N_13010);
and U13963 (N_13963,N_12358,N_13498);
nand U13964 (N_13964,N_12396,N_12303);
nand U13965 (N_13965,N_13386,N_12985);
or U13966 (N_13966,N_13146,N_12824);
nand U13967 (N_13967,N_13253,N_12185);
or U13968 (N_13968,N_12863,N_13109);
nor U13969 (N_13969,N_12888,N_12446);
nand U13970 (N_13970,N_13434,N_13095);
nor U13971 (N_13971,N_12866,N_12194);
nand U13972 (N_13972,N_13317,N_12212);
nand U13973 (N_13973,N_13487,N_12833);
or U13974 (N_13974,N_13096,N_13182);
or U13975 (N_13975,N_12797,N_13025);
or U13976 (N_13976,N_13381,N_13169);
and U13977 (N_13977,N_13392,N_13174);
nand U13978 (N_13978,N_12632,N_12073);
or U13979 (N_13979,N_12123,N_12196);
and U13980 (N_13980,N_13064,N_13087);
and U13981 (N_13981,N_12205,N_12529);
nand U13982 (N_13982,N_13359,N_12647);
nand U13983 (N_13983,N_12159,N_12946);
and U13984 (N_13984,N_12999,N_12747);
or U13985 (N_13985,N_13342,N_12876);
nor U13986 (N_13986,N_12148,N_12973);
nand U13987 (N_13987,N_12573,N_12133);
nand U13988 (N_13988,N_12167,N_13470);
or U13989 (N_13989,N_12469,N_12436);
nor U13990 (N_13990,N_12857,N_12155);
or U13991 (N_13991,N_12169,N_12059);
nor U13992 (N_13992,N_12808,N_12042);
xnor U13993 (N_13993,N_12092,N_12729);
nand U13994 (N_13994,N_12118,N_13368);
and U13995 (N_13995,N_12445,N_12273);
or U13996 (N_13996,N_13251,N_12982);
or U13997 (N_13997,N_12969,N_13326);
nor U13998 (N_13998,N_13044,N_13012);
nor U13999 (N_13999,N_13300,N_13055);
and U14000 (N_14000,N_12356,N_12441);
nand U14001 (N_14001,N_12432,N_13056);
nor U14002 (N_14002,N_13357,N_13478);
nand U14003 (N_14003,N_12368,N_12409);
and U14004 (N_14004,N_12658,N_12304);
or U14005 (N_14005,N_12836,N_13333);
and U14006 (N_14006,N_12785,N_12019);
nor U14007 (N_14007,N_12723,N_13364);
or U14008 (N_14008,N_12285,N_12766);
and U14009 (N_14009,N_12043,N_12805);
and U14010 (N_14010,N_12675,N_13407);
and U14011 (N_14011,N_13015,N_12890);
and U14012 (N_14012,N_13428,N_13203);
nor U14013 (N_14013,N_12597,N_13196);
or U14014 (N_14014,N_12295,N_12851);
nor U14015 (N_14015,N_13367,N_12802);
xnor U14016 (N_14016,N_12104,N_12298);
nor U14017 (N_14017,N_12848,N_12918);
and U14018 (N_14018,N_12784,N_12286);
nor U14019 (N_14019,N_12974,N_12847);
and U14020 (N_14020,N_12369,N_12195);
nand U14021 (N_14021,N_13250,N_12966);
and U14022 (N_14022,N_12569,N_13177);
and U14023 (N_14023,N_12125,N_12894);
or U14024 (N_14024,N_13173,N_13394);
or U14025 (N_14025,N_13472,N_12732);
nor U14026 (N_14026,N_12009,N_13353);
and U14027 (N_14027,N_13323,N_12674);
or U14028 (N_14028,N_12001,N_12769);
or U14029 (N_14029,N_13239,N_13303);
or U14030 (N_14030,N_13031,N_12501);
nand U14031 (N_14031,N_13497,N_12970);
or U14032 (N_14032,N_13320,N_12752);
or U14033 (N_14033,N_12942,N_12949);
nand U14034 (N_14034,N_12892,N_12140);
nand U14035 (N_14035,N_12508,N_12046);
or U14036 (N_14036,N_12908,N_12323);
and U14037 (N_14037,N_12047,N_13252);
nand U14038 (N_14038,N_12397,N_13218);
nand U14039 (N_14039,N_13414,N_12865);
and U14040 (N_14040,N_12681,N_13464);
nor U14041 (N_14041,N_13168,N_12428);
or U14042 (N_14042,N_12227,N_12128);
nand U14043 (N_14043,N_12079,N_12913);
or U14044 (N_14044,N_12164,N_12962);
nor U14045 (N_14045,N_12748,N_12427);
nor U14046 (N_14046,N_12025,N_12697);
nand U14047 (N_14047,N_12071,N_12618);
nand U14048 (N_14048,N_13077,N_12896);
nand U14049 (N_14049,N_12036,N_13334);
or U14050 (N_14050,N_13234,N_13437);
nand U14051 (N_14051,N_12471,N_12481);
nor U14052 (N_14052,N_13230,N_12696);
or U14053 (N_14053,N_12332,N_13018);
or U14054 (N_14054,N_13385,N_12202);
and U14055 (N_14055,N_13191,N_13376);
nand U14056 (N_14056,N_12972,N_12572);
or U14057 (N_14057,N_12667,N_12884);
nand U14058 (N_14058,N_13249,N_13379);
nor U14059 (N_14059,N_12986,N_12022);
xnor U14060 (N_14060,N_12099,N_12403);
nand U14061 (N_14061,N_12221,N_13149);
xnor U14062 (N_14062,N_12216,N_12340);
nor U14063 (N_14063,N_13099,N_12978);
nor U14064 (N_14064,N_12312,N_12951);
nor U14065 (N_14065,N_12649,N_12490);
nor U14066 (N_14066,N_12103,N_12731);
or U14067 (N_14067,N_12663,N_12365);
or U14068 (N_14068,N_12039,N_12274);
and U14069 (N_14069,N_12906,N_12013);
or U14070 (N_14070,N_12139,N_13032);
or U14071 (N_14071,N_12271,N_12520);
nand U14072 (N_14072,N_12448,N_13490);
nor U14073 (N_14073,N_13448,N_12823);
or U14074 (N_14074,N_12989,N_12678);
nand U14075 (N_14075,N_13489,N_12599);
nor U14076 (N_14076,N_12383,N_12788);
nor U14077 (N_14077,N_13265,N_13402);
nor U14078 (N_14078,N_12038,N_12129);
and U14079 (N_14079,N_12927,N_12668);
xnor U14080 (N_14080,N_12188,N_13285);
or U14081 (N_14081,N_12248,N_13435);
or U14082 (N_14082,N_12745,N_13242);
or U14083 (N_14083,N_13162,N_12387);
and U14084 (N_14084,N_13331,N_12172);
or U14085 (N_14085,N_12706,N_13237);
or U14086 (N_14086,N_13164,N_13081);
nor U14087 (N_14087,N_12622,N_13279);
or U14088 (N_14088,N_13075,N_12011);
nor U14089 (N_14089,N_13132,N_12834);
or U14090 (N_14090,N_13499,N_13486);
and U14091 (N_14091,N_12588,N_12881);
and U14092 (N_14092,N_13241,N_13329);
nor U14093 (N_14093,N_13444,N_12277);
nor U14094 (N_14094,N_12812,N_12281);
and U14095 (N_14095,N_13436,N_12602);
nor U14096 (N_14096,N_13100,N_13222);
xor U14097 (N_14097,N_13355,N_12620);
nor U14098 (N_14098,N_12345,N_13256);
or U14099 (N_14099,N_12730,N_12958);
and U14100 (N_14100,N_12313,N_12839);
and U14101 (N_14101,N_12550,N_12463);
or U14102 (N_14102,N_12971,N_13111);
and U14103 (N_14103,N_13372,N_12265);
or U14104 (N_14104,N_13276,N_12778);
nand U14105 (N_14105,N_12361,N_12754);
nor U14106 (N_14106,N_12806,N_13439);
and U14107 (N_14107,N_12832,N_12329);
nor U14108 (N_14108,N_12178,N_13001);
or U14109 (N_14109,N_12577,N_12666);
or U14110 (N_14110,N_13063,N_12828);
nand U14111 (N_14111,N_12088,N_12454);
nand U14112 (N_14112,N_12135,N_12883);
and U14113 (N_14113,N_13079,N_12779);
xor U14114 (N_14114,N_13126,N_12053);
nand U14115 (N_14115,N_12183,N_12138);
nand U14116 (N_14116,N_13002,N_12415);
or U14117 (N_14117,N_13311,N_12669);
nor U14118 (N_14118,N_12293,N_13352);
nor U14119 (N_14119,N_13481,N_12840);
nand U14120 (N_14120,N_12684,N_12781);
nor U14121 (N_14121,N_13441,N_13299);
nand U14122 (N_14122,N_12916,N_12334);
nor U14123 (N_14123,N_12643,N_12052);
and U14124 (N_14124,N_12548,N_12910);
nand U14125 (N_14125,N_12181,N_12268);
nor U14126 (N_14126,N_12761,N_12402);
and U14127 (N_14127,N_13445,N_12855);
xnor U14128 (N_14128,N_12177,N_12414);
or U14129 (N_14129,N_12613,N_12458);
or U14130 (N_14130,N_12161,N_13009);
nor U14131 (N_14131,N_12173,N_13067);
or U14132 (N_14132,N_13066,N_12283);
nand U14133 (N_14133,N_13346,N_12553);
or U14134 (N_14134,N_13151,N_12659);
nor U14135 (N_14135,N_12584,N_13071);
or U14136 (N_14136,N_12932,N_12767);
and U14137 (N_14137,N_12230,N_13391);
nand U14138 (N_14138,N_12278,N_12592);
nand U14139 (N_14139,N_13106,N_13141);
nand U14140 (N_14140,N_12425,N_12276);
nor U14141 (N_14141,N_12246,N_12439);
nand U14142 (N_14142,N_12144,N_13369);
nor U14143 (N_14143,N_12267,N_12065);
nand U14144 (N_14144,N_12120,N_13325);
and U14145 (N_14145,N_12701,N_13232);
or U14146 (N_14146,N_13354,N_13304);
or U14147 (N_14147,N_12699,N_12204);
and U14148 (N_14148,N_12086,N_12111);
and U14149 (N_14149,N_13133,N_13037);
and U14150 (N_14150,N_12262,N_12114);
and U14151 (N_14151,N_13080,N_13185);
nand U14152 (N_14152,N_12305,N_12244);
nand U14153 (N_14153,N_12717,N_12488);
nand U14154 (N_14154,N_12089,N_12486);
nand U14155 (N_14155,N_12931,N_13371);
nor U14156 (N_14156,N_13496,N_13217);
nand U14157 (N_14157,N_13184,N_13043);
and U14158 (N_14158,N_12174,N_12694);
nand U14159 (N_14159,N_13330,N_12854);
nand U14160 (N_14160,N_12270,N_13270);
xor U14161 (N_14161,N_13202,N_13447);
nor U14162 (N_14162,N_12134,N_12822);
nand U14163 (N_14163,N_12759,N_12095);
and U14164 (N_14164,N_12016,N_13396);
and U14165 (N_14165,N_12473,N_12941);
and U14166 (N_14166,N_12226,N_12853);
nor U14167 (N_14167,N_12306,N_13220);
xor U14168 (N_14168,N_12562,N_12438);
nand U14169 (N_14169,N_12735,N_12002);
nand U14170 (N_14170,N_12449,N_12521);
nand U14171 (N_14171,N_12540,N_12774);
and U14172 (N_14172,N_12749,N_13123);
nand U14173 (N_14173,N_12665,N_12080);
nor U14174 (N_14174,N_12707,N_13118);
xor U14175 (N_14175,N_12483,N_13384);
nor U14176 (N_14176,N_12641,N_12024);
and U14177 (N_14177,N_12789,N_12657);
and U14178 (N_14178,N_13209,N_12838);
nor U14179 (N_14179,N_12199,N_13340);
or U14180 (N_14180,N_12815,N_13113);
or U14181 (N_14181,N_12233,N_13038);
or U14182 (N_14182,N_13052,N_12821);
and U14183 (N_14183,N_12116,N_12416);
xnor U14184 (N_14184,N_12909,N_12389);
nor U14185 (N_14185,N_12768,N_12565);
and U14186 (N_14186,N_12899,N_12258);
or U14187 (N_14187,N_12629,N_12990);
nor U14188 (N_14188,N_12879,N_12085);
nor U14189 (N_14189,N_13495,N_13479);
and U14190 (N_14190,N_12049,N_13443);
or U14191 (N_14191,N_13440,N_12837);
and U14192 (N_14192,N_12690,N_13308);
or U14193 (N_14193,N_12157,N_12398);
or U14194 (N_14194,N_13373,N_13358);
nor U14195 (N_14195,N_12776,N_12096);
nand U14196 (N_14196,N_13366,N_12698);
or U14197 (N_14197,N_12628,N_12994);
and U14198 (N_14198,N_13199,N_12284);
xnor U14199 (N_14199,N_12637,N_12279);
nand U14200 (N_14200,N_12350,N_12108);
or U14201 (N_14201,N_12758,N_13310);
nor U14202 (N_14202,N_12783,N_12536);
or U14203 (N_14203,N_12355,N_12482);
nor U14204 (N_14204,N_12795,N_12367);
or U14205 (N_14205,N_13438,N_13221);
nor U14206 (N_14206,N_12734,N_13183);
nand U14207 (N_14207,N_12097,N_13287);
nand U14208 (N_14208,N_12869,N_12453);
nand U14209 (N_14209,N_12517,N_13035);
xor U14210 (N_14210,N_12484,N_12315);
or U14211 (N_14211,N_12920,N_13363);
nand U14212 (N_14212,N_12130,N_12831);
nor U14213 (N_14213,N_12600,N_12474);
nor U14214 (N_14214,N_12843,N_13057);
or U14215 (N_14215,N_12044,N_13458);
nand U14216 (N_14216,N_13462,N_13051);
nand U14217 (N_14217,N_13207,N_12057);
xor U14218 (N_14218,N_12460,N_12408);
nand U14219 (N_14219,N_13452,N_13365);
or U14220 (N_14220,N_13461,N_12492);
nand U14221 (N_14221,N_12380,N_12733);
xor U14222 (N_14222,N_12522,N_12560);
or U14223 (N_14223,N_12242,N_12539);
or U14224 (N_14224,N_12497,N_12030);
nand U14225 (N_14225,N_12670,N_12810);
nand U14226 (N_14226,N_12106,N_13124);
and U14227 (N_14227,N_13054,N_12191);
nand U14228 (N_14228,N_13236,N_12081);
xor U14229 (N_14229,N_13161,N_12714);
nor U14230 (N_14230,N_12817,N_12393);
nor U14231 (N_14231,N_12715,N_12190);
nor U14232 (N_14232,N_12919,N_12594);
and U14233 (N_14233,N_13374,N_12137);
nand U14234 (N_14234,N_13069,N_13309);
and U14235 (N_14235,N_12938,N_13344);
nand U14236 (N_14236,N_13398,N_12773);
xnor U14237 (N_14237,N_13175,N_12006);
nor U14238 (N_14238,N_12621,N_12370);
or U14239 (N_14239,N_13388,N_12603);
and U14240 (N_14240,N_13137,N_12718);
and U14241 (N_14241,N_12470,N_12430);
or U14242 (N_14242,N_12598,N_12462);
or U14243 (N_14243,N_13277,N_12545);
and U14244 (N_14244,N_12564,N_12998);
nand U14245 (N_14245,N_12162,N_12328);
or U14246 (N_14246,N_13475,N_13180);
and U14247 (N_14247,N_13257,N_13139);
nor U14248 (N_14248,N_12711,N_12929);
nand U14249 (N_14249,N_12326,N_12100);
or U14250 (N_14250,N_12224,N_12132);
and U14251 (N_14251,N_12092,N_12712);
or U14252 (N_14252,N_12045,N_12292);
or U14253 (N_14253,N_12621,N_12546);
xnor U14254 (N_14254,N_12765,N_13037);
nand U14255 (N_14255,N_12040,N_12738);
and U14256 (N_14256,N_13197,N_12639);
xnor U14257 (N_14257,N_12797,N_12756);
xnor U14258 (N_14258,N_13093,N_12327);
or U14259 (N_14259,N_12745,N_12370);
nor U14260 (N_14260,N_12709,N_12276);
xnor U14261 (N_14261,N_12609,N_13087);
nor U14262 (N_14262,N_12160,N_13491);
nand U14263 (N_14263,N_13037,N_13488);
and U14264 (N_14264,N_13426,N_12186);
or U14265 (N_14265,N_13080,N_12544);
and U14266 (N_14266,N_12032,N_12358);
or U14267 (N_14267,N_12828,N_13227);
nand U14268 (N_14268,N_13229,N_12440);
or U14269 (N_14269,N_13039,N_13460);
nand U14270 (N_14270,N_13478,N_12487);
and U14271 (N_14271,N_12198,N_12196);
nor U14272 (N_14272,N_12878,N_12890);
and U14273 (N_14273,N_13372,N_12008);
nor U14274 (N_14274,N_12996,N_13435);
or U14275 (N_14275,N_12161,N_13402);
nand U14276 (N_14276,N_12011,N_12501);
nand U14277 (N_14277,N_13148,N_12941);
nand U14278 (N_14278,N_12191,N_12119);
xor U14279 (N_14279,N_12636,N_12690);
nand U14280 (N_14280,N_12921,N_12591);
or U14281 (N_14281,N_13238,N_12506);
nor U14282 (N_14282,N_12758,N_12899);
nand U14283 (N_14283,N_13493,N_12426);
xor U14284 (N_14284,N_12083,N_12013);
and U14285 (N_14285,N_12735,N_12733);
nand U14286 (N_14286,N_12016,N_12639);
or U14287 (N_14287,N_12568,N_13056);
nor U14288 (N_14288,N_12547,N_12644);
nor U14289 (N_14289,N_13453,N_13109);
and U14290 (N_14290,N_13496,N_12853);
and U14291 (N_14291,N_12777,N_12936);
nor U14292 (N_14292,N_12772,N_12845);
and U14293 (N_14293,N_12025,N_12597);
or U14294 (N_14294,N_13436,N_13278);
nor U14295 (N_14295,N_12606,N_12871);
nor U14296 (N_14296,N_13383,N_13486);
or U14297 (N_14297,N_13259,N_13051);
nor U14298 (N_14298,N_13034,N_12360);
nand U14299 (N_14299,N_12219,N_12125);
nor U14300 (N_14300,N_13232,N_12829);
nand U14301 (N_14301,N_12289,N_12903);
and U14302 (N_14302,N_12039,N_12633);
or U14303 (N_14303,N_13115,N_12790);
nor U14304 (N_14304,N_12805,N_12955);
and U14305 (N_14305,N_12089,N_13071);
nor U14306 (N_14306,N_13239,N_13364);
nor U14307 (N_14307,N_13306,N_12366);
and U14308 (N_14308,N_13189,N_12158);
or U14309 (N_14309,N_12212,N_12590);
nand U14310 (N_14310,N_13250,N_12672);
or U14311 (N_14311,N_13247,N_12044);
or U14312 (N_14312,N_13486,N_13039);
nor U14313 (N_14313,N_13255,N_13385);
nand U14314 (N_14314,N_12596,N_13171);
or U14315 (N_14315,N_13429,N_12214);
and U14316 (N_14316,N_13309,N_12920);
and U14317 (N_14317,N_12335,N_12552);
nand U14318 (N_14318,N_12473,N_12917);
xor U14319 (N_14319,N_12784,N_13008);
nor U14320 (N_14320,N_12824,N_12084);
nor U14321 (N_14321,N_12052,N_12116);
or U14322 (N_14322,N_13084,N_12519);
nor U14323 (N_14323,N_12217,N_12251);
nor U14324 (N_14324,N_12356,N_13479);
and U14325 (N_14325,N_12654,N_12729);
nor U14326 (N_14326,N_12503,N_12560);
nor U14327 (N_14327,N_13175,N_12427);
or U14328 (N_14328,N_12793,N_13194);
nor U14329 (N_14329,N_12175,N_13448);
nor U14330 (N_14330,N_13442,N_12265);
nand U14331 (N_14331,N_12642,N_13230);
and U14332 (N_14332,N_12775,N_13003);
and U14333 (N_14333,N_13155,N_12877);
nor U14334 (N_14334,N_12049,N_13055);
or U14335 (N_14335,N_12622,N_13012);
nand U14336 (N_14336,N_13312,N_12975);
and U14337 (N_14337,N_12841,N_12378);
and U14338 (N_14338,N_13370,N_12459);
and U14339 (N_14339,N_12080,N_12643);
or U14340 (N_14340,N_13153,N_12291);
and U14341 (N_14341,N_13032,N_12823);
nor U14342 (N_14342,N_13423,N_12458);
nand U14343 (N_14343,N_13124,N_12122);
or U14344 (N_14344,N_12984,N_12330);
xnor U14345 (N_14345,N_13053,N_12387);
or U14346 (N_14346,N_13451,N_13425);
nor U14347 (N_14347,N_12843,N_13330);
nor U14348 (N_14348,N_12259,N_12382);
nor U14349 (N_14349,N_13151,N_12263);
or U14350 (N_14350,N_12463,N_12470);
nor U14351 (N_14351,N_12886,N_13253);
nor U14352 (N_14352,N_12847,N_13440);
nand U14353 (N_14353,N_12400,N_12265);
or U14354 (N_14354,N_12448,N_12651);
nor U14355 (N_14355,N_13077,N_12657);
or U14356 (N_14356,N_12883,N_13132);
nor U14357 (N_14357,N_12136,N_13356);
nor U14358 (N_14358,N_12995,N_12110);
or U14359 (N_14359,N_12725,N_12104);
xnor U14360 (N_14360,N_13110,N_12772);
nand U14361 (N_14361,N_12802,N_12281);
nor U14362 (N_14362,N_13099,N_12547);
nor U14363 (N_14363,N_12600,N_13108);
and U14364 (N_14364,N_12103,N_12883);
or U14365 (N_14365,N_13249,N_12378);
and U14366 (N_14366,N_12561,N_13362);
and U14367 (N_14367,N_12611,N_13337);
and U14368 (N_14368,N_12856,N_13266);
or U14369 (N_14369,N_13323,N_13311);
or U14370 (N_14370,N_13474,N_13230);
and U14371 (N_14371,N_13054,N_13124);
xnor U14372 (N_14372,N_12409,N_13324);
nor U14373 (N_14373,N_12654,N_12959);
and U14374 (N_14374,N_12644,N_13450);
or U14375 (N_14375,N_12758,N_13265);
or U14376 (N_14376,N_12787,N_12681);
nand U14377 (N_14377,N_12496,N_12687);
nor U14378 (N_14378,N_12028,N_13072);
nor U14379 (N_14379,N_13107,N_12004);
and U14380 (N_14380,N_13381,N_12649);
nor U14381 (N_14381,N_13427,N_12855);
nand U14382 (N_14382,N_13199,N_12762);
or U14383 (N_14383,N_12308,N_13024);
and U14384 (N_14384,N_12107,N_12589);
or U14385 (N_14385,N_12940,N_13151);
and U14386 (N_14386,N_12731,N_12978);
and U14387 (N_14387,N_13312,N_12277);
and U14388 (N_14388,N_13086,N_12289);
nor U14389 (N_14389,N_12167,N_12567);
nand U14390 (N_14390,N_12240,N_12190);
or U14391 (N_14391,N_12763,N_13229);
nor U14392 (N_14392,N_13242,N_12943);
nand U14393 (N_14393,N_13073,N_12932);
or U14394 (N_14394,N_13420,N_13373);
nor U14395 (N_14395,N_12282,N_13342);
nor U14396 (N_14396,N_12292,N_13389);
nor U14397 (N_14397,N_12503,N_12402);
or U14398 (N_14398,N_12035,N_13224);
nor U14399 (N_14399,N_13332,N_12152);
and U14400 (N_14400,N_13459,N_12450);
or U14401 (N_14401,N_12667,N_12630);
and U14402 (N_14402,N_12262,N_13008);
and U14403 (N_14403,N_12680,N_13471);
xnor U14404 (N_14404,N_13244,N_12995);
and U14405 (N_14405,N_12045,N_13285);
and U14406 (N_14406,N_13302,N_12233);
nor U14407 (N_14407,N_12718,N_13494);
and U14408 (N_14408,N_12116,N_12211);
and U14409 (N_14409,N_12439,N_12583);
or U14410 (N_14410,N_12556,N_12362);
or U14411 (N_14411,N_12293,N_13072);
or U14412 (N_14412,N_13094,N_13301);
nand U14413 (N_14413,N_13192,N_13207);
and U14414 (N_14414,N_13270,N_12685);
and U14415 (N_14415,N_13378,N_13051);
nand U14416 (N_14416,N_12207,N_12343);
nor U14417 (N_14417,N_13487,N_13055);
nand U14418 (N_14418,N_12644,N_12329);
nor U14419 (N_14419,N_12636,N_13123);
and U14420 (N_14420,N_13350,N_12168);
nand U14421 (N_14421,N_12997,N_12016);
nand U14422 (N_14422,N_13485,N_13281);
or U14423 (N_14423,N_13437,N_12314);
or U14424 (N_14424,N_13373,N_12234);
nand U14425 (N_14425,N_12514,N_13114);
nor U14426 (N_14426,N_12380,N_13177);
nand U14427 (N_14427,N_12430,N_13488);
nand U14428 (N_14428,N_12916,N_13472);
and U14429 (N_14429,N_13315,N_13134);
or U14430 (N_14430,N_12670,N_13061);
nor U14431 (N_14431,N_13428,N_13351);
and U14432 (N_14432,N_13025,N_12566);
and U14433 (N_14433,N_12187,N_12327);
xor U14434 (N_14434,N_12457,N_12677);
nand U14435 (N_14435,N_12470,N_12273);
or U14436 (N_14436,N_12602,N_13493);
or U14437 (N_14437,N_13465,N_12275);
or U14438 (N_14438,N_12764,N_12786);
xnor U14439 (N_14439,N_12380,N_13156);
and U14440 (N_14440,N_12591,N_13362);
nand U14441 (N_14441,N_12200,N_12016);
xnor U14442 (N_14442,N_12931,N_12075);
and U14443 (N_14443,N_13374,N_12022);
and U14444 (N_14444,N_12973,N_13051);
nand U14445 (N_14445,N_13376,N_12141);
and U14446 (N_14446,N_13330,N_12605);
and U14447 (N_14447,N_12531,N_12196);
nand U14448 (N_14448,N_13350,N_12051);
nand U14449 (N_14449,N_12947,N_12718);
nand U14450 (N_14450,N_13307,N_12356);
and U14451 (N_14451,N_12959,N_13410);
and U14452 (N_14452,N_12179,N_12080);
or U14453 (N_14453,N_13409,N_12682);
xnor U14454 (N_14454,N_13124,N_12924);
xnor U14455 (N_14455,N_12235,N_13259);
or U14456 (N_14456,N_13096,N_13319);
nand U14457 (N_14457,N_12151,N_12424);
nand U14458 (N_14458,N_12376,N_12773);
and U14459 (N_14459,N_13475,N_12094);
nor U14460 (N_14460,N_12799,N_12625);
or U14461 (N_14461,N_12639,N_13248);
or U14462 (N_14462,N_12929,N_12564);
nand U14463 (N_14463,N_12953,N_12096);
nand U14464 (N_14464,N_12973,N_12555);
nor U14465 (N_14465,N_13082,N_13470);
or U14466 (N_14466,N_12093,N_12229);
and U14467 (N_14467,N_12295,N_12718);
or U14468 (N_14468,N_12804,N_12222);
nor U14469 (N_14469,N_12723,N_12378);
and U14470 (N_14470,N_13217,N_12268);
or U14471 (N_14471,N_12142,N_13295);
xor U14472 (N_14472,N_13265,N_12354);
or U14473 (N_14473,N_12810,N_12951);
nor U14474 (N_14474,N_12985,N_13039);
nor U14475 (N_14475,N_12208,N_12619);
and U14476 (N_14476,N_12761,N_12133);
or U14477 (N_14477,N_12980,N_12188);
or U14478 (N_14478,N_12935,N_12279);
xor U14479 (N_14479,N_12060,N_12297);
or U14480 (N_14480,N_13374,N_12012);
and U14481 (N_14481,N_12932,N_12958);
xor U14482 (N_14482,N_13138,N_12760);
nand U14483 (N_14483,N_12157,N_12246);
and U14484 (N_14484,N_12695,N_12114);
nand U14485 (N_14485,N_12569,N_12406);
nand U14486 (N_14486,N_12729,N_12638);
nand U14487 (N_14487,N_12794,N_12855);
nand U14488 (N_14488,N_12187,N_12810);
nand U14489 (N_14489,N_12324,N_12221);
nand U14490 (N_14490,N_12111,N_13398);
nand U14491 (N_14491,N_12624,N_13220);
and U14492 (N_14492,N_13295,N_13181);
nand U14493 (N_14493,N_12929,N_13345);
and U14494 (N_14494,N_12868,N_12192);
xor U14495 (N_14495,N_12118,N_12293);
or U14496 (N_14496,N_12612,N_13354);
nor U14497 (N_14497,N_12635,N_12525);
nand U14498 (N_14498,N_12867,N_12955);
nand U14499 (N_14499,N_12715,N_12883);
and U14500 (N_14500,N_12599,N_13113);
nor U14501 (N_14501,N_12719,N_13230);
xor U14502 (N_14502,N_13106,N_12773);
and U14503 (N_14503,N_12898,N_12293);
nand U14504 (N_14504,N_12059,N_13157);
and U14505 (N_14505,N_13255,N_12400);
nor U14506 (N_14506,N_12838,N_12342);
or U14507 (N_14507,N_12451,N_12352);
nand U14508 (N_14508,N_12082,N_12002);
nor U14509 (N_14509,N_13419,N_12979);
or U14510 (N_14510,N_12605,N_12737);
nand U14511 (N_14511,N_13220,N_12269);
and U14512 (N_14512,N_12066,N_12083);
nand U14513 (N_14513,N_12978,N_13461);
and U14514 (N_14514,N_12184,N_13265);
and U14515 (N_14515,N_12686,N_12921);
or U14516 (N_14516,N_12911,N_12707);
and U14517 (N_14517,N_13454,N_13481);
nor U14518 (N_14518,N_12548,N_12468);
xor U14519 (N_14519,N_12917,N_13366);
and U14520 (N_14520,N_12697,N_12259);
xnor U14521 (N_14521,N_12161,N_12282);
nand U14522 (N_14522,N_12518,N_12220);
and U14523 (N_14523,N_12506,N_12574);
nor U14524 (N_14524,N_13001,N_13274);
nor U14525 (N_14525,N_13111,N_12774);
and U14526 (N_14526,N_13202,N_12275);
or U14527 (N_14527,N_13317,N_13197);
or U14528 (N_14528,N_12431,N_13100);
and U14529 (N_14529,N_12252,N_13407);
nand U14530 (N_14530,N_13191,N_13035);
nor U14531 (N_14531,N_12156,N_12195);
nand U14532 (N_14532,N_12280,N_13220);
nand U14533 (N_14533,N_13053,N_13338);
nand U14534 (N_14534,N_13327,N_12997);
nand U14535 (N_14535,N_13160,N_13203);
or U14536 (N_14536,N_12211,N_12942);
nand U14537 (N_14537,N_13065,N_12966);
and U14538 (N_14538,N_12713,N_12354);
or U14539 (N_14539,N_12525,N_13091);
nand U14540 (N_14540,N_12072,N_12112);
or U14541 (N_14541,N_12107,N_13260);
and U14542 (N_14542,N_13090,N_12169);
or U14543 (N_14543,N_13424,N_13426);
nand U14544 (N_14544,N_12837,N_12846);
nor U14545 (N_14545,N_13301,N_13064);
nand U14546 (N_14546,N_12769,N_12553);
nand U14547 (N_14547,N_12365,N_13391);
xnor U14548 (N_14548,N_12048,N_13416);
nor U14549 (N_14549,N_12038,N_12110);
nor U14550 (N_14550,N_12207,N_12529);
or U14551 (N_14551,N_13410,N_13466);
and U14552 (N_14552,N_12293,N_13292);
nand U14553 (N_14553,N_12558,N_13195);
nand U14554 (N_14554,N_12939,N_12391);
and U14555 (N_14555,N_12706,N_12799);
nand U14556 (N_14556,N_12070,N_12915);
or U14557 (N_14557,N_12257,N_12639);
nand U14558 (N_14558,N_12687,N_12377);
nor U14559 (N_14559,N_13319,N_13036);
or U14560 (N_14560,N_13050,N_12324);
nor U14561 (N_14561,N_12622,N_13083);
or U14562 (N_14562,N_13198,N_13408);
nor U14563 (N_14563,N_12967,N_12629);
nand U14564 (N_14564,N_12420,N_12351);
nor U14565 (N_14565,N_12254,N_13168);
nand U14566 (N_14566,N_12942,N_13073);
nand U14567 (N_14567,N_13331,N_12216);
xnor U14568 (N_14568,N_13149,N_12356);
nand U14569 (N_14569,N_12542,N_12102);
nor U14570 (N_14570,N_12689,N_12762);
and U14571 (N_14571,N_12518,N_12267);
or U14572 (N_14572,N_13089,N_12347);
nand U14573 (N_14573,N_13350,N_13023);
nand U14574 (N_14574,N_13356,N_12728);
nor U14575 (N_14575,N_13428,N_12165);
or U14576 (N_14576,N_13169,N_12895);
xnor U14577 (N_14577,N_12435,N_12752);
nand U14578 (N_14578,N_12531,N_12921);
and U14579 (N_14579,N_13167,N_12946);
nor U14580 (N_14580,N_13110,N_12010);
or U14581 (N_14581,N_13057,N_13487);
xor U14582 (N_14582,N_13437,N_13193);
and U14583 (N_14583,N_12365,N_13390);
or U14584 (N_14584,N_12763,N_13217);
nand U14585 (N_14585,N_12353,N_12792);
nand U14586 (N_14586,N_13418,N_12485);
nand U14587 (N_14587,N_12604,N_12166);
and U14588 (N_14588,N_13058,N_12403);
and U14589 (N_14589,N_12179,N_12568);
xor U14590 (N_14590,N_13062,N_12390);
nor U14591 (N_14591,N_12027,N_13065);
xnor U14592 (N_14592,N_12150,N_13425);
xnor U14593 (N_14593,N_12953,N_12186);
and U14594 (N_14594,N_12502,N_12251);
and U14595 (N_14595,N_12886,N_13111);
nand U14596 (N_14596,N_12817,N_12458);
nand U14597 (N_14597,N_12064,N_12984);
and U14598 (N_14598,N_12105,N_13002);
and U14599 (N_14599,N_12349,N_12375);
nor U14600 (N_14600,N_13189,N_12137);
or U14601 (N_14601,N_12457,N_12332);
and U14602 (N_14602,N_12342,N_12373);
xor U14603 (N_14603,N_13076,N_12161);
or U14604 (N_14604,N_13441,N_12489);
and U14605 (N_14605,N_12688,N_13044);
and U14606 (N_14606,N_12884,N_13096);
and U14607 (N_14607,N_12774,N_12186);
or U14608 (N_14608,N_13141,N_13367);
and U14609 (N_14609,N_12338,N_12560);
nor U14610 (N_14610,N_13038,N_12271);
nor U14611 (N_14611,N_12105,N_12246);
nand U14612 (N_14612,N_12155,N_13230);
nor U14613 (N_14613,N_13461,N_13337);
or U14614 (N_14614,N_13052,N_12040);
and U14615 (N_14615,N_12926,N_12540);
or U14616 (N_14616,N_12150,N_12507);
or U14617 (N_14617,N_13477,N_12649);
nand U14618 (N_14618,N_12116,N_12290);
or U14619 (N_14619,N_12688,N_13345);
nand U14620 (N_14620,N_13310,N_13330);
nand U14621 (N_14621,N_12552,N_12214);
or U14622 (N_14622,N_12606,N_12710);
and U14623 (N_14623,N_13050,N_13214);
nand U14624 (N_14624,N_12463,N_13498);
xnor U14625 (N_14625,N_12146,N_12052);
and U14626 (N_14626,N_13430,N_12646);
nand U14627 (N_14627,N_12590,N_12928);
nor U14628 (N_14628,N_12636,N_13288);
xnor U14629 (N_14629,N_12414,N_12315);
nand U14630 (N_14630,N_12913,N_13210);
or U14631 (N_14631,N_13294,N_12080);
nand U14632 (N_14632,N_12818,N_13056);
or U14633 (N_14633,N_12622,N_13233);
nor U14634 (N_14634,N_13451,N_12291);
and U14635 (N_14635,N_12655,N_13239);
nand U14636 (N_14636,N_12214,N_12123);
nand U14637 (N_14637,N_13346,N_13332);
nand U14638 (N_14638,N_13227,N_12494);
nor U14639 (N_14639,N_13277,N_12577);
and U14640 (N_14640,N_12743,N_13416);
nand U14641 (N_14641,N_13338,N_13292);
and U14642 (N_14642,N_12432,N_12100);
nor U14643 (N_14643,N_12013,N_13110);
nand U14644 (N_14644,N_13162,N_13237);
nand U14645 (N_14645,N_12802,N_13407);
nand U14646 (N_14646,N_12181,N_13247);
nand U14647 (N_14647,N_12956,N_13408);
nor U14648 (N_14648,N_12306,N_13071);
and U14649 (N_14649,N_13079,N_13491);
nor U14650 (N_14650,N_12946,N_12427);
nor U14651 (N_14651,N_12734,N_12533);
and U14652 (N_14652,N_13058,N_12836);
nor U14653 (N_14653,N_12322,N_12575);
nand U14654 (N_14654,N_12229,N_12236);
or U14655 (N_14655,N_12316,N_12027);
nor U14656 (N_14656,N_13193,N_13062);
nor U14657 (N_14657,N_12148,N_13214);
nor U14658 (N_14658,N_12976,N_12284);
nand U14659 (N_14659,N_13246,N_12891);
nor U14660 (N_14660,N_12258,N_13018);
nand U14661 (N_14661,N_12857,N_12123);
or U14662 (N_14662,N_12870,N_13067);
xnor U14663 (N_14663,N_12607,N_13495);
nand U14664 (N_14664,N_13475,N_12769);
xnor U14665 (N_14665,N_12309,N_13464);
nor U14666 (N_14666,N_13041,N_12061);
or U14667 (N_14667,N_12278,N_12726);
nor U14668 (N_14668,N_13359,N_12797);
nand U14669 (N_14669,N_13317,N_13058);
and U14670 (N_14670,N_12289,N_13454);
or U14671 (N_14671,N_12984,N_13317);
or U14672 (N_14672,N_12029,N_12328);
nor U14673 (N_14673,N_12989,N_12112);
xor U14674 (N_14674,N_12820,N_12631);
nor U14675 (N_14675,N_12961,N_12523);
or U14676 (N_14676,N_12697,N_13077);
and U14677 (N_14677,N_12279,N_12368);
xnor U14678 (N_14678,N_12746,N_12801);
and U14679 (N_14679,N_13276,N_12297);
nand U14680 (N_14680,N_12208,N_13032);
and U14681 (N_14681,N_13215,N_13167);
or U14682 (N_14682,N_13226,N_12346);
or U14683 (N_14683,N_13397,N_13281);
nand U14684 (N_14684,N_12984,N_12615);
or U14685 (N_14685,N_13470,N_12065);
nor U14686 (N_14686,N_12651,N_12262);
nand U14687 (N_14687,N_12222,N_12971);
and U14688 (N_14688,N_13073,N_12855);
xor U14689 (N_14689,N_13427,N_13465);
xor U14690 (N_14690,N_13295,N_12385);
nor U14691 (N_14691,N_13410,N_13171);
xnor U14692 (N_14692,N_12371,N_13283);
nor U14693 (N_14693,N_12510,N_12872);
nor U14694 (N_14694,N_13137,N_12014);
or U14695 (N_14695,N_12558,N_13484);
and U14696 (N_14696,N_12437,N_12907);
nor U14697 (N_14697,N_12624,N_13042);
and U14698 (N_14698,N_12824,N_13371);
or U14699 (N_14699,N_12404,N_12698);
nand U14700 (N_14700,N_12225,N_13206);
and U14701 (N_14701,N_13492,N_12694);
nand U14702 (N_14702,N_12252,N_12126);
or U14703 (N_14703,N_12539,N_12512);
and U14704 (N_14704,N_13077,N_12653);
and U14705 (N_14705,N_12331,N_12242);
xor U14706 (N_14706,N_12154,N_12684);
xor U14707 (N_14707,N_12534,N_13294);
nand U14708 (N_14708,N_12886,N_12484);
nand U14709 (N_14709,N_13433,N_13112);
and U14710 (N_14710,N_12351,N_12151);
and U14711 (N_14711,N_12944,N_13122);
and U14712 (N_14712,N_13414,N_12675);
nand U14713 (N_14713,N_12278,N_12620);
nor U14714 (N_14714,N_12373,N_13383);
nor U14715 (N_14715,N_12152,N_12505);
and U14716 (N_14716,N_12972,N_12801);
and U14717 (N_14717,N_12132,N_12066);
xor U14718 (N_14718,N_12296,N_12821);
and U14719 (N_14719,N_12457,N_12568);
nor U14720 (N_14720,N_12078,N_12701);
nand U14721 (N_14721,N_12696,N_12542);
or U14722 (N_14722,N_13343,N_12486);
and U14723 (N_14723,N_13081,N_12254);
or U14724 (N_14724,N_13416,N_12390);
or U14725 (N_14725,N_12848,N_12373);
or U14726 (N_14726,N_12000,N_13205);
nor U14727 (N_14727,N_13111,N_12630);
or U14728 (N_14728,N_12220,N_13409);
and U14729 (N_14729,N_13063,N_12340);
or U14730 (N_14730,N_12385,N_12580);
nor U14731 (N_14731,N_12419,N_13143);
and U14732 (N_14732,N_12218,N_12162);
nor U14733 (N_14733,N_12073,N_12243);
nand U14734 (N_14734,N_12930,N_13400);
xor U14735 (N_14735,N_13010,N_12912);
nand U14736 (N_14736,N_12075,N_12369);
nor U14737 (N_14737,N_12121,N_13065);
or U14738 (N_14738,N_13007,N_12329);
nor U14739 (N_14739,N_12532,N_12463);
or U14740 (N_14740,N_12780,N_12905);
or U14741 (N_14741,N_13147,N_12508);
nor U14742 (N_14742,N_12027,N_13010);
nor U14743 (N_14743,N_13240,N_13425);
nor U14744 (N_14744,N_13048,N_13322);
nand U14745 (N_14745,N_12072,N_12260);
nand U14746 (N_14746,N_13262,N_12718);
and U14747 (N_14747,N_12272,N_12964);
nor U14748 (N_14748,N_12194,N_13014);
nor U14749 (N_14749,N_12189,N_12419);
and U14750 (N_14750,N_13325,N_12783);
nor U14751 (N_14751,N_13417,N_12254);
nand U14752 (N_14752,N_12351,N_12678);
nand U14753 (N_14753,N_13328,N_12526);
or U14754 (N_14754,N_12359,N_12122);
and U14755 (N_14755,N_13387,N_12390);
nand U14756 (N_14756,N_12732,N_12522);
nor U14757 (N_14757,N_12501,N_12673);
nor U14758 (N_14758,N_13469,N_12393);
nand U14759 (N_14759,N_12764,N_12462);
nand U14760 (N_14760,N_12717,N_12435);
and U14761 (N_14761,N_12574,N_12726);
nor U14762 (N_14762,N_12730,N_12079);
and U14763 (N_14763,N_12245,N_12763);
nor U14764 (N_14764,N_13115,N_12832);
nand U14765 (N_14765,N_12136,N_12736);
and U14766 (N_14766,N_12310,N_12758);
nand U14767 (N_14767,N_13196,N_12020);
nor U14768 (N_14768,N_13209,N_13243);
and U14769 (N_14769,N_12423,N_12473);
and U14770 (N_14770,N_12702,N_12993);
or U14771 (N_14771,N_12136,N_12420);
nand U14772 (N_14772,N_12609,N_13301);
and U14773 (N_14773,N_12106,N_13275);
nor U14774 (N_14774,N_12185,N_13288);
xor U14775 (N_14775,N_12068,N_13269);
nor U14776 (N_14776,N_13448,N_12322);
nor U14777 (N_14777,N_12180,N_12543);
nor U14778 (N_14778,N_13302,N_12210);
nor U14779 (N_14779,N_13151,N_12091);
and U14780 (N_14780,N_13454,N_13369);
nand U14781 (N_14781,N_12601,N_13170);
nor U14782 (N_14782,N_12799,N_12203);
or U14783 (N_14783,N_13104,N_12379);
xnor U14784 (N_14784,N_12006,N_12319);
nor U14785 (N_14785,N_13420,N_13381);
and U14786 (N_14786,N_12531,N_13205);
nor U14787 (N_14787,N_12436,N_13040);
and U14788 (N_14788,N_13481,N_12178);
nand U14789 (N_14789,N_12494,N_13249);
xor U14790 (N_14790,N_12031,N_12278);
or U14791 (N_14791,N_12261,N_12566);
nand U14792 (N_14792,N_12307,N_13461);
nor U14793 (N_14793,N_12669,N_13260);
nor U14794 (N_14794,N_13277,N_12162);
nor U14795 (N_14795,N_13482,N_12777);
nor U14796 (N_14796,N_13022,N_12041);
and U14797 (N_14797,N_12882,N_12534);
or U14798 (N_14798,N_12110,N_12761);
or U14799 (N_14799,N_13261,N_13069);
or U14800 (N_14800,N_12301,N_12606);
nor U14801 (N_14801,N_12734,N_13094);
or U14802 (N_14802,N_12052,N_13445);
nor U14803 (N_14803,N_12890,N_12434);
xor U14804 (N_14804,N_13462,N_12922);
nor U14805 (N_14805,N_12664,N_13414);
and U14806 (N_14806,N_13066,N_13140);
nand U14807 (N_14807,N_12057,N_12886);
nor U14808 (N_14808,N_12809,N_13107);
or U14809 (N_14809,N_13101,N_13419);
nor U14810 (N_14810,N_13497,N_12265);
nor U14811 (N_14811,N_13376,N_12288);
and U14812 (N_14812,N_12037,N_12450);
or U14813 (N_14813,N_12142,N_12624);
or U14814 (N_14814,N_12988,N_12983);
nand U14815 (N_14815,N_13131,N_13496);
and U14816 (N_14816,N_12955,N_12475);
nor U14817 (N_14817,N_12298,N_13403);
nor U14818 (N_14818,N_12383,N_12325);
nor U14819 (N_14819,N_12394,N_12841);
or U14820 (N_14820,N_13241,N_13226);
xor U14821 (N_14821,N_12638,N_12946);
and U14822 (N_14822,N_12693,N_12940);
and U14823 (N_14823,N_12832,N_12789);
or U14824 (N_14824,N_12584,N_12451);
or U14825 (N_14825,N_13370,N_12298);
nor U14826 (N_14826,N_12404,N_12937);
nand U14827 (N_14827,N_13485,N_12441);
and U14828 (N_14828,N_13357,N_12029);
or U14829 (N_14829,N_12707,N_12265);
nand U14830 (N_14830,N_13340,N_12966);
nand U14831 (N_14831,N_12348,N_12719);
and U14832 (N_14832,N_12757,N_12701);
xor U14833 (N_14833,N_12282,N_13449);
nor U14834 (N_14834,N_12819,N_13131);
and U14835 (N_14835,N_12496,N_12414);
and U14836 (N_14836,N_12406,N_12683);
and U14837 (N_14837,N_12829,N_12807);
or U14838 (N_14838,N_12553,N_13215);
and U14839 (N_14839,N_12864,N_12005);
nor U14840 (N_14840,N_12037,N_12957);
nor U14841 (N_14841,N_13299,N_12112);
or U14842 (N_14842,N_13384,N_13306);
nand U14843 (N_14843,N_13104,N_13327);
and U14844 (N_14844,N_13255,N_13291);
nand U14845 (N_14845,N_13306,N_13425);
xnor U14846 (N_14846,N_12900,N_13063);
nand U14847 (N_14847,N_13171,N_12501);
and U14848 (N_14848,N_12289,N_12319);
or U14849 (N_14849,N_12017,N_13370);
nor U14850 (N_14850,N_12455,N_12976);
or U14851 (N_14851,N_12004,N_12896);
and U14852 (N_14852,N_12934,N_12634);
nand U14853 (N_14853,N_13041,N_12606);
nor U14854 (N_14854,N_13010,N_12694);
and U14855 (N_14855,N_12166,N_13189);
nor U14856 (N_14856,N_12047,N_12963);
xor U14857 (N_14857,N_12225,N_13348);
xnor U14858 (N_14858,N_12851,N_12484);
and U14859 (N_14859,N_12956,N_12272);
nand U14860 (N_14860,N_12671,N_13441);
xnor U14861 (N_14861,N_13397,N_12059);
nand U14862 (N_14862,N_13429,N_12623);
or U14863 (N_14863,N_12464,N_12638);
and U14864 (N_14864,N_13050,N_12093);
nor U14865 (N_14865,N_12145,N_13379);
or U14866 (N_14866,N_12369,N_12401);
or U14867 (N_14867,N_12747,N_13242);
nor U14868 (N_14868,N_12496,N_13351);
xor U14869 (N_14869,N_12630,N_12621);
and U14870 (N_14870,N_12591,N_12239);
nand U14871 (N_14871,N_13207,N_12911);
nor U14872 (N_14872,N_12931,N_13290);
or U14873 (N_14873,N_13247,N_12210);
nor U14874 (N_14874,N_12096,N_12696);
nor U14875 (N_14875,N_12457,N_12553);
xnor U14876 (N_14876,N_12396,N_13411);
and U14877 (N_14877,N_12516,N_13094);
nor U14878 (N_14878,N_13310,N_12838);
nor U14879 (N_14879,N_12626,N_12884);
and U14880 (N_14880,N_12374,N_12606);
nor U14881 (N_14881,N_12076,N_12340);
nand U14882 (N_14882,N_13323,N_13035);
nor U14883 (N_14883,N_12325,N_12915);
nand U14884 (N_14884,N_12161,N_13197);
nor U14885 (N_14885,N_12704,N_13401);
nor U14886 (N_14886,N_12570,N_13272);
or U14887 (N_14887,N_13001,N_13406);
nor U14888 (N_14888,N_12692,N_12596);
or U14889 (N_14889,N_13282,N_12697);
or U14890 (N_14890,N_12316,N_12303);
nand U14891 (N_14891,N_13255,N_13068);
nor U14892 (N_14892,N_13421,N_12309);
or U14893 (N_14893,N_13304,N_12405);
nor U14894 (N_14894,N_12210,N_12963);
nand U14895 (N_14895,N_13121,N_12031);
or U14896 (N_14896,N_12266,N_13362);
and U14897 (N_14897,N_12180,N_12074);
nor U14898 (N_14898,N_12591,N_13468);
nor U14899 (N_14899,N_13097,N_12247);
nand U14900 (N_14900,N_12662,N_13181);
nand U14901 (N_14901,N_12411,N_13471);
nor U14902 (N_14902,N_12201,N_13065);
nand U14903 (N_14903,N_12785,N_12393);
or U14904 (N_14904,N_12917,N_13057);
nand U14905 (N_14905,N_12443,N_12431);
nor U14906 (N_14906,N_12896,N_12707);
and U14907 (N_14907,N_12888,N_12925);
nor U14908 (N_14908,N_12987,N_12083);
xor U14909 (N_14909,N_13414,N_13393);
nand U14910 (N_14910,N_12528,N_12068);
nand U14911 (N_14911,N_13219,N_13106);
or U14912 (N_14912,N_13301,N_12148);
and U14913 (N_14913,N_12572,N_12686);
nand U14914 (N_14914,N_13047,N_13438);
nand U14915 (N_14915,N_12653,N_12572);
nor U14916 (N_14916,N_13116,N_12919);
nand U14917 (N_14917,N_12519,N_12515);
nand U14918 (N_14918,N_12782,N_12578);
or U14919 (N_14919,N_13331,N_13472);
and U14920 (N_14920,N_13245,N_13149);
nor U14921 (N_14921,N_13222,N_13077);
or U14922 (N_14922,N_13414,N_13233);
and U14923 (N_14923,N_12280,N_12990);
nand U14924 (N_14924,N_12377,N_13036);
nand U14925 (N_14925,N_12531,N_12312);
xor U14926 (N_14926,N_12599,N_12216);
and U14927 (N_14927,N_12495,N_13494);
or U14928 (N_14928,N_12750,N_12998);
nor U14929 (N_14929,N_12796,N_12778);
and U14930 (N_14930,N_12358,N_13461);
nand U14931 (N_14931,N_12395,N_13453);
and U14932 (N_14932,N_13086,N_13307);
and U14933 (N_14933,N_13012,N_12847);
and U14934 (N_14934,N_13103,N_12817);
and U14935 (N_14935,N_12713,N_12661);
or U14936 (N_14936,N_12240,N_12428);
nor U14937 (N_14937,N_12159,N_12030);
nand U14938 (N_14938,N_13022,N_12169);
nor U14939 (N_14939,N_12648,N_12855);
nand U14940 (N_14940,N_13122,N_12371);
xnor U14941 (N_14941,N_13484,N_12789);
or U14942 (N_14942,N_12133,N_12706);
and U14943 (N_14943,N_12271,N_13280);
and U14944 (N_14944,N_13022,N_13283);
nand U14945 (N_14945,N_12330,N_13065);
nor U14946 (N_14946,N_12168,N_12159);
nand U14947 (N_14947,N_13199,N_12553);
nand U14948 (N_14948,N_12444,N_12126);
or U14949 (N_14949,N_12621,N_12906);
xor U14950 (N_14950,N_13073,N_12448);
nand U14951 (N_14951,N_12362,N_12792);
or U14952 (N_14952,N_12972,N_12733);
nand U14953 (N_14953,N_12259,N_12377);
or U14954 (N_14954,N_12883,N_12397);
and U14955 (N_14955,N_12889,N_13245);
nor U14956 (N_14956,N_12066,N_12865);
or U14957 (N_14957,N_12208,N_12612);
nor U14958 (N_14958,N_12964,N_12718);
nor U14959 (N_14959,N_12026,N_13259);
or U14960 (N_14960,N_12750,N_12721);
nor U14961 (N_14961,N_12292,N_12913);
nor U14962 (N_14962,N_13242,N_12825);
nor U14963 (N_14963,N_13052,N_13104);
and U14964 (N_14964,N_12524,N_12322);
nand U14965 (N_14965,N_12366,N_12446);
or U14966 (N_14966,N_12714,N_12817);
and U14967 (N_14967,N_12809,N_12677);
or U14968 (N_14968,N_12936,N_12143);
and U14969 (N_14969,N_12285,N_13021);
and U14970 (N_14970,N_12436,N_12714);
xnor U14971 (N_14971,N_12622,N_12461);
and U14972 (N_14972,N_13351,N_12925);
and U14973 (N_14973,N_13289,N_12456);
or U14974 (N_14974,N_12056,N_13483);
nand U14975 (N_14975,N_13020,N_13380);
or U14976 (N_14976,N_12410,N_12615);
and U14977 (N_14977,N_12570,N_12543);
and U14978 (N_14978,N_13032,N_13146);
nor U14979 (N_14979,N_12203,N_12412);
or U14980 (N_14980,N_12689,N_12224);
and U14981 (N_14981,N_13356,N_12541);
nor U14982 (N_14982,N_12270,N_13470);
xnor U14983 (N_14983,N_13286,N_13060);
or U14984 (N_14984,N_12695,N_13465);
and U14985 (N_14985,N_13499,N_12297);
or U14986 (N_14986,N_12866,N_12806);
nand U14987 (N_14987,N_12747,N_12771);
nand U14988 (N_14988,N_12617,N_12084);
nor U14989 (N_14989,N_12562,N_13255);
nor U14990 (N_14990,N_13484,N_12998);
or U14991 (N_14991,N_12939,N_12037);
xnor U14992 (N_14992,N_12652,N_12873);
nand U14993 (N_14993,N_12107,N_13041);
nor U14994 (N_14994,N_13334,N_12089);
or U14995 (N_14995,N_13085,N_12187);
and U14996 (N_14996,N_12706,N_12707);
xor U14997 (N_14997,N_12665,N_13471);
and U14998 (N_14998,N_12439,N_12636);
and U14999 (N_14999,N_13391,N_12354);
or UO_0 (O_0,N_13583,N_13543);
nor UO_1 (O_1,N_14801,N_14774);
nor UO_2 (O_2,N_14080,N_13709);
or UO_3 (O_3,N_14876,N_14564);
or UO_4 (O_4,N_13814,N_13915);
and UO_5 (O_5,N_14936,N_14174);
and UO_6 (O_6,N_13878,N_13750);
or UO_7 (O_7,N_13995,N_14879);
or UO_8 (O_8,N_13538,N_14541);
nor UO_9 (O_9,N_13504,N_14413);
or UO_10 (O_10,N_14820,N_14953);
nor UO_11 (O_11,N_14793,N_14993);
xnor UO_12 (O_12,N_13888,N_13766);
nand UO_13 (O_13,N_13974,N_14481);
or UO_14 (O_14,N_14750,N_14212);
or UO_15 (O_15,N_14385,N_13778);
and UO_16 (O_16,N_14300,N_13639);
nand UO_17 (O_17,N_13862,N_14173);
xnor UO_18 (O_18,N_14365,N_14051);
or UO_19 (O_19,N_13875,N_13674);
nand UO_20 (O_20,N_13847,N_13670);
nor UO_21 (O_21,N_14943,N_13932);
nand UO_22 (O_22,N_13746,N_14473);
or UO_23 (O_23,N_14699,N_14949);
nor UO_24 (O_24,N_14797,N_14600);
or UO_25 (O_25,N_14015,N_14304);
or UO_26 (O_26,N_13514,N_14122);
xor UO_27 (O_27,N_14898,N_14239);
or UO_28 (O_28,N_13937,N_13672);
and UO_29 (O_29,N_14794,N_14031);
and UO_30 (O_30,N_14809,N_14107);
or UO_31 (O_31,N_13662,N_14922);
nor UO_32 (O_32,N_14914,N_14892);
or UO_33 (O_33,N_14146,N_14233);
or UO_34 (O_34,N_14204,N_13957);
and UO_35 (O_35,N_14241,N_14288);
nor UO_36 (O_36,N_13757,N_13555);
nand UO_37 (O_37,N_14136,N_14802);
and UO_38 (O_38,N_14361,N_14836);
nand UO_39 (O_39,N_13767,N_13809);
and UO_40 (O_40,N_13864,N_14917);
nor UO_41 (O_41,N_14553,N_14590);
nor UO_42 (O_42,N_13892,N_14334);
nor UO_43 (O_43,N_14569,N_13935);
or UO_44 (O_44,N_13702,N_13721);
nand UO_45 (O_45,N_14965,N_14097);
xnor UO_46 (O_46,N_14971,N_13596);
or UO_47 (O_47,N_13681,N_14065);
nand UO_48 (O_48,N_14333,N_14562);
nand UO_49 (O_49,N_13752,N_14527);
or UO_50 (O_50,N_13890,N_14745);
and UO_51 (O_51,N_14504,N_13677);
and UO_52 (O_52,N_14372,N_14501);
and UO_53 (O_53,N_13887,N_14113);
nor UO_54 (O_54,N_14132,N_14624);
or UO_55 (O_55,N_14875,N_14651);
xnor UO_56 (O_56,N_14225,N_14613);
nor UO_57 (O_57,N_14604,N_14664);
nand UO_58 (O_58,N_14535,N_14418);
or UO_59 (O_59,N_13874,N_14768);
nor UO_60 (O_60,N_14099,N_14157);
or UO_61 (O_61,N_14566,N_14608);
or UO_62 (O_62,N_13943,N_14770);
and UO_63 (O_63,N_13779,N_14800);
and UO_64 (O_64,N_14773,N_14321);
nand UO_65 (O_65,N_14865,N_14027);
or UO_66 (O_66,N_13810,N_13865);
or UO_67 (O_67,N_13613,N_14798);
or UO_68 (O_68,N_14899,N_14596);
and UO_69 (O_69,N_14355,N_14838);
xnor UO_70 (O_70,N_14658,N_14140);
or UO_71 (O_71,N_14280,N_13925);
and UO_72 (O_72,N_14787,N_13858);
or UO_73 (O_73,N_14359,N_14395);
or UO_74 (O_74,N_13747,N_14509);
and UO_75 (O_75,N_13838,N_14606);
nand UO_76 (O_76,N_14062,N_14673);
nand UO_77 (O_77,N_14337,N_13740);
and UO_78 (O_78,N_14450,N_14919);
nor UO_79 (O_79,N_14435,N_14048);
nor UO_80 (O_80,N_13870,N_13671);
and UO_81 (O_81,N_14725,N_14669);
nor UO_82 (O_82,N_14013,N_14442);
and UO_83 (O_83,N_13904,N_14232);
and UO_84 (O_84,N_14551,N_13611);
nor UO_85 (O_85,N_14292,N_14859);
nand UO_86 (O_86,N_14188,N_14490);
or UO_87 (O_87,N_14989,N_14880);
and UO_88 (O_88,N_13930,N_14528);
or UO_89 (O_89,N_13617,N_13537);
or UO_90 (O_90,N_14368,N_13969);
nand UO_91 (O_91,N_14381,N_14067);
nor UO_92 (O_92,N_14915,N_14681);
and UO_93 (O_93,N_14530,N_13685);
and UO_94 (O_94,N_14247,N_13627);
and UO_95 (O_95,N_14180,N_14369);
xnor UO_96 (O_96,N_14694,N_13768);
xor UO_97 (O_97,N_13642,N_14616);
nor UO_98 (O_98,N_14317,N_13563);
or UO_99 (O_99,N_14710,N_14257);
and UO_100 (O_100,N_14677,N_13907);
nor UO_101 (O_101,N_13595,N_14955);
nand UO_102 (O_102,N_14384,N_14558);
xor UO_103 (O_103,N_13698,N_14127);
or UO_104 (O_104,N_14702,N_13895);
nand UO_105 (O_105,N_13513,N_13986);
xor UO_106 (O_106,N_13713,N_14701);
nand UO_107 (O_107,N_14035,N_14390);
nor UO_108 (O_108,N_14828,N_14692);
nand UO_109 (O_109,N_13808,N_14546);
nand UO_110 (O_110,N_14073,N_13585);
nor UO_111 (O_111,N_13552,N_14069);
and UO_112 (O_112,N_14082,N_14370);
or UO_113 (O_113,N_14867,N_13645);
or UO_114 (O_114,N_13851,N_13817);
or UO_115 (O_115,N_14056,N_13620);
nand UO_116 (O_116,N_14499,N_14716);
or UO_117 (O_117,N_13822,N_13773);
nand UO_118 (O_118,N_13812,N_14078);
xnor UO_119 (O_119,N_14106,N_14312);
nor UO_120 (O_120,N_13553,N_14563);
or UO_121 (O_121,N_14030,N_13931);
xor UO_122 (O_122,N_14290,N_13661);
nand UO_123 (O_123,N_13604,N_14962);
or UO_124 (O_124,N_14308,N_13738);
nor UO_125 (O_125,N_14485,N_13632);
nand UO_126 (O_126,N_13988,N_14626);
or UO_127 (O_127,N_14724,N_14025);
nor UO_128 (O_128,N_14958,N_13997);
nand UO_129 (O_129,N_14167,N_13722);
or UO_130 (O_130,N_13868,N_13519);
or UO_131 (O_131,N_14416,N_14218);
nor UO_132 (O_132,N_14900,N_14124);
or UO_133 (O_133,N_14561,N_13684);
or UO_134 (O_134,N_13544,N_14869);
nor UO_135 (O_135,N_13560,N_14843);
or UO_136 (O_136,N_13983,N_14789);
or UO_137 (O_137,N_14480,N_13918);
and UO_138 (O_138,N_13723,N_14448);
or UO_139 (O_139,N_14647,N_14941);
nand UO_140 (O_140,N_14456,N_14686);
and UO_141 (O_141,N_14471,N_14006);
nor UO_142 (O_142,N_14906,N_14454);
nor UO_143 (O_143,N_14482,N_13708);
and UO_144 (O_144,N_14657,N_14761);
xor UO_145 (O_145,N_14438,N_14091);
and UO_146 (O_146,N_14367,N_13625);
nand UO_147 (O_147,N_14555,N_13554);
nand UO_148 (O_148,N_13760,N_14594);
and UO_149 (O_149,N_14848,N_14742);
nand UO_150 (O_150,N_13732,N_14327);
and UO_151 (O_151,N_14133,N_13717);
or UO_152 (O_152,N_13697,N_14617);
nor UO_153 (O_153,N_14937,N_14428);
xnor UO_154 (O_154,N_14753,N_14574);
nor UO_155 (O_155,N_13994,N_14469);
or UO_156 (O_156,N_14245,N_13827);
and UO_157 (O_157,N_14165,N_13704);
nand UO_158 (O_158,N_13512,N_14851);
nand UO_159 (O_159,N_13984,N_14697);
nor UO_160 (O_160,N_14881,N_14659);
or UO_161 (O_161,N_14644,N_14197);
or UO_162 (O_162,N_14039,N_13855);
nor UO_163 (O_163,N_13557,N_14723);
nand UO_164 (O_164,N_14003,N_14618);
or UO_165 (O_165,N_14074,N_14058);
nor UO_166 (O_166,N_14226,N_14883);
or UO_167 (O_167,N_13755,N_14947);
nand UO_168 (O_168,N_13777,N_14084);
nand UO_169 (O_169,N_14829,N_14315);
and UO_170 (O_170,N_14534,N_14096);
and UO_171 (O_171,N_13608,N_13578);
and UO_172 (O_172,N_14302,N_14459);
nor UO_173 (O_173,N_14072,N_14391);
or UO_174 (O_174,N_14727,N_14804);
nand UO_175 (O_175,N_13761,N_14264);
nor UO_176 (O_176,N_13794,N_14913);
nor UO_177 (O_177,N_14595,N_14895);
or UO_178 (O_178,N_14762,N_13837);
nand UO_179 (O_179,N_14511,N_14224);
and UO_180 (O_180,N_13790,N_13597);
xnor UO_181 (O_181,N_14837,N_14000);
and UO_182 (O_182,N_14890,N_14776);
xnor UO_183 (O_183,N_13819,N_14852);
or UO_184 (O_184,N_14529,N_14984);
nand UO_185 (O_185,N_14926,N_14044);
nand UO_186 (O_186,N_14183,N_14491);
and UO_187 (O_187,N_14293,N_14230);
nor UO_188 (O_188,N_14156,N_14001);
xnor UO_189 (O_189,N_14688,N_13891);
nor UO_190 (O_190,N_14741,N_14620);
and UO_191 (O_191,N_14634,N_14863);
and UO_192 (O_192,N_14743,N_14275);
and UO_193 (O_193,N_14130,N_14670);
nor UO_194 (O_194,N_14537,N_14495);
xnor UO_195 (O_195,N_13866,N_13582);
nor UO_196 (O_196,N_14076,N_14665);
xnor UO_197 (O_197,N_14477,N_13700);
xnor UO_198 (O_198,N_14734,N_14389);
or UO_199 (O_199,N_14324,N_13961);
nor UO_200 (O_200,N_14143,N_14339);
xnor UO_201 (O_201,N_14238,N_13971);
nand UO_202 (O_202,N_14930,N_14749);
nor UO_203 (O_203,N_13775,N_13881);
nand UO_204 (O_204,N_14289,N_14593);
nand UO_205 (O_205,N_13791,N_14053);
nand UO_206 (O_206,N_13970,N_14968);
xnor UO_207 (O_207,N_13899,N_14799);
or UO_208 (O_208,N_13852,N_14318);
or UO_209 (O_209,N_13978,N_14924);
nand UO_210 (O_210,N_14497,N_14503);
xnor UO_211 (O_211,N_14022,N_14311);
nand UO_212 (O_212,N_13824,N_14353);
nor UO_213 (O_213,N_14754,N_14427);
xor UO_214 (O_214,N_14316,N_14861);
or UO_215 (O_215,N_14629,N_13889);
or UO_216 (O_216,N_13876,N_14378);
and UO_217 (O_217,N_14720,N_14653);
nand UO_218 (O_218,N_14446,N_14672);
nand UO_219 (O_219,N_14273,N_13926);
nor UO_220 (O_220,N_14933,N_14980);
and UO_221 (O_221,N_14410,N_13561);
and UO_222 (O_222,N_13962,N_14840);
or UO_223 (O_223,N_14627,N_14708);
nand UO_224 (O_224,N_13712,N_13618);
or UO_225 (O_225,N_14813,N_14005);
nand UO_226 (O_226,N_14897,N_14747);
nor UO_227 (O_227,N_13831,N_14777);
nand UO_228 (O_228,N_13676,N_14190);
or UO_229 (O_229,N_14252,N_14085);
or UO_230 (O_230,N_14194,N_13534);
nor UO_231 (O_231,N_13748,N_14407);
xor UO_232 (O_232,N_14995,N_14307);
nand UO_233 (O_233,N_14319,N_13707);
and UO_234 (O_234,N_14896,N_14376);
xnor UO_235 (O_235,N_13829,N_14976);
xor UO_236 (O_236,N_14795,N_14236);
or UO_237 (O_237,N_14019,N_14573);
and UO_238 (O_238,N_14102,N_14021);
or UO_239 (O_239,N_13951,N_13637);
nand UO_240 (O_240,N_13913,N_14847);
or UO_241 (O_241,N_13694,N_14717);
nor UO_242 (O_242,N_14791,N_14115);
nand UO_243 (O_243,N_13525,N_14117);
nand UO_244 (O_244,N_14575,N_14826);
or UO_245 (O_245,N_13634,N_14927);
and UO_246 (O_246,N_14584,N_13678);
or UO_247 (O_247,N_13638,N_14109);
and UO_248 (O_248,N_14655,N_13541);
xnor UO_249 (O_249,N_14952,N_14916);
nor UO_250 (O_250,N_14360,N_14228);
and UO_251 (O_251,N_13664,N_13692);
nor UO_252 (O_252,N_14583,N_14274);
nand UO_253 (O_253,N_14888,N_14248);
or UO_254 (O_254,N_13735,N_14542);
nor UO_255 (O_255,N_14012,N_13830);
and UO_256 (O_256,N_13584,N_14344);
xnor UO_257 (O_257,N_14493,N_13523);
and UO_258 (O_258,N_14401,N_14277);
nand UO_259 (O_259,N_14145,N_14163);
nor UO_260 (O_260,N_14964,N_14974);
or UO_261 (O_261,N_13614,N_14223);
or UO_262 (O_262,N_14790,N_14332);
nand UO_263 (O_263,N_13844,N_14784);
nor UO_264 (O_264,N_13762,N_13739);
and UO_265 (O_265,N_13653,N_13575);
and UO_266 (O_266,N_13548,N_14816);
xnor UO_267 (O_267,N_13857,N_14287);
nor UO_268 (O_268,N_14008,N_13576);
nand UO_269 (O_269,N_13823,N_14028);
nor UO_270 (O_270,N_14077,N_14862);
nor UO_271 (O_271,N_14782,N_14671);
nand UO_272 (O_272,N_14020,N_13649);
or UO_273 (O_273,N_13743,N_14712);
or UO_274 (O_274,N_13797,N_14766);
or UO_275 (O_275,N_13912,N_14556);
or UO_276 (O_276,N_14217,N_14599);
nand UO_277 (O_277,N_14153,N_14550);
or UO_278 (O_278,N_13689,N_14063);
xor UO_279 (O_279,N_14415,N_13648);
or UO_280 (O_280,N_14079,N_13947);
xnor UO_281 (O_281,N_14181,N_14615);
and UO_282 (O_282,N_13569,N_13622);
or UO_283 (O_283,N_14641,N_13641);
or UO_284 (O_284,N_14612,N_13528);
and UO_285 (O_285,N_14703,N_13659);
and UO_286 (O_286,N_13594,N_14767);
nor UO_287 (O_287,N_14904,N_14685);
xnor UO_288 (O_288,N_14886,N_14577);
nand UO_289 (O_289,N_14975,N_14630);
nand UO_290 (O_290,N_14948,N_14162);
or UO_291 (O_291,N_14954,N_14040);
or UO_292 (O_292,N_13900,N_14193);
nand UO_293 (O_293,N_14540,N_14487);
nor UO_294 (O_294,N_14780,N_14329);
or UO_295 (O_295,N_13897,N_14873);
nor UO_296 (O_296,N_13894,N_13610);
or UO_297 (O_297,N_14352,N_13896);
xnor UO_298 (O_298,N_14320,N_14341);
and UO_299 (O_299,N_14309,N_13950);
xor UO_300 (O_300,N_13908,N_14160);
and UO_301 (O_301,N_13651,N_14614);
or UO_302 (O_302,N_14945,N_14400);
or UO_303 (O_303,N_13564,N_14377);
xnor UO_304 (O_304,N_13501,N_14402);
xor UO_305 (O_305,N_14760,N_13964);
nand UO_306 (O_306,N_13796,N_13898);
nor UO_307 (O_307,N_14757,N_14220);
nand UO_308 (O_308,N_13787,N_14739);
or UO_309 (O_309,N_14923,N_14981);
xnor UO_310 (O_310,N_13929,N_14696);
nor UO_311 (O_311,N_14414,N_14882);
nand UO_312 (O_312,N_14552,N_14387);
or UO_313 (O_313,N_13631,N_13588);
or UO_314 (O_314,N_14322,N_14089);
nand UO_315 (O_315,N_14137,N_14269);
nand UO_316 (O_316,N_14810,N_13774);
nor UO_317 (O_317,N_14819,N_13522);
nor UO_318 (O_318,N_14706,N_14885);
nor UO_319 (O_319,N_13607,N_14314);
nand UO_320 (O_320,N_14397,N_13656);
and UO_321 (O_321,N_14521,N_14066);
nor UO_322 (O_322,N_14973,N_14354);
nand UO_323 (O_323,N_13658,N_13644);
or UO_324 (O_324,N_14514,N_13784);
or UO_325 (O_325,N_14205,N_14198);
nor UO_326 (O_326,N_13826,N_14538);
or UO_327 (O_327,N_14796,N_14938);
and UO_328 (O_328,N_14570,N_14211);
or UO_329 (O_329,N_13630,N_14603);
or UO_330 (O_330,N_13598,N_13903);
nor UO_331 (O_331,N_14411,N_14166);
or UO_332 (O_332,N_14931,N_13628);
or UO_333 (O_333,N_14272,N_14656);
or UO_334 (O_334,N_14421,N_14479);
or UO_335 (O_335,N_13567,N_14364);
nor UO_336 (O_336,N_13696,N_14271);
nand UO_337 (O_337,N_14437,N_14484);
or UO_338 (O_338,N_14925,N_14513);
and UO_339 (O_339,N_13799,N_13780);
or UO_340 (O_340,N_14689,N_14158);
and UO_341 (O_341,N_14472,N_14187);
nand UO_342 (O_342,N_14977,N_14347);
nor UO_343 (O_343,N_14565,N_13815);
or UO_344 (O_344,N_13990,N_13516);
nand UO_345 (O_345,N_14866,N_13643);
and UO_346 (O_346,N_14719,N_14023);
nand UO_347 (O_347,N_13728,N_14894);
nor UO_348 (O_348,N_14523,N_14213);
and UO_349 (O_349,N_14940,N_14609);
or UO_350 (O_350,N_13813,N_13727);
nor UO_351 (O_351,N_14932,N_14823);
xor UO_352 (O_352,N_14786,N_14464);
nand UO_353 (O_353,N_13916,N_14687);
xnor UO_354 (O_354,N_14281,N_14854);
or UO_355 (O_355,N_13612,N_14821);
or UO_356 (O_356,N_14441,N_14519);
nor UO_357 (O_357,N_14970,N_14999);
or UO_358 (O_358,N_14060,N_14474);
or UO_359 (O_359,N_14335,N_13836);
and UO_360 (O_360,N_14219,N_14726);
xor UO_361 (O_361,N_14986,N_14602);
or UO_362 (O_362,N_14557,N_13921);
nand UO_363 (O_363,N_14476,N_13909);
and UO_364 (O_364,N_14141,N_13940);
and UO_365 (O_365,N_13781,N_14921);
or UO_366 (O_366,N_14095,N_14496);
nor UO_367 (O_367,N_14215,N_14452);
or UO_368 (O_368,N_14234,N_14559);
nand UO_369 (O_369,N_14123,N_13959);
nor UO_370 (O_370,N_14253,N_13860);
nor UO_371 (O_371,N_14568,N_14751);
xor UO_372 (O_372,N_14972,N_14532);
and UO_373 (O_373,N_14346,N_14845);
or UO_374 (O_374,N_14830,N_14149);
or UO_375 (O_375,N_14805,N_13803);
or UO_376 (O_376,N_13952,N_13589);
or UO_377 (O_377,N_13764,N_14803);
or UO_378 (O_378,N_13871,N_14508);
xnor UO_379 (O_379,N_13724,N_14822);
nand UO_380 (O_380,N_14990,N_14874);
xnor UO_381 (O_381,N_14114,N_13505);
nand UO_382 (O_382,N_14910,N_14808);
and UO_383 (O_383,N_14992,N_14147);
xor UO_384 (O_384,N_14765,N_13811);
or UO_385 (O_385,N_14522,N_13953);
or UO_386 (O_386,N_13786,N_13845);
nor UO_387 (O_387,N_14591,N_13849);
nand UO_388 (O_388,N_13510,N_13686);
nor UO_389 (O_389,N_13906,N_14038);
nand UO_390 (O_390,N_14052,N_13835);
and UO_391 (O_391,N_13869,N_14817);
xor UO_392 (O_392,N_14486,N_13745);
nand UO_393 (O_393,N_14049,N_13683);
or UO_394 (O_394,N_14285,N_13795);
nand UO_395 (O_395,N_14439,N_13967);
and UO_396 (O_396,N_14718,N_14029);
or UO_397 (O_397,N_14177,N_14134);
nand UO_398 (O_398,N_13705,N_13734);
nor UO_399 (O_399,N_14018,N_14889);
nand UO_400 (O_400,N_13882,N_13821);
nor UO_401 (O_401,N_14560,N_13591);
nor UO_402 (O_402,N_14891,N_14175);
or UO_403 (O_403,N_14963,N_13518);
or UO_404 (O_404,N_14849,N_13539);
or UO_405 (O_405,N_13919,N_14887);
or UO_406 (O_406,N_14547,N_14957);
and UO_407 (O_407,N_14978,N_14011);
nand UO_408 (O_408,N_14094,N_14383);
nor UO_409 (O_409,N_14988,N_13503);
or UO_410 (O_410,N_13818,N_13893);
nor UO_411 (O_411,N_14375,N_13675);
xnor UO_412 (O_412,N_13652,N_14126);
nand UO_413 (O_413,N_13979,N_14168);
xor UO_414 (O_414,N_13936,N_13825);
and UO_415 (O_415,N_13633,N_14396);
and UO_416 (O_416,N_14358,N_13859);
and UO_417 (O_417,N_13885,N_14444);
nor UO_418 (O_418,N_14267,N_13843);
or UO_419 (O_419,N_14336,N_13565);
and UO_420 (O_420,N_14036,N_14545);
nor UO_421 (O_421,N_13980,N_14934);
or UO_422 (O_422,N_14240,N_14150);
xor UO_423 (O_423,N_13600,N_13958);
nor UO_424 (O_424,N_14764,N_14858);
nor UO_425 (O_425,N_14152,N_13527);
nand UO_426 (O_426,N_14108,N_13792);
and UO_427 (O_427,N_13788,N_14299);
and UO_428 (O_428,N_14404,N_13731);
and UO_429 (O_429,N_14192,N_14398);
nor UO_430 (O_430,N_13949,N_14246);
and UO_431 (O_431,N_13854,N_13730);
nor UO_432 (O_432,N_13945,N_14517);
nand UO_433 (O_433,N_14092,N_13793);
and UO_434 (O_434,N_14667,N_14161);
nand UO_435 (O_435,N_14735,N_14884);
nand UO_436 (O_436,N_14666,N_14393);
nand UO_437 (O_437,N_14250,N_13636);
or UO_438 (O_438,N_14462,N_13573);
nor UO_439 (O_439,N_14251,N_14216);
nor UO_440 (O_440,N_13580,N_14244);
and UO_441 (O_441,N_14740,N_14942);
and UO_442 (O_442,N_14242,N_13832);
nand UO_443 (O_443,N_14356,N_13763);
nor UO_444 (O_444,N_13842,N_13867);
nand UO_445 (O_445,N_14675,N_14331);
nor UO_446 (O_446,N_14055,N_14643);
nor UO_447 (O_447,N_14901,N_14283);
nand UO_448 (O_448,N_13593,N_13574);
nand UO_449 (O_449,N_13695,N_14179);
xnor UO_450 (O_450,N_14700,N_14016);
or UO_451 (O_451,N_14661,N_13839);
nand UO_452 (O_452,N_14775,N_14721);
and UO_453 (O_453,N_13587,N_14195);
nor UO_454 (O_454,N_13693,N_14433);
nand UO_455 (O_455,N_14772,N_14640);
nand UO_456 (O_456,N_14409,N_14405);
nand UO_457 (O_457,N_13954,N_14424);
and UO_458 (O_458,N_13993,N_14440);
nand UO_459 (O_459,N_14057,N_14632);
or UO_460 (O_460,N_14961,N_13846);
xor UO_461 (O_461,N_14908,N_13540);
nor UO_462 (O_462,N_13798,N_14297);
and UO_463 (O_463,N_14690,N_14576);
nand UO_464 (O_464,N_14121,N_13883);
and UO_465 (O_465,N_14350,N_13547);
or UO_466 (O_466,N_14009,N_14182);
nor UO_467 (O_467,N_13725,N_14492);
nand UO_468 (O_468,N_13920,N_14373);
xor UO_469 (O_469,N_13989,N_14579);
nand UO_470 (O_470,N_13960,N_14142);
or UO_471 (O_471,N_13556,N_14905);
xnor UO_472 (O_472,N_13816,N_14844);
or UO_473 (O_473,N_13942,N_14728);
nor UO_474 (O_474,N_14680,N_14505);
and UO_475 (O_475,N_14068,N_14746);
nor UO_476 (O_476,N_13529,N_14572);
or UO_477 (O_477,N_14323,N_13669);
and UO_478 (O_478,N_14588,N_14510);
nand UO_479 (O_479,N_14357,N_14607);
nand UO_480 (O_480,N_13850,N_14169);
and UO_481 (O_481,N_14148,N_13769);
and UO_482 (O_482,N_14419,N_13647);
or UO_483 (O_483,N_14209,N_14516);
and UO_484 (O_484,N_14825,N_13783);
nor UO_485 (O_485,N_13619,N_13714);
or UO_486 (O_486,N_13879,N_13741);
or UO_487 (O_487,N_14266,N_14944);
nand UO_488 (O_488,N_14270,N_14709);
and UO_489 (O_489,N_14758,N_14155);
nor UO_490 (O_490,N_13756,N_14737);
xor UO_491 (O_491,N_14120,N_14868);
and UO_492 (O_492,N_13679,N_13657);
nor UO_493 (O_493,N_13710,N_13917);
nor UO_494 (O_494,N_14164,N_13688);
nand UO_495 (O_495,N_13806,N_14154);
xnor UO_496 (O_496,N_14105,N_14682);
or UO_497 (O_497,N_13736,N_13535);
nand UO_498 (O_498,N_13733,N_14351);
and UO_499 (O_499,N_14104,N_13663);
nand UO_500 (O_500,N_14589,N_13640);
nor UO_501 (O_501,N_14646,N_14468);
nor UO_502 (O_502,N_14619,N_14420);
nand UO_503 (O_503,N_14711,N_14792);
nor UO_504 (O_504,N_13549,N_14112);
nand UO_505 (O_505,N_14636,N_13515);
xnor UO_506 (O_506,N_14610,N_14637);
nand UO_507 (O_507,N_13840,N_13690);
and UO_508 (O_508,N_14601,N_13626);
or UO_509 (O_509,N_13910,N_13880);
nand UO_510 (O_510,N_13603,N_14611);
and UO_511 (O_511,N_14831,N_14276);
and UO_512 (O_512,N_14581,N_13841);
and UO_513 (O_513,N_14278,N_14445);
and UO_514 (O_514,N_14841,N_14969);
or UO_515 (O_515,N_14412,N_13524);
and UO_516 (O_516,N_14585,N_13623);
nor UO_517 (O_517,N_13615,N_14447);
or UO_518 (O_518,N_13744,N_14432);
nor UO_519 (O_519,N_14779,N_13687);
nand UO_520 (O_520,N_13765,N_13772);
or UO_521 (O_521,N_14306,N_13570);
nand UO_522 (O_522,N_14348,N_14678);
xnor UO_523 (O_523,N_14732,N_14118);
or UO_524 (O_524,N_14186,N_14536);
nor UO_525 (O_525,N_13807,N_14191);
nand UO_526 (O_526,N_14343,N_14531);
or UO_527 (O_527,N_14363,N_14507);
or UO_528 (O_528,N_13771,N_14037);
and UO_529 (O_529,N_13972,N_14325);
and UO_530 (O_530,N_14781,N_14778);
nor UO_531 (O_531,N_13530,N_13938);
nand UO_532 (O_532,N_13872,N_13718);
nor UO_533 (O_533,N_13532,N_14729);
or UO_534 (O_534,N_13550,N_14024);
nand UO_535 (O_535,N_14684,N_14263);
or UO_536 (O_536,N_13719,N_13665);
xor UO_537 (O_537,N_14683,N_14338);
or UO_538 (O_538,N_14128,N_14034);
or UO_539 (O_539,N_14693,N_13861);
or UO_540 (O_540,N_14047,N_14451);
xnor UO_541 (O_541,N_14059,N_14827);
and UO_542 (O_542,N_13551,N_14214);
or UO_543 (O_543,N_13701,N_14045);
nor UO_544 (O_544,N_13737,N_14648);
or UO_545 (O_545,N_13965,N_13699);
nor UO_546 (O_546,N_14458,N_13800);
nand UO_547 (O_547,N_13616,N_14301);
or UO_548 (O_548,N_14835,N_14070);
nand UO_549 (O_549,N_14434,N_14371);
nand UO_550 (O_550,N_14582,N_14135);
nor UO_551 (O_551,N_14979,N_14633);
or UO_552 (O_552,N_13956,N_14403);
nor UO_553 (O_553,N_13602,N_14983);
or UO_554 (O_554,N_14928,N_14254);
nand UO_555 (O_555,N_14548,N_14465);
nor UO_556 (O_556,N_13828,N_14506);
or UO_557 (O_557,N_14533,N_13706);
or UO_558 (O_558,N_14642,N_14785);
xor UO_559 (O_559,N_14380,N_14625);
nand UO_560 (O_560,N_14255,N_14959);
nor UO_561 (O_561,N_14086,N_14935);
and UO_562 (O_562,N_14834,N_14093);
nor UO_563 (O_563,N_14623,N_14631);
nand UO_564 (O_564,N_14125,N_14679);
and UO_565 (O_565,N_14567,N_14259);
nor UO_566 (O_566,N_14707,N_14704);
or UO_567 (O_567,N_14026,N_13914);
and UO_568 (O_568,N_14676,N_14587);
or UO_569 (O_569,N_14176,N_13691);
and UO_570 (O_570,N_13902,N_14478);
nand UO_571 (O_571,N_14518,N_13715);
nand UO_572 (O_572,N_14399,N_14443);
and UO_573 (O_573,N_14628,N_14151);
or UO_574 (O_574,N_14422,N_14303);
nor UO_575 (O_575,N_14083,N_13782);
or UO_576 (O_576,N_14635,N_14014);
xnor UO_577 (O_577,N_14081,N_13654);
nand UO_578 (O_578,N_14695,N_14206);
and UO_579 (O_579,N_14842,N_14116);
nor UO_580 (O_580,N_14996,N_14663);
and UO_581 (O_581,N_13577,N_14714);
nand UO_582 (O_582,N_14621,N_14870);
nor UO_583 (O_583,N_13933,N_13856);
xor UO_584 (O_584,N_14202,N_14172);
nand UO_585 (O_585,N_14806,N_14296);
and UO_586 (O_586,N_13834,N_14466);
nand UO_587 (O_587,N_13968,N_14249);
nand UO_588 (O_588,N_13606,N_14771);
and UO_589 (O_589,N_14966,N_14453);
nand UO_590 (O_590,N_13758,N_14812);
xor UO_591 (O_591,N_14131,N_13801);
nor UO_592 (O_592,N_14738,N_14429);
nand UO_593 (O_593,N_14298,N_14200);
or UO_594 (O_594,N_13922,N_14227);
and UO_595 (O_595,N_13507,N_14903);
nor UO_596 (O_596,N_14877,N_14998);
and UO_597 (O_597,N_14388,N_13533);
xor UO_598 (O_598,N_14041,N_13629);
or UO_599 (O_599,N_14071,N_14101);
nand UO_600 (O_600,N_13963,N_14184);
or UO_601 (O_601,N_14605,N_13590);
and UO_602 (O_602,N_13749,N_14649);
or UO_603 (O_603,N_13601,N_14208);
nor UO_604 (O_604,N_14543,N_14436);
nand UO_605 (O_605,N_13500,N_14460);
xnor UO_606 (O_606,N_13517,N_14262);
nor UO_607 (O_607,N_14736,N_13973);
and UO_608 (O_608,N_13572,N_14032);
nand UO_609 (O_609,N_14455,N_14342);
and UO_610 (O_610,N_13966,N_13599);
or UO_611 (O_611,N_14909,N_14201);
and UO_612 (O_612,N_13877,N_13511);
or UO_613 (O_613,N_13581,N_14652);
and UO_614 (O_614,N_14850,N_14502);
nor UO_615 (O_615,N_14406,N_14956);
nand UO_616 (O_616,N_14294,N_13873);
nor UO_617 (O_617,N_14002,N_13998);
nand UO_618 (O_618,N_14853,N_14129);
nor UO_619 (O_619,N_13562,N_14500);
nand UO_620 (O_620,N_14987,N_14043);
and UO_621 (O_621,N_13673,N_14902);
or UO_622 (O_622,N_14878,N_14730);
nor UO_623 (O_623,N_14488,N_13977);
nand UO_624 (O_624,N_13502,N_13621);
and UO_625 (O_625,N_13624,N_14064);
and UO_626 (O_626,N_14638,N_14713);
nor UO_627 (O_627,N_14457,N_14982);
nor UO_628 (O_628,N_13545,N_14010);
and UO_629 (O_629,N_14857,N_14744);
nor UO_630 (O_630,N_14467,N_14295);
nand UO_631 (O_631,N_13655,N_14178);
nor UO_632 (O_632,N_14960,N_13999);
and UO_633 (O_633,N_14261,N_14991);
or UO_634 (O_634,N_13720,N_13526);
nor UO_635 (O_635,N_13660,N_14715);
xor UO_636 (O_636,N_13884,N_14814);
and UO_637 (O_637,N_14098,N_14475);
xor UO_638 (O_638,N_14571,N_13901);
or UO_639 (O_639,N_14515,N_14139);
or UO_640 (O_640,N_13742,N_14090);
or UO_641 (O_641,N_13716,N_14386);
or UO_642 (O_642,N_14622,N_13558);
or UO_643 (O_643,N_14382,N_14752);
or UO_644 (O_644,N_14660,N_13955);
nor UO_645 (O_645,N_14119,N_14592);
nand UO_646 (O_646,N_14811,N_13776);
xor UO_647 (O_647,N_14203,N_14408);
nand UO_648 (O_648,N_14379,N_13759);
nor UO_649 (O_649,N_13939,N_14196);
and UO_650 (O_650,N_13886,N_14313);
nor UO_651 (O_651,N_14939,N_13566);
nor UO_652 (O_652,N_14430,N_14833);
and UO_653 (O_653,N_14832,N_14668);
nand UO_654 (O_654,N_14075,N_14985);
nand UO_655 (O_655,N_14731,N_13754);
or UO_656 (O_656,N_14967,N_14872);
nor UO_657 (O_657,N_14839,N_14645);
or UO_658 (O_658,N_14907,N_14815);
nand UO_659 (O_659,N_13975,N_13646);
nand UO_660 (O_660,N_13927,N_14291);
and UO_661 (O_661,N_14756,N_14512);
or UO_662 (O_662,N_14498,N_13981);
nand UO_663 (O_663,N_14580,N_14763);
nor UO_664 (O_664,N_14256,N_14691);
and UO_665 (O_665,N_14286,N_14705);
or UO_666 (O_666,N_13976,N_14463);
nor UO_667 (O_667,N_13992,N_13520);
or UO_668 (O_668,N_14994,N_13911);
nand UO_669 (O_669,N_14310,N_14951);
or UO_670 (O_670,N_14586,N_14759);
nor UO_671 (O_671,N_13579,N_13650);
or UO_672 (O_672,N_14918,N_14426);
or UO_673 (O_673,N_14210,N_14258);
nand UO_674 (O_674,N_14138,N_14345);
nor UO_675 (O_675,N_14349,N_14394);
nor UO_676 (O_676,N_14860,N_14470);
xnor UO_677 (O_677,N_13934,N_14417);
and UO_678 (O_678,N_14366,N_13991);
nand UO_679 (O_679,N_13753,N_13905);
nand UO_680 (O_680,N_14265,N_14461);
or UO_681 (O_681,N_14237,N_14755);
or UO_682 (O_682,N_14674,N_14362);
and UO_683 (O_683,N_14549,N_13635);
or UO_684 (O_684,N_13542,N_14017);
and UO_685 (O_685,N_14554,N_13833);
xnor UO_686 (O_686,N_14856,N_14698);
or UO_687 (O_687,N_14061,N_13928);
or UO_688 (O_688,N_14520,N_14392);
or UO_689 (O_689,N_13667,N_13751);
and UO_690 (O_690,N_14004,N_13531);
and UO_691 (O_691,N_13571,N_14088);
and UO_692 (O_692,N_14100,N_14733);
or UO_693 (O_693,N_14110,N_14231);
nor UO_694 (O_694,N_14207,N_13682);
nor UO_695 (O_695,N_14243,N_14374);
nor UO_696 (O_696,N_14046,N_13609);
and UO_697 (O_697,N_14929,N_14111);
nand UO_698 (O_698,N_14159,N_14783);
or UO_699 (O_699,N_14425,N_13785);
nor UO_700 (O_700,N_13804,N_13820);
or UO_701 (O_701,N_14222,N_14722);
nor UO_702 (O_702,N_13944,N_13546);
nor UO_703 (O_703,N_14748,N_14449);
and UO_704 (O_704,N_13802,N_14946);
nor UO_705 (O_705,N_14007,N_14284);
and UO_706 (O_706,N_14911,N_14189);
and UO_707 (O_707,N_13509,N_14103);
or UO_708 (O_708,N_13711,N_14578);
nand UO_709 (O_709,N_13506,N_13703);
and UO_710 (O_710,N_14654,N_14260);
and UO_711 (O_711,N_14871,N_14639);
xnor UO_712 (O_712,N_13941,N_14539);
nand UO_713 (O_713,N_13536,N_13924);
nand UO_714 (O_714,N_14340,N_14912);
nor UO_715 (O_715,N_14268,N_13605);
nor UO_716 (O_716,N_14221,N_13726);
nor UO_717 (O_717,N_13985,N_14185);
nand UO_718 (O_718,N_14650,N_13521);
or UO_719 (O_719,N_14235,N_13592);
and UO_720 (O_720,N_13789,N_13668);
nor UO_721 (O_721,N_13982,N_14864);
nand UO_722 (O_722,N_13848,N_14328);
nand UO_723 (O_723,N_14524,N_14997);
nand UO_724 (O_724,N_14920,N_13586);
or UO_725 (O_725,N_13805,N_14855);
nand UO_726 (O_726,N_14597,N_13853);
xor UO_727 (O_727,N_13948,N_14087);
and UO_728 (O_728,N_14305,N_14483);
or UO_729 (O_729,N_14489,N_14279);
nand UO_730 (O_730,N_13559,N_14171);
nand UO_731 (O_731,N_13863,N_14769);
or UO_732 (O_732,N_14423,N_14846);
nand UO_733 (O_733,N_14807,N_14282);
or UO_734 (O_734,N_14170,N_13729);
nand UO_735 (O_735,N_14950,N_14330);
nand UO_736 (O_736,N_14544,N_14054);
nand UO_737 (O_737,N_14525,N_14526);
nand UO_738 (O_738,N_14431,N_13996);
nor UO_739 (O_739,N_13666,N_13508);
nor UO_740 (O_740,N_14788,N_14598);
nor UO_741 (O_741,N_13568,N_13770);
nor UO_742 (O_742,N_14199,N_14824);
or UO_743 (O_743,N_14494,N_14818);
and UO_744 (O_744,N_14662,N_13987);
or UO_745 (O_745,N_14042,N_13946);
nor UO_746 (O_746,N_14050,N_13680);
nor UO_747 (O_747,N_14893,N_14229);
nor UO_748 (O_748,N_14144,N_14326);
nand UO_749 (O_749,N_14033,N_13923);
nand UO_750 (O_750,N_13621,N_13807);
or UO_751 (O_751,N_13872,N_14232);
nand UO_752 (O_752,N_13643,N_14043);
or UO_753 (O_753,N_13620,N_14736);
or UO_754 (O_754,N_14282,N_14784);
nand UO_755 (O_755,N_13974,N_13784);
nand UO_756 (O_756,N_14056,N_14388);
xor UO_757 (O_757,N_14211,N_14059);
nand UO_758 (O_758,N_13587,N_13715);
or UO_759 (O_759,N_14804,N_14677);
nand UO_760 (O_760,N_13516,N_14377);
or UO_761 (O_761,N_14064,N_14302);
nand UO_762 (O_762,N_14331,N_13524);
and UO_763 (O_763,N_13514,N_14876);
or UO_764 (O_764,N_14549,N_13807);
or UO_765 (O_765,N_14839,N_13587);
nand UO_766 (O_766,N_14634,N_14645);
nand UO_767 (O_767,N_14192,N_14484);
and UO_768 (O_768,N_14330,N_14609);
nor UO_769 (O_769,N_14641,N_14496);
and UO_770 (O_770,N_14981,N_13978);
nor UO_771 (O_771,N_13581,N_13521);
nand UO_772 (O_772,N_13530,N_14720);
or UO_773 (O_773,N_13978,N_14758);
or UO_774 (O_774,N_14535,N_14679);
or UO_775 (O_775,N_13580,N_14246);
nor UO_776 (O_776,N_14501,N_13979);
and UO_777 (O_777,N_13970,N_14370);
nor UO_778 (O_778,N_13808,N_14793);
or UO_779 (O_779,N_13979,N_13765);
nand UO_780 (O_780,N_14694,N_13654);
and UO_781 (O_781,N_13529,N_14579);
nand UO_782 (O_782,N_13873,N_14983);
nand UO_783 (O_783,N_13985,N_13691);
or UO_784 (O_784,N_13739,N_13693);
nand UO_785 (O_785,N_14482,N_14675);
nand UO_786 (O_786,N_14864,N_13706);
nand UO_787 (O_787,N_13562,N_14009);
nor UO_788 (O_788,N_13881,N_13664);
nor UO_789 (O_789,N_14867,N_14183);
nor UO_790 (O_790,N_14178,N_14160);
xnor UO_791 (O_791,N_14836,N_13995);
xnor UO_792 (O_792,N_14165,N_14908);
nand UO_793 (O_793,N_14670,N_14032);
nand UO_794 (O_794,N_14787,N_14502);
and UO_795 (O_795,N_14776,N_13523);
and UO_796 (O_796,N_14467,N_14462);
nand UO_797 (O_797,N_14312,N_14814);
nand UO_798 (O_798,N_14743,N_13698);
nor UO_799 (O_799,N_13853,N_13883);
xor UO_800 (O_800,N_13966,N_13821);
xor UO_801 (O_801,N_13945,N_14860);
nor UO_802 (O_802,N_14760,N_14266);
nand UO_803 (O_803,N_14150,N_14371);
and UO_804 (O_804,N_14964,N_14102);
and UO_805 (O_805,N_14194,N_14103);
and UO_806 (O_806,N_14652,N_14265);
nand UO_807 (O_807,N_14279,N_13763);
nand UO_808 (O_808,N_14695,N_13599);
nor UO_809 (O_809,N_13873,N_13584);
nor UO_810 (O_810,N_14063,N_14923);
nand UO_811 (O_811,N_14484,N_14294);
xnor UO_812 (O_812,N_13951,N_14321);
or UO_813 (O_813,N_13535,N_13873);
nand UO_814 (O_814,N_13599,N_13920);
nand UO_815 (O_815,N_13711,N_14809);
and UO_816 (O_816,N_13731,N_13611);
nand UO_817 (O_817,N_14171,N_13942);
nand UO_818 (O_818,N_14664,N_13682);
nor UO_819 (O_819,N_14641,N_13647);
nand UO_820 (O_820,N_13820,N_14058);
and UO_821 (O_821,N_13551,N_14624);
or UO_822 (O_822,N_13888,N_13765);
nand UO_823 (O_823,N_14375,N_14458);
nor UO_824 (O_824,N_13785,N_14564);
nand UO_825 (O_825,N_14592,N_14276);
nand UO_826 (O_826,N_14232,N_14531);
nor UO_827 (O_827,N_14508,N_14928);
nand UO_828 (O_828,N_13846,N_14456);
or UO_829 (O_829,N_14468,N_14445);
xnor UO_830 (O_830,N_14265,N_14813);
and UO_831 (O_831,N_14013,N_14601);
nor UO_832 (O_832,N_14970,N_13782);
nor UO_833 (O_833,N_14872,N_13642);
nand UO_834 (O_834,N_14135,N_14519);
nand UO_835 (O_835,N_13793,N_13668);
nand UO_836 (O_836,N_13799,N_13617);
and UO_837 (O_837,N_13977,N_14570);
or UO_838 (O_838,N_13608,N_14483);
nand UO_839 (O_839,N_14947,N_14929);
or UO_840 (O_840,N_14982,N_13974);
or UO_841 (O_841,N_13622,N_14254);
nor UO_842 (O_842,N_14187,N_14495);
nand UO_843 (O_843,N_13907,N_13612);
nor UO_844 (O_844,N_13699,N_14581);
and UO_845 (O_845,N_14043,N_14865);
nand UO_846 (O_846,N_14689,N_13576);
nor UO_847 (O_847,N_14356,N_14536);
or UO_848 (O_848,N_14901,N_14638);
and UO_849 (O_849,N_14778,N_13603);
or UO_850 (O_850,N_14207,N_14586);
and UO_851 (O_851,N_14059,N_13977);
nand UO_852 (O_852,N_14154,N_13514);
nand UO_853 (O_853,N_13939,N_13953);
and UO_854 (O_854,N_14544,N_14822);
nand UO_855 (O_855,N_14968,N_14367);
nor UO_856 (O_856,N_14914,N_13912);
nor UO_857 (O_857,N_13926,N_14059);
nor UO_858 (O_858,N_13722,N_14386);
or UO_859 (O_859,N_14221,N_14244);
nand UO_860 (O_860,N_14710,N_14457);
xnor UO_861 (O_861,N_14300,N_14650);
nand UO_862 (O_862,N_14947,N_13726);
nor UO_863 (O_863,N_13865,N_14175);
xor UO_864 (O_864,N_14916,N_14583);
or UO_865 (O_865,N_14609,N_13876);
or UO_866 (O_866,N_14171,N_14284);
nand UO_867 (O_867,N_13899,N_14123);
or UO_868 (O_868,N_14948,N_14575);
and UO_869 (O_869,N_14904,N_14171);
and UO_870 (O_870,N_14920,N_14851);
and UO_871 (O_871,N_14625,N_14382);
nand UO_872 (O_872,N_14769,N_14585);
nand UO_873 (O_873,N_13990,N_14261);
nand UO_874 (O_874,N_14574,N_13856);
or UO_875 (O_875,N_13632,N_13978);
and UO_876 (O_876,N_14293,N_13722);
and UO_877 (O_877,N_14885,N_14391);
nand UO_878 (O_878,N_14546,N_13987);
and UO_879 (O_879,N_14576,N_14278);
xor UO_880 (O_880,N_14566,N_13732);
nand UO_881 (O_881,N_13662,N_14999);
nand UO_882 (O_882,N_14377,N_13574);
nor UO_883 (O_883,N_13917,N_14219);
nand UO_884 (O_884,N_13735,N_14401);
nor UO_885 (O_885,N_13824,N_14011);
nor UO_886 (O_886,N_14016,N_14967);
and UO_887 (O_887,N_14093,N_14459);
nor UO_888 (O_888,N_14135,N_14970);
or UO_889 (O_889,N_14186,N_13800);
or UO_890 (O_890,N_14583,N_14813);
nor UO_891 (O_891,N_13667,N_14738);
or UO_892 (O_892,N_14234,N_13932);
and UO_893 (O_893,N_14774,N_14621);
or UO_894 (O_894,N_13793,N_14924);
or UO_895 (O_895,N_13970,N_14590);
nand UO_896 (O_896,N_14287,N_14371);
nand UO_897 (O_897,N_14352,N_14920);
nor UO_898 (O_898,N_13924,N_14488);
or UO_899 (O_899,N_13844,N_14949);
and UO_900 (O_900,N_14457,N_14868);
and UO_901 (O_901,N_13750,N_14035);
nand UO_902 (O_902,N_14249,N_14616);
and UO_903 (O_903,N_14205,N_14893);
and UO_904 (O_904,N_13828,N_14028);
and UO_905 (O_905,N_14504,N_14260);
nor UO_906 (O_906,N_13635,N_14828);
xor UO_907 (O_907,N_14554,N_14801);
nand UO_908 (O_908,N_13869,N_14093);
and UO_909 (O_909,N_13690,N_14416);
nor UO_910 (O_910,N_14925,N_13605);
nor UO_911 (O_911,N_13896,N_14931);
or UO_912 (O_912,N_14513,N_14239);
and UO_913 (O_913,N_14613,N_13716);
xnor UO_914 (O_914,N_13702,N_14926);
and UO_915 (O_915,N_14059,N_14085);
nand UO_916 (O_916,N_14473,N_13868);
xnor UO_917 (O_917,N_13913,N_13933);
xnor UO_918 (O_918,N_14626,N_14891);
nor UO_919 (O_919,N_14424,N_14910);
nor UO_920 (O_920,N_14252,N_13649);
or UO_921 (O_921,N_14217,N_14716);
or UO_922 (O_922,N_14226,N_13628);
nor UO_923 (O_923,N_13710,N_14633);
nor UO_924 (O_924,N_13574,N_13641);
nor UO_925 (O_925,N_14513,N_14291);
nand UO_926 (O_926,N_14101,N_13938);
nand UO_927 (O_927,N_14595,N_14680);
nand UO_928 (O_928,N_13907,N_14610);
xor UO_929 (O_929,N_14187,N_14543);
xor UO_930 (O_930,N_14502,N_14375);
and UO_931 (O_931,N_13845,N_14421);
xnor UO_932 (O_932,N_14764,N_14438);
nand UO_933 (O_933,N_13685,N_14314);
nand UO_934 (O_934,N_14927,N_13767);
and UO_935 (O_935,N_14434,N_14046);
nand UO_936 (O_936,N_14490,N_14180);
or UO_937 (O_937,N_13626,N_13589);
nor UO_938 (O_938,N_13596,N_13584);
nand UO_939 (O_939,N_13595,N_14362);
and UO_940 (O_940,N_13990,N_13844);
nor UO_941 (O_941,N_14969,N_14592);
and UO_942 (O_942,N_14365,N_13938);
nand UO_943 (O_943,N_14237,N_13947);
and UO_944 (O_944,N_13844,N_13550);
nor UO_945 (O_945,N_14933,N_13622);
nor UO_946 (O_946,N_13538,N_13773);
or UO_947 (O_947,N_14327,N_14205);
nor UO_948 (O_948,N_14814,N_14369);
nand UO_949 (O_949,N_14625,N_14387);
and UO_950 (O_950,N_14315,N_14563);
or UO_951 (O_951,N_14792,N_14665);
and UO_952 (O_952,N_14028,N_13650);
xnor UO_953 (O_953,N_13854,N_13699);
xnor UO_954 (O_954,N_13748,N_14037);
or UO_955 (O_955,N_14199,N_14818);
nor UO_956 (O_956,N_13676,N_14323);
xnor UO_957 (O_957,N_14029,N_13848);
nand UO_958 (O_958,N_14255,N_14977);
nor UO_959 (O_959,N_14150,N_14137);
nand UO_960 (O_960,N_13648,N_14762);
nand UO_961 (O_961,N_14662,N_13780);
and UO_962 (O_962,N_14610,N_13668);
and UO_963 (O_963,N_14749,N_13977);
nor UO_964 (O_964,N_13688,N_14322);
nor UO_965 (O_965,N_14539,N_14850);
nand UO_966 (O_966,N_14555,N_14173);
or UO_967 (O_967,N_14003,N_14079);
and UO_968 (O_968,N_14483,N_13945);
nand UO_969 (O_969,N_14944,N_14646);
and UO_970 (O_970,N_14578,N_13750);
nor UO_971 (O_971,N_14513,N_14248);
nand UO_972 (O_972,N_14851,N_13883);
nor UO_973 (O_973,N_14871,N_13624);
nand UO_974 (O_974,N_14158,N_14893);
nor UO_975 (O_975,N_14178,N_14239);
or UO_976 (O_976,N_14415,N_13878);
and UO_977 (O_977,N_13616,N_14438);
or UO_978 (O_978,N_13811,N_13565);
or UO_979 (O_979,N_14677,N_14071);
xor UO_980 (O_980,N_14915,N_14096);
and UO_981 (O_981,N_14975,N_14055);
or UO_982 (O_982,N_13985,N_13568);
or UO_983 (O_983,N_14827,N_14368);
xnor UO_984 (O_984,N_14081,N_13650);
xnor UO_985 (O_985,N_13556,N_14896);
or UO_986 (O_986,N_13903,N_14435);
and UO_987 (O_987,N_14112,N_13690);
nand UO_988 (O_988,N_14741,N_14912);
or UO_989 (O_989,N_14306,N_14619);
nand UO_990 (O_990,N_14236,N_14835);
and UO_991 (O_991,N_13763,N_14364);
xnor UO_992 (O_992,N_13895,N_14685);
and UO_993 (O_993,N_14210,N_14310);
and UO_994 (O_994,N_14005,N_14945);
or UO_995 (O_995,N_13609,N_14469);
and UO_996 (O_996,N_13572,N_14957);
nor UO_997 (O_997,N_13894,N_14861);
nor UO_998 (O_998,N_13732,N_13989);
xnor UO_999 (O_999,N_13758,N_13606);
and UO_1000 (O_1000,N_13522,N_14991);
nand UO_1001 (O_1001,N_14008,N_14581);
nor UO_1002 (O_1002,N_13715,N_13915);
nor UO_1003 (O_1003,N_14708,N_14938);
or UO_1004 (O_1004,N_14232,N_13730);
nand UO_1005 (O_1005,N_14667,N_14938);
nor UO_1006 (O_1006,N_14308,N_14316);
or UO_1007 (O_1007,N_13799,N_14414);
or UO_1008 (O_1008,N_13852,N_13862);
and UO_1009 (O_1009,N_13556,N_13761);
nor UO_1010 (O_1010,N_14098,N_13511);
xnor UO_1011 (O_1011,N_14689,N_14804);
or UO_1012 (O_1012,N_14090,N_14405);
nand UO_1013 (O_1013,N_14708,N_14462);
and UO_1014 (O_1014,N_14886,N_14218);
nand UO_1015 (O_1015,N_14385,N_14584);
nor UO_1016 (O_1016,N_14125,N_14424);
nand UO_1017 (O_1017,N_13813,N_13778);
or UO_1018 (O_1018,N_13775,N_14340);
or UO_1019 (O_1019,N_14104,N_14042);
nand UO_1020 (O_1020,N_13621,N_14365);
nand UO_1021 (O_1021,N_14489,N_14114);
nor UO_1022 (O_1022,N_13813,N_14750);
nor UO_1023 (O_1023,N_13810,N_13760);
nand UO_1024 (O_1024,N_14422,N_14958);
or UO_1025 (O_1025,N_14014,N_14338);
or UO_1026 (O_1026,N_14566,N_14311);
or UO_1027 (O_1027,N_14410,N_14888);
nand UO_1028 (O_1028,N_14608,N_14489);
and UO_1029 (O_1029,N_14962,N_14786);
nand UO_1030 (O_1030,N_14590,N_14576);
nor UO_1031 (O_1031,N_14153,N_14465);
xor UO_1032 (O_1032,N_13641,N_14533);
or UO_1033 (O_1033,N_13721,N_14425);
nand UO_1034 (O_1034,N_14258,N_14419);
or UO_1035 (O_1035,N_14110,N_14095);
or UO_1036 (O_1036,N_14810,N_14905);
or UO_1037 (O_1037,N_14204,N_13578);
nor UO_1038 (O_1038,N_13854,N_14985);
nor UO_1039 (O_1039,N_13747,N_14423);
and UO_1040 (O_1040,N_13950,N_14764);
xnor UO_1041 (O_1041,N_14842,N_14984);
or UO_1042 (O_1042,N_14444,N_14539);
or UO_1043 (O_1043,N_13911,N_14683);
nand UO_1044 (O_1044,N_14714,N_13780);
and UO_1045 (O_1045,N_14431,N_14547);
or UO_1046 (O_1046,N_14090,N_14551);
and UO_1047 (O_1047,N_13905,N_14168);
nand UO_1048 (O_1048,N_13890,N_14512);
nor UO_1049 (O_1049,N_14560,N_14954);
and UO_1050 (O_1050,N_13744,N_14791);
nor UO_1051 (O_1051,N_13524,N_14761);
or UO_1052 (O_1052,N_14693,N_14555);
nand UO_1053 (O_1053,N_14766,N_14368);
xnor UO_1054 (O_1054,N_14045,N_14100);
nor UO_1055 (O_1055,N_14563,N_14024);
nand UO_1056 (O_1056,N_14449,N_14690);
or UO_1057 (O_1057,N_14711,N_14404);
and UO_1058 (O_1058,N_13986,N_14399);
or UO_1059 (O_1059,N_13978,N_14323);
and UO_1060 (O_1060,N_13840,N_13980);
or UO_1061 (O_1061,N_14494,N_14010);
nor UO_1062 (O_1062,N_13951,N_13557);
nand UO_1063 (O_1063,N_13685,N_14173);
or UO_1064 (O_1064,N_14042,N_14475);
or UO_1065 (O_1065,N_14973,N_14789);
nor UO_1066 (O_1066,N_13775,N_14911);
and UO_1067 (O_1067,N_13883,N_13800);
or UO_1068 (O_1068,N_13771,N_13815);
and UO_1069 (O_1069,N_14595,N_13768);
or UO_1070 (O_1070,N_14490,N_14166);
or UO_1071 (O_1071,N_13688,N_14207);
nand UO_1072 (O_1072,N_14538,N_14983);
and UO_1073 (O_1073,N_13567,N_14526);
nor UO_1074 (O_1074,N_13501,N_14351);
or UO_1075 (O_1075,N_13654,N_13820);
nand UO_1076 (O_1076,N_14204,N_13600);
or UO_1077 (O_1077,N_13641,N_13635);
xnor UO_1078 (O_1078,N_14171,N_14407);
xor UO_1079 (O_1079,N_14765,N_14591);
or UO_1080 (O_1080,N_14867,N_13782);
nor UO_1081 (O_1081,N_14126,N_14336);
nand UO_1082 (O_1082,N_14162,N_14702);
nand UO_1083 (O_1083,N_14059,N_13530);
and UO_1084 (O_1084,N_14604,N_14510);
or UO_1085 (O_1085,N_14675,N_14688);
nand UO_1086 (O_1086,N_14201,N_13748);
or UO_1087 (O_1087,N_14868,N_13566);
nor UO_1088 (O_1088,N_13525,N_14072);
nand UO_1089 (O_1089,N_13602,N_14228);
or UO_1090 (O_1090,N_14644,N_13616);
or UO_1091 (O_1091,N_14772,N_14265);
nand UO_1092 (O_1092,N_14245,N_14059);
nor UO_1093 (O_1093,N_14948,N_14126);
or UO_1094 (O_1094,N_14194,N_14961);
and UO_1095 (O_1095,N_14382,N_13756);
nand UO_1096 (O_1096,N_14562,N_13868);
nand UO_1097 (O_1097,N_14848,N_14075);
or UO_1098 (O_1098,N_13718,N_14619);
or UO_1099 (O_1099,N_14940,N_14886);
nor UO_1100 (O_1100,N_14927,N_14854);
xnor UO_1101 (O_1101,N_14222,N_14256);
and UO_1102 (O_1102,N_14335,N_13967);
xnor UO_1103 (O_1103,N_14302,N_13563);
nor UO_1104 (O_1104,N_14550,N_13581);
xnor UO_1105 (O_1105,N_13843,N_13921);
xnor UO_1106 (O_1106,N_14226,N_14928);
and UO_1107 (O_1107,N_14351,N_14088);
nand UO_1108 (O_1108,N_14784,N_14291);
or UO_1109 (O_1109,N_14775,N_13645);
and UO_1110 (O_1110,N_14764,N_13676);
nor UO_1111 (O_1111,N_14971,N_13513);
nand UO_1112 (O_1112,N_14250,N_14161);
and UO_1113 (O_1113,N_13750,N_14062);
and UO_1114 (O_1114,N_14280,N_13541);
nor UO_1115 (O_1115,N_14995,N_14370);
or UO_1116 (O_1116,N_14483,N_14185);
or UO_1117 (O_1117,N_13606,N_14963);
nor UO_1118 (O_1118,N_14918,N_14868);
or UO_1119 (O_1119,N_14424,N_14577);
nor UO_1120 (O_1120,N_14250,N_14470);
or UO_1121 (O_1121,N_14626,N_14572);
and UO_1122 (O_1122,N_13540,N_13629);
nor UO_1123 (O_1123,N_13715,N_14292);
and UO_1124 (O_1124,N_14665,N_14515);
nor UO_1125 (O_1125,N_14808,N_13651);
nand UO_1126 (O_1126,N_13611,N_14905);
and UO_1127 (O_1127,N_14745,N_13535);
and UO_1128 (O_1128,N_14698,N_14901);
or UO_1129 (O_1129,N_14442,N_13744);
nand UO_1130 (O_1130,N_14049,N_14541);
xor UO_1131 (O_1131,N_14458,N_14155);
nor UO_1132 (O_1132,N_14757,N_14402);
nor UO_1133 (O_1133,N_14837,N_13668);
or UO_1134 (O_1134,N_13584,N_14727);
or UO_1135 (O_1135,N_13547,N_13573);
nor UO_1136 (O_1136,N_14793,N_14806);
xor UO_1137 (O_1137,N_13706,N_13591);
and UO_1138 (O_1138,N_14405,N_14278);
or UO_1139 (O_1139,N_14957,N_14044);
or UO_1140 (O_1140,N_13830,N_14937);
xor UO_1141 (O_1141,N_14299,N_14275);
nor UO_1142 (O_1142,N_14531,N_14181);
nor UO_1143 (O_1143,N_13929,N_14598);
nor UO_1144 (O_1144,N_13766,N_14316);
or UO_1145 (O_1145,N_14891,N_14096);
nand UO_1146 (O_1146,N_14194,N_14240);
nor UO_1147 (O_1147,N_14980,N_13932);
nand UO_1148 (O_1148,N_13850,N_14601);
and UO_1149 (O_1149,N_14949,N_14118);
or UO_1150 (O_1150,N_14439,N_13875);
and UO_1151 (O_1151,N_14480,N_14893);
nor UO_1152 (O_1152,N_14318,N_14749);
or UO_1153 (O_1153,N_14576,N_13939);
nor UO_1154 (O_1154,N_13890,N_13622);
nand UO_1155 (O_1155,N_14367,N_14221);
or UO_1156 (O_1156,N_14605,N_13771);
nand UO_1157 (O_1157,N_14187,N_14992);
nor UO_1158 (O_1158,N_14167,N_14881);
and UO_1159 (O_1159,N_13712,N_14884);
and UO_1160 (O_1160,N_13734,N_14724);
and UO_1161 (O_1161,N_13778,N_13924);
xnor UO_1162 (O_1162,N_14566,N_14881);
nand UO_1163 (O_1163,N_14206,N_13792);
and UO_1164 (O_1164,N_13571,N_14773);
nand UO_1165 (O_1165,N_14996,N_14034);
and UO_1166 (O_1166,N_14700,N_13746);
and UO_1167 (O_1167,N_14044,N_14936);
or UO_1168 (O_1168,N_13524,N_14373);
nand UO_1169 (O_1169,N_13861,N_14443);
nand UO_1170 (O_1170,N_14383,N_14891);
nand UO_1171 (O_1171,N_13928,N_14357);
or UO_1172 (O_1172,N_14270,N_13533);
nand UO_1173 (O_1173,N_14025,N_14743);
or UO_1174 (O_1174,N_14551,N_13927);
or UO_1175 (O_1175,N_14090,N_13729);
and UO_1176 (O_1176,N_14489,N_14424);
and UO_1177 (O_1177,N_13739,N_13942);
nand UO_1178 (O_1178,N_14528,N_13510);
nor UO_1179 (O_1179,N_13944,N_14329);
nor UO_1180 (O_1180,N_14701,N_14559);
xor UO_1181 (O_1181,N_13985,N_13660);
or UO_1182 (O_1182,N_14425,N_14740);
nor UO_1183 (O_1183,N_14697,N_14012);
nor UO_1184 (O_1184,N_13823,N_14373);
nand UO_1185 (O_1185,N_14808,N_13825);
or UO_1186 (O_1186,N_14714,N_13552);
or UO_1187 (O_1187,N_14416,N_14701);
or UO_1188 (O_1188,N_13752,N_14909);
or UO_1189 (O_1189,N_13897,N_14302);
and UO_1190 (O_1190,N_13576,N_14601);
nor UO_1191 (O_1191,N_14065,N_14840);
xor UO_1192 (O_1192,N_14010,N_14513);
or UO_1193 (O_1193,N_14074,N_13727);
nand UO_1194 (O_1194,N_14648,N_13912);
or UO_1195 (O_1195,N_13603,N_14911);
or UO_1196 (O_1196,N_14836,N_13671);
nand UO_1197 (O_1197,N_14789,N_14232);
nand UO_1198 (O_1198,N_14434,N_14503);
nor UO_1199 (O_1199,N_13517,N_13623);
nand UO_1200 (O_1200,N_14263,N_14711);
and UO_1201 (O_1201,N_14491,N_14768);
nand UO_1202 (O_1202,N_13785,N_14479);
and UO_1203 (O_1203,N_14471,N_14890);
nor UO_1204 (O_1204,N_14401,N_13519);
and UO_1205 (O_1205,N_13514,N_14343);
or UO_1206 (O_1206,N_13528,N_14321);
nand UO_1207 (O_1207,N_14255,N_13673);
and UO_1208 (O_1208,N_14463,N_14972);
nor UO_1209 (O_1209,N_14249,N_13701);
or UO_1210 (O_1210,N_14978,N_14582);
and UO_1211 (O_1211,N_13664,N_13502);
and UO_1212 (O_1212,N_14555,N_13779);
nor UO_1213 (O_1213,N_13881,N_14925);
nor UO_1214 (O_1214,N_14466,N_14119);
nor UO_1215 (O_1215,N_14573,N_14449);
nand UO_1216 (O_1216,N_14025,N_14078);
or UO_1217 (O_1217,N_13979,N_13634);
or UO_1218 (O_1218,N_14375,N_14464);
nand UO_1219 (O_1219,N_14610,N_13671);
nand UO_1220 (O_1220,N_14496,N_14140);
nor UO_1221 (O_1221,N_14903,N_14748);
nor UO_1222 (O_1222,N_13777,N_13756);
xnor UO_1223 (O_1223,N_13849,N_13796);
and UO_1224 (O_1224,N_13514,N_13908);
and UO_1225 (O_1225,N_14724,N_13655);
and UO_1226 (O_1226,N_14735,N_14581);
nand UO_1227 (O_1227,N_14266,N_14819);
or UO_1228 (O_1228,N_14996,N_14238);
or UO_1229 (O_1229,N_13889,N_13732);
nand UO_1230 (O_1230,N_14050,N_13689);
or UO_1231 (O_1231,N_13702,N_14034);
nor UO_1232 (O_1232,N_14212,N_13907);
or UO_1233 (O_1233,N_14855,N_14578);
nand UO_1234 (O_1234,N_14962,N_14629);
nand UO_1235 (O_1235,N_14519,N_13580);
nand UO_1236 (O_1236,N_14827,N_13647);
nand UO_1237 (O_1237,N_13594,N_14870);
nand UO_1238 (O_1238,N_14485,N_14145);
or UO_1239 (O_1239,N_14247,N_13537);
nor UO_1240 (O_1240,N_13967,N_13702);
or UO_1241 (O_1241,N_14693,N_13796);
nor UO_1242 (O_1242,N_13711,N_14385);
nand UO_1243 (O_1243,N_13907,N_13584);
or UO_1244 (O_1244,N_14931,N_13663);
and UO_1245 (O_1245,N_13674,N_14631);
nand UO_1246 (O_1246,N_14915,N_14422);
nor UO_1247 (O_1247,N_14819,N_14148);
and UO_1248 (O_1248,N_13824,N_13952);
nor UO_1249 (O_1249,N_14415,N_13881);
or UO_1250 (O_1250,N_14336,N_14045);
nor UO_1251 (O_1251,N_14878,N_14339);
nor UO_1252 (O_1252,N_14343,N_14724);
nor UO_1253 (O_1253,N_14306,N_13530);
nand UO_1254 (O_1254,N_14082,N_14194);
nor UO_1255 (O_1255,N_14459,N_14315);
nor UO_1256 (O_1256,N_13726,N_14641);
nor UO_1257 (O_1257,N_13575,N_13700);
nand UO_1258 (O_1258,N_13984,N_14758);
nor UO_1259 (O_1259,N_14278,N_14806);
nand UO_1260 (O_1260,N_13989,N_14062);
and UO_1261 (O_1261,N_14872,N_14935);
nor UO_1262 (O_1262,N_13724,N_14437);
nand UO_1263 (O_1263,N_14334,N_14517);
nor UO_1264 (O_1264,N_14651,N_14559);
nor UO_1265 (O_1265,N_14788,N_14523);
nor UO_1266 (O_1266,N_14408,N_14828);
or UO_1267 (O_1267,N_14040,N_14375);
and UO_1268 (O_1268,N_14269,N_13816);
nand UO_1269 (O_1269,N_14282,N_13650);
and UO_1270 (O_1270,N_14554,N_14224);
nand UO_1271 (O_1271,N_13520,N_13552);
nor UO_1272 (O_1272,N_13545,N_14046);
nand UO_1273 (O_1273,N_13557,N_14828);
or UO_1274 (O_1274,N_14775,N_14766);
nand UO_1275 (O_1275,N_14842,N_14820);
and UO_1276 (O_1276,N_14232,N_13928);
or UO_1277 (O_1277,N_14041,N_13581);
nor UO_1278 (O_1278,N_14038,N_14486);
and UO_1279 (O_1279,N_13719,N_14320);
nor UO_1280 (O_1280,N_13936,N_14842);
nand UO_1281 (O_1281,N_14474,N_13641);
or UO_1282 (O_1282,N_14340,N_14187);
nor UO_1283 (O_1283,N_14842,N_14841);
xnor UO_1284 (O_1284,N_14304,N_14194);
nor UO_1285 (O_1285,N_13863,N_14882);
nand UO_1286 (O_1286,N_13846,N_13920);
or UO_1287 (O_1287,N_13706,N_14023);
nor UO_1288 (O_1288,N_13812,N_14970);
nand UO_1289 (O_1289,N_13876,N_14488);
xor UO_1290 (O_1290,N_14440,N_14806);
xor UO_1291 (O_1291,N_13831,N_14460);
nand UO_1292 (O_1292,N_14175,N_13698);
or UO_1293 (O_1293,N_14036,N_14946);
nand UO_1294 (O_1294,N_14903,N_14302);
and UO_1295 (O_1295,N_14509,N_13811);
nand UO_1296 (O_1296,N_14572,N_13633);
and UO_1297 (O_1297,N_13607,N_14204);
and UO_1298 (O_1298,N_14454,N_14950);
and UO_1299 (O_1299,N_14948,N_14430);
xor UO_1300 (O_1300,N_13990,N_14184);
and UO_1301 (O_1301,N_13836,N_13699);
nor UO_1302 (O_1302,N_14323,N_14836);
xor UO_1303 (O_1303,N_14585,N_14215);
or UO_1304 (O_1304,N_14985,N_14301);
nor UO_1305 (O_1305,N_14061,N_14234);
and UO_1306 (O_1306,N_13518,N_14194);
xnor UO_1307 (O_1307,N_14509,N_13952);
nor UO_1308 (O_1308,N_14770,N_14541);
xor UO_1309 (O_1309,N_14018,N_14884);
or UO_1310 (O_1310,N_14568,N_14694);
and UO_1311 (O_1311,N_14588,N_14779);
nand UO_1312 (O_1312,N_14625,N_13627);
nor UO_1313 (O_1313,N_14466,N_14631);
nand UO_1314 (O_1314,N_13642,N_14453);
and UO_1315 (O_1315,N_14225,N_14735);
xnor UO_1316 (O_1316,N_13648,N_13878);
nor UO_1317 (O_1317,N_13620,N_13667);
nor UO_1318 (O_1318,N_14051,N_14423);
nand UO_1319 (O_1319,N_14855,N_13868);
nor UO_1320 (O_1320,N_13518,N_14167);
nand UO_1321 (O_1321,N_13795,N_13835);
or UO_1322 (O_1322,N_13717,N_14621);
or UO_1323 (O_1323,N_13576,N_14403);
nor UO_1324 (O_1324,N_13790,N_13910);
or UO_1325 (O_1325,N_14478,N_13807);
or UO_1326 (O_1326,N_14344,N_14379);
nand UO_1327 (O_1327,N_13850,N_14465);
or UO_1328 (O_1328,N_14827,N_13596);
or UO_1329 (O_1329,N_14246,N_14425);
or UO_1330 (O_1330,N_14938,N_14975);
and UO_1331 (O_1331,N_14957,N_14219);
nand UO_1332 (O_1332,N_13565,N_14050);
nand UO_1333 (O_1333,N_14849,N_14588);
nand UO_1334 (O_1334,N_14061,N_13556);
and UO_1335 (O_1335,N_13606,N_13636);
nor UO_1336 (O_1336,N_14593,N_14282);
and UO_1337 (O_1337,N_13569,N_14803);
nand UO_1338 (O_1338,N_14152,N_13584);
nand UO_1339 (O_1339,N_13967,N_14951);
nor UO_1340 (O_1340,N_13833,N_14994);
or UO_1341 (O_1341,N_14391,N_14783);
nor UO_1342 (O_1342,N_14353,N_14224);
and UO_1343 (O_1343,N_14327,N_14180);
and UO_1344 (O_1344,N_14410,N_14252);
or UO_1345 (O_1345,N_13884,N_14850);
nand UO_1346 (O_1346,N_14838,N_13991);
nand UO_1347 (O_1347,N_14880,N_14372);
or UO_1348 (O_1348,N_14121,N_14872);
or UO_1349 (O_1349,N_13721,N_14618);
or UO_1350 (O_1350,N_13587,N_13884);
xnor UO_1351 (O_1351,N_14521,N_13677);
nand UO_1352 (O_1352,N_14920,N_14329);
or UO_1353 (O_1353,N_14786,N_14700);
xor UO_1354 (O_1354,N_14013,N_13950);
xor UO_1355 (O_1355,N_13852,N_14558);
nand UO_1356 (O_1356,N_13925,N_14353);
or UO_1357 (O_1357,N_14122,N_14571);
xor UO_1358 (O_1358,N_14073,N_14725);
and UO_1359 (O_1359,N_13501,N_14695);
or UO_1360 (O_1360,N_14665,N_14884);
nand UO_1361 (O_1361,N_13946,N_14011);
or UO_1362 (O_1362,N_14487,N_14746);
nand UO_1363 (O_1363,N_14817,N_14509);
xor UO_1364 (O_1364,N_13897,N_13963);
and UO_1365 (O_1365,N_14783,N_13766);
nand UO_1366 (O_1366,N_13884,N_13915);
or UO_1367 (O_1367,N_14000,N_13687);
and UO_1368 (O_1368,N_13567,N_14654);
and UO_1369 (O_1369,N_14355,N_14705);
or UO_1370 (O_1370,N_14021,N_13787);
nand UO_1371 (O_1371,N_14161,N_13552);
and UO_1372 (O_1372,N_14868,N_14766);
xnor UO_1373 (O_1373,N_14878,N_13739);
nand UO_1374 (O_1374,N_13766,N_13877);
nor UO_1375 (O_1375,N_14318,N_13634);
nor UO_1376 (O_1376,N_14400,N_13736);
nand UO_1377 (O_1377,N_14539,N_13819);
xnor UO_1378 (O_1378,N_14267,N_13830);
nand UO_1379 (O_1379,N_13712,N_14338);
nand UO_1380 (O_1380,N_14431,N_13833);
and UO_1381 (O_1381,N_14719,N_13839);
nand UO_1382 (O_1382,N_13662,N_13797);
or UO_1383 (O_1383,N_14885,N_13605);
nor UO_1384 (O_1384,N_14851,N_13736);
nor UO_1385 (O_1385,N_13764,N_14456);
nand UO_1386 (O_1386,N_14837,N_14068);
xor UO_1387 (O_1387,N_14197,N_14975);
nor UO_1388 (O_1388,N_13522,N_14298);
or UO_1389 (O_1389,N_14664,N_14319);
and UO_1390 (O_1390,N_13523,N_13870);
nor UO_1391 (O_1391,N_14200,N_14290);
or UO_1392 (O_1392,N_14376,N_14986);
nand UO_1393 (O_1393,N_14277,N_14686);
nand UO_1394 (O_1394,N_14149,N_14643);
or UO_1395 (O_1395,N_14838,N_14986);
and UO_1396 (O_1396,N_14511,N_14921);
nand UO_1397 (O_1397,N_13604,N_14866);
or UO_1398 (O_1398,N_14167,N_14718);
and UO_1399 (O_1399,N_13992,N_14895);
or UO_1400 (O_1400,N_13779,N_14904);
or UO_1401 (O_1401,N_14584,N_14512);
nand UO_1402 (O_1402,N_14175,N_14522);
and UO_1403 (O_1403,N_13943,N_13552);
xnor UO_1404 (O_1404,N_13925,N_14678);
nor UO_1405 (O_1405,N_13770,N_13900);
or UO_1406 (O_1406,N_13605,N_13550);
nor UO_1407 (O_1407,N_13506,N_14438);
nand UO_1408 (O_1408,N_14506,N_13756);
and UO_1409 (O_1409,N_13803,N_13604);
nand UO_1410 (O_1410,N_14198,N_13689);
or UO_1411 (O_1411,N_14289,N_13646);
and UO_1412 (O_1412,N_14335,N_14867);
nand UO_1413 (O_1413,N_13803,N_13963);
and UO_1414 (O_1414,N_13646,N_13710);
nand UO_1415 (O_1415,N_14784,N_14675);
and UO_1416 (O_1416,N_14642,N_13883);
xor UO_1417 (O_1417,N_14969,N_14708);
nor UO_1418 (O_1418,N_13581,N_13737);
xor UO_1419 (O_1419,N_13516,N_14398);
or UO_1420 (O_1420,N_14878,N_13774);
nor UO_1421 (O_1421,N_13567,N_13588);
nor UO_1422 (O_1422,N_13640,N_14508);
nor UO_1423 (O_1423,N_14850,N_14621);
nand UO_1424 (O_1424,N_14417,N_14311);
or UO_1425 (O_1425,N_14963,N_14472);
nand UO_1426 (O_1426,N_14221,N_14326);
xnor UO_1427 (O_1427,N_14022,N_14302);
or UO_1428 (O_1428,N_14751,N_14302);
nand UO_1429 (O_1429,N_14694,N_14522);
and UO_1430 (O_1430,N_14326,N_14668);
and UO_1431 (O_1431,N_13733,N_13790);
nor UO_1432 (O_1432,N_14987,N_14115);
or UO_1433 (O_1433,N_14829,N_13757);
xnor UO_1434 (O_1434,N_14901,N_14013);
or UO_1435 (O_1435,N_14996,N_13868);
nor UO_1436 (O_1436,N_14181,N_14485);
nor UO_1437 (O_1437,N_14953,N_13954);
and UO_1438 (O_1438,N_14476,N_14993);
nor UO_1439 (O_1439,N_13680,N_13684);
nand UO_1440 (O_1440,N_14885,N_14172);
or UO_1441 (O_1441,N_14335,N_14600);
and UO_1442 (O_1442,N_13588,N_14236);
and UO_1443 (O_1443,N_14688,N_14339);
nand UO_1444 (O_1444,N_14455,N_13756);
xor UO_1445 (O_1445,N_13957,N_14722);
nor UO_1446 (O_1446,N_13589,N_14932);
and UO_1447 (O_1447,N_14311,N_13897);
nor UO_1448 (O_1448,N_14854,N_14746);
nor UO_1449 (O_1449,N_13538,N_14468);
nor UO_1450 (O_1450,N_14139,N_14306);
xnor UO_1451 (O_1451,N_14358,N_14952);
or UO_1452 (O_1452,N_14466,N_14943);
xnor UO_1453 (O_1453,N_14727,N_14854);
or UO_1454 (O_1454,N_14822,N_14142);
and UO_1455 (O_1455,N_14142,N_14062);
nand UO_1456 (O_1456,N_14274,N_13998);
and UO_1457 (O_1457,N_14103,N_14232);
and UO_1458 (O_1458,N_14903,N_14614);
nand UO_1459 (O_1459,N_14428,N_14605);
nand UO_1460 (O_1460,N_14430,N_13844);
and UO_1461 (O_1461,N_13509,N_14183);
xor UO_1462 (O_1462,N_14316,N_14420);
nor UO_1463 (O_1463,N_14035,N_13804);
nand UO_1464 (O_1464,N_14067,N_14191);
nand UO_1465 (O_1465,N_14761,N_14714);
or UO_1466 (O_1466,N_14732,N_13874);
nor UO_1467 (O_1467,N_13612,N_14913);
and UO_1468 (O_1468,N_13653,N_13957);
or UO_1469 (O_1469,N_14522,N_14184);
nor UO_1470 (O_1470,N_14947,N_13724);
nor UO_1471 (O_1471,N_14796,N_14941);
xor UO_1472 (O_1472,N_13786,N_13549);
nand UO_1473 (O_1473,N_14773,N_14171);
nand UO_1474 (O_1474,N_14852,N_14982);
or UO_1475 (O_1475,N_14683,N_14699);
xnor UO_1476 (O_1476,N_14400,N_14918);
and UO_1477 (O_1477,N_14880,N_14227);
and UO_1478 (O_1478,N_13977,N_14035);
or UO_1479 (O_1479,N_14645,N_14764);
nand UO_1480 (O_1480,N_14664,N_14924);
and UO_1481 (O_1481,N_14623,N_13592);
nand UO_1482 (O_1482,N_13833,N_14587);
nor UO_1483 (O_1483,N_14110,N_14297);
nand UO_1484 (O_1484,N_14228,N_14546);
or UO_1485 (O_1485,N_13900,N_14824);
nor UO_1486 (O_1486,N_14876,N_13825);
nand UO_1487 (O_1487,N_14325,N_14447);
or UO_1488 (O_1488,N_14266,N_13645);
or UO_1489 (O_1489,N_13554,N_13926);
or UO_1490 (O_1490,N_13982,N_13528);
or UO_1491 (O_1491,N_13854,N_13949);
xor UO_1492 (O_1492,N_14519,N_14029);
or UO_1493 (O_1493,N_14276,N_14363);
nor UO_1494 (O_1494,N_13861,N_13681);
and UO_1495 (O_1495,N_13716,N_13625);
nand UO_1496 (O_1496,N_13952,N_14662);
or UO_1497 (O_1497,N_14741,N_14572);
nor UO_1498 (O_1498,N_13807,N_14330);
or UO_1499 (O_1499,N_13938,N_14657);
and UO_1500 (O_1500,N_13909,N_14450);
or UO_1501 (O_1501,N_14282,N_13750);
xor UO_1502 (O_1502,N_14159,N_14882);
xor UO_1503 (O_1503,N_14912,N_14406);
nand UO_1504 (O_1504,N_14079,N_14405);
nand UO_1505 (O_1505,N_14161,N_13530);
xnor UO_1506 (O_1506,N_14388,N_13593);
nor UO_1507 (O_1507,N_14699,N_14304);
or UO_1508 (O_1508,N_14600,N_14380);
nor UO_1509 (O_1509,N_14988,N_13622);
and UO_1510 (O_1510,N_14387,N_14660);
nand UO_1511 (O_1511,N_13622,N_13956);
nor UO_1512 (O_1512,N_14457,N_13901);
xor UO_1513 (O_1513,N_14482,N_14046);
xor UO_1514 (O_1514,N_13744,N_14214);
nand UO_1515 (O_1515,N_14426,N_14959);
or UO_1516 (O_1516,N_13844,N_13933);
nand UO_1517 (O_1517,N_13982,N_14769);
xor UO_1518 (O_1518,N_13649,N_13768);
nor UO_1519 (O_1519,N_13560,N_13898);
or UO_1520 (O_1520,N_14085,N_14595);
and UO_1521 (O_1521,N_13593,N_13935);
xnor UO_1522 (O_1522,N_14537,N_14496);
or UO_1523 (O_1523,N_14072,N_14218);
and UO_1524 (O_1524,N_13763,N_14262);
and UO_1525 (O_1525,N_14433,N_14323);
or UO_1526 (O_1526,N_13665,N_14491);
or UO_1527 (O_1527,N_13555,N_14619);
nand UO_1528 (O_1528,N_14937,N_13941);
and UO_1529 (O_1529,N_14856,N_13564);
nand UO_1530 (O_1530,N_14708,N_14798);
nand UO_1531 (O_1531,N_14313,N_14352);
nor UO_1532 (O_1532,N_14914,N_14415);
or UO_1533 (O_1533,N_13533,N_13852);
nand UO_1534 (O_1534,N_14527,N_14916);
or UO_1535 (O_1535,N_14670,N_14106);
or UO_1536 (O_1536,N_14154,N_13870);
nor UO_1537 (O_1537,N_14595,N_14658);
nor UO_1538 (O_1538,N_14787,N_13743);
or UO_1539 (O_1539,N_14393,N_14062);
nand UO_1540 (O_1540,N_14024,N_14828);
nor UO_1541 (O_1541,N_14407,N_14353);
nor UO_1542 (O_1542,N_14450,N_14790);
nand UO_1543 (O_1543,N_13937,N_13718);
or UO_1544 (O_1544,N_14390,N_14374);
nor UO_1545 (O_1545,N_14692,N_14996);
or UO_1546 (O_1546,N_14873,N_14914);
and UO_1547 (O_1547,N_14439,N_13981);
and UO_1548 (O_1548,N_14826,N_14470);
and UO_1549 (O_1549,N_14723,N_13545);
nor UO_1550 (O_1550,N_14723,N_13653);
and UO_1551 (O_1551,N_14851,N_14169);
nor UO_1552 (O_1552,N_14968,N_14897);
nand UO_1553 (O_1553,N_14978,N_14955);
nand UO_1554 (O_1554,N_14927,N_14246);
xnor UO_1555 (O_1555,N_14776,N_14683);
and UO_1556 (O_1556,N_14618,N_14050);
nand UO_1557 (O_1557,N_14483,N_14298);
nor UO_1558 (O_1558,N_14241,N_14894);
nor UO_1559 (O_1559,N_13763,N_13740);
xnor UO_1560 (O_1560,N_13678,N_13983);
or UO_1561 (O_1561,N_13788,N_14112);
and UO_1562 (O_1562,N_14495,N_13964);
and UO_1563 (O_1563,N_14559,N_14428);
and UO_1564 (O_1564,N_14550,N_13649);
nor UO_1565 (O_1565,N_14984,N_14820);
and UO_1566 (O_1566,N_14694,N_14331);
nand UO_1567 (O_1567,N_14001,N_13536);
nand UO_1568 (O_1568,N_14337,N_13659);
and UO_1569 (O_1569,N_14647,N_13569);
or UO_1570 (O_1570,N_13947,N_14531);
nand UO_1571 (O_1571,N_14498,N_13919);
nor UO_1572 (O_1572,N_14007,N_14157);
nor UO_1573 (O_1573,N_13980,N_14740);
or UO_1574 (O_1574,N_14088,N_14219);
xor UO_1575 (O_1575,N_14442,N_14603);
nand UO_1576 (O_1576,N_13891,N_13970);
nor UO_1577 (O_1577,N_13807,N_14741);
nor UO_1578 (O_1578,N_14030,N_13734);
or UO_1579 (O_1579,N_14625,N_14463);
xor UO_1580 (O_1580,N_14840,N_14497);
nand UO_1581 (O_1581,N_13682,N_13668);
nor UO_1582 (O_1582,N_14087,N_13779);
or UO_1583 (O_1583,N_14182,N_14279);
and UO_1584 (O_1584,N_14642,N_14486);
or UO_1585 (O_1585,N_14781,N_14471);
nand UO_1586 (O_1586,N_14572,N_13549);
and UO_1587 (O_1587,N_13922,N_14574);
nor UO_1588 (O_1588,N_13802,N_14697);
or UO_1589 (O_1589,N_14056,N_13963);
xnor UO_1590 (O_1590,N_13588,N_13517);
nand UO_1591 (O_1591,N_14063,N_14460);
and UO_1592 (O_1592,N_13844,N_14492);
nor UO_1593 (O_1593,N_14051,N_13969);
and UO_1594 (O_1594,N_13946,N_14665);
or UO_1595 (O_1595,N_14942,N_14488);
nand UO_1596 (O_1596,N_14195,N_13671);
xor UO_1597 (O_1597,N_14246,N_13597);
and UO_1598 (O_1598,N_14217,N_14913);
xnor UO_1599 (O_1599,N_13928,N_14459);
nor UO_1600 (O_1600,N_13555,N_14465);
and UO_1601 (O_1601,N_14972,N_14670);
nor UO_1602 (O_1602,N_13978,N_14405);
or UO_1603 (O_1603,N_13698,N_14140);
or UO_1604 (O_1604,N_13562,N_14889);
nand UO_1605 (O_1605,N_13539,N_14417);
nand UO_1606 (O_1606,N_14770,N_13522);
nor UO_1607 (O_1607,N_13661,N_14473);
and UO_1608 (O_1608,N_13892,N_13638);
or UO_1609 (O_1609,N_13783,N_13995);
and UO_1610 (O_1610,N_13810,N_14090);
nand UO_1611 (O_1611,N_14879,N_14068);
nor UO_1612 (O_1612,N_14369,N_13644);
nor UO_1613 (O_1613,N_13590,N_14436);
and UO_1614 (O_1614,N_13773,N_14163);
and UO_1615 (O_1615,N_14371,N_14246);
or UO_1616 (O_1616,N_14885,N_13759);
or UO_1617 (O_1617,N_14939,N_14264);
nor UO_1618 (O_1618,N_14080,N_14264);
and UO_1619 (O_1619,N_14802,N_14494);
xor UO_1620 (O_1620,N_13547,N_14235);
nor UO_1621 (O_1621,N_14720,N_14865);
nor UO_1622 (O_1622,N_13527,N_14254);
nor UO_1623 (O_1623,N_14172,N_14871);
and UO_1624 (O_1624,N_14270,N_14189);
and UO_1625 (O_1625,N_14456,N_14371);
and UO_1626 (O_1626,N_13658,N_14941);
and UO_1627 (O_1627,N_14376,N_14958);
nor UO_1628 (O_1628,N_14652,N_13813);
xor UO_1629 (O_1629,N_14090,N_13538);
nand UO_1630 (O_1630,N_14713,N_14908);
nor UO_1631 (O_1631,N_14468,N_14963);
nor UO_1632 (O_1632,N_14623,N_14513);
nand UO_1633 (O_1633,N_13936,N_14987);
nor UO_1634 (O_1634,N_14578,N_14183);
or UO_1635 (O_1635,N_14422,N_14745);
xnor UO_1636 (O_1636,N_13716,N_14088);
nand UO_1637 (O_1637,N_14938,N_14097);
nand UO_1638 (O_1638,N_13627,N_14896);
or UO_1639 (O_1639,N_14467,N_14409);
xor UO_1640 (O_1640,N_13939,N_14550);
nor UO_1641 (O_1641,N_14746,N_13522);
nor UO_1642 (O_1642,N_14242,N_14126);
and UO_1643 (O_1643,N_14207,N_13552);
nor UO_1644 (O_1644,N_14734,N_14233);
and UO_1645 (O_1645,N_14685,N_13630);
nor UO_1646 (O_1646,N_13681,N_13951);
xor UO_1647 (O_1647,N_13900,N_14065);
and UO_1648 (O_1648,N_13794,N_14598);
nand UO_1649 (O_1649,N_13789,N_13921);
or UO_1650 (O_1650,N_14717,N_14104);
or UO_1651 (O_1651,N_14191,N_13896);
nor UO_1652 (O_1652,N_14796,N_14275);
nand UO_1653 (O_1653,N_13593,N_13561);
or UO_1654 (O_1654,N_13850,N_14551);
nor UO_1655 (O_1655,N_13652,N_13867);
nor UO_1656 (O_1656,N_14901,N_13536);
and UO_1657 (O_1657,N_14551,N_14309);
nand UO_1658 (O_1658,N_14756,N_13766);
nand UO_1659 (O_1659,N_14236,N_13887);
nand UO_1660 (O_1660,N_14198,N_13751);
or UO_1661 (O_1661,N_13869,N_14949);
or UO_1662 (O_1662,N_13840,N_13525);
nand UO_1663 (O_1663,N_14759,N_14161);
or UO_1664 (O_1664,N_13735,N_13670);
or UO_1665 (O_1665,N_14318,N_14826);
nor UO_1666 (O_1666,N_14785,N_14786);
nand UO_1667 (O_1667,N_13797,N_14848);
or UO_1668 (O_1668,N_13714,N_14768);
or UO_1669 (O_1669,N_14641,N_14447);
or UO_1670 (O_1670,N_14063,N_14038);
nor UO_1671 (O_1671,N_14409,N_14555);
and UO_1672 (O_1672,N_13933,N_13646);
xor UO_1673 (O_1673,N_14673,N_14901);
xnor UO_1674 (O_1674,N_14836,N_14358);
nor UO_1675 (O_1675,N_14790,N_14335);
nand UO_1676 (O_1676,N_14979,N_14234);
xor UO_1677 (O_1677,N_14867,N_14974);
and UO_1678 (O_1678,N_13835,N_14607);
and UO_1679 (O_1679,N_14141,N_13645);
nand UO_1680 (O_1680,N_14510,N_14173);
and UO_1681 (O_1681,N_14658,N_14779);
xor UO_1682 (O_1682,N_14116,N_14665);
or UO_1683 (O_1683,N_14960,N_13570);
or UO_1684 (O_1684,N_14887,N_14057);
nand UO_1685 (O_1685,N_14821,N_14037);
nor UO_1686 (O_1686,N_13933,N_13895);
xor UO_1687 (O_1687,N_14158,N_13742);
nand UO_1688 (O_1688,N_13780,N_13622);
or UO_1689 (O_1689,N_13934,N_14955);
nand UO_1690 (O_1690,N_13864,N_14972);
nor UO_1691 (O_1691,N_13729,N_14092);
and UO_1692 (O_1692,N_14378,N_14458);
nand UO_1693 (O_1693,N_14548,N_13777);
nand UO_1694 (O_1694,N_14543,N_14891);
and UO_1695 (O_1695,N_14984,N_13748);
nor UO_1696 (O_1696,N_13729,N_14401);
or UO_1697 (O_1697,N_14432,N_14332);
nand UO_1698 (O_1698,N_14136,N_13728);
or UO_1699 (O_1699,N_13661,N_14765);
or UO_1700 (O_1700,N_14120,N_14376);
xnor UO_1701 (O_1701,N_13941,N_13575);
xnor UO_1702 (O_1702,N_14755,N_14436);
and UO_1703 (O_1703,N_14888,N_13802);
and UO_1704 (O_1704,N_14239,N_13711);
and UO_1705 (O_1705,N_13891,N_14519);
and UO_1706 (O_1706,N_14623,N_14536);
nand UO_1707 (O_1707,N_13979,N_14735);
and UO_1708 (O_1708,N_14780,N_14406);
or UO_1709 (O_1709,N_14946,N_14210);
nand UO_1710 (O_1710,N_14772,N_14022);
or UO_1711 (O_1711,N_13757,N_13582);
nand UO_1712 (O_1712,N_14960,N_14757);
xor UO_1713 (O_1713,N_13756,N_14301);
nor UO_1714 (O_1714,N_14214,N_14913);
and UO_1715 (O_1715,N_13501,N_13931);
nand UO_1716 (O_1716,N_14904,N_13835);
and UO_1717 (O_1717,N_14864,N_13572);
and UO_1718 (O_1718,N_14516,N_14068);
or UO_1719 (O_1719,N_14279,N_13521);
or UO_1720 (O_1720,N_14243,N_13917);
and UO_1721 (O_1721,N_13692,N_14386);
nand UO_1722 (O_1722,N_14343,N_14799);
xnor UO_1723 (O_1723,N_14817,N_14057);
or UO_1724 (O_1724,N_13584,N_13703);
nor UO_1725 (O_1725,N_14108,N_13829);
and UO_1726 (O_1726,N_14031,N_14687);
xnor UO_1727 (O_1727,N_13671,N_13884);
nand UO_1728 (O_1728,N_13822,N_14509);
and UO_1729 (O_1729,N_13839,N_13702);
nor UO_1730 (O_1730,N_13802,N_14614);
or UO_1731 (O_1731,N_14587,N_13537);
or UO_1732 (O_1732,N_13814,N_14479);
and UO_1733 (O_1733,N_14954,N_14524);
and UO_1734 (O_1734,N_13636,N_14784);
nand UO_1735 (O_1735,N_13894,N_13916);
nor UO_1736 (O_1736,N_14482,N_14543);
and UO_1737 (O_1737,N_14719,N_14467);
and UO_1738 (O_1738,N_14869,N_14360);
or UO_1739 (O_1739,N_14524,N_14078);
nor UO_1740 (O_1740,N_13669,N_14850);
nand UO_1741 (O_1741,N_14766,N_13555);
and UO_1742 (O_1742,N_14385,N_14501);
nor UO_1743 (O_1743,N_13813,N_14481);
xor UO_1744 (O_1744,N_14135,N_14459);
and UO_1745 (O_1745,N_13615,N_14836);
or UO_1746 (O_1746,N_14085,N_14858);
or UO_1747 (O_1747,N_14333,N_14433);
nor UO_1748 (O_1748,N_13657,N_14228);
and UO_1749 (O_1749,N_14401,N_14553);
nand UO_1750 (O_1750,N_14762,N_14421);
nand UO_1751 (O_1751,N_14602,N_14284);
nand UO_1752 (O_1752,N_14833,N_14127);
and UO_1753 (O_1753,N_14677,N_14516);
nor UO_1754 (O_1754,N_14594,N_14420);
nor UO_1755 (O_1755,N_13628,N_14789);
nand UO_1756 (O_1756,N_14759,N_13869);
nand UO_1757 (O_1757,N_14722,N_14906);
or UO_1758 (O_1758,N_14854,N_14086);
and UO_1759 (O_1759,N_14777,N_14963);
nand UO_1760 (O_1760,N_14148,N_13988);
nor UO_1761 (O_1761,N_13808,N_14146);
nor UO_1762 (O_1762,N_14892,N_14508);
or UO_1763 (O_1763,N_14863,N_14965);
nor UO_1764 (O_1764,N_14804,N_14611);
xor UO_1765 (O_1765,N_14592,N_14279);
nand UO_1766 (O_1766,N_14548,N_13522);
or UO_1767 (O_1767,N_14796,N_14922);
or UO_1768 (O_1768,N_14807,N_14666);
xnor UO_1769 (O_1769,N_14699,N_14277);
or UO_1770 (O_1770,N_13947,N_14793);
nor UO_1771 (O_1771,N_14617,N_14731);
or UO_1772 (O_1772,N_14949,N_13888);
nand UO_1773 (O_1773,N_14597,N_13895);
and UO_1774 (O_1774,N_14185,N_14827);
nand UO_1775 (O_1775,N_13601,N_13897);
and UO_1776 (O_1776,N_14221,N_14868);
nand UO_1777 (O_1777,N_14338,N_14335);
and UO_1778 (O_1778,N_14316,N_14952);
nand UO_1779 (O_1779,N_14787,N_13976);
and UO_1780 (O_1780,N_13821,N_14645);
or UO_1781 (O_1781,N_14179,N_14419);
nor UO_1782 (O_1782,N_14882,N_14051);
and UO_1783 (O_1783,N_14831,N_14350);
xor UO_1784 (O_1784,N_14368,N_13668);
nand UO_1785 (O_1785,N_14032,N_14682);
and UO_1786 (O_1786,N_13644,N_14057);
and UO_1787 (O_1787,N_14759,N_14844);
and UO_1788 (O_1788,N_14083,N_13816);
nand UO_1789 (O_1789,N_13514,N_13594);
nor UO_1790 (O_1790,N_14553,N_13699);
nand UO_1791 (O_1791,N_14007,N_14008);
or UO_1792 (O_1792,N_14789,N_14032);
or UO_1793 (O_1793,N_14682,N_14200);
or UO_1794 (O_1794,N_13847,N_13974);
or UO_1795 (O_1795,N_14021,N_13779);
nor UO_1796 (O_1796,N_14381,N_14361);
and UO_1797 (O_1797,N_13502,N_14718);
or UO_1798 (O_1798,N_14907,N_13691);
and UO_1799 (O_1799,N_13580,N_14953);
nor UO_1800 (O_1800,N_13987,N_14397);
nand UO_1801 (O_1801,N_14095,N_14364);
nor UO_1802 (O_1802,N_14889,N_14936);
nor UO_1803 (O_1803,N_14810,N_14930);
nand UO_1804 (O_1804,N_14549,N_14931);
nand UO_1805 (O_1805,N_13587,N_13691);
or UO_1806 (O_1806,N_14584,N_14573);
xor UO_1807 (O_1807,N_13503,N_14434);
xor UO_1808 (O_1808,N_14290,N_14296);
nor UO_1809 (O_1809,N_13775,N_14101);
and UO_1810 (O_1810,N_13521,N_14484);
nor UO_1811 (O_1811,N_14245,N_14089);
or UO_1812 (O_1812,N_14620,N_14734);
and UO_1813 (O_1813,N_13657,N_14749);
and UO_1814 (O_1814,N_14955,N_14525);
and UO_1815 (O_1815,N_14955,N_13687);
and UO_1816 (O_1816,N_14789,N_14637);
and UO_1817 (O_1817,N_13697,N_13843);
and UO_1818 (O_1818,N_14407,N_13849);
nor UO_1819 (O_1819,N_14893,N_14925);
nand UO_1820 (O_1820,N_14773,N_14744);
nor UO_1821 (O_1821,N_13914,N_14495);
or UO_1822 (O_1822,N_14937,N_14421);
nand UO_1823 (O_1823,N_13690,N_14283);
nor UO_1824 (O_1824,N_14428,N_14274);
xor UO_1825 (O_1825,N_14563,N_14606);
nand UO_1826 (O_1826,N_14086,N_13533);
nor UO_1827 (O_1827,N_14595,N_14520);
and UO_1828 (O_1828,N_14289,N_14975);
and UO_1829 (O_1829,N_13552,N_13813);
nand UO_1830 (O_1830,N_14192,N_14389);
nand UO_1831 (O_1831,N_14160,N_14479);
nand UO_1832 (O_1832,N_13522,N_14902);
or UO_1833 (O_1833,N_13919,N_14774);
and UO_1834 (O_1834,N_14098,N_13956);
or UO_1835 (O_1835,N_14078,N_13845);
nor UO_1836 (O_1836,N_13821,N_13854);
nor UO_1837 (O_1837,N_14528,N_14229);
and UO_1838 (O_1838,N_14738,N_14383);
or UO_1839 (O_1839,N_13820,N_13856);
nand UO_1840 (O_1840,N_14717,N_13509);
nor UO_1841 (O_1841,N_13581,N_14653);
nand UO_1842 (O_1842,N_14686,N_14690);
and UO_1843 (O_1843,N_13994,N_13947);
or UO_1844 (O_1844,N_13816,N_14333);
nand UO_1845 (O_1845,N_13609,N_14975);
xor UO_1846 (O_1846,N_13951,N_13567);
nand UO_1847 (O_1847,N_14103,N_14138);
nand UO_1848 (O_1848,N_13781,N_13752);
nor UO_1849 (O_1849,N_14162,N_13729);
and UO_1850 (O_1850,N_14857,N_13827);
nor UO_1851 (O_1851,N_14711,N_14101);
nor UO_1852 (O_1852,N_13516,N_14400);
or UO_1853 (O_1853,N_14717,N_14289);
or UO_1854 (O_1854,N_13833,N_13537);
nand UO_1855 (O_1855,N_13948,N_14390);
xnor UO_1856 (O_1856,N_13806,N_13738);
and UO_1857 (O_1857,N_14690,N_13980);
xnor UO_1858 (O_1858,N_14600,N_14256);
nor UO_1859 (O_1859,N_14631,N_14319);
and UO_1860 (O_1860,N_14385,N_14079);
nand UO_1861 (O_1861,N_14750,N_14474);
nand UO_1862 (O_1862,N_14557,N_14628);
nand UO_1863 (O_1863,N_14309,N_14829);
nor UO_1864 (O_1864,N_13933,N_13617);
or UO_1865 (O_1865,N_14878,N_14468);
or UO_1866 (O_1866,N_14197,N_14021);
nor UO_1867 (O_1867,N_14829,N_13687);
nand UO_1868 (O_1868,N_13791,N_13776);
nand UO_1869 (O_1869,N_13708,N_14044);
or UO_1870 (O_1870,N_14434,N_14500);
or UO_1871 (O_1871,N_13648,N_14745);
or UO_1872 (O_1872,N_14571,N_14812);
nand UO_1873 (O_1873,N_14567,N_14613);
nor UO_1874 (O_1874,N_13708,N_14067);
nand UO_1875 (O_1875,N_13734,N_14779);
and UO_1876 (O_1876,N_14295,N_14860);
and UO_1877 (O_1877,N_14634,N_13558);
nand UO_1878 (O_1878,N_14014,N_14879);
and UO_1879 (O_1879,N_14763,N_13536);
xnor UO_1880 (O_1880,N_14244,N_13736);
xnor UO_1881 (O_1881,N_14207,N_13781);
nor UO_1882 (O_1882,N_13672,N_14984);
nand UO_1883 (O_1883,N_14810,N_14827);
and UO_1884 (O_1884,N_14557,N_13805);
nor UO_1885 (O_1885,N_14614,N_13670);
xnor UO_1886 (O_1886,N_14072,N_14843);
or UO_1887 (O_1887,N_14319,N_14787);
nor UO_1888 (O_1888,N_14465,N_14367);
or UO_1889 (O_1889,N_13747,N_13880);
nor UO_1890 (O_1890,N_13659,N_13803);
and UO_1891 (O_1891,N_14209,N_13838);
nand UO_1892 (O_1892,N_14577,N_14432);
or UO_1893 (O_1893,N_14604,N_14712);
nand UO_1894 (O_1894,N_14291,N_14183);
nand UO_1895 (O_1895,N_14909,N_14116);
and UO_1896 (O_1896,N_14311,N_14744);
or UO_1897 (O_1897,N_14106,N_13821);
and UO_1898 (O_1898,N_13830,N_13509);
and UO_1899 (O_1899,N_14544,N_14236);
and UO_1900 (O_1900,N_14946,N_14814);
nand UO_1901 (O_1901,N_14656,N_14830);
nor UO_1902 (O_1902,N_13549,N_13953);
or UO_1903 (O_1903,N_14071,N_14755);
and UO_1904 (O_1904,N_14658,N_14107);
xor UO_1905 (O_1905,N_13920,N_14895);
nand UO_1906 (O_1906,N_14402,N_14005);
xor UO_1907 (O_1907,N_14025,N_14595);
and UO_1908 (O_1908,N_14043,N_13751);
and UO_1909 (O_1909,N_13798,N_14841);
nor UO_1910 (O_1910,N_14778,N_14142);
nand UO_1911 (O_1911,N_13970,N_14577);
nor UO_1912 (O_1912,N_14342,N_13805);
nor UO_1913 (O_1913,N_14656,N_14707);
and UO_1914 (O_1914,N_13951,N_13701);
nor UO_1915 (O_1915,N_14000,N_14543);
nor UO_1916 (O_1916,N_14888,N_14935);
or UO_1917 (O_1917,N_14288,N_13690);
xnor UO_1918 (O_1918,N_13841,N_14963);
or UO_1919 (O_1919,N_14706,N_14646);
and UO_1920 (O_1920,N_13689,N_14373);
nand UO_1921 (O_1921,N_14598,N_13667);
nand UO_1922 (O_1922,N_14902,N_14224);
nor UO_1923 (O_1923,N_14217,N_14476);
nor UO_1924 (O_1924,N_13642,N_14701);
or UO_1925 (O_1925,N_14939,N_13792);
or UO_1926 (O_1926,N_14781,N_13878);
nor UO_1927 (O_1927,N_14693,N_14835);
or UO_1928 (O_1928,N_13749,N_14373);
and UO_1929 (O_1929,N_13606,N_14690);
and UO_1930 (O_1930,N_14144,N_14354);
nor UO_1931 (O_1931,N_14204,N_14002);
nand UO_1932 (O_1932,N_14874,N_13919);
or UO_1933 (O_1933,N_14792,N_14427);
and UO_1934 (O_1934,N_14848,N_14903);
nor UO_1935 (O_1935,N_14864,N_14524);
nand UO_1936 (O_1936,N_14461,N_14873);
nor UO_1937 (O_1937,N_14498,N_14196);
nor UO_1938 (O_1938,N_14233,N_14489);
and UO_1939 (O_1939,N_14663,N_14904);
nand UO_1940 (O_1940,N_14841,N_13887);
and UO_1941 (O_1941,N_14718,N_13890);
nand UO_1942 (O_1942,N_13900,N_13659);
nand UO_1943 (O_1943,N_13663,N_14122);
nand UO_1944 (O_1944,N_14140,N_13714);
nor UO_1945 (O_1945,N_14093,N_14657);
or UO_1946 (O_1946,N_14012,N_14991);
or UO_1947 (O_1947,N_14928,N_13929);
nor UO_1948 (O_1948,N_13629,N_14425);
nand UO_1949 (O_1949,N_14512,N_14884);
or UO_1950 (O_1950,N_14541,N_13501);
or UO_1951 (O_1951,N_13744,N_14351);
nor UO_1952 (O_1952,N_13649,N_14277);
nor UO_1953 (O_1953,N_14621,N_13613);
or UO_1954 (O_1954,N_14492,N_14281);
nor UO_1955 (O_1955,N_14229,N_13673);
nor UO_1956 (O_1956,N_13917,N_13747);
and UO_1957 (O_1957,N_14505,N_14007);
nor UO_1958 (O_1958,N_14164,N_13902);
nor UO_1959 (O_1959,N_14073,N_14528);
nand UO_1960 (O_1960,N_14400,N_14602);
nor UO_1961 (O_1961,N_13951,N_14930);
and UO_1962 (O_1962,N_13985,N_14855);
or UO_1963 (O_1963,N_14107,N_13989);
and UO_1964 (O_1964,N_13898,N_14726);
or UO_1965 (O_1965,N_14125,N_14213);
and UO_1966 (O_1966,N_13781,N_14742);
nand UO_1967 (O_1967,N_14936,N_14949);
or UO_1968 (O_1968,N_14317,N_14184);
nor UO_1969 (O_1969,N_13873,N_14220);
or UO_1970 (O_1970,N_14337,N_14914);
and UO_1971 (O_1971,N_13958,N_14599);
and UO_1972 (O_1972,N_14590,N_14532);
and UO_1973 (O_1973,N_14200,N_14704);
and UO_1974 (O_1974,N_13972,N_14714);
or UO_1975 (O_1975,N_14723,N_13977);
and UO_1976 (O_1976,N_14402,N_14930);
or UO_1977 (O_1977,N_13670,N_14256);
nor UO_1978 (O_1978,N_14920,N_14193);
and UO_1979 (O_1979,N_13700,N_13710);
and UO_1980 (O_1980,N_14038,N_14365);
nand UO_1981 (O_1981,N_13588,N_14097);
xnor UO_1982 (O_1982,N_13602,N_14155);
and UO_1983 (O_1983,N_14974,N_14860);
and UO_1984 (O_1984,N_14915,N_14617);
and UO_1985 (O_1985,N_14333,N_13613);
xor UO_1986 (O_1986,N_14796,N_14220);
nor UO_1987 (O_1987,N_14760,N_13587);
or UO_1988 (O_1988,N_14084,N_14442);
nand UO_1989 (O_1989,N_13789,N_13950);
or UO_1990 (O_1990,N_13523,N_13815);
nor UO_1991 (O_1991,N_14994,N_14765);
and UO_1992 (O_1992,N_14747,N_13567);
or UO_1993 (O_1993,N_14319,N_14399);
nand UO_1994 (O_1994,N_14208,N_14983);
and UO_1995 (O_1995,N_14559,N_14811);
nand UO_1996 (O_1996,N_14338,N_13671);
or UO_1997 (O_1997,N_14884,N_13739);
or UO_1998 (O_1998,N_13992,N_14414);
xor UO_1999 (O_1999,N_14477,N_14104);
endmodule