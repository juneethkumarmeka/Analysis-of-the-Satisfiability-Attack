module basic_2000_20000_2500_100_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1734,In_1609);
and U1 (N_1,In_1404,In_2);
and U2 (N_2,In_523,In_520);
or U3 (N_3,In_880,In_917);
or U4 (N_4,In_1464,In_668);
or U5 (N_5,In_1361,In_40);
and U6 (N_6,In_1653,In_1661);
xnor U7 (N_7,In_255,In_1953);
and U8 (N_8,In_715,In_1075);
nand U9 (N_9,In_103,In_406);
xor U10 (N_10,In_1593,In_1660);
nand U11 (N_11,In_1515,In_1927);
or U12 (N_12,In_1316,In_1973);
nor U13 (N_13,In_730,In_979);
xnor U14 (N_14,In_1360,In_345);
and U15 (N_15,In_1638,In_1039);
nor U16 (N_16,In_1059,In_497);
xor U17 (N_17,In_1477,In_450);
xor U18 (N_18,In_1233,In_618);
or U19 (N_19,In_667,In_813);
or U20 (N_20,In_1824,In_1339);
nor U21 (N_21,In_1941,In_1952);
xnor U22 (N_22,In_1525,In_1028);
nor U23 (N_23,In_205,In_1350);
or U24 (N_24,In_1860,In_1586);
nand U25 (N_25,In_1365,In_1706);
or U26 (N_26,In_401,In_432);
and U27 (N_27,In_1109,In_1167);
xor U28 (N_28,In_1409,In_1117);
or U29 (N_29,In_485,In_570);
and U30 (N_30,In_1490,In_1536);
or U31 (N_31,In_1532,In_1169);
nor U32 (N_32,In_1074,In_1429);
xnor U33 (N_33,In_816,In_1567);
xnor U34 (N_34,In_1862,In_1018);
nand U35 (N_35,In_514,In_734);
nor U36 (N_36,In_1312,In_419);
and U37 (N_37,In_984,In_1946);
nor U38 (N_38,In_745,In_1118);
and U39 (N_39,In_1032,In_73);
nor U40 (N_40,In_1622,In_1043);
or U41 (N_41,In_384,In_886);
nor U42 (N_42,In_688,In_1817);
nor U43 (N_43,In_1015,In_814);
or U44 (N_44,In_772,In_1331);
xnor U45 (N_45,In_1217,In_6);
nor U46 (N_46,In_1507,In_1308);
and U47 (N_47,In_1003,In_716);
xnor U48 (N_48,In_575,In_1034);
or U49 (N_49,In_186,In_1443);
nand U50 (N_50,In_1066,In_607);
nand U51 (N_51,In_689,In_1592);
or U52 (N_52,In_1940,In_128);
and U53 (N_53,In_1403,In_858);
xnor U54 (N_54,In_791,In_195);
or U55 (N_55,In_1989,In_92);
or U56 (N_56,In_1480,In_673);
nand U57 (N_57,In_1575,In_1235);
and U58 (N_58,In_1643,In_974);
xnor U59 (N_59,In_1799,In_1207);
nand U60 (N_60,In_1992,In_988);
xnor U61 (N_61,In_489,In_764);
or U62 (N_62,In_147,In_1256);
nand U63 (N_63,In_633,In_962);
nand U64 (N_64,In_758,In_1195);
nand U65 (N_65,In_926,In_473);
or U66 (N_66,In_582,In_242);
and U67 (N_67,In_903,In_1280);
nand U68 (N_68,In_249,In_1296);
or U69 (N_69,In_1017,In_621);
nor U70 (N_70,In_1483,In_185);
and U71 (N_71,In_49,In_1760);
nand U72 (N_72,In_1197,In_878);
nand U73 (N_73,In_1267,In_496);
and U74 (N_74,In_663,In_1372);
nor U75 (N_75,In_228,In_1944);
nand U76 (N_76,In_1617,In_1655);
or U77 (N_77,In_961,In_1964);
or U78 (N_78,In_1438,In_261);
nand U79 (N_79,In_1485,In_1423);
nor U80 (N_80,In_580,In_91);
nor U81 (N_81,In_150,In_889);
xnor U82 (N_82,In_339,In_1722);
or U83 (N_83,In_341,In_1460);
and U84 (N_84,In_1090,In_1237);
nor U85 (N_85,In_742,In_708);
or U86 (N_86,In_653,In_1792);
xor U87 (N_87,In_1300,In_76);
nand U88 (N_88,In_0,In_146);
and U89 (N_89,In_366,In_600);
nand U90 (N_90,In_1373,In_113);
nand U91 (N_91,In_241,In_1902);
and U92 (N_92,In_971,In_1950);
nor U93 (N_93,In_1291,In_1226);
or U94 (N_94,In_246,In_324);
nor U95 (N_95,In_565,In_284);
nor U96 (N_96,In_1664,In_180);
and U97 (N_97,In_7,In_546);
nand U98 (N_98,In_1837,In_1975);
or U99 (N_99,In_426,In_1275);
and U100 (N_100,In_944,In_477);
nand U101 (N_101,In_1475,In_1619);
or U102 (N_102,In_528,In_1108);
or U103 (N_103,In_1642,In_38);
nor U104 (N_104,In_1138,In_17);
xnor U105 (N_105,In_447,In_1590);
nand U106 (N_106,In_695,In_63);
xor U107 (N_107,In_1796,In_1220);
xor U108 (N_108,In_817,In_19);
xor U109 (N_109,In_1910,In_1002);
nor U110 (N_110,In_1347,In_394);
nand U111 (N_111,In_1891,In_18);
or U112 (N_112,In_910,In_414);
and U113 (N_113,In_389,In_1768);
nor U114 (N_114,In_1131,In_1029);
and U115 (N_115,In_1582,In_1440);
nor U116 (N_116,In_1835,In_1345);
and U117 (N_117,In_435,In_1355);
xnor U118 (N_118,In_549,In_885);
nand U119 (N_119,In_482,In_374);
nor U120 (N_120,In_1542,In_1095);
or U121 (N_121,In_1496,In_1925);
and U122 (N_122,In_1875,In_529);
nand U123 (N_123,In_112,In_1265);
nor U124 (N_124,In_844,In_397);
xor U125 (N_125,In_297,In_1659);
xor U126 (N_126,In_1165,In_1382);
nand U127 (N_127,In_1246,In_1588);
nor U128 (N_128,In_665,In_662);
nand U129 (N_129,In_392,In_196);
and U130 (N_130,In_90,In_1182);
nor U131 (N_131,In_1897,In_1122);
xnor U132 (N_132,In_101,In_198);
xor U133 (N_133,In_1299,In_1119);
nand U134 (N_134,In_991,In_1321);
and U135 (N_135,In_586,In_1302);
nor U136 (N_136,In_1949,In_651);
nor U137 (N_137,In_1405,In_942);
xor U138 (N_138,In_1729,In_761);
xor U139 (N_139,In_171,In_760);
nand U140 (N_140,In_627,In_382);
nand U141 (N_141,In_1545,In_61);
nand U142 (N_142,In_177,In_157);
and U143 (N_143,In_1569,In_1080);
nand U144 (N_144,In_613,In_958);
and U145 (N_145,In_1395,In_1811);
nor U146 (N_146,In_1273,In_47);
or U147 (N_147,In_1600,In_1036);
nand U148 (N_148,In_288,In_1363);
nand U149 (N_149,In_1132,In_1529);
xor U150 (N_150,In_1863,In_768);
and U151 (N_151,In_1635,In_1644);
nor U152 (N_152,In_960,In_1434);
xor U153 (N_153,In_1271,In_254);
xor U154 (N_154,In_1114,In_915);
nor U155 (N_155,In_1936,In_1063);
xnor U156 (N_156,In_1621,In_1868);
and U157 (N_157,In_1625,In_1371);
xnor U158 (N_158,In_1081,In_1505);
xnor U159 (N_159,In_1924,In_1758);
nor U160 (N_160,In_1879,In_1392);
or U161 (N_161,In_1848,In_151);
and U162 (N_162,In_932,In_1938);
or U163 (N_163,In_1603,In_1213);
nor U164 (N_164,In_1412,In_1918);
and U165 (N_165,In_963,In_1394);
xnor U166 (N_166,In_812,In_1324);
or U167 (N_167,In_58,In_1473);
nand U168 (N_168,In_108,In_271);
xnor U169 (N_169,In_1761,In_609);
xnor U170 (N_170,In_1315,In_747);
and U171 (N_171,In_1309,In_1987);
xnor U172 (N_172,In_115,In_457);
nand U173 (N_173,In_415,In_1945);
xor U174 (N_174,In_1612,In_332);
or U175 (N_175,In_204,In_1608);
nand U176 (N_176,In_359,In_1222);
and U177 (N_177,In_1719,In_1769);
or U178 (N_178,In_798,In_980);
and U179 (N_179,In_1839,In_978);
xor U180 (N_180,In_1783,In_311);
and U181 (N_181,In_107,In_1931);
nor U182 (N_182,In_1135,In_1693);
xnor U183 (N_183,In_96,In_320);
or U184 (N_184,In_1516,In_1911);
nor U185 (N_185,In_133,In_1709);
nand U186 (N_186,In_57,In_1127);
xor U187 (N_187,In_162,In_1539);
or U188 (N_188,In_358,In_5);
xor U189 (N_189,In_285,In_1393);
nor U190 (N_190,In_492,In_1107);
or U191 (N_191,In_871,In_806);
nor U192 (N_192,In_129,In_1886);
or U193 (N_193,In_568,In_1115);
xnor U194 (N_194,In_276,In_1461);
or U195 (N_195,In_1223,In_620);
or U196 (N_196,In_774,In_503);
nand U197 (N_197,In_1319,In_1607);
nand U198 (N_198,In_20,In_1162);
and U199 (N_199,In_1375,In_1128);
xnor U200 (N_200,In_344,In_1976);
nor U201 (N_201,N_147,In_1654);
or U202 (N_202,In_243,In_175);
xnor U203 (N_203,In_879,In_1069);
nand U204 (N_204,In_220,N_56);
and U205 (N_205,N_155,In_1183);
or U206 (N_206,In_495,In_1203);
nand U207 (N_207,In_1947,N_153);
and U208 (N_208,In_1113,In_111);
and U209 (N_209,In_398,In_1663);
or U210 (N_210,In_1164,In_362);
nand U211 (N_211,N_137,N_73);
and U212 (N_212,In_323,In_280);
nor U213 (N_213,In_1045,In_617);
nand U214 (N_214,In_1673,N_55);
nand U215 (N_215,In_982,In_14);
nand U216 (N_216,In_1136,In_1882);
xnor U217 (N_217,In_50,In_676);
and U218 (N_218,In_1088,N_198);
xnor U219 (N_219,In_1874,In_661);
xnor U220 (N_220,In_628,In_685);
xor U221 (N_221,In_1996,In_1776);
or U222 (N_222,In_1951,In_1210);
or U223 (N_223,In_411,In_1431);
nor U224 (N_224,N_154,In_1422);
and U225 (N_225,In_1180,In_997);
nor U226 (N_226,In_1909,In_490);
and U227 (N_227,In_512,In_702);
xnor U228 (N_228,In_703,In_911);
and U229 (N_229,In_315,In_1142);
nand U230 (N_230,In_318,N_35);
or U231 (N_231,In_959,In_170);
and U232 (N_232,In_1419,In_863);
and U233 (N_233,In_937,In_1913);
nor U234 (N_234,In_85,In_51);
nor U235 (N_235,In_1895,In_1982);
nand U236 (N_236,In_1492,N_152);
xor U237 (N_237,In_52,In_1804);
nand U238 (N_238,In_691,In_552);
xnor U239 (N_239,In_522,In_780);
and U240 (N_240,In_418,In_1818);
nor U241 (N_241,In_827,In_598);
and U242 (N_242,N_196,In_1692);
or U243 (N_243,In_1921,In_588);
and U244 (N_244,In_902,In_521);
and U245 (N_245,N_53,In_28);
nor U246 (N_246,N_89,In_215);
nor U247 (N_247,In_310,In_648);
nor U248 (N_248,In_1675,In_1322);
nor U249 (N_249,In_1894,In_1008);
nor U250 (N_250,In_1899,N_103);
xor U251 (N_251,In_131,N_145);
nor U252 (N_252,In_1967,In_483);
xor U253 (N_253,In_706,N_7);
or U254 (N_254,In_348,In_957);
or U255 (N_255,In_722,In_1342);
or U256 (N_256,N_114,In_856);
nand U257 (N_257,In_829,In_919);
nand U258 (N_258,In_652,N_20);
or U259 (N_259,In_638,In_501);
xor U260 (N_260,In_104,In_31);
nand U261 (N_261,In_1741,In_563);
or U262 (N_262,In_591,In_712);
nor U263 (N_263,In_106,In_1543);
nor U264 (N_264,In_548,In_1881);
or U265 (N_265,In_1914,In_1933);
nor U266 (N_266,In_144,In_1649);
xnor U267 (N_267,In_785,In_1518);
and U268 (N_268,In_983,In_1867);
or U269 (N_269,In_1500,In_1971);
nor U270 (N_270,N_72,In_674);
xnor U271 (N_271,In_1010,In_1501);
nor U272 (N_272,In_1616,In_262);
and U273 (N_273,In_1187,In_237);
or U274 (N_274,In_1819,In_649);
or U275 (N_275,In_796,In_1055);
nor U276 (N_276,In_1990,In_566);
or U277 (N_277,In_535,N_36);
nand U278 (N_278,In_230,In_584);
or U279 (N_279,In_838,In_1742);
xnor U280 (N_280,N_101,In_361);
xor U281 (N_281,In_936,In_410);
xnor U282 (N_282,In_1629,N_118);
and U283 (N_283,In_235,In_302);
xnor U284 (N_284,In_165,In_1610);
xor U285 (N_285,In_644,In_66);
or U286 (N_286,In_1561,In_1687);
nor U287 (N_287,In_119,In_777);
or U288 (N_288,In_300,In_1301);
nand U289 (N_289,In_1842,In_1449);
or U290 (N_290,In_338,In_850);
or U291 (N_291,In_1620,In_1831);
and U292 (N_292,In_923,In_1006);
or U293 (N_293,In_1147,In_855);
nor U294 (N_294,In_173,In_1292);
and U295 (N_295,In_1563,N_49);
or U296 (N_296,In_508,In_1077);
nor U297 (N_297,In_905,In_947);
or U298 (N_298,N_128,In_352);
xor U299 (N_299,In_378,In_659);
xnor U300 (N_300,N_117,In_1685);
xor U301 (N_301,In_216,In_75);
nand U302 (N_302,In_1573,In_1853);
xnor U303 (N_303,N_14,In_191);
nand U304 (N_304,In_809,In_218);
nand U305 (N_305,In_1452,In_612);
or U306 (N_306,In_1704,In_705);
nor U307 (N_307,In_429,In_328);
nor U308 (N_308,In_1820,In_1474);
xor U309 (N_309,N_184,In_183);
nand U310 (N_310,In_142,In_370);
xnor U311 (N_311,In_553,In_1259);
or U312 (N_312,In_141,In_1058);
nor U313 (N_313,N_95,In_966);
nand U314 (N_314,In_547,In_287);
xnor U315 (N_315,In_1723,In_1454);
xnor U316 (N_316,N_186,In_172);
and U317 (N_317,In_1656,In_1979);
xor U318 (N_318,In_1790,In_1668);
or U319 (N_319,In_1215,In_1359);
nand U320 (N_320,In_1714,In_763);
xor U321 (N_321,In_805,In_1155);
or U322 (N_322,In_1143,In_1966);
nor U323 (N_323,In_124,In_1937);
nand U324 (N_324,In_46,N_140);
nor U325 (N_325,In_687,In_1040);
xor U326 (N_326,N_38,In_309);
nand U327 (N_327,In_594,In_655);
or U328 (N_328,In_901,In_1627);
and U329 (N_329,In_1427,In_1019);
and U330 (N_330,In_1439,In_53);
nand U331 (N_331,In_1823,In_1070);
or U332 (N_332,In_654,In_1623);
xnor U333 (N_333,In_1725,In_1572);
nor U334 (N_334,In_381,In_1367);
and U335 (N_335,In_724,In_1060);
and U336 (N_336,In_1067,In_964);
or U337 (N_337,In_632,In_577);
or U338 (N_338,In_301,In_630);
xnor U339 (N_339,In_386,In_290);
nor U340 (N_340,In_631,In_679);
or U341 (N_341,In_1794,In_336);
nand U342 (N_342,In_1777,In_445);
and U343 (N_343,In_610,In_86);
nor U344 (N_344,In_1387,In_412);
or U345 (N_345,In_446,In_405);
and U346 (N_346,In_459,In_240);
and U347 (N_347,In_666,In_792);
and U348 (N_348,In_1340,In_321);
nand U349 (N_349,In_727,N_163);
xnor U350 (N_350,In_1711,In_68);
xor U351 (N_351,In_795,In_505);
and U352 (N_352,In_833,In_1772);
or U353 (N_353,In_232,In_1836);
nand U354 (N_354,N_115,In_1857);
nor U355 (N_355,In_1056,In_42);
or U356 (N_356,In_1896,In_1468);
nand U357 (N_357,In_458,In_898);
or U358 (N_358,In_1998,N_173);
nand U359 (N_359,N_88,In_286);
xnor U360 (N_360,In_488,In_291);
nor U361 (N_361,In_298,In_826);
and U362 (N_362,In_484,In_71);
nand U363 (N_363,In_1024,In_894);
or U364 (N_364,In_752,In_343);
and U365 (N_365,In_1883,In_1606);
and U366 (N_366,In_1733,N_194);
nand U367 (N_367,In_1369,In_1374);
nor U368 (N_368,N_54,In_1806);
and U369 (N_369,In_1922,In_1228);
nor U370 (N_370,In_1385,In_765);
xor U371 (N_371,In_1171,In_1327);
nand U372 (N_372,In_1021,In_449);
nor U373 (N_373,In_436,In_767);
and U374 (N_374,In_1576,In_1802);
or U375 (N_375,In_634,In_313);
nand U376 (N_376,In_434,In_684);
and U377 (N_377,In_95,In_864);
xnor U378 (N_378,In_1391,In_1686);
nor U379 (N_379,In_744,In_1281);
xor U380 (N_380,N_27,In_1049);
and U381 (N_381,In_35,In_1759);
nor U382 (N_382,In_1329,In_943);
nor U383 (N_383,N_187,In_1465);
xor U384 (N_384,In_189,N_97);
nand U385 (N_385,In_754,In_1242);
or U386 (N_386,In_201,In_1803);
xnor U387 (N_387,N_109,In_714);
xor U388 (N_388,In_1912,In_1814);
or U389 (N_389,In_56,In_1232);
nor U390 (N_390,N_43,N_148);
and U391 (N_391,In_887,In_1807);
nor U392 (N_392,In_1145,In_1481);
xor U393 (N_393,In_1889,In_208);
and U394 (N_394,In_1159,In_1175);
xnor U395 (N_395,In_1991,In_606);
and U396 (N_396,In_1849,In_1014);
nor U397 (N_397,In_1270,In_1652);
xnor U398 (N_398,In_1445,In_1601);
xor U399 (N_399,In_578,In_1585);
nor U400 (N_400,N_286,In_1141);
and U401 (N_401,In_428,N_372);
nand U402 (N_402,N_328,In_1702);
xnor U403 (N_403,In_611,In_1718);
xor U404 (N_404,In_801,N_255);
or U405 (N_405,In_671,N_363);
and U406 (N_406,In_461,In_1358);
xor U407 (N_407,In_895,In_30);
or U408 (N_408,In_1176,In_1864);
nor U409 (N_409,N_245,N_8);
nor U410 (N_410,In_1731,In_1876);
nand U411 (N_411,In_1512,In_1958);
xor U412 (N_412,In_1757,In_1514);
nor U413 (N_413,In_1815,In_1954);
nand U414 (N_414,In_1389,In_466);
or U415 (N_415,In_1245,In_1337);
nor U416 (N_416,N_60,In_1243);
xnor U417 (N_417,In_604,In_1216);
nand U418 (N_418,In_707,In_1682);
nand U419 (N_419,In_1137,In_1188);
nand U420 (N_420,In_1283,In_1230);
and U421 (N_421,In_550,In_585);
and U422 (N_422,In_89,In_1917);
xor U423 (N_423,In_527,In_102);
and U424 (N_424,In_1851,N_300);
nor U425 (N_425,In_1707,In_592);
nor U426 (N_426,In_395,In_1866);
and U427 (N_427,In_718,In_27);
nor U428 (N_428,In_70,N_231);
xnor U429 (N_429,In_193,In_933);
and U430 (N_430,In_1435,In_1061);
or U431 (N_431,In_1763,N_271);
xnor U432 (N_432,In_454,In_1437);
or U433 (N_433,In_1844,In_599);
nand U434 (N_434,In_1482,In_741);
nor U435 (N_435,N_5,In_1139);
nor U436 (N_436,In_77,In_1578);
xor U437 (N_437,In_1751,In_1306);
nor U438 (N_438,In_1364,In_319);
nand U439 (N_439,In_815,In_272);
and U440 (N_440,In_1221,In_379);
nor U441 (N_441,In_929,N_358);
nor U442 (N_442,In_1878,N_383);
and U443 (N_443,In_408,In_1559);
nand U444 (N_444,In_509,In_1209);
nand U445 (N_445,In_203,In_664);
nor U446 (N_446,In_1808,N_268);
or U447 (N_447,N_377,N_37);
or U448 (N_448,In_1286,N_181);
nand U449 (N_449,In_176,In_993);
xor U450 (N_450,In_373,In_872);
or U451 (N_451,In_799,In_790);
xnor U452 (N_452,N_297,In_645);
and U453 (N_453,In_1052,N_1);
or U454 (N_454,N_4,In_1318);
or U455 (N_455,In_1873,N_249);
and U456 (N_456,In_1701,In_1614);
nand U457 (N_457,In_135,In_697);
nor U458 (N_458,In_899,In_1037);
or U459 (N_459,N_360,In_1589);
and U460 (N_460,In_955,In_569);
and U461 (N_461,In_1547,In_371);
nor U462 (N_462,N_176,In_1082);
and U463 (N_463,In_1968,In_375);
and U464 (N_464,In_140,In_656);
and U465 (N_465,In_681,In_1890);
or U466 (N_466,N_243,In_1755);
nand U467 (N_467,In_1700,In_1255);
and U468 (N_468,In_1277,In_1710);
and U469 (N_469,N_208,In_562);
or U470 (N_470,In_1420,In_896);
nand U471 (N_471,In_1970,In_1198);
xnor U472 (N_472,N_336,In_55);
nor U473 (N_473,N_345,In_802);
and U474 (N_474,In_1830,N_279);
and U475 (N_475,In_749,In_781);
xnor U476 (N_476,In_884,In_940);
or U477 (N_477,In_818,In_1756);
nor U478 (N_478,In_1923,N_121);
or U479 (N_479,In_1746,In_245);
or U480 (N_480,In_1352,In_1444);
and U481 (N_481,In_1747,In_267);
xor U482 (N_482,In_1597,In_1007);
or U483 (N_483,In_629,In_945);
nand U484 (N_484,In_1681,In_867);
nand U485 (N_485,In_480,In_756);
xnor U486 (N_486,N_64,In_169);
and U487 (N_487,In_238,In_1076);
and U488 (N_488,In_350,N_303);
or U489 (N_489,N_256,N_394);
or U490 (N_490,In_253,In_1083);
nor U491 (N_491,In_1871,N_151);
xor U492 (N_492,N_385,N_91);
or U493 (N_493,N_110,In_1489);
xnor U494 (N_494,In_922,In_1456);
and U495 (N_495,In_670,N_149);
and U496 (N_496,In_221,In_478);
nor U497 (N_497,In_158,In_194);
or U498 (N_498,In_1522,In_1520);
and U499 (N_499,In_746,In_1027);
xnor U500 (N_500,In_474,N_304);
and U501 (N_501,In_558,In_560);
nor U502 (N_502,In_640,N_99);
or U503 (N_503,N_223,In_701);
or U504 (N_504,In_986,In_1750);
and U505 (N_505,In_743,In_387);
xor U506 (N_506,In_1079,N_254);
nand U507 (N_507,In_54,N_326);
and U508 (N_508,In_259,In_1676);
or U509 (N_509,In_377,N_357);
or U510 (N_510,In_973,In_1289);
nand U511 (N_511,N_212,In_244);
or U512 (N_512,In_1624,In_507);
xor U513 (N_513,N_391,In_1721);
nand U514 (N_514,In_468,In_493);
nand U515 (N_515,In_179,In_37);
nand U516 (N_516,In_1715,In_476);
nand U517 (N_517,In_1541,In_1898);
and U518 (N_518,In_1553,In_1749);
or U519 (N_519,In_1744,In_834);
nor U520 (N_520,In_1430,In_1411);
xor U521 (N_521,N_314,In_322);
xnor U522 (N_522,In_865,N_388);
nor U523 (N_523,In_388,N_275);
nand U524 (N_524,In_1287,N_39);
nand U525 (N_525,In_64,In_912);
nor U526 (N_526,N_356,N_227);
xor U527 (N_527,N_119,In_433);
and U528 (N_528,In_1905,N_193);
xor U529 (N_529,In_308,In_1782);
or U530 (N_530,In_1407,In_427);
or U531 (N_531,In_462,In_1035);
nand U532 (N_532,In_1956,In_1272);
nand U533 (N_533,In_808,In_425);
nand U534 (N_534,In_417,In_479);
or U535 (N_535,In_1200,N_12);
and U536 (N_536,N_312,In_537);
nand U537 (N_537,In_353,N_277);
nand U538 (N_538,In_60,N_146);
nor U539 (N_539,In_1151,In_317);
nor U540 (N_540,N_384,In_1695);
nand U541 (N_541,N_387,In_1821);
nor U542 (N_542,In_1577,In_1678);
xor U543 (N_543,In_1859,In_1294);
and U544 (N_544,N_290,In_1907);
or U545 (N_545,N_71,In_740);
xnor U546 (N_546,In_1647,In_1730);
nor U547 (N_547,In_360,In_1789);
nand U548 (N_548,In_539,In_72);
and U549 (N_549,In_890,In_1551);
and U550 (N_550,In_506,N_348);
nor U551 (N_551,In_1307,In_823);
nand U552 (N_552,In_1338,In_1314);
and U553 (N_553,N_29,In_316);
nor U554 (N_554,In_1432,N_334);
or U555 (N_555,In_1540,In_351);
nor U556 (N_556,In_1838,In_900);
nand U557 (N_557,In_985,N_66);
xor U558 (N_558,In_587,In_16);
xnor U559 (N_559,In_536,In_266);
nor U560 (N_560,In_713,In_1455);
xnor U561 (N_561,In_187,In_729);
or U562 (N_562,N_63,N_127);
xor U563 (N_563,In_182,In_399);
nand U564 (N_564,In_327,In_1775);
and U565 (N_565,N_232,N_397);
and U566 (N_566,In_1166,N_267);
or U567 (N_567,N_138,In_12);
or U568 (N_568,In_987,In_1205);
and U569 (N_569,N_332,N_33);
nand U570 (N_570,N_156,In_364);
nand U571 (N_571,In_1671,In_1381);
and U572 (N_572,In_642,In_110);
xnor U573 (N_573,In_441,In_1795);
nand U574 (N_574,N_24,In_888);
xor U575 (N_575,In_1304,In_1988);
and U576 (N_576,In_1089,N_278);
xnor U577 (N_577,In_1986,In_1800);
xnor U578 (N_578,In_168,In_602);
xnor U579 (N_579,N_369,N_122);
nand U580 (N_580,In_100,In_1810);
nand U581 (N_581,N_58,In_524);
or U582 (N_582,In_1099,In_1713);
nand U583 (N_583,N_78,In_1587);
nand U584 (N_584,In_167,In_927);
nor U585 (N_585,In_1133,In_538);
nand U586 (N_586,In_1549,In_438);
and U587 (N_587,In_635,In_442);
nand U588 (N_588,N_320,In_1502);
or U589 (N_589,In_130,In_571);
and U590 (N_590,In_851,In_1100);
xnor U591 (N_591,In_1667,N_28);
and U592 (N_592,In_561,In_800);
nor U593 (N_593,In_148,In_857);
xor U594 (N_594,In_1841,In_197);
xnor U595 (N_595,In_616,N_355);
and U596 (N_596,In_1865,In_581);
xnor U597 (N_597,In_213,In_1376);
or U598 (N_598,N_298,In_1765);
xor U599 (N_599,In_989,N_65);
nand U600 (N_600,In_1517,In_624);
or U601 (N_601,N_477,In_114);
or U602 (N_602,In_334,N_506);
xor U603 (N_603,In_601,In_891);
nor U604 (N_604,In_1016,In_346);
or U605 (N_605,N_185,In_1650);
or U606 (N_606,In_876,N_414);
nor U607 (N_607,In_750,In_1106);
and U608 (N_608,N_234,In_950);
and U609 (N_609,N_491,N_505);
xor U610 (N_610,In_534,In_83);
and U611 (N_611,N_90,In_573);
nand U612 (N_612,N_226,In_1054);
xnor U613 (N_613,In_1646,N_375);
nor U614 (N_614,N_46,N_503);
and U615 (N_615,In_751,In_660);
xor U616 (N_616,In_759,In_1383);
nand U617 (N_617,N_253,In_1186);
or U618 (N_618,In_831,In_916);
xor U619 (N_619,In_968,N_159);
or U620 (N_620,N_474,In_283);
and U621 (N_621,N_190,In_143);
and U622 (N_622,N_516,N_217);
and U623 (N_623,In_636,In_1679);
nand U624 (N_624,In_1633,N_459);
xnor U625 (N_625,In_1584,In_1253);
nand U626 (N_626,N_273,In_1112);
and U627 (N_627,In_576,In_717);
nand U628 (N_628,In_544,In_728);
nor U629 (N_629,In_1330,In_212);
nor U630 (N_630,N_573,In_1708);
xnor U631 (N_631,In_1703,N_510);
nor U632 (N_632,In_1249,In_1125);
nor U633 (N_633,In_1858,In_1877);
nand U634 (N_634,N_433,In_248);
nand U635 (N_635,N_429,In_1552);
nand U636 (N_636,N_507,In_210);
and U637 (N_637,In_1916,In_934);
nand U638 (N_638,In_270,In_1639);
xor U639 (N_639,In_1884,In_1596);
or U640 (N_640,In_1154,In_597);
nand U641 (N_641,N_228,In_1985);
nor U642 (N_642,In_564,N_106);
and U643 (N_643,In_1771,N_235);
xnor U644 (N_644,N_577,In_1179);
or U645 (N_645,In_1450,In_498);
xor U646 (N_646,In_1144,In_1981);
xnor U647 (N_647,In_625,In_1472);
and U648 (N_648,N_554,N_411);
xor U649 (N_649,In_1193,N_430);
and U650 (N_650,N_265,In_209);
xor U651 (N_651,In_1738,In_1870);
nand U652 (N_652,In_626,In_1995);
or U653 (N_653,N_295,In_1670);
nand U654 (N_654,N_352,In_605);
nor U655 (N_655,In_1328,In_992);
nand U656 (N_656,N_269,In_643);
nand U657 (N_657,In_861,In_614);
or U658 (N_658,In_682,In_672);
nand U659 (N_659,In_619,N_296);
nand U660 (N_660,In_1994,N_415);
nor U661 (N_661,In_1446,In_1284);
and U662 (N_662,In_1261,N_359);
xor U663 (N_663,In_1469,In_710);
and U664 (N_664,In_1504,In_949);
or U665 (N_665,In_1199,In_491);
or U666 (N_666,In_1105,N_435);
and U667 (N_667,N_465,In_1538);
nor U668 (N_668,N_439,N_45);
and U669 (N_669,In_1962,In_200);
and U670 (N_670,In_152,In_1666);
nand U671 (N_671,N_381,In_853);
xor U672 (N_672,N_487,In_646);
or U673 (N_673,N_242,In_1948);
or U674 (N_674,N_583,In_385);
nand U675 (N_675,N_287,N_51);
nor U676 (N_676,In_84,N_313);
nand U677 (N_677,In_1963,In_10);
nor U678 (N_678,In_424,In_1762);
and U679 (N_679,In_1892,In_23);
and U680 (N_680,In_939,In_87);
nor U681 (N_681,N_3,In_69);
nand U682 (N_682,In_866,In_207);
nor U683 (N_683,In_1684,In_822);
or U684 (N_684,In_1390,In_1303);
and U685 (N_685,N_250,In_946);
and U686 (N_686,N_26,In_517);
nor U687 (N_687,In_1983,N_371);
or U688 (N_688,In_413,In_154);
nor U689 (N_689,In_1084,In_1826);
nand U690 (N_690,In_1279,N_424);
nand U691 (N_691,In_709,In_1126);
or U692 (N_692,N_306,In_1124);
nor U693 (N_693,In_1615,N_570);
nand U694 (N_694,In_1556,In_1523);
nand U695 (N_695,N_454,In_1274);
nand U696 (N_696,In_1349,N_83);
nand U697 (N_697,N_165,N_307);
xnor U698 (N_698,N_319,N_571);
and U699 (N_699,In_1146,In_1042);
nand U700 (N_700,In_1011,N_123);
nor U701 (N_701,In_786,In_1097);
xnor U702 (N_702,In_1293,In_641);
xor U703 (N_703,N_220,N_511);
xnor U704 (N_704,N_467,N_131);
xnor U705 (N_705,N_308,N_175);
or U706 (N_706,In_907,In_1173);
nor U707 (N_707,In_1023,In_789);
nor U708 (N_708,N_251,N_349);
xnor U709 (N_709,N_260,In_526);
xnor U710 (N_710,In_1250,N_338);
and U711 (N_711,N_421,In_1344);
nand U712 (N_712,In_423,N_504);
and U713 (N_713,N_162,In_440);
and U714 (N_714,N_518,N_233);
nor U715 (N_715,In_545,N_224);
or U716 (N_716,In_421,N_406);
or U717 (N_717,N_453,In_1634);
nor U718 (N_718,In_1263,In_821);
nor U719 (N_719,In_726,In_797);
xnor U720 (N_720,N_537,In_263);
nor U721 (N_721,N_142,In_1202);
nor U722 (N_722,In_1120,In_515);
or U723 (N_723,In_277,N_263);
and U724 (N_724,N_426,In_1348);
and U725 (N_725,N_393,N_502);
nand U726 (N_726,In_188,In_1739);
xor U727 (N_727,N_32,N_498);
xor U728 (N_728,N_546,In_731);
nor U729 (N_729,N_480,N_100);
or U730 (N_730,In_567,N_317);
or U731 (N_731,In_773,N_309);
nor U732 (N_732,In_693,In_782);
or U733 (N_733,In_1479,In_1594);
or U734 (N_734,In_1424,In_269);
nand U735 (N_735,In_437,In_1103);
nor U736 (N_736,In_1508,N_206);
nand U737 (N_737,In_439,N_538);
or U738 (N_738,N_460,In_502);
nor U739 (N_739,N_353,In_893);
nor U740 (N_740,In_848,In_307);
and U741 (N_741,In_525,In_139);
nor U742 (N_742,In_1051,In_803);
or U743 (N_743,N_361,In_1506);
or U744 (N_744,N_321,In_825);
xor U745 (N_745,In_1961,In_1726);
xor U746 (N_746,N_404,In_1929);
xor U747 (N_747,N_22,N_434);
nand U748 (N_748,In_1311,N_366);
nor U749 (N_749,N_130,N_134);
xor U750 (N_750,In_1528,In_970);
xor U751 (N_751,In_225,N_9);
nor U752 (N_752,N_327,N_266);
and U753 (N_753,In_1388,In_1960);
xnor U754 (N_754,N_447,In_965);
and U755 (N_755,In_329,N_335);
xor U756 (N_756,In_1869,In_256);
xor U757 (N_757,In_804,In_909);
xor U758 (N_758,In_347,In_1410);
or U759 (N_759,In_583,N_178);
xnor U760 (N_760,In_274,N_284);
nor U761 (N_761,In_1503,N_105);
nand U762 (N_762,In_1827,In_1357);
nor U763 (N_763,In_1662,In_303);
nor U764 (N_764,N_386,In_1185);
nand U765 (N_765,In_1129,In_1156);
or U766 (N_766,In_153,N_364);
nand U767 (N_767,In_80,In_299);
or U768 (N_768,In_98,In_1781);
and U769 (N_769,In_1724,In_1415);
nand U770 (N_770,In_1158,In_1290);
nand U771 (N_771,In_279,In_1697);
and U772 (N_772,In_1801,In_416);
xnor U773 (N_773,In_79,In_794);
nor U774 (N_774,In_1712,N_579);
xor U775 (N_775,N_76,In_680);
nand U776 (N_776,In_383,In_1591);
nand U777 (N_777,In_513,In_1062);
and U778 (N_778,In_1368,N_331);
nor U779 (N_779,N_259,N_210);
and U780 (N_780,In_331,In_1688);
nand U781 (N_781,In_1417,N_497);
nor U782 (N_782,In_810,N_378);
or U783 (N_783,In_1334,In_67);
or U784 (N_784,In_704,N_293);
or U785 (N_785,N_77,In_1057);
or U786 (N_786,In_1451,N_456);
and U787 (N_787,In_1254,N_392);
nand U788 (N_788,N_270,In_306);
nand U789 (N_789,In_1571,In_1778);
xor U790 (N_790,In_555,In_686);
nand U791 (N_791,In_1231,In_404);
and U792 (N_792,In_1696,In_48);
xnor U793 (N_793,N_466,N_365);
xor U794 (N_794,In_914,In_499);
xor U795 (N_795,In_390,In_1386);
and U796 (N_796,N_339,N_552);
and U797 (N_797,In_1453,In_1641);
nor U798 (N_798,In_1192,In_1053);
nor U799 (N_799,In_1754,In_1764);
and U800 (N_800,In_1478,N_241);
or U801 (N_801,N_713,In_456);
nor U802 (N_802,N_662,In_463);
or U803 (N_803,N_722,N_778);
nor U804 (N_804,N_428,N_591);
and U805 (N_805,In_1904,N_168);
xnor U806 (N_806,N_794,In_1674);
xor U807 (N_807,N_527,N_323);
nand U808 (N_808,In_1787,N_195);
and U809 (N_809,N_61,In_1096);
nand U810 (N_810,N_171,In_1012);
nand U811 (N_811,In_1524,N_139);
xor U812 (N_812,In_860,N_600);
nand U813 (N_813,In_1579,In_675);
nand U814 (N_814,In_843,N_292);
nand U815 (N_815,N_731,N_79);
and U816 (N_816,N_455,N_702);
nand U817 (N_817,N_410,In_1598);
and U818 (N_818,In_1104,N_747);
nor U819 (N_819,In_1570,N_344);
xnor U820 (N_820,In_1872,In_637);
and U821 (N_821,N_606,N_274);
xor U822 (N_822,N_17,N_347);
or U823 (N_823,In_1980,In_771);
nand U824 (N_824,In_1025,In_1736);
and U825 (N_825,In_981,In_1786);
nand U826 (N_826,In_542,N_325);
xnor U827 (N_827,In_967,In_206);
xnor U828 (N_828,In_1880,In_1224);
xnor U829 (N_829,In_1022,N_795);
nand U830 (N_830,In_181,In_82);
nand U831 (N_831,In_1728,N_125);
nand U832 (N_832,N_136,In_775);
xor U833 (N_833,N_788,N_225);
nand U834 (N_834,N_765,In_1611);
nor U835 (N_835,N_655,N_663);
and U836 (N_836,N_564,N_451);
xor U837 (N_837,In_1797,N_170);
nor U838 (N_838,In_948,In_1631);
xor U839 (N_839,N_593,In_314);
or U840 (N_840,In_1190,N_532);
nand U841 (N_841,N_108,In_913);
nor U842 (N_842,N_568,N_486);
or U843 (N_843,N_699,N_337);
xnor U844 (N_844,N_555,In_1400);
nand U845 (N_845,N_512,N_86);
nor U846 (N_846,In_531,In_748);
nor U847 (N_847,In_951,N_412);
nand U848 (N_848,N_230,In_120);
nor U849 (N_849,In_26,N_749);
nor U850 (N_850,N_449,In_842);
nand U851 (N_851,In_1773,N_437);
xnor U852 (N_852,In_1238,In_779);
or U853 (N_853,N_793,In_1978);
or U854 (N_854,In_1380,N_221);
nand U855 (N_855,In_1645,In_551);
xor U856 (N_856,In_1402,N_534);
nand U857 (N_857,In_1753,In_832);
nand U858 (N_858,In_1397,In_121);
or U859 (N_859,In_931,In_1068);
nor U860 (N_860,In_293,In_369);
xor U861 (N_861,N_672,In_994);
xnor U862 (N_862,In_1534,In_356);
nand U863 (N_863,N_706,N_634);
or U864 (N_864,N_322,In_975);
nor U865 (N_865,In_696,In_236);
and U866 (N_866,N_315,N_436);
or U867 (N_867,N_744,In_1934);
and U868 (N_868,In_260,In_1554);
nand U869 (N_869,In_1047,In_199);
xnor U870 (N_870,N_614,N_422);
and U871 (N_871,N_350,N_183);
or U872 (N_872,In_164,N_282);
nor U873 (N_873,In_1805,In_1384);
nand U874 (N_874,In_78,N_612);
and U875 (N_875,In_1580,N_262);
nor U876 (N_876,N_276,In_1343);
or U877 (N_877,N_535,N_701);
xor U878 (N_878,N_657,N_346);
nor U879 (N_879,N_721,In_400);
or U880 (N_880,N_729,In_122);
nand U881 (N_881,In_1698,N_705);
or U882 (N_882,N_646,In_753);
and U883 (N_883,In_239,N_515);
xnor U884 (N_884,N_373,N_677);
nand U885 (N_885,In_393,In_1229);
and U886 (N_886,In_123,N_541);
or U887 (N_887,N_494,In_720);
nand U888 (N_888,N_252,In_1533);
xnor U889 (N_889,N_616,In_282);
and U890 (N_890,In_1565,In_990);
nor U891 (N_891,In_93,In_1845);
or U892 (N_892,N_755,In_711);
nand U893 (N_893,In_226,In_1163);
or U894 (N_894,In_739,In_925);
or U895 (N_895,N_343,In_1408);
xnor U896 (N_896,In_1251,In_1377);
and U897 (N_897,N_520,In_1252);
or U898 (N_898,In_1665,In_1943);
xor U899 (N_899,N_272,In_783);
nor U900 (N_900,In_572,In_1476);
and U901 (N_901,In_1885,In_1211);
or U902 (N_902,N_628,N_797);
nand U903 (N_903,In_793,N_608);
and U904 (N_904,In_1241,In_721);
or U905 (N_905,In_723,In_1048);
or U906 (N_906,N_601,N_696);
or U907 (N_907,In_1442,In_1766);
nor U908 (N_908,In_304,N_81);
nor U909 (N_909,In_1288,In_1448);
xor U910 (N_910,In_669,N_660);
nand U911 (N_911,N_751,In_1908);
or U912 (N_912,In_1326,In_88);
nand U913 (N_913,In_1926,N_528);
and U914 (N_914,In_1001,N_746);
or U915 (N_915,In_1993,N_605);
nand U916 (N_916,N_627,In_543);
xnor U917 (N_917,N_737,In_1418);
and U918 (N_918,N_724,N_620);
nor U919 (N_919,N_768,In_1737);
or U920 (N_920,In_935,In_956);
and U921 (N_921,N_222,N_120);
or U922 (N_922,In_219,N_246);
or U923 (N_923,N_580,N_425);
and U924 (N_924,In_1930,In_109);
or U925 (N_925,In_1149,N_398);
nand U926 (N_926,In_1091,N_642);
xor U927 (N_927,N_670,N_586);
or U928 (N_928,N_470,In_875);
nor U929 (N_929,In_1101,N_111);
or U930 (N_930,In_1194,In_1903);
nand U931 (N_931,In_1148,N_407);
xnor U932 (N_932,In_579,In_852);
nor U933 (N_933,In_1599,N_219);
nand U934 (N_934,In_846,N_141);
nor U935 (N_935,In_1341,In_380);
nand U936 (N_936,In_1581,In_1511);
nor U937 (N_937,In_1566,In_1401);
nand U938 (N_938,N_75,N_21);
and U939 (N_939,In_658,In_155);
xor U940 (N_940,In_920,In_367);
nand U941 (N_941,In_325,N_257);
xor U942 (N_942,In_1855,In_1493);
and U943 (N_943,N_403,In_873);
nand U944 (N_944,In_1191,In_1583);
nor U945 (N_945,N_569,N_318);
nor U946 (N_946,In_1098,In_460);
nor U947 (N_947,In_229,In_1208);
and U948 (N_948,In_1735,In_1847);
or U949 (N_949,N_654,N_710);
and U950 (N_950,In_735,In_921);
nor U951 (N_951,In_1219,N_621);
nand U952 (N_952,In_340,N_578);
nand U953 (N_953,N_787,In_1513);
nand U954 (N_954,N_550,In_770);
xor U955 (N_955,N_485,In_1041);
nor U956 (N_956,In_1406,N_182);
nor U957 (N_957,N_561,In_1004);
xnor U958 (N_958,In_897,In_1470);
or U959 (N_959,In_1677,N_19);
xor U960 (N_960,N_67,N_659);
xor U961 (N_961,In_830,N_248);
xnor U962 (N_962,N_215,In_4);
nor U963 (N_963,N_595,N_305);
nor U964 (N_964,In_683,In_839);
nand U965 (N_965,In_1033,In_622);
or U966 (N_966,N_758,In_762);
xnor U967 (N_967,In_81,N_13);
and U968 (N_968,In_1065,In_1240);
nor U969 (N_969,N_418,N_777);
xnor U970 (N_970,In_273,In_1888);
and U971 (N_971,N_689,N_102);
and U972 (N_972,In_1336,In_117);
nand U973 (N_973,In_1323,In_1637);
or U974 (N_974,In_1791,N_11);
xnor U975 (N_975,In_1788,In_1071);
xor U976 (N_976,In_217,N_158);
and U977 (N_977,N_540,In_1398);
and U978 (N_978,In_45,In_1378);
and U979 (N_979,N_548,N_549);
or U980 (N_980,N_693,In_1168);
nand U981 (N_981,In_354,N_563);
xnor U982 (N_982,N_590,N_280);
or U983 (N_983,In_1030,N_201);
xor U984 (N_984,N_779,N_690);
and U985 (N_985,In_264,In_1499);
and U986 (N_986,In_766,N_790);
nor U987 (N_987,N_237,In_1833);
nor U988 (N_988,In_559,In_540);
and U989 (N_989,N_484,In_976);
nand U990 (N_990,In_1560,N_633);
and U991 (N_991,In_132,In_174);
xor U992 (N_992,In_1521,In_1699);
nand U993 (N_993,In_737,N_771);
nor U994 (N_994,In_1013,In_1784);
or U995 (N_995,In_99,N_592);
and U996 (N_996,In_1,In_1928);
or U997 (N_997,In_126,In_1564);
and U998 (N_998,In_234,In_251);
xor U999 (N_999,In_678,In_1262);
or U1000 (N_1000,N_735,N_639);
and U1001 (N_1001,In_1498,N_855);
nand U1002 (N_1002,In_1557,N_819);
xnor U1003 (N_1003,In_137,In_1752);
nor U1004 (N_1004,In_1310,N_643);
and U1005 (N_1005,In_422,In_977);
nand U1006 (N_1006,In_275,N_889);
nor U1007 (N_1007,N_602,N_458);
nand U1008 (N_1008,In_1793,N_958);
xor U1009 (N_1009,N_964,N_409);
nor U1010 (N_1010,N_133,In_1038);
xor U1011 (N_1011,In_516,In_32);
or U1012 (N_1012,In_1550,In_725);
nor U1013 (N_1013,N_971,In_1957);
or U1014 (N_1014,N_483,N_342);
nor U1015 (N_1015,In_738,In_1005);
and U1016 (N_1016,N_47,In_1000);
xor U1017 (N_1017,In_1236,N_866);
nor U1018 (N_1018,N_870,In_1562);
xor U1019 (N_1019,In_337,N_144);
xor U1020 (N_1020,In_1248,N_299);
nand U1021 (N_1021,N_878,In_1093);
or U1022 (N_1022,N_963,In_335);
nand U1023 (N_1023,N_104,N_961);
nand U1024 (N_1024,N_551,N_70);
or U1025 (N_1025,N_995,N_200);
nand U1026 (N_1026,N_860,In_1239);
xor U1027 (N_1027,N_468,N_741);
nor U1028 (N_1028,In_1177,N_463);
nand U1029 (N_1029,N_653,N_446);
nand U1030 (N_1030,N_985,N_330);
nor U1031 (N_1031,In_1974,N_539);
and U1032 (N_1032,N_34,N_74);
xnor U1033 (N_1033,In_954,N_417);
nor U1034 (N_1034,N_974,N_980);
nor U1035 (N_1035,In_1157,N_444);
xnor U1036 (N_1036,In_1509,In_820);
nand U1037 (N_1037,N_786,In_184);
nor U1038 (N_1038,N_523,N_843);
or U1039 (N_1039,In_1537,In_1530);
nor U1040 (N_1040,N_685,In_333);
and U1041 (N_1041,N_390,N_871);
and U1042 (N_1042,N_783,N_695);
or U1043 (N_1043,N_824,In_1494);
xor U1044 (N_1044,In_1413,N_805);
and U1045 (N_1045,In_1269,N_977);
nand U1046 (N_1046,N_941,N_869);
nand U1047 (N_1047,In_41,N_770);
nand U1048 (N_1048,In_1266,N_769);
nor U1049 (N_1049,N_82,N_522);
and U1050 (N_1050,In_1285,In_999);
nor U1051 (N_1051,In_1214,N_396);
xor U1052 (N_1052,In_1969,In_883);
and U1053 (N_1053,N_830,N_681);
xor U1054 (N_1054,N_2,N_845);
xor U1055 (N_1055,N_427,In_574);
xnor U1056 (N_1056,N_675,N_825);
and U1057 (N_1057,In_1297,In_481);
and U1058 (N_1058,N_461,N_838);
and U1059 (N_1059,N_906,In_1856);
nor U1060 (N_1060,N_567,N_953);
nor U1061 (N_1061,N_789,N_23);
xnor U1062 (N_1062,N_687,N_405);
xnor U1063 (N_1063,In_224,N_949);
xnor U1064 (N_1064,N_723,N_658);
and U1065 (N_1065,In_995,N_604);
or U1066 (N_1066,In_1094,N_93);
or U1067 (N_1067,N_898,In_281);
nor U1068 (N_1068,N_189,In_1399);
nor U1069 (N_1069,In_1351,N_529);
and U1070 (N_1070,In_227,N_400);
xnor U1071 (N_1071,In_1428,N_374);
nor U1072 (N_1072,N_59,N_822);
nand U1073 (N_1073,In_590,In_1110);
nor U1074 (N_1074,In_1370,In_1354);
and U1075 (N_1075,In_1843,N_736);
xnor U1076 (N_1076,In_268,N_536);
nor U1077 (N_1077,N_909,In_1196);
xnor U1078 (N_1078,N_626,In_1134);
xor U1079 (N_1079,In_854,N_25);
and U1080 (N_1080,In_1900,N_207);
nor U1081 (N_1081,N_890,N_966);
nor U1082 (N_1082,N_288,N_913);
xor U1083 (N_1083,N_939,In_202);
or U1084 (N_1084,N_928,In_11);
or U1085 (N_1085,N_833,In_1745);
or U1086 (N_1086,N_98,In_1335);
or U1087 (N_1087,In_252,In_402);
and U1088 (N_1088,In_1484,N_135);
nor U1089 (N_1089,In_650,N_730);
nand U1090 (N_1090,In_1111,In_1640);
nor U1091 (N_1091,N_164,N_918);
nor U1092 (N_1092,N_553,N_865);
and U1093 (N_1093,N_969,In_1595);
nand U1094 (N_1094,N_665,In_593);
nor U1095 (N_1095,N_341,In_1206);
and U1096 (N_1096,In_1626,N_885);
or U1097 (N_1097,N_933,In_1657);
and U1098 (N_1098,In_116,N_711);
nand U1099 (N_1099,N_756,N_792);
xor U1100 (N_1100,N_811,In_467);
xor U1101 (N_1101,In_1332,In_647);
or U1102 (N_1102,In_1487,N_873);
nor U1103 (N_1103,In_487,In_1201);
nor U1104 (N_1104,In_882,In_1227);
xnor U1105 (N_1105,N_942,N_509);
nand U1106 (N_1106,N_946,N_442);
xor U1107 (N_1107,N_840,In_1816);
xor U1108 (N_1108,N_748,In_1244);
nand U1109 (N_1109,N_401,N_817);
nand U1110 (N_1110,In_1346,N_698);
or U1111 (N_1111,N_764,In_841);
and U1112 (N_1112,N_543,In_1906);
xnor U1113 (N_1113,N_806,N_340);
or U1114 (N_1114,In_452,N_851);
or U1115 (N_1115,N_598,In_1832);
xnor U1116 (N_1116,N_700,N_482);
nor U1117 (N_1117,N_647,N_513);
nand U1118 (N_1118,N_462,In_1716);
or U1119 (N_1119,N_798,In_1212);
nor U1120 (N_1120,N_707,In_1161);
nor U1121 (N_1121,In_530,N_624);
or U1122 (N_1122,In_1471,In_700);
or U1123 (N_1123,N_229,In_13);
nand U1124 (N_1124,In_25,In_1123);
or U1125 (N_1125,N_772,In_470);
nor U1126 (N_1126,In_1121,In_1046);
nand U1127 (N_1127,In_1218,In_556);
nor U1128 (N_1128,N_818,In_904);
nand U1129 (N_1129,N_925,In_589);
or U1130 (N_1130,N_982,N_413);
and U1131 (N_1131,N_472,N_519);
or U1132 (N_1132,N_908,N_804);
xor U1133 (N_1133,N_471,In_39);
xor U1134 (N_1134,N_129,N_760);
and U1135 (N_1135,N_191,In_1630);
nor U1136 (N_1136,In_1078,In_1463);
nor U1137 (N_1137,In_368,N_547);
and U1138 (N_1138,N_380,N_452);
nor U1139 (N_1139,In_1767,N_882);
and U1140 (N_1140,N_499,N_214);
xor U1141 (N_1141,N_395,N_87);
xor U1142 (N_1142,In_1278,N_572);
or U1143 (N_1143,N_929,In_1264);
nor U1144 (N_1144,In_326,N_937);
nor U1145 (N_1145,N_581,N_893);
or U1146 (N_1146,N_857,N_618);
or U1147 (N_1147,In_1379,In_1009);
nor U1148 (N_1148,N_517,N_999);
and U1149 (N_1149,In_1433,N_720);
nor U1150 (N_1150,N_703,N_683);
or U1151 (N_1151,In_836,In_1854);
xor U1152 (N_1152,In_278,N_574);
and U1153 (N_1153,N_919,N_907);
or U1154 (N_1154,N_754,In_214);
nor U1155 (N_1155,N_850,In_778);
xnor U1156 (N_1156,N_708,N_849);
or U1157 (N_1157,In_1669,In_952);
nand U1158 (N_1158,N_960,N_562);
and U1159 (N_1159,N_478,N_611);
nand U1160 (N_1160,N_836,In_391);
and U1161 (N_1161,In_1462,In_1268);
nor U1162 (N_1162,In_494,N_954);
nor U1163 (N_1163,In_1648,N_967);
and U1164 (N_1164,In_250,N_691);
and U1165 (N_1165,N_774,In_1458);
or U1166 (N_1166,In_1809,In_869);
xnor U1167 (N_1167,In_1932,In_1680);
and U1168 (N_1168,N_947,In_924);
nand U1169 (N_1169,N_679,N_203);
and U1170 (N_1170,In_1846,In_1258);
nor U1171 (N_1171,N_496,N_661);
nor U1172 (N_1172,N_861,N_715);
nor U1173 (N_1173,In_1690,N_416);
nand U1174 (N_1174,In_623,N_419);
and U1175 (N_1175,N_879,In_118);
nand U1176 (N_1176,N_493,N_10);
or U1177 (N_1177,N_514,In_15);
xnor U1178 (N_1178,N_962,N_874);
xnor U1179 (N_1179,N_169,N_476);
nand U1180 (N_1180,N_533,N_495);
or U1181 (N_1181,N_886,N_752);
or U1182 (N_1182,In_1467,In_211);
nor U1183 (N_1183,N_853,N_934);
or U1184 (N_1184,N_209,In_1574);
xnor U1185 (N_1185,N_188,In_1295);
and U1186 (N_1186,N_565,N_868);
nand U1187 (N_1187,In_603,In_615);
nand U1188 (N_1188,N_738,N_972);
nor U1189 (N_1189,In_1972,In_231);
and U1190 (N_1190,N_489,N_952);
nand U1191 (N_1191,N_166,In_1636);
nand U1192 (N_1192,N_438,N_852);
nor U1193 (N_1193,N_884,N_781);
xor U1194 (N_1194,N_559,N_989);
xnor U1195 (N_1195,In_677,In_1829);
nand U1196 (N_1196,N_160,N_566);
or U1197 (N_1197,In_1320,N_799);
and U1198 (N_1198,N_370,N_902);
nor U1199 (N_1199,N_809,N_932);
xnor U1200 (N_1200,In_1526,N_40);
nand U1201 (N_1201,In_930,In_1740);
and U1202 (N_1202,N_1036,N_475);
or U1203 (N_1203,N_1107,N_1026);
and U1204 (N_1204,In_1901,N_892);
nand U1205 (N_1205,N_441,N_997);
nor U1206 (N_1206,N_998,N_957);
xor U1207 (N_1207,N_1160,In_1939);
nor U1208 (N_1208,N_704,In_475);
nor U1209 (N_1209,In_1325,N_636);
and U1210 (N_1210,N_473,In_292);
and U1211 (N_1211,N_638,N_1148);
nand U1212 (N_1212,In_1366,In_1535);
or U1213 (N_1213,N_1114,N_940);
and U1214 (N_1214,N_648,In_1919);
or U1215 (N_1215,N_992,In_733);
nand U1216 (N_1216,N_1195,N_367);
and U1217 (N_1217,N_718,In_736);
nand U1218 (N_1218,In_1915,In_192);
nor U1219 (N_1219,N_450,In_127);
and U1220 (N_1220,N_920,N_1186);
xnor U1221 (N_1221,N_1055,N_94);
nor U1222 (N_1222,N_585,In_160);
or U1223 (N_1223,In_1447,N_1139);
nor U1224 (N_1224,N_1091,N_1196);
nor U1225 (N_1225,N_667,In_469);
xor U1226 (N_1226,In_265,N_1115);
or U1227 (N_1227,In_1181,N_557);
and U1228 (N_1228,N_1120,In_1189);
xnor U1229 (N_1229,In_1087,N_1079);
nand U1230 (N_1230,N_244,N_766);
nand U1231 (N_1231,N_211,N_1169);
nor U1232 (N_1232,N_1156,In_1425);
nand U1233 (N_1233,N_132,N_1146);
nor U1234 (N_1234,N_525,N_684);
or U1235 (N_1235,N_740,In_396);
or U1236 (N_1236,N_1138,N_651);
nand U1237 (N_1237,N_1178,N_1183);
and U1238 (N_1238,N_1048,N_1113);
and U1239 (N_1239,N_44,In_787);
or U1240 (N_1240,In_1732,N_859);
nor U1241 (N_1241,In_247,N_281);
xor U1242 (N_1242,N_829,N_686);
nor U1243 (N_1243,In_163,N_1135);
or U1244 (N_1244,N_915,N_1167);
nand U1245 (N_1245,N_1124,N_931);
xnor U1246 (N_1246,N_1053,In_62);
nand U1247 (N_1247,N_782,N_1064);
nor U1248 (N_1248,N_236,In_1257);
and U1249 (N_1249,N_978,In_1605);
nor U1250 (N_1250,N_1110,N_944);
xor U1251 (N_1251,N_938,N_694);
nor U1252 (N_1252,N_1180,N_1157);
or U1253 (N_1253,N_1105,N_481);
or U1254 (N_1254,N_842,N_238);
and U1255 (N_1255,In_1672,N_1073);
nor U1256 (N_1256,N_1188,In_464);
nor U1257 (N_1257,N_656,N_1025);
nand U1258 (N_1258,In_65,In_1774);
nand U1259 (N_1259,N_1068,N_50);
or U1260 (N_1260,N_1061,N_1019);
xnor U1261 (N_1261,In_312,N_1090);
or U1262 (N_1262,N_1016,N_1087);
or U1263 (N_1263,N_864,In_1770);
nand U1264 (N_1264,N_291,In_355);
and U1265 (N_1265,N_542,N_1027);
xnor U1266 (N_1266,In_1044,N_351);
nand U1267 (N_1267,N_814,N_285);
xor U1268 (N_1268,N_1150,In_59);
nor U1269 (N_1269,N_1123,In_444);
or U1270 (N_1270,N_167,N_1082);
or U1271 (N_1271,In_1632,In_1497);
xnor U1272 (N_1272,In_1510,N_955);
and U1273 (N_1273,In_1152,N_1075);
nand U1274 (N_1274,N_432,In_472);
xnor U1275 (N_1275,N_921,N_68);
nor U1276 (N_1276,In_145,In_596);
and U1277 (N_1277,N_1021,N_739);
xor U1278 (N_1278,In_1282,In_877);
and U1279 (N_1279,In_1225,N_1006);
nand U1280 (N_1280,N_530,In_161);
nor U1281 (N_1281,In_918,N_1175);
nand U1282 (N_1282,In_972,N_983);
xnor U1283 (N_1283,In_74,N_431);
nand U1284 (N_1284,N_1088,N_311);
xnor U1285 (N_1285,N_831,N_1171);
nand U1286 (N_1286,In_533,N_1086);
nand U1287 (N_1287,N_524,N_950);
xnor U1288 (N_1288,In_1683,N_1130);
or U1289 (N_1289,N_1190,N_197);
or U1290 (N_1290,N_666,N_800);
nor U1291 (N_1291,N_1097,N_1126);
nand U1292 (N_1292,N_791,In_807);
or U1293 (N_1293,In_138,N_732);
xnor U1294 (N_1294,N_92,N_177);
and U1295 (N_1295,N_1029,N_1103);
or U1296 (N_1296,In_1491,N_987);
nand U1297 (N_1297,In_1085,N_981);
and U1298 (N_1298,N_899,N_1118);
xnor U1299 (N_1299,N_420,In_430);
nand U1300 (N_1300,N_440,N_1051);
and U1301 (N_1301,N_1059,In_998);
or U1302 (N_1302,In_557,N_1046);
nor U1303 (N_1303,In_1628,N_1166);
or U1304 (N_1304,N_112,N_1039);
and U1305 (N_1305,N_776,N_1003);
nand U1306 (N_1306,In_33,N_464);
xnor U1307 (N_1307,In_1893,In_541);
and U1308 (N_1308,In_837,In_1935);
xor U1309 (N_1309,In_784,N_1035);
and U1310 (N_1310,N_688,N_179);
xnor U1311 (N_1311,N_607,N_1065);
nor U1312 (N_1312,N_1095,N_302);
or U1313 (N_1313,In_692,N_1037);
nor U1314 (N_1314,N_883,N_69);
or U1315 (N_1315,N_1049,In_1072);
and U1316 (N_1316,N_1134,N_988);
nor U1317 (N_1317,N_1099,N_1008);
xnor U1318 (N_1318,N_379,N_1161);
nor U1319 (N_1319,In_3,In_9);
or U1320 (N_1320,N_216,N_594);
and U1321 (N_1321,N_1185,In_455);
or U1322 (N_1322,N_1163,In_363);
or U1323 (N_1323,N_1033,In_105);
nand U1324 (N_1324,N_725,N_753);
xnor U1325 (N_1325,In_1178,In_1965);
nand U1326 (N_1326,N_1176,In_443);
or U1327 (N_1327,N_1078,In_1527);
nor U1328 (N_1328,In_448,N_880);
and U1329 (N_1329,N_816,In_233);
and U1330 (N_1330,In_1955,In_1495);
or U1331 (N_1331,N_862,In_257);
xnor U1332 (N_1332,In_1887,N_1104);
nor U1333 (N_1333,N_1085,N_761);
nor U1334 (N_1334,N_979,N_784);
nand U1335 (N_1335,In_1531,In_1812);
or U1336 (N_1336,N_975,In_1026);
and U1337 (N_1337,N_490,In_928);
or U1338 (N_1338,In_1086,In_1317);
nor U1339 (N_1339,N_205,N_1152);
or U1340 (N_1340,N_823,In_372);
xnor U1341 (N_1341,N_1162,N_1158);
or U1342 (N_1342,In_453,N_1141);
nor U1343 (N_1343,N_1108,In_1834);
and U1344 (N_1344,In_1050,In_97);
or U1345 (N_1345,In_451,In_1798);
nor U1346 (N_1346,In_1184,N_767);
or U1347 (N_1347,In_365,In_22);
nor U1348 (N_1348,In_1544,N_759);
and U1349 (N_1349,N_1121,In_1850);
and U1350 (N_1350,In_1743,In_1172);
and U1351 (N_1351,In_330,In_166);
nand U1352 (N_1352,N_1147,N_714);
nor U1353 (N_1353,N_808,In_34);
nand U1354 (N_1354,N_113,N_1045);
xor U1355 (N_1355,In_941,In_1546);
nor U1356 (N_1356,N_1024,N_157);
or U1357 (N_1357,In_21,In_719);
nor U1358 (N_1358,N_588,N_1000);
or U1359 (N_1359,N_560,In_24);
and U1360 (N_1360,N_1013,N_763);
and U1361 (N_1361,In_1276,In_403);
xnor U1362 (N_1362,In_1825,N_1077);
or U1363 (N_1363,In_1705,N_294);
or U1364 (N_1364,N_630,N_1101);
nor U1365 (N_1365,N_1014,N_1071);
xor U1366 (N_1366,In_431,In_1828);
xnor U1367 (N_1367,N_973,N_673);
or U1368 (N_1368,N_834,In_1153);
or U1369 (N_1369,In_1313,In_1779);
and U1370 (N_1370,N_1012,N_1153);
xnor U1371 (N_1371,In_376,N_846);
xnor U1372 (N_1372,N_526,N_1094);
xnor U1373 (N_1373,N_1112,N_1170);
nor U1374 (N_1374,N_1067,N_30);
nand U1375 (N_1375,In_532,In_1568);
xnor U1376 (N_1376,In_289,In_1486);
nor U1377 (N_1377,In_840,In_1618);
nand U1378 (N_1378,In_953,In_1920);
and U1379 (N_1379,N_1084,N_1032);
and U1380 (N_1380,N_1005,N_810);
and U1381 (N_1381,N_18,N_854);
xnor U1382 (N_1382,N_1187,In_294);
or U1383 (N_1383,In_511,N_1042);
or U1384 (N_1384,In_892,N_649);
xor U1385 (N_1385,N_872,In_1466);
nand U1386 (N_1386,In_828,N_903);
or U1387 (N_1387,N_1004,N_927);
or U1388 (N_1388,N_1001,N_641);
nor U1389 (N_1389,N_1122,In_1140);
nor U1390 (N_1390,N_1142,N_996);
or U1391 (N_1391,In_1997,N_617);
and U1392 (N_1392,In_94,N_1154);
or U1393 (N_1393,In_554,N_881);
nand U1394 (N_1394,N_1117,N_408);
or U1395 (N_1395,In_1396,N_558);
nor U1396 (N_1396,N_1136,In_349);
xnor U1397 (N_1397,In_1558,N_1145);
nor U1398 (N_1398,In_1333,N_664);
xor U1399 (N_1399,In_1780,In_1519);
xor U1400 (N_1400,N_1174,N_1314);
nand U1401 (N_1401,N_1320,N_1106);
xnor U1402 (N_1402,N_986,N_968);
nand U1403 (N_1403,N_813,N_619);
nand U1404 (N_1404,In_136,N_1253);
nor U1405 (N_1405,N_959,N_1379);
or U1406 (N_1406,N_492,N_41);
and U1407 (N_1407,In_518,N_1207);
nor U1408 (N_1408,N_905,N_301);
nor U1409 (N_1409,N_1248,N_1260);
or U1410 (N_1410,In_471,N_1302);
xnor U1411 (N_1411,N_6,N_1089);
xnor U1412 (N_1412,N_863,N_240);
and U1413 (N_1413,N_743,N_757);
and U1414 (N_1414,N_1391,N_1301);
nor U1415 (N_1415,N_1374,N_1072);
or U1416 (N_1416,N_1334,N_213);
nand U1417 (N_1417,N_956,N_935);
nor U1418 (N_1418,N_1289,N_1274);
nor U1419 (N_1419,N_719,N_1393);
and U1420 (N_1420,N_1265,N_644);
or U1421 (N_1421,N_310,In_694);
nor U1422 (N_1422,N_597,N_124);
or U1423 (N_1423,N_0,N_1214);
nand U1424 (N_1424,N_1096,N_1266);
or U1425 (N_1425,In_1959,N_382);
or U1426 (N_1426,N_891,N_801);
nor U1427 (N_1427,N_1222,N_1354);
xnor U1428 (N_1428,In_159,N_1366);
nand U1429 (N_1429,N_750,In_1459);
nor U1430 (N_1430,In_769,N_1382);
xor U1431 (N_1431,N_837,In_657);
nor U1432 (N_1432,N_1198,N_1387);
nand U1433 (N_1433,In_1174,N_218);
nor U1434 (N_1434,N_1213,N_922);
and U1435 (N_1435,N_80,N_15);
and U1436 (N_1436,N_1116,N_821);
nand U1437 (N_1437,In_1694,N_1250);
nand U1438 (N_1438,N_264,In_870);
nand U1439 (N_1439,N_1295,N_1346);
or U1440 (N_1440,N_1237,In_1813);
xor U1441 (N_1441,N_1165,N_1337);
nor U1442 (N_1442,N_1203,N_1344);
and U1443 (N_1443,N_894,In_996);
nand U1444 (N_1444,N_637,In_420);
xor U1445 (N_1445,N_1234,In_500);
xnor U1446 (N_1446,In_1298,In_1852);
or U1447 (N_1447,In_906,N_733);
nor U1448 (N_1448,N_1212,N_1321);
nand U1449 (N_1449,In_698,N_1342);
xnor U1450 (N_1450,N_1256,N_858);
xnor U1451 (N_1451,N_1276,N_1364);
or U1452 (N_1452,N_1329,In_1840);
nand U1453 (N_1453,N_1197,N_1298);
nand U1454 (N_1454,N_1371,N_16);
xor U1455 (N_1455,N_202,N_1284);
xor U1456 (N_1456,N_469,N_775);
nor U1457 (N_1457,N_1223,In_969);
nand U1458 (N_1458,N_1381,N_1128);
xor U1459 (N_1459,N_1217,In_862);
and U1460 (N_1460,N_1319,N_457);
nand U1461 (N_1461,N_1209,N_671);
nand U1462 (N_1462,N_640,N_1394);
xnor U1463 (N_1463,N_832,N_912);
xor U1464 (N_1464,N_984,In_938);
xor U1465 (N_1465,N_900,N_1098);
nand U1466 (N_1466,In_222,N_1297);
xor U1467 (N_1467,In_1073,N_1351);
xnor U1468 (N_1468,N_1338,N_1306);
or U1469 (N_1469,In_1436,N_1249);
and U1470 (N_1470,In_1130,N_1247);
nand U1471 (N_1471,N_174,N_1129);
nand U1472 (N_1472,In_296,N_807);
nor U1473 (N_1473,N_1312,N_1375);
nand U1474 (N_1474,In_819,In_44);
or U1475 (N_1475,N_1370,N_1263);
or U1476 (N_1476,N_1277,In_1717);
xor U1477 (N_1477,N_1125,N_1058);
and U1478 (N_1478,N_1293,N_1041);
and U1479 (N_1479,N_1015,In_811);
xor U1480 (N_1480,In_1691,N_603);
or U1481 (N_1481,In_1356,N_584);
nand U1482 (N_1482,N_1020,N_914);
nand U1483 (N_1483,N_1324,N_1007);
nand U1484 (N_1484,In_465,N_623);
xor U1485 (N_1485,N_1056,N_1385);
nand U1486 (N_1486,N_116,N_1205);
nor U1487 (N_1487,N_1300,N_1144);
nand U1488 (N_1488,N_1189,N_1261);
nor U1489 (N_1489,N_1328,N_1357);
nand U1490 (N_1490,N_1349,In_190);
nand U1491 (N_1491,N_1360,N_423);
and U1492 (N_1492,N_1184,N_930);
and U1493 (N_1493,N_531,N_1243);
nor U1494 (N_1494,N_1119,N_1347);
nor U1495 (N_1495,N_1283,N_1373);
and U1496 (N_1496,In_1102,N_1164);
nor U1497 (N_1497,In_1416,N_1398);
and U1498 (N_1498,In_1977,In_1150);
and U1499 (N_1499,N_1386,N_712);
xnor U1500 (N_1500,N_610,N_726);
and U1501 (N_1501,N_1202,In_868);
or U1502 (N_1502,N_1307,N_1229);
and U1503 (N_1503,N_1057,N_1368);
xor U1504 (N_1504,N_994,N_1356);
xnor U1505 (N_1505,N_289,N_1390);
or U1506 (N_1506,N_544,N_674);
nand U1507 (N_1507,N_1155,In_1170);
and U1508 (N_1508,N_545,N_1228);
nor U1509 (N_1509,N_1038,N_596);
nand U1510 (N_1510,In_847,In_1160);
nand U1511 (N_1511,N_609,N_1350);
and U1512 (N_1512,N_827,In_1260);
nand U1513 (N_1513,N_1081,In_1727);
or U1514 (N_1514,N_150,N_1377);
nand U1515 (N_1515,N_1285,N_1227);
xor U1516 (N_1516,N_1028,N_1052);
xor U1517 (N_1517,N_329,N_1362);
xor U1518 (N_1518,N_1290,N_1221);
xor U1519 (N_1519,N_1127,N_1384);
and U1520 (N_1520,In_1602,N_1233);
and U1521 (N_1521,In_1362,N_877);
xor U1522 (N_1522,N_815,N_1367);
or U1523 (N_1523,N_625,In_1785);
or U1524 (N_1524,N_1255,N_826);
nor U1525 (N_1525,N_1009,N_1030);
xor U1526 (N_1526,N_48,N_1100);
nor U1527 (N_1527,N_283,N_448);
nand U1528 (N_1528,N_1199,N_1313);
nor U1529 (N_1529,N_1047,N_1218);
or U1530 (N_1530,N_875,N_1335);
xor U1531 (N_1531,In_8,N_1259);
or U1532 (N_1532,In_608,N_1040);
or U1533 (N_1533,In_1353,N_1280);
or U1534 (N_1534,N_1365,N_376);
xor U1535 (N_1535,N_247,N_258);
nor U1536 (N_1536,N_1339,N_402);
nor U1537 (N_1537,N_635,N_1010);
nand U1538 (N_1538,N_820,N_333);
nor U1539 (N_1539,In_1555,In_1414);
and U1540 (N_1540,N_1252,N_1181);
nand U1541 (N_1541,N_745,N_1241);
nor U1542 (N_1542,N_887,N_1341);
xnor U1543 (N_1543,In_258,N_645);
xor U1544 (N_1544,N_1389,N_1232);
and U1545 (N_1545,N_1193,N_508);
nor U1546 (N_1546,In_788,In_156);
nor U1547 (N_1547,N_1240,N_1017);
and U1548 (N_1548,N_1294,In_149);
xnor U1549 (N_1549,N_1192,N_521);
or U1550 (N_1550,N_1327,N_324);
nand U1551 (N_1551,N_443,N_1083);
nand U1552 (N_1552,N_1137,N_389);
and U1553 (N_1553,N_501,In_1421);
nor U1554 (N_1554,N_1069,In_1613);
nand U1555 (N_1555,N_629,N_1299);
or U1556 (N_1556,N_896,N_678);
nand U1557 (N_1557,N_1044,N_943);
nor U1558 (N_1558,In_1720,N_1262);
xor U1559 (N_1559,In_881,N_1022);
and U1560 (N_1560,N_1254,N_632);
and U1561 (N_1561,N_841,N_1323);
nor U1562 (N_1562,In_1457,In_849);
nand U1563 (N_1563,N_734,N_848);
xnor U1564 (N_1564,In_1861,N_945);
nor U1565 (N_1565,N_1143,N_576);
nor U1566 (N_1566,N_1031,N_901);
or U1567 (N_1567,N_1269,N_803);
or U1568 (N_1568,N_844,In_510);
nor U1569 (N_1569,N_1279,N_1278);
or U1570 (N_1570,N_682,In_305);
xor U1571 (N_1571,N_936,N_62);
or U1572 (N_1572,In_504,N_582);
nand U1573 (N_1573,N_1268,N_1288);
nand U1574 (N_1574,N_1235,N_895);
xnor U1575 (N_1575,N_1210,N_1109);
xnor U1576 (N_1576,N_1219,N_1080);
and U1577 (N_1577,N_976,In_1305);
xor U1578 (N_1578,N_785,N_52);
xnor U1579 (N_1579,In_486,N_1273);
nor U1580 (N_1580,N_500,N_1132);
and U1581 (N_1581,In_1984,N_1182);
xor U1582 (N_1582,N_1034,In_1426);
nor U1583 (N_1583,N_917,N_1332);
nand U1584 (N_1584,N_96,In_1204);
xor U1585 (N_1585,In_1441,N_924);
nand U1586 (N_1586,N_615,N_399);
nand U1587 (N_1587,N_1063,N_1206);
nand U1588 (N_1588,In_845,In_1689);
or U1589 (N_1589,N_1242,N_1348);
nand U1590 (N_1590,N_1244,In_407);
nor U1591 (N_1591,N_488,In_342);
nand U1592 (N_1592,N_1246,N_676);
nand U1593 (N_1593,In_757,In_1604);
xnor U1594 (N_1594,N_1194,N_368);
nand U1595 (N_1595,N_847,N_727);
nor U1596 (N_1596,N_1272,N_1216);
nor U1597 (N_1597,N_1316,N_796);
nor U1598 (N_1598,N_856,N_1076);
or U1599 (N_1599,N_161,In_1658);
and U1600 (N_1600,N_1588,N_1515);
or U1601 (N_1601,In_1234,N_192);
or U1602 (N_1602,N_1435,N_1447);
and U1603 (N_1603,N_1554,N_42);
xor U1604 (N_1604,N_1440,N_1343);
xor U1605 (N_1605,N_835,N_897);
nand U1606 (N_1606,N_1565,N_1405);
nor U1607 (N_1607,N_1423,N_1510);
and U1608 (N_1608,In_1488,N_1359);
nand U1609 (N_1609,N_1023,N_1540);
nand U1610 (N_1610,N_1408,N_1446);
or U1611 (N_1611,N_1455,N_965);
nor U1612 (N_1612,N_1491,N_1545);
xor U1613 (N_1613,N_709,N_31);
xnor U1614 (N_1614,N_1534,N_1204);
or U1615 (N_1615,N_1431,In_295);
and U1616 (N_1616,N_1011,In_29);
and U1617 (N_1617,N_172,N_1475);
or U1618 (N_1618,N_1522,In_732);
nand U1619 (N_1619,N_1506,N_911);
and U1620 (N_1620,N_1133,In_595);
nand U1621 (N_1621,N_1562,In_699);
xor U1622 (N_1622,N_1597,N_1102);
nand U1623 (N_1623,N_1492,N_1043);
xor U1624 (N_1624,N_1572,N_910);
xnor U1625 (N_1625,N_1512,N_1002);
nand U1626 (N_1626,In_639,N_1392);
and U1627 (N_1627,N_1231,N_1518);
and U1628 (N_1628,N_1050,N_1589);
xor U1629 (N_1629,N_1401,N_1383);
and U1630 (N_1630,N_1548,N_1201);
nor U1631 (N_1631,N_1418,N_1448);
and U1632 (N_1632,N_1521,N_1535);
nand U1633 (N_1633,N_680,N_951);
xnor U1634 (N_1634,N_1587,N_1457);
or U1635 (N_1635,N_1483,N_1497);
nand U1636 (N_1636,N_1404,N_1411);
nor U1637 (N_1637,N_1333,N_1578);
or U1638 (N_1638,N_1480,N_180);
and U1639 (N_1639,N_668,N_261);
and U1640 (N_1640,N_1464,N_888);
and U1641 (N_1641,N_1225,In_1064);
and U1642 (N_1642,In_43,N_1159);
nand U1643 (N_1643,N_1476,N_1507);
xor U1644 (N_1644,N_126,N_1511);
nor U1645 (N_1645,N_1286,N_1317);
nand U1646 (N_1646,N_199,N_589);
or U1647 (N_1647,N_1442,N_1353);
nand U1648 (N_1648,N_1358,N_1558);
nand U1649 (N_1649,In_1651,N_1478);
nor U1650 (N_1650,N_1264,N_1211);
nand U1651 (N_1651,N_1437,In_1092);
or U1652 (N_1652,N_1490,N_1528);
and U1653 (N_1653,N_669,N_1598);
or U1654 (N_1654,N_1474,N_1520);
xnor U1655 (N_1655,N_1179,N_1585);
nor U1656 (N_1656,N_1477,N_1361);
or U1657 (N_1657,N_717,N_1586);
xnor U1658 (N_1658,N_1527,N_1533);
or U1659 (N_1659,In_859,N_948);
or U1660 (N_1660,In_1748,N_1516);
xnor U1661 (N_1661,N_1482,N_1458);
xor U1662 (N_1662,N_923,N_1131);
and U1663 (N_1663,In_1247,N_1060);
xor U1664 (N_1664,N_1326,In_874);
or U1665 (N_1665,N_1593,N_1525);
or U1666 (N_1666,N_1267,N_1168);
and U1667 (N_1667,N_1574,N_1336);
or U1668 (N_1668,N_1581,N_1547);
nand U1669 (N_1669,N_1413,N_697);
or U1670 (N_1670,N_1399,N_1462);
nor U1671 (N_1671,N_1544,N_728);
xnor U1672 (N_1672,N_1257,N_1546);
nor U1673 (N_1673,N_1526,N_1173);
nand U1674 (N_1674,N_1303,N_1239);
or U1675 (N_1675,N_1465,N_1496);
and U1676 (N_1676,N_1503,N_990);
nor U1677 (N_1677,N_1275,N_1538);
nor U1678 (N_1678,N_1509,N_1400);
xnor U1679 (N_1679,N_1236,N_1556);
nand U1680 (N_1680,N_1270,N_1456);
or U1681 (N_1681,N_1550,N_1555);
nand U1682 (N_1682,N_1433,N_716);
nand U1683 (N_1683,N_1582,N_1524);
nor U1684 (N_1684,N_991,N_1310);
xor U1685 (N_1685,N_1472,N_1463);
or U1686 (N_1686,N_613,N_1479);
nor U1687 (N_1687,N_1568,N_1070);
nor U1688 (N_1688,N_1559,In_755);
and U1689 (N_1689,In_409,N_1372);
xor U1690 (N_1690,N_1466,N_316);
or U1691 (N_1691,N_1592,N_1498);
nand U1692 (N_1692,N_1066,In_1116);
or U1693 (N_1693,N_652,N_1577);
nand U1694 (N_1694,N_970,N_1151);
or U1695 (N_1695,N_1410,N_1473);
xnor U1696 (N_1696,N_1517,N_1595);
xnor U1697 (N_1697,In_178,N_1426);
nand U1698 (N_1698,N_1549,N_1495);
and U1699 (N_1699,N_1191,In_776);
xor U1700 (N_1700,N_1018,In_125);
nor U1701 (N_1701,N_1226,In_519);
nand U1702 (N_1702,N_1493,N_1397);
and U1703 (N_1703,N_1484,N_1331);
nand U1704 (N_1704,N_1530,N_1443);
nand U1705 (N_1705,N_575,N_1599);
nor U1706 (N_1706,N_1315,N_1238);
nand U1707 (N_1707,N_1571,N_1460);
or U1708 (N_1708,N_1092,N_1432);
nand U1709 (N_1709,N_1318,In_1031);
and U1710 (N_1710,N_1407,N_85);
or U1711 (N_1711,N_1563,N_1296);
nand U1712 (N_1712,N_1591,N_1486);
nand U1713 (N_1713,N_1224,N_1489);
and U1714 (N_1714,N_1420,N_1501);
xor U1715 (N_1715,N_1566,In_690);
or U1716 (N_1716,N_1459,N_1552);
or U1717 (N_1717,N_1468,N_773);
xor U1718 (N_1718,N_1355,N_1580);
xor U1719 (N_1719,N_1519,N_1414);
and U1720 (N_1720,N_1287,N_1430);
nand U1721 (N_1721,N_1541,N_993);
xor U1722 (N_1722,N_1412,N_1093);
xor U1723 (N_1723,N_1230,N_1502);
or U1724 (N_1724,N_239,N_1363);
nor U1725 (N_1725,N_1454,N_1445);
nor U1726 (N_1726,N_1395,N_692);
nand U1727 (N_1727,N_1505,In_134);
and U1728 (N_1728,N_1513,N_1451);
nor U1729 (N_1729,N_1471,N_1245);
xor U1730 (N_1730,N_1149,In_1548);
xnor U1731 (N_1731,N_1322,In_36);
nor U1732 (N_1732,N_1499,N_1584);
nand U1733 (N_1733,N_650,N_57);
nand U1734 (N_1734,N_1258,N_1564);
and U1735 (N_1735,N_1380,In_1822);
nor U1736 (N_1736,N_1500,N_1352);
nor U1737 (N_1737,In_835,N_1396);
xor U1738 (N_1738,N_1543,N_916);
and U1739 (N_1739,N_1345,N_1402);
and U1740 (N_1740,N_1304,N_802);
nor U1741 (N_1741,N_1325,N_1531);
and U1742 (N_1742,N_1438,N_904);
xor U1743 (N_1743,N_1376,N_1330);
or U1744 (N_1744,N_742,N_1583);
nor U1745 (N_1745,N_354,N_1388);
nor U1746 (N_1746,N_1208,N_1409);
xor U1747 (N_1747,N_762,N_926);
nand U1748 (N_1748,N_1282,N_479);
nand U1749 (N_1749,N_1470,In_223);
nor U1750 (N_1750,N_1421,N_1441);
xnor U1751 (N_1751,N_1569,N_1429);
nand U1752 (N_1752,N_1292,N_1439);
or U1753 (N_1753,N_1140,N_839);
nand U1754 (N_1754,N_1532,N_1449);
xnor U1755 (N_1755,N_362,N_1419);
nand U1756 (N_1756,N_1428,N_1415);
or U1757 (N_1757,N_812,N_1579);
nand U1758 (N_1758,N_204,N_1485);
and U1759 (N_1759,N_1557,N_1271);
nand U1760 (N_1760,N_1529,N_1369);
and U1761 (N_1761,N_1573,N_1074);
nor U1762 (N_1762,N_1054,N_1417);
and U1763 (N_1763,N_1427,N_1575);
or U1764 (N_1764,N_1453,N_1305);
and U1765 (N_1765,N_622,In_1020);
nor U1766 (N_1766,N_1536,N_84);
and U1767 (N_1767,N_1488,N_1561);
and U1768 (N_1768,N_1570,N_1403);
and U1769 (N_1769,In_824,N_1281);
xor U1770 (N_1770,N_780,N_1514);
and U1771 (N_1771,N_143,N_1537);
nand U1772 (N_1772,In_357,N_1450);
nand U1773 (N_1773,N_876,N_1215);
or U1774 (N_1774,N_1481,N_1291);
nor U1775 (N_1775,N_1172,N_1553);
xnor U1776 (N_1776,N_1560,N_631);
and U1777 (N_1777,N_1177,N_828);
or U1778 (N_1778,N_1504,N_1111);
or U1779 (N_1779,N_1434,N_1424);
or U1780 (N_1780,N_1425,N_1200);
nor U1781 (N_1781,N_1406,N_1461);
or U1782 (N_1782,In_908,N_1452);
xnor U1783 (N_1783,N_1309,In_1999);
and U1784 (N_1784,N_1487,N_1444);
and U1785 (N_1785,N_1340,N_1308);
xor U1786 (N_1786,N_599,N_1539);
and U1787 (N_1787,N_1551,N_1467);
nor U1788 (N_1788,N_1508,N_1494);
and U1789 (N_1789,N_1567,N_1220);
nor U1790 (N_1790,N_1576,N_1542);
xnor U1791 (N_1791,N_1062,In_1942);
or U1792 (N_1792,N_1523,N_867);
nand U1793 (N_1793,N_1311,N_587);
xor U1794 (N_1794,N_1251,N_1590);
or U1795 (N_1795,N_1422,N_1469);
xnor U1796 (N_1796,N_1596,N_107);
and U1797 (N_1797,N_445,N_556);
xor U1798 (N_1798,N_1594,N_1416);
nor U1799 (N_1799,N_1436,N_1378);
nand U1800 (N_1800,N_1771,N_1790);
xor U1801 (N_1801,N_1751,N_1735);
nand U1802 (N_1802,N_1776,N_1770);
nand U1803 (N_1803,N_1747,N_1797);
and U1804 (N_1804,N_1772,N_1664);
xor U1805 (N_1805,N_1684,N_1625);
and U1806 (N_1806,N_1673,N_1713);
nor U1807 (N_1807,N_1662,N_1659);
and U1808 (N_1808,N_1666,N_1697);
nand U1809 (N_1809,N_1668,N_1781);
and U1810 (N_1810,N_1779,N_1694);
xnor U1811 (N_1811,N_1628,N_1686);
nand U1812 (N_1812,N_1765,N_1729);
nor U1813 (N_1813,N_1602,N_1691);
nand U1814 (N_1814,N_1639,N_1665);
and U1815 (N_1815,N_1792,N_1796);
xnor U1816 (N_1816,N_1682,N_1646);
and U1817 (N_1817,N_1676,N_1726);
xor U1818 (N_1818,N_1670,N_1657);
nand U1819 (N_1819,N_1623,N_1611);
nor U1820 (N_1820,N_1711,N_1741);
or U1821 (N_1821,N_1632,N_1702);
nand U1822 (N_1822,N_1614,N_1718);
or U1823 (N_1823,N_1696,N_1672);
nor U1824 (N_1824,N_1638,N_1758);
nand U1825 (N_1825,N_1620,N_1653);
nor U1826 (N_1826,N_1730,N_1685);
xor U1827 (N_1827,N_1734,N_1783);
nand U1828 (N_1828,N_1701,N_1642);
and U1829 (N_1829,N_1759,N_1608);
nor U1830 (N_1830,N_1724,N_1645);
nand U1831 (N_1831,N_1733,N_1615);
xnor U1832 (N_1832,N_1660,N_1667);
or U1833 (N_1833,N_1731,N_1703);
xor U1834 (N_1834,N_1795,N_1762);
xnor U1835 (N_1835,N_1785,N_1798);
xor U1836 (N_1836,N_1763,N_1761);
nand U1837 (N_1837,N_1725,N_1777);
and U1838 (N_1838,N_1636,N_1606);
or U1839 (N_1839,N_1786,N_1788);
xor U1840 (N_1840,N_1656,N_1743);
nor U1841 (N_1841,N_1610,N_1768);
or U1842 (N_1842,N_1603,N_1706);
nor U1843 (N_1843,N_1756,N_1669);
xor U1844 (N_1844,N_1630,N_1720);
nand U1845 (N_1845,N_1654,N_1683);
and U1846 (N_1846,N_1722,N_1626);
or U1847 (N_1847,N_1704,N_1717);
xor U1848 (N_1848,N_1690,N_1738);
xor U1849 (N_1849,N_1641,N_1681);
nand U1850 (N_1850,N_1742,N_1732);
nand U1851 (N_1851,N_1671,N_1794);
or U1852 (N_1852,N_1631,N_1647);
and U1853 (N_1853,N_1661,N_1746);
xor U1854 (N_1854,N_1616,N_1739);
nor U1855 (N_1855,N_1736,N_1752);
and U1856 (N_1856,N_1708,N_1687);
nand U1857 (N_1857,N_1754,N_1799);
nor U1858 (N_1858,N_1760,N_1705);
nand U1859 (N_1859,N_1793,N_1658);
or U1860 (N_1860,N_1710,N_1714);
and U1861 (N_1861,N_1605,N_1663);
and U1862 (N_1862,N_1778,N_1688);
or U1863 (N_1863,N_1774,N_1728);
nor U1864 (N_1864,N_1692,N_1755);
nand U1865 (N_1865,N_1624,N_1753);
or U1866 (N_1866,N_1723,N_1695);
xor U1867 (N_1867,N_1745,N_1601);
nor U1868 (N_1868,N_1627,N_1727);
nor U1869 (N_1869,N_1679,N_1600);
xor U1870 (N_1870,N_1675,N_1634);
xor U1871 (N_1871,N_1775,N_1643);
xnor U1872 (N_1872,N_1716,N_1749);
xnor U1873 (N_1873,N_1678,N_1782);
xnor U1874 (N_1874,N_1640,N_1650);
nor U1875 (N_1875,N_1621,N_1607);
or U1876 (N_1876,N_1791,N_1644);
or U1877 (N_1877,N_1712,N_1709);
xnor U1878 (N_1878,N_1674,N_1612);
nor U1879 (N_1879,N_1748,N_1744);
or U1880 (N_1880,N_1764,N_1617);
xnor U1881 (N_1881,N_1707,N_1689);
and U1882 (N_1882,N_1757,N_1719);
xor U1883 (N_1883,N_1699,N_1789);
or U1884 (N_1884,N_1773,N_1700);
xnor U1885 (N_1885,N_1784,N_1649);
xor U1886 (N_1886,N_1780,N_1740);
and U1887 (N_1887,N_1619,N_1613);
or U1888 (N_1888,N_1787,N_1635);
nor U1889 (N_1889,N_1651,N_1769);
or U1890 (N_1890,N_1637,N_1609);
nand U1891 (N_1891,N_1677,N_1767);
nor U1892 (N_1892,N_1648,N_1652);
xor U1893 (N_1893,N_1604,N_1633);
xor U1894 (N_1894,N_1715,N_1766);
or U1895 (N_1895,N_1680,N_1698);
nor U1896 (N_1896,N_1750,N_1629);
nand U1897 (N_1897,N_1618,N_1737);
nor U1898 (N_1898,N_1693,N_1655);
xnor U1899 (N_1899,N_1622,N_1721);
nand U1900 (N_1900,N_1746,N_1791);
and U1901 (N_1901,N_1617,N_1725);
xor U1902 (N_1902,N_1785,N_1646);
and U1903 (N_1903,N_1753,N_1730);
nor U1904 (N_1904,N_1686,N_1664);
nand U1905 (N_1905,N_1791,N_1647);
xor U1906 (N_1906,N_1776,N_1715);
xnor U1907 (N_1907,N_1719,N_1703);
nor U1908 (N_1908,N_1770,N_1700);
nand U1909 (N_1909,N_1773,N_1645);
nor U1910 (N_1910,N_1788,N_1618);
and U1911 (N_1911,N_1625,N_1624);
nor U1912 (N_1912,N_1679,N_1653);
nand U1913 (N_1913,N_1706,N_1768);
nand U1914 (N_1914,N_1613,N_1685);
xor U1915 (N_1915,N_1754,N_1756);
and U1916 (N_1916,N_1710,N_1784);
nand U1917 (N_1917,N_1644,N_1790);
nand U1918 (N_1918,N_1753,N_1610);
or U1919 (N_1919,N_1709,N_1718);
nor U1920 (N_1920,N_1773,N_1706);
xnor U1921 (N_1921,N_1720,N_1714);
nor U1922 (N_1922,N_1645,N_1732);
nor U1923 (N_1923,N_1656,N_1626);
or U1924 (N_1924,N_1643,N_1613);
xor U1925 (N_1925,N_1701,N_1750);
and U1926 (N_1926,N_1673,N_1697);
and U1927 (N_1927,N_1640,N_1682);
nand U1928 (N_1928,N_1684,N_1681);
and U1929 (N_1929,N_1738,N_1661);
and U1930 (N_1930,N_1776,N_1638);
xor U1931 (N_1931,N_1637,N_1756);
or U1932 (N_1932,N_1750,N_1666);
or U1933 (N_1933,N_1710,N_1791);
and U1934 (N_1934,N_1748,N_1669);
nand U1935 (N_1935,N_1613,N_1681);
and U1936 (N_1936,N_1789,N_1654);
xor U1937 (N_1937,N_1663,N_1686);
and U1938 (N_1938,N_1676,N_1759);
nor U1939 (N_1939,N_1674,N_1631);
xor U1940 (N_1940,N_1634,N_1667);
and U1941 (N_1941,N_1755,N_1673);
or U1942 (N_1942,N_1705,N_1759);
or U1943 (N_1943,N_1656,N_1726);
or U1944 (N_1944,N_1673,N_1771);
nand U1945 (N_1945,N_1782,N_1778);
or U1946 (N_1946,N_1702,N_1674);
and U1947 (N_1947,N_1652,N_1665);
and U1948 (N_1948,N_1709,N_1784);
xor U1949 (N_1949,N_1775,N_1710);
nor U1950 (N_1950,N_1764,N_1695);
or U1951 (N_1951,N_1641,N_1753);
nor U1952 (N_1952,N_1666,N_1712);
and U1953 (N_1953,N_1725,N_1685);
nor U1954 (N_1954,N_1758,N_1749);
nand U1955 (N_1955,N_1685,N_1673);
xnor U1956 (N_1956,N_1716,N_1720);
and U1957 (N_1957,N_1735,N_1764);
xnor U1958 (N_1958,N_1731,N_1682);
xnor U1959 (N_1959,N_1783,N_1788);
or U1960 (N_1960,N_1754,N_1791);
and U1961 (N_1961,N_1615,N_1640);
nand U1962 (N_1962,N_1730,N_1769);
or U1963 (N_1963,N_1657,N_1635);
or U1964 (N_1964,N_1760,N_1660);
and U1965 (N_1965,N_1796,N_1780);
xor U1966 (N_1966,N_1622,N_1756);
and U1967 (N_1967,N_1704,N_1694);
nor U1968 (N_1968,N_1757,N_1630);
or U1969 (N_1969,N_1712,N_1763);
xor U1970 (N_1970,N_1660,N_1601);
or U1971 (N_1971,N_1766,N_1795);
and U1972 (N_1972,N_1713,N_1615);
nor U1973 (N_1973,N_1654,N_1721);
or U1974 (N_1974,N_1782,N_1679);
xor U1975 (N_1975,N_1605,N_1718);
nor U1976 (N_1976,N_1765,N_1799);
or U1977 (N_1977,N_1676,N_1705);
and U1978 (N_1978,N_1720,N_1660);
xnor U1979 (N_1979,N_1632,N_1601);
nor U1980 (N_1980,N_1726,N_1729);
or U1981 (N_1981,N_1685,N_1770);
or U1982 (N_1982,N_1751,N_1697);
and U1983 (N_1983,N_1640,N_1717);
xnor U1984 (N_1984,N_1765,N_1625);
and U1985 (N_1985,N_1762,N_1730);
xor U1986 (N_1986,N_1754,N_1619);
or U1987 (N_1987,N_1768,N_1657);
nand U1988 (N_1988,N_1642,N_1644);
nor U1989 (N_1989,N_1673,N_1705);
xnor U1990 (N_1990,N_1614,N_1646);
and U1991 (N_1991,N_1670,N_1600);
nor U1992 (N_1992,N_1638,N_1799);
or U1993 (N_1993,N_1707,N_1731);
or U1994 (N_1994,N_1788,N_1676);
nor U1995 (N_1995,N_1713,N_1775);
or U1996 (N_1996,N_1612,N_1768);
or U1997 (N_1997,N_1670,N_1651);
xor U1998 (N_1998,N_1630,N_1756);
nor U1999 (N_1999,N_1671,N_1634);
nor U2000 (N_2000,N_1825,N_1899);
and U2001 (N_2001,N_1816,N_1819);
xnor U2002 (N_2002,N_1911,N_1834);
xor U2003 (N_2003,N_1939,N_1809);
and U2004 (N_2004,N_1996,N_1821);
or U2005 (N_2005,N_1919,N_1949);
and U2006 (N_2006,N_1833,N_1804);
xor U2007 (N_2007,N_1995,N_1893);
nand U2008 (N_2008,N_1997,N_1922);
and U2009 (N_2009,N_1965,N_1993);
or U2010 (N_2010,N_1946,N_1843);
nor U2011 (N_2011,N_1879,N_1916);
nor U2012 (N_2012,N_1813,N_1971);
nor U2013 (N_2013,N_1953,N_1978);
nand U2014 (N_2014,N_1865,N_1969);
or U2015 (N_2015,N_1906,N_1944);
nand U2016 (N_2016,N_1923,N_1989);
or U2017 (N_2017,N_1856,N_1930);
or U2018 (N_2018,N_1991,N_1839);
xnor U2019 (N_2019,N_1961,N_1942);
xor U2020 (N_2020,N_1860,N_1814);
nand U2021 (N_2021,N_1844,N_1847);
or U2022 (N_2022,N_1849,N_1895);
and U2023 (N_2023,N_1818,N_1884);
or U2024 (N_2024,N_1917,N_1842);
nand U2025 (N_2025,N_1886,N_1876);
or U2026 (N_2026,N_1940,N_1905);
and U2027 (N_2027,N_1822,N_1963);
nand U2028 (N_2028,N_1948,N_1840);
nand U2029 (N_2029,N_1875,N_1850);
or U2030 (N_2030,N_1950,N_1861);
xor U2031 (N_2031,N_1897,N_1921);
nand U2032 (N_2032,N_1907,N_1896);
xnor U2033 (N_2033,N_1877,N_1970);
nand U2034 (N_2034,N_1885,N_1859);
and U2035 (N_2035,N_1867,N_1951);
and U2036 (N_2036,N_1932,N_1851);
nand U2037 (N_2037,N_1976,N_1864);
nor U2038 (N_2038,N_1880,N_1947);
and U2039 (N_2039,N_1881,N_1854);
xnor U2040 (N_2040,N_1824,N_1988);
nor U2041 (N_2041,N_1987,N_1898);
nand U2042 (N_2042,N_1831,N_1964);
nand U2043 (N_2043,N_1980,N_1914);
and U2044 (N_2044,N_1926,N_1928);
or U2045 (N_2045,N_1841,N_1887);
and U2046 (N_2046,N_1832,N_1852);
xor U2047 (N_2047,N_1837,N_1869);
nor U2048 (N_2048,N_1909,N_1938);
nand U2049 (N_2049,N_1853,N_1800);
nand U2050 (N_2050,N_1845,N_1977);
or U2051 (N_2051,N_1857,N_1878);
nor U2052 (N_2052,N_1998,N_1983);
nor U2053 (N_2053,N_1966,N_1812);
or U2054 (N_2054,N_1913,N_1872);
and U2055 (N_2055,N_1962,N_1858);
and U2056 (N_2056,N_1904,N_1918);
nand U2057 (N_2057,N_1943,N_1890);
xor U2058 (N_2058,N_1982,N_1945);
or U2059 (N_2059,N_1915,N_1894);
nor U2060 (N_2060,N_1836,N_1941);
xnor U2061 (N_2061,N_1830,N_1929);
nand U2062 (N_2062,N_1810,N_1855);
and U2063 (N_2063,N_1954,N_1925);
nor U2064 (N_2064,N_1817,N_1827);
or U2065 (N_2065,N_1972,N_1815);
and U2066 (N_2066,N_1957,N_1870);
and U2067 (N_2067,N_1912,N_1927);
xnor U2068 (N_2068,N_1882,N_1900);
or U2069 (N_2069,N_1955,N_1888);
or U2070 (N_2070,N_1873,N_1807);
nand U2071 (N_2071,N_1935,N_1958);
and U2072 (N_2072,N_1868,N_1892);
or U2073 (N_2073,N_1986,N_1866);
nand U2074 (N_2074,N_1838,N_1826);
nand U2075 (N_2075,N_1973,N_1979);
nand U2076 (N_2076,N_1863,N_1828);
nor U2077 (N_2077,N_1975,N_1981);
nand U2078 (N_2078,N_1937,N_1967);
or U2079 (N_2079,N_1903,N_1801);
nand U2080 (N_2080,N_1891,N_1985);
and U2081 (N_2081,N_1811,N_1823);
xnor U2082 (N_2082,N_1910,N_1999);
nor U2083 (N_2083,N_1902,N_1901);
nor U2084 (N_2084,N_1862,N_1803);
xnor U2085 (N_2085,N_1920,N_1924);
and U2086 (N_2086,N_1805,N_1933);
or U2087 (N_2087,N_1874,N_1934);
nand U2088 (N_2088,N_1931,N_1883);
nor U2089 (N_2089,N_1848,N_1956);
or U2090 (N_2090,N_1952,N_1806);
xor U2091 (N_2091,N_1889,N_1820);
xnor U2092 (N_2092,N_1968,N_1992);
or U2093 (N_2093,N_1829,N_1994);
xnor U2094 (N_2094,N_1960,N_1990);
nor U2095 (N_2095,N_1984,N_1871);
and U2096 (N_2096,N_1846,N_1936);
nor U2097 (N_2097,N_1908,N_1808);
nand U2098 (N_2098,N_1959,N_1835);
nand U2099 (N_2099,N_1802,N_1974);
and U2100 (N_2100,N_1818,N_1906);
nand U2101 (N_2101,N_1908,N_1973);
xor U2102 (N_2102,N_1966,N_1950);
or U2103 (N_2103,N_1948,N_1982);
nand U2104 (N_2104,N_1878,N_1901);
nand U2105 (N_2105,N_1823,N_1942);
xor U2106 (N_2106,N_1998,N_1952);
or U2107 (N_2107,N_1886,N_1821);
nand U2108 (N_2108,N_1875,N_1999);
nor U2109 (N_2109,N_1847,N_1853);
nand U2110 (N_2110,N_1902,N_1918);
nor U2111 (N_2111,N_1897,N_1833);
nor U2112 (N_2112,N_1821,N_1964);
and U2113 (N_2113,N_1918,N_1896);
nand U2114 (N_2114,N_1967,N_1893);
xor U2115 (N_2115,N_1997,N_1886);
nor U2116 (N_2116,N_1898,N_1934);
and U2117 (N_2117,N_1824,N_1844);
nor U2118 (N_2118,N_1958,N_1962);
or U2119 (N_2119,N_1915,N_1883);
nor U2120 (N_2120,N_1957,N_1950);
and U2121 (N_2121,N_1811,N_1981);
nor U2122 (N_2122,N_1973,N_1969);
or U2123 (N_2123,N_1983,N_1984);
nand U2124 (N_2124,N_1812,N_1984);
nand U2125 (N_2125,N_1885,N_1889);
xnor U2126 (N_2126,N_1833,N_1914);
and U2127 (N_2127,N_1842,N_1853);
nor U2128 (N_2128,N_1820,N_1877);
or U2129 (N_2129,N_1874,N_1891);
nand U2130 (N_2130,N_1947,N_1802);
and U2131 (N_2131,N_1816,N_1978);
nor U2132 (N_2132,N_1968,N_1910);
nand U2133 (N_2133,N_1935,N_1839);
xnor U2134 (N_2134,N_1874,N_1830);
and U2135 (N_2135,N_1966,N_1878);
xor U2136 (N_2136,N_1918,N_1934);
and U2137 (N_2137,N_1883,N_1947);
nand U2138 (N_2138,N_1953,N_1827);
xor U2139 (N_2139,N_1835,N_1942);
xor U2140 (N_2140,N_1816,N_1976);
nor U2141 (N_2141,N_1984,N_1891);
or U2142 (N_2142,N_1939,N_1810);
nand U2143 (N_2143,N_1912,N_1896);
xor U2144 (N_2144,N_1802,N_1849);
nand U2145 (N_2145,N_1903,N_1978);
and U2146 (N_2146,N_1992,N_1983);
nor U2147 (N_2147,N_1840,N_1921);
xnor U2148 (N_2148,N_1871,N_1941);
and U2149 (N_2149,N_1811,N_1936);
and U2150 (N_2150,N_1986,N_1819);
xor U2151 (N_2151,N_1835,N_1824);
or U2152 (N_2152,N_1927,N_1805);
and U2153 (N_2153,N_1822,N_1973);
xor U2154 (N_2154,N_1990,N_1995);
and U2155 (N_2155,N_1992,N_1964);
nand U2156 (N_2156,N_1968,N_1979);
xor U2157 (N_2157,N_1898,N_1902);
nand U2158 (N_2158,N_1809,N_1868);
nor U2159 (N_2159,N_1958,N_1971);
and U2160 (N_2160,N_1948,N_1827);
nand U2161 (N_2161,N_1813,N_1825);
or U2162 (N_2162,N_1846,N_1875);
nor U2163 (N_2163,N_1965,N_1961);
nor U2164 (N_2164,N_1804,N_1840);
xnor U2165 (N_2165,N_1841,N_1804);
nand U2166 (N_2166,N_1842,N_1966);
nor U2167 (N_2167,N_1852,N_1937);
or U2168 (N_2168,N_1933,N_1926);
nor U2169 (N_2169,N_1876,N_1827);
nand U2170 (N_2170,N_1980,N_1956);
nand U2171 (N_2171,N_1965,N_1825);
xor U2172 (N_2172,N_1809,N_1808);
xor U2173 (N_2173,N_1899,N_1861);
nor U2174 (N_2174,N_1802,N_1801);
xor U2175 (N_2175,N_1952,N_1951);
or U2176 (N_2176,N_1951,N_1810);
nor U2177 (N_2177,N_1879,N_1825);
and U2178 (N_2178,N_1831,N_1901);
and U2179 (N_2179,N_1854,N_1829);
xor U2180 (N_2180,N_1808,N_1964);
and U2181 (N_2181,N_1872,N_1844);
xnor U2182 (N_2182,N_1939,N_1947);
nor U2183 (N_2183,N_1924,N_1838);
xnor U2184 (N_2184,N_1925,N_1871);
and U2185 (N_2185,N_1972,N_1981);
nand U2186 (N_2186,N_1964,N_1885);
and U2187 (N_2187,N_1800,N_1938);
or U2188 (N_2188,N_1860,N_1818);
or U2189 (N_2189,N_1841,N_1907);
and U2190 (N_2190,N_1845,N_1882);
nand U2191 (N_2191,N_1939,N_1896);
nand U2192 (N_2192,N_1999,N_1991);
nor U2193 (N_2193,N_1867,N_1844);
xor U2194 (N_2194,N_1938,N_1990);
and U2195 (N_2195,N_1839,N_1903);
xnor U2196 (N_2196,N_1922,N_1897);
and U2197 (N_2197,N_1827,N_1894);
xor U2198 (N_2198,N_1898,N_1880);
nor U2199 (N_2199,N_1939,N_1948);
nor U2200 (N_2200,N_2100,N_2083);
and U2201 (N_2201,N_2085,N_2109);
or U2202 (N_2202,N_2144,N_2098);
nand U2203 (N_2203,N_2192,N_2147);
nor U2204 (N_2204,N_2034,N_2165);
nand U2205 (N_2205,N_2045,N_2102);
nand U2206 (N_2206,N_2078,N_2017);
xor U2207 (N_2207,N_2193,N_2051);
xnor U2208 (N_2208,N_2068,N_2152);
nor U2209 (N_2209,N_2110,N_2107);
and U2210 (N_2210,N_2059,N_2028);
xor U2211 (N_2211,N_2025,N_2127);
nor U2212 (N_2212,N_2148,N_2096);
xnor U2213 (N_2213,N_2125,N_2174);
or U2214 (N_2214,N_2021,N_2139);
xor U2215 (N_2215,N_2114,N_2159);
or U2216 (N_2216,N_2189,N_2044);
nor U2217 (N_2217,N_2160,N_2095);
xor U2218 (N_2218,N_2116,N_2119);
and U2219 (N_2219,N_2161,N_2141);
nand U2220 (N_2220,N_2128,N_2185);
or U2221 (N_2221,N_2060,N_2167);
nand U2222 (N_2222,N_2092,N_2108);
nand U2223 (N_2223,N_2040,N_2093);
and U2224 (N_2224,N_2135,N_2081);
and U2225 (N_2225,N_2063,N_2099);
and U2226 (N_2226,N_2074,N_2122);
or U2227 (N_2227,N_2084,N_2169);
xnor U2228 (N_2228,N_2073,N_2052);
nor U2229 (N_2229,N_2010,N_2123);
and U2230 (N_2230,N_2055,N_2146);
nand U2231 (N_2231,N_2187,N_2004);
xor U2232 (N_2232,N_2130,N_2050);
or U2233 (N_2233,N_2039,N_2069);
and U2234 (N_2234,N_2168,N_2163);
nor U2235 (N_2235,N_2032,N_2138);
and U2236 (N_2236,N_2105,N_2140);
nand U2237 (N_2237,N_2196,N_2118);
or U2238 (N_2238,N_2019,N_2006);
xnor U2239 (N_2239,N_2000,N_2106);
nand U2240 (N_2240,N_2191,N_2067);
and U2241 (N_2241,N_2178,N_2070);
nor U2242 (N_2242,N_2183,N_2195);
nand U2243 (N_2243,N_2120,N_2077);
nand U2244 (N_2244,N_2053,N_2037);
xor U2245 (N_2245,N_2023,N_2090);
nand U2246 (N_2246,N_2186,N_2031);
nor U2247 (N_2247,N_2132,N_2065);
nand U2248 (N_2248,N_2143,N_2057);
and U2249 (N_2249,N_2011,N_2030);
nand U2250 (N_2250,N_2166,N_2181);
xor U2251 (N_2251,N_2058,N_2054);
or U2252 (N_2252,N_2008,N_2171);
nor U2253 (N_2253,N_2104,N_2071);
and U2254 (N_2254,N_2082,N_2033);
and U2255 (N_2255,N_2134,N_2164);
or U2256 (N_2256,N_2026,N_2027);
and U2257 (N_2257,N_2066,N_2190);
xnor U2258 (N_2258,N_2042,N_2015);
xnor U2259 (N_2259,N_2126,N_2177);
and U2260 (N_2260,N_2086,N_2005);
nor U2261 (N_2261,N_2087,N_2182);
and U2262 (N_2262,N_2124,N_2080);
nand U2263 (N_2263,N_2101,N_2153);
xor U2264 (N_2264,N_2188,N_2016);
or U2265 (N_2265,N_2115,N_2041);
or U2266 (N_2266,N_2079,N_2009);
or U2267 (N_2267,N_2014,N_2001);
nand U2268 (N_2268,N_2049,N_2097);
and U2269 (N_2269,N_2003,N_2076);
nor U2270 (N_2270,N_2111,N_2064);
and U2271 (N_2271,N_2088,N_2173);
nand U2272 (N_2272,N_2117,N_2133);
xnor U2273 (N_2273,N_2020,N_2103);
xor U2274 (N_2274,N_2157,N_2137);
nand U2275 (N_2275,N_2175,N_2154);
xor U2276 (N_2276,N_2151,N_2091);
or U2277 (N_2277,N_2022,N_2170);
or U2278 (N_2278,N_2024,N_2047);
nand U2279 (N_2279,N_2046,N_2094);
and U2280 (N_2280,N_2029,N_2018);
or U2281 (N_2281,N_2197,N_2150);
nand U2282 (N_2282,N_2198,N_2036);
and U2283 (N_2283,N_2129,N_2038);
or U2284 (N_2284,N_2136,N_2179);
nor U2285 (N_2285,N_2199,N_2131);
nand U2286 (N_2286,N_2149,N_2113);
xnor U2287 (N_2287,N_2043,N_2156);
or U2288 (N_2288,N_2112,N_2002);
or U2289 (N_2289,N_2012,N_2158);
nor U2290 (N_2290,N_2142,N_2176);
and U2291 (N_2291,N_2013,N_2048);
nor U2292 (N_2292,N_2062,N_2075);
and U2293 (N_2293,N_2155,N_2184);
and U2294 (N_2294,N_2180,N_2061);
or U2295 (N_2295,N_2007,N_2121);
nand U2296 (N_2296,N_2056,N_2172);
xor U2297 (N_2297,N_2194,N_2162);
nand U2298 (N_2298,N_2072,N_2089);
nand U2299 (N_2299,N_2035,N_2145);
or U2300 (N_2300,N_2071,N_2156);
nor U2301 (N_2301,N_2158,N_2097);
xor U2302 (N_2302,N_2149,N_2129);
and U2303 (N_2303,N_2036,N_2173);
and U2304 (N_2304,N_2101,N_2050);
nor U2305 (N_2305,N_2175,N_2078);
and U2306 (N_2306,N_2167,N_2109);
nor U2307 (N_2307,N_2051,N_2158);
and U2308 (N_2308,N_2197,N_2145);
xor U2309 (N_2309,N_2132,N_2048);
or U2310 (N_2310,N_2188,N_2163);
nor U2311 (N_2311,N_2189,N_2192);
xnor U2312 (N_2312,N_2197,N_2192);
or U2313 (N_2313,N_2125,N_2188);
xnor U2314 (N_2314,N_2192,N_2103);
xor U2315 (N_2315,N_2094,N_2091);
or U2316 (N_2316,N_2065,N_2052);
xor U2317 (N_2317,N_2136,N_2142);
xor U2318 (N_2318,N_2198,N_2197);
nand U2319 (N_2319,N_2078,N_2134);
and U2320 (N_2320,N_2170,N_2162);
or U2321 (N_2321,N_2046,N_2181);
or U2322 (N_2322,N_2011,N_2171);
and U2323 (N_2323,N_2163,N_2121);
or U2324 (N_2324,N_2131,N_2048);
or U2325 (N_2325,N_2165,N_2073);
xnor U2326 (N_2326,N_2072,N_2106);
xor U2327 (N_2327,N_2101,N_2057);
nand U2328 (N_2328,N_2192,N_2090);
xnor U2329 (N_2329,N_2001,N_2032);
nor U2330 (N_2330,N_2117,N_2067);
or U2331 (N_2331,N_2120,N_2187);
nand U2332 (N_2332,N_2183,N_2158);
xor U2333 (N_2333,N_2015,N_2126);
or U2334 (N_2334,N_2128,N_2058);
and U2335 (N_2335,N_2128,N_2051);
nor U2336 (N_2336,N_2176,N_2068);
nor U2337 (N_2337,N_2127,N_2035);
and U2338 (N_2338,N_2003,N_2091);
or U2339 (N_2339,N_2170,N_2002);
xnor U2340 (N_2340,N_2192,N_2066);
or U2341 (N_2341,N_2152,N_2148);
xnor U2342 (N_2342,N_2170,N_2061);
xnor U2343 (N_2343,N_2177,N_2066);
and U2344 (N_2344,N_2171,N_2051);
xor U2345 (N_2345,N_2000,N_2129);
or U2346 (N_2346,N_2126,N_2074);
and U2347 (N_2347,N_2138,N_2009);
or U2348 (N_2348,N_2177,N_2036);
nor U2349 (N_2349,N_2000,N_2029);
and U2350 (N_2350,N_2132,N_2010);
nor U2351 (N_2351,N_2197,N_2039);
and U2352 (N_2352,N_2014,N_2052);
xor U2353 (N_2353,N_2154,N_2146);
xor U2354 (N_2354,N_2120,N_2176);
and U2355 (N_2355,N_2142,N_2099);
xor U2356 (N_2356,N_2193,N_2151);
nand U2357 (N_2357,N_2116,N_2184);
nand U2358 (N_2358,N_2009,N_2042);
and U2359 (N_2359,N_2021,N_2150);
nor U2360 (N_2360,N_2157,N_2163);
and U2361 (N_2361,N_2135,N_2173);
or U2362 (N_2362,N_2163,N_2005);
or U2363 (N_2363,N_2114,N_2028);
xnor U2364 (N_2364,N_2178,N_2002);
nand U2365 (N_2365,N_2189,N_2069);
and U2366 (N_2366,N_2190,N_2111);
nor U2367 (N_2367,N_2182,N_2191);
and U2368 (N_2368,N_2181,N_2151);
or U2369 (N_2369,N_2140,N_2097);
nor U2370 (N_2370,N_2018,N_2174);
nor U2371 (N_2371,N_2031,N_2135);
nor U2372 (N_2372,N_2140,N_2142);
and U2373 (N_2373,N_2044,N_2051);
nor U2374 (N_2374,N_2050,N_2060);
or U2375 (N_2375,N_2089,N_2135);
nand U2376 (N_2376,N_2112,N_2172);
nand U2377 (N_2377,N_2133,N_2127);
nor U2378 (N_2378,N_2070,N_2089);
or U2379 (N_2379,N_2155,N_2121);
and U2380 (N_2380,N_2019,N_2109);
xor U2381 (N_2381,N_2039,N_2143);
xor U2382 (N_2382,N_2021,N_2075);
and U2383 (N_2383,N_2112,N_2050);
nand U2384 (N_2384,N_2078,N_2099);
xor U2385 (N_2385,N_2118,N_2083);
and U2386 (N_2386,N_2005,N_2028);
nand U2387 (N_2387,N_2142,N_2052);
nor U2388 (N_2388,N_2073,N_2187);
nor U2389 (N_2389,N_2035,N_2190);
nand U2390 (N_2390,N_2133,N_2136);
xnor U2391 (N_2391,N_2126,N_2025);
nor U2392 (N_2392,N_2070,N_2046);
or U2393 (N_2393,N_2146,N_2169);
nand U2394 (N_2394,N_2102,N_2139);
nor U2395 (N_2395,N_2093,N_2132);
xor U2396 (N_2396,N_2005,N_2049);
and U2397 (N_2397,N_2125,N_2154);
nand U2398 (N_2398,N_2136,N_2093);
and U2399 (N_2399,N_2008,N_2014);
and U2400 (N_2400,N_2281,N_2203);
nand U2401 (N_2401,N_2246,N_2316);
xnor U2402 (N_2402,N_2223,N_2217);
nand U2403 (N_2403,N_2250,N_2233);
or U2404 (N_2404,N_2371,N_2215);
nor U2405 (N_2405,N_2294,N_2358);
or U2406 (N_2406,N_2380,N_2280);
nand U2407 (N_2407,N_2328,N_2231);
nor U2408 (N_2408,N_2276,N_2266);
or U2409 (N_2409,N_2355,N_2286);
nor U2410 (N_2410,N_2315,N_2390);
xnor U2411 (N_2411,N_2287,N_2319);
xnor U2412 (N_2412,N_2327,N_2339);
and U2413 (N_2413,N_2394,N_2277);
nand U2414 (N_2414,N_2296,N_2384);
and U2415 (N_2415,N_2353,N_2222);
and U2416 (N_2416,N_2317,N_2270);
nor U2417 (N_2417,N_2208,N_2377);
xor U2418 (N_2418,N_2392,N_2200);
or U2419 (N_2419,N_2299,N_2360);
nand U2420 (N_2420,N_2209,N_2366);
or U2421 (N_2421,N_2261,N_2282);
nand U2422 (N_2422,N_2364,N_2235);
xnor U2423 (N_2423,N_2341,N_2201);
and U2424 (N_2424,N_2206,N_2304);
nor U2425 (N_2425,N_2300,N_2307);
xor U2426 (N_2426,N_2376,N_2374);
and U2427 (N_2427,N_2338,N_2228);
nor U2428 (N_2428,N_2290,N_2239);
xor U2429 (N_2429,N_2369,N_2254);
nor U2430 (N_2430,N_2278,N_2202);
and U2431 (N_2431,N_2324,N_2245);
or U2432 (N_2432,N_2237,N_2361);
xor U2433 (N_2433,N_2314,N_2313);
xnor U2434 (N_2434,N_2257,N_2382);
xnor U2435 (N_2435,N_2321,N_2230);
xor U2436 (N_2436,N_2214,N_2252);
xor U2437 (N_2437,N_2344,N_2213);
xnor U2438 (N_2438,N_2308,N_2323);
nor U2439 (N_2439,N_2351,N_2306);
xor U2440 (N_2440,N_2352,N_2204);
and U2441 (N_2441,N_2275,N_2375);
nor U2442 (N_2442,N_2309,N_2258);
nand U2443 (N_2443,N_2342,N_2301);
nor U2444 (N_2444,N_2332,N_2368);
xnor U2445 (N_2445,N_2381,N_2349);
and U2446 (N_2446,N_2350,N_2320);
or U2447 (N_2447,N_2397,N_2329);
and U2448 (N_2448,N_2210,N_2372);
nor U2449 (N_2449,N_2216,N_2391);
xnor U2450 (N_2450,N_2262,N_2291);
or U2451 (N_2451,N_2386,N_2395);
xor U2452 (N_2452,N_2265,N_2220);
xor U2453 (N_2453,N_2205,N_2263);
and U2454 (N_2454,N_2365,N_2370);
nor U2455 (N_2455,N_2343,N_2256);
nor U2456 (N_2456,N_2221,N_2243);
and U2457 (N_2457,N_2336,N_2357);
nand U2458 (N_2458,N_2273,N_2248);
nand U2459 (N_2459,N_2219,N_2312);
xor U2460 (N_2460,N_2292,N_2242);
nand U2461 (N_2461,N_2211,N_2305);
or U2462 (N_2462,N_2387,N_2331);
nor U2463 (N_2463,N_2251,N_2333);
xor U2464 (N_2464,N_2389,N_2247);
xnor U2465 (N_2465,N_2367,N_2269);
nand U2466 (N_2466,N_2227,N_2378);
xnor U2467 (N_2467,N_2383,N_2334);
nor U2468 (N_2468,N_2385,N_2249);
or U2469 (N_2469,N_2373,N_2288);
nor U2470 (N_2470,N_2293,N_2234);
xor U2471 (N_2471,N_2298,N_2302);
nand U2472 (N_2472,N_2264,N_2311);
nand U2473 (N_2473,N_2255,N_2253);
or U2474 (N_2474,N_2303,N_2363);
nand U2475 (N_2475,N_2326,N_2347);
nand U2476 (N_2476,N_2325,N_2346);
and U2477 (N_2477,N_2297,N_2229);
or U2478 (N_2478,N_2348,N_2318);
xnor U2479 (N_2479,N_2285,N_2225);
nand U2480 (N_2480,N_2212,N_2388);
and U2481 (N_2481,N_2268,N_2218);
or U2482 (N_2482,N_2354,N_2335);
and U2483 (N_2483,N_2398,N_2232);
nand U2484 (N_2484,N_2345,N_2272);
or U2485 (N_2485,N_2244,N_2362);
nand U2486 (N_2486,N_2289,N_2284);
nand U2487 (N_2487,N_2340,N_2322);
nand U2488 (N_2488,N_2260,N_2379);
or U2489 (N_2489,N_2356,N_2267);
and U2490 (N_2490,N_2274,N_2279);
nand U2491 (N_2491,N_2241,N_2359);
nand U2492 (N_2492,N_2271,N_2399);
and U2493 (N_2493,N_2337,N_2207);
nor U2494 (N_2494,N_2283,N_2238);
or U2495 (N_2495,N_2259,N_2295);
xnor U2496 (N_2496,N_2224,N_2240);
nand U2497 (N_2497,N_2236,N_2393);
xnor U2498 (N_2498,N_2330,N_2310);
or U2499 (N_2499,N_2226,N_2396);
xnor U2500 (N_2500,N_2332,N_2379);
and U2501 (N_2501,N_2340,N_2298);
nand U2502 (N_2502,N_2295,N_2356);
xnor U2503 (N_2503,N_2284,N_2222);
nor U2504 (N_2504,N_2327,N_2367);
nor U2505 (N_2505,N_2352,N_2393);
nand U2506 (N_2506,N_2302,N_2359);
nor U2507 (N_2507,N_2211,N_2324);
and U2508 (N_2508,N_2286,N_2203);
and U2509 (N_2509,N_2213,N_2238);
nor U2510 (N_2510,N_2306,N_2391);
nand U2511 (N_2511,N_2331,N_2270);
nor U2512 (N_2512,N_2275,N_2277);
nand U2513 (N_2513,N_2380,N_2249);
and U2514 (N_2514,N_2376,N_2346);
nand U2515 (N_2515,N_2268,N_2209);
and U2516 (N_2516,N_2281,N_2383);
and U2517 (N_2517,N_2315,N_2231);
or U2518 (N_2518,N_2251,N_2296);
nor U2519 (N_2519,N_2339,N_2237);
xnor U2520 (N_2520,N_2311,N_2284);
and U2521 (N_2521,N_2290,N_2302);
nor U2522 (N_2522,N_2316,N_2249);
xnor U2523 (N_2523,N_2237,N_2281);
xor U2524 (N_2524,N_2267,N_2284);
xnor U2525 (N_2525,N_2309,N_2361);
nor U2526 (N_2526,N_2382,N_2225);
nand U2527 (N_2527,N_2370,N_2254);
or U2528 (N_2528,N_2229,N_2247);
nor U2529 (N_2529,N_2309,N_2359);
nand U2530 (N_2530,N_2259,N_2262);
xor U2531 (N_2531,N_2268,N_2204);
xnor U2532 (N_2532,N_2291,N_2259);
nor U2533 (N_2533,N_2229,N_2232);
nor U2534 (N_2534,N_2286,N_2388);
nand U2535 (N_2535,N_2215,N_2254);
and U2536 (N_2536,N_2298,N_2228);
or U2537 (N_2537,N_2295,N_2202);
or U2538 (N_2538,N_2340,N_2385);
nand U2539 (N_2539,N_2314,N_2349);
and U2540 (N_2540,N_2229,N_2361);
and U2541 (N_2541,N_2379,N_2210);
or U2542 (N_2542,N_2369,N_2392);
or U2543 (N_2543,N_2238,N_2354);
and U2544 (N_2544,N_2224,N_2387);
and U2545 (N_2545,N_2223,N_2205);
nand U2546 (N_2546,N_2339,N_2379);
nand U2547 (N_2547,N_2320,N_2270);
xnor U2548 (N_2548,N_2347,N_2233);
and U2549 (N_2549,N_2311,N_2273);
xor U2550 (N_2550,N_2387,N_2379);
or U2551 (N_2551,N_2272,N_2238);
or U2552 (N_2552,N_2385,N_2279);
or U2553 (N_2553,N_2247,N_2298);
nand U2554 (N_2554,N_2286,N_2297);
nor U2555 (N_2555,N_2228,N_2272);
nand U2556 (N_2556,N_2378,N_2203);
nor U2557 (N_2557,N_2382,N_2343);
or U2558 (N_2558,N_2288,N_2340);
nand U2559 (N_2559,N_2204,N_2209);
nand U2560 (N_2560,N_2365,N_2368);
or U2561 (N_2561,N_2248,N_2235);
and U2562 (N_2562,N_2399,N_2303);
nor U2563 (N_2563,N_2297,N_2324);
or U2564 (N_2564,N_2238,N_2362);
nor U2565 (N_2565,N_2270,N_2377);
and U2566 (N_2566,N_2347,N_2319);
nand U2567 (N_2567,N_2218,N_2302);
or U2568 (N_2568,N_2341,N_2324);
xnor U2569 (N_2569,N_2218,N_2390);
or U2570 (N_2570,N_2293,N_2254);
and U2571 (N_2571,N_2221,N_2352);
xor U2572 (N_2572,N_2348,N_2234);
and U2573 (N_2573,N_2304,N_2382);
nor U2574 (N_2574,N_2210,N_2217);
and U2575 (N_2575,N_2271,N_2305);
or U2576 (N_2576,N_2310,N_2341);
xnor U2577 (N_2577,N_2263,N_2387);
xnor U2578 (N_2578,N_2211,N_2250);
xnor U2579 (N_2579,N_2390,N_2295);
nand U2580 (N_2580,N_2295,N_2367);
xnor U2581 (N_2581,N_2399,N_2317);
nand U2582 (N_2582,N_2224,N_2399);
and U2583 (N_2583,N_2217,N_2364);
nand U2584 (N_2584,N_2288,N_2250);
xor U2585 (N_2585,N_2347,N_2320);
and U2586 (N_2586,N_2369,N_2312);
xnor U2587 (N_2587,N_2280,N_2270);
xnor U2588 (N_2588,N_2244,N_2398);
xor U2589 (N_2589,N_2361,N_2397);
nand U2590 (N_2590,N_2320,N_2395);
or U2591 (N_2591,N_2222,N_2215);
or U2592 (N_2592,N_2293,N_2306);
xor U2593 (N_2593,N_2291,N_2329);
xnor U2594 (N_2594,N_2343,N_2372);
xor U2595 (N_2595,N_2323,N_2389);
nand U2596 (N_2596,N_2395,N_2335);
and U2597 (N_2597,N_2398,N_2309);
nor U2598 (N_2598,N_2267,N_2379);
xnor U2599 (N_2599,N_2284,N_2361);
or U2600 (N_2600,N_2407,N_2414);
and U2601 (N_2601,N_2455,N_2532);
and U2602 (N_2602,N_2551,N_2528);
or U2603 (N_2603,N_2484,N_2411);
nor U2604 (N_2604,N_2596,N_2480);
nor U2605 (N_2605,N_2542,N_2423);
xor U2606 (N_2606,N_2545,N_2451);
nand U2607 (N_2607,N_2440,N_2519);
nand U2608 (N_2608,N_2550,N_2594);
nor U2609 (N_2609,N_2406,N_2487);
xnor U2610 (N_2610,N_2462,N_2522);
xor U2611 (N_2611,N_2489,N_2497);
xnor U2612 (N_2612,N_2500,N_2570);
nand U2613 (N_2613,N_2453,N_2482);
nor U2614 (N_2614,N_2585,N_2424);
xnor U2615 (N_2615,N_2485,N_2595);
or U2616 (N_2616,N_2456,N_2588);
xnor U2617 (N_2617,N_2464,N_2427);
xnor U2618 (N_2618,N_2574,N_2428);
xnor U2619 (N_2619,N_2520,N_2573);
nand U2620 (N_2620,N_2513,N_2576);
nor U2621 (N_2621,N_2527,N_2465);
and U2622 (N_2622,N_2511,N_2418);
or U2623 (N_2623,N_2472,N_2599);
nor U2624 (N_2624,N_2442,N_2447);
nor U2625 (N_2625,N_2559,N_2557);
xnor U2626 (N_2626,N_2530,N_2494);
and U2627 (N_2627,N_2581,N_2476);
nand U2628 (N_2628,N_2473,N_2549);
and U2629 (N_2629,N_2562,N_2499);
nor U2630 (N_2630,N_2420,N_2400);
or U2631 (N_2631,N_2431,N_2401);
xor U2632 (N_2632,N_2516,N_2533);
and U2633 (N_2633,N_2521,N_2583);
nor U2634 (N_2634,N_2531,N_2556);
xor U2635 (N_2635,N_2564,N_2432);
and U2636 (N_2636,N_2569,N_2470);
xor U2637 (N_2637,N_2589,N_2537);
and U2638 (N_2638,N_2460,N_2415);
or U2639 (N_2639,N_2449,N_2430);
nand U2640 (N_2640,N_2512,N_2477);
or U2641 (N_2641,N_2468,N_2547);
or U2642 (N_2642,N_2571,N_2553);
nor U2643 (N_2643,N_2446,N_2546);
and U2644 (N_2644,N_2538,N_2509);
nor U2645 (N_2645,N_2548,N_2412);
and U2646 (N_2646,N_2541,N_2567);
nand U2647 (N_2647,N_2426,N_2558);
nor U2648 (N_2648,N_2490,N_2591);
or U2649 (N_2649,N_2598,N_2421);
xor U2650 (N_2650,N_2526,N_2529);
nand U2651 (N_2651,N_2404,N_2444);
or U2652 (N_2652,N_2555,N_2517);
xnor U2653 (N_2653,N_2560,N_2425);
nor U2654 (N_2654,N_2552,N_2579);
nand U2655 (N_2655,N_2506,N_2413);
xor U2656 (N_2656,N_2498,N_2448);
xnor U2657 (N_2657,N_2445,N_2496);
nand U2658 (N_2658,N_2503,N_2405);
and U2659 (N_2659,N_2514,N_2403);
or U2660 (N_2660,N_2469,N_2419);
nor U2661 (N_2661,N_2486,N_2593);
nand U2662 (N_2662,N_2481,N_2474);
or U2663 (N_2663,N_2438,N_2586);
nand U2664 (N_2664,N_2536,N_2441);
xnor U2665 (N_2665,N_2454,N_2572);
nand U2666 (N_2666,N_2433,N_2587);
nor U2667 (N_2667,N_2535,N_2483);
nor U2668 (N_2668,N_2510,N_2458);
nand U2669 (N_2669,N_2478,N_2515);
or U2670 (N_2670,N_2452,N_2410);
and U2671 (N_2671,N_2543,N_2439);
nand U2672 (N_2672,N_2457,N_2568);
xor U2673 (N_2673,N_2492,N_2577);
nor U2674 (N_2674,N_2554,N_2539);
nand U2675 (N_2675,N_2408,N_2409);
and U2676 (N_2676,N_2580,N_2436);
and U2677 (N_2677,N_2566,N_2563);
and U2678 (N_2678,N_2402,N_2450);
and U2679 (N_2679,N_2504,N_2467);
nand U2680 (N_2680,N_2479,N_2501);
xnor U2681 (N_2681,N_2435,N_2561);
and U2682 (N_2682,N_2459,N_2544);
nand U2683 (N_2683,N_2488,N_2523);
nand U2684 (N_2684,N_2422,N_2493);
nand U2685 (N_2685,N_2417,N_2524);
or U2686 (N_2686,N_2584,N_2592);
nand U2687 (N_2687,N_2495,N_2590);
nand U2688 (N_2688,N_2475,N_2534);
and U2689 (N_2689,N_2463,N_2491);
or U2690 (N_2690,N_2525,N_2505);
or U2691 (N_2691,N_2578,N_2471);
nand U2692 (N_2692,N_2461,N_2540);
nor U2693 (N_2693,N_2416,N_2597);
or U2694 (N_2694,N_2565,N_2466);
and U2695 (N_2695,N_2437,N_2507);
nor U2696 (N_2696,N_2508,N_2502);
or U2697 (N_2697,N_2429,N_2518);
or U2698 (N_2698,N_2443,N_2434);
and U2699 (N_2699,N_2575,N_2582);
nor U2700 (N_2700,N_2507,N_2478);
nand U2701 (N_2701,N_2484,N_2572);
and U2702 (N_2702,N_2418,N_2460);
and U2703 (N_2703,N_2527,N_2499);
nor U2704 (N_2704,N_2462,N_2537);
nor U2705 (N_2705,N_2525,N_2450);
nor U2706 (N_2706,N_2416,N_2426);
nand U2707 (N_2707,N_2554,N_2525);
and U2708 (N_2708,N_2545,N_2548);
nand U2709 (N_2709,N_2567,N_2464);
nand U2710 (N_2710,N_2587,N_2428);
nor U2711 (N_2711,N_2534,N_2547);
nand U2712 (N_2712,N_2479,N_2458);
nor U2713 (N_2713,N_2447,N_2587);
and U2714 (N_2714,N_2471,N_2511);
nand U2715 (N_2715,N_2467,N_2545);
or U2716 (N_2716,N_2559,N_2469);
nand U2717 (N_2717,N_2528,N_2426);
nor U2718 (N_2718,N_2586,N_2598);
and U2719 (N_2719,N_2595,N_2467);
nand U2720 (N_2720,N_2498,N_2591);
xor U2721 (N_2721,N_2417,N_2493);
nor U2722 (N_2722,N_2504,N_2440);
nor U2723 (N_2723,N_2580,N_2575);
nor U2724 (N_2724,N_2462,N_2499);
nand U2725 (N_2725,N_2556,N_2564);
xnor U2726 (N_2726,N_2584,N_2596);
or U2727 (N_2727,N_2464,N_2446);
or U2728 (N_2728,N_2582,N_2512);
nor U2729 (N_2729,N_2461,N_2488);
nor U2730 (N_2730,N_2513,N_2452);
nand U2731 (N_2731,N_2530,N_2495);
nor U2732 (N_2732,N_2589,N_2533);
xor U2733 (N_2733,N_2561,N_2492);
nand U2734 (N_2734,N_2454,N_2544);
xnor U2735 (N_2735,N_2547,N_2594);
nor U2736 (N_2736,N_2476,N_2497);
nor U2737 (N_2737,N_2545,N_2537);
nor U2738 (N_2738,N_2522,N_2597);
nand U2739 (N_2739,N_2544,N_2507);
nand U2740 (N_2740,N_2591,N_2508);
xor U2741 (N_2741,N_2465,N_2562);
and U2742 (N_2742,N_2583,N_2529);
nor U2743 (N_2743,N_2471,N_2559);
xor U2744 (N_2744,N_2477,N_2484);
or U2745 (N_2745,N_2416,N_2439);
nand U2746 (N_2746,N_2579,N_2508);
nor U2747 (N_2747,N_2516,N_2452);
and U2748 (N_2748,N_2450,N_2570);
and U2749 (N_2749,N_2497,N_2501);
nand U2750 (N_2750,N_2579,N_2471);
nor U2751 (N_2751,N_2503,N_2423);
xnor U2752 (N_2752,N_2414,N_2486);
and U2753 (N_2753,N_2534,N_2464);
nand U2754 (N_2754,N_2509,N_2573);
and U2755 (N_2755,N_2542,N_2580);
xnor U2756 (N_2756,N_2488,N_2566);
xor U2757 (N_2757,N_2440,N_2517);
nor U2758 (N_2758,N_2429,N_2452);
or U2759 (N_2759,N_2488,N_2546);
or U2760 (N_2760,N_2491,N_2579);
and U2761 (N_2761,N_2557,N_2446);
and U2762 (N_2762,N_2452,N_2526);
nand U2763 (N_2763,N_2404,N_2464);
nor U2764 (N_2764,N_2469,N_2431);
and U2765 (N_2765,N_2556,N_2501);
nor U2766 (N_2766,N_2528,N_2576);
nor U2767 (N_2767,N_2495,N_2429);
and U2768 (N_2768,N_2449,N_2477);
xor U2769 (N_2769,N_2533,N_2401);
nand U2770 (N_2770,N_2581,N_2538);
and U2771 (N_2771,N_2591,N_2579);
nand U2772 (N_2772,N_2481,N_2558);
nand U2773 (N_2773,N_2407,N_2549);
or U2774 (N_2774,N_2517,N_2464);
and U2775 (N_2775,N_2468,N_2513);
and U2776 (N_2776,N_2563,N_2591);
nor U2777 (N_2777,N_2535,N_2401);
xor U2778 (N_2778,N_2434,N_2446);
and U2779 (N_2779,N_2529,N_2491);
xor U2780 (N_2780,N_2592,N_2511);
nor U2781 (N_2781,N_2527,N_2537);
nor U2782 (N_2782,N_2545,N_2424);
xor U2783 (N_2783,N_2403,N_2490);
nor U2784 (N_2784,N_2587,N_2482);
and U2785 (N_2785,N_2553,N_2408);
nand U2786 (N_2786,N_2446,N_2477);
and U2787 (N_2787,N_2513,N_2589);
nand U2788 (N_2788,N_2527,N_2463);
and U2789 (N_2789,N_2456,N_2436);
xnor U2790 (N_2790,N_2475,N_2457);
nand U2791 (N_2791,N_2513,N_2594);
nand U2792 (N_2792,N_2570,N_2432);
and U2793 (N_2793,N_2545,N_2436);
and U2794 (N_2794,N_2583,N_2472);
or U2795 (N_2795,N_2593,N_2434);
or U2796 (N_2796,N_2558,N_2401);
or U2797 (N_2797,N_2567,N_2423);
and U2798 (N_2798,N_2446,N_2528);
nand U2799 (N_2799,N_2470,N_2465);
xnor U2800 (N_2800,N_2617,N_2737);
nor U2801 (N_2801,N_2791,N_2687);
xnor U2802 (N_2802,N_2764,N_2674);
and U2803 (N_2803,N_2732,N_2779);
or U2804 (N_2804,N_2606,N_2718);
or U2805 (N_2805,N_2782,N_2781);
and U2806 (N_2806,N_2641,N_2616);
nand U2807 (N_2807,N_2780,N_2642);
and U2808 (N_2808,N_2766,N_2620);
or U2809 (N_2809,N_2660,N_2638);
nor U2810 (N_2810,N_2646,N_2786);
xnor U2811 (N_2811,N_2662,N_2688);
or U2812 (N_2812,N_2767,N_2651);
nand U2813 (N_2813,N_2715,N_2668);
nand U2814 (N_2814,N_2736,N_2719);
nand U2815 (N_2815,N_2725,N_2701);
or U2816 (N_2816,N_2756,N_2792);
or U2817 (N_2817,N_2644,N_2773);
or U2818 (N_2818,N_2771,N_2699);
xor U2819 (N_2819,N_2640,N_2671);
nand U2820 (N_2820,N_2664,N_2613);
and U2821 (N_2821,N_2768,N_2735);
nor U2822 (N_2822,N_2635,N_2793);
nand U2823 (N_2823,N_2637,N_2716);
xor U2824 (N_2824,N_2627,N_2709);
and U2825 (N_2825,N_2626,N_2794);
xnor U2826 (N_2826,N_2631,N_2708);
nand U2827 (N_2827,N_2698,N_2747);
and U2828 (N_2828,N_2785,N_2745);
and U2829 (N_2829,N_2624,N_2649);
or U2830 (N_2830,N_2653,N_2705);
xor U2831 (N_2831,N_2661,N_2691);
or U2832 (N_2832,N_2695,N_2740);
xnor U2833 (N_2833,N_2618,N_2743);
nor U2834 (N_2834,N_2645,N_2729);
nor U2835 (N_2835,N_2765,N_2752);
nand U2836 (N_2836,N_2778,N_2721);
or U2837 (N_2837,N_2774,N_2741);
xor U2838 (N_2838,N_2723,N_2656);
nand U2839 (N_2839,N_2733,N_2692);
or U2840 (N_2840,N_2703,N_2672);
or U2841 (N_2841,N_2726,N_2652);
nor U2842 (N_2842,N_2681,N_2684);
nor U2843 (N_2843,N_2742,N_2760);
xnor U2844 (N_2844,N_2798,N_2679);
or U2845 (N_2845,N_2738,N_2647);
nor U2846 (N_2846,N_2685,N_2763);
and U2847 (N_2847,N_2704,N_2728);
or U2848 (N_2848,N_2609,N_2682);
nor U2849 (N_2849,N_2675,N_2625);
and U2850 (N_2850,N_2734,N_2673);
nor U2851 (N_2851,N_2724,N_2677);
xor U2852 (N_2852,N_2607,N_2796);
xor U2853 (N_2853,N_2711,N_2602);
or U2854 (N_2854,N_2623,N_2659);
nor U2855 (N_2855,N_2758,N_2690);
xnor U2856 (N_2856,N_2759,N_2762);
and U2857 (N_2857,N_2789,N_2730);
or U2858 (N_2858,N_2600,N_2648);
and U2859 (N_2859,N_2717,N_2658);
and U2860 (N_2860,N_2761,N_2731);
nand U2861 (N_2861,N_2754,N_2670);
xor U2862 (N_2862,N_2669,N_2694);
or U2863 (N_2863,N_2707,N_2621);
and U2864 (N_2864,N_2689,N_2755);
and U2865 (N_2865,N_2615,N_2632);
nor U2866 (N_2866,N_2628,N_2784);
or U2867 (N_2867,N_2693,N_2601);
or U2868 (N_2868,N_2770,N_2788);
and U2869 (N_2869,N_2706,N_2797);
xnor U2870 (N_2870,N_2619,N_2769);
nor U2871 (N_2871,N_2787,N_2722);
xor U2872 (N_2872,N_2795,N_2714);
and U2873 (N_2873,N_2614,N_2700);
nor U2874 (N_2874,N_2712,N_2612);
xnor U2875 (N_2875,N_2739,N_2633);
nor U2876 (N_2876,N_2697,N_2680);
and U2877 (N_2877,N_2799,N_2750);
or U2878 (N_2878,N_2643,N_2744);
or U2879 (N_2879,N_2654,N_2683);
and U2880 (N_2880,N_2678,N_2753);
or U2881 (N_2881,N_2696,N_2751);
or U2882 (N_2882,N_2710,N_2790);
and U2883 (N_2883,N_2757,N_2629);
or U2884 (N_2884,N_2655,N_2639);
or U2885 (N_2885,N_2727,N_2604);
nand U2886 (N_2886,N_2746,N_2657);
xnor U2887 (N_2887,N_2666,N_2776);
nor U2888 (N_2888,N_2720,N_2686);
nor U2889 (N_2889,N_2611,N_2777);
nand U2890 (N_2890,N_2610,N_2713);
nand U2891 (N_2891,N_2702,N_2605);
nor U2892 (N_2892,N_2603,N_2676);
or U2893 (N_2893,N_2783,N_2772);
xor U2894 (N_2894,N_2749,N_2634);
nor U2895 (N_2895,N_2667,N_2622);
or U2896 (N_2896,N_2608,N_2663);
nand U2897 (N_2897,N_2636,N_2748);
nand U2898 (N_2898,N_2775,N_2630);
nand U2899 (N_2899,N_2665,N_2650);
or U2900 (N_2900,N_2756,N_2631);
and U2901 (N_2901,N_2673,N_2755);
or U2902 (N_2902,N_2761,N_2790);
xnor U2903 (N_2903,N_2650,N_2711);
and U2904 (N_2904,N_2715,N_2759);
and U2905 (N_2905,N_2635,N_2692);
nand U2906 (N_2906,N_2687,N_2741);
nand U2907 (N_2907,N_2753,N_2751);
xor U2908 (N_2908,N_2741,N_2724);
nand U2909 (N_2909,N_2755,N_2697);
or U2910 (N_2910,N_2636,N_2752);
nand U2911 (N_2911,N_2600,N_2791);
xnor U2912 (N_2912,N_2714,N_2685);
xnor U2913 (N_2913,N_2661,N_2628);
and U2914 (N_2914,N_2633,N_2745);
xor U2915 (N_2915,N_2723,N_2778);
and U2916 (N_2916,N_2683,N_2704);
nand U2917 (N_2917,N_2731,N_2708);
nor U2918 (N_2918,N_2613,N_2669);
or U2919 (N_2919,N_2761,N_2717);
and U2920 (N_2920,N_2662,N_2622);
nand U2921 (N_2921,N_2671,N_2735);
or U2922 (N_2922,N_2645,N_2617);
and U2923 (N_2923,N_2630,N_2731);
or U2924 (N_2924,N_2649,N_2777);
and U2925 (N_2925,N_2633,N_2642);
or U2926 (N_2926,N_2618,N_2789);
nor U2927 (N_2927,N_2626,N_2738);
nand U2928 (N_2928,N_2610,N_2716);
nor U2929 (N_2929,N_2601,N_2795);
nor U2930 (N_2930,N_2795,N_2687);
and U2931 (N_2931,N_2785,N_2698);
nor U2932 (N_2932,N_2608,N_2671);
or U2933 (N_2933,N_2716,N_2643);
nand U2934 (N_2934,N_2633,N_2681);
nand U2935 (N_2935,N_2732,N_2676);
xor U2936 (N_2936,N_2671,N_2600);
nand U2937 (N_2937,N_2612,N_2637);
nor U2938 (N_2938,N_2742,N_2779);
xor U2939 (N_2939,N_2671,N_2771);
xnor U2940 (N_2940,N_2608,N_2699);
xnor U2941 (N_2941,N_2624,N_2703);
and U2942 (N_2942,N_2771,N_2719);
nor U2943 (N_2943,N_2704,N_2652);
or U2944 (N_2944,N_2711,N_2702);
xnor U2945 (N_2945,N_2786,N_2672);
nor U2946 (N_2946,N_2784,N_2615);
nor U2947 (N_2947,N_2740,N_2775);
xnor U2948 (N_2948,N_2679,N_2673);
nor U2949 (N_2949,N_2753,N_2666);
and U2950 (N_2950,N_2761,N_2626);
nand U2951 (N_2951,N_2619,N_2668);
nor U2952 (N_2952,N_2730,N_2764);
or U2953 (N_2953,N_2618,N_2776);
xnor U2954 (N_2954,N_2709,N_2741);
and U2955 (N_2955,N_2660,N_2615);
or U2956 (N_2956,N_2763,N_2603);
nor U2957 (N_2957,N_2769,N_2651);
xor U2958 (N_2958,N_2641,N_2612);
or U2959 (N_2959,N_2671,N_2795);
and U2960 (N_2960,N_2722,N_2737);
or U2961 (N_2961,N_2639,N_2712);
or U2962 (N_2962,N_2731,N_2684);
and U2963 (N_2963,N_2644,N_2767);
nor U2964 (N_2964,N_2664,N_2681);
and U2965 (N_2965,N_2682,N_2620);
and U2966 (N_2966,N_2726,N_2693);
and U2967 (N_2967,N_2764,N_2738);
nand U2968 (N_2968,N_2756,N_2667);
nor U2969 (N_2969,N_2677,N_2604);
nor U2970 (N_2970,N_2693,N_2621);
and U2971 (N_2971,N_2670,N_2741);
or U2972 (N_2972,N_2614,N_2663);
xnor U2973 (N_2973,N_2726,N_2783);
xor U2974 (N_2974,N_2643,N_2763);
xor U2975 (N_2975,N_2652,N_2709);
xor U2976 (N_2976,N_2737,N_2694);
and U2977 (N_2977,N_2629,N_2651);
nand U2978 (N_2978,N_2658,N_2679);
xor U2979 (N_2979,N_2771,N_2797);
xor U2980 (N_2980,N_2675,N_2689);
nand U2981 (N_2981,N_2619,N_2788);
nand U2982 (N_2982,N_2794,N_2607);
nand U2983 (N_2983,N_2671,N_2624);
xnor U2984 (N_2984,N_2777,N_2609);
nor U2985 (N_2985,N_2772,N_2621);
nor U2986 (N_2986,N_2752,N_2601);
nor U2987 (N_2987,N_2631,N_2635);
nand U2988 (N_2988,N_2619,N_2779);
nor U2989 (N_2989,N_2648,N_2740);
or U2990 (N_2990,N_2728,N_2692);
xnor U2991 (N_2991,N_2661,N_2655);
xnor U2992 (N_2992,N_2623,N_2690);
xor U2993 (N_2993,N_2682,N_2686);
nand U2994 (N_2994,N_2660,N_2619);
xnor U2995 (N_2995,N_2713,N_2677);
xnor U2996 (N_2996,N_2664,N_2666);
and U2997 (N_2997,N_2605,N_2748);
or U2998 (N_2998,N_2765,N_2769);
nor U2999 (N_2999,N_2756,N_2668);
nand U3000 (N_3000,N_2920,N_2820);
nor U3001 (N_3001,N_2833,N_2861);
nand U3002 (N_3002,N_2911,N_2814);
nor U3003 (N_3003,N_2853,N_2808);
or U3004 (N_3004,N_2866,N_2869);
xnor U3005 (N_3005,N_2857,N_2870);
nand U3006 (N_3006,N_2899,N_2862);
nor U3007 (N_3007,N_2888,N_2977);
nand U3008 (N_3008,N_2889,N_2971);
xnor U3009 (N_3009,N_2882,N_2886);
and U3010 (N_3010,N_2878,N_2944);
and U3011 (N_3011,N_2828,N_2923);
xor U3012 (N_3012,N_2938,N_2915);
and U3013 (N_3013,N_2917,N_2969);
nor U3014 (N_3014,N_2956,N_2932);
and U3015 (N_3015,N_2848,N_2876);
nand U3016 (N_3016,N_2895,N_2945);
and U3017 (N_3017,N_2877,N_2805);
and U3018 (N_3018,N_2991,N_2872);
or U3019 (N_3019,N_2906,N_2830);
nor U3020 (N_3020,N_2841,N_2806);
xnor U3021 (N_3021,N_2874,N_2840);
nor U3022 (N_3022,N_2968,N_2901);
and U3023 (N_3023,N_2890,N_2897);
and U3024 (N_3024,N_2912,N_2910);
or U3025 (N_3025,N_2918,N_2999);
nor U3026 (N_3026,N_2967,N_2865);
or U3027 (N_3027,N_2824,N_2936);
nor U3028 (N_3028,N_2942,N_2834);
nand U3029 (N_3029,N_2998,N_2827);
and U3030 (N_3030,N_2950,N_2948);
nor U3031 (N_3031,N_2851,N_2823);
nor U3032 (N_3032,N_2815,N_2850);
nor U3033 (N_3033,N_2957,N_2859);
and U3034 (N_3034,N_2990,N_2963);
or U3035 (N_3035,N_2843,N_2913);
nor U3036 (N_3036,N_2852,N_2896);
nand U3037 (N_3037,N_2994,N_2856);
nor U3038 (N_3038,N_2826,N_2854);
nand U3039 (N_3039,N_2930,N_2993);
xnor U3040 (N_3040,N_2953,N_2844);
xnor U3041 (N_3041,N_2959,N_2952);
and U3042 (N_3042,N_2831,N_2846);
or U3043 (N_3043,N_2811,N_2928);
or U3044 (N_3044,N_2845,N_2997);
or U3045 (N_3045,N_2821,N_2892);
xor U3046 (N_3046,N_2960,N_2801);
xor U3047 (N_3047,N_2898,N_2875);
or U3048 (N_3048,N_2987,N_2809);
nand U3049 (N_3049,N_2972,N_2829);
and U3050 (N_3050,N_2868,N_2939);
or U3051 (N_3051,N_2907,N_2937);
or U3052 (N_3052,N_2849,N_2817);
nor U3053 (N_3053,N_2836,N_2926);
and U3054 (N_3054,N_2954,N_2961);
xnor U3055 (N_3055,N_2943,N_2985);
xor U3056 (N_3056,N_2976,N_2946);
nor U3057 (N_3057,N_2981,N_2973);
nand U3058 (N_3058,N_2904,N_2916);
nand U3059 (N_3059,N_2884,N_2842);
nor U3060 (N_3060,N_2992,N_2964);
or U3061 (N_3061,N_2982,N_2940);
nand U3062 (N_3062,N_2858,N_2934);
xor U3063 (N_3063,N_2812,N_2995);
nand U3064 (N_3064,N_2965,N_2908);
xor U3065 (N_3065,N_2947,N_2933);
xnor U3066 (N_3066,N_2909,N_2838);
nor U3067 (N_3067,N_2983,N_2979);
and U3068 (N_3068,N_2873,N_2921);
or U3069 (N_3069,N_2879,N_2860);
nor U3070 (N_3070,N_2837,N_2804);
and U3071 (N_3071,N_2864,N_2881);
nor U3072 (N_3072,N_2941,N_2986);
nand U3073 (N_3073,N_2871,N_2810);
nor U3074 (N_3074,N_2887,N_2825);
nand U3075 (N_3075,N_2978,N_2914);
or U3076 (N_3076,N_2818,N_2835);
xor U3077 (N_3077,N_2925,N_2816);
nand U3078 (N_3078,N_2894,N_2927);
or U3079 (N_3079,N_2891,N_2931);
xnor U3080 (N_3080,N_2974,N_2919);
and U3081 (N_3081,N_2807,N_2955);
and U3082 (N_3082,N_2867,N_2832);
nand U3083 (N_3083,N_2819,N_2970);
nand U3084 (N_3084,N_2893,N_2822);
or U3085 (N_3085,N_2975,N_2996);
nand U3086 (N_3086,N_2855,N_2839);
nand U3087 (N_3087,N_2924,N_2813);
xor U3088 (N_3088,N_2929,N_2988);
nor U3089 (N_3089,N_2958,N_2951);
and U3090 (N_3090,N_2863,N_2900);
or U3091 (N_3091,N_2800,N_2949);
nand U3092 (N_3092,N_2966,N_2802);
or U3093 (N_3093,N_2989,N_2984);
nand U3094 (N_3094,N_2883,N_2962);
xnor U3095 (N_3095,N_2903,N_2905);
or U3096 (N_3096,N_2885,N_2847);
nand U3097 (N_3097,N_2922,N_2803);
xor U3098 (N_3098,N_2880,N_2902);
nor U3099 (N_3099,N_2980,N_2935);
xnor U3100 (N_3100,N_2835,N_2918);
and U3101 (N_3101,N_2946,N_2877);
and U3102 (N_3102,N_2950,N_2804);
xnor U3103 (N_3103,N_2869,N_2947);
xnor U3104 (N_3104,N_2887,N_2901);
nand U3105 (N_3105,N_2836,N_2904);
xnor U3106 (N_3106,N_2875,N_2894);
nand U3107 (N_3107,N_2993,N_2951);
and U3108 (N_3108,N_2933,N_2816);
xnor U3109 (N_3109,N_2955,N_2856);
xnor U3110 (N_3110,N_2897,N_2881);
or U3111 (N_3111,N_2803,N_2911);
xnor U3112 (N_3112,N_2905,N_2968);
nand U3113 (N_3113,N_2894,N_2985);
xnor U3114 (N_3114,N_2901,N_2885);
or U3115 (N_3115,N_2801,N_2993);
nor U3116 (N_3116,N_2984,N_2981);
nor U3117 (N_3117,N_2966,N_2801);
nor U3118 (N_3118,N_2981,N_2905);
nor U3119 (N_3119,N_2885,N_2844);
nand U3120 (N_3120,N_2921,N_2959);
and U3121 (N_3121,N_2913,N_2962);
or U3122 (N_3122,N_2800,N_2816);
or U3123 (N_3123,N_2930,N_2803);
and U3124 (N_3124,N_2810,N_2854);
or U3125 (N_3125,N_2884,N_2825);
or U3126 (N_3126,N_2965,N_2856);
xnor U3127 (N_3127,N_2821,N_2914);
nor U3128 (N_3128,N_2948,N_2828);
nand U3129 (N_3129,N_2882,N_2896);
xnor U3130 (N_3130,N_2928,N_2838);
or U3131 (N_3131,N_2800,N_2879);
or U3132 (N_3132,N_2954,N_2963);
nor U3133 (N_3133,N_2946,N_2866);
and U3134 (N_3134,N_2900,N_2818);
and U3135 (N_3135,N_2947,N_2969);
nand U3136 (N_3136,N_2911,N_2979);
and U3137 (N_3137,N_2963,N_2983);
or U3138 (N_3138,N_2896,N_2961);
and U3139 (N_3139,N_2873,N_2972);
nand U3140 (N_3140,N_2952,N_2948);
or U3141 (N_3141,N_2806,N_2811);
nand U3142 (N_3142,N_2894,N_2907);
xor U3143 (N_3143,N_2860,N_2949);
nor U3144 (N_3144,N_2904,N_2882);
nand U3145 (N_3145,N_2985,N_2846);
or U3146 (N_3146,N_2822,N_2868);
xor U3147 (N_3147,N_2830,N_2964);
or U3148 (N_3148,N_2824,N_2926);
nand U3149 (N_3149,N_2841,N_2911);
nor U3150 (N_3150,N_2955,N_2878);
and U3151 (N_3151,N_2821,N_2804);
xnor U3152 (N_3152,N_2877,N_2942);
or U3153 (N_3153,N_2800,N_2922);
xor U3154 (N_3154,N_2802,N_2972);
nand U3155 (N_3155,N_2961,N_2977);
nor U3156 (N_3156,N_2879,N_2912);
and U3157 (N_3157,N_2912,N_2962);
nand U3158 (N_3158,N_2930,N_2914);
nand U3159 (N_3159,N_2866,N_2803);
nor U3160 (N_3160,N_2856,N_2951);
nand U3161 (N_3161,N_2940,N_2926);
nand U3162 (N_3162,N_2803,N_2906);
xor U3163 (N_3163,N_2952,N_2939);
or U3164 (N_3164,N_2947,N_2887);
nand U3165 (N_3165,N_2946,N_2861);
or U3166 (N_3166,N_2914,N_2912);
xor U3167 (N_3167,N_2986,N_2939);
nand U3168 (N_3168,N_2991,N_2801);
and U3169 (N_3169,N_2939,N_2931);
and U3170 (N_3170,N_2917,N_2864);
nand U3171 (N_3171,N_2801,N_2900);
or U3172 (N_3172,N_2871,N_2999);
and U3173 (N_3173,N_2955,N_2949);
nor U3174 (N_3174,N_2894,N_2853);
nand U3175 (N_3175,N_2923,N_2884);
nand U3176 (N_3176,N_2975,N_2947);
nand U3177 (N_3177,N_2836,N_2980);
nand U3178 (N_3178,N_2856,N_2804);
or U3179 (N_3179,N_2938,N_2900);
nor U3180 (N_3180,N_2810,N_2940);
or U3181 (N_3181,N_2833,N_2929);
or U3182 (N_3182,N_2843,N_2949);
xnor U3183 (N_3183,N_2903,N_2816);
xor U3184 (N_3184,N_2941,N_2801);
and U3185 (N_3185,N_2908,N_2956);
or U3186 (N_3186,N_2834,N_2816);
or U3187 (N_3187,N_2801,N_2819);
nor U3188 (N_3188,N_2936,N_2981);
and U3189 (N_3189,N_2967,N_2942);
nor U3190 (N_3190,N_2894,N_2850);
nand U3191 (N_3191,N_2973,N_2993);
or U3192 (N_3192,N_2824,N_2922);
xor U3193 (N_3193,N_2837,N_2960);
nor U3194 (N_3194,N_2825,N_2997);
nor U3195 (N_3195,N_2931,N_2817);
nand U3196 (N_3196,N_2855,N_2865);
or U3197 (N_3197,N_2964,N_2894);
nor U3198 (N_3198,N_2989,N_2893);
nor U3199 (N_3199,N_2958,N_2835);
nor U3200 (N_3200,N_3065,N_3100);
xnor U3201 (N_3201,N_3165,N_3046);
xor U3202 (N_3202,N_3185,N_3011);
nor U3203 (N_3203,N_3194,N_3150);
nand U3204 (N_3204,N_3197,N_3168);
nand U3205 (N_3205,N_3171,N_3107);
nand U3206 (N_3206,N_3014,N_3003);
or U3207 (N_3207,N_3018,N_3085);
or U3208 (N_3208,N_3053,N_3006);
xor U3209 (N_3209,N_3143,N_3129);
and U3210 (N_3210,N_3043,N_3009);
and U3211 (N_3211,N_3012,N_3141);
xor U3212 (N_3212,N_3158,N_3170);
and U3213 (N_3213,N_3159,N_3049);
nor U3214 (N_3214,N_3115,N_3090);
or U3215 (N_3215,N_3123,N_3041);
nor U3216 (N_3216,N_3054,N_3106);
or U3217 (N_3217,N_3163,N_3005);
nand U3218 (N_3218,N_3152,N_3146);
xnor U3219 (N_3219,N_3151,N_3110);
or U3220 (N_3220,N_3089,N_3099);
nor U3221 (N_3221,N_3020,N_3160);
or U3222 (N_3222,N_3112,N_3025);
and U3223 (N_3223,N_3064,N_3186);
or U3224 (N_3224,N_3010,N_3148);
and U3225 (N_3225,N_3173,N_3080);
and U3226 (N_3226,N_3071,N_3029);
xor U3227 (N_3227,N_3078,N_3136);
and U3228 (N_3228,N_3062,N_3017);
and U3229 (N_3229,N_3030,N_3183);
nand U3230 (N_3230,N_3027,N_3153);
nor U3231 (N_3231,N_3061,N_3087);
xnor U3232 (N_3232,N_3121,N_3024);
nand U3233 (N_3233,N_3075,N_3134);
xnor U3234 (N_3234,N_3188,N_3164);
and U3235 (N_3235,N_3082,N_3138);
or U3236 (N_3236,N_3108,N_3162);
xor U3237 (N_3237,N_3016,N_3036);
or U3238 (N_3238,N_3147,N_3149);
nand U3239 (N_3239,N_3069,N_3076);
nand U3240 (N_3240,N_3066,N_3126);
nand U3241 (N_3241,N_3023,N_3144);
nor U3242 (N_3242,N_3072,N_3093);
and U3243 (N_3243,N_3068,N_3174);
or U3244 (N_3244,N_3088,N_3033);
xor U3245 (N_3245,N_3119,N_3133);
nor U3246 (N_3246,N_3103,N_3037);
xor U3247 (N_3247,N_3028,N_3092);
or U3248 (N_3248,N_3105,N_3137);
nor U3249 (N_3249,N_3187,N_3145);
nand U3250 (N_3250,N_3081,N_3169);
nand U3251 (N_3251,N_3074,N_3191);
nor U3252 (N_3252,N_3180,N_3077);
nand U3253 (N_3253,N_3166,N_3083);
and U3254 (N_3254,N_3142,N_3155);
or U3255 (N_3255,N_3199,N_3007);
nand U3256 (N_3256,N_3176,N_3032);
nor U3257 (N_3257,N_3084,N_3095);
nor U3258 (N_3258,N_3038,N_3048);
nor U3259 (N_3259,N_3052,N_3125);
xnor U3260 (N_3260,N_3157,N_3161);
xor U3261 (N_3261,N_3022,N_3198);
or U3262 (N_3262,N_3127,N_3175);
or U3263 (N_3263,N_3113,N_3190);
and U3264 (N_3264,N_3111,N_3139);
nand U3265 (N_3265,N_3177,N_3181);
and U3266 (N_3266,N_3130,N_3086);
nand U3267 (N_3267,N_3104,N_3102);
and U3268 (N_3268,N_3091,N_3118);
nand U3269 (N_3269,N_3040,N_3096);
or U3270 (N_3270,N_3067,N_3109);
xnor U3271 (N_3271,N_3044,N_3192);
nor U3272 (N_3272,N_3013,N_3124);
nor U3273 (N_3273,N_3117,N_3196);
and U3274 (N_3274,N_3034,N_3042);
xor U3275 (N_3275,N_3131,N_3132);
nand U3276 (N_3276,N_3179,N_3008);
and U3277 (N_3277,N_3114,N_3097);
xnor U3278 (N_3278,N_3098,N_3116);
nand U3279 (N_3279,N_3128,N_3002);
nand U3280 (N_3280,N_3178,N_3156);
nor U3281 (N_3281,N_3055,N_3059);
xor U3282 (N_3282,N_3057,N_3172);
or U3283 (N_3283,N_3001,N_3039);
nor U3284 (N_3284,N_3045,N_3050);
nand U3285 (N_3285,N_3094,N_3167);
or U3286 (N_3286,N_3079,N_3193);
or U3287 (N_3287,N_3140,N_3000);
and U3288 (N_3288,N_3019,N_3135);
xor U3289 (N_3289,N_3004,N_3051);
and U3290 (N_3290,N_3060,N_3026);
nand U3291 (N_3291,N_3122,N_3063);
nand U3292 (N_3292,N_3015,N_3101);
or U3293 (N_3293,N_3035,N_3154);
nand U3294 (N_3294,N_3195,N_3056);
or U3295 (N_3295,N_3184,N_3058);
nor U3296 (N_3296,N_3073,N_3031);
or U3297 (N_3297,N_3189,N_3021);
nor U3298 (N_3298,N_3120,N_3070);
nor U3299 (N_3299,N_3182,N_3047);
xnor U3300 (N_3300,N_3162,N_3138);
or U3301 (N_3301,N_3121,N_3063);
or U3302 (N_3302,N_3100,N_3024);
or U3303 (N_3303,N_3052,N_3104);
xor U3304 (N_3304,N_3114,N_3042);
nand U3305 (N_3305,N_3110,N_3028);
or U3306 (N_3306,N_3048,N_3191);
and U3307 (N_3307,N_3147,N_3174);
nor U3308 (N_3308,N_3189,N_3003);
nand U3309 (N_3309,N_3110,N_3194);
nand U3310 (N_3310,N_3087,N_3068);
nor U3311 (N_3311,N_3125,N_3133);
xor U3312 (N_3312,N_3082,N_3150);
and U3313 (N_3313,N_3032,N_3072);
nand U3314 (N_3314,N_3103,N_3068);
and U3315 (N_3315,N_3104,N_3094);
or U3316 (N_3316,N_3116,N_3128);
and U3317 (N_3317,N_3187,N_3161);
xnor U3318 (N_3318,N_3189,N_3078);
or U3319 (N_3319,N_3162,N_3086);
nand U3320 (N_3320,N_3029,N_3164);
nand U3321 (N_3321,N_3183,N_3173);
or U3322 (N_3322,N_3000,N_3093);
nand U3323 (N_3323,N_3083,N_3151);
and U3324 (N_3324,N_3069,N_3170);
or U3325 (N_3325,N_3088,N_3067);
or U3326 (N_3326,N_3034,N_3072);
and U3327 (N_3327,N_3140,N_3176);
xor U3328 (N_3328,N_3058,N_3116);
xor U3329 (N_3329,N_3017,N_3009);
nand U3330 (N_3330,N_3074,N_3023);
nor U3331 (N_3331,N_3195,N_3085);
and U3332 (N_3332,N_3173,N_3056);
xor U3333 (N_3333,N_3150,N_3123);
or U3334 (N_3334,N_3058,N_3130);
and U3335 (N_3335,N_3168,N_3118);
or U3336 (N_3336,N_3128,N_3009);
nor U3337 (N_3337,N_3049,N_3178);
nor U3338 (N_3338,N_3076,N_3188);
nand U3339 (N_3339,N_3177,N_3013);
nor U3340 (N_3340,N_3173,N_3015);
nor U3341 (N_3341,N_3152,N_3138);
xor U3342 (N_3342,N_3073,N_3161);
nor U3343 (N_3343,N_3075,N_3182);
and U3344 (N_3344,N_3130,N_3153);
and U3345 (N_3345,N_3175,N_3177);
and U3346 (N_3346,N_3129,N_3102);
or U3347 (N_3347,N_3084,N_3025);
or U3348 (N_3348,N_3117,N_3126);
nor U3349 (N_3349,N_3143,N_3083);
xnor U3350 (N_3350,N_3106,N_3164);
xnor U3351 (N_3351,N_3093,N_3170);
nand U3352 (N_3352,N_3149,N_3007);
and U3353 (N_3353,N_3163,N_3172);
xor U3354 (N_3354,N_3016,N_3131);
or U3355 (N_3355,N_3199,N_3025);
nand U3356 (N_3356,N_3021,N_3056);
and U3357 (N_3357,N_3025,N_3056);
nand U3358 (N_3358,N_3042,N_3049);
xor U3359 (N_3359,N_3160,N_3126);
or U3360 (N_3360,N_3132,N_3192);
or U3361 (N_3361,N_3028,N_3016);
or U3362 (N_3362,N_3155,N_3064);
xor U3363 (N_3363,N_3170,N_3101);
xnor U3364 (N_3364,N_3094,N_3120);
xnor U3365 (N_3365,N_3129,N_3192);
nor U3366 (N_3366,N_3125,N_3014);
or U3367 (N_3367,N_3024,N_3079);
and U3368 (N_3368,N_3090,N_3028);
nor U3369 (N_3369,N_3113,N_3058);
and U3370 (N_3370,N_3017,N_3000);
and U3371 (N_3371,N_3164,N_3099);
nor U3372 (N_3372,N_3100,N_3171);
and U3373 (N_3373,N_3047,N_3183);
and U3374 (N_3374,N_3064,N_3013);
and U3375 (N_3375,N_3152,N_3150);
xnor U3376 (N_3376,N_3142,N_3151);
or U3377 (N_3377,N_3185,N_3042);
nand U3378 (N_3378,N_3142,N_3092);
xnor U3379 (N_3379,N_3012,N_3113);
nor U3380 (N_3380,N_3145,N_3061);
and U3381 (N_3381,N_3006,N_3077);
nand U3382 (N_3382,N_3174,N_3096);
and U3383 (N_3383,N_3048,N_3034);
nand U3384 (N_3384,N_3003,N_3193);
xnor U3385 (N_3385,N_3053,N_3192);
and U3386 (N_3386,N_3082,N_3005);
and U3387 (N_3387,N_3066,N_3142);
or U3388 (N_3388,N_3011,N_3038);
nand U3389 (N_3389,N_3063,N_3037);
and U3390 (N_3390,N_3009,N_3055);
nand U3391 (N_3391,N_3002,N_3045);
and U3392 (N_3392,N_3031,N_3101);
nor U3393 (N_3393,N_3199,N_3056);
nor U3394 (N_3394,N_3149,N_3059);
nand U3395 (N_3395,N_3089,N_3015);
or U3396 (N_3396,N_3005,N_3144);
and U3397 (N_3397,N_3003,N_3186);
nor U3398 (N_3398,N_3106,N_3170);
nand U3399 (N_3399,N_3118,N_3128);
xor U3400 (N_3400,N_3292,N_3247);
or U3401 (N_3401,N_3223,N_3351);
xnor U3402 (N_3402,N_3248,N_3375);
and U3403 (N_3403,N_3296,N_3327);
nor U3404 (N_3404,N_3206,N_3253);
or U3405 (N_3405,N_3383,N_3340);
nor U3406 (N_3406,N_3262,N_3257);
and U3407 (N_3407,N_3322,N_3236);
and U3408 (N_3408,N_3226,N_3214);
nand U3409 (N_3409,N_3337,N_3398);
nor U3410 (N_3410,N_3303,N_3225);
or U3411 (N_3411,N_3323,N_3205);
or U3412 (N_3412,N_3355,N_3361);
nor U3413 (N_3413,N_3356,N_3370);
nor U3414 (N_3414,N_3250,N_3229);
nor U3415 (N_3415,N_3260,N_3343);
or U3416 (N_3416,N_3273,N_3228);
xnor U3417 (N_3417,N_3231,N_3338);
xor U3418 (N_3418,N_3298,N_3268);
nand U3419 (N_3419,N_3334,N_3290);
nand U3420 (N_3420,N_3215,N_3316);
nor U3421 (N_3421,N_3332,N_3300);
or U3422 (N_3422,N_3299,N_3382);
xnor U3423 (N_3423,N_3364,N_3384);
or U3424 (N_3424,N_3310,N_3251);
or U3425 (N_3425,N_3208,N_3376);
nand U3426 (N_3426,N_3213,N_3246);
nor U3427 (N_3427,N_3220,N_3278);
or U3428 (N_3428,N_3390,N_3272);
or U3429 (N_3429,N_3365,N_3305);
xnor U3430 (N_3430,N_3385,N_3238);
nand U3431 (N_3431,N_3200,N_3313);
xnor U3432 (N_3432,N_3397,N_3325);
nand U3433 (N_3433,N_3302,N_3319);
and U3434 (N_3434,N_3381,N_3359);
nor U3435 (N_3435,N_3221,N_3371);
and U3436 (N_3436,N_3308,N_3212);
and U3437 (N_3437,N_3263,N_3341);
nor U3438 (N_3438,N_3367,N_3222);
nand U3439 (N_3439,N_3320,N_3387);
nor U3440 (N_3440,N_3346,N_3318);
nand U3441 (N_3441,N_3286,N_3315);
xnor U3442 (N_3442,N_3269,N_3288);
xor U3443 (N_3443,N_3211,N_3209);
and U3444 (N_3444,N_3216,N_3306);
and U3445 (N_3445,N_3349,N_3330);
and U3446 (N_3446,N_3396,N_3307);
xor U3447 (N_3447,N_3333,N_3280);
nand U3448 (N_3448,N_3287,N_3284);
nand U3449 (N_3449,N_3264,N_3389);
or U3450 (N_3450,N_3274,N_3378);
nand U3451 (N_3451,N_3276,N_3369);
or U3452 (N_3452,N_3230,N_3244);
and U3453 (N_3453,N_3345,N_3314);
nor U3454 (N_3454,N_3358,N_3350);
nand U3455 (N_3455,N_3394,N_3321);
nand U3456 (N_3456,N_3353,N_3224);
xnor U3457 (N_3457,N_3277,N_3399);
and U3458 (N_3458,N_3283,N_3347);
nand U3459 (N_3459,N_3372,N_3336);
nor U3460 (N_3460,N_3218,N_3261);
or U3461 (N_3461,N_3344,N_3291);
nand U3462 (N_3462,N_3258,N_3335);
nor U3463 (N_3463,N_3379,N_3328);
nor U3464 (N_3464,N_3324,N_3219);
and U3465 (N_3465,N_3282,N_3256);
nor U3466 (N_3466,N_3309,N_3210);
xor U3467 (N_3467,N_3240,N_3392);
or U3468 (N_3468,N_3342,N_3326);
or U3469 (N_3469,N_3239,N_3254);
xnor U3470 (N_3470,N_3373,N_3203);
xnor U3471 (N_3471,N_3279,N_3204);
nand U3472 (N_3472,N_3304,N_3255);
or U3473 (N_3473,N_3377,N_3386);
xnor U3474 (N_3474,N_3252,N_3360);
nor U3475 (N_3475,N_3395,N_3391);
xnor U3476 (N_3476,N_3301,N_3388);
or U3477 (N_3477,N_3235,N_3232);
and U3478 (N_3478,N_3234,N_3352);
nand U3479 (N_3479,N_3317,N_3297);
or U3480 (N_3480,N_3201,N_3339);
nor U3481 (N_3481,N_3366,N_3241);
or U3482 (N_3482,N_3259,N_3265);
nor U3483 (N_3483,N_3202,N_3271);
nor U3484 (N_3484,N_3362,N_3281);
nor U3485 (N_3485,N_3207,N_3233);
nor U3486 (N_3486,N_3294,N_3237);
nand U3487 (N_3487,N_3311,N_3374);
nand U3488 (N_3488,N_3393,N_3293);
and U3489 (N_3489,N_3275,N_3354);
nor U3490 (N_3490,N_3329,N_3331);
nand U3491 (N_3491,N_3295,N_3363);
or U3492 (N_3492,N_3243,N_3348);
nor U3493 (N_3493,N_3289,N_3368);
and U3494 (N_3494,N_3242,N_3312);
nor U3495 (N_3495,N_3227,N_3270);
or U3496 (N_3496,N_3357,N_3249);
xnor U3497 (N_3497,N_3285,N_3267);
and U3498 (N_3498,N_3245,N_3217);
or U3499 (N_3499,N_3380,N_3266);
and U3500 (N_3500,N_3355,N_3269);
and U3501 (N_3501,N_3381,N_3210);
nor U3502 (N_3502,N_3304,N_3272);
nor U3503 (N_3503,N_3282,N_3305);
and U3504 (N_3504,N_3200,N_3317);
xnor U3505 (N_3505,N_3270,N_3342);
nor U3506 (N_3506,N_3210,N_3261);
nand U3507 (N_3507,N_3354,N_3394);
xnor U3508 (N_3508,N_3366,N_3295);
and U3509 (N_3509,N_3389,N_3262);
xnor U3510 (N_3510,N_3385,N_3247);
or U3511 (N_3511,N_3303,N_3226);
or U3512 (N_3512,N_3345,N_3216);
and U3513 (N_3513,N_3325,N_3323);
nand U3514 (N_3514,N_3293,N_3268);
nor U3515 (N_3515,N_3286,N_3262);
nand U3516 (N_3516,N_3204,N_3381);
or U3517 (N_3517,N_3377,N_3332);
or U3518 (N_3518,N_3328,N_3301);
or U3519 (N_3519,N_3274,N_3257);
or U3520 (N_3520,N_3255,N_3201);
and U3521 (N_3521,N_3321,N_3276);
nand U3522 (N_3522,N_3391,N_3325);
or U3523 (N_3523,N_3338,N_3395);
nor U3524 (N_3524,N_3239,N_3377);
and U3525 (N_3525,N_3219,N_3320);
xor U3526 (N_3526,N_3240,N_3209);
nor U3527 (N_3527,N_3329,N_3323);
nand U3528 (N_3528,N_3356,N_3376);
nand U3529 (N_3529,N_3310,N_3340);
nor U3530 (N_3530,N_3374,N_3361);
or U3531 (N_3531,N_3226,N_3223);
and U3532 (N_3532,N_3256,N_3291);
and U3533 (N_3533,N_3301,N_3234);
or U3534 (N_3534,N_3339,N_3220);
and U3535 (N_3535,N_3291,N_3263);
nand U3536 (N_3536,N_3262,N_3302);
or U3537 (N_3537,N_3207,N_3276);
nor U3538 (N_3538,N_3394,N_3308);
nor U3539 (N_3539,N_3289,N_3388);
or U3540 (N_3540,N_3287,N_3239);
xor U3541 (N_3541,N_3346,N_3330);
and U3542 (N_3542,N_3215,N_3257);
or U3543 (N_3543,N_3258,N_3271);
nor U3544 (N_3544,N_3342,N_3203);
or U3545 (N_3545,N_3290,N_3203);
or U3546 (N_3546,N_3311,N_3283);
and U3547 (N_3547,N_3292,N_3346);
nand U3548 (N_3548,N_3389,N_3268);
nand U3549 (N_3549,N_3342,N_3208);
nor U3550 (N_3550,N_3300,N_3216);
nor U3551 (N_3551,N_3396,N_3332);
or U3552 (N_3552,N_3202,N_3240);
nand U3553 (N_3553,N_3313,N_3333);
nand U3554 (N_3554,N_3277,N_3238);
and U3555 (N_3555,N_3369,N_3214);
nor U3556 (N_3556,N_3224,N_3227);
and U3557 (N_3557,N_3236,N_3229);
nand U3558 (N_3558,N_3331,N_3252);
xnor U3559 (N_3559,N_3273,N_3339);
nand U3560 (N_3560,N_3258,N_3201);
or U3561 (N_3561,N_3233,N_3292);
or U3562 (N_3562,N_3218,N_3359);
nand U3563 (N_3563,N_3268,N_3381);
xnor U3564 (N_3564,N_3253,N_3385);
or U3565 (N_3565,N_3314,N_3247);
and U3566 (N_3566,N_3359,N_3317);
nor U3567 (N_3567,N_3219,N_3225);
nor U3568 (N_3568,N_3351,N_3218);
nand U3569 (N_3569,N_3347,N_3354);
and U3570 (N_3570,N_3338,N_3274);
nand U3571 (N_3571,N_3369,N_3347);
nand U3572 (N_3572,N_3232,N_3305);
nor U3573 (N_3573,N_3317,N_3329);
and U3574 (N_3574,N_3272,N_3395);
and U3575 (N_3575,N_3256,N_3391);
or U3576 (N_3576,N_3393,N_3302);
and U3577 (N_3577,N_3204,N_3202);
and U3578 (N_3578,N_3397,N_3262);
or U3579 (N_3579,N_3275,N_3227);
xnor U3580 (N_3580,N_3236,N_3238);
nor U3581 (N_3581,N_3319,N_3278);
or U3582 (N_3582,N_3341,N_3209);
nor U3583 (N_3583,N_3325,N_3266);
and U3584 (N_3584,N_3302,N_3347);
nor U3585 (N_3585,N_3379,N_3283);
nand U3586 (N_3586,N_3380,N_3206);
xnor U3587 (N_3587,N_3347,N_3212);
and U3588 (N_3588,N_3213,N_3386);
or U3589 (N_3589,N_3231,N_3359);
nor U3590 (N_3590,N_3282,N_3286);
xnor U3591 (N_3591,N_3305,N_3394);
nor U3592 (N_3592,N_3308,N_3386);
and U3593 (N_3593,N_3219,N_3304);
nand U3594 (N_3594,N_3268,N_3380);
xnor U3595 (N_3595,N_3211,N_3312);
or U3596 (N_3596,N_3345,N_3213);
nand U3597 (N_3597,N_3271,N_3234);
nand U3598 (N_3598,N_3223,N_3365);
nand U3599 (N_3599,N_3346,N_3293);
and U3600 (N_3600,N_3444,N_3574);
nor U3601 (N_3601,N_3402,N_3523);
or U3602 (N_3602,N_3504,N_3415);
or U3603 (N_3603,N_3485,N_3406);
nor U3604 (N_3604,N_3526,N_3508);
nand U3605 (N_3605,N_3422,N_3491);
xor U3606 (N_3606,N_3404,N_3528);
xor U3607 (N_3607,N_3442,N_3494);
or U3608 (N_3608,N_3515,N_3496);
xnor U3609 (N_3609,N_3545,N_3581);
xor U3610 (N_3610,N_3423,N_3480);
xnor U3611 (N_3611,N_3409,N_3567);
nor U3612 (N_3612,N_3456,N_3419);
xnor U3613 (N_3613,N_3553,N_3594);
xor U3614 (N_3614,N_3477,N_3489);
nand U3615 (N_3615,N_3461,N_3583);
or U3616 (N_3616,N_3450,N_3519);
and U3617 (N_3617,N_3412,N_3546);
or U3618 (N_3618,N_3452,N_3591);
nor U3619 (N_3619,N_3410,N_3454);
and U3620 (N_3620,N_3598,N_3414);
or U3621 (N_3621,N_3467,N_3441);
and U3622 (N_3622,N_3436,N_3498);
xor U3623 (N_3623,N_3476,N_3455);
nor U3624 (N_3624,N_3405,N_3503);
or U3625 (N_3625,N_3544,N_3522);
and U3626 (N_3626,N_3554,N_3472);
or U3627 (N_3627,N_3537,N_3445);
nor U3628 (N_3628,N_3536,N_3524);
nand U3629 (N_3629,N_3408,N_3400);
nor U3630 (N_3630,N_3509,N_3425);
nand U3631 (N_3631,N_3540,N_3571);
nor U3632 (N_3632,N_3453,N_3507);
or U3633 (N_3633,N_3428,N_3527);
xnor U3634 (N_3634,N_3584,N_3449);
nor U3635 (N_3635,N_3587,N_3438);
nand U3636 (N_3636,N_3579,N_3474);
xor U3637 (N_3637,N_3520,N_3578);
and U3638 (N_3638,N_3559,N_3557);
xnor U3639 (N_3639,N_3435,N_3471);
nand U3640 (N_3640,N_3586,N_3532);
and U3641 (N_3641,N_3563,N_3403);
or U3642 (N_3642,N_3458,N_3466);
xor U3643 (N_3643,N_3549,N_3552);
or U3644 (N_3644,N_3413,N_3473);
and U3645 (N_3645,N_3558,N_3575);
nor U3646 (N_3646,N_3470,N_3529);
xor U3647 (N_3647,N_3533,N_3421);
or U3648 (N_3648,N_3514,N_3463);
nand U3649 (N_3649,N_3577,N_3501);
xnor U3650 (N_3650,N_3551,N_3426);
nand U3651 (N_3651,N_3430,N_3550);
or U3652 (N_3652,N_3411,N_3510);
nand U3653 (N_3653,N_3490,N_3561);
nor U3654 (N_3654,N_3499,N_3418);
and U3655 (N_3655,N_3506,N_3599);
and U3656 (N_3656,N_3566,N_3596);
nor U3657 (N_3657,N_3542,N_3483);
and U3658 (N_3658,N_3431,N_3565);
or U3659 (N_3659,N_3478,N_3416);
or U3660 (N_3660,N_3525,N_3459);
or U3661 (N_3661,N_3429,N_3502);
or U3662 (N_3662,N_3576,N_3541);
xnor U3663 (N_3663,N_3548,N_3481);
nor U3664 (N_3664,N_3569,N_3464);
or U3665 (N_3665,N_3447,N_3517);
or U3666 (N_3666,N_3564,N_3488);
and U3667 (N_3667,N_3516,N_3448);
and U3668 (N_3668,N_3432,N_3512);
nor U3669 (N_3669,N_3420,N_3484);
and U3670 (N_3670,N_3457,N_3497);
nor U3671 (N_3671,N_3595,N_3547);
nand U3672 (N_3672,N_3437,N_3534);
nor U3673 (N_3673,N_3585,N_3556);
nand U3674 (N_3674,N_3590,N_3588);
nor U3675 (N_3675,N_3487,N_3479);
xor U3676 (N_3676,N_3492,N_3500);
and U3677 (N_3677,N_3424,N_3568);
xnor U3678 (N_3678,N_3562,N_3593);
or U3679 (N_3679,N_3535,N_3469);
nor U3680 (N_3680,N_3417,N_3531);
or U3681 (N_3681,N_3407,N_3592);
nand U3682 (N_3682,N_3589,N_3538);
xnor U3683 (N_3683,N_3427,N_3475);
nor U3684 (N_3684,N_3539,N_3434);
nor U3685 (N_3685,N_3468,N_3433);
nor U3686 (N_3686,N_3495,N_3513);
and U3687 (N_3687,N_3570,N_3401);
nor U3688 (N_3688,N_3560,N_3597);
nand U3689 (N_3689,N_3572,N_3573);
or U3690 (N_3690,N_3482,N_3443);
nor U3691 (N_3691,N_3486,N_3582);
nand U3692 (N_3692,N_3505,N_3518);
xnor U3693 (N_3693,N_3511,N_3555);
nand U3694 (N_3694,N_3439,N_3460);
nor U3695 (N_3695,N_3451,N_3521);
and U3696 (N_3696,N_3493,N_3543);
or U3697 (N_3697,N_3465,N_3462);
or U3698 (N_3698,N_3446,N_3530);
and U3699 (N_3699,N_3580,N_3440);
nor U3700 (N_3700,N_3505,N_3503);
nand U3701 (N_3701,N_3464,N_3568);
xor U3702 (N_3702,N_3455,N_3420);
xnor U3703 (N_3703,N_3526,N_3547);
and U3704 (N_3704,N_3542,N_3554);
nand U3705 (N_3705,N_3511,N_3491);
nor U3706 (N_3706,N_3520,N_3448);
xnor U3707 (N_3707,N_3514,N_3526);
or U3708 (N_3708,N_3484,N_3490);
and U3709 (N_3709,N_3562,N_3503);
xnor U3710 (N_3710,N_3468,N_3415);
xor U3711 (N_3711,N_3407,N_3591);
xnor U3712 (N_3712,N_3539,N_3424);
or U3713 (N_3713,N_3564,N_3593);
or U3714 (N_3714,N_3509,N_3429);
and U3715 (N_3715,N_3447,N_3479);
nor U3716 (N_3716,N_3552,N_3432);
xnor U3717 (N_3717,N_3525,N_3424);
nor U3718 (N_3718,N_3488,N_3415);
xor U3719 (N_3719,N_3575,N_3482);
and U3720 (N_3720,N_3444,N_3596);
nor U3721 (N_3721,N_3541,N_3490);
xor U3722 (N_3722,N_3417,N_3569);
xor U3723 (N_3723,N_3564,N_3574);
and U3724 (N_3724,N_3470,N_3581);
and U3725 (N_3725,N_3502,N_3436);
nand U3726 (N_3726,N_3474,N_3592);
nor U3727 (N_3727,N_3421,N_3577);
nor U3728 (N_3728,N_3507,N_3458);
nand U3729 (N_3729,N_3421,N_3405);
xor U3730 (N_3730,N_3507,N_3530);
nand U3731 (N_3731,N_3591,N_3428);
or U3732 (N_3732,N_3586,N_3453);
xor U3733 (N_3733,N_3425,N_3528);
xnor U3734 (N_3734,N_3483,N_3461);
nor U3735 (N_3735,N_3502,N_3527);
xor U3736 (N_3736,N_3464,N_3514);
nand U3737 (N_3737,N_3404,N_3406);
xnor U3738 (N_3738,N_3514,N_3537);
or U3739 (N_3739,N_3529,N_3498);
nor U3740 (N_3740,N_3424,N_3548);
and U3741 (N_3741,N_3421,N_3581);
nor U3742 (N_3742,N_3508,N_3510);
xor U3743 (N_3743,N_3572,N_3551);
and U3744 (N_3744,N_3577,N_3466);
and U3745 (N_3745,N_3599,N_3491);
and U3746 (N_3746,N_3401,N_3592);
nand U3747 (N_3747,N_3527,N_3444);
nor U3748 (N_3748,N_3573,N_3542);
xor U3749 (N_3749,N_3535,N_3455);
nor U3750 (N_3750,N_3472,N_3507);
nor U3751 (N_3751,N_3482,N_3537);
nand U3752 (N_3752,N_3561,N_3500);
and U3753 (N_3753,N_3465,N_3444);
and U3754 (N_3754,N_3548,N_3549);
xor U3755 (N_3755,N_3543,N_3554);
and U3756 (N_3756,N_3544,N_3425);
or U3757 (N_3757,N_3429,N_3507);
or U3758 (N_3758,N_3535,N_3473);
xor U3759 (N_3759,N_3516,N_3541);
nor U3760 (N_3760,N_3575,N_3530);
and U3761 (N_3761,N_3589,N_3553);
nor U3762 (N_3762,N_3454,N_3510);
nor U3763 (N_3763,N_3516,N_3442);
nand U3764 (N_3764,N_3404,N_3551);
and U3765 (N_3765,N_3506,N_3482);
xnor U3766 (N_3766,N_3597,N_3583);
xnor U3767 (N_3767,N_3519,N_3506);
or U3768 (N_3768,N_3400,N_3474);
and U3769 (N_3769,N_3502,N_3469);
and U3770 (N_3770,N_3470,N_3532);
and U3771 (N_3771,N_3443,N_3455);
xor U3772 (N_3772,N_3475,N_3563);
or U3773 (N_3773,N_3426,N_3425);
and U3774 (N_3774,N_3479,N_3522);
nor U3775 (N_3775,N_3445,N_3435);
nand U3776 (N_3776,N_3588,N_3474);
and U3777 (N_3777,N_3479,N_3558);
and U3778 (N_3778,N_3528,N_3426);
and U3779 (N_3779,N_3567,N_3586);
nor U3780 (N_3780,N_3595,N_3470);
nand U3781 (N_3781,N_3529,N_3489);
and U3782 (N_3782,N_3462,N_3438);
xor U3783 (N_3783,N_3503,N_3539);
nor U3784 (N_3784,N_3500,N_3579);
and U3785 (N_3785,N_3539,N_3488);
nor U3786 (N_3786,N_3554,N_3461);
nor U3787 (N_3787,N_3442,N_3562);
nand U3788 (N_3788,N_3573,N_3552);
nor U3789 (N_3789,N_3597,N_3413);
and U3790 (N_3790,N_3446,N_3407);
or U3791 (N_3791,N_3524,N_3587);
nor U3792 (N_3792,N_3540,N_3445);
xnor U3793 (N_3793,N_3476,N_3556);
xor U3794 (N_3794,N_3543,N_3549);
xnor U3795 (N_3795,N_3518,N_3465);
nor U3796 (N_3796,N_3509,N_3524);
nand U3797 (N_3797,N_3410,N_3400);
and U3798 (N_3798,N_3598,N_3454);
or U3799 (N_3799,N_3597,N_3578);
nand U3800 (N_3800,N_3700,N_3604);
nor U3801 (N_3801,N_3768,N_3716);
nand U3802 (N_3802,N_3729,N_3738);
nand U3803 (N_3803,N_3735,N_3777);
nor U3804 (N_3804,N_3708,N_3649);
nor U3805 (N_3805,N_3681,N_3781);
nand U3806 (N_3806,N_3683,N_3602);
nand U3807 (N_3807,N_3614,N_3761);
and U3808 (N_3808,N_3692,N_3611);
nand U3809 (N_3809,N_3736,N_3728);
or U3810 (N_3810,N_3770,N_3744);
nand U3811 (N_3811,N_3685,N_3607);
or U3812 (N_3812,N_3684,N_3663);
nand U3813 (N_3813,N_3665,N_3751);
xor U3814 (N_3814,N_3620,N_3757);
or U3815 (N_3815,N_3606,N_3696);
and U3816 (N_3816,N_3627,N_3646);
and U3817 (N_3817,N_3706,N_3662);
and U3818 (N_3818,N_3730,N_3689);
or U3819 (N_3819,N_3724,N_3687);
xor U3820 (N_3820,N_3609,N_3623);
xnor U3821 (N_3821,N_3795,N_3746);
nand U3822 (N_3822,N_3670,N_3721);
nor U3823 (N_3823,N_3766,N_3686);
and U3824 (N_3824,N_3650,N_3617);
and U3825 (N_3825,N_3771,N_3625);
xnor U3826 (N_3826,N_3657,N_3763);
and U3827 (N_3827,N_3743,N_3754);
and U3828 (N_3828,N_3671,N_3626);
and U3829 (N_3829,N_3737,N_3705);
and U3830 (N_3830,N_3679,N_3747);
xnor U3831 (N_3831,N_3764,N_3673);
nor U3832 (N_3832,N_3655,N_3613);
nor U3833 (N_3833,N_3622,N_3600);
and U3834 (N_3834,N_3779,N_3739);
xnor U3835 (N_3835,N_3782,N_3616);
nor U3836 (N_3836,N_3661,N_3642);
nor U3837 (N_3837,N_3722,N_3667);
nor U3838 (N_3838,N_3758,N_3698);
or U3839 (N_3839,N_3715,N_3636);
nand U3840 (N_3840,N_3783,N_3731);
nor U3841 (N_3841,N_3794,N_3629);
and U3842 (N_3842,N_3682,N_3760);
and U3843 (N_3843,N_3668,N_3714);
xor U3844 (N_3844,N_3778,N_3759);
or U3845 (N_3845,N_3612,N_3719);
and U3846 (N_3846,N_3718,N_3651);
nand U3847 (N_3847,N_3666,N_3643);
nor U3848 (N_3848,N_3704,N_3769);
nor U3849 (N_3849,N_3713,N_3740);
and U3850 (N_3850,N_3695,N_3745);
nor U3851 (N_3851,N_3669,N_3619);
xnor U3852 (N_3852,N_3653,N_3753);
xnor U3853 (N_3853,N_3628,N_3780);
nand U3854 (N_3854,N_3690,N_3772);
and U3855 (N_3855,N_3697,N_3791);
xnor U3856 (N_3856,N_3785,N_3790);
nand U3857 (N_3857,N_3725,N_3637);
nand U3858 (N_3858,N_3752,N_3788);
xnor U3859 (N_3859,N_3678,N_3784);
nand U3860 (N_3860,N_3688,N_3710);
and U3861 (N_3861,N_3796,N_3797);
or U3862 (N_3862,N_3773,N_3787);
nand U3863 (N_3863,N_3749,N_3762);
and U3864 (N_3864,N_3630,N_3798);
xnor U3865 (N_3865,N_3717,N_3632);
xor U3866 (N_3866,N_3742,N_3644);
xnor U3867 (N_3867,N_3755,N_3634);
or U3868 (N_3868,N_3645,N_3635);
and U3869 (N_3869,N_3654,N_3647);
and U3870 (N_3870,N_3641,N_3767);
nor U3871 (N_3871,N_3618,N_3638);
xor U3872 (N_3872,N_3733,N_3691);
or U3873 (N_3873,N_3723,N_3775);
or U3874 (N_3874,N_3660,N_3658);
and U3875 (N_3875,N_3776,N_3610);
and U3876 (N_3876,N_3701,N_3789);
nor U3877 (N_3877,N_3792,N_3608);
nor U3878 (N_3878,N_3605,N_3656);
and U3879 (N_3879,N_3674,N_3709);
nor U3880 (N_3880,N_3799,N_3659);
nand U3881 (N_3881,N_3741,N_3726);
or U3882 (N_3882,N_3615,N_3711);
and U3883 (N_3883,N_3676,N_3664);
or U3884 (N_3884,N_3786,N_3748);
nor U3885 (N_3885,N_3750,N_3631);
and U3886 (N_3886,N_3699,N_3702);
nand U3887 (N_3887,N_3672,N_3793);
xor U3888 (N_3888,N_3774,N_3680);
xnor U3889 (N_3889,N_3756,N_3639);
and U3890 (N_3890,N_3727,N_3734);
or U3891 (N_3891,N_3732,N_3675);
and U3892 (N_3892,N_3633,N_3694);
xor U3893 (N_3893,N_3601,N_3640);
and U3894 (N_3894,N_3677,N_3648);
nor U3895 (N_3895,N_3720,N_3603);
and U3896 (N_3896,N_3652,N_3712);
nor U3897 (N_3897,N_3703,N_3693);
or U3898 (N_3898,N_3765,N_3624);
and U3899 (N_3899,N_3707,N_3621);
or U3900 (N_3900,N_3795,N_3606);
nor U3901 (N_3901,N_3600,N_3760);
nand U3902 (N_3902,N_3755,N_3720);
xnor U3903 (N_3903,N_3718,N_3672);
nor U3904 (N_3904,N_3630,N_3710);
nor U3905 (N_3905,N_3669,N_3607);
nor U3906 (N_3906,N_3788,N_3767);
nor U3907 (N_3907,N_3764,N_3651);
and U3908 (N_3908,N_3614,N_3603);
or U3909 (N_3909,N_3674,N_3794);
or U3910 (N_3910,N_3785,N_3796);
xor U3911 (N_3911,N_3744,N_3653);
or U3912 (N_3912,N_3741,N_3746);
xor U3913 (N_3913,N_3740,N_3605);
xor U3914 (N_3914,N_3730,N_3633);
nor U3915 (N_3915,N_3711,N_3710);
nand U3916 (N_3916,N_3639,N_3761);
xor U3917 (N_3917,N_3631,N_3730);
xor U3918 (N_3918,N_3722,N_3727);
xnor U3919 (N_3919,N_3678,N_3795);
and U3920 (N_3920,N_3752,N_3691);
nand U3921 (N_3921,N_3754,N_3747);
nand U3922 (N_3922,N_3611,N_3605);
xnor U3923 (N_3923,N_3759,N_3770);
nor U3924 (N_3924,N_3613,N_3774);
nand U3925 (N_3925,N_3620,N_3656);
nand U3926 (N_3926,N_3601,N_3605);
nand U3927 (N_3927,N_3672,N_3678);
nand U3928 (N_3928,N_3720,N_3600);
or U3929 (N_3929,N_3750,N_3603);
xnor U3930 (N_3930,N_3651,N_3645);
or U3931 (N_3931,N_3624,N_3616);
nand U3932 (N_3932,N_3750,N_3725);
and U3933 (N_3933,N_3639,N_3648);
nor U3934 (N_3934,N_3769,N_3714);
nand U3935 (N_3935,N_3633,N_3620);
nand U3936 (N_3936,N_3776,N_3682);
nor U3937 (N_3937,N_3739,N_3713);
xnor U3938 (N_3938,N_3609,N_3799);
nand U3939 (N_3939,N_3765,N_3675);
nand U3940 (N_3940,N_3697,N_3784);
and U3941 (N_3941,N_3648,N_3759);
nor U3942 (N_3942,N_3790,N_3736);
nor U3943 (N_3943,N_3714,N_3751);
xor U3944 (N_3944,N_3698,N_3607);
nor U3945 (N_3945,N_3685,N_3797);
and U3946 (N_3946,N_3794,N_3764);
nor U3947 (N_3947,N_3636,N_3610);
and U3948 (N_3948,N_3747,N_3781);
and U3949 (N_3949,N_3739,N_3603);
xnor U3950 (N_3950,N_3745,N_3728);
or U3951 (N_3951,N_3728,N_3603);
nand U3952 (N_3952,N_3769,N_3632);
nor U3953 (N_3953,N_3690,N_3644);
or U3954 (N_3954,N_3743,N_3670);
and U3955 (N_3955,N_3719,N_3737);
nor U3956 (N_3956,N_3736,N_3610);
or U3957 (N_3957,N_3710,N_3697);
nand U3958 (N_3958,N_3757,N_3787);
xnor U3959 (N_3959,N_3683,N_3725);
nor U3960 (N_3960,N_3746,N_3727);
xor U3961 (N_3961,N_3648,N_3619);
or U3962 (N_3962,N_3736,N_3717);
xor U3963 (N_3963,N_3738,N_3678);
xnor U3964 (N_3964,N_3778,N_3791);
nor U3965 (N_3965,N_3780,N_3646);
or U3966 (N_3966,N_3619,N_3771);
nand U3967 (N_3967,N_3727,N_3642);
nor U3968 (N_3968,N_3660,N_3644);
xor U3969 (N_3969,N_3694,N_3650);
or U3970 (N_3970,N_3710,N_3616);
and U3971 (N_3971,N_3636,N_3656);
nand U3972 (N_3972,N_3671,N_3698);
nand U3973 (N_3973,N_3706,N_3711);
nor U3974 (N_3974,N_3720,N_3799);
or U3975 (N_3975,N_3614,N_3650);
nand U3976 (N_3976,N_3633,N_3678);
xnor U3977 (N_3977,N_3732,N_3678);
nand U3978 (N_3978,N_3662,N_3734);
nor U3979 (N_3979,N_3743,N_3733);
nand U3980 (N_3980,N_3676,N_3626);
nand U3981 (N_3981,N_3738,N_3653);
nor U3982 (N_3982,N_3627,N_3711);
or U3983 (N_3983,N_3768,N_3625);
or U3984 (N_3984,N_3753,N_3618);
xnor U3985 (N_3985,N_3748,N_3681);
nand U3986 (N_3986,N_3733,N_3735);
nand U3987 (N_3987,N_3641,N_3728);
and U3988 (N_3988,N_3636,N_3764);
nor U3989 (N_3989,N_3689,N_3657);
and U3990 (N_3990,N_3753,N_3716);
and U3991 (N_3991,N_3605,N_3641);
nor U3992 (N_3992,N_3769,N_3785);
xor U3993 (N_3993,N_3740,N_3636);
nand U3994 (N_3994,N_3792,N_3727);
xor U3995 (N_3995,N_3782,N_3706);
and U3996 (N_3996,N_3712,N_3631);
xnor U3997 (N_3997,N_3764,N_3606);
xnor U3998 (N_3998,N_3755,N_3601);
nor U3999 (N_3999,N_3676,N_3723);
nor U4000 (N_4000,N_3932,N_3933);
or U4001 (N_4001,N_3982,N_3956);
and U4002 (N_4002,N_3818,N_3941);
or U4003 (N_4003,N_3986,N_3963);
nor U4004 (N_4004,N_3997,N_3931);
or U4005 (N_4005,N_3924,N_3875);
or U4006 (N_4006,N_3883,N_3993);
and U4007 (N_4007,N_3939,N_3836);
nor U4008 (N_4008,N_3965,N_3915);
nor U4009 (N_4009,N_3888,N_3848);
xnor U4010 (N_4010,N_3847,N_3944);
xnor U4011 (N_4011,N_3830,N_3892);
and U4012 (N_4012,N_3996,N_3910);
xnor U4013 (N_4013,N_3887,N_3907);
xnor U4014 (N_4014,N_3948,N_3897);
nor U4015 (N_4015,N_3821,N_3958);
nand U4016 (N_4016,N_3951,N_3813);
and U4017 (N_4017,N_3994,N_3942);
and U4018 (N_4018,N_3878,N_3876);
xor U4019 (N_4019,N_3985,N_3834);
or U4020 (N_4020,N_3843,N_3862);
nand U4021 (N_4021,N_3952,N_3937);
xnor U4022 (N_4022,N_3844,N_3842);
or U4023 (N_4023,N_3895,N_3811);
nand U4024 (N_4024,N_3970,N_3850);
nor U4025 (N_4025,N_3854,N_3868);
or U4026 (N_4026,N_3992,N_3901);
xor U4027 (N_4027,N_3858,N_3825);
nor U4028 (N_4028,N_3804,N_3886);
xor U4029 (N_4029,N_3802,N_3855);
and U4030 (N_4030,N_3954,N_3906);
nor U4031 (N_4031,N_3926,N_3999);
or U4032 (N_4032,N_3968,N_3902);
xor U4033 (N_4033,N_3927,N_3989);
or U4034 (N_4034,N_3814,N_3874);
or U4035 (N_4035,N_3820,N_3950);
or U4036 (N_4036,N_3987,N_3961);
xnor U4037 (N_4037,N_3881,N_3940);
or U4038 (N_4038,N_3998,N_3810);
or U4039 (N_4039,N_3803,N_3863);
and U4040 (N_4040,N_3935,N_3864);
nand U4041 (N_4041,N_3984,N_3879);
and U4042 (N_4042,N_3816,N_3943);
and U4043 (N_4043,N_3974,N_3909);
nand U4044 (N_4044,N_3930,N_3872);
xnor U4045 (N_4045,N_3938,N_3914);
xor U4046 (N_4046,N_3819,N_3817);
or U4047 (N_4047,N_3849,N_3953);
xnor U4048 (N_4048,N_3894,N_3882);
nand U4049 (N_4049,N_3826,N_3934);
or U4050 (N_4050,N_3976,N_3905);
and U4051 (N_4051,N_3801,N_3981);
nor U4052 (N_4052,N_3977,N_3920);
nand U4053 (N_4053,N_3846,N_3807);
xnor U4054 (N_4054,N_3947,N_3918);
and U4055 (N_4055,N_3966,N_3979);
nor U4056 (N_4056,N_3923,N_3859);
nor U4057 (N_4057,N_3957,N_3911);
xor U4058 (N_4058,N_3867,N_3871);
or U4059 (N_4059,N_3988,N_3845);
or U4060 (N_4060,N_3959,N_3978);
or U4061 (N_4061,N_3936,N_3928);
xnor U4062 (N_4062,N_3949,N_3912);
or U4063 (N_4063,N_3833,N_3870);
nand U4064 (N_4064,N_3873,N_3835);
or U4065 (N_4065,N_3971,N_3960);
nand U4066 (N_4066,N_3929,N_3964);
nand U4067 (N_4067,N_3917,N_3896);
xor U4068 (N_4068,N_3857,N_3840);
or U4069 (N_4069,N_3808,N_3913);
nor U4070 (N_4070,N_3823,N_3856);
nand U4071 (N_4071,N_3921,N_3893);
and U4072 (N_4072,N_3962,N_3908);
xnor U4073 (N_4073,N_3925,N_3973);
xnor U4074 (N_4074,N_3824,N_3812);
nor U4075 (N_4075,N_3860,N_3865);
nand U4076 (N_4076,N_3831,N_3869);
nand U4077 (N_4077,N_3891,N_3991);
nand U4078 (N_4078,N_3827,N_3919);
and U4079 (N_4079,N_3829,N_3898);
or U4080 (N_4080,N_3955,N_3877);
nor U4081 (N_4081,N_3828,N_3916);
xor U4082 (N_4082,N_3885,N_3975);
or U4083 (N_4083,N_3815,N_3851);
or U4084 (N_4084,N_3967,N_3866);
xor U4085 (N_4085,N_3889,N_3800);
xor U4086 (N_4086,N_3890,N_3990);
and U4087 (N_4087,N_3903,N_3852);
nand U4088 (N_4088,N_3822,N_3884);
nand U4089 (N_4089,N_3809,N_3945);
and U4090 (N_4090,N_3922,N_3980);
or U4091 (N_4091,N_3904,N_3995);
nor U4092 (N_4092,N_3880,N_3838);
or U4093 (N_4093,N_3805,N_3969);
nor U4094 (N_4094,N_3900,N_3972);
nand U4095 (N_4095,N_3853,N_3832);
xnor U4096 (N_4096,N_3861,N_3946);
xor U4097 (N_4097,N_3839,N_3899);
or U4098 (N_4098,N_3983,N_3837);
or U4099 (N_4099,N_3841,N_3806);
and U4100 (N_4100,N_3903,N_3971);
and U4101 (N_4101,N_3824,N_3884);
and U4102 (N_4102,N_3914,N_3802);
and U4103 (N_4103,N_3883,N_3930);
or U4104 (N_4104,N_3923,N_3800);
xnor U4105 (N_4105,N_3925,N_3857);
xnor U4106 (N_4106,N_3834,N_3941);
or U4107 (N_4107,N_3842,N_3836);
or U4108 (N_4108,N_3886,N_3854);
nand U4109 (N_4109,N_3812,N_3979);
and U4110 (N_4110,N_3825,N_3804);
or U4111 (N_4111,N_3877,N_3956);
or U4112 (N_4112,N_3894,N_3916);
or U4113 (N_4113,N_3953,N_3869);
and U4114 (N_4114,N_3964,N_3873);
nand U4115 (N_4115,N_3931,N_3980);
xnor U4116 (N_4116,N_3981,N_3873);
and U4117 (N_4117,N_3982,N_3938);
nor U4118 (N_4118,N_3834,N_3966);
nand U4119 (N_4119,N_3820,N_3907);
xnor U4120 (N_4120,N_3867,N_3991);
xnor U4121 (N_4121,N_3876,N_3861);
nor U4122 (N_4122,N_3858,N_3997);
nand U4123 (N_4123,N_3905,N_3834);
or U4124 (N_4124,N_3831,N_3983);
and U4125 (N_4125,N_3964,N_3837);
xor U4126 (N_4126,N_3978,N_3952);
or U4127 (N_4127,N_3843,N_3974);
xor U4128 (N_4128,N_3922,N_3835);
or U4129 (N_4129,N_3861,N_3888);
or U4130 (N_4130,N_3824,N_3911);
nand U4131 (N_4131,N_3825,N_3855);
nor U4132 (N_4132,N_3845,N_3882);
nor U4133 (N_4133,N_3862,N_3847);
nand U4134 (N_4134,N_3830,N_3801);
nand U4135 (N_4135,N_3806,N_3915);
and U4136 (N_4136,N_3830,N_3926);
nand U4137 (N_4137,N_3960,N_3947);
or U4138 (N_4138,N_3817,N_3884);
nor U4139 (N_4139,N_3921,N_3959);
nor U4140 (N_4140,N_3817,N_3997);
xor U4141 (N_4141,N_3995,N_3916);
or U4142 (N_4142,N_3835,N_3973);
nor U4143 (N_4143,N_3883,N_3947);
nand U4144 (N_4144,N_3944,N_3905);
nor U4145 (N_4145,N_3955,N_3829);
nand U4146 (N_4146,N_3903,N_3871);
nor U4147 (N_4147,N_3845,N_3937);
xor U4148 (N_4148,N_3901,N_3985);
or U4149 (N_4149,N_3838,N_3992);
xor U4150 (N_4150,N_3956,N_3943);
nor U4151 (N_4151,N_3966,N_3812);
nor U4152 (N_4152,N_3976,N_3810);
or U4153 (N_4153,N_3852,N_3942);
nor U4154 (N_4154,N_3961,N_3865);
and U4155 (N_4155,N_3975,N_3959);
nor U4156 (N_4156,N_3981,N_3893);
xor U4157 (N_4157,N_3944,N_3930);
xor U4158 (N_4158,N_3934,N_3916);
nand U4159 (N_4159,N_3999,N_3868);
or U4160 (N_4160,N_3851,N_3982);
or U4161 (N_4161,N_3894,N_3998);
xor U4162 (N_4162,N_3872,N_3937);
xor U4163 (N_4163,N_3904,N_3851);
xor U4164 (N_4164,N_3943,N_3967);
nand U4165 (N_4165,N_3833,N_3805);
and U4166 (N_4166,N_3967,N_3858);
nor U4167 (N_4167,N_3926,N_3890);
nand U4168 (N_4168,N_3985,N_3923);
nand U4169 (N_4169,N_3867,N_3926);
xor U4170 (N_4170,N_3832,N_3880);
xor U4171 (N_4171,N_3937,N_3877);
xnor U4172 (N_4172,N_3918,N_3929);
or U4173 (N_4173,N_3969,N_3821);
xnor U4174 (N_4174,N_3808,N_3935);
or U4175 (N_4175,N_3855,N_3927);
nor U4176 (N_4176,N_3998,N_3890);
nand U4177 (N_4177,N_3948,N_3993);
xor U4178 (N_4178,N_3974,N_3953);
and U4179 (N_4179,N_3845,N_3945);
xnor U4180 (N_4180,N_3922,N_3974);
nand U4181 (N_4181,N_3996,N_3894);
or U4182 (N_4182,N_3973,N_3819);
or U4183 (N_4183,N_3994,N_3963);
nor U4184 (N_4184,N_3908,N_3965);
xor U4185 (N_4185,N_3916,N_3856);
xor U4186 (N_4186,N_3856,N_3983);
nor U4187 (N_4187,N_3925,N_3948);
nand U4188 (N_4188,N_3911,N_3860);
nor U4189 (N_4189,N_3898,N_3958);
xnor U4190 (N_4190,N_3853,N_3819);
xor U4191 (N_4191,N_3977,N_3816);
or U4192 (N_4192,N_3922,N_3801);
xnor U4193 (N_4193,N_3874,N_3907);
nand U4194 (N_4194,N_3856,N_3808);
nand U4195 (N_4195,N_3856,N_3817);
and U4196 (N_4196,N_3987,N_3870);
nand U4197 (N_4197,N_3951,N_3896);
nand U4198 (N_4198,N_3912,N_3885);
or U4199 (N_4199,N_3866,N_3812);
xor U4200 (N_4200,N_4058,N_4110);
nor U4201 (N_4201,N_4017,N_4103);
or U4202 (N_4202,N_4127,N_4179);
xnor U4203 (N_4203,N_4027,N_4093);
xnor U4204 (N_4204,N_4186,N_4141);
nor U4205 (N_4205,N_4134,N_4196);
nand U4206 (N_4206,N_4004,N_4096);
and U4207 (N_4207,N_4031,N_4144);
nor U4208 (N_4208,N_4166,N_4094);
xnor U4209 (N_4209,N_4131,N_4097);
or U4210 (N_4210,N_4139,N_4048);
and U4211 (N_4211,N_4156,N_4039);
or U4212 (N_4212,N_4188,N_4162);
and U4213 (N_4213,N_4165,N_4145);
nor U4214 (N_4214,N_4148,N_4065);
xor U4215 (N_4215,N_4088,N_4064);
or U4216 (N_4216,N_4137,N_4069);
nand U4217 (N_4217,N_4068,N_4067);
nand U4218 (N_4218,N_4072,N_4199);
xor U4219 (N_4219,N_4119,N_4149);
nor U4220 (N_4220,N_4182,N_4029);
or U4221 (N_4221,N_4085,N_4078);
xnor U4222 (N_4222,N_4124,N_4183);
xnor U4223 (N_4223,N_4007,N_4089);
nor U4224 (N_4224,N_4087,N_4066);
xor U4225 (N_4225,N_4011,N_4126);
or U4226 (N_4226,N_4147,N_4041);
nand U4227 (N_4227,N_4063,N_4138);
or U4228 (N_4228,N_4121,N_4042);
or U4229 (N_4229,N_4032,N_4151);
nor U4230 (N_4230,N_4043,N_4136);
nand U4231 (N_4231,N_4009,N_4189);
xnor U4232 (N_4232,N_4035,N_4080);
xor U4233 (N_4233,N_4142,N_4173);
nand U4234 (N_4234,N_4023,N_4164);
nor U4235 (N_4235,N_4167,N_4140);
or U4236 (N_4236,N_4014,N_4114);
and U4237 (N_4237,N_4192,N_4033);
xor U4238 (N_4238,N_4160,N_4047);
or U4239 (N_4239,N_4018,N_4163);
xor U4240 (N_4240,N_4062,N_4109);
and U4241 (N_4241,N_4025,N_4132);
and U4242 (N_4242,N_4100,N_4120);
xor U4243 (N_4243,N_4024,N_4115);
nor U4244 (N_4244,N_4090,N_4129);
and U4245 (N_4245,N_4026,N_4150);
or U4246 (N_4246,N_4037,N_4015);
or U4247 (N_4247,N_4020,N_4154);
nor U4248 (N_4248,N_4059,N_4193);
nand U4249 (N_4249,N_4116,N_4102);
or U4250 (N_4250,N_4071,N_4169);
xnor U4251 (N_4251,N_4074,N_4195);
or U4252 (N_4252,N_4181,N_4045);
or U4253 (N_4253,N_4101,N_4191);
or U4254 (N_4254,N_4197,N_4055);
xnor U4255 (N_4255,N_4010,N_4112);
xor U4256 (N_4256,N_4170,N_4174);
and U4257 (N_4257,N_4036,N_4046);
nand U4258 (N_4258,N_4187,N_4133);
and U4259 (N_4259,N_4185,N_4028);
nand U4260 (N_4260,N_4057,N_4083);
or U4261 (N_4261,N_4146,N_4070);
nor U4262 (N_4262,N_4034,N_4177);
or U4263 (N_4263,N_4107,N_4002);
nand U4264 (N_4264,N_4001,N_4184);
xnor U4265 (N_4265,N_4003,N_4051);
and U4266 (N_4266,N_4082,N_4022);
nor U4267 (N_4267,N_4128,N_4111);
nor U4268 (N_4268,N_4198,N_4008);
xor U4269 (N_4269,N_4081,N_4157);
and U4270 (N_4270,N_4076,N_4038);
or U4271 (N_4271,N_4021,N_4168);
or U4272 (N_4272,N_4152,N_4049);
nor U4273 (N_4273,N_4180,N_4105);
and U4274 (N_4274,N_4000,N_4079);
and U4275 (N_4275,N_4158,N_4099);
nand U4276 (N_4276,N_4084,N_4143);
xnor U4277 (N_4277,N_4077,N_4125);
or U4278 (N_4278,N_4104,N_4012);
xnor U4279 (N_4279,N_4175,N_4019);
nand U4280 (N_4280,N_4050,N_4153);
or U4281 (N_4281,N_4060,N_4005);
nor U4282 (N_4282,N_4052,N_4118);
nand U4283 (N_4283,N_4054,N_4098);
and U4284 (N_4284,N_4095,N_4030);
or U4285 (N_4285,N_4123,N_4106);
nor U4286 (N_4286,N_4172,N_4092);
nand U4287 (N_4287,N_4006,N_4061);
or U4288 (N_4288,N_4122,N_4075);
nor U4289 (N_4289,N_4091,N_4056);
and U4290 (N_4290,N_4016,N_4113);
nand U4291 (N_4291,N_4108,N_4053);
xor U4292 (N_4292,N_4117,N_4044);
and U4293 (N_4293,N_4040,N_4135);
nor U4294 (N_4294,N_4161,N_4130);
or U4295 (N_4295,N_4171,N_4155);
and U4296 (N_4296,N_4190,N_4013);
or U4297 (N_4297,N_4086,N_4176);
nor U4298 (N_4298,N_4194,N_4159);
or U4299 (N_4299,N_4178,N_4073);
xor U4300 (N_4300,N_4176,N_4160);
nand U4301 (N_4301,N_4110,N_4019);
or U4302 (N_4302,N_4075,N_4052);
or U4303 (N_4303,N_4143,N_4021);
and U4304 (N_4304,N_4193,N_4006);
nor U4305 (N_4305,N_4045,N_4158);
or U4306 (N_4306,N_4014,N_4035);
and U4307 (N_4307,N_4033,N_4112);
or U4308 (N_4308,N_4161,N_4094);
and U4309 (N_4309,N_4044,N_4063);
or U4310 (N_4310,N_4195,N_4153);
xor U4311 (N_4311,N_4025,N_4103);
nand U4312 (N_4312,N_4043,N_4095);
xnor U4313 (N_4313,N_4015,N_4087);
nand U4314 (N_4314,N_4188,N_4116);
nor U4315 (N_4315,N_4074,N_4112);
nand U4316 (N_4316,N_4185,N_4001);
and U4317 (N_4317,N_4058,N_4108);
and U4318 (N_4318,N_4064,N_4187);
xnor U4319 (N_4319,N_4196,N_4008);
and U4320 (N_4320,N_4037,N_4183);
nand U4321 (N_4321,N_4096,N_4195);
or U4322 (N_4322,N_4176,N_4106);
and U4323 (N_4323,N_4016,N_4051);
nor U4324 (N_4324,N_4019,N_4033);
nand U4325 (N_4325,N_4016,N_4115);
and U4326 (N_4326,N_4169,N_4017);
nand U4327 (N_4327,N_4134,N_4193);
nand U4328 (N_4328,N_4013,N_4149);
or U4329 (N_4329,N_4189,N_4102);
nand U4330 (N_4330,N_4092,N_4023);
or U4331 (N_4331,N_4048,N_4117);
nor U4332 (N_4332,N_4068,N_4008);
or U4333 (N_4333,N_4172,N_4174);
nor U4334 (N_4334,N_4091,N_4133);
and U4335 (N_4335,N_4110,N_4188);
xor U4336 (N_4336,N_4094,N_4035);
nor U4337 (N_4337,N_4056,N_4122);
or U4338 (N_4338,N_4009,N_4139);
and U4339 (N_4339,N_4018,N_4167);
nor U4340 (N_4340,N_4082,N_4128);
xnor U4341 (N_4341,N_4136,N_4065);
or U4342 (N_4342,N_4043,N_4091);
and U4343 (N_4343,N_4032,N_4076);
and U4344 (N_4344,N_4019,N_4015);
nand U4345 (N_4345,N_4074,N_4130);
nand U4346 (N_4346,N_4185,N_4007);
and U4347 (N_4347,N_4061,N_4136);
and U4348 (N_4348,N_4156,N_4196);
nand U4349 (N_4349,N_4109,N_4102);
nor U4350 (N_4350,N_4086,N_4039);
and U4351 (N_4351,N_4048,N_4194);
or U4352 (N_4352,N_4125,N_4123);
xor U4353 (N_4353,N_4117,N_4015);
xor U4354 (N_4354,N_4071,N_4143);
or U4355 (N_4355,N_4065,N_4165);
nor U4356 (N_4356,N_4176,N_4035);
nor U4357 (N_4357,N_4091,N_4164);
nor U4358 (N_4358,N_4064,N_4089);
nand U4359 (N_4359,N_4031,N_4121);
and U4360 (N_4360,N_4044,N_4198);
xnor U4361 (N_4361,N_4167,N_4083);
and U4362 (N_4362,N_4085,N_4196);
xnor U4363 (N_4363,N_4119,N_4126);
nand U4364 (N_4364,N_4006,N_4154);
or U4365 (N_4365,N_4127,N_4056);
xor U4366 (N_4366,N_4173,N_4048);
xor U4367 (N_4367,N_4068,N_4045);
nand U4368 (N_4368,N_4089,N_4004);
or U4369 (N_4369,N_4016,N_4124);
xnor U4370 (N_4370,N_4190,N_4023);
or U4371 (N_4371,N_4128,N_4118);
xnor U4372 (N_4372,N_4112,N_4066);
xor U4373 (N_4373,N_4150,N_4153);
or U4374 (N_4374,N_4154,N_4190);
nand U4375 (N_4375,N_4081,N_4144);
xnor U4376 (N_4376,N_4026,N_4030);
xor U4377 (N_4377,N_4047,N_4082);
nor U4378 (N_4378,N_4030,N_4147);
nor U4379 (N_4379,N_4078,N_4179);
xor U4380 (N_4380,N_4032,N_4094);
or U4381 (N_4381,N_4073,N_4183);
nor U4382 (N_4382,N_4078,N_4150);
and U4383 (N_4383,N_4081,N_4150);
nor U4384 (N_4384,N_4118,N_4085);
and U4385 (N_4385,N_4128,N_4000);
nor U4386 (N_4386,N_4015,N_4028);
nor U4387 (N_4387,N_4104,N_4169);
nor U4388 (N_4388,N_4122,N_4074);
or U4389 (N_4389,N_4115,N_4083);
xnor U4390 (N_4390,N_4128,N_4001);
nor U4391 (N_4391,N_4054,N_4061);
and U4392 (N_4392,N_4075,N_4148);
xnor U4393 (N_4393,N_4130,N_4065);
or U4394 (N_4394,N_4178,N_4063);
nor U4395 (N_4395,N_4086,N_4055);
xnor U4396 (N_4396,N_4009,N_4032);
and U4397 (N_4397,N_4127,N_4175);
nand U4398 (N_4398,N_4173,N_4100);
and U4399 (N_4399,N_4098,N_4190);
xor U4400 (N_4400,N_4330,N_4394);
and U4401 (N_4401,N_4329,N_4347);
and U4402 (N_4402,N_4375,N_4289);
or U4403 (N_4403,N_4351,N_4396);
nor U4404 (N_4404,N_4264,N_4243);
nand U4405 (N_4405,N_4383,N_4292);
nand U4406 (N_4406,N_4341,N_4311);
and U4407 (N_4407,N_4381,N_4284);
or U4408 (N_4408,N_4236,N_4260);
xor U4409 (N_4409,N_4258,N_4397);
xnor U4410 (N_4410,N_4328,N_4234);
or U4411 (N_4411,N_4248,N_4353);
nor U4412 (N_4412,N_4392,N_4358);
nand U4413 (N_4413,N_4269,N_4232);
or U4414 (N_4414,N_4220,N_4349);
xnor U4415 (N_4415,N_4245,N_4265);
or U4416 (N_4416,N_4348,N_4251);
nand U4417 (N_4417,N_4281,N_4227);
xnor U4418 (N_4418,N_4354,N_4224);
xor U4419 (N_4419,N_4223,N_4386);
nand U4420 (N_4420,N_4308,N_4313);
or U4421 (N_4421,N_4202,N_4395);
or U4422 (N_4422,N_4315,N_4293);
nand U4423 (N_4423,N_4212,N_4334);
and U4424 (N_4424,N_4365,N_4273);
and U4425 (N_4425,N_4327,N_4255);
nand U4426 (N_4426,N_4305,N_4237);
xnor U4427 (N_4427,N_4343,N_4373);
xnor U4428 (N_4428,N_4244,N_4302);
or U4429 (N_4429,N_4210,N_4299);
xnor U4430 (N_4430,N_4340,N_4211);
nor U4431 (N_4431,N_4221,N_4204);
and U4432 (N_4432,N_4275,N_4217);
nand U4433 (N_4433,N_4271,N_4320);
xnor U4434 (N_4434,N_4377,N_4356);
and U4435 (N_4435,N_4268,N_4256);
xnor U4436 (N_4436,N_4254,N_4231);
xnor U4437 (N_4437,N_4247,N_4378);
and U4438 (N_4438,N_4310,N_4279);
nand U4439 (N_4439,N_4372,N_4208);
or U4440 (N_4440,N_4357,N_4287);
and U4441 (N_4441,N_4298,N_4309);
xnor U4442 (N_4442,N_4282,N_4389);
xor U4443 (N_4443,N_4288,N_4295);
nor U4444 (N_4444,N_4263,N_4338);
and U4445 (N_4445,N_4376,N_4222);
and U4446 (N_4446,N_4316,N_4304);
and U4447 (N_4447,N_4359,N_4344);
or U4448 (N_4448,N_4242,N_4390);
or U4449 (N_4449,N_4207,N_4214);
xnor U4450 (N_4450,N_4339,N_4352);
and U4451 (N_4451,N_4253,N_4215);
nor U4452 (N_4452,N_4333,N_4262);
nor U4453 (N_4453,N_4350,N_4380);
nand U4454 (N_4454,N_4206,N_4259);
and U4455 (N_4455,N_4387,N_4246);
nor U4456 (N_4456,N_4306,N_4361);
and U4457 (N_4457,N_4364,N_4280);
nand U4458 (N_4458,N_4388,N_4294);
or U4459 (N_4459,N_4297,N_4270);
and U4460 (N_4460,N_4382,N_4216);
and U4461 (N_4461,N_4307,N_4285);
or U4462 (N_4462,N_4209,N_4355);
or U4463 (N_4463,N_4398,N_4366);
xor U4464 (N_4464,N_4301,N_4367);
or U4465 (N_4465,N_4391,N_4290);
and U4466 (N_4466,N_4213,N_4321);
xor U4467 (N_4467,N_4267,N_4374);
xor U4468 (N_4468,N_4399,N_4252);
xnor U4469 (N_4469,N_4261,N_4379);
nand U4470 (N_4470,N_4337,N_4368);
or U4471 (N_4471,N_4226,N_4230);
xnor U4472 (N_4472,N_4362,N_4276);
nor U4473 (N_4473,N_4312,N_4371);
and U4474 (N_4474,N_4239,N_4238);
nor U4475 (N_4475,N_4385,N_4323);
and U4476 (N_4476,N_4336,N_4228);
nand U4477 (N_4477,N_4240,N_4277);
nand U4478 (N_4478,N_4300,N_4286);
or U4479 (N_4479,N_4283,N_4278);
xor U4480 (N_4480,N_4331,N_4219);
and U4481 (N_4481,N_4393,N_4314);
and U4482 (N_4482,N_4225,N_4235);
or U4483 (N_4483,N_4274,N_4325);
nor U4484 (N_4484,N_4241,N_4324);
or U4485 (N_4485,N_4266,N_4384);
xnor U4486 (N_4486,N_4257,N_4370);
nand U4487 (N_4487,N_4345,N_4332);
nor U4488 (N_4488,N_4360,N_4346);
xor U4489 (N_4489,N_4205,N_4326);
xnor U4490 (N_4490,N_4318,N_4272);
xor U4491 (N_4491,N_4303,N_4335);
or U4492 (N_4492,N_4203,N_4342);
and U4493 (N_4493,N_4250,N_4229);
or U4494 (N_4494,N_4201,N_4200);
xor U4495 (N_4495,N_4218,N_4317);
nor U4496 (N_4496,N_4369,N_4363);
or U4497 (N_4497,N_4322,N_4233);
xor U4498 (N_4498,N_4319,N_4296);
nor U4499 (N_4499,N_4249,N_4291);
xnor U4500 (N_4500,N_4270,N_4329);
or U4501 (N_4501,N_4374,N_4286);
nand U4502 (N_4502,N_4284,N_4203);
nor U4503 (N_4503,N_4250,N_4222);
xnor U4504 (N_4504,N_4257,N_4251);
and U4505 (N_4505,N_4317,N_4333);
and U4506 (N_4506,N_4331,N_4241);
nor U4507 (N_4507,N_4275,N_4353);
nor U4508 (N_4508,N_4375,N_4225);
xor U4509 (N_4509,N_4288,N_4323);
xor U4510 (N_4510,N_4318,N_4391);
and U4511 (N_4511,N_4394,N_4368);
xnor U4512 (N_4512,N_4258,N_4393);
nand U4513 (N_4513,N_4229,N_4294);
and U4514 (N_4514,N_4395,N_4356);
nand U4515 (N_4515,N_4346,N_4318);
nor U4516 (N_4516,N_4205,N_4214);
nand U4517 (N_4517,N_4310,N_4204);
nand U4518 (N_4518,N_4234,N_4308);
or U4519 (N_4519,N_4239,N_4377);
or U4520 (N_4520,N_4234,N_4357);
or U4521 (N_4521,N_4332,N_4341);
and U4522 (N_4522,N_4368,N_4280);
and U4523 (N_4523,N_4348,N_4374);
or U4524 (N_4524,N_4275,N_4227);
nand U4525 (N_4525,N_4330,N_4227);
xor U4526 (N_4526,N_4347,N_4233);
xnor U4527 (N_4527,N_4235,N_4322);
xnor U4528 (N_4528,N_4219,N_4276);
and U4529 (N_4529,N_4345,N_4324);
or U4530 (N_4530,N_4392,N_4310);
or U4531 (N_4531,N_4246,N_4281);
and U4532 (N_4532,N_4241,N_4337);
or U4533 (N_4533,N_4256,N_4318);
nor U4534 (N_4534,N_4366,N_4327);
and U4535 (N_4535,N_4376,N_4342);
and U4536 (N_4536,N_4375,N_4238);
xnor U4537 (N_4537,N_4288,N_4279);
or U4538 (N_4538,N_4210,N_4288);
or U4539 (N_4539,N_4274,N_4284);
and U4540 (N_4540,N_4230,N_4209);
nor U4541 (N_4541,N_4317,N_4342);
nand U4542 (N_4542,N_4317,N_4239);
xnor U4543 (N_4543,N_4327,N_4245);
or U4544 (N_4544,N_4200,N_4282);
nor U4545 (N_4545,N_4375,N_4348);
and U4546 (N_4546,N_4383,N_4296);
nor U4547 (N_4547,N_4301,N_4260);
nand U4548 (N_4548,N_4329,N_4385);
or U4549 (N_4549,N_4300,N_4296);
nand U4550 (N_4550,N_4211,N_4301);
or U4551 (N_4551,N_4242,N_4298);
nor U4552 (N_4552,N_4348,N_4309);
nand U4553 (N_4553,N_4397,N_4267);
xor U4554 (N_4554,N_4254,N_4252);
nand U4555 (N_4555,N_4398,N_4376);
and U4556 (N_4556,N_4243,N_4354);
nor U4557 (N_4557,N_4351,N_4273);
nand U4558 (N_4558,N_4315,N_4305);
xor U4559 (N_4559,N_4233,N_4222);
nand U4560 (N_4560,N_4291,N_4207);
or U4561 (N_4561,N_4253,N_4384);
nor U4562 (N_4562,N_4316,N_4378);
nand U4563 (N_4563,N_4234,N_4394);
nand U4564 (N_4564,N_4240,N_4217);
xor U4565 (N_4565,N_4201,N_4320);
nor U4566 (N_4566,N_4310,N_4272);
nor U4567 (N_4567,N_4276,N_4251);
xnor U4568 (N_4568,N_4303,N_4289);
or U4569 (N_4569,N_4266,N_4393);
nand U4570 (N_4570,N_4223,N_4289);
xnor U4571 (N_4571,N_4296,N_4370);
nand U4572 (N_4572,N_4214,N_4377);
or U4573 (N_4573,N_4326,N_4262);
nor U4574 (N_4574,N_4386,N_4317);
nor U4575 (N_4575,N_4252,N_4209);
nand U4576 (N_4576,N_4345,N_4278);
or U4577 (N_4577,N_4280,N_4305);
nor U4578 (N_4578,N_4253,N_4210);
nand U4579 (N_4579,N_4260,N_4360);
and U4580 (N_4580,N_4254,N_4282);
or U4581 (N_4581,N_4326,N_4255);
nor U4582 (N_4582,N_4309,N_4356);
nor U4583 (N_4583,N_4243,N_4294);
and U4584 (N_4584,N_4258,N_4291);
or U4585 (N_4585,N_4321,N_4386);
and U4586 (N_4586,N_4261,N_4340);
and U4587 (N_4587,N_4329,N_4292);
xnor U4588 (N_4588,N_4231,N_4394);
and U4589 (N_4589,N_4377,N_4326);
and U4590 (N_4590,N_4385,N_4306);
xnor U4591 (N_4591,N_4313,N_4334);
nor U4592 (N_4592,N_4260,N_4314);
and U4593 (N_4593,N_4316,N_4214);
and U4594 (N_4594,N_4278,N_4297);
nand U4595 (N_4595,N_4293,N_4365);
nand U4596 (N_4596,N_4309,N_4368);
and U4597 (N_4597,N_4289,N_4313);
and U4598 (N_4598,N_4325,N_4212);
nor U4599 (N_4599,N_4328,N_4364);
or U4600 (N_4600,N_4553,N_4479);
nand U4601 (N_4601,N_4575,N_4513);
nor U4602 (N_4602,N_4542,N_4555);
xnor U4603 (N_4603,N_4449,N_4533);
xor U4604 (N_4604,N_4564,N_4403);
nand U4605 (N_4605,N_4476,N_4493);
nand U4606 (N_4606,N_4524,N_4537);
or U4607 (N_4607,N_4576,N_4484);
or U4608 (N_4608,N_4486,N_4574);
xnor U4609 (N_4609,N_4531,N_4535);
nand U4610 (N_4610,N_4458,N_4468);
xnor U4611 (N_4611,N_4415,N_4587);
nor U4612 (N_4612,N_4578,N_4507);
xor U4613 (N_4613,N_4448,N_4580);
nor U4614 (N_4614,N_4552,N_4459);
nor U4615 (N_4615,N_4536,N_4501);
nor U4616 (N_4616,N_4592,N_4579);
nand U4617 (N_4617,N_4433,N_4447);
nor U4618 (N_4618,N_4420,N_4526);
xor U4619 (N_4619,N_4521,N_4510);
xor U4620 (N_4620,N_4401,N_4566);
nor U4621 (N_4621,N_4584,N_4583);
nor U4622 (N_4622,N_4556,N_4503);
or U4623 (N_4623,N_4421,N_4512);
and U4624 (N_4624,N_4546,N_4416);
or U4625 (N_4625,N_4430,N_4487);
xor U4626 (N_4626,N_4500,N_4464);
and U4627 (N_4627,N_4425,N_4434);
nand U4628 (N_4628,N_4429,N_4432);
nand U4629 (N_4629,N_4582,N_4499);
nand U4630 (N_4630,N_4558,N_4515);
and U4631 (N_4631,N_4411,N_4427);
or U4632 (N_4632,N_4522,N_4494);
or U4633 (N_4633,N_4469,N_4591);
nand U4634 (N_4634,N_4561,N_4593);
nor U4635 (N_4635,N_4492,N_4439);
nand U4636 (N_4636,N_4454,N_4456);
xor U4637 (N_4637,N_4490,N_4473);
xor U4638 (N_4638,N_4443,N_4481);
nor U4639 (N_4639,N_4423,N_4463);
or U4640 (N_4640,N_4409,N_4498);
nand U4641 (N_4641,N_4400,N_4404);
nor U4642 (N_4642,N_4485,N_4445);
nand U4643 (N_4643,N_4441,N_4457);
nand U4644 (N_4644,N_4569,N_4532);
and U4645 (N_4645,N_4589,N_4428);
nand U4646 (N_4646,N_4444,N_4568);
and U4647 (N_4647,N_4563,N_4547);
or U4648 (N_4648,N_4470,N_4545);
or U4649 (N_4649,N_4525,N_4517);
or U4650 (N_4650,N_4405,N_4406);
or U4651 (N_4651,N_4534,N_4529);
and U4652 (N_4652,N_4482,N_4418);
or U4653 (N_4653,N_4549,N_4557);
or U4654 (N_4654,N_4573,N_4502);
and U4655 (N_4655,N_4410,N_4407);
xnor U4656 (N_4656,N_4431,N_4570);
or U4657 (N_4657,N_4596,N_4541);
nor U4658 (N_4658,N_4472,N_4426);
nor U4659 (N_4659,N_4554,N_4504);
nand U4660 (N_4660,N_4523,N_4436);
xnor U4661 (N_4661,N_4539,N_4412);
or U4662 (N_4662,N_4478,N_4413);
or U4663 (N_4663,N_4508,N_4594);
or U4664 (N_4664,N_4419,N_4424);
nor U4665 (N_4665,N_4506,N_4550);
nor U4666 (N_4666,N_4471,N_4437);
and U4667 (N_4667,N_4442,N_4511);
nand U4668 (N_4668,N_4586,N_4450);
nand U4669 (N_4669,N_4475,N_4514);
xor U4670 (N_4670,N_4598,N_4435);
xnor U4671 (N_4671,N_4519,N_4571);
nand U4672 (N_4672,N_4474,N_4477);
nor U4673 (N_4673,N_4581,N_4453);
nor U4674 (N_4674,N_4543,N_4562);
nand U4675 (N_4675,N_4527,N_4544);
or U4676 (N_4676,N_4572,N_4483);
or U4677 (N_4677,N_4565,N_4597);
nand U4678 (N_4678,N_4461,N_4496);
or U4679 (N_4679,N_4438,N_4462);
xnor U4680 (N_4680,N_4455,N_4588);
or U4681 (N_4681,N_4567,N_4414);
nor U4682 (N_4682,N_4599,N_4466);
xor U4683 (N_4683,N_4590,N_4538);
xnor U4684 (N_4684,N_4467,N_4460);
and U4685 (N_4685,N_4402,N_4509);
and U4686 (N_4686,N_4530,N_4548);
or U4687 (N_4687,N_4465,N_4528);
and U4688 (N_4688,N_4497,N_4559);
and U4689 (N_4689,N_4540,N_4505);
nor U4690 (N_4690,N_4495,N_4417);
nand U4691 (N_4691,N_4489,N_4577);
and U4692 (N_4692,N_4585,N_4491);
or U4693 (N_4693,N_4520,N_4422);
or U4694 (N_4694,N_4446,N_4560);
xor U4695 (N_4695,N_4488,N_4452);
xor U4696 (N_4696,N_4516,N_4551);
and U4697 (N_4697,N_4440,N_4408);
or U4698 (N_4698,N_4451,N_4480);
nor U4699 (N_4699,N_4518,N_4595);
nand U4700 (N_4700,N_4441,N_4518);
or U4701 (N_4701,N_4541,N_4576);
or U4702 (N_4702,N_4505,N_4454);
nand U4703 (N_4703,N_4463,N_4411);
nor U4704 (N_4704,N_4401,N_4596);
or U4705 (N_4705,N_4551,N_4448);
xnor U4706 (N_4706,N_4461,N_4444);
nand U4707 (N_4707,N_4548,N_4420);
or U4708 (N_4708,N_4571,N_4548);
xnor U4709 (N_4709,N_4464,N_4476);
and U4710 (N_4710,N_4582,N_4502);
and U4711 (N_4711,N_4481,N_4433);
nor U4712 (N_4712,N_4524,N_4528);
xnor U4713 (N_4713,N_4482,N_4425);
xor U4714 (N_4714,N_4559,N_4410);
xnor U4715 (N_4715,N_4508,N_4411);
nor U4716 (N_4716,N_4445,N_4539);
xnor U4717 (N_4717,N_4573,N_4474);
xor U4718 (N_4718,N_4435,N_4568);
or U4719 (N_4719,N_4521,N_4551);
nand U4720 (N_4720,N_4534,N_4542);
and U4721 (N_4721,N_4480,N_4514);
and U4722 (N_4722,N_4420,N_4502);
and U4723 (N_4723,N_4571,N_4488);
nor U4724 (N_4724,N_4541,N_4579);
and U4725 (N_4725,N_4548,N_4453);
nand U4726 (N_4726,N_4476,N_4505);
and U4727 (N_4727,N_4507,N_4526);
and U4728 (N_4728,N_4454,N_4591);
nor U4729 (N_4729,N_4541,N_4559);
nor U4730 (N_4730,N_4519,N_4561);
or U4731 (N_4731,N_4530,N_4524);
xor U4732 (N_4732,N_4423,N_4451);
or U4733 (N_4733,N_4472,N_4573);
nor U4734 (N_4734,N_4547,N_4576);
or U4735 (N_4735,N_4472,N_4513);
and U4736 (N_4736,N_4480,N_4590);
xnor U4737 (N_4737,N_4435,N_4402);
xor U4738 (N_4738,N_4556,N_4438);
or U4739 (N_4739,N_4451,N_4588);
xor U4740 (N_4740,N_4452,N_4413);
and U4741 (N_4741,N_4471,N_4497);
or U4742 (N_4742,N_4442,N_4462);
nand U4743 (N_4743,N_4425,N_4562);
nand U4744 (N_4744,N_4522,N_4476);
and U4745 (N_4745,N_4427,N_4436);
or U4746 (N_4746,N_4568,N_4460);
xor U4747 (N_4747,N_4511,N_4565);
and U4748 (N_4748,N_4483,N_4570);
nand U4749 (N_4749,N_4511,N_4559);
or U4750 (N_4750,N_4411,N_4477);
or U4751 (N_4751,N_4590,N_4553);
nor U4752 (N_4752,N_4429,N_4430);
and U4753 (N_4753,N_4503,N_4404);
and U4754 (N_4754,N_4534,N_4585);
nor U4755 (N_4755,N_4567,N_4550);
nand U4756 (N_4756,N_4466,N_4439);
and U4757 (N_4757,N_4400,N_4449);
nand U4758 (N_4758,N_4515,N_4470);
xor U4759 (N_4759,N_4481,N_4590);
or U4760 (N_4760,N_4595,N_4596);
and U4761 (N_4761,N_4521,N_4483);
xor U4762 (N_4762,N_4565,N_4560);
and U4763 (N_4763,N_4548,N_4559);
nor U4764 (N_4764,N_4412,N_4501);
nand U4765 (N_4765,N_4553,N_4533);
nand U4766 (N_4766,N_4411,N_4437);
nand U4767 (N_4767,N_4545,N_4583);
or U4768 (N_4768,N_4500,N_4466);
nor U4769 (N_4769,N_4509,N_4455);
nor U4770 (N_4770,N_4534,N_4484);
nand U4771 (N_4771,N_4508,N_4553);
or U4772 (N_4772,N_4526,N_4403);
and U4773 (N_4773,N_4536,N_4438);
and U4774 (N_4774,N_4504,N_4457);
xnor U4775 (N_4775,N_4412,N_4483);
or U4776 (N_4776,N_4533,N_4583);
nor U4777 (N_4777,N_4541,N_4457);
xnor U4778 (N_4778,N_4430,N_4451);
xor U4779 (N_4779,N_4412,N_4500);
and U4780 (N_4780,N_4526,N_4581);
and U4781 (N_4781,N_4463,N_4551);
or U4782 (N_4782,N_4502,N_4564);
xnor U4783 (N_4783,N_4593,N_4481);
xor U4784 (N_4784,N_4473,N_4546);
nand U4785 (N_4785,N_4589,N_4479);
and U4786 (N_4786,N_4549,N_4540);
nand U4787 (N_4787,N_4559,N_4596);
nor U4788 (N_4788,N_4403,N_4546);
nand U4789 (N_4789,N_4423,N_4434);
or U4790 (N_4790,N_4575,N_4598);
nand U4791 (N_4791,N_4404,N_4569);
nand U4792 (N_4792,N_4588,N_4447);
xnor U4793 (N_4793,N_4439,N_4427);
or U4794 (N_4794,N_4499,N_4583);
nor U4795 (N_4795,N_4517,N_4403);
and U4796 (N_4796,N_4506,N_4464);
xnor U4797 (N_4797,N_4498,N_4501);
and U4798 (N_4798,N_4560,N_4407);
nor U4799 (N_4799,N_4596,N_4419);
or U4800 (N_4800,N_4703,N_4764);
nand U4801 (N_4801,N_4604,N_4719);
nor U4802 (N_4802,N_4619,N_4665);
or U4803 (N_4803,N_4605,N_4661);
nor U4804 (N_4804,N_4628,N_4639);
xor U4805 (N_4805,N_4797,N_4648);
xor U4806 (N_4806,N_4730,N_4629);
nand U4807 (N_4807,N_4622,N_4603);
xor U4808 (N_4808,N_4744,N_4708);
nor U4809 (N_4809,N_4717,N_4620);
xnor U4810 (N_4810,N_4615,N_4611);
or U4811 (N_4811,N_4613,N_4711);
nor U4812 (N_4812,N_4642,N_4669);
nor U4813 (N_4813,N_4728,N_4671);
nor U4814 (N_4814,N_4678,N_4631);
and U4815 (N_4815,N_4656,N_4636);
nor U4816 (N_4816,N_4659,N_4610);
or U4817 (N_4817,N_4601,N_4732);
nor U4818 (N_4818,N_4767,N_4640);
or U4819 (N_4819,N_4667,N_4758);
or U4820 (N_4820,N_4684,N_4726);
xnor U4821 (N_4821,N_4761,N_4743);
nor U4822 (N_4822,N_4774,N_4664);
and U4823 (N_4823,N_4710,N_4783);
and U4824 (N_4824,N_4676,N_4614);
and U4825 (N_4825,N_4692,N_4793);
nor U4826 (N_4826,N_4714,N_4704);
or U4827 (N_4827,N_4696,N_4653);
nand U4828 (N_4828,N_4736,N_4715);
and U4829 (N_4829,N_4757,N_4759);
nand U4830 (N_4830,N_4722,N_4779);
xnor U4831 (N_4831,N_4649,N_4763);
nand U4832 (N_4832,N_4673,N_4784);
or U4833 (N_4833,N_4788,N_4695);
or U4834 (N_4834,N_4750,N_4637);
nand U4835 (N_4835,N_4655,N_4638);
nand U4836 (N_4836,N_4632,N_4724);
or U4837 (N_4837,N_4652,N_4794);
and U4838 (N_4838,N_4712,N_4626);
nor U4839 (N_4839,N_4699,N_4738);
and U4840 (N_4840,N_4641,N_4694);
or U4841 (N_4841,N_4618,N_4729);
nand U4842 (N_4842,N_4721,N_4624);
nand U4843 (N_4843,N_4630,N_4787);
or U4844 (N_4844,N_4709,N_4700);
nand U4845 (N_4845,N_4775,N_4792);
nor U4846 (N_4846,N_4755,N_4677);
and U4847 (N_4847,N_4682,N_4791);
or U4848 (N_4848,N_4731,N_4737);
and U4849 (N_4849,N_4786,N_4658);
or U4850 (N_4850,N_4644,N_4675);
or U4851 (N_4851,N_4609,N_4606);
nand U4852 (N_4852,N_4685,N_4718);
xor U4853 (N_4853,N_4735,N_4600);
or U4854 (N_4854,N_4725,N_4698);
and U4855 (N_4855,N_4691,N_4681);
or U4856 (N_4856,N_4765,N_4771);
or U4857 (N_4857,N_4789,N_4634);
and U4858 (N_4858,N_4660,N_4742);
and U4859 (N_4859,N_4790,N_4690);
nor U4860 (N_4860,N_4727,N_4772);
and U4861 (N_4861,N_4666,N_4777);
and U4862 (N_4862,N_4706,N_4720);
xnor U4863 (N_4863,N_4657,N_4770);
and U4864 (N_4864,N_4668,N_4650);
or U4865 (N_4865,N_4608,N_4780);
or U4866 (N_4866,N_4689,N_4693);
nand U4867 (N_4867,N_4651,N_4623);
or U4868 (N_4868,N_4785,N_4746);
xnor U4869 (N_4869,N_4745,N_4798);
nor U4870 (N_4870,N_4633,N_4716);
nor U4871 (N_4871,N_4756,N_4751);
nand U4872 (N_4872,N_4672,N_4662);
and U4873 (N_4873,N_4663,N_4747);
nand U4874 (N_4874,N_4625,N_4697);
and U4875 (N_4875,N_4748,N_4768);
or U4876 (N_4876,N_4760,N_4753);
nand U4877 (N_4877,N_4733,N_4707);
and U4878 (N_4878,N_4713,N_4687);
nor U4879 (N_4879,N_4602,N_4635);
xnor U4880 (N_4880,N_4754,N_4766);
nand U4881 (N_4881,N_4647,N_4702);
or U4882 (N_4882,N_4739,N_4627);
nand U4883 (N_4883,N_4607,N_4616);
or U4884 (N_4884,N_4781,N_4769);
or U4885 (N_4885,N_4643,N_4645);
or U4886 (N_4886,N_4778,N_4680);
and U4887 (N_4887,N_4782,N_4674);
nand U4888 (N_4888,N_4621,N_4762);
or U4889 (N_4889,N_4670,N_4795);
xnor U4890 (N_4890,N_4646,N_4799);
nor U4891 (N_4891,N_4749,N_4723);
xor U4892 (N_4892,N_4741,N_4705);
nor U4893 (N_4893,N_4686,N_4688);
nor U4894 (N_4894,N_4654,N_4752);
nand U4895 (N_4895,N_4683,N_4612);
xnor U4896 (N_4896,N_4773,N_4734);
nand U4897 (N_4897,N_4740,N_4679);
xnor U4898 (N_4898,N_4776,N_4796);
nor U4899 (N_4899,N_4617,N_4701);
xor U4900 (N_4900,N_4616,N_4650);
and U4901 (N_4901,N_4647,N_4768);
nor U4902 (N_4902,N_4792,N_4664);
xnor U4903 (N_4903,N_4604,N_4720);
nor U4904 (N_4904,N_4728,N_4732);
xnor U4905 (N_4905,N_4626,N_4631);
nand U4906 (N_4906,N_4684,N_4689);
nand U4907 (N_4907,N_4649,N_4731);
or U4908 (N_4908,N_4670,N_4662);
xor U4909 (N_4909,N_4726,N_4670);
nand U4910 (N_4910,N_4776,N_4637);
nor U4911 (N_4911,N_4675,N_4626);
and U4912 (N_4912,N_4635,N_4775);
xor U4913 (N_4913,N_4776,N_4765);
and U4914 (N_4914,N_4700,N_4627);
nand U4915 (N_4915,N_4714,N_4790);
nand U4916 (N_4916,N_4681,N_4706);
nor U4917 (N_4917,N_4774,N_4700);
or U4918 (N_4918,N_4608,N_4615);
xor U4919 (N_4919,N_4687,N_4788);
and U4920 (N_4920,N_4701,N_4716);
or U4921 (N_4921,N_4659,N_4654);
or U4922 (N_4922,N_4604,N_4648);
nand U4923 (N_4923,N_4622,N_4772);
xor U4924 (N_4924,N_4729,N_4607);
or U4925 (N_4925,N_4713,N_4712);
xnor U4926 (N_4926,N_4622,N_4604);
nand U4927 (N_4927,N_4657,N_4621);
and U4928 (N_4928,N_4702,N_4785);
xnor U4929 (N_4929,N_4689,N_4630);
xnor U4930 (N_4930,N_4784,N_4663);
nor U4931 (N_4931,N_4616,N_4711);
xor U4932 (N_4932,N_4796,N_4764);
or U4933 (N_4933,N_4710,N_4607);
nor U4934 (N_4934,N_4704,N_4692);
nand U4935 (N_4935,N_4694,N_4678);
or U4936 (N_4936,N_4600,N_4652);
or U4937 (N_4937,N_4645,N_4612);
or U4938 (N_4938,N_4683,N_4664);
xnor U4939 (N_4939,N_4713,N_4770);
or U4940 (N_4940,N_4739,N_4665);
or U4941 (N_4941,N_4654,N_4604);
nor U4942 (N_4942,N_4645,N_4716);
and U4943 (N_4943,N_4667,N_4783);
nand U4944 (N_4944,N_4792,N_4611);
and U4945 (N_4945,N_4797,N_4728);
or U4946 (N_4946,N_4636,N_4685);
or U4947 (N_4947,N_4762,N_4613);
xor U4948 (N_4948,N_4687,N_4751);
xnor U4949 (N_4949,N_4632,N_4677);
nand U4950 (N_4950,N_4788,N_4670);
and U4951 (N_4951,N_4757,N_4641);
nor U4952 (N_4952,N_4653,N_4628);
or U4953 (N_4953,N_4798,N_4728);
or U4954 (N_4954,N_4725,N_4640);
or U4955 (N_4955,N_4729,N_4705);
nor U4956 (N_4956,N_4635,N_4695);
or U4957 (N_4957,N_4601,N_4724);
and U4958 (N_4958,N_4788,N_4677);
nand U4959 (N_4959,N_4729,N_4629);
nand U4960 (N_4960,N_4700,N_4619);
nor U4961 (N_4961,N_4702,N_4725);
nor U4962 (N_4962,N_4618,N_4779);
nand U4963 (N_4963,N_4612,N_4662);
and U4964 (N_4964,N_4655,N_4775);
nor U4965 (N_4965,N_4735,N_4713);
and U4966 (N_4966,N_4793,N_4636);
nor U4967 (N_4967,N_4683,N_4672);
and U4968 (N_4968,N_4600,N_4678);
and U4969 (N_4969,N_4773,N_4641);
nor U4970 (N_4970,N_4678,N_4614);
nor U4971 (N_4971,N_4621,N_4770);
nor U4972 (N_4972,N_4752,N_4641);
or U4973 (N_4973,N_4727,N_4669);
nor U4974 (N_4974,N_4775,N_4621);
nand U4975 (N_4975,N_4696,N_4607);
nor U4976 (N_4976,N_4739,N_4793);
and U4977 (N_4977,N_4711,N_4676);
xor U4978 (N_4978,N_4662,N_4642);
and U4979 (N_4979,N_4709,N_4658);
xnor U4980 (N_4980,N_4643,N_4617);
xor U4981 (N_4981,N_4772,N_4643);
or U4982 (N_4982,N_4736,N_4616);
or U4983 (N_4983,N_4663,N_4666);
xnor U4984 (N_4984,N_4627,N_4691);
nand U4985 (N_4985,N_4619,N_4608);
xor U4986 (N_4986,N_4745,N_4692);
or U4987 (N_4987,N_4708,N_4667);
xor U4988 (N_4988,N_4787,N_4623);
and U4989 (N_4989,N_4786,N_4634);
nor U4990 (N_4990,N_4722,N_4784);
nor U4991 (N_4991,N_4650,N_4700);
nor U4992 (N_4992,N_4768,N_4744);
xor U4993 (N_4993,N_4649,N_4715);
nor U4994 (N_4994,N_4652,N_4717);
nor U4995 (N_4995,N_4724,N_4696);
nand U4996 (N_4996,N_4732,N_4765);
or U4997 (N_4997,N_4612,N_4685);
and U4998 (N_4998,N_4690,N_4741);
nor U4999 (N_4999,N_4640,N_4728);
nand U5000 (N_5000,N_4916,N_4847);
and U5001 (N_5001,N_4911,N_4863);
and U5002 (N_5002,N_4907,N_4944);
or U5003 (N_5003,N_4921,N_4992);
nor U5004 (N_5004,N_4945,N_4958);
xor U5005 (N_5005,N_4895,N_4966);
nor U5006 (N_5006,N_4811,N_4902);
nand U5007 (N_5007,N_4814,N_4901);
and U5008 (N_5008,N_4951,N_4939);
nand U5009 (N_5009,N_4934,N_4953);
nand U5010 (N_5010,N_4829,N_4931);
nor U5011 (N_5011,N_4917,N_4969);
nand U5012 (N_5012,N_4869,N_4873);
xnor U5013 (N_5013,N_4808,N_4820);
and U5014 (N_5014,N_4982,N_4899);
nor U5015 (N_5015,N_4920,N_4856);
nand U5016 (N_5016,N_4868,N_4844);
nor U5017 (N_5017,N_4974,N_4976);
or U5018 (N_5018,N_4827,N_4851);
nor U5019 (N_5019,N_4849,N_4874);
nor U5020 (N_5020,N_4935,N_4922);
xnor U5021 (N_5021,N_4812,N_4967);
nand U5022 (N_5022,N_4908,N_4854);
xnor U5023 (N_5023,N_4978,N_4848);
nand U5024 (N_5024,N_4815,N_4893);
or U5025 (N_5025,N_4857,N_4823);
xnor U5026 (N_5026,N_4800,N_4970);
xor U5027 (N_5027,N_4865,N_4889);
nor U5028 (N_5028,N_4906,N_4980);
nor U5029 (N_5029,N_4930,N_4880);
xnor U5030 (N_5030,N_4938,N_4825);
and U5031 (N_5031,N_4943,N_4954);
nor U5032 (N_5032,N_4843,N_4955);
nand U5033 (N_5033,N_4990,N_4948);
nand U5034 (N_5034,N_4875,N_4833);
or U5035 (N_5035,N_4836,N_4983);
nand U5036 (N_5036,N_4923,N_4932);
nor U5037 (N_5037,N_4961,N_4821);
xor U5038 (N_5038,N_4971,N_4898);
and U5039 (N_5039,N_4852,N_4828);
or U5040 (N_5040,N_4834,N_4929);
and U5041 (N_5041,N_4846,N_4817);
nand U5042 (N_5042,N_4919,N_4926);
and U5043 (N_5043,N_4986,N_4877);
or U5044 (N_5044,N_4896,N_4999);
and U5045 (N_5045,N_4981,N_4830);
nand U5046 (N_5046,N_4946,N_4872);
or U5047 (N_5047,N_4816,N_4909);
nand U5048 (N_5048,N_4855,N_4995);
and U5049 (N_5049,N_4883,N_4933);
xnor U5050 (N_5050,N_4915,N_4850);
nor U5051 (N_5051,N_4910,N_4997);
or U5052 (N_5052,N_4949,N_4960);
and U5053 (N_5053,N_4904,N_4888);
or U5054 (N_5054,N_4905,N_4801);
and U5055 (N_5055,N_4831,N_4975);
xnor U5056 (N_5056,N_4842,N_4818);
and U5057 (N_5057,N_4835,N_4963);
xor U5058 (N_5058,N_4839,N_4998);
or U5059 (N_5059,N_4804,N_4845);
nor U5060 (N_5060,N_4840,N_4870);
nor U5061 (N_5061,N_4903,N_4973);
xor U5062 (N_5062,N_4913,N_4957);
xnor U5063 (N_5063,N_4996,N_4994);
nor U5064 (N_5064,N_4802,N_4887);
nor U5065 (N_5065,N_4882,N_4824);
and U5066 (N_5066,N_4853,N_4928);
and U5067 (N_5067,N_4891,N_4940);
or U5068 (N_5068,N_4988,N_4984);
xor U5069 (N_5069,N_4805,N_4861);
xor U5070 (N_5070,N_4807,N_4806);
nor U5071 (N_5071,N_4810,N_4964);
nor U5072 (N_5072,N_4878,N_4952);
nor U5073 (N_5073,N_4876,N_4987);
and U5074 (N_5074,N_4979,N_4881);
xor U5075 (N_5075,N_4838,N_4819);
or U5076 (N_5076,N_4860,N_4965);
or U5077 (N_5077,N_4900,N_4947);
xor U5078 (N_5078,N_4858,N_4826);
nor U5079 (N_5079,N_4942,N_4822);
nand U5080 (N_5080,N_4841,N_4859);
nand U5081 (N_5081,N_4937,N_4989);
xnor U5082 (N_5082,N_4912,N_4832);
xnor U5083 (N_5083,N_4866,N_4941);
or U5084 (N_5084,N_4879,N_4925);
or U5085 (N_5085,N_4936,N_4977);
or U5086 (N_5086,N_4914,N_4972);
nor U5087 (N_5087,N_4885,N_4837);
nand U5088 (N_5088,N_4886,N_4884);
nand U5089 (N_5089,N_4950,N_4985);
nand U5090 (N_5090,N_4993,N_4809);
and U5091 (N_5091,N_4897,N_4864);
nor U5092 (N_5092,N_4959,N_4862);
or U5093 (N_5093,N_4918,N_4871);
nor U5094 (N_5094,N_4894,N_4813);
nand U5095 (N_5095,N_4867,N_4956);
nor U5096 (N_5096,N_4962,N_4892);
or U5097 (N_5097,N_4803,N_4927);
and U5098 (N_5098,N_4924,N_4890);
and U5099 (N_5099,N_4968,N_4991);
or U5100 (N_5100,N_4896,N_4924);
xnor U5101 (N_5101,N_4998,N_4892);
xnor U5102 (N_5102,N_4855,N_4968);
or U5103 (N_5103,N_4936,N_4952);
nor U5104 (N_5104,N_4819,N_4989);
nor U5105 (N_5105,N_4862,N_4920);
or U5106 (N_5106,N_4849,N_4972);
and U5107 (N_5107,N_4984,N_4807);
and U5108 (N_5108,N_4815,N_4806);
xor U5109 (N_5109,N_4806,N_4845);
nor U5110 (N_5110,N_4887,N_4980);
or U5111 (N_5111,N_4907,N_4901);
xor U5112 (N_5112,N_4818,N_4957);
nand U5113 (N_5113,N_4913,N_4822);
or U5114 (N_5114,N_4800,N_4807);
and U5115 (N_5115,N_4947,N_4897);
and U5116 (N_5116,N_4836,N_4929);
and U5117 (N_5117,N_4847,N_4976);
xor U5118 (N_5118,N_4929,N_4965);
or U5119 (N_5119,N_4971,N_4870);
xor U5120 (N_5120,N_4928,N_4986);
nand U5121 (N_5121,N_4982,N_4984);
or U5122 (N_5122,N_4834,N_4904);
xor U5123 (N_5123,N_4853,N_4936);
xor U5124 (N_5124,N_4959,N_4813);
xor U5125 (N_5125,N_4925,N_4822);
nor U5126 (N_5126,N_4863,N_4985);
and U5127 (N_5127,N_4826,N_4958);
nand U5128 (N_5128,N_4898,N_4956);
xnor U5129 (N_5129,N_4847,N_4991);
nand U5130 (N_5130,N_4989,N_4839);
or U5131 (N_5131,N_4988,N_4997);
nand U5132 (N_5132,N_4854,N_4872);
xnor U5133 (N_5133,N_4811,N_4992);
nand U5134 (N_5134,N_4826,N_4815);
xnor U5135 (N_5135,N_4838,N_4961);
and U5136 (N_5136,N_4935,N_4916);
xor U5137 (N_5137,N_4916,N_4879);
xnor U5138 (N_5138,N_4944,N_4921);
xor U5139 (N_5139,N_4855,N_4842);
nand U5140 (N_5140,N_4970,N_4946);
nand U5141 (N_5141,N_4970,N_4806);
xor U5142 (N_5142,N_4841,N_4850);
nor U5143 (N_5143,N_4954,N_4868);
or U5144 (N_5144,N_4976,N_4922);
and U5145 (N_5145,N_4951,N_4962);
nand U5146 (N_5146,N_4904,N_4820);
nand U5147 (N_5147,N_4811,N_4874);
nand U5148 (N_5148,N_4836,N_4812);
xor U5149 (N_5149,N_4821,N_4829);
or U5150 (N_5150,N_4951,N_4975);
xnor U5151 (N_5151,N_4994,N_4872);
xor U5152 (N_5152,N_4982,N_4968);
nor U5153 (N_5153,N_4942,N_4978);
and U5154 (N_5154,N_4964,N_4951);
nor U5155 (N_5155,N_4808,N_4968);
and U5156 (N_5156,N_4961,N_4801);
and U5157 (N_5157,N_4860,N_4974);
and U5158 (N_5158,N_4873,N_4810);
or U5159 (N_5159,N_4834,N_4824);
and U5160 (N_5160,N_4987,N_4952);
and U5161 (N_5161,N_4929,N_4899);
or U5162 (N_5162,N_4994,N_4812);
xor U5163 (N_5163,N_4890,N_4943);
and U5164 (N_5164,N_4818,N_4809);
xor U5165 (N_5165,N_4992,N_4999);
or U5166 (N_5166,N_4881,N_4803);
xnor U5167 (N_5167,N_4811,N_4894);
nand U5168 (N_5168,N_4878,N_4825);
nor U5169 (N_5169,N_4802,N_4973);
nand U5170 (N_5170,N_4981,N_4875);
nor U5171 (N_5171,N_4927,N_4931);
nor U5172 (N_5172,N_4938,N_4823);
xnor U5173 (N_5173,N_4897,N_4814);
or U5174 (N_5174,N_4817,N_4890);
nand U5175 (N_5175,N_4840,N_4832);
xor U5176 (N_5176,N_4847,N_4814);
nand U5177 (N_5177,N_4934,N_4834);
nor U5178 (N_5178,N_4838,N_4897);
xnor U5179 (N_5179,N_4858,N_4945);
nor U5180 (N_5180,N_4917,N_4869);
and U5181 (N_5181,N_4888,N_4818);
xnor U5182 (N_5182,N_4915,N_4914);
and U5183 (N_5183,N_4994,N_4800);
xnor U5184 (N_5184,N_4840,N_4978);
nand U5185 (N_5185,N_4918,N_4874);
nand U5186 (N_5186,N_4963,N_4987);
xor U5187 (N_5187,N_4915,N_4881);
or U5188 (N_5188,N_4976,N_4999);
xnor U5189 (N_5189,N_4857,N_4991);
nor U5190 (N_5190,N_4963,N_4934);
xor U5191 (N_5191,N_4821,N_4916);
xnor U5192 (N_5192,N_4806,N_4950);
xor U5193 (N_5193,N_4898,N_4980);
and U5194 (N_5194,N_4964,N_4927);
and U5195 (N_5195,N_4963,N_4843);
and U5196 (N_5196,N_4875,N_4806);
xnor U5197 (N_5197,N_4930,N_4809);
nand U5198 (N_5198,N_4962,N_4813);
nor U5199 (N_5199,N_4888,N_4898);
xor U5200 (N_5200,N_5057,N_5111);
nor U5201 (N_5201,N_5121,N_5064);
or U5202 (N_5202,N_5136,N_5054);
or U5203 (N_5203,N_5062,N_5135);
nor U5204 (N_5204,N_5080,N_5053);
xor U5205 (N_5205,N_5011,N_5046);
nor U5206 (N_5206,N_5138,N_5106);
nor U5207 (N_5207,N_5079,N_5134);
or U5208 (N_5208,N_5008,N_5021);
or U5209 (N_5209,N_5002,N_5000);
nor U5210 (N_5210,N_5048,N_5124);
xnor U5211 (N_5211,N_5098,N_5063);
xor U5212 (N_5212,N_5003,N_5049);
or U5213 (N_5213,N_5118,N_5151);
nor U5214 (N_5214,N_5092,N_5009);
or U5215 (N_5215,N_5035,N_5109);
nor U5216 (N_5216,N_5018,N_5116);
and U5217 (N_5217,N_5091,N_5084);
xor U5218 (N_5218,N_5101,N_5094);
or U5219 (N_5219,N_5089,N_5119);
xnor U5220 (N_5220,N_5174,N_5031);
nand U5221 (N_5221,N_5073,N_5176);
nor U5222 (N_5222,N_5037,N_5122);
xnor U5223 (N_5223,N_5085,N_5065);
nand U5224 (N_5224,N_5162,N_5165);
nor U5225 (N_5225,N_5032,N_5188);
nand U5226 (N_5226,N_5113,N_5019);
nor U5227 (N_5227,N_5158,N_5010);
nor U5228 (N_5228,N_5128,N_5038);
or U5229 (N_5229,N_5168,N_5072);
or U5230 (N_5230,N_5159,N_5088);
or U5231 (N_5231,N_5114,N_5017);
or U5232 (N_5232,N_5105,N_5086);
or U5233 (N_5233,N_5099,N_5133);
or U5234 (N_5234,N_5082,N_5026);
or U5235 (N_5235,N_5153,N_5110);
or U5236 (N_5236,N_5148,N_5044);
nand U5237 (N_5237,N_5163,N_5130);
and U5238 (N_5238,N_5075,N_5173);
xnor U5239 (N_5239,N_5071,N_5093);
and U5240 (N_5240,N_5103,N_5042);
nor U5241 (N_5241,N_5183,N_5160);
xor U5242 (N_5242,N_5050,N_5115);
nand U5243 (N_5243,N_5125,N_5014);
nor U5244 (N_5244,N_5152,N_5081);
nor U5245 (N_5245,N_5137,N_5095);
xnor U5246 (N_5246,N_5020,N_5144);
nor U5247 (N_5247,N_5164,N_5024);
nand U5248 (N_5248,N_5146,N_5161);
nand U5249 (N_5249,N_5004,N_5051);
xnor U5250 (N_5250,N_5061,N_5142);
and U5251 (N_5251,N_5154,N_5023);
xnor U5252 (N_5252,N_5198,N_5043);
nor U5253 (N_5253,N_5007,N_5132);
or U5254 (N_5254,N_5172,N_5123);
xnor U5255 (N_5255,N_5140,N_5139);
nor U5256 (N_5256,N_5108,N_5199);
or U5257 (N_5257,N_5070,N_5025);
nor U5258 (N_5258,N_5177,N_5193);
nand U5259 (N_5259,N_5087,N_5040);
nor U5260 (N_5260,N_5191,N_5060);
or U5261 (N_5261,N_5022,N_5083);
nor U5262 (N_5262,N_5141,N_5156);
xor U5263 (N_5263,N_5066,N_5001);
or U5264 (N_5264,N_5147,N_5102);
xor U5265 (N_5265,N_5036,N_5126);
or U5266 (N_5266,N_5196,N_5030);
or U5267 (N_5267,N_5096,N_5068);
nand U5268 (N_5268,N_5131,N_5190);
or U5269 (N_5269,N_5005,N_5155);
nand U5270 (N_5270,N_5013,N_5166);
xnor U5271 (N_5271,N_5117,N_5169);
and U5272 (N_5272,N_5077,N_5041);
xnor U5273 (N_5273,N_5112,N_5034);
and U5274 (N_5274,N_5170,N_5090);
or U5275 (N_5275,N_5069,N_5027);
or U5276 (N_5276,N_5186,N_5055);
nor U5277 (N_5277,N_5180,N_5167);
nand U5278 (N_5278,N_5184,N_5143);
and U5279 (N_5279,N_5100,N_5074);
xor U5280 (N_5280,N_5047,N_5059);
nor U5281 (N_5281,N_5076,N_5012);
xor U5282 (N_5282,N_5120,N_5197);
nand U5283 (N_5283,N_5078,N_5187);
xor U5284 (N_5284,N_5097,N_5181);
nand U5285 (N_5285,N_5028,N_5039);
or U5286 (N_5286,N_5045,N_5058);
nor U5287 (N_5287,N_5016,N_5006);
or U5288 (N_5288,N_5171,N_5056);
xor U5289 (N_5289,N_5175,N_5015);
nor U5290 (N_5290,N_5189,N_5052);
xor U5291 (N_5291,N_5029,N_5033);
xor U5292 (N_5292,N_5145,N_5179);
nand U5293 (N_5293,N_5178,N_5107);
nor U5294 (N_5294,N_5067,N_5192);
or U5295 (N_5295,N_5150,N_5129);
and U5296 (N_5296,N_5195,N_5104);
xnor U5297 (N_5297,N_5182,N_5185);
nand U5298 (N_5298,N_5157,N_5149);
nand U5299 (N_5299,N_5127,N_5194);
nor U5300 (N_5300,N_5152,N_5000);
or U5301 (N_5301,N_5150,N_5156);
nor U5302 (N_5302,N_5109,N_5176);
nand U5303 (N_5303,N_5193,N_5008);
or U5304 (N_5304,N_5175,N_5118);
or U5305 (N_5305,N_5084,N_5165);
nand U5306 (N_5306,N_5132,N_5082);
nor U5307 (N_5307,N_5103,N_5051);
xor U5308 (N_5308,N_5109,N_5085);
xnor U5309 (N_5309,N_5005,N_5046);
xnor U5310 (N_5310,N_5160,N_5094);
xnor U5311 (N_5311,N_5028,N_5171);
nor U5312 (N_5312,N_5089,N_5173);
nand U5313 (N_5313,N_5025,N_5120);
nor U5314 (N_5314,N_5023,N_5185);
nand U5315 (N_5315,N_5127,N_5049);
xor U5316 (N_5316,N_5085,N_5128);
xor U5317 (N_5317,N_5023,N_5117);
nand U5318 (N_5318,N_5159,N_5052);
nor U5319 (N_5319,N_5021,N_5063);
nand U5320 (N_5320,N_5161,N_5121);
nand U5321 (N_5321,N_5129,N_5072);
or U5322 (N_5322,N_5127,N_5164);
or U5323 (N_5323,N_5114,N_5065);
nor U5324 (N_5324,N_5177,N_5121);
nand U5325 (N_5325,N_5073,N_5013);
nor U5326 (N_5326,N_5129,N_5144);
and U5327 (N_5327,N_5106,N_5162);
xor U5328 (N_5328,N_5017,N_5003);
nor U5329 (N_5329,N_5116,N_5166);
or U5330 (N_5330,N_5079,N_5177);
nand U5331 (N_5331,N_5058,N_5167);
and U5332 (N_5332,N_5054,N_5189);
and U5333 (N_5333,N_5003,N_5027);
or U5334 (N_5334,N_5121,N_5019);
or U5335 (N_5335,N_5073,N_5185);
and U5336 (N_5336,N_5098,N_5166);
nand U5337 (N_5337,N_5108,N_5055);
xor U5338 (N_5338,N_5121,N_5136);
nor U5339 (N_5339,N_5010,N_5128);
nand U5340 (N_5340,N_5008,N_5077);
nor U5341 (N_5341,N_5195,N_5187);
nand U5342 (N_5342,N_5198,N_5196);
nor U5343 (N_5343,N_5192,N_5078);
nor U5344 (N_5344,N_5054,N_5027);
nand U5345 (N_5345,N_5100,N_5096);
xor U5346 (N_5346,N_5162,N_5016);
nor U5347 (N_5347,N_5077,N_5138);
nor U5348 (N_5348,N_5165,N_5067);
or U5349 (N_5349,N_5009,N_5144);
nand U5350 (N_5350,N_5011,N_5128);
nor U5351 (N_5351,N_5127,N_5024);
or U5352 (N_5352,N_5190,N_5069);
nand U5353 (N_5353,N_5144,N_5140);
or U5354 (N_5354,N_5111,N_5023);
and U5355 (N_5355,N_5025,N_5034);
and U5356 (N_5356,N_5069,N_5096);
or U5357 (N_5357,N_5013,N_5010);
or U5358 (N_5358,N_5087,N_5070);
nor U5359 (N_5359,N_5131,N_5011);
xor U5360 (N_5360,N_5010,N_5075);
or U5361 (N_5361,N_5166,N_5143);
nor U5362 (N_5362,N_5077,N_5192);
nor U5363 (N_5363,N_5065,N_5023);
nand U5364 (N_5364,N_5110,N_5080);
nor U5365 (N_5365,N_5170,N_5175);
nand U5366 (N_5366,N_5082,N_5112);
and U5367 (N_5367,N_5164,N_5080);
or U5368 (N_5368,N_5022,N_5088);
and U5369 (N_5369,N_5032,N_5127);
or U5370 (N_5370,N_5095,N_5132);
and U5371 (N_5371,N_5010,N_5090);
nor U5372 (N_5372,N_5099,N_5145);
nand U5373 (N_5373,N_5163,N_5111);
or U5374 (N_5374,N_5194,N_5022);
and U5375 (N_5375,N_5197,N_5185);
xnor U5376 (N_5376,N_5035,N_5080);
xor U5377 (N_5377,N_5104,N_5084);
nand U5378 (N_5378,N_5114,N_5022);
nand U5379 (N_5379,N_5037,N_5113);
nand U5380 (N_5380,N_5171,N_5089);
xor U5381 (N_5381,N_5023,N_5165);
xor U5382 (N_5382,N_5007,N_5051);
and U5383 (N_5383,N_5104,N_5021);
xnor U5384 (N_5384,N_5026,N_5016);
and U5385 (N_5385,N_5047,N_5014);
nor U5386 (N_5386,N_5025,N_5176);
nor U5387 (N_5387,N_5097,N_5116);
xor U5388 (N_5388,N_5167,N_5041);
xnor U5389 (N_5389,N_5041,N_5106);
nand U5390 (N_5390,N_5040,N_5076);
xor U5391 (N_5391,N_5127,N_5123);
nor U5392 (N_5392,N_5036,N_5109);
and U5393 (N_5393,N_5133,N_5044);
and U5394 (N_5394,N_5132,N_5188);
nor U5395 (N_5395,N_5126,N_5178);
or U5396 (N_5396,N_5003,N_5018);
and U5397 (N_5397,N_5150,N_5161);
and U5398 (N_5398,N_5082,N_5086);
xor U5399 (N_5399,N_5138,N_5120);
or U5400 (N_5400,N_5309,N_5398);
nor U5401 (N_5401,N_5242,N_5281);
nand U5402 (N_5402,N_5363,N_5364);
xor U5403 (N_5403,N_5257,N_5290);
nor U5404 (N_5404,N_5211,N_5213);
and U5405 (N_5405,N_5395,N_5357);
and U5406 (N_5406,N_5342,N_5314);
and U5407 (N_5407,N_5323,N_5367);
nor U5408 (N_5408,N_5391,N_5380);
xnor U5409 (N_5409,N_5236,N_5254);
nand U5410 (N_5410,N_5249,N_5266);
or U5411 (N_5411,N_5372,N_5389);
nor U5412 (N_5412,N_5350,N_5235);
and U5413 (N_5413,N_5221,N_5298);
or U5414 (N_5414,N_5279,N_5346);
and U5415 (N_5415,N_5286,N_5304);
xnor U5416 (N_5416,N_5358,N_5243);
nor U5417 (N_5417,N_5273,N_5351);
and U5418 (N_5418,N_5397,N_5225);
nor U5419 (N_5419,N_5245,N_5277);
xnor U5420 (N_5420,N_5370,N_5232);
or U5421 (N_5421,N_5217,N_5202);
xor U5422 (N_5422,N_5344,N_5335);
nand U5423 (N_5423,N_5271,N_5373);
xnor U5424 (N_5424,N_5348,N_5231);
nand U5425 (N_5425,N_5310,N_5208);
and U5426 (N_5426,N_5387,N_5359);
xor U5427 (N_5427,N_5296,N_5341);
and U5428 (N_5428,N_5285,N_5333);
xnor U5429 (N_5429,N_5276,N_5321);
xnor U5430 (N_5430,N_5331,N_5270);
nor U5431 (N_5431,N_5238,N_5218);
nand U5432 (N_5432,N_5369,N_5345);
or U5433 (N_5433,N_5239,N_5379);
and U5434 (N_5434,N_5396,N_5262);
xor U5435 (N_5435,N_5265,N_5337);
nor U5436 (N_5436,N_5340,N_5360);
or U5437 (N_5437,N_5224,N_5216);
nand U5438 (N_5438,N_5206,N_5301);
nor U5439 (N_5439,N_5317,N_5205);
or U5440 (N_5440,N_5347,N_5336);
xor U5441 (N_5441,N_5220,N_5252);
and U5442 (N_5442,N_5300,N_5280);
or U5443 (N_5443,N_5201,N_5316);
nor U5444 (N_5444,N_5219,N_5390);
or U5445 (N_5445,N_5349,N_5318);
or U5446 (N_5446,N_5308,N_5263);
xnor U5447 (N_5447,N_5203,N_5385);
xnor U5448 (N_5448,N_5320,N_5269);
and U5449 (N_5449,N_5394,N_5393);
xnor U5450 (N_5450,N_5366,N_5223);
nand U5451 (N_5451,N_5388,N_5361);
nor U5452 (N_5452,N_5294,N_5334);
or U5453 (N_5453,N_5303,N_5275);
nand U5454 (N_5454,N_5392,N_5283);
and U5455 (N_5455,N_5255,N_5315);
nand U5456 (N_5456,N_5375,N_5326);
xor U5457 (N_5457,N_5258,N_5291);
and U5458 (N_5458,N_5332,N_5297);
nand U5459 (N_5459,N_5227,N_5233);
and U5460 (N_5460,N_5378,N_5377);
nor U5461 (N_5461,N_5311,N_5259);
nor U5462 (N_5462,N_5246,N_5287);
nor U5463 (N_5463,N_5325,N_5302);
nor U5464 (N_5464,N_5295,N_5228);
nand U5465 (N_5465,N_5278,N_5204);
nand U5466 (N_5466,N_5237,N_5288);
nor U5467 (N_5467,N_5212,N_5305);
and U5468 (N_5468,N_5247,N_5328);
nand U5469 (N_5469,N_5374,N_5244);
nand U5470 (N_5470,N_5306,N_5312);
and U5471 (N_5471,N_5207,N_5319);
nand U5472 (N_5472,N_5368,N_5248);
or U5473 (N_5473,N_5329,N_5355);
or U5474 (N_5474,N_5362,N_5322);
xnor U5475 (N_5475,N_5324,N_5230);
xor U5476 (N_5476,N_5253,N_5313);
and U5477 (N_5477,N_5381,N_5338);
nor U5478 (N_5478,N_5274,N_5339);
xnor U5479 (N_5479,N_5251,N_5356);
xnor U5480 (N_5480,N_5384,N_5327);
nand U5481 (N_5481,N_5352,N_5267);
and U5482 (N_5482,N_5222,N_5354);
xor U5483 (N_5483,N_5376,N_5382);
nor U5484 (N_5484,N_5256,N_5282);
nand U5485 (N_5485,N_5289,N_5365);
and U5486 (N_5486,N_5260,N_5272);
xor U5487 (N_5487,N_5353,N_5307);
xnor U5488 (N_5488,N_5261,N_5299);
and U5489 (N_5489,N_5399,N_5241);
xnor U5490 (N_5490,N_5200,N_5209);
xnor U5491 (N_5491,N_5383,N_5292);
nand U5492 (N_5492,N_5343,N_5240);
or U5493 (N_5493,N_5330,N_5264);
or U5494 (N_5494,N_5226,N_5210);
nand U5495 (N_5495,N_5284,N_5250);
xor U5496 (N_5496,N_5234,N_5268);
nand U5497 (N_5497,N_5229,N_5386);
nand U5498 (N_5498,N_5215,N_5293);
and U5499 (N_5499,N_5214,N_5371);
xnor U5500 (N_5500,N_5301,N_5238);
or U5501 (N_5501,N_5354,N_5390);
xor U5502 (N_5502,N_5204,N_5373);
nand U5503 (N_5503,N_5217,N_5326);
xor U5504 (N_5504,N_5377,N_5275);
nor U5505 (N_5505,N_5236,N_5348);
and U5506 (N_5506,N_5201,N_5385);
and U5507 (N_5507,N_5269,N_5347);
or U5508 (N_5508,N_5347,N_5328);
nor U5509 (N_5509,N_5294,N_5276);
nor U5510 (N_5510,N_5356,N_5319);
xor U5511 (N_5511,N_5230,N_5323);
xnor U5512 (N_5512,N_5279,N_5321);
nand U5513 (N_5513,N_5252,N_5377);
nor U5514 (N_5514,N_5262,N_5216);
or U5515 (N_5515,N_5320,N_5321);
xor U5516 (N_5516,N_5232,N_5328);
or U5517 (N_5517,N_5375,N_5258);
xor U5518 (N_5518,N_5271,N_5205);
and U5519 (N_5519,N_5269,N_5330);
nand U5520 (N_5520,N_5295,N_5359);
or U5521 (N_5521,N_5320,N_5270);
nor U5522 (N_5522,N_5299,N_5318);
and U5523 (N_5523,N_5214,N_5288);
xnor U5524 (N_5524,N_5245,N_5375);
xnor U5525 (N_5525,N_5392,N_5231);
nor U5526 (N_5526,N_5266,N_5390);
xnor U5527 (N_5527,N_5213,N_5314);
or U5528 (N_5528,N_5307,N_5384);
or U5529 (N_5529,N_5389,N_5267);
and U5530 (N_5530,N_5355,N_5354);
and U5531 (N_5531,N_5213,N_5283);
nand U5532 (N_5532,N_5222,N_5328);
or U5533 (N_5533,N_5307,N_5376);
or U5534 (N_5534,N_5252,N_5200);
and U5535 (N_5535,N_5204,N_5221);
nand U5536 (N_5536,N_5319,N_5216);
nor U5537 (N_5537,N_5356,N_5381);
nand U5538 (N_5538,N_5269,N_5389);
xor U5539 (N_5539,N_5332,N_5325);
nand U5540 (N_5540,N_5270,N_5349);
nand U5541 (N_5541,N_5371,N_5317);
xor U5542 (N_5542,N_5335,N_5217);
xor U5543 (N_5543,N_5340,N_5350);
xnor U5544 (N_5544,N_5395,N_5254);
and U5545 (N_5545,N_5305,N_5338);
nor U5546 (N_5546,N_5347,N_5335);
nand U5547 (N_5547,N_5318,N_5245);
nand U5548 (N_5548,N_5274,N_5307);
xnor U5549 (N_5549,N_5364,N_5247);
and U5550 (N_5550,N_5288,N_5236);
and U5551 (N_5551,N_5368,N_5327);
xnor U5552 (N_5552,N_5225,N_5273);
xnor U5553 (N_5553,N_5245,N_5276);
or U5554 (N_5554,N_5255,N_5252);
and U5555 (N_5555,N_5229,N_5282);
nand U5556 (N_5556,N_5270,N_5295);
xor U5557 (N_5557,N_5229,N_5334);
xnor U5558 (N_5558,N_5390,N_5363);
or U5559 (N_5559,N_5222,N_5269);
or U5560 (N_5560,N_5350,N_5206);
nand U5561 (N_5561,N_5257,N_5374);
and U5562 (N_5562,N_5290,N_5292);
xor U5563 (N_5563,N_5333,N_5368);
xnor U5564 (N_5564,N_5284,N_5215);
and U5565 (N_5565,N_5288,N_5386);
xnor U5566 (N_5566,N_5381,N_5388);
or U5567 (N_5567,N_5306,N_5237);
nand U5568 (N_5568,N_5313,N_5384);
xnor U5569 (N_5569,N_5208,N_5248);
xor U5570 (N_5570,N_5303,N_5325);
or U5571 (N_5571,N_5201,N_5312);
and U5572 (N_5572,N_5291,N_5398);
nand U5573 (N_5573,N_5374,N_5248);
and U5574 (N_5574,N_5247,N_5376);
nor U5575 (N_5575,N_5306,N_5258);
or U5576 (N_5576,N_5232,N_5392);
nor U5577 (N_5577,N_5227,N_5277);
xor U5578 (N_5578,N_5277,N_5285);
xnor U5579 (N_5579,N_5396,N_5365);
or U5580 (N_5580,N_5312,N_5246);
nand U5581 (N_5581,N_5212,N_5332);
and U5582 (N_5582,N_5394,N_5346);
and U5583 (N_5583,N_5223,N_5238);
nand U5584 (N_5584,N_5239,N_5275);
xnor U5585 (N_5585,N_5262,N_5363);
nor U5586 (N_5586,N_5261,N_5390);
or U5587 (N_5587,N_5369,N_5351);
or U5588 (N_5588,N_5384,N_5230);
or U5589 (N_5589,N_5334,N_5340);
and U5590 (N_5590,N_5282,N_5346);
or U5591 (N_5591,N_5203,N_5246);
or U5592 (N_5592,N_5283,N_5210);
or U5593 (N_5593,N_5345,N_5387);
nand U5594 (N_5594,N_5309,N_5268);
or U5595 (N_5595,N_5381,N_5223);
or U5596 (N_5596,N_5324,N_5315);
nor U5597 (N_5597,N_5361,N_5334);
nand U5598 (N_5598,N_5383,N_5243);
and U5599 (N_5599,N_5286,N_5386);
nand U5600 (N_5600,N_5530,N_5432);
nand U5601 (N_5601,N_5431,N_5547);
or U5602 (N_5602,N_5414,N_5582);
nor U5603 (N_5603,N_5444,N_5552);
xor U5604 (N_5604,N_5509,N_5579);
or U5605 (N_5605,N_5409,N_5571);
or U5606 (N_5606,N_5482,N_5485);
or U5607 (N_5607,N_5452,N_5425);
nand U5608 (N_5608,N_5551,N_5540);
nor U5609 (N_5609,N_5463,N_5575);
nand U5610 (N_5610,N_5440,N_5422);
and U5611 (N_5611,N_5439,N_5528);
or U5612 (N_5612,N_5558,N_5402);
or U5613 (N_5613,N_5459,N_5597);
or U5614 (N_5614,N_5549,N_5531);
or U5615 (N_5615,N_5487,N_5462);
nand U5616 (N_5616,N_5416,N_5455);
xnor U5617 (N_5617,N_5460,N_5553);
and U5618 (N_5618,N_5491,N_5546);
xor U5619 (N_5619,N_5594,N_5591);
or U5620 (N_5620,N_5534,N_5433);
xor U5621 (N_5621,N_5410,N_5492);
nand U5622 (N_5622,N_5458,N_5541);
and U5623 (N_5623,N_5511,N_5488);
and U5624 (N_5624,N_5465,N_5523);
or U5625 (N_5625,N_5415,N_5419);
nor U5626 (N_5626,N_5464,N_5420);
or U5627 (N_5627,N_5484,N_5477);
nor U5628 (N_5628,N_5426,N_5461);
nor U5629 (N_5629,N_5527,N_5581);
nor U5630 (N_5630,N_5468,N_5479);
nand U5631 (N_5631,N_5471,N_5505);
nor U5632 (N_5632,N_5430,N_5584);
or U5633 (N_5633,N_5407,N_5595);
xnor U5634 (N_5634,N_5489,N_5542);
and U5635 (N_5635,N_5588,N_5580);
nand U5636 (N_5636,N_5457,N_5536);
xor U5637 (N_5637,N_5500,N_5592);
xnor U5638 (N_5638,N_5490,N_5445);
nor U5639 (N_5639,N_5454,N_5599);
or U5640 (N_5640,N_5586,N_5532);
or U5641 (N_5641,N_5565,N_5400);
nor U5642 (N_5642,N_5548,N_5495);
or U5643 (N_5643,N_5418,N_5576);
xor U5644 (N_5644,N_5494,N_5429);
and U5645 (N_5645,N_5556,N_5486);
nand U5646 (N_5646,N_5545,N_5568);
or U5647 (N_5647,N_5435,N_5449);
or U5648 (N_5648,N_5503,N_5470);
xor U5649 (N_5649,N_5537,N_5519);
nand U5650 (N_5650,N_5434,N_5535);
nor U5651 (N_5651,N_5517,N_5555);
or U5652 (N_5652,N_5590,N_5467);
and U5653 (N_5653,N_5559,N_5564);
or U5654 (N_5654,N_5566,N_5498);
xnor U5655 (N_5655,N_5557,N_5501);
or U5656 (N_5656,N_5572,N_5596);
or U5657 (N_5657,N_5474,N_5480);
nor U5658 (N_5658,N_5521,N_5543);
nor U5659 (N_5659,N_5447,N_5522);
or U5660 (N_5660,N_5413,N_5450);
nand U5661 (N_5661,N_5421,N_5401);
nand U5662 (N_5662,N_5404,N_5436);
and U5663 (N_5663,N_5518,N_5563);
or U5664 (N_5664,N_5411,N_5403);
nand U5665 (N_5665,N_5526,N_5504);
xnor U5666 (N_5666,N_5512,N_5524);
xnor U5667 (N_5667,N_5438,N_5507);
and U5668 (N_5668,N_5550,N_5508);
and U5669 (N_5669,N_5441,N_5483);
or U5670 (N_5670,N_5497,N_5473);
nor U5671 (N_5671,N_5481,N_5446);
xor U5672 (N_5672,N_5456,N_5520);
xnor U5673 (N_5673,N_5562,N_5587);
or U5674 (N_5674,N_5516,N_5573);
xor U5675 (N_5675,N_5408,N_5442);
or U5676 (N_5676,N_5589,N_5499);
nand U5677 (N_5677,N_5514,N_5560);
xor U5678 (N_5678,N_5448,N_5478);
xor U5679 (N_5679,N_5510,N_5513);
xnor U5680 (N_5680,N_5574,N_5443);
nand U5681 (N_5681,N_5515,N_5506);
or U5682 (N_5682,N_5525,N_5585);
nor U5683 (N_5683,N_5598,N_5593);
nor U5684 (N_5684,N_5405,N_5437);
nand U5685 (N_5685,N_5554,N_5539);
nor U5686 (N_5686,N_5469,N_5502);
or U5687 (N_5687,N_5544,N_5428);
and U5688 (N_5688,N_5577,N_5496);
nor U5689 (N_5689,N_5412,N_5570);
nand U5690 (N_5690,N_5451,N_5423);
nand U5691 (N_5691,N_5561,N_5466);
and U5692 (N_5692,N_5578,N_5476);
nand U5693 (N_5693,N_5583,N_5475);
or U5694 (N_5694,N_5533,N_5567);
or U5695 (N_5695,N_5417,N_5424);
or U5696 (N_5696,N_5493,N_5406);
xor U5697 (N_5697,N_5538,N_5427);
xor U5698 (N_5698,N_5569,N_5472);
nand U5699 (N_5699,N_5529,N_5453);
nor U5700 (N_5700,N_5466,N_5482);
nand U5701 (N_5701,N_5417,N_5443);
or U5702 (N_5702,N_5537,N_5465);
xor U5703 (N_5703,N_5561,N_5412);
xor U5704 (N_5704,N_5519,N_5458);
and U5705 (N_5705,N_5520,N_5540);
and U5706 (N_5706,N_5494,N_5516);
or U5707 (N_5707,N_5443,N_5480);
nor U5708 (N_5708,N_5562,N_5442);
xnor U5709 (N_5709,N_5558,N_5409);
or U5710 (N_5710,N_5439,N_5593);
nor U5711 (N_5711,N_5409,N_5542);
nand U5712 (N_5712,N_5513,N_5451);
and U5713 (N_5713,N_5525,N_5549);
xnor U5714 (N_5714,N_5590,N_5574);
or U5715 (N_5715,N_5409,N_5488);
nand U5716 (N_5716,N_5448,N_5462);
and U5717 (N_5717,N_5504,N_5568);
and U5718 (N_5718,N_5497,N_5492);
nand U5719 (N_5719,N_5571,N_5556);
nand U5720 (N_5720,N_5433,N_5400);
nand U5721 (N_5721,N_5477,N_5444);
nor U5722 (N_5722,N_5441,N_5492);
or U5723 (N_5723,N_5429,N_5415);
or U5724 (N_5724,N_5480,N_5563);
or U5725 (N_5725,N_5573,N_5558);
xnor U5726 (N_5726,N_5414,N_5436);
and U5727 (N_5727,N_5556,N_5404);
nand U5728 (N_5728,N_5536,N_5581);
or U5729 (N_5729,N_5569,N_5412);
nand U5730 (N_5730,N_5510,N_5583);
or U5731 (N_5731,N_5599,N_5535);
or U5732 (N_5732,N_5520,N_5450);
or U5733 (N_5733,N_5573,N_5457);
and U5734 (N_5734,N_5492,N_5475);
nor U5735 (N_5735,N_5530,N_5531);
nand U5736 (N_5736,N_5548,N_5438);
xor U5737 (N_5737,N_5420,N_5415);
and U5738 (N_5738,N_5505,N_5484);
nand U5739 (N_5739,N_5545,N_5517);
and U5740 (N_5740,N_5487,N_5509);
xor U5741 (N_5741,N_5494,N_5404);
nand U5742 (N_5742,N_5429,N_5580);
xor U5743 (N_5743,N_5486,N_5580);
or U5744 (N_5744,N_5400,N_5500);
or U5745 (N_5745,N_5535,N_5528);
nand U5746 (N_5746,N_5485,N_5407);
nor U5747 (N_5747,N_5445,N_5566);
and U5748 (N_5748,N_5450,N_5515);
and U5749 (N_5749,N_5535,N_5427);
xor U5750 (N_5750,N_5570,N_5411);
and U5751 (N_5751,N_5525,N_5599);
and U5752 (N_5752,N_5433,N_5441);
xor U5753 (N_5753,N_5570,N_5485);
or U5754 (N_5754,N_5467,N_5452);
nand U5755 (N_5755,N_5436,N_5506);
and U5756 (N_5756,N_5490,N_5525);
nor U5757 (N_5757,N_5415,N_5553);
and U5758 (N_5758,N_5510,N_5534);
nand U5759 (N_5759,N_5409,N_5597);
xnor U5760 (N_5760,N_5531,N_5577);
xor U5761 (N_5761,N_5593,N_5580);
nand U5762 (N_5762,N_5442,N_5599);
nor U5763 (N_5763,N_5428,N_5506);
xor U5764 (N_5764,N_5554,N_5512);
or U5765 (N_5765,N_5402,N_5478);
xnor U5766 (N_5766,N_5540,N_5539);
nor U5767 (N_5767,N_5460,N_5546);
nand U5768 (N_5768,N_5474,N_5402);
and U5769 (N_5769,N_5424,N_5580);
nand U5770 (N_5770,N_5504,N_5508);
nor U5771 (N_5771,N_5426,N_5422);
nand U5772 (N_5772,N_5451,N_5553);
and U5773 (N_5773,N_5583,N_5420);
xor U5774 (N_5774,N_5550,N_5545);
nor U5775 (N_5775,N_5565,N_5595);
or U5776 (N_5776,N_5499,N_5400);
nor U5777 (N_5777,N_5572,N_5414);
nor U5778 (N_5778,N_5491,N_5502);
nor U5779 (N_5779,N_5436,N_5400);
and U5780 (N_5780,N_5427,N_5510);
xor U5781 (N_5781,N_5479,N_5577);
and U5782 (N_5782,N_5453,N_5476);
and U5783 (N_5783,N_5467,N_5510);
and U5784 (N_5784,N_5403,N_5576);
xnor U5785 (N_5785,N_5546,N_5429);
and U5786 (N_5786,N_5410,N_5423);
and U5787 (N_5787,N_5540,N_5565);
nand U5788 (N_5788,N_5468,N_5552);
nand U5789 (N_5789,N_5481,N_5571);
or U5790 (N_5790,N_5597,N_5501);
nor U5791 (N_5791,N_5421,N_5458);
or U5792 (N_5792,N_5549,N_5471);
or U5793 (N_5793,N_5509,N_5491);
nand U5794 (N_5794,N_5534,N_5455);
nor U5795 (N_5795,N_5440,N_5415);
nand U5796 (N_5796,N_5434,N_5551);
or U5797 (N_5797,N_5519,N_5536);
nand U5798 (N_5798,N_5468,N_5533);
or U5799 (N_5799,N_5592,N_5400);
nand U5800 (N_5800,N_5778,N_5735);
nor U5801 (N_5801,N_5671,N_5741);
nand U5802 (N_5802,N_5694,N_5618);
and U5803 (N_5803,N_5784,N_5701);
or U5804 (N_5804,N_5779,N_5617);
and U5805 (N_5805,N_5691,N_5733);
or U5806 (N_5806,N_5670,N_5685);
and U5807 (N_5807,N_5751,N_5697);
nor U5808 (N_5808,N_5602,N_5660);
nor U5809 (N_5809,N_5608,N_5677);
nor U5810 (N_5810,N_5659,N_5758);
xnor U5811 (N_5811,N_5661,N_5773);
and U5812 (N_5812,N_5668,N_5774);
and U5813 (N_5813,N_5795,N_5787);
nand U5814 (N_5814,N_5702,N_5706);
nand U5815 (N_5815,N_5639,N_5652);
nor U5816 (N_5816,N_5768,N_5745);
or U5817 (N_5817,N_5698,N_5709);
nand U5818 (N_5818,N_5720,N_5616);
and U5819 (N_5819,N_5646,N_5610);
and U5820 (N_5820,N_5667,N_5793);
nor U5821 (N_5821,N_5693,N_5759);
nor U5822 (N_5822,N_5719,N_5731);
and U5823 (N_5823,N_5713,N_5603);
nor U5824 (N_5824,N_5664,N_5750);
nand U5825 (N_5825,N_5765,N_5654);
or U5826 (N_5826,N_5782,N_5786);
or U5827 (N_5827,N_5715,N_5681);
nand U5828 (N_5828,N_5658,N_5737);
and U5829 (N_5829,N_5615,N_5754);
or U5830 (N_5830,N_5682,N_5637);
nor U5831 (N_5831,N_5675,N_5647);
xor U5832 (N_5832,N_5730,N_5755);
nor U5833 (N_5833,N_5767,N_5743);
nor U5834 (N_5834,N_5649,N_5764);
and U5835 (N_5835,N_5714,N_5680);
and U5836 (N_5836,N_5729,N_5601);
xnor U5837 (N_5837,N_5742,N_5666);
nand U5838 (N_5838,N_5699,N_5689);
or U5839 (N_5839,N_5789,N_5611);
and U5840 (N_5840,N_5609,N_5688);
nor U5841 (N_5841,N_5716,N_5732);
and U5842 (N_5842,N_5704,N_5656);
or U5843 (N_5843,N_5695,N_5636);
nand U5844 (N_5844,N_5757,N_5629);
or U5845 (N_5845,N_5738,N_5727);
and U5846 (N_5846,N_5711,N_5781);
and U5847 (N_5847,N_5674,N_5631);
and U5848 (N_5848,N_5687,N_5790);
and U5849 (N_5849,N_5628,N_5621);
nor U5850 (N_5850,N_5799,N_5606);
nand U5851 (N_5851,N_5769,N_5683);
and U5852 (N_5852,N_5605,N_5613);
nand U5853 (N_5853,N_5644,N_5663);
nor U5854 (N_5854,N_5756,N_5722);
xnor U5855 (N_5855,N_5712,N_5627);
nand U5856 (N_5856,N_5726,N_5638);
xor U5857 (N_5857,N_5771,N_5734);
or U5858 (N_5858,N_5665,N_5770);
xnor U5859 (N_5859,N_5761,N_5672);
xor U5860 (N_5860,N_5622,N_5619);
and U5861 (N_5861,N_5673,N_5696);
or U5862 (N_5862,N_5653,N_5788);
xor U5863 (N_5863,N_5752,N_5728);
or U5864 (N_5864,N_5783,N_5798);
nand U5865 (N_5865,N_5650,N_5797);
and U5866 (N_5866,N_5643,N_5717);
nand U5867 (N_5867,N_5600,N_5703);
xor U5868 (N_5868,N_5725,N_5707);
nand U5869 (N_5869,N_5791,N_5633);
nand U5870 (N_5870,N_5692,N_5724);
or U5871 (N_5871,N_5744,N_5642);
nor U5872 (N_5872,N_5669,N_5777);
nand U5873 (N_5873,N_5641,N_5657);
xor U5874 (N_5874,N_5655,N_5651);
nor U5875 (N_5875,N_5753,N_5705);
or U5876 (N_5876,N_5700,N_5676);
xor U5877 (N_5877,N_5645,N_5746);
and U5878 (N_5878,N_5766,N_5625);
and U5879 (N_5879,N_5775,N_5772);
or U5880 (N_5880,N_5624,N_5678);
nand U5881 (N_5881,N_5635,N_5612);
and U5882 (N_5882,N_5785,N_5634);
nor U5883 (N_5883,N_5760,N_5747);
or U5884 (N_5884,N_5762,N_5690);
nor U5885 (N_5885,N_5796,N_5718);
or U5886 (N_5886,N_5736,N_5632);
nand U5887 (N_5887,N_5614,N_5684);
and U5888 (N_5888,N_5620,N_5749);
nor U5889 (N_5889,N_5604,N_5648);
nor U5890 (N_5890,N_5623,N_5739);
and U5891 (N_5891,N_5607,N_5630);
nor U5892 (N_5892,N_5662,N_5763);
xor U5893 (N_5893,N_5748,N_5776);
nor U5894 (N_5894,N_5708,N_5721);
and U5895 (N_5895,N_5723,N_5780);
nor U5896 (N_5896,N_5686,N_5792);
nor U5897 (N_5897,N_5740,N_5640);
nand U5898 (N_5898,N_5794,N_5679);
nand U5899 (N_5899,N_5710,N_5626);
xnor U5900 (N_5900,N_5733,N_5769);
xor U5901 (N_5901,N_5689,N_5663);
xor U5902 (N_5902,N_5643,N_5798);
nand U5903 (N_5903,N_5735,N_5689);
nand U5904 (N_5904,N_5674,N_5601);
nand U5905 (N_5905,N_5683,N_5799);
nor U5906 (N_5906,N_5620,N_5773);
and U5907 (N_5907,N_5621,N_5757);
or U5908 (N_5908,N_5794,N_5625);
and U5909 (N_5909,N_5706,N_5614);
nor U5910 (N_5910,N_5774,N_5731);
or U5911 (N_5911,N_5781,N_5615);
xnor U5912 (N_5912,N_5603,N_5768);
nand U5913 (N_5913,N_5797,N_5748);
nand U5914 (N_5914,N_5722,N_5668);
xnor U5915 (N_5915,N_5724,N_5723);
or U5916 (N_5916,N_5763,N_5679);
xnor U5917 (N_5917,N_5725,N_5669);
xor U5918 (N_5918,N_5662,N_5696);
nor U5919 (N_5919,N_5786,N_5603);
or U5920 (N_5920,N_5650,N_5706);
nand U5921 (N_5921,N_5794,N_5610);
xor U5922 (N_5922,N_5690,N_5634);
or U5923 (N_5923,N_5799,N_5722);
nand U5924 (N_5924,N_5759,N_5764);
and U5925 (N_5925,N_5637,N_5764);
nand U5926 (N_5926,N_5756,N_5600);
nor U5927 (N_5927,N_5732,N_5734);
xor U5928 (N_5928,N_5613,N_5603);
nand U5929 (N_5929,N_5737,N_5728);
nor U5930 (N_5930,N_5724,N_5666);
xnor U5931 (N_5931,N_5715,N_5782);
xnor U5932 (N_5932,N_5699,N_5760);
xnor U5933 (N_5933,N_5622,N_5793);
and U5934 (N_5934,N_5667,N_5679);
nand U5935 (N_5935,N_5603,N_5662);
nand U5936 (N_5936,N_5674,N_5723);
nand U5937 (N_5937,N_5641,N_5600);
nor U5938 (N_5938,N_5735,N_5605);
or U5939 (N_5939,N_5736,N_5785);
or U5940 (N_5940,N_5708,N_5682);
nand U5941 (N_5941,N_5727,N_5773);
and U5942 (N_5942,N_5786,N_5752);
and U5943 (N_5943,N_5787,N_5638);
or U5944 (N_5944,N_5790,N_5640);
xnor U5945 (N_5945,N_5688,N_5636);
and U5946 (N_5946,N_5735,N_5757);
xnor U5947 (N_5947,N_5630,N_5735);
xor U5948 (N_5948,N_5791,N_5636);
xor U5949 (N_5949,N_5630,N_5611);
and U5950 (N_5950,N_5756,N_5715);
nor U5951 (N_5951,N_5677,N_5623);
nand U5952 (N_5952,N_5642,N_5703);
and U5953 (N_5953,N_5620,N_5640);
xor U5954 (N_5954,N_5651,N_5745);
xor U5955 (N_5955,N_5681,N_5793);
or U5956 (N_5956,N_5677,N_5707);
or U5957 (N_5957,N_5692,N_5725);
and U5958 (N_5958,N_5705,N_5749);
or U5959 (N_5959,N_5704,N_5624);
xnor U5960 (N_5960,N_5636,N_5664);
nor U5961 (N_5961,N_5690,N_5714);
xor U5962 (N_5962,N_5644,N_5669);
or U5963 (N_5963,N_5679,N_5649);
nor U5964 (N_5964,N_5612,N_5609);
xor U5965 (N_5965,N_5684,N_5669);
nor U5966 (N_5966,N_5621,N_5687);
nand U5967 (N_5967,N_5645,N_5758);
xor U5968 (N_5968,N_5605,N_5752);
xnor U5969 (N_5969,N_5602,N_5643);
nand U5970 (N_5970,N_5774,N_5781);
nand U5971 (N_5971,N_5721,N_5630);
nand U5972 (N_5972,N_5639,N_5683);
or U5973 (N_5973,N_5739,N_5759);
or U5974 (N_5974,N_5682,N_5756);
and U5975 (N_5975,N_5711,N_5611);
xnor U5976 (N_5976,N_5737,N_5675);
or U5977 (N_5977,N_5707,N_5689);
nor U5978 (N_5978,N_5692,N_5701);
xor U5979 (N_5979,N_5653,N_5778);
and U5980 (N_5980,N_5755,N_5726);
xor U5981 (N_5981,N_5632,N_5764);
and U5982 (N_5982,N_5645,N_5799);
nor U5983 (N_5983,N_5740,N_5656);
or U5984 (N_5984,N_5755,N_5767);
nor U5985 (N_5985,N_5660,N_5673);
or U5986 (N_5986,N_5602,N_5745);
xor U5987 (N_5987,N_5666,N_5760);
nor U5988 (N_5988,N_5684,N_5790);
nand U5989 (N_5989,N_5643,N_5760);
nand U5990 (N_5990,N_5760,N_5754);
or U5991 (N_5991,N_5723,N_5618);
or U5992 (N_5992,N_5645,N_5652);
or U5993 (N_5993,N_5736,N_5676);
xor U5994 (N_5994,N_5679,N_5775);
or U5995 (N_5995,N_5735,N_5742);
or U5996 (N_5996,N_5720,N_5631);
nor U5997 (N_5997,N_5710,N_5736);
xor U5998 (N_5998,N_5746,N_5614);
nand U5999 (N_5999,N_5781,N_5717);
and U6000 (N_6000,N_5925,N_5841);
xor U6001 (N_6001,N_5859,N_5945);
or U6002 (N_6002,N_5939,N_5931);
and U6003 (N_6003,N_5904,N_5873);
and U6004 (N_6004,N_5979,N_5840);
nor U6005 (N_6005,N_5932,N_5962);
or U6006 (N_6006,N_5902,N_5888);
or U6007 (N_6007,N_5834,N_5814);
xor U6008 (N_6008,N_5960,N_5848);
nor U6009 (N_6009,N_5894,N_5938);
or U6010 (N_6010,N_5920,N_5967);
nor U6011 (N_6011,N_5849,N_5850);
nor U6012 (N_6012,N_5874,N_5852);
or U6013 (N_6013,N_5838,N_5919);
or U6014 (N_6014,N_5989,N_5918);
and U6015 (N_6015,N_5959,N_5993);
and U6016 (N_6016,N_5804,N_5858);
nor U6017 (N_6017,N_5926,N_5826);
nor U6018 (N_6018,N_5942,N_5875);
and U6019 (N_6019,N_5806,N_5997);
or U6020 (N_6020,N_5803,N_5981);
and U6021 (N_6021,N_5909,N_5820);
and U6022 (N_6022,N_5941,N_5955);
and U6023 (N_6023,N_5897,N_5907);
nor U6024 (N_6024,N_5936,N_5827);
or U6025 (N_6025,N_5843,N_5898);
nand U6026 (N_6026,N_5802,N_5893);
nand U6027 (N_6027,N_5978,N_5952);
nand U6028 (N_6028,N_5985,N_5801);
nor U6029 (N_6029,N_5964,N_5924);
nand U6030 (N_6030,N_5851,N_5805);
nor U6031 (N_6031,N_5903,N_5928);
and U6032 (N_6032,N_5914,N_5881);
and U6033 (N_6033,N_5998,N_5988);
xnor U6034 (N_6034,N_5976,N_5863);
and U6035 (N_6035,N_5808,N_5934);
nand U6036 (N_6036,N_5974,N_5867);
nor U6037 (N_6037,N_5910,N_5922);
xnor U6038 (N_6038,N_5870,N_5807);
or U6039 (N_6039,N_5833,N_5800);
nand U6040 (N_6040,N_5865,N_5895);
nor U6041 (N_6041,N_5946,N_5930);
or U6042 (N_6042,N_5882,N_5809);
and U6043 (N_6043,N_5958,N_5856);
nor U6044 (N_6044,N_5823,N_5966);
nor U6045 (N_6045,N_5994,N_5995);
and U6046 (N_6046,N_5821,N_5825);
nand U6047 (N_6047,N_5970,N_5868);
or U6048 (N_6048,N_5954,N_5975);
nor U6049 (N_6049,N_5855,N_5908);
xnor U6050 (N_6050,N_5982,N_5861);
nor U6051 (N_6051,N_5933,N_5877);
nor U6052 (N_6052,N_5886,N_5832);
or U6053 (N_6053,N_5857,N_5990);
nand U6054 (N_6054,N_5890,N_5937);
nand U6055 (N_6055,N_5829,N_5984);
xor U6056 (N_6056,N_5973,N_5923);
nand U6057 (N_6057,N_5911,N_5847);
nor U6058 (N_6058,N_5815,N_5983);
nor U6059 (N_6059,N_5817,N_5810);
or U6060 (N_6060,N_5912,N_5862);
or U6061 (N_6061,N_5916,N_5921);
nand U6062 (N_6062,N_5830,N_5950);
nor U6063 (N_6063,N_5831,N_5980);
or U6064 (N_6064,N_5949,N_5813);
nor U6065 (N_6065,N_5883,N_5819);
xor U6066 (N_6066,N_5889,N_5887);
and U6067 (N_6067,N_5951,N_5835);
nor U6068 (N_6068,N_5953,N_5824);
nand U6069 (N_6069,N_5977,N_5876);
or U6070 (N_6070,N_5869,N_5822);
or U6071 (N_6071,N_5992,N_5961);
or U6072 (N_6072,N_5818,N_5996);
xnor U6073 (N_6073,N_5811,N_5844);
nor U6074 (N_6074,N_5812,N_5971);
and U6075 (N_6075,N_5956,N_5836);
nand U6076 (N_6076,N_5884,N_5905);
or U6077 (N_6077,N_5854,N_5880);
or U6078 (N_6078,N_5846,N_5943);
nand U6079 (N_6079,N_5842,N_5947);
xor U6080 (N_6080,N_5871,N_5900);
or U6081 (N_6081,N_5866,N_5816);
or U6082 (N_6082,N_5944,N_5853);
nor U6083 (N_6083,N_5927,N_5987);
and U6084 (N_6084,N_5906,N_5878);
xnor U6085 (N_6085,N_5972,N_5899);
nand U6086 (N_6086,N_5913,N_5940);
and U6087 (N_6087,N_5935,N_5968);
and U6088 (N_6088,N_5872,N_5929);
xnor U6089 (N_6089,N_5845,N_5901);
nor U6090 (N_6090,N_5948,N_5969);
xor U6091 (N_6091,N_5986,N_5837);
nor U6092 (N_6092,N_5915,N_5999);
nor U6093 (N_6093,N_5963,N_5965);
or U6094 (N_6094,N_5839,N_5892);
nor U6095 (N_6095,N_5879,N_5885);
nand U6096 (N_6096,N_5957,N_5917);
nand U6097 (N_6097,N_5991,N_5896);
nand U6098 (N_6098,N_5891,N_5864);
or U6099 (N_6099,N_5828,N_5860);
and U6100 (N_6100,N_5914,N_5953);
xnor U6101 (N_6101,N_5925,N_5959);
xnor U6102 (N_6102,N_5882,N_5877);
and U6103 (N_6103,N_5889,N_5965);
nor U6104 (N_6104,N_5904,N_5990);
nor U6105 (N_6105,N_5928,N_5955);
or U6106 (N_6106,N_5976,N_5857);
nand U6107 (N_6107,N_5877,N_5981);
xor U6108 (N_6108,N_5981,N_5929);
and U6109 (N_6109,N_5841,N_5913);
nand U6110 (N_6110,N_5853,N_5912);
or U6111 (N_6111,N_5899,N_5908);
nor U6112 (N_6112,N_5928,N_5992);
nand U6113 (N_6113,N_5919,N_5835);
or U6114 (N_6114,N_5860,N_5867);
or U6115 (N_6115,N_5875,N_5804);
or U6116 (N_6116,N_5865,N_5978);
nor U6117 (N_6117,N_5949,N_5833);
nand U6118 (N_6118,N_5983,N_5891);
and U6119 (N_6119,N_5851,N_5862);
nand U6120 (N_6120,N_5824,N_5831);
and U6121 (N_6121,N_5912,N_5953);
or U6122 (N_6122,N_5905,N_5879);
xnor U6123 (N_6123,N_5870,N_5803);
nor U6124 (N_6124,N_5937,N_5882);
and U6125 (N_6125,N_5937,N_5945);
or U6126 (N_6126,N_5810,N_5813);
nand U6127 (N_6127,N_5803,N_5914);
and U6128 (N_6128,N_5986,N_5823);
xnor U6129 (N_6129,N_5925,N_5806);
nor U6130 (N_6130,N_5917,N_5827);
or U6131 (N_6131,N_5965,N_5816);
and U6132 (N_6132,N_5812,N_5861);
and U6133 (N_6133,N_5836,N_5885);
nor U6134 (N_6134,N_5809,N_5914);
xnor U6135 (N_6135,N_5925,N_5901);
nand U6136 (N_6136,N_5894,N_5827);
nand U6137 (N_6137,N_5802,N_5805);
and U6138 (N_6138,N_5950,N_5983);
nand U6139 (N_6139,N_5920,N_5942);
nor U6140 (N_6140,N_5868,N_5976);
xor U6141 (N_6141,N_5895,N_5977);
xor U6142 (N_6142,N_5998,N_5935);
nand U6143 (N_6143,N_5983,N_5864);
nor U6144 (N_6144,N_5997,N_5849);
nor U6145 (N_6145,N_5980,N_5994);
nand U6146 (N_6146,N_5923,N_5801);
xnor U6147 (N_6147,N_5806,N_5899);
nor U6148 (N_6148,N_5917,N_5842);
xor U6149 (N_6149,N_5840,N_5923);
nor U6150 (N_6150,N_5912,N_5906);
xor U6151 (N_6151,N_5976,N_5947);
nor U6152 (N_6152,N_5807,N_5894);
and U6153 (N_6153,N_5986,N_5872);
or U6154 (N_6154,N_5804,N_5867);
nand U6155 (N_6155,N_5831,N_5822);
nand U6156 (N_6156,N_5877,N_5813);
nand U6157 (N_6157,N_5984,N_5852);
nor U6158 (N_6158,N_5928,N_5906);
xnor U6159 (N_6159,N_5870,N_5867);
and U6160 (N_6160,N_5874,N_5882);
xor U6161 (N_6161,N_5960,N_5985);
xor U6162 (N_6162,N_5810,N_5822);
or U6163 (N_6163,N_5863,N_5856);
nand U6164 (N_6164,N_5800,N_5940);
nor U6165 (N_6165,N_5836,N_5978);
and U6166 (N_6166,N_5857,N_5930);
nor U6167 (N_6167,N_5840,N_5812);
xor U6168 (N_6168,N_5931,N_5906);
nand U6169 (N_6169,N_5889,N_5830);
nand U6170 (N_6170,N_5815,N_5820);
xor U6171 (N_6171,N_5851,N_5921);
nand U6172 (N_6172,N_5845,N_5959);
nor U6173 (N_6173,N_5824,N_5843);
and U6174 (N_6174,N_5883,N_5892);
and U6175 (N_6175,N_5991,N_5897);
or U6176 (N_6176,N_5851,N_5941);
xor U6177 (N_6177,N_5833,N_5933);
or U6178 (N_6178,N_5953,N_5964);
nand U6179 (N_6179,N_5926,N_5843);
or U6180 (N_6180,N_5920,N_5944);
nand U6181 (N_6181,N_5948,N_5991);
and U6182 (N_6182,N_5837,N_5926);
and U6183 (N_6183,N_5955,N_5906);
nand U6184 (N_6184,N_5894,N_5820);
or U6185 (N_6185,N_5979,N_5908);
nor U6186 (N_6186,N_5960,N_5926);
xor U6187 (N_6187,N_5926,N_5800);
and U6188 (N_6188,N_5831,N_5845);
nor U6189 (N_6189,N_5867,N_5958);
xor U6190 (N_6190,N_5982,N_5853);
nand U6191 (N_6191,N_5920,N_5822);
xor U6192 (N_6192,N_5938,N_5890);
and U6193 (N_6193,N_5980,N_5894);
xor U6194 (N_6194,N_5928,N_5897);
nor U6195 (N_6195,N_5936,N_5914);
and U6196 (N_6196,N_5872,N_5842);
or U6197 (N_6197,N_5830,N_5918);
xnor U6198 (N_6198,N_5810,N_5840);
or U6199 (N_6199,N_5814,N_5819);
xor U6200 (N_6200,N_6177,N_6079);
xnor U6201 (N_6201,N_6111,N_6087);
nor U6202 (N_6202,N_6114,N_6071);
and U6203 (N_6203,N_6026,N_6005);
nand U6204 (N_6204,N_6162,N_6044);
nor U6205 (N_6205,N_6067,N_6041);
nand U6206 (N_6206,N_6115,N_6070);
nor U6207 (N_6207,N_6133,N_6054);
or U6208 (N_6208,N_6091,N_6003);
and U6209 (N_6209,N_6029,N_6163);
xnor U6210 (N_6210,N_6009,N_6098);
nand U6211 (N_6211,N_6117,N_6051);
nor U6212 (N_6212,N_6132,N_6097);
xnor U6213 (N_6213,N_6096,N_6072);
nand U6214 (N_6214,N_6088,N_6123);
nand U6215 (N_6215,N_6021,N_6170);
and U6216 (N_6216,N_6038,N_6167);
nand U6217 (N_6217,N_6083,N_6049);
xnor U6218 (N_6218,N_6158,N_6105);
or U6219 (N_6219,N_6034,N_6090);
nand U6220 (N_6220,N_6145,N_6122);
nor U6221 (N_6221,N_6025,N_6116);
nand U6222 (N_6222,N_6140,N_6064);
and U6223 (N_6223,N_6012,N_6135);
xor U6224 (N_6224,N_6148,N_6171);
xnor U6225 (N_6225,N_6164,N_6166);
xor U6226 (N_6226,N_6196,N_6042);
nand U6227 (N_6227,N_6010,N_6008);
or U6228 (N_6228,N_6182,N_6048);
nand U6229 (N_6229,N_6121,N_6033);
nand U6230 (N_6230,N_6022,N_6094);
nor U6231 (N_6231,N_6059,N_6195);
nand U6232 (N_6232,N_6173,N_6189);
and U6233 (N_6233,N_6018,N_6153);
nand U6234 (N_6234,N_6134,N_6046);
or U6235 (N_6235,N_6076,N_6032);
xor U6236 (N_6236,N_6047,N_6027);
nor U6237 (N_6237,N_6089,N_6178);
or U6238 (N_6238,N_6040,N_6118);
xnor U6239 (N_6239,N_6077,N_6084);
xor U6240 (N_6240,N_6110,N_6066);
nand U6241 (N_6241,N_6000,N_6169);
and U6242 (N_6242,N_6053,N_6081);
xor U6243 (N_6243,N_6001,N_6131);
or U6244 (N_6244,N_6073,N_6113);
nor U6245 (N_6245,N_6043,N_6057);
or U6246 (N_6246,N_6139,N_6062);
xnor U6247 (N_6247,N_6128,N_6108);
nand U6248 (N_6248,N_6037,N_6102);
nor U6249 (N_6249,N_6172,N_6011);
nand U6250 (N_6250,N_6179,N_6138);
nand U6251 (N_6251,N_6156,N_6058);
xnor U6252 (N_6252,N_6019,N_6099);
nor U6253 (N_6253,N_6017,N_6020);
nand U6254 (N_6254,N_6186,N_6106);
or U6255 (N_6255,N_6126,N_6095);
nor U6256 (N_6256,N_6119,N_6112);
nand U6257 (N_6257,N_6100,N_6143);
xor U6258 (N_6258,N_6154,N_6120);
and U6259 (N_6259,N_6176,N_6183);
or U6260 (N_6260,N_6074,N_6002);
and U6261 (N_6261,N_6109,N_6060);
xor U6262 (N_6262,N_6146,N_6157);
and U6263 (N_6263,N_6104,N_6069);
xor U6264 (N_6264,N_6006,N_6150);
xnor U6265 (N_6265,N_6129,N_6015);
xor U6266 (N_6266,N_6082,N_6155);
xor U6267 (N_6267,N_6192,N_6004);
and U6268 (N_6268,N_6013,N_6039);
nand U6269 (N_6269,N_6050,N_6152);
nand U6270 (N_6270,N_6107,N_6068);
nand U6271 (N_6271,N_6103,N_6188);
xor U6272 (N_6272,N_6144,N_6194);
nand U6273 (N_6273,N_6045,N_6080);
or U6274 (N_6274,N_6198,N_6078);
xor U6275 (N_6275,N_6190,N_6030);
and U6276 (N_6276,N_6055,N_6165);
and U6277 (N_6277,N_6056,N_6185);
and U6278 (N_6278,N_6136,N_6007);
nor U6279 (N_6279,N_6160,N_6197);
nor U6280 (N_6280,N_6149,N_6101);
or U6281 (N_6281,N_6085,N_6024);
xor U6282 (N_6282,N_6187,N_6065);
and U6283 (N_6283,N_6191,N_6125);
nand U6284 (N_6284,N_6052,N_6061);
or U6285 (N_6285,N_6174,N_6016);
nor U6286 (N_6286,N_6075,N_6124);
or U6287 (N_6287,N_6147,N_6142);
xnor U6288 (N_6288,N_6181,N_6175);
or U6289 (N_6289,N_6130,N_6093);
nor U6290 (N_6290,N_6063,N_6180);
nor U6291 (N_6291,N_6036,N_6199);
or U6292 (N_6292,N_6127,N_6023);
xnor U6293 (N_6293,N_6086,N_6151);
xnor U6294 (N_6294,N_6168,N_6184);
and U6295 (N_6295,N_6161,N_6092);
nor U6296 (N_6296,N_6193,N_6014);
xnor U6297 (N_6297,N_6141,N_6035);
nor U6298 (N_6298,N_6031,N_6159);
xnor U6299 (N_6299,N_6028,N_6137);
and U6300 (N_6300,N_6123,N_6192);
nand U6301 (N_6301,N_6082,N_6132);
or U6302 (N_6302,N_6156,N_6108);
nor U6303 (N_6303,N_6101,N_6058);
nand U6304 (N_6304,N_6014,N_6062);
nor U6305 (N_6305,N_6050,N_6145);
xor U6306 (N_6306,N_6028,N_6062);
xor U6307 (N_6307,N_6187,N_6013);
nor U6308 (N_6308,N_6000,N_6182);
xnor U6309 (N_6309,N_6045,N_6193);
nor U6310 (N_6310,N_6170,N_6002);
nor U6311 (N_6311,N_6153,N_6098);
nand U6312 (N_6312,N_6057,N_6073);
and U6313 (N_6313,N_6029,N_6125);
nor U6314 (N_6314,N_6165,N_6169);
and U6315 (N_6315,N_6174,N_6025);
xor U6316 (N_6316,N_6094,N_6037);
nand U6317 (N_6317,N_6115,N_6024);
and U6318 (N_6318,N_6072,N_6140);
xor U6319 (N_6319,N_6012,N_6027);
nor U6320 (N_6320,N_6115,N_6061);
and U6321 (N_6321,N_6110,N_6121);
or U6322 (N_6322,N_6112,N_6067);
nand U6323 (N_6323,N_6172,N_6091);
or U6324 (N_6324,N_6142,N_6103);
xor U6325 (N_6325,N_6011,N_6010);
xor U6326 (N_6326,N_6107,N_6141);
xor U6327 (N_6327,N_6020,N_6154);
nand U6328 (N_6328,N_6180,N_6119);
nand U6329 (N_6329,N_6112,N_6104);
nor U6330 (N_6330,N_6197,N_6147);
xor U6331 (N_6331,N_6040,N_6171);
xnor U6332 (N_6332,N_6107,N_6189);
nor U6333 (N_6333,N_6166,N_6118);
nor U6334 (N_6334,N_6188,N_6184);
nand U6335 (N_6335,N_6123,N_6143);
and U6336 (N_6336,N_6014,N_6103);
and U6337 (N_6337,N_6064,N_6004);
xnor U6338 (N_6338,N_6037,N_6078);
or U6339 (N_6339,N_6170,N_6011);
or U6340 (N_6340,N_6104,N_6132);
xnor U6341 (N_6341,N_6122,N_6133);
or U6342 (N_6342,N_6087,N_6019);
xor U6343 (N_6343,N_6087,N_6069);
nand U6344 (N_6344,N_6128,N_6182);
or U6345 (N_6345,N_6092,N_6075);
and U6346 (N_6346,N_6008,N_6004);
and U6347 (N_6347,N_6132,N_6153);
nor U6348 (N_6348,N_6165,N_6120);
nand U6349 (N_6349,N_6062,N_6117);
nand U6350 (N_6350,N_6004,N_6024);
nand U6351 (N_6351,N_6037,N_6199);
nand U6352 (N_6352,N_6138,N_6094);
xor U6353 (N_6353,N_6175,N_6100);
and U6354 (N_6354,N_6113,N_6020);
nand U6355 (N_6355,N_6198,N_6062);
nor U6356 (N_6356,N_6042,N_6001);
and U6357 (N_6357,N_6169,N_6154);
nor U6358 (N_6358,N_6188,N_6169);
and U6359 (N_6359,N_6182,N_6104);
xnor U6360 (N_6360,N_6023,N_6093);
or U6361 (N_6361,N_6164,N_6160);
and U6362 (N_6362,N_6034,N_6040);
nand U6363 (N_6363,N_6159,N_6094);
or U6364 (N_6364,N_6183,N_6136);
and U6365 (N_6365,N_6101,N_6031);
and U6366 (N_6366,N_6093,N_6013);
or U6367 (N_6367,N_6014,N_6033);
xnor U6368 (N_6368,N_6185,N_6005);
and U6369 (N_6369,N_6018,N_6170);
nor U6370 (N_6370,N_6041,N_6072);
xnor U6371 (N_6371,N_6074,N_6000);
or U6372 (N_6372,N_6002,N_6027);
nand U6373 (N_6373,N_6185,N_6067);
and U6374 (N_6374,N_6124,N_6186);
nor U6375 (N_6375,N_6028,N_6080);
nor U6376 (N_6376,N_6129,N_6178);
xor U6377 (N_6377,N_6092,N_6085);
or U6378 (N_6378,N_6051,N_6025);
or U6379 (N_6379,N_6179,N_6144);
xnor U6380 (N_6380,N_6075,N_6091);
nand U6381 (N_6381,N_6148,N_6105);
xnor U6382 (N_6382,N_6197,N_6095);
or U6383 (N_6383,N_6186,N_6133);
nor U6384 (N_6384,N_6110,N_6080);
nor U6385 (N_6385,N_6015,N_6168);
xnor U6386 (N_6386,N_6053,N_6101);
nand U6387 (N_6387,N_6086,N_6141);
and U6388 (N_6388,N_6113,N_6169);
and U6389 (N_6389,N_6117,N_6053);
xnor U6390 (N_6390,N_6124,N_6192);
nand U6391 (N_6391,N_6026,N_6123);
and U6392 (N_6392,N_6152,N_6001);
nor U6393 (N_6393,N_6005,N_6119);
xnor U6394 (N_6394,N_6102,N_6018);
nor U6395 (N_6395,N_6119,N_6139);
nor U6396 (N_6396,N_6129,N_6049);
xnor U6397 (N_6397,N_6070,N_6150);
xnor U6398 (N_6398,N_6094,N_6043);
xnor U6399 (N_6399,N_6160,N_6138);
nand U6400 (N_6400,N_6268,N_6265);
nor U6401 (N_6401,N_6296,N_6360);
and U6402 (N_6402,N_6217,N_6373);
and U6403 (N_6403,N_6233,N_6229);
or U6404 (N_6404,N_6234,N_6276);
xor U6405 (N_6405,N_6204,N_6330);
or U6406 (N_6406,N_6374,N_6208);
nor U6407 (N_6407,N_6206,N_6361);
nor U6408 (N_6408,N_6307,N_6396);
nor U6409 (N_6409,N_6242,N_6272);
nor U6410 (N_6410,N_6212,N_6261);
nor U6411 (N_6411,N_6209,N_6291);
and U6412 (N_6412,N_6326,N_6294);
nor U6413 (N_6413,N_6375,N_6232);
xnor U6414 (N_6414,N_6200,N_6213);
nand U6415 (N_6415,N_6335,N_6344);
nor U6416 (N_6416,N_6301,N_6399);
xor U6417 (N_6417,N_6304,N_6219);
and U6418 (N_6418,N_6257,N_6271);
or U6419 (N_6419,N_6231,N_6324);
xor U6420 (N_6420,N_6255,N_6349);
and U6421 (N_6421,N_6220,N_6273);
xor U6422 (N_6422,N_6207,N_6252);
and U6423 (N_6423,N_6286,N_6254);
nand U6424 (N_6424,N_6394,N_6302);
or U6425 (N_6425,N_6323,N_6318);
xnor U6426 (N_6426,N_6211,N_6227);
nor U6427 (N_6427,N_6263,N_6228);
nand U6428 (N_6428,N_6230,N_6262);
and U6429 (N_6429,N_6292,N_6325);
and U6430 (N_6430,N_6285,N_6300);
nand U6431 (N_6431,N_6346,N_6366);
nand U6432 (N_6432,N_6266,N_6303);
or U6433 (N_6433,N_6202,N_6372);
and U6434 (N_6434,N_6218,N_6259);
xor U6435 (N_6435,N_6389,N_6369);
or U6436 (N_6436,N_6215,N_6336);
or U6437 (N_6437,N_6249,N_6363);
and U6438 (N_6438,N_6264,N_6226);
and U6439 (N_6439,N_6310,N_6332);
or U6440 (N_6440,N_6327,N_6260);
or U6441 (N_6441,N_6224,N_6378);
nor U6442 (N_6442,N_6253,N_6290);
nor U6443 (N_6443,N_6312,N_6392);
or U6444 (N_6444,N_6376,N_6250);
nor U6445 (N_6445,N_6240,N_6279);
nand U6446 (N_6446,N_6222,N_6345);
nand U6447 (N_6447,N_6289,N_6277);
and U6448 (N_6448,N_6306,N_6316);
and U6449 (N_6449,N_6241,N_6239);
or U6450 (N_6450,N_6317,N_6393);
nand U6451 (N_6451,N_6319,N_6334);
xor U6452 (N_6452,N_6367,N_6347);
or U6453 (N_6453,N_6371,N_6269);
nor U6454 (N_6454,N_6390,N_6362);
xnor U6455 (N_6455,N_6275,N_6343);
nor U6456 (N_6456,N_6225,N_6237);
and U6457 (N_6457,N_6246,N_6256);
nand U6458 (N_6458,N_6337,N_6270);
nand U6459 (N_6459,N_6288,N_6247);
nor U6460 (N_6460,N_6251,N_6315);
nor U6461 (N_6461,N_6358,N_6287);
nand U6462 (N_6462,N_6383,N_6221);
xor U6463 (N_6463,N_6258,N_6329);
nor U6464 (N_6464,N_6314,N_6340);
or U6465 (N_6465,N_6210,N_6278);
or U6466 (N_6466,N_6380,N_6235);
or U6467 (N_6467,N_6320,N_6243);
or U6468 (N_6468,N_6350,N_6395);
xor U6469 (N_6469,N_6223,N_6384);
nand U6470 (N_6470,N_6348,N_6398);
xnor U6471 (N_6471,N_6352,N_6311);
nor U6472 (N_6472,N_6391,N_6297);
or U6473 (N_6473,N_6322,N_6245);
nor U6474 (N_6474,N_6248,N_6370);
xor U6475 (N_6475,N_6355,N_6201);
nand U6476 (N_6476,N_6244,N_6293);
and U6477 (N_6477,N_6341,N_6216);
nand U6478 (N_6478,N_6354,N_6282);
and U6479 (N_6479,N_6353,N_6357);
nor U6480 (N_6480,N_6313,N_6281);
or U6481 (N_6481,N_6342,N_6379);
and U6482 (N_6482,N_6205,N_6267);
or U6483 (N_6483,N_6386,N_6356);
nand U6484 (N_6484,N_6280,N_6236);
and U6485 (N_6485,N_6397,N_6321);
xor U6486 (N_6486,N_6203,N_6339);
and U6487 (N_6487,N_6238,N_6364);
xnor U6488 (N_6488,N_6385,N_6328);
nand U6489 (N_6489,N_6331,N_6284);
and U6490 (N_6490,N_6381,N_6308);
or U6491 (N_6491,N_6333,N_6295);
or U6492 (N_6492,N_6351,N_6274);
or U6493 (N_6493,N_6359,N_6298);
nand U6494 (N_6494,N_6338,N_6309);
nand U6495 (N_6495,N_6388,N_6365);
nor U6496 (N_6496,N_6299,N_6387);
or U6497 (N_6497,N_6377,N_6305);
nand U6498 (N_6498,N_6382,N_6214);
nor U6499 (N_6499,N_6368,N_6283);
nand U6500 (N_6500,N_6254,N_6317);
nand U6501 (N_6501,N_6354,N_6226);
nand U6502 (N_6502,N_6396,N_6315);
and U6503 (N_6503,N_6384,N_6282);
nor U6504 (N_6504,N_6240,N_6306);
nor U6505 (N_6505,N_6327,N_6323);
nor U6506 (N_6506,N_6209,N_6274);
nand U6507 (N_6507,N_6365,N_6342);
nor U6508 (N_6508,N_6255,N_6210);
nor U6509 (N_6509,N_6374,N_6220);
xor U6510 (N_6510,N_6221,N_6360);
or U6511 (N_6511,N_6223,N_6372);
xor U6512 (N_6512,N_6216,N_6328);
xnor U6513 (N_6513,N_6289,N_6398);
nor U6514 (N_6514,N_6387,N_6342);
or U6515 (N_6515,N_6335,N_6323);
and U6516 (N_6516,N_6277,N_6340);
xnor U6517 (N_6517,N_6275,N_6391);
and U6518 (N_6518,N_6355,N_6306);
xor U6519 (N_6519,N_6361,N_6228);
nand U6520 (N_6520,N_6235,N_6232);
nor U6521 (N_6521,N_6284,N_6380);
and U6522 (N_6522,N_6291,N_6342);
nor U6523 (N_6523,N_6368,N_6202);
and U6524 (N_6524,N_6313,N_6245);
nand U6525 (N_6525,N_6206,N_6207);
nor U6526 (N_6526,N_6278,N_6388);
nor U6527 (N_6527,N_6201,N_6261);
nand U6528 (N_6528,N_6368,N_6323);
nand U6529 (N_6529,N_6284,N_6292);
nor U6530 (N_6530,N_6365,N_6241);
nand U6531 (N_6531,N_6345,N_6391);
or U6532 (N_6532,N_6243,N_6271);
or U6533 (N_6533,N_6220,N_6348);
and U6534 (N_6534,N_6305,N_6244);
nor U6535 (N_6535,N_6316,N_6209);
nor U6536 (N_6536,N_6235,N_6281);
xor U6537 (N_6537,N_6273,N_6211);
and U6538 (N_6538,N_6313,N_6209);
nor U6539 (N_6539,N_6211,N_6394);
xnor U6540 (N_6540,N_6244,N_6295);
nor U6541 (N_6541,N_6202,N_6325);
nor U6542 (N_6542,N_6238,N_6318);
and U6543 (N_6543,N_6232,N_6284);
nor U6544 (N_6544,N_6311,N_6371);
or U6545 (N_6545,N_6278,N_6318);
nor U6546 (N_6546,N_6333,N_6366);
or U6547 (N_6547,N_6266,N_6212);
and U6548 (N_6548,N_6331,N_6249);
nor U6549 (N_6549,N_6282,N_6281);
nor U6550 (N_6550,N_6385,N_6214);
nor U6551 (N_6551,N_6340,N_6354);
xnor U6552 (N_6552,N_6253,N_6233);
or U6553 (N_6553,N_6339,N_6326);
nand U6554 (N_6554,N_6257,N_6242);
nor U6555 (N_6555,N_6307,N_6391);
xor U6556 (N_6556,N_6230,N_6368);
or U6557 (N_6557,N_6330,N_6289);
xor U6558 (N_6558,N_6230,N_6247);
nand U6559 (N_6559,N_6374,N_6299);
or U6560 (N_6560,N_6287,N_6361);
and U6561 (N_6561,N_6360,N_6229);
xor U6562 (N_6562,N_6236,N_6248);
and U6563 (N_6563,N_6284,N_6254);
and U6564 (N_6564,N_6320,N_6354);
xor U6565 (N_6565,N_6360,N_6267);
nand U6566 (N_6566,N_6300,N_6269);
or U6567 (N_6567,N_6344,N_6326);
nor U6568 (N_6568,N_6337,N_6392);
xor U6569 (N_6569,N_6217,N_6371);
or U6570 (N_6570,N_6237,N_6317);
or U6571 (N_6571,N_6359,N_6382);
nor U6572 (N_6572,N_6309,N_6316);
nand U6573 (N_6573,N_6398,N_6318);
or U6574 (N_6574,N_6241,N_6207);
and U6575 (N_6575,N_6349,N_6332);
or U6576 (N_6576,N_6279,N_6377);
xnor U6577 (N_6577,N_6398,N_6389);
xor U6578 (N_6578,N_6210,N_6392);
xnor U6579 (N_6579,N_6214,N_6254);
xnor U6580 (N_6580,N_6238,N_6243);
nand U6581 (N_6581,N_6280,N_6253);
xnor U6582 (N_6582,N_6353,N_6392);
and U6583 (N_6583,N_6203,N_6357);
and U6584 (N_6584,N_6278,N_6225);
or U6585 (N_6585,N_6238,N_6323);
and U6586 (N_6586,N_6391,N_6251);
and U6587 (N_6587,N_6214,N_6396);
nand U6588 (N_6588,N_6320,N_6387);
xor U6589 (N_6589,N_6252,N_6382);
nor U6590 (N_6590,N_6311,N_6284);
nand U6591 (N_6591,N_6307,N_6315);
nor U6592 (N_6592,N_6350,N_6291);
nand U6593 (N_6593,N_6345,N_6375);
or U6594 (N_6594,N_6367,N_6212);
xor U6595 (N_6595,N_6222,N_6212);
or U6596 (N_6596,N_6348,N_6296);
nand U6597 (N_6597,N_6348,N_6332);
xnor U6598 (N_6598,N_6386,N_6395);
nor U6599 (N_6599,N_6348,N_6202);
or U6600 (N_6600,N_6526,N_6524);
xor U6601 (N_6601,N_6588,N_6574);
and U6602 (N_6602,N_6506,N_6494);
nor U6603 (N_6603,N_6453,N_6587);
xnor U6604 (N_6604,N_6468,N_6551);
and U6605 (N_6605,N_6461,N_6420);
and U6606 (N_6606,N_6415,N_6408);
and U6607 (N_6607,N_6573,N_6424);
or U6608 (N_6608,N_6592,N_6417);
xnor U6609 (N_6609,N_6426,N_6463);
nand U6610 (N_6610,N_6473,N_6590);
nand U6611 (N_6611,N_6513,N_6517);
nand U6612 (N_6612,N_6534,N_6540);
nor U6613 (N_6613,N_6501,N_6432);
xor U6614 (N_6614,N_6570,N_6509);
or U6615 (N_6615,N_6487,N_6403);
nand U6616 (N_6616,N_6446,N_6455);
xnor U6617 (N_6617,N_6401,N_6405);
nor U6618 (N_6618,N_6596,N_6423);
xnor U6619 (N_6619,N_6488,N_6482);
or U6620 (N_6620,N_6560,N_6436);
and U6621 (N_6621,N_6476,N_6443);
and U6622 (N_6622,N_6594,N_6537);
nor U6623 (N_6623,N_6456,N_6515);
xnor U6624 (N_6624,N_6445,N_6581);
or U6625 (N_6625,N_6421,N_6577);
xor U6626 (N_6626,N_6410,N_6564);
xnor U6627 (N_6627,N_6505,N_6585);
nand U6628 (N_6628,N_6595,N_6532);
nand U6629 (N_6629,N_6498,N_6460);
nor U6630 (N_6630,N_6510,N_6580);
nand U6631 (N_6631,N_6583,N_6449);
and U6632 (N_6632,N_6496,N_6416);
nand U6633 (N_6633,N_6550,N_6531);
nor U6634 (N_6634,N_6520,N_6504);
and U6635 (N_6635,N_6589,N_6427);
or U6636 (N_6636,N_6434,N_6459);
and U6637 (N_6637,N_6544,N_6452);
or U6638 (N_6638,N_6500,N_6447);
nand U6639 (N_6639,N_6441,N_6430);
or U6640 (N_6640,N_6571,N_6565);
or U6641 (N_6641,N_6419,N_6418);
xnor U6642 (N_6642,N_6439,N_6562);
or U6643 (N_6643,N_6527,N_6507);
nor U6644 (N_6644,N_6425,N_6539);
nor U6645 (N_6645,N_6413,N_6518);
nor U6646 (N_6646,N_6475,N_6428);
and U6647 (N_6647,N_6516,N_6591);
or U6648 (N_6648,N_6542,N_6598);
xor U6649 (N_6649,N_6549,N_6490);
and U6650 (N_6650,N_6559,N_6552);
and U6651 (N_6651,N_6554,N_6533);
nor U6652 (N_6652,N_6512,N_6569);
nand U6653 (N_6653,N_6438,N_6566);
or U6654 (N_6654,N_6572,N_6511);
and U6655 (N_6655,N_6508,N_6404);
or U6656 (N_6656,N_6450,N_6499);
xnor U6657 (N_6657,N_6458,N_6502);
nand U6658 (N_6658,N_6529,N_6448);
xnor U6659 (N_6659,N_6547,N_6546);
and U6660 (N_6660,N_6422,N_6462);
and U6661 (N_6661,N_6479,N_6567);
or U6662 (N_6662,N_6480,N_6470);
xnor U6663 (N_6663,N_6525,N_6535);
nand U6664 (N_6664,N_6451,N_6530);
nor U6665 (N_6665,N_6582,N_6429);
xnor U6666 (N_6666,N_6521,N_6556);
nand U6667 (N_6667,N_6483,N_6599);
xor U6668 (N_6668,N_6523,N_6486);
or U6669 (N_6669,N_6503,N_6561);
xor U6670 (N_6670,N_6522,N_6548);
nor U6671 (N_6671,N_6444,N_6440);
or U6672 (N_6672,N_6497,N_6514);
and U6673 (N_6673,N_6563,N_6584);
xor U6674 (N_6674,N_6545,N_6491);
and U6675 (N_6675,N_6400,N_6579);
nor U6676 (N_6676,N_6536,N_6412);
and U6677 (N_6677,N_6465,N_6492);
and U6678 (N_6678,N_6578,N_6469);
or U6679 (N_6679,N_6407,N_6457);
and U6680 (N_6680,N_6485,N_6568);
and U6681 (N_6681,N_6555,N_6484);
nor U6682 (N_6682,N_6543,N_6402);
and U6683 (N_6683,N_6528,N_6467);
nor U6684 (N_6684,N_6409,N_6454);
xor U6685 (N_6685,N_6466,N_6433);
nor U6686 (N_6686,N_6541,N_6414);
nor U6687 (N_6687,N_6593,N_6575);
nand U6688 (N_6688,N_6478,N_6411);
nand U6689 (N_6689,N_6495,N_6558);
and U6690 (N_6690,N_6435,N_6474);
or U6691 (N_6691,N_6597,N_6553);
or U6692 (N_6692,N_6489,N_6493);
and U6693 (N_6693,N_6471,N_6586);
xnor U6694 (N_6694,N_6538,N_6472);
and U6695 (N_6695,N_6481,N_6406);
or U6696 (N_6696,N_6557,N_6442);
xnor U6697 (N_6697,N_6464,N_6431);
and U6698 (N_6698,N_6437,N_6519);
or U6699 (N_6699,N_6477,N_6576);
or U6700 (N_6700,N_6548,N_6443);
nand U6701 (N_6701,N_6542,N_6506);
xnor U6702 (N_6702,N_6446,N_6464);
nor U6703 (N_6703,N_6595,N_6437);
nand U6704 (N_6704,N_6539,N_6414);
or U6705 (N_6705,N_6480,N_6424);
xnor U6706 (N_6706,N_6401,N_6465);
or U6707 (N_6707,N_6492,N_6472);
nor U6708 (N_6708,N_6598,N_6565);
and U6709 (N_6709,N_6545,N_6441);
and U6710 (N_6710,N_6415,N_6580);
or U6711 (N_6711,N_6513,N_6424);
xor U6712 (N_6712,N_6411,N_6474);
and U6713 (N_6713,N_6559,N_6505);
nand U6714 (N_6714,N_6526,N_6416);
and U6715 (N_6715,N_6599,N_6406);
xor U6716 (N_6716,N_6540,N_6524);
or U6717 (N_6717,N_6439,N_6598);
xor U6718 (N_6718,N_6421,N_6550);
nand U6719 (N_6719,N_6454,N_6574);
or U6720 (N_6720,N_6581,N_6595);
nand U6721 (N_6721,N_6549,N_6410);
and U6722 (N_6722,N_6567,N_6594);
nand U6723 (N_6723,N_6537,N_6541);
nor U6724 (N_6724,N_6446,N_6426);
and U6725 (N_6725,N_6497,N_6549);
and U6726 (N_6726,N_6552,N_6445);
nand U6727 (N_6727,N_6516,N_6506);
nand U6728 (N_6728,N_6421,N_6407);
nand U6729 (N_6729,N_6530,N_6472);
nor U6730 (N_6730,N_6541,N_6515);
xnor U6731 (N_6731,N_6462,N_6554);
or U6732 (N_6732,N_6453,N_6501);
xor U6733 (N_6733,N_6424,N_6559);
or U6734 (N_6734,N_6561,N_6474);
or U6735 (N_6735,N_6484,N_6464);
or U6736 (N_6736,N_6473,N_6424);
and U6737 (N_6737,N_6552,N_6428);
xor U6738 (N_6738,N_6569,N_6413);
nand U6739 (N_6739,N_6481,N_6403);
or U6740 (N_6740,N_6439,N_6557);
nor U6741 (N_6741,N_6587,N_6553);
and U6742 (N_6742,N_6513,N_6512);
and U6743 (N_6743,N_6555,N_6584);
nand U6744 (N_6744,N_6509,N_6581);
and U6745 (N_6745,N_6532,N_6588);
nand U6746 (N_6746,N_6566,N_6464);
or U6747 (N_6747,N_6422,N_6596);
nor U6748 (N_6748,N_6423,N_6536);
and U6749 (N_6749,N_6432,N_6438);
nor U6750 (N_6750,N_6561,N_6497);
or U6751 (N_6751,N_6553,N_6404);
nand U6752 (N_6752,N_6592,N_6508);
xor U6753 (N_6753,N_6482,N_6484);
nor U6754 (N_6754,N_6521,N_6465);
or U6755 (N_6755,N_6480,N_6528);
xnor U6756 (N_6756,N_6556,N_6446);
or U6757 (N_6757,N_6597,N_6562);
and U6758 (N_6758,N_6409,N_6493);
or U6759 (N_6759,N_6515,N_6559);
nand U6760 (N_6760,N_6440,N_6579);
or U6761 (N_6761,N_6511,N_6555);
nand U6762 (N_6762,N_6412,N_6472);
and U6763 (N_6763,N_6447,N_6574);
or U6764 (N_6764,N_6440,N_6582);
xor U6765 (N_6765,N_6439,N_6414);
nand U6766 (N_6766,N_6572,N_6472);
nor U6767 (N_6767,N_6519,N_6568);
and U6768 (N_6768,N_6462,N_6525);
nor U6769 (N_6769,N_6455,N_6581);
and U6770 (N_6770,N_6531,N_6464);
nand U6771 (N_6771,N_6592,N_6436);
nand U6772 (N_6772,N_6546,N_6515);
nand U6773 (N_6773,N_6453,N_6536);
nor U6774 (N_6774,N_6576,N_6561);
and U6775 (N_6775,N_6400,N_6547);
xor U6776 (N_6776,N_6514,N_6504);
xor U6777 (N_6777,N_6407,N_6596);
xnor U6778 (N_6778,N_6546,N_6519);
nand U6779 (N_6779,N_6454,N_6485);
and U6780 (N_6780,N_6468,N_6407);
nor U6781 (N_6781,N_6449,N_6446);
nand U6782 (N_6782,N_6503,N_6506);
nand U6783 (N_6783,N_6549,N_6579);
nor U6784 (N_6784,N_6547,N_6580);
or U6785 (N_6785,N_6587,N_6578);
nand U6786 (N_6786,N_6506,N_6559);
nor U6787 (N_6787,N_6556,N_6596);
nand U6788 (N_6788,N_6464,N_6418);
xnor U6789 (N_6789,N_6404,N_6590);
nor U6790 (N_6790,N_6581,N_6474);
nor U6791 (N_6791,N_6426,N_6400);
and U6792 (N_6792,N_6527,N_6592);
nor U6793 (N_6793,N_6581,N_6471);
or U6794 (N_6794,N_6490,N_6467);
or U6795 (N_6795,N_6433,N_6545);
xnor U6796 (N_6796,N_6467,N_6511);
nand U6797 (N_6797,N_6491,N_6598);
or U6798 (N_6798,N_6463,N_6567);
nand U6799 (N_6799,N_6459,N_6538);
xor U6800 (N_6800,N_6620,N_6738);
nand U6801 (N_6801,N_6607,N_6700);
xor U6802 (N_6802,N_6729,N_6712);
nor U6803 (N_6803,N_6682,N_6716);
and U6804 (N_6804,N_6749,N_6667);
nand U6805 (N_6805,N_6727,N_6675);
nand U6806 (N_6806,N_6775,N_6792);
xnor U6807 (N_6807,N_6782,N_6717);
nor U6808 (N_6808,N_6784,N_6760);
or U6809 (N_6809,N_6646,N_6605);
or U6810 (N_6810,N_6608,N_6707);
nor U6811 (N_6811,N_6691,N_6703);
and U6812 (N_6812,N_6609,N_6614);
nand U6813 (N_6813,N_6699,N_6649);
xnor U6814 (N_6814,N_6690,N_6741);
and U6815 (N_6815,N_6789,N_6721);
xor U6816 (N_6816,N_6602,N_6683);
xnor U6817 (N_6817,N_6610,N_6659);
xnor U6818 (N_6818,N_6632,N_6623);
and U6819 (N_6819,N_6654,N_6704);
nor U6820 (N_6820,N_6677,N_6627);
or U6821 (N_6821,N_6714,N_6655);
nor U6822 (N_6822,N_6747,N_6636);
nor U6823 (N_6823,N_6731,N_6778);
or U6824 (N_6824,N_6656,N_6761);
and U6825 (N_6825,N_6612,N_6722);
nand U6826 (N_6826,N_6743,N_6777);
nand U6827 (N_6827,N_6748,N_6611);
nand U6828 (N_6828,N_6763,N_6668);
nand U6829 (N_6829,N_6658,N_6652);
and U6830 (N_6830,N_6781,N_6637);
nand U6831 (N_6831,N_6757,N_6660);
or U6832 (N_6832,N_6641,N_6693);
nand U6833 (N_6833,N_6679,N_6633);
nand U6834 (N_6834,N_6663,N_6681);
nand U6835 (N_6835,N_6680,N_6732);
and U6836 (N_6836,N_6750,N_6671);
nor U6837 (N_6837,N_6766,N_6715);
or U6838 (N_6838,N_6796,N_6643);
xor U6839 (N_6839,N_6774,N_6689);
xor U6840 (N_6840,N_6711,N_6634);
or U6841 (N_6841,N_6698,N_6669);
nor U6842 (N_6842,N_6769,N_6670);
and U6843 (N_6843,N_6735,N_6780);
or U6844 (N_6844,N_6773,N_6734);
xnor U6845 (N_6845,N_6606,N_6739);
or U6846 (N_6846,N_6710,N_6648);
nand U6847 (N_6847,N_6666,N_6793);
or U6848 (N_6848,N_6752,N_6702);
xnor U6849 (N_6849,N_6708,N_6779);
xnor U6850 (N_6850,N_6754,N_6764);
nand U6851 (N_6851,N_6744,N_6728);
or U6852 (N_6852,N_6687,N_6737);
nand U6853 (N_6853,N_6684,N_6706);
nor U6854 (N_6854,N_6695,N_6650);
nor U6855 (N_6855,N_6613,N_6762);
nor U6856 (N_6856,N_6767,N_6621);
and U6857 (N_6857,N_6628,N_6657);
or U6858 (N_6858,N_6726,N_6644);
nand U6859 (N_6859,N_6746,N_6725);
nor U6860 (N_6860,N_6783,N_6630);
xor U6861 (N_6861,N_6645,N_6616);
or U6862 (N_6862,N_6753,N_6603);
xnor U6863 (N_6863,N_6665,N_6673);
nor U6864 (N_6864,N_6791,N_6758);
and U6865 (N_6865,N_6629,N_6799);
nor U6866 (N_6866,N_6601,N_6709);
xnor U6867 (N_6867,N_6686,N_6697);
nor U6868 (N_6868,N_6730,N_6619);
nor U6869 (N_6869,N_6759,N_6676);
nor U6870 (N_6870,N_6647,N_6639);
nand U6871 (N_6871,N_6776,N_6705);
and U6872 (N_6872,N_6640,N_6622);
and U6873 (N_6873,N_6724,N_6771);
xnor U6874 (N_6874,N_6788,N_6718);
xnor U6875 (N_6875,N_6742,N_6625);
nand U6876 (N_6876,N_6626,N_6794);
xor U6877 (N_6877,N_6790,N_6756);
and U6878 (N_6878,N_6664,N_6785);
nor U6879 (N_6879,N_6642,N_6713);
xor U6880 (N_6880,N_6768,N_6678);
or U6881 (N_6881,N_6662,N_6631);
xnor U6882 (N_6882,N_6618,N_6600);
nor U6883 (N_6883,N_6604,N_6795);
xnor U6884 (N_6884,N_6653,N_6615);
or U6885 (N_6885,N_6798,N_6736);
nor U6886 (N_6886,N_6692,N_6701);
nor U6887 (N_6887,N_6638,N_6772);
or U6888 (N_6888,N_6765,N_6694);
xor U6889 (N_6889,N_6733,N_6688);
or U6890 (N_6890,N_6745,N_6797);
nor U6891 (N_6891,N_6651,N_6740);
nor U6892 (N_6892,N_6770,N_6674);
nand U6893 (N_6893,N_6787,N_6720);
and U6894 (N_6894,N_6751,N_6723);
nor U6895 (N_6895,N_6635,N_6617);
nand U6896 (N_6896,N_6661,N_6672);
xnor U6897 (N_6897,N_6624,N_6755);
nand U6898 (N_6898,N_6696,N_6786);
nand U6899 (N_6899,N_6685,N_6719);
and U6900 (N_6900,N_6719,N_6743);
nor U6901 (N_6901,N_6655,N_6748);
and U6902 (N_6902,N_6729,N_6753);
or U6903 (N_6903,N_6678,N_6747);
or U6904 (N_6904,N_6656,N_6637);
nor U6905 (N_6905,N_6787,N_6723);
or U6906 (N_6906,N_6663,N_6743);
and U6907 (N_6907,N_6723,N_6678);
nand U6908 (N_6908,N_6774,N_6707);
or U6909 (N_6909,N_6785,N_6606);
nand U6910 (N_6910,N_6607,N_6720);
or U6911 (N_6911,N_6657,N_6680);
and U6912 (N_6912,N_6694,N_6781);
and U6913 (N_6913,N_6675,N_6786);
and U6914 (N_6914,N_6794,N_6686);
nand U6915 (N_6915,N_6667,N_6620);
nor U6916 (N_6916,N_6680,N_6652);
nand U6917 (N_6917,N_6758,N_6770);
nor U6918 (N_6918,N_6674,N_6645);
nor U6919 (N_6919,N_6648,N_6690);
xor U6920 (N_6920,N_6629,N_6705);
nand U6921 (N_6921,N_6661,N_6667);
or U6922 (N_6922,N_6677,N_6617);
xor U6923 (N_6923,N_6658,N_6751);
nor U6924 (N_6924,N_6709,N_6728);
and U6925 (N_6925,N_6605,N_6743);
or U6926 (N_6926,N_6640,N_6752);
nor U6927 (N_6927,N_6721,N_6791);
xnor U6928 (N_6928,N_6753,N_6715);
or U6929 (N_6929,N_6648,N_6746);
and U6930 (N_6930,N_6789,N_6686);
nor U6931 (N_6931,N_6799,N_6641);
nor U6932 (N_6932,N_6620,N_6720);
and U6933 (N_6933,N_6707,N_6776);
nand U6934 (N_6934,N_6670,N_6673);
xnor U6935 (N_6935,N_6666,N_6764);
or U6936 (N_6936,N_6731,N_6746);
and U6937 (N_6937,N_6649,N_6654);
or U6938 (N_6938,N_6653,N_6703);
or U6939 (N_6939,N_6676,N_6762);
nand U6940 (N_6940,N_6681,N_6700);
or U6941 (N_6941,N_6633,N_6667);
and U6942 (N_6942,N_6744,N_6652);
or U6943 (N_6943,N_6737,N_6782);
nand U6944 (N_6944,N_6721,N_6679);
or U6945 (N_6945,N_6787,N_6799);
nand U6946 (N_6946,N_6783,N_6733);
and U6947 (N_6947,N_6758,N_6620);
nand U6948 (N_6948,N_6649,N_6652);
nand U6949 (N_6949,N_6751,N_6654);
xnor U6950 (N_6950,N_6763,N_6768);
and U6951 (N_6951,N_6674,N_6683);
nand U6952 (N_6952,N_6679,N_6777);
or U6953 (N_6953,N_6731,N_6782);
and U6954 (N_6954,N_6619,N_6728);
or U6955 (N_6955,N_6612,N_6728);
nor U6956 (N_6956,N_6790,N_6686);
nor U6957 (N_6957,N_6694,N_6721);
and U6958 (N_6958,N_6779,N_6661);
nand U6959 (N_6959,N_6713,N_6609);
xor U6960 (N_6960,N_6629,N_6783);
and U6961 (N_6961,N_6762,N_6693);
nand U6962 (N_6962,N_6718,N_6703);
xor U6963 (N_6963,N_6720,N_6632);
xnor U6964 (N_6964,N_6654,N_6682);
nand U6965 (N_6965,N_6705,N_6701);
nor U6966 (N_6966,N_6767,N_6787);
nand U6967 (N_6967,N_6772,N_6687);
or U6968 (N_6968,N_6773,N_6677);
nand U6969 (N_6969,N_6799,N_6608);
nor U6970 (N_6970,N_6622,N_6685);
or U6971 (N_6971,N_6613,N_6783);
and U6972 (N_6972,N_6759,N_6655);
nor U6973 (N_6973,N_6605,N_6785);
or U6974 (N_6974,N_6741,N_6703);
and U6975 (N_6975,N_6636,N_6631);
nand U6976 (N_6976,N_6617,N_6611);
and U6977 (N_6977,N_6679,N_6768);
nor U6978 (N_6978,N_6663,N_6762);
nand U6979 (N_6979,N_6715,N_6683);
or U6980 (N_6980,N_6697,N_6640);
xor U6981 (N_6981,N_6756,N_6673);
and U6982 (N_6982,N_6761,N_6719);
xor U6983 (N_6983,N_6677,N_6792);
nand U6984 (N_6984,N_6661,N_6721);
nor U6985 (N_6985,N_6650,N_6727);
and U6986 (N_6986,N_6675,N_6718);
nand U6987 (N_6987,N_6657,N_6669);
or U6988 (N_6988,N_6797,N_6652);
nor U6989 (N_6989,N_6731,N_6701);
nand U6990 (N_6990,N_6646,N_6728);
xor U6991 (N_6991,N_6763,N_6790);
nand U6992 (N_6992,N_6671,N_6725);
nor U6993 (N_6993,N_6719,N_6769);
xor U6994 (N_6994,N_6734,N_6614);
nor U6995 (N_6995,N_6600,N_6792);
and U6996 (N_6996,N_6778,N_6614);
nand U6997 (N_6997,N_6681,N_6628);
and U6998 (N_6998,N_6740,N_6793);
xor U6999 (N_6999,N_6765,N_6669);
nand U7000 (N_7000,N_6883,N_6924);
and U7001 (N_7001,N_6820,N_6806);
nor U7002 (N_7002,N_6918,N_6972);
xnor U7003 (N_7003,N_6931,N_6919);
or U7004 (N_7004,N_6967,N_6963);
xnor U7005 (N_7005,N_6921,N_6953);
and U7006 (N_7006,N_6897,N_6940);
nor U7007 (N_7007,N_6923,N_6976);
nand U7008 (N_7008,N_6999,N_6836);
or U7009 (N_7009,N_6929,N_6930);
or U7010 (N_7010,N_6908,N_6888);
or U7011 (N_7011,N_6823,N_6941);
nor U7012 (N_7012,N_6948,N_6973);
nand U7013 (N_7013,N_6893,N_6814);
xor U7014 (N_7014,N_6861,N_6950);
nor U7015 (N_7015,N_6865,N_6828);
xor U7016 (N_7016,N_6896,N_6933);
nor U7017 (N_7017,N_6880,N_6899);
or U7018 (N_7018,N_6977,N_6834);
nand U7019 (N_7019,N_6832,N_6954);
nand U7020 (N_7020,N_6885,N_6879);
or U7021 (N_7021,N_6909,N_6847);
nand U7022 (N_7022,N_6824,N_6975);
nand U7023 (N_7023,N_6803,N_6958);
nand U7024 (N_7024,N_6943,N_6938);
xnor U7025 (N_7025,N_6868,N_6856);
nand U7026 (N_7026,N_6978,N_6959);
and U7027 (N_7027,N_6960,N_6934);
or U7028 (N_7028,N_6990,N_6985);
nor U7029 (N_7029,N_6882,N_6872);
and U7030 (N_7030,N_6851,N_6966);
nand U7031 (N_7031,N_6901,N_6840);
nor U7032 (N_7032,N_6887,N_6982);
nor U7033 (N_7033,N_6859,N_6889);
xnor U7034 (N_7034,N_6854,N_6841);
xor U7035 (N_7035,N_6855,N_6810);
nor U7036 (N_7036,N_6970,N_6905);
or U7037 (N_7037,N_6819,N_6964);
and U7038 (N_7038,N_6808,N_6804);
and U7039 (N_7039,N_6912,N_6936);
or U7040 (N_7040,N_6831,N_6875);
xor U7041 (N_7041,N_6987,N_6955);
xnor U7042 (N_7042,N_6946,N_6894);
xnor U7043 (N_7043,N_6986,N_6989);
xnor U7044 (N_7044,N_6971,N_6914);
xnor U7045 (N_7045,N_6805,N_6816);
or U7046 (N_7046,N_6947,N_6874);
and U7047 (N_7047,N_6926,N_6980);
and U7048 (N_7048,N_6838,N_6815);
and U7049 (N_7049,N_6956,N_6829);
nor U7050 (N_7050,N_6807,N_6939);
nor U7051 (N_7051,N_6965,N_6925);
nor U7052 (N_7052,N_6818,N_6949);
nor U7053 (N_7053,N_6913,N_6988);
xnor U7054 (N_7054,N_6864,N_6845);
or U7055 (N_7055,N_6866,N_6857);
nor U7056 (N_7056,N_6998,N_6904);
and U7057 (N_7057,N_6813,N_6871);
nand U7058 (N_7058,N_6898,N_6962);
and U7059 (N_7059,N_6830,N_6932);
or U7060 (N_7060,N_6983,N_6846);
and U7061 (N_7061,N_6825,N_6993);
nor U7062 (N_7062,N_6812,N_6863);
nand U7063 (N_7063,N_6811,N_6860);
nor U7064 (N_7064,N_6911,N_6944);
nand U7065 (N_7065,N_6850,N_6844);
and U7066 (N_7066,N_6867,N_6835);
nor U7067 (N_7067,N_6994,N_6800);
or U7068 (N_7068,N_6881,N_6809);
and U7069 (N_7069,N_6878,N_6848);
xor U7070 (N_7070,N_6886,N_6992);
or U7071 (N_7071,N_6906,N_6821);
nor U7072 (N_7072,N_6991,N_6951);
nand U7073 (N_7073,N_6843,N_6849);
or U7074 (N_7074,N_6979,N_6927);
and U7075 (N_7075,N_6969,N_6961);
nand U7076 (N_7076,N_6877,N_6942);
nor U7077 (N_7077,N_6890,N_6833);
nor U7078 (N_7078,N_6839,N_6826);
nor U7079 (N_7079,N_6917,N_6922);
or U7080 (N_7080,N_6900,N_6876);
or U7081 (N_7081,N_6891,N_6916);
nor U7082 (N_7082,N_6827,N_6995);
or U7083 (N_7083,N_6935,N_6974);
xor U7084 (N_7084,N_6915,N_6873);
or U7085 (N_7085,N_6920,N_6895);
nand U7086 (N_7086,N_6869,N_6822);
or U7087 (N_7087,N_6907,N_6801);
xnor U7088 (N_7088,N_6937,N_6903);
nand U7089 (N_7089,N_6981,N_6858);
and U7090 (N_7090,N_6945,N_6802);
or U7091 (N_7091,N_6870,N_6928);
and U7092 (N_7092,N_6910,N_6996);
nor U7093 (N_7093,N_6984,N_6997);
nand U7094 (N_7094,N_6817,N_6952);
nand U7095 (N_7095,N_6884,N_6957);
or U7096 (N_7096,N_6842,N_6853);
xor U7097 (N_7097,N_6862,N_6892);
nor U7098 (N_7098,N_6837,N_6852);
and U7099 (N_7099,N_6902,N_6968);
xor U7100 (N_7100,N_6943,N_6874);
or U7101 (N_7101,N_6945,N_6841);
nor U7102 (N_7102,N_6906,N_6869);
or U7103 (N_7103,N_6806,N_6988);
and U7104 (N_7104,N_6889,N_6981);
and U7105 (N_7105,N_6933,N_6909);
or U7106 (N_7106,N_6931,N_6817);
and U7107 (N_7107,N_6868,N_6992);
or U7108 (N_7108,N_6991,N_6899);
nor U7109 (N_7109,N_6817,N_6962);
or U7110 (N_7110,N_6914,N_6893);
nand U7111 (N_7111,N_6861,N_6896);
nand U7112 (N_7112,N_6891,N_6802);
xor U7113 (N_7113,N_6821,N_6844);
nand U7114 (N_7114,N_6939,N_6827);
xnor U7115 (N_7115,N_6857,N_6947);
xor U7116 (N_7116,N_6821,N_6953);
nand U7117 (N_7117,N_6814,N_6927);
and U7118 (N_7118,N_6914,N_6993);
or U7119 (N_7119,N_6888,N_6814);
nor U7120 (N_7120,N_6921,N_6943);
and U7121 (N_7121,N_6890,N_6829);
nand U7122 (N_7122,N_6996,N_6850);
nor U7123 (N_7123,N_6967,N_6861);
nand U7124 (N_7124,N_6964,N_6874);
xnor U7125 (N_7125,N_6903,N_6876);
xnor U7126 (N_7126,N_6837,N_6832);
and U7127 (N_7127,N_6865,N_6905);
xor U7128 (N_7128,N_6807,N_6954);
nor U7129 (N_7129,N_6951,N_6834);
nand U7130 (N_7130,N_6960,N_6998);
or U7131 (N_7131,N_6908,N_6901);
and U7132 (N_7132,N_6871,N_6875);
or U7133 (N_7133,N_6857,N_6888);
nor U7134 (N_7134,N_6868,N_6854);
or U7135 (N_7135,N_6887,N_6872);
nor U7136 (N_7136,N_6806,N_6812);
xnor U7137 (N_7137,N_6984,N_6994);
nand U7138 (N_7138,N_6907,N_6845);
nor U7139 (N_7139,N_6973,N_6874);
or U7140 (N_7140,N_6985,N_6873);
or U7141 (N_7141,N_6876,N_6913);
xnor U7142 (N_7142,N_6808,N_6811);
or U7143 (N_7143,N_6869,N_6889);
nand U7144 (N_7144,N_6961,N_6880);
nand U7145 (N_7145,N_6927,N_6948);
xor U7146 (N_7146,N_6915,N_6874);
or U7147 (N_7147,N_6935,N_6844);
or U7148 (N_7148,N_6804,N_6933);
and U7149 (N_7149,N_6877,N_6921);
xnor U7150 (N_7150,N_6875,N_6988);
nand U7151 (N_7151,N_6940,N_6914);
and U7152 (N_7152,N_6895,N_6826);
and U7153 (N_7153,N_6862,N_6969);
and U7154 (N_7154,N_6833,N_6987);
or U7155 (N_7155,N_6983,N_6916);
nor U7156 (N_7156,N_6981,N_6845);
or U7157 (N_7157,N_6990,N_6837);
or U7158 (N_7158,N_6974,N_6854);
nor U7159 (N_7159,N_6912,N_6862);
and U7160 (N_7160,N_6963,N_6809);
or U7161 (N_7161,N_6910,N_6921);
xnor U7162 (N_7162,N_6933,N_6818);
nor U7163 (N_7163,N_6950,N_6918);
or U7164 (N_7164,N_6871,N_6806);
nand U7165 (N_7165,N_6819,N_6857);
nand U7166 (N_7166,N_6810,N_6816);
nand U7167 (N_7167,N_6921,N_6995);
xor U7168 (N_7168,N_6811,N_6968);
or U7169 (N_7169,N_6856,N_6860);
or U7170 (N_7170,N_6921,N_6982);
nand U7171 (N_7171,N_6974,N_6942);
xnor U7172 (N_7172,N_6927,N_6959);
or U7173 (N_7173,N_6955,N_6885);
xor U7174 (N_7174,N_6948,N_6920);
xnor U7175 (N_7175,N_6896,N_6986);
or U7176 (N_7176,N_6800,N_6989);
or U7177 (N_7177,N_6967,N_6825);
or U7178 (N_7178,N_6952,N_6832);
and U7179 (N_7179,N_6871,N_6966);
and U7180 (N_7180,N_6966,N_6890);
xor U7181 (N_7181,N_6872,N_6987);
and U7182 (N_7182,N_6809,N_6836);
and U7183 (N_7183,N_6943,N_6995);
or U7184 (N_7184,N_6980,N_6976);
nand U7185 (N_7185,N_6930,N_6873);
nor U7186 (N_7186,N_6961,N_6895);
and U7187 (N_7187,N_6964,N_6924);
or U7188 (N_7188,N_6862,N_6926);
and U7189 (N_7189,N_6846,N_6903);
xor U7190 (N_7190,N_6996,N_6861);
and U7191 (N_7191,N_6924,N_6935);
xnor U7192 (N_7192,N_6915,N_6938);
or U7193 (N_7193,N_6955,N_6867);
or U7194 (N_7194,N_6933,N_6848);
nor U7195 (N_7195,N_6828,N_6968);
xnor U7196 (N_7196,N_6929,N_6920);
or U7197 (N_7197,N_6869,N_6939);
and U7198 (N_7198,N_6806,N_6961);
xor U7199 (N_7199,N_6816,N_6820);
or U7200 (N_7200,N_7119,N_7032);
nor U7201 (N_7201,N_7002,N_7038);
or U7202 (N_7202,N_7074,N_7188);
nor U7203 (N_7203,N_7116,N_7010);
or U7204 (N_7204,N_7181,N_7077);
xnor U7205 (N_7205,N_7072,N_7034);
xnor U7206 (N_7206,N_7155,N_7021);
and U7207 (N_7207,N_7138,N_7024);
and U7208 (N_7208,N_7030,N_7102);
and U7209 (N_7209,N_7054,N_7125);
xor U7210 (N_7210,N_7170,N_7092);
xnor U7211 (N_7211,N_7109,N_7189);
xnor U7212 (N_7212,N_7104,N_7123);
or U7213 (N_7213,N_7106,N_7046);
xnor U7214 (N_7214,N_7001,N_7137);
and U7215 (N_7215,N_7005,N_7084);
and U7216 (N_7216,N_7169,N_7168);
xor U7217 (N_7217,N_7112,N_7012);
xnor U7218 (N_7218,N_7060,N_7057);
nor U7219 (N_7219,N_7105,N_7098);
nor U7220 (N_7220,N_7113,N_7041);
xor U7221 (N_7221,N_7176,N_7075);
or U7222 (N_7222,N_7033,N_7108);
and U7223 (N_7223,N_7122,N_7114);
nor U7224 (N_7224,N_7083,N_7047);
and U7225 (N_7225,N_7146,N_7040);
xor U7226 (N_7226,N_7199,N_7088);
or U7227 (N_7227,N_7147,N_7071);
and U7228 (N_7228,N_7027,N_7049);
or U7229 (N_7229,N_7174,N_7016);
nor U7230 (N_7230,N_7158,N_7141);
nand U7231 (N_7231,N_7026,N_7070);
nor U7232 (N_7232,N_7140,N_7079);
nand U7233 (N_7233,N_7179,N_7187);
and U7234 (N_7234,N_7096,N_7035);
xnor U7235 (N_7235,N_7148,N_7023);
and U7236 (N_7236,N_7042,N_7044);
nor U7237 (N_7237,N_7110,N_7097);
nand U7238 (N_7238,N_7194,N_7180);
xor U7239 (N_7239,N_7173,N_7101);
xor U7240 (N_7240,N_7019,N_7153);
nor U7241 (N_7241,N_7061,N_7099);
xor U7242 (N_7242,N_7025,N_7080);
nor U7243 (N_7243,N_7091,N_7185);
or U7244 (N_7244,N_7161,N_7050);
and U7245 (N_7245,N_7053,N_7095);
or U7246 (N_7246,N_7039,N_7118);
or U7247 (N_7247,N_7190,N_7196);
or U7248 (N_7248,N_7064,N_7182);
and U7249 (N_7249,N_7059,N_7089);
and U7250 (N_7250,N_7036,N_7076);
nand U7251 (N_7251,N_7197,N_7150);
nand U7252 (N_7252,N_7166,N_7031);
nor U7253 (N_7253,N_7029,N_7164);
nor U7254 (N_7254,N_7062,N_7045);
or U7255 (N_7255,N_7154,N_7011);
nor U7256 (N_7256,N_7120,N_7127);
or U7257 (N_7257,N_7171,N_7142);
and U7258 (N_7258,N_7094,N_7100);
xor U7259 (N_7259,N_7165,N_7145);
nor U7260 (N_7260,N_7022,N_7160);
xor U7261 (N_7261,N_7191,N_7115);
nand U7262 (N_7262,N_7067,N_7193);
xor U7263 (N_7263,N_7186,N_7149);
xor U7264 (N_7264,N_7015,N_7066);
xnor U7265 (N_7265,N_7058,N_7135);
or U7266 (N_7266,N_7167,N_7082);
nor U7267 (N_7267,N_7052,N_7133);
nand U7268 (N_7268,N_7048,N_7007);
nand U7269 (N_7269,N_7131,N_7004);
or U7270 (N_7270,N_7132,N_7136);
nor U7271 (N_7271,N_7018,N_7008);
and U7272 (N_7272,N_7183,N_7159);
or U7273 (N_7273,N_7056,N_7198);
or U7274 (N_7274,N_7014,N_7134);
xnor U7275 (N_7275,N_7144,N_7121);
and U7276 (N_7276,N_7009,N_7003);
or U7277 (N_7277,N_7163,N_7090);
and U7278 (N_7278,N_7028,N_7107);
nor U7279 (N_7279,N_7051,N_7178);
or U7280 (N_7280,N_7085,N_7065);
xnor U7281 (N_7281,N_7006,N_7017);
and U7282 (N_7282,N_7124,N_7143);
xnor U7283 (N_7283,N_7020,N_7093);
nand U7284 (N_7284,N_7117,N_7037);
nand U7285 (N_7285,N_7055,N_7078);
xnor U7286 (N_7286,N_7043,N_7103);
and U7287 (N_7287,N_7175,N_7184);
nand U7288 (N_7288,N_7000,N_7152);
xor U7289 (N_7289,N_7069,N_7156);
nand U7290 (N_7290,N_7111,N_7068);
nor U7291 (N_7291,N_7087,N_7013);
or U7292 (N_7292,N_7162,N_7177);
and U7293 (N_7293,N_7129,N_7192);
xnor U7294 (N_7294,N_7126,N_7139);
xnor U7295 (N_7295,N_7130,N_7081);
or U7296 (N_7296,N_7128,N_7073);
or U7297 (N_7297,N_7157,N_7063);
nand U7298 (N_7298,N_7172,N_7086);
and U7299 (N_7299,N_7151,N_7195);
xnor U7300 (N_7300,N_7193,N_7074);
nor U7301 (N_7301,N_7074,N_7103);
nor U7302 (N_7302,N_7141,N_7182);
xor U7303 (N_7303,N_7087,N_7005);
or U7304 (N_7304,N_7169,N_7105);
nor U7305 (N_7305,N_7192,N_7138);
nand U7306 (N_7306,N_7125,N_7120);
xnor U7307 (N_7307,N_7067,N_7081);
or U7308 (N_7308,N_7057,N_7068);
or U7309 (N_7309,N_7112,N_7145);
or U7310 (N_7310,N_7015,N_7057);
nand U7311 (N_7311,N_7120,N_7058);
nand U7312 (N_7312,N_7010,N_7130);
or U7313 (N_7313,N_7044,N_7137);
and U7314 (N_7314,N_7036,N_7034);
nor U7315 (N_7315,N_7166,N_7115);
or U7316 (N_7316,N_7069,N_7035);
xor U7317 (N_7317,N_7023,N_7048);
nor U7318 (N_7318,N_7145,N_7189);
or U7319 (N_7319,N_7078,N_7113);
nand U7320 (N_7320,N_7080,N_7167);
and U7321 (N_7321,N_7064,N_7052);
and U7322 (N_7322,N_7081,N_7141);
nor U7323 (N_7323,N_7176,N_7185);
xor U7324 (N_7324,N_7076,N_7121);
nand U7325 (N_7325,N_7066,N_7080);
and U7326 (N_7326,N_7196,N_7156);
and U7327 (N_7327,N_7031,N_7065);
and U7328 (N_7328,N_7168,N_7083);
nand U7329 (N_7329,N_7034,N_7021);
or U7330 (N_7330,N_7040,N_7019);
and U7331 (N_7331,N_7117,N_7064);
and U7332 (N_7332,N_7005,N_7198);
nand U7333 (N_7333,N_7090,N_7096);
nor U7334 (N_7334,N_7176,N_7181);
nand U7335 (N_7335,N_7098,N_7022);
and U7336 (N_7336,N_7115,N_7101);
nand U7337 (N_7337,N_7150,N_7038);
and U7338 (N_7338,N_7147,N_7142);
nand U7339 (N_7339,N_7021,N_7129);
or U7340 (N_7340,N_7076,N_7067);
and U7341 (N_7341,N_7176,N_7030);
xor U7342 (N_7342,N_7122,N_7048);
xnor U7343 (N_7343,N_7083,N_7196);
and U7344 (N_7344,N_7126,N_7086);
and U7345 (N_7345,N_7166,N_7000);
xor U7346 (N_7346,N_7175,N_7071);
xor U7347 (N_7347,N_7105,N_7020);
or U7348 (N_7348,N_7068,N_7129);
and U7349 (N_7349,N_7040,N_7005);
xor U7350 (N_7350,N_7007,N_7173);
nor U7351 (N_7351,N_7130,N_7072);
or U7352 (N_7352,N_7191,N_7006);
xnor U7353 (N_7353,N_7078,N_7012);
nand U7354 (N_7354,N_7088,N_7106);
or U7355 (N_7355,N_7175,N_7157);
nand U7356 (N_7356,N_7085,N_7075);
and U7357 (N_7357,N_7050,N_7020);
xor U7358 (N_7358,N_7111,N_7088);
or U7359 (N_7359,N_7161,N_7020);
xnor U7360 (N_7360,N_7169,N_7137);
and U7361 (N_7361,N_7181,N_7125);
nand U7362 (N_7362,N_7027,N_7022);
xor U7363 (N_7363,N_7093,N_7034);
nand U7364 (N_7364,N_7100,N_7022);
and U7365 (N_7365,N_7176,N_7010);
nor U7366 (N_7366,N_7169,N_7018);
nand U7367 (N_7367,N_7086,N_7154);
or U7368 (N_7368,N_7014,N_7132);
nor U7369 (N_7369,N_7128,N_7173);
nand U7370 (N_7370,N_7039,N_7137);
nor U7371 (N_7371,N_7084,N_7000);
nor U7372 (N_7372,N_7159,N_7077);
or U7373 (N_7373,N_7026,N_7147);
and U7374 (N_7374,N_7160,N_7027);
nand U7375 (N_7375,N_7062,N_7197);
xnor U7376 (N_7376,N_7071,N_7004);
and U7377 (N_7377,N_7085,N_7000);
xnor U7378 (N_7378,N_7170,N_7172);
xnor U7379 (N_7379,N_7184,N_7081);
nand U7380 (N_7380,N_7044,N_7007);
and U7381 (N_7381,N_7050,N_7088);
and U7382 (N_7382,N_7063,N_7029);
nand U7383 (N_7383,N_7014,N_7016);
xor U7384 (N_7384,N_7046,N_7077);
nor U7385 (N_7385,N_7022,N_7162);
nor U7386 (N_7386,N_7147,N_7062);
xor U7387 (N_7387,N_7016,N_7062);
or U7388 (N_7388,N_7104,N_7081);
and U7389 (N_7389,N_7004,N_7022);
or U7390 (N_7390,N_7001,N_7125);
and U7391 (N_7391,N_7117,N_7085);
nand U7392 (N_7392,N_7123,N_7133);
or U7393 (N_7393,N_7064,N_7151);
and U7394 (N_7394,N_7190,N_7047);
and U7395 (N_7395,N_7049,N_7193);
or U7396 (N_7396,N_7123,N_7030);
and U7397 (N_7397,N_7187,N_7091);
nor U7398 (N_7398,N_7150,N_7177);
and U7399 (N_7399,N_7084,N_7125);
nand U7400 (N_7400,N_7224,N_7389);
or U7401 (N_7401,N_7331,N_7368);
or U7402 (N_7402,N_7307,N_7325);
or U7403 (N_7403,N_7254,N_7223);
or U7404 (N_7404,N_7210,N_7298);
nand U7405 (N_7405,N_7329,N_7317);
nand U7406 (N_7406,N_7211,N_7270);
and U7407 (N_7407,N_7232,N_7381);
and U7408 (N_7408,N_7302,N_7393);
and U7409 (N_7409,N_7280,N_7205);
nor U7410 (N_7410,N_7345,N_7225);
nor U7411 (N_7411,N_7263,N_7286);
nor U7412 (N_7412,N_7228,N_7367);
nand U7413 (N_7413,N_7332,N_7249);
xor U7414 (N_7414,N_7314,N_7274);
or U7415 (N_7415,N_7388,N_7230);
nor U7416 (N_7416,N_7337,N_7273);
nor U7417 (N_7417,N_7374,N_7242);
nor U7418 (N_7418,N_7271,N_7354);
xor U7419 (N_7419,N_7304,N_7236);
xnor U7420 (N_7420,N_7220,N_7204);
nor U7421 (N_7421,N_7378,N_7330);
nor U7422 (N_7422,N_7216,N_7221);
nand U7423 (N_7423,N_7247,N_7371);
nor U7424 (N_7424,N_7260,N_7217);
nor U7425 (N_7425,N_7311,N_7310);
or U7426 (N_7426,N_7227,N_7305);
nand U7427 (N_7427,N_7200,N_7276);
or U7428 (N_7428,N_7398,N_7320);
xnor U7429 (N_7429,N_7278,N_7243);
and U7430 (N_7430,N_7350,N_7246);
xnor U7431 (N_7431,N_7362,N_7285);
xnor U7432 (N_7432,N_7341,N_7312);
nor U7433 (N_7433,N_7358,N_7370);
and U7434 (N_7434,N_7335,N_7293);
nand U7435 (N_7435,N_7372,N_7322);
xor U7436 (N_7436,N_7279,N_7303);
and U7437 (N_7437,N_7252,N_7256);
xor U7438 (N_7438,N_7299,N_7399);
xor U7439 (N_7439,N_7283,N_7219);
xor U7440 (N_7440,N_7364,N_7376);
and U7441 (N_7441,N_7385,N_7347);
or U7442 (N_7442,N_7288,N_7353);
or U7443 (N_7443,N_7379,N_7231);
or U7444 (N_7444,N_7318,N_7396);
xor U7445 (N_7445,N_7208,N_7218);
or U7446 (N_7446,N_7319,N_7295);
nor U7447 (N_7447,N_7309,N_7222);
or U7448 (N_7448,N_7262,N_7386);
and U7449 (N_7449,N_7214,N_7206);
or U7450 (N_7450,N_7382,N_7296);
xor U7451 (N_7451,N_7383,N_7248);
and U7452 (N_7452,N_7292,N_7290);
xor U7453 (N_7453,N_7234,N_7342);
nand U7454 (N_7454,N_7306,N_7377);
and U7455 (N_7455,N_7265,N_7259);
nor U7456 (N_7456,N_7201,N_7255);
nor U7457 (N_7457,N_7373,N_7245);
or U7458 (N_7458,N_7360,N_7326);
nor U7459 (N_7459,N_7300,N_7355);
and U7460 (N_7460,N_7375,N_7343);
nor U7461 (N_7461,N_7387,N_7384);
nand U7462 (N_7462,N_7363,N_7229);
xor U7463 (N_7463,N_7284,N_7261);
xnor U7464 (N_7464,N_7277,N_7338);
nor U7465 (N_7465,N_7324,N_7287);
nor U7466 (N_7466,N_7395,N_7357);
nand U7467 (N_7467,N_7275,N_7351);
xnor U7468 (N_7468,N_7334,N_7281);
nor U7469 (N_7469,N_7207,N_7313);
xor U7470 (N_7470,N_7202,N_7380);
nand U7471 (N_7471,N_7289,N_7253);
nor U7472 (N_7472,N_7282,N_7203);
and U7473 (N_7473,N_7267,N_7369);
nand U7474 (N_7474,N_7348,N_7333);
or U7475 (N_7475,N_7241,N_7215);
xor U7476 (N_7476,N_7336,N_7321);
nor U7477 (N_7477,N_7327,N_7258);
xnor U7478 (N_7478,N_7239,N_7365);
xnor U7479 (N_7479,N_7339,N_7268);
xnor U7480 (N_7480,N_7257,N_7328);
nor U7481 (N_7481,N_7244,N_7294);
nand U7482 (N_7482,N_7344,N_7359);
xnor U7483 (N_7483,N_7301,N_7392);
and U7484 (N_7484,N_7361,N_7397);
and U7485 (N_7485,N_7356,N_7352);
and U7486 (N_7486,N_7390,N_7269);
and U7487 (N_7487,N_7366,N_7272);
nor U7488 (N_7488,N_7235,N_7212);
or U7489 (N_7489,N_7233,N_7323);
nor U7490 (N_7490,N_7349,N_7240);
xor U7491 (N_7491,N_7291,N_7308);
and U7492 (N_7492,N_7266,N_7340);
xnor U7493 (N_7493,N_7226,N_7209);
xnor U7494 (N_7494,N_7316,N_7251);
nand U7495 (N_7495,N_7264,N_7315);
or U7496 (N_7496,N_7297,N_7394);
xnor U7497 (N_7497,N_7250,N_7391);
or U7498 (N_7498,N_7346,N_7237);
and U7499 (N_7499,N_7238,N_7213);
and U7500 (N_7500,N_7388,N_7218);
or U7501 (N_7501,N_7227,N_7302);
or U7502 (N_7502,N_7275,N_7313);
nor U7503 (N_7503,N_7363,N_7285);
xnor U7504 (N_7504,N_7298,N_7306);
nor U7505 (N_7505,N_7366,N_7256);
or U7506 (N_7506,N_7335,N_7316);
nor U7507 (N_7507,N_7321,N_7309);
xnor U7508 (N_7508,N_7234,N_7291);
nand U7509 (N_7509,N_7384,N_7222);
xnor U7510 (N_7510,N_7387,N_7314);
or U7511 (N_7511,N_7213,N_7203);
nor U7512 (N_7512,N_7344,N_7293);
or U7513 (N_7513,N_7207,N_7378);
or U7514 (N_7514,N_7222,N_7365);
nor U7515 (N_7515,N_7215,N_7382);
nor U7516 (N_7516,N_7381,N_7305);
or U7517 (N_7517,N_7273,N_7244);
and U7518 (N_7518,N_7397,N_7313);
and U7519 (N_7519,N_7206,N_7337);
and U7520 (N_7520,N_7270,N_7379);
or U7521 (N_7521,N_7233,N_7274);
nor U7522 (N_7522,N_7319,N_7282);
xor U7523 (N_7523,N_7309,N_7377);
or U7524 (N_7524,N_7396,N_7271);
or U7525 (N_7525,N_7266,N_7310);
xnor U7526 (N_7526,N_7310,N_7378);
nand U7527 (N_7527,N_7395,N_7293);
xnor U7528 (N_7528,N_7326,N_7389);
nand U7529 (N_7529,N_7261,N_7227);
or U7530 (N_7530,N_7378,N_7347);
and U7531 (N_7531,N_7348,N_7336);
or U7532 (N_7532,N_7320,N_7227);
xor U7533 (N_7533,N_7265,N_7393);
and U7534 (N_7534,N_7362,N_7289);
xor U7535 (N_7535,N_7398,N_7305);
and U7536 (N_7536,N_7399,N_7348);
xor U7537 (N_7537,N_7336,N_7271);
nor U7538 (N_7538,N_7231,N_7251);
xnor U7539 (N_7539,N_7280,N_7287);
xor U7540 (N_7540,N_7255,N_7340);
and U7541 (N_7541,N_7231,N_7355);
nand U7542 (N_7542,N_7242,N_7366);
and U7543 (N_7543,N_7311,N_7262);
xnor U7544 (N_7544,N_7356,N_7223);
nor U7545 (N_7545,N_7346,N_7376);
or U7546 (N_7546,N_7295,N_7274);
nor U7547 (N_7547,N_7257,N_7252);
and U7548 (N_7548,N_7398,N_7342);
nand U7549 (N_7549,N_7361,N_7356);
nor U7550 (N_7550,N_7209,N_7332);
nand U7551 (N_7551,N_7368,N_7332);
and U7552 (N_7552,N_7390,N_7386);
xor U7553 (N_7553,N_7266,N_7316);
or U7554 (N_7554,N_7366,N_7302);
xnor U7555 (N_7555,N_7246,N_7371);
nand U7556 (N_7556,N_7378,N_7300);
nand U7557 (N_7557,N_7293,N_7386);
xnor U7558 (N_7558,N_7205,N_7394);
xnor U7559 (N_7559,N_7326,N_7256);
nor U7560 (N_7560,N_7208,N_7206);
xnor U7561 (N_7561,N_7201,N_7368);
and U7562 (N_7562,N_7310,N_7206);
nand U7563 (N_7563,N_7378,N_7249);
xor U7564 (N_7564,N_7207,N_7271);
or U7565 (N_7565,N_7391,N_7226);
nand U7566 (N_7566,N_7279,N_7276);
nor U7567 (N_7567,N_7220,N_7380);
and U7568 (N_7568,N_7297,N_7300);
nand U7569 (N_7569,N_7263,N_7207);
nor U7570 (N_7570,N_7392,N_7296);
xnor U7571 (N_7571,N_7270,N_7394);
or U7572 (N_7572,N_7399,N_7330);
xor U7573 (N_7573,N_7325,N_7330);
nor U7574 (N_7574,N_7362,N_7385);
or U7575 (N_7575,N_7397,N_7201);
and U7576 (N_7576,N_7357,N_7386);
nor U7577 (N_7577,N_7290,N_7281);
nand U7578 (N_7578,N_7326,N_7343);
and U7579 (N_7579,N_7316,N_7225);
nor U7580 (N_7580,N_7228,N_7314);
and U7581 (N_7581,N_7312,N_7394);
xnor U7582 (N_7582,N_7300,N_7348);
nand U7583 (N_7583,N_7369,N_7233);
xnor U7584 (N_7584,N_7399,N_7395);
nor U7585 (N_7585,N_7241,N_7335);
nand U7586 (N_7586,N_7210,N_7281);
xnor U7587 (N_7587,N_7326,N_7385);
xnor U7588 (N_7588,N_7329,N_7399);
and U7589 (N_7589,N_7300,N_7206);
and U7590 (N_7590,N_7204,N_7297);
xor U7591 (N_7591,N_7299,N_7258);
xnor U7592 (N_7592,N_7366,N_7320);
xnor U7593 (N_7593,N_7211,N_7308);
nor U7594 (N_7594,N_7385,N_7243);
or U7595 (N_7595,N_7393,N_7267);
nor U7596 (N_7596,N_7360,N_7237);
and U7597 (N_7597,N_7391,N_7349);
and U7598 (N_7598,N_7235,N_7381);
and U7599 (N_7599,N_7395,N_7312);
nor U7600 (N_7600,N_7456,N_7536);
and U7601 (N_7601,N_7596,N_7426);
or U7602 (N_7602,N_7447,N_7494);
nor U7603 (N_7603,N_7419,N_7488);
nor U7604 (N_7604,N_7427,N_7436);
xor U7605 (N_7605,N_7515,N_7554);
and U7606 (N_7606,N_7444,N_7583);
and U7607 (N_7607,N_7483,N_7527);
xnor U7608 (N_7608,N_7428,N_7418);
xnor U7609 (N_7609,N_7566,N_7533);
nor U7610 (N_7610,N_7517,N_7534);
or U7611 (N_7611,N_7597,N_7469);
or U7612 (N_7612,N_7518,N_7595);
nand U7613 (N_7613,N_7409,N_7516);
and U7614 (N_7614,N_7522,N_7430);
and U7615 (N_7615,N_7450,N_7460);
nor U7616 (N_7616,N_7570,N_7417);
nor U7617 (N_7617,N_7452,N_7551);
or U7618 (N_7618,N_7415,N_7402);
xnor U7619 (N_7619,N_7586,N_7470);
xnor U7620 (N_7620,N_7558,N_7520);
nor U7621 (N_7621,N_7414,N_7569);
and U7622 (N_7622,N_7521,N_7571);
or U7623 (N_7623,N_7529,N_7504);
nor U7624 (N_7624,N_7584,N_7467);
and U7625 (N_7625,N_7526,N_7464);
or U7626 (N_7626,N_7547,N_7400);
nand U7627 (N_7627,N_7519,N_7545);
and U7628 (N_7628,N_7446,N_7514);
xnor U7629 (N_7629,N_7429,N_7531);
nand U7630 (N_7630,N_7567,N_7535);
or U7631 (N_7631,N_7579,N_7591);
nor U7632 (N_7632,N_7482,N_7538);
xnor U7633 (N_7633,N_7537,N_7562);
and U7634 (N_7634,N_7403,N_7421);
nor U7635 (N_7635,N_7552,N_7497);
nor U7636 (N_7636,N_7445,N_7512);
xnor U7637 (N_7637,N_7471,N_7561);
nor U7638 (N_7638,N_7466,N_7424);
and U7639 (N_7639,N_7524,N_7443);
nor U7640 (N_7640,N_7434,N_7523);
and U7641 (N_7641,N_7498,N_7573);
or U7642 (N_7642,N_7543,N_7412);
nor U7643 (N_7643,N_7506,N_7416);
nand U7644 (N_7644,N_7599,N_7493);
or U7645 (N_7645,N_7431,N_7578);
nand U7646 (N_7646,N_7441,N_7559);
xnor U7647 (N_7647,N_7574,N_7541);
or U7648 (N_7648,N_7475,N_7525);
nor U7649 (N_7649,N_7411,N_7565);
xor U7650 (N_7650,N_7576,N_7598);
nand U7651 (N_7651,N_7496,N_7438);
or U7652 (N_7652,N_7433,N_7503);
xor U7653 (N_7653,N_7481,N_7413);
or U7654 (N_7654,N_7492,N_7407);
or U7655 (N_7655,N_7468,N_7457);
nand U7656 (N_7656,N_7401,N_7485);
nand U7657 (N_7657,N_7592,N_7508);
or U7658 (N_7658,N_7474,N_7472);
and U7659 (N_7659,N_7404,N_7440);
nand U7660 (N_7660,N_7449,N_7575);
nor U7661 (N_7661,N_7486,N_7422);
and U7662 (N_7662,N_7563,N_7513);
nor U7663 (N_7663,N_7442,N_7410);
nand U7664 (N_7664,N_7490,N_7408);
xor U7665 (N_7665,N_7476,N_7487);
or U7666 (N_7666,N_7581,N_7458);
and U7667 (N_7667,N_7502,N_7590);
or U7668 (N_7668,N_7580,N_7477);
xor U7669 (N_7669,N_7555,N_7405);
and U7670 (N_7670,N_7439,N_7448);
or U7671 (N_7671,N_7509,N_7451);
and U7672 (N_7672,N_7585,N_7546);
xor U7673 (N_7673,N_7489,N_7540);
and U7674 (N_7674,N_7507,N_7530);
nor U7675 (N_7675,N_7589,N_7454);
xor U7676 (N_7676,N_7553,N_7594);
xor U7677 (N_7677,N_7453,N_7588);
nand U7678 (N_7678,N_7501,N_7587);
xnor U7679 (N_7679,N_7511,N_7532);
xnor U7680 (N_7680,N_7455,N_7564);
nor U7681 (N_7681,N_7542,N_7425);
or U7682 (N_7682,N_7495,N_7510);
xnor U7683 (N_7683,N_7593,N_7465);
and U7684 (N_7684,N_7550,N_7459);
xnor U7685 (N_7685,N_7572,N_7461);
or U7686 (N_7686,N_7528,N_7491);
nor U7687 (N_7687,N_7505,N_7479);
or U7688 (N_7688,N_7557,N_7544);
and U7689 (N_7689,N_7473,N_7480);
and U7690 (N_7690,N_7539,N_7582);
or U7691 (N_7691,N_7560,N_7462);
nand U7692 (N_7692,N_7548,N_7499);
nand U7693 (N_7693,N_7500,N_7423);
or U7694 (N_7694,N_7577,N_7478);
xnor U7695 (N_7695,N_7549,N_7406);
xor U7696 (N_7696,N_7568,N_7463);
and U7697 (N_7697,N_7420,N_7435);
nor U7698 (N_7698,N_7484,N_7437);
nand U7699 (N_7699,N_7432,N_7556);
and U7700 (N_7700,N_7459,N_7569);
and U7701 (N_7701,N_7560,N_7544);
nand U7702 (N_7702,N_7591,N_7562);
and U7703 (N_7703,N_7509,N_7582);
xnor U7704 (N_7704,N_7501,N_7583);
or U7705 (N_7705,N_7499,N_7478);
or U7706 (N_7706,N_7441,N_7430);
nand U7707 (N_7707,N_7449,N_7542);
and U7708 (N_7708,N_7563,N_7493);
nand U7709 (N_7709,N_7594,N_7555);
nand U7710 (N_7710,N_7440,N_7484);
nand U7711 (N_7711,N_7494,N_7449);
and U7712 (N_7712,N_7433,N_7513);
or U7713 (N_7713,N_7456,N_7564);
xor U7714 (N_7714,N_7590,N_7413);
nand U7715 (N_7715,N_7481,N_7404);
nor U7716 (N_7716,N_7598,N_7469);
nand U7717 (N_7717,N_7435,N_7503);
and U7718 (N_7718,N_7434,N_7527);
xnor U7719 (N_7719,N_7579,N_7447);
nand U7720 (N_7720,N_7498,N_7441);
nand U7721 (N_7721,N_7563,N_7578);
nand U7722 (N_7722,N_7598,N_7487);
nand U7723 (N_7723,N_7432,N_7511);
and U7724 (N_7724,N_7491,N_7408);
or U7725 (N_7725,N_7414,N_7422);
nand U7726 (N_7726,N_7520,N_7459);
or U7727 (N_7727,N_7501,N_7487);
nand U7728 (N_7728,N_7488,N_7530);
nand U7729 (N_7729,N_7566,N_7551);
nor U7730 (N_7730,N_7405,N_7572);
nor U7731 (N_7731,N_7580,N_7517);
xnor U7732 (N_7732,N_7557,N_7504);
and U7733 (N_7733,N_7439,N_7517);
and U7734 (N_7734,N_7483,N_7512);
nand U7735 (N_7735,N_7488,N_7583);
and U7736 (N_7736,N_7589,N_7464);
nor U7737 (N_7737,N_7423,N_7482);
nor U7738 (N_7738,N_7566,N_7498);
nand U7739 (N_7739,N_7537,N_7557);
and U7740 (N_7740,N_7467,N_7423);
nor U7741 (N_7741,N_7508,N_7516);
nand U7742 (N_7742,N_7570,N_7510);
nor U7743 (N_7743,N_7527,N_7459);
xnor U7744 (N_7744,N_7458,N_7426);
xnor U7745 (N_7745,N_7428,N_7543);
nand U7746 (N_7746,N_7597,N_7519);
nand U7747 (N_7747,N_7522,N_7419);
xor U7748 (N_7748,N_7405,N_7416);
xnor U7749 (N_7749,N_7562,N_7430);
xor U7750 (N_7750,N_7460,N_7427);
nor U7751 (N_7751,N_7580,N_7570);
nand U7752 (N_7752,N_7506,N_7432);
or U7753 (N_7753,N_7519,N_7475);
or U7754 (N_7754,N_7539,N_7414);
nor U7755 (N_7755,N_7537,N_7561);
xnor U7756 (N_7756,N_7594,N_7515);
nor U7757 (N_7757,N_7564,N_7521);
and U7758 (N_7758,N_7405,N_7484);
or U7759 (N_7759,N_7509,N_7470);
nand U7760 (N_7760,N_7461,N_7569);
or U7761 (N_7761,N_7446,N_7584);
xnor U7762 (N_7762,N_7543,N_7432);
xor U7763 (N_7763,N_7555,N_7523);
and U7764 (N_7764,N_7415,N_7454);
nand U7765 (N_7765,N_7408,N_7435);
xor U7766 (N_7766,N_7436,N_7526);
xor U7767 (N_7767,N_7422,N_7473);
xor U7768 (N_7768,N_7434,N_7548);
and U7769 (N_7769,N_7433,N_7521);
nor U7770 (N_7770,N_7419,N_7446);
xor U7771 (N_7771,N_7469,N_7453);
nand U7772 (N_7772,N_7573,N_7516);
nand U7773 (N_7773,N_7557,N_7455);
xor U7774 (N_7774,N_7527,N_7559);
or U7775 (N_7775,N_7497,N_7506);
and U7776 (N_7776,N_7402,N_7442);
nor U7777 (N_7777,N_7525,N_7431);
nand U7778 (N_7778,N_7587,N_7465);
xor U7779 (N_7779,N_7583,N_7404);
xor U7780 (N_7780,N_7496,N_7490);
nand U7781 (N_7781,N_7557,N_7506);
xnor U7782 (N_7782,N_7572,N_7599);
xor U7783 (N_7783,N_7502,N_7505);
nand U7784 (N_7784,N_7549,N_7519);
or U7785 (N_7785,N_7449,N_7530);
or U7786 (N_7786,N_7446,N_7437);
xor U7787 (N_7787,N_7527,N_7489);
or U7788 (N_7788,N_7487,N_7508);
or U7789 (N_7789,N_7433,N_7529);
nor U7790 (N_7790,N_7498,N_7521);
xor U7791 (N_7791,N_7503,N_7572);
nand U7792 (N_7792,N_7424,N_7552);
and U7793 (N_7793,N_7427,N_7520);
or U7794 (N_7794,N_7435,N_7443);
and U7795 (N_7795,N_7462,N_7555);
nand U7796 (N_7796,N_7408,N_7495);
or U7797 (N_7797,N_7438,N_7480);
and U7798 (N_7798,N_7439,N_7554);
or U7799 (N_7799,N_7417,N_7473);
or U7800 (N_7800,N_7690,N_7643);
nor U7801 (N_7801,N_7608,N_7761);
nand U7802 (N_7802,N_7655,N_7730);
xor U7803 (N_7803,N_7654,N_7718);
nor U7804 (N_7804,N_7788,N_7689);
nor U7805 (N_7805,N_7602,N_7701);
nand U7806 (N_7806,N_7716,N_7710);
nor U7807 (N_7807,N_7630,N_7627);
nand U7808 (N_7808,N_7721,N_7691);
xnor U7809 (N_7809,N_7603,N_7644);
nand U7810 (N_7810,N_7767,N_7723);
xnor U7811 (N_7811,N_7660,N_7645);
and U7812 (N_7812,N_7686,N_7757);
nand U7813 (N_7813,N_7684,N_7613);
or U7814 (N_7814,N_7799,N_7623);
xor U7815 (N_7815,N_7778,N_7614);
nand U7816 (N_7816,N_7620,N_7739);
and U7817 (N_7817,N_7752,N_7753);
nor U7818 (N_7818,N_7781,N_7766);
xor U7819 (N_7819,N_7783,N_7798);
nand U7820 (N_7820,N_7657,N_7708);
nor U7821 (N_7821,N_7683,N_7679);
nor U7822 (N_7822,N_7735,N_7707);
nand U7823 (N_7823,N_7664,N_7764);
nand U7824 (N_7824,N_7626,N_7652);
or U7825 (N_7825,N_7647,N_7715);
nor U7826 (N_7826,N_7675,N_7725);
nand U7827 (N_7827,N_7604,N_7663);
nor U7828 (N_7828,N_7750,N_7661);
or U7829 (N_7829,N_7672,N_7616);
or U7830 (N_7830,N_7702,N_7659);
nor U7831 (N_7831,N_7688,N_7697);
nand U7832 (N_7832,N_7617,N_7698);
nand U7833 (N_7833,N_7703,N_7605);
nor U7834 (N_7834,N_7745,N_7769);
nor U7835 (N_7835,N_7796,N_7726);
or U7836 (N_7836,N_7736,N_7685);
or U7837 (N_7837,N_7775,N_7768);
or U7838 (N_7838,N_7622,N_7633);
xnor U7839 (N_7839,N_7743,N_7607);
nand U7840 (N_7840,N_7674,N_7747);
or U7841 (N_7841,N_7741,N_7787);
nor U7842 (N_7842,N_7774,N_7760);
and U7843 (N_7843,N_7722,N_7662);
and U7844 (N_7844,N_7668,N_7621);
xor U7845 (N_7845,N_7610,N_7635);
or U7846 (N_7846,N_7665,N_7628);
and U7847 (N_7847,N_7667,N_7648);
xor U7848 (N_7848,N_7714,N_7680);
nor U7849 (N_7849,N_7777,N_7794);
or U7850 (N_7850,N_7719,N_7651);
or U7851 (N_7851,N_7656,N_7780);
or U7852 (N_7852,N_7713,N_7770);
and U7853 (N_7853,N_7776,N_7748);
nand U7854 (N_7854,N_7749,N_7638);
nand U7855 (N_7855,N_7612,N_7600);
and U7856 (N_7856,N_7677,N_7789);
and U7857 (N_7857,N_7609,N_7695);
nand U7858 (N_7858,N_7694,N_7792);
or U7859 (N_7859,N_7731,N_7636);
xor U7860 (N_7860,N_7673,N_7717);
nand U7861 (N_7861,N_7797,N_7693);
or U7862 (N_7862,N_7692,N_7737);
or U7863 (N_7863,N_7759,N_7709);
or U7864 (N_7864,N_7642,N_7790);
xor U7865 (N_7865,N_7649,N_7639);
or U7866 (N_7866,N_7740,N_7763);
nand U7867 (N_7867,N_7640,N_7772);
xor U7868 (N_7868,N_7729,N_7720);
xnor U7869 (N_7869,N_7733,N_7724);
nand U7870 (N_7870,N_7625,N_7754);
xnor U7871 (N_7871,N_7751,N_7629);
or U7872 (N_7872,N_7670,N_7732);
xor U7873 (N_7873,N_7618,N_7742);
nor U7874 (N_7874,N_7744,N_7678);
nor U7875 (N_7875,N_7773,N_7706);
or U7876 (N_7876,N_7637,N_7681);
nand U7877 (N_7877,N_7671,N_7632);
and U7878 (N_7878,N_7765,N_7728);
and U7879 (N_7879,N_7624,N_7791);
nor U7880 (N_7880,N_7606,N_7687);
nor U7881 (N_7881,N_7711,N_7666);
or U7882 (N_7882,N_7696,N_7615);
or U7883 (N_7883,N_7619,N_7793);
and U7884 (N_7884,N_7611,N_7653);
nand U7885 (N_7885,N_7756,N_7727);
or U7886 (N_7886,N_7704,N_7634);
or U7887 (N_7887,N_7631,N_7669);
and U7888 (N_7888,N_7779,N_7786);
xnor U7889 (N_7889,N_7782,N_7705);
or U7890 (N_7890,N_7601,N_7762);
or U7891 (N_7891,N_7699,N_7682);
nand U7892 (N_7892,N_7785,N_7784);
and U7893 (N_7893,N_7755,N_7771);
nand U7894 (N_7894,N_7700,N_7646);
nand U7895 (N_7895,N_7734,N_7676);
and U7896 (N_7896,N_7746,N_7658);
nor U7897 (N_7897,N_7795,N_7738);
or U7898 (N_7898,N_7641,N_7712);
xnor U7899 (N_7899,N_7650,N_7758);
and U7900 (N_7900,N_7681,N_7685);
and U7901 (N_7901,N_7701,N_7783);
or U7902 (N_7902,N_7788,N_7774);
xor U7903 (N_7903,N_7713,N_7693);
nand U7904 (N_7904,N_7652,N_7704);
and U7905 (N_7905,N_7775,N_7650);
nor U7906 (N_7906,N_7641,N_7701);
nor U7907 (N_7907,N_7716,N_7780);
xor U7908 (N_7908,N_7668,N_7797);
or U7909 (N_7909,N_7758,N_7633);
nand U7910 (N_7910,N_7786,N_7665);
and U7911 (N_7911,N_7678,N_7653);
nand U7912 (N_7912,N_7671,N_7773);
xnor U7913 (N_7913,N_7695,N_7697);
nand U7914 (N_7914,N_7626,N_7641);
nand U7915 (N_7915,N_7661,N_7668);
nand U7916 (N_7916,N_7666,N_7730);
xor U7917 (N_7917,N_7775,N_7655);
nand U7918 (N_7918,N_7642,N_7707);
nor U7919 (N_7919,N_7698,N_7795);
and U7920 (N_7920,N_7788,N_7703);
nand U7921 (N_7921,N_7743,N_7794);
xnor U7922 (N_7922,N_7783,N_7623);
nand U7923 (N_7923,N_7652,N_7766);
and U7924 (N_7924,N_7670,N_7656);
or U7925 (N_7925,N_7798,N_7705);
nand U7926 (N_7926,N_7708,N_7633);
nor U7927 (N_7927,N_7634,N_7645);
xor U7928 (N_7928,N_7751,N_7768);
xor U7929 (N_7929,N_7703,N_7661);
xnor U7930 (N_7930,N_7630,N_7624);
xor U7931 (N_7931,N_7776,N_7628);
xor U7932 (N_7932,N_7651,N_7780);
nand U7933 (N_7933,N_7616,N_7775);
nand U7934 (N_7934,N_7785,N_7636);
nor U7935 (N_7935,N_7748,N_7754);
xor U7936 (N_7936,N_7699,N_7654);
and U7937 (N_7937,N_7641,N_7713);
and U7938 (N_7938,N_7606,N_7629);
and U7939 (N_7939,N_7603,N_7732);
xor U7940 (N_7940,N_7664,N_7659);
or U7941 (N_7941,N_7655,N_7748);
and U7942 (N_7942,N_7734,N_7793);
nor U7943 (N_7943,N_7781,N_7605);
and U7944 (N_7944,N_7691,N_7669);
or U7945 (N_7945,N_7728,N_7704);
xnor U7946 (N_7946,N_7760,N_7726);
or U7947 (N_7947,N_7711,N_7799);
nor U7948 (N_7948,N_7729,N_7743);
xor U7949 (N_7949,N_7783,N_7679);
nor U7950 (N_7950,N_7729,N_7638);
nor U7951 (N_7951,N_7666,N_7739);
or U7952 (N_7952,N_7624,N_7799);
nor U7953 (N_7953,N_7763,N_7614);
and U7954 (N_7954,N_7669,N_7700);
nor U7955 (N_7955,N_7778,N_7716);
nor U7956 (N_7956,N_7620,N_7740);
nand U7957 (N_7957,N_7775,N_7719);
and U7958 (N_7958,N_7747,N_7653);
nand U7959 (N_7959,N_7630,N_7644);
or U7960 (N_7960,N_7698,N_7750);
or U7961 (N_7961,N_7718,N_7776);
and U7962 (N_7962,N_7697,N_7635);
and U7963 (N_7963,N_7759,N_7677);
and U7964 (N_7964,N_7720,N_7794);
and U7965 (N_7965,N_7691,N_7624);
or U7966 (N_7966,N_7692,N_7610);
nand U7967 (N_7967,N_7697,N_7650);
nand U7968 (N_7968,N_7709,N_7744);
nor U7969 (N_7969,N_7642,N_7751);
or U7970 (N_7970,N_7740,N_7658);
nand U7971 (N_7971,N_7780,N_7672);
and U7972 (N_7972,N_7724,N_7630);
or U7973 (N_7973,N_7610,N_7670);
xor U7974 (N_7974,N_7718,N_7626);
nand U7975 (N_7975,N_7756,N_7655);
xnor U7976 (N_7976,N_7733,N_7710);
nor U7977 (N_7977,N_7754,N_7605);
and U7978 (N_7978,N_7640,N_7628);
and U7979 (N_7979,N_7677,N_7725);
xor U7980 (N_7980,N_7646,N_7792);
or U7981 (N_7981,N_7657,N_7734);
nor U7982 (N_7982,N_7680,N_7646);
or U7983 (N_7983,N_7724,N_7703);
nand U7984 (N_7984,N_7749,N_7601);
nand U7985 (N_7985,N_7757,N_7608);
xor U7986 (N_7986,N_7613,N_7672);
xnor U7987 (N_7987,N_7752,N_7724);
xnor U7988 (N_7988,N_7696,N_7636);
or U7989 (N_7989,N_7650,N_7730);
or U7990 (N_7990,N_7655,N_7678);
nor U7991 (N_7991,N_7612,N_7610);
nor U7992 (N_7992,N_7732,N_7654);
nand U7993 (N_7993,N_7621,N_7613);
and U7994 (N_7994,N_7753,N_7729);
xnor U7995 (N_7995,N_7628,N_7789);
or U7996 (N_7996,N_7799,N_7712);
nor U7997 (N_7997,N_7739,N_7673);
and U7998 (N_7998,N_7747,N_7739);
or U7999 (N_7999,N_7728,N_7644);
xnor U8000 (N_8000,N_7914,N_7879);
xor U8001 (N_8001,N_7943,N_7971);
and U8002 (N_8002,N_7855,N_7836);
and U8003 (N_8003,N_7816,N_7933);
and U8004 (N_8004,N_7987,N_7944);
xnor U8005 (N_8005,N_7883,N_7962);
nand U8006 (N_8006,N_7911,N_7957);
nor U8007 (N_8007,N_7849,N_7876);
xnor U8008 (N_8008,N_7824,N_7845);
xor U8009 (N_8009,N_7959,N_7838);
or U8010 (N_8010,N_7837,N_7819);
and U8011 (N_8011,N_7830,N_7897);
or U8012 (N_8012,N_7844,N_7878);
nor U8013 (N_8013,N_7827,N_7823);
nand U8014 (N_8014,N_7865,N_7867);
xnor U8015 (N_8015,N_7986,N_7997);
nor U8016 (N_8016,N_7817,N_7941);
xor U8017 (N_8017,N_7832,N_7800);
nor U8018 (N_8018,N_7809,N_7864);
xnor U8019 (N_8019,N_7893,N_7952);
or U8020 (N_8020,N_7834,N_7811);
xor U8021 (N_8021,N_7961,N_7805);
and U8022 (N_8022,N_7906,N_7821);
and U8023 (N_8023,N_7991,N_7826);
xnor U8024 (N_8024,N_7807,N_7888);
xor U8025 (N_8025,N_7982,N_7940);
xor U8026 (N_8026,N_7927,N_7998);
or U8027 (N_8027,N_7868,N_7907);
nand U8028 (N_8028,N_7917,N_7808);
and U8029 (N_8029,N_7963,N_7995);
nand U8030 (N_8030,N_7956,N_7992);
xnor U8031 (N_8031,N_7895,N_7901);
nor U8032 (N_8032,N_7884,N_7846);
or U8033 (N_8033,N_7885,N_7916);
xnor U8034 (N_8034,N_7904,N_7835);
and U8035 (N_8035,N_7890,N_7841);
and U8036 (N_8036,N_7825,N_7881);
nand U8037 (N_8037,N_7951,N_7905);
nand U8038 (N_8038,N_7856,N_7833);
nor U8039 (N_8039,N_7934,N_7980);
nor U8040 (N_8040,N_7978,N_7908);
nor U8041 (N_8041,N_7975,N_7863);
or U8042 (N_8042,N_7853,N_7814);
and U8043 (N_8043,N_7938,N_7960);
or U8044 (N_8044,N_7994,N_7874);
and U8045 (N_8045,N_7894,N_7887);
xnor U8046 (N_8046,N_7953,N_7964);
and U8047 (N_8047,N_7872,N_7926);
or U8048 (N_8048,N_7966,N_7913);
xor U8049 (N_8049,N_7965,N_7851);
nand U8050 (N_8050,N_7810,N_7985);
or U8051 (N_8051,N_7979,N_7948);
and U8052 (N_8052,N_7939,N_7873);
or U8053 (N_8053,N_7972,N_7974);
xnor U8054 (N_8054,N_7892,N_7869);
nand U8055 (N_8055,N_7932,N_7918);
nand U8056 (N_8056,N_7988,N_7920);
nand U8057 (N_8057,N_7896,N_7942);
and U8058 (N_8058,N_7928,N_7950);
and U8059 (N_8059,N_7839,N_7970);
or U8060 (N_8060,N_7822,N_7949);
and U8061 (N_8061,N_7870,N_7871);
nand U8062 (N_8062,N_7898,N_7945);
and U8063 (N_8063,N_7858,N_7983);
nor U8064 (N_8064,N_7804,N_7806);
or U8065 (N_8065,N_7848,N_7921);
nand U8066 (N_8066,N_7912,N_7860);
xor U8067 (N_8067,N_7947,N_7925);
and U8068 (N_8068,N_7857,N_7854);
and U8069 (N_8069,N_7954,N_7996);
xor U8070 (N_8070,N_7803,N_7910);
or U8071 (N_8071,N_7984,N_7900);
or U8072 (N_8072,N_7882,N_7877);
xor U8073 (N_8073,N_7842,N_7831);
xor U8074 (N_8074,N_7958,N_7875);
xor U8075 (N_8075,N_7802,N_7899);
nand U8076 (N_8076,N_7955,N_7852);
nor U8077 (N_8077,N_7866,N_7989);
nand U8078 (N_8078,N_7843,N_7936);
nor U8079 (N_8079,N_7930,N_7993);
nand U8080 (N_8080,N_7880,N_7915);
xor U8081 (N_8081,N_7861,N_7840);
xnor U8082 (N_8082,N_7967,N_7922);
and U8083 (N_8083,N_7862,N_7981);
xor U8084 (N_8084,N_7847,N_7999);
xor U8085 (N_8085,N_7923,N_7815);
or U8086 (N_8086,N_7903,N_7976);
nor U8087 (N_8087,N_7891,N_7969);
xor U8088 (N_8088,N_7924,N_7889);
nor U8089 (N_8089,N_7829,N_7973);
and U8090 (N_8090,N_7812,N_7818);
nand U8091 (N_8091,N_7937,N_7929);
nor U8092 (N_8092,N_7828,N_7935);
xnor U8093 (N_8093,N_7968,N_7990);
or U8094 (N_8094,N_7919,N_7813);
nand U8095 (N_8095,N_7886,N_7977);
and U8096 (N_8096,N_7801,N_7902);
and U8097 (N_8097,N_7820,N_7909);
nor U8098 (N_8098,N_7931,N_7850);
nor U8099 (N_8099,N_7859,N_7946);
nor U8100 (N_8100,N_7932,N_7837);
and U8101 (N_8101,N_7857,N_7981);
nor U8102 (N_8102,N_7901,N_7873);
xnor U8103 (N_8103,N_7895,N_7855);
and U8104 (N_8104,N_7992,N_7857);
xnor U8105 (N_8105,N_7897,N_7915);
or U8106 (N_8106,N_7832,N_7917);
nor U8107 (N_8107,N_7989,N_7874);
and U8108 (N_8108,N_7903,N_7978);
and U8109 (N_8109,N_7860,N_7934);
nand U8110 (N_8110,N_7844,N_7812);
nor U8111 (N_8111,N_7841,N_7861);
nand U8112 (N_8112,N_7805,N_7871);
or U8113 (N_8113,N_7818,N_7868);
and U8114 (N_8114,N_7851,N_7922);
or U8115 (N_8115,N_7937,N_7933);
nor U8116 (N_8116,N_7888,N_7923);
xor U8117 (N_8117,N_7889,N_7835);
xor U8118 (N_8118,N_7813,N_7992);
and U8119 (N_8119,N_7924,N_7822);
nor U8120 (N_8120,N_7963,N_7807);
nand U8121 (N_8121,N_7984,N_7907);
xnor U8122 (N_8122,N_7802,N_7827);
and U8123 (N_8123,N_7949,N_7859);
and U8124 (N_8124,N_7841,N_7870);
nor U8125 (N_8125,N_7817,N_7848);
nor U8126 (N_8126,N_7838,N_7989);
xor U8127 (N_8127,N_7883,N_7945);
nor U8128 (N_8128,N_7823,N_7922);
xor U8129 (N_8129,N_7886,N_7976);
nor U8130 (N_8130,N_7967,N_7899);
nor U8131 (N_8131,N_7826,N_7888);
xor U8132 (N_8132,N_7881,N_7987);
or U8133 (N_8133,N_7822,N_7937);
and U8134 (N_8134,N_7999,N_7883);
xor U8135 (N_8135,N_7805,N_7842);
or U8136 (N_8136,N_7910,N_7957);
and U8137 (N_8137,N_7901,N_7976);
or U8138 (N_8138,N_7814,N_7832);
nor U8139 (N_8139,N_7859,N_7927);
or U8140 (N_8140,N_7947,N_7943);
nor U8141 (N_8141,N_7995,N_7844);
nor U8142 (N_8142,N_7948,N_7893);
nand U8143 (N_8143,N_7910,N_7886);
and U8144 (N_8144,N_7954,N_7801);
nand U8145 (N_8145,N_7832,N_7860);
and U8146 (N_8146,N_7831,N_7896);
or U8147 (N_8147,N_7934,N_7887);
or U8148 (N_8148,N_7814,N_7951);
xnor U8149 (N_8149,N_7886,N_7919);
and U8150 (N_8150,N_7853,N_7988);
and U8151 (N_8151,N_7917,N_7915);
nor U8152 (N_8152,N_7951,N_7989);
nor U8153 (N_8153,N_7936,N_7998);
nor U8154 (N_8154,N_7812,N_7824);
nor U8155 (N_8155,N_7992,N_7920);
nand U8156 (N_8156,N_7872,N_7896);
xnor U8157 (N_8157,N_7808,N_7939);
nor U8158 (N_8158,N_7807,N_7961);
and U8159 (N_8159,N_7800,N_7908);
nand U8160 (N_8160,N_7835,N_7891);
xnor U8161 (N_8161,N_7853,N_7968);
nand U8162 (N_8162,N_7835,N_7993);
or U8163 (N_8163,N_7811,N_7827);
or U8164 (N_8164,N_7823,N_7880);
or U8165 (N_8165,N_7933,N_7849);
or U8166 (N_8166,N_7845,N_7916);
and U8167 (N_8167,N_7834,N_7853);
nand U8168 (N_8168,N_7856,N_7949);
nand U8169 (N_8169,N_7961,N_7915);
or U8170 (N_8170,N_7900,N_7874);
nand U8171 (N_8171,N_7898,N_7948);
nand U8172 (N_8172,N_7932,N_7870);
xnor U8173 (N_8173,N_7827,N_7883);
nor U8174 (N_8174,N_7979,N_7868);
and U8175 (N_8175,N_7911,N_7804);
or U8176 (N_8176,N_7858,N_7848);
or U8177 (N_8177,N_7885,N_7884);
and U8178 (N_8178,N_7873,N_7813);
xnor U8179 (N_8179,N_7987,N_7886);
nor U8180 (N_8180,N_7805,N_7807);
or U8181 (N_8181,N_7923,N_7860);
nor U8182 (N_8182,N_7847,N_7940);
nor U8183 (N_8183,N_7958,N_7959);
nor U8184 (N_8184,N_7913,N_7926);
nand U8185 (N_8185,N_7884,N_7839);
or U8186 (N_8186,N_7820,N_7915);
or U8187 (N_8187,N_7932,N_7813);
and U8188 (N_8188,N_7919,N_7991);
or U8189 (N_8189,N_7852,N_7901);
and U8190 (N_8190,N_7830,N_7958);
nand U8191 (N_8191,N_7903,N_7850);
and U8192 (N_8192,N_7816,N_7840);
and U8193 (N_8193,N_7881,N_7918);
nor U8194 (N_8194,N_7931,N_7963);
or U8195 (N_8195,N_7830,N_7937);
nor U8196 (N_8196,N_7825,N_7806);
and U8197 (N_8197,N_7945,N_7894);
and U8198 (N_8198,N_7984,N_7892);
nor U8199 (N_8199,N_7825,N_7974);
xnor U8200 (N_8200,N_8121,N_8072);
nand U8201 (N_8201,N_8026,N_8103);
xor U8202 (N_8202,N_8166,N_8064);
nor U8203 (N_8203,N_8015,N_8045);
xor U8204 (N_8204,N_8136,N_8177);
nand U8205 (N_8205,N_8046,N_8100);
and U8206 (N_8206,N_8194,N_8153);
or U8207 (N_8207,N_8092,N_8041);
or U8208 (N_8208,N_8089,N_8071);
or U8209 (N_8209,N_8066,N_8178);
xor U8210 (N_8210,N_8016,N_8059);
xnor U8211 (N_8211,N_8032,N_8101);
nor U8212 (N_8212,N_8138,N_8055);
xnor U8213 (N_8213,N_8165,N_8148);
nand U8214 (N_8214,N_8003,N_8083);
nor U8215 (N_8215,N_8102,N_8078);
and U8216 (N_8216,N_8181,N_8035);
nor U8217 (N_8217,N_8004,N_8063);
nand U8218 (N_8218,N_8118,N_8114);
nor U8219 (N_8219,N_8091,N_8110);
nand U8220 (N_8220,N_8030,N_8180);
nand U8221 (N_8221,N_8196,N_8008);
and U8222 (N_8222,N_8053,N_8157);
and U8223 (N_8223,N_8014,N_8124);
nand U8224 (N_8224,N_8172,N_8179);
xnor U8225 (N_8225,N_8067,N_8129);
or U8226 (N_8226,N_8060,N_8068);
or U8227 (N_8227,N_8189,N_8186);
nor U8228 (N_8228,N_8176,N_8077);
nand U8229 (N_8229,N_8022,N_8144);
or U8230 (N_8230,N_8141,N_8013);
nand U8231 (N_8231,N_8043,N_8169);
nand U8232 (N_8232,N_8161,N_8007);
nand U8233 (N_8233,N_8019,N_8048);
and U8234 (N_8234,N_8006,N_8074);
and U8235 (N_8235,N_8168,N_8096);
xnor U8236 (N_8236,N_8106,N_8122);
and U8237 (N_8237,N_8088,N_8198);
nand U8238 (N_8238,N_8054,N_8162);
or U8239 (N_8239,N_8051,N_8012);
or U8240 (N_8240,N_8135,N_8057);
xor U8241 (N_8241,N_8164,N_8084);
and U8242 (N_8242,N_8197,N_8065);
and U8243 (N_8243,N_8159,N_8037);
xnor U8244 (N_8244,N_8115,N_8143);
and U8245 (N_8245,N_8107,N_8123);
xnor U8246 (N_8246,N_8093,N_8131);
and U8247 (N_8247,N_8052,N_8005);
or U8248 (N_8248,N_8024,N_8020);
or U8249 (N_8249,N_8113,N_8021);
or U8250 (N_8250,N_8128,N_8011);
or U8251 (N_8251,N_8191,N_8098);
xnor U8252 (N_8252,N_8025,N_8170);
xnor U8253 (N_8253,N_8152,N_8192);
xnor U8254 (N_8254,N_8033,N_8139);
and U8255 (N_8255,N_8105,N_8119);
and U8256 (N_8256,N_8151,N_8116);
nor U8257 (N_8257,N_8183,N_8187);
and U8258 (N_8258,N_8023,N_8109);
nor U8259 (N_8259,N_8185,N_8050);
xnor U8260 (N_8260,N_8079,N_8049);
xor U8261 (N_8261,N_8167,N_8097);
nand U8262 (N_8262,N_8156,N_8018);
or U8263 (N_8263,N_8146,N_8163);
xnor U8264 (N_8264,N_8087,N_8058);
xor U8265 (N_8265,N_8062,N_8145);
xnor U8266 (N_8266,N_8160,N_8171);
nand U8267 (N_8267,N_8133,N_8134);
or U8268 (N_8268,N_8081,N_8061);
nand U8269 (N_8269,N_8154,N_8042);
and U8270 (N_8270,N_8111,N_8056);
nor U8271 (N_8271,N_8044,N_8190);
and U8272 (N_8272,N_8127,N_8099);
xnor U8273 (N_8273,N_8070,N_8104);
or U8274 (N_8274,N_8150,N_8142);
nand U8275 (N_8275,N_8080,N_8094);
nand U8276 (N_8276,N_8175,N_8010);
xnor U8277 (N_8277,N_8195,N_8090);
xor U8278 (N_8278,N_8085,N_8149);
xnor U8279 (N_8279,N_8188,N_8073);
nand U8280 (N_8280,N_8147,N_8029);
xor U8281 (N_8281,N_8038,N_8193);
nor U8282 (N_8282,N_8112,N_8155);
xnor U8283 (N_8283,N_8001,N_8182);
nand U8284 (N_8284,N_8076,N_8158);
nor U8285 (N_8285,N_8027,N_8017);
nand U8286 (N_8286,N_8125,N_8184);
xnor U8287 (N_8287,N_8126,N_8137);
xnor U8288 (N_8288,N_8120,N_8117);
nand U8289 (N_8289,N_8095,N_8108);
xor U8290 (N_8290,N_8036,N_8002);
xnor U8291 (N_8291,N_8174,N_8075);
nand U8292 (N_8292,N_8199,N_8130);
or U8293 (N_8293,N_8000,N_8034);
and U8294 (N_8294,N_8132,N_8028);
xor U8295 (N_8295,N_8040,N_8086);
or U8296 (N_8296,N_8173,N_8140);
xnor U8297 (N_8297,N_8082,N_8039);
and U8298 (N_8298,N_8031,N_8069);
nand U8299 (N_8299,N_8047,N_8009);
nor U8300 (N_8300,N_8082,N_8194);
xor U8301 (N_8301,N_8100,N_8055);
nor U8302 (N_8302,N_8168,N_8138);
xor U8303 (N_8303,N_8112,N_8016);
nor U8304 (N_8304,N_8128,N_8117);
xnor U8305 (N_8305,N_8141,N_8047);
nor U8306 (N_8306,N_8105,N_8172);
nand U8307 (N_8307,N_8106,N_8169);
nor U8308 (N_8308,N_8023,N_8085);
or U8309 (N_8309,N_8074,N_8099);
xnor U8310 (N_8310,N_8082,N_8115);
or U8311 (N_8311,N_8044,N_8194);
nand U8312 (N_8312,N_8171,N_8101);
or U8313 (N_8313,N_8182,N_8039);
xor U8314 (N_8314,N_8191,N_8044);
and U8315 (N_8315,N_8042,N_8090);
or U8316 (N_8316,N_8105,N_8124);
and U8317 (N_8317,N_8073,N_8183);
nand U8318 (N_8318,N_8004,N_8008);
nor U8319 (N_8319,N_8174,N_8113);
or U8320 (N_8320,N_8178,N_8026);
nor U8321 (N_8321,N_8122,N_8165);
or U8322 (N_8322,N_8093,N_8172);
nor U8323 (N_8323,N_8126,N_8099);
and U8324 (N_8324,N_8056,N_8023);
nand U8325 (N_8325,N_8136,N_8125);
or U8326 (N_8326,N_8120,N_8070);
nor U8327 (N_8327,N_8001,N_8087);
nor U8328 (N_8328,N_8001,N_8006);
or U8329 (N_8329,N_8176,N_8168);
and U8330 (N_8330,N_8006,N_8180);
nand U8331 (N_8331,N_8198,N_8186);
nor U8332 (N_8332,N_8199,N_8106);
nor U8333 (N_8333,N_8101,N_8130);
nand U8334 (N_8334,N_8050,N_8082);
nand U8335 (N_8335,N_8123,N_8011);
xnor U8336 (N_8336,N_8174,N_8015);
or U8337 (N_8337,N_8121,N_8168);
and U8338 (N_8338,N_8004,N_8199);
or U8339 (N_8339,N_8147,N_8069);
and U8340 (N_8340,N_8128,N_8181);
nand U8341 (N_8341,N_8186,N_8143);
xnor U8342 (N_8342,N_8087,N_8064);
nor U8343 (N_8343,N_8190,N_8090);
or U8344 (N_8344,N_8043,N_8074);
and U8345 (N_8345,N_8005,N_8006);
nor U8346 (N_8346,N_8087,N_8091);
nand U8347 (N_8347,N_8091,N_8096);
and U8348 (N_8348,N_8122,N_8000);
xor U8349 (N_8349,N_8034,N_8110);
nor U8350 (N_8350,N_8043,N_8123);
xnor U8351 (N_8351,N_8075,N_8140);
nand U8352 (N_8352,N_8123,N_8064);
xnor U8353 (N_8353,N_8017,N_8154);
or U8354 (N_8354,N_8030,N_8039);
and U8355 (N_8355,N_8068,N_8007);
xor U8356 (N_8356,N_8167,N_8008);
or U8357 (N_8357,N_8174,N_8029);
or U8358 (N_8358,N_8111,N_8172);
or U8359 (N_8359,N_8161,N_8148);
nand U8360 (N_8360,N_8023,N_8107);
and U8361 (N_8361,N_8026,N_8068);
or U8362 (N_8362,N_8122,N_8031);
nor U8363 (N_8363,N_8114,N_8160);
nand U8364 (N_8364,N_8186,N_8137);
nor U8365 (N_8365,N_8032,N_8134);
nand U8366 (N_8366,N_8153,N_8189);
nand U8367 (N_8367,N_8177,N_8061);
and U8368 (N_8368,N_8153,N_8165);
or U8369 (N_8369,N_8117,N_8061);
and U8370 (N_8370,N_8036,N_8123);
nor U8371 (N_8371,N_8054,N_8006);
xnor U8372 (N_8372,N_8040,N_8129);
or U8373 (N_8373,N_8081,N_8106);
xor U8374 (N_8374,N_8197,N_8014);
nor U8375 (N_8375,N_8187,N_8003);
and U8376 (N_8376,N_8097,N_8074);
or U8377 (N_8377,N_8105,N_8082);
or U8378 (N_8378,N_8186,N_8171);
nand U8379 (N_8379,N_8103,N_8014);
nand U8380 (N_8380,N_8051,N_8139);
and U8381 (N_8381,N_8054,N_8130);
or U8382 (N_8382,N_8198,N_8106);
and U8383 (N_8383,N_8059,N_8063);
or U8384 (N_8384,N_8170,N_8069);
and U8385 (N_8385,N_8171,N_8028);
and U8386 (N_8386,N_8156,N_8183);
and U8387 (N_8387,N_8009,N_8167);
xor U8388 (N_8388,N_8036,N_8100);
or U8389 (N_8389,N_8029,N_8036);
or U8390 (N_8390,N_8012,N_8189);
and U8391 (N_8391,N_8116,N_8181);
nand U8392 (N_8392,N_8023,N_8027);
and U8393 (N_8393,N_8086,N_8097);
xnor U8394 (N_8394,N_8106,N_8056);
nand U8395 (N_8395,N_8068,N_8028);
and U8396 (N_8396,N_8115,N_8033);
nor U8397 (N_8397,N_8162,N_8025);
or U8398 (N_8398,N_8137,N_8175);
and U8399 (N_8399,N_8197,N_8049);
nor U8400 (N_8400,N_8390,N_8269);
and U8401 (N_8401,N_8253,N_8371);
and U8402 (N_8402,N_8359,N_8207);
and U8403 (N_8403,N_8339,N_8388);
nand U8404 (N_8404,N_8322,N_8232);
nor U8405 (N_8405,N_8356,N_8396);
or U8406 (N_8406,N_8330,N_8280);
or U8407 (N_8407,N_8291,N_8226);
nand U8408 (N_8408,N_8398,N_8294);
or U8409 (N_8409,N_8346,N_8315);
and U8410 (N_8410,N_8362,N_8209);
xnor U8411 (N_8411,N_8320,N_8235);
nand U8412 (N_8412,N_8213,N_8336);
nor U8413 (N_8413,N_8224,N_8313);
xnor U8414 (N_8414,N_8208,N_8205);
nor U8415 (N_8415,N_8278,N_8331);
or U8416 (N_8416,N_8355,N_8364);
or U8417 (N_8417,N_8317,N_8361);
or U8418 (N_8418,N_8251,N_8324);
and U8419 (N_8419,N_8289,N_8379);
nor U8420 (N_8420,N_8263,N_8271);
or U8421 (N_8421,N_8333,N_8395);
nand U8422 (N_8422,N_8214,N_8329);
and U8423 (N_8423,N_8301,N_8340);
nor U8424 (N_8424,N_8374,N_8257);
nand U8425 (N_8425,N_8375,N_8350);
xor U8426 (N_8426,N_8286,N_8325);
nand U8427 (N_8427,N_8391,N_8200);
and U8428 (N_8428,N_8243,N_8316);
nand U8429 (N_8429,N_8268,N_8255);
and U8430 (N_8430,N_8277,N_8247);
and U8431 (N_8431,N_8245,N_8399);
nand U8432 (N_8432,N_8272,N_8292);
or U8433 (N_8433,N_8264,N_8354);
or U8434 (N_8434,N_8326,N_8260);
or U8435 (N_8435,N_8394,N_8385);
xnor U8436 (N_8436,N_8293,N_8261);
xor U8437 (N_8437,N_8380,N_8341);
xnor U8438 (N_8438,N_8363,N_8296);
or U8439 (N_8439,N_8229,N_8281);
and U8440 (N_8440,N_8351,N_8382);
xor U8441 (N_8441,N_8206,N_8332);
or U8442 (N_8442,N_8383,N_8344);
xor U8443 (N_8443,N_8220,N_8233);
nor U8444 (N_8444,N_8276,N_8254);
nor U8445 (N_8445,N_8231,N_8303);
nand U8446 (N_8446,N_8307,N_8347);
or U8447 (N_8447,N_8310,N_8252);
nand U8448 (N_8448,N_8211,N_8241);
nand U8449 (N_8449,N_8262,N_8397);
or U8450 (N_8450,N_8216,N_8290);
or U8451 (N_8451,N_8321,N_8323);
nor U8452 (N_8452,N_8284,N_8210);
and U8453 (N_8453,N_8314,N_8370);
xnor U8454 (N_8454,N_8393,N_8308);
or U8455 (N_8455,N_8368,N_8228);
or U8456 (N_8456,N_8256,N_8360);
xor U8457 (N_8457,N_8299,N_8223);
xor U8458 (N_8458,N_8345,N_8297);
nor U8459 (N_8459,N_8352,N_8369);
nand U8460 (N_8460,N_8300,N_8239);
or U8461 (N_8461,N_8236,N_8295);
and U8462 (N_8462,N_8338,N_8377);
and U8463 (N_8463,N_8240,N_8217);
xnor U8464 (N_8464,N_8367,N_8203);
and U8465 (N_8465,N_8378,N_8201);
xnor U8466 (N_8466,N_8312,N_8365);
and U8467 (N_8467,N_8334,N_8244);
or U8468 (N_8468,N_8304,N_8282);
nand U8469 (N_8469,N_8234,N_8242);
and U8470 (N_8470,N_8267,N_8249);
nor U8471 (N_8471,N_8238,N_8221);
nor U8472 (N_8472,N_8298,N_8342);
xor U8473 (N_8473,N_8204,N_8202);
nand U8474 (N_8474,N_8358,N_8285);
nor U8475 (N_8475,N_8337,N_8353);
nor U8476 (N_8476,N_8265,N_8215);
nand U8477 (N_8477,N_8250,N_8230);
xor U8478 (N_8478,N_8237,N_8246);
or U8479 (N_8479,N_8318,N_8283);
nor U8480 (N_8480,N_8335,N_8381);
nor U8481 (N_8481,N_8259,N_8389);
or U8482 (N_8482,N_8349,N_8366);
and U8483 (N_8483,N_8386,N_8387);
nor U8484 (N_8484,N_8273,N_8258);
xor U8485 (N_8485,N_8219,N_8279);
xor U8486 (N_8486,N_8225,N_8376);
nand U8487 (N_8487,N_8343,N_8372);
and U8488 (N_8488,N_8227,N_8328);
and U8489 (N_8489,N_8306,N_8274);
and U8490 (N_8490,N_8248,N_8392);
and U8491 (N_8491,N_8348,N_8288);
nand U8492 (N_8492,N_8319,N_8357);
or U8493 (N_8493,N_8384,N_8373);
xor U8494 (N_8494,N_8327,N_8302);
nand U8495 (N_8495,N_8311,N_8309);
nor U8496 (N_8496,N_8218,N_8222);
xor U8497 (N_8497,N_8212,N_8270);
nand U8498 (N_8498,N_8266,N_8275);
xor U8499 (N_8499,N_8287,N_8305);
xnor U8500 (N_8500,N_8263,N_8293);
xnor U8501 (N_8501,N_8274,N_8367);
and U8502 (N_8502,N_8298,N_8334);
nor U8503 (N_8503,N_8286,N_8323);
nand U8504 (N_8504,N_8320,N_8313);
and U8505 (N_8505,N_8300,N_8282);
and U8506 (N_8506,N_8365,N_8212);
xnor U8507 (N_8507,N_8379,N_8237);
and U8508 (N_8508,N_8299,N_8246);
or U8509 (N_8509,N_8287,N_8388);
or U8510 (N_8510,N_8209,N_8335);
nor U8511 (N_8511,N_8302,N_8291);
xor U8512 (N_8512,N_8325,N_8354);
and U8513 (N_8513,N_8312,N_8202);
nand U8514 (N_8514,N_8241,N_8355);
nor U8515 (N_8515,N_8361,N_8314);
and U8516 (N_8516,N_8313,N_8384);
and U8517 (N_8517,N_8213,N_8256);
nor U8518 (N_8518,N_8207,N_8380);
or U8519 (N_8519,N_8203,N_8399);
or U8520 (N_8520,N_8343,N_8234);
xnor U8521 (N_8521,N_8231,N_8221);
xnor U8522 (N_8522,N_8272,N_8377);
and U8523 (N_8523,N_8301,N_8218);
nand U8524 (N_8524,N_8202,N_8337);
nor U8525 (N_8525,N_8381,N_8376);
xor U8526 (N_8526,N_8296,N_8232);
and U8527 (N_8527,N_8327,N_8273);
nand U8528 (N_8528,N_8254,N_8356);
or U8529 (N_8529,N_8349,N_8378);
nand U8530 (N_8530,N_8326,N_8217);
xnor U8531 (N_8531,N_8397,N_8209);
or U8532 (N_8532,N_8257,N_8369);
and U8533 (N_8533,N_8359,N_8302);
or U8534 (N_8534,N_8288,N_8347);
nand U8535 (N_8535,N_8238,N_8260);
and U8536 (N_8536,N_8222,N_8337);
or U8537 (N_8537,N_8250,N_8267);
and U8538 (N_8538,N_8205,N_8261);
or U8539 (N_8539,N_8234,N_8337);
and U8540 (N_8540,N_8320,N_8262);
nand U8541 (N_8541,N_8289,N_8370);
nand U8542 (N_8542,N_8379,N_8340);
xnor U8543 (N_8543,N_8258,N_8337);
and U8544 (N_8544,N_8221,N_8342);
xor U8545 (N_8545,N_8259,N_8252);
nand U8546 (N_8546,N_8342,N_8305);
or U8547 (N_8547,N_8326,N_8371);
or U8548 (N_8548,N_8218,N_8368);
nand U8549 (N_8549,N_8278,N_8296);
xor U8550 (N_8550,N_8309,N_8396);
nor U8551 (N_8551,N_8361,N_8217);
and U8552 (N_8552,N_8219,N_8370);
nor U8553 (N_8553,N_8351,N_8376);
nand U8554 (N_8554,N_8335,N_8232);
or U8555 (N_8555,N_8327,N_8334);
or U8556 (N_8556,N_8229,N_8237);
or U8557 (N_8557,N_8339,N_8321);
nand U8558 (N_8558,N_8282,N_8246);
nor U8559 (N_8559,N_8295,N_8293);
and U8560 (N_8560,N_8399,N_8273);
nand U8561 (N_8561,N_8249,N_8212);
and U8562 (N_8562,N_8282,N_8258);
nand U8563 (N_8563,N_8251,N_8240);
nor U8564 (N_8564,N_8357,N_8381);
or U8565 (N_8565,N_8214,N_8327);
nor U8566 (N_8566,N_8398,N_8317);
and U8567 (N_8567,N_8258,N_8360);
xnor U8568 (N_8568,N_8392,N_8275);
nand U8569 (N_8569,N_8277,N_8367);
and U8570 (N_8570,N_8206,N_8211);
nor U8571 (N_8571,N_8306,N_8203);
nand U8572 (N_8572,N_8340,N_8231);
nor U8573 (N_8573,N_8240,N_8218);
and U8574 (N_8574,N_8300,N_8381);
nand U8575 (N_8575,N_8383,N_8311);
xor U8576 (N_8576,N_8327,N_8270);
nand U8577 (N_8577,N_8381,N_8382);
or U8578 (N_8578,N_8296,N_8325);
or U8579 (N_8579,N_8257,N_8287);
and U8580 (N_8580,N_8202,N_8398);
nand U8581 (N_8581,N_8230,N_8321);
xor U8582 (N_8582,N_8399,N_8330);
or U8583 (N_8583,N_8367,N_8223);
nand U8584 (N_8584,N_8248,N_8200);
nor U8585 (N_8585,N_8264,N_8339);
nor U8586 (N_8586,N_8253,N_8357);
or U8587 (N_8587,N_8361,N_8323);
nand U8588 (N_8588,N_8331,N_8388);
nand U8589 (N_8589,N_8362,N_8227);
and U8590 (N_8590,N_8244,N_8380);
or U8591 (N_8591,N_8325,N_8201);
or U8592 (N_8592,N_8301,N_8332);
nor U8593 (N_8593,N_8366,N_8342);
xnor U8594 (N_8594,N_8259,N_8292);
nand U8595 (N_8595,N_8224,N_8328);
nand U8596 (N_8596,N_8256,N_8384);
nand U8597 (N_8597,N_8396,N_8351);
nand U8598 (N_8598,N_8311,N_8357);
nor U8599 (N_8599,N_8340,N_8367);
nand U8600 (N_8600,N_8475,N_8581);
nand U8601 (N_8601,N_8479,N_8425);
xnor U8602 (N_8602,N_8582,N_8433);
xnor U8603 (N_8603,N_8457,N_8494);
and U8604 (N_8604,N_8504,N_8445);
or U8605 (N_8605,N_8472,N_8554);
xnor U8606 (N_8606,N_8573,N_8567);
or U8607 (N_8607,N_8420,N_8414);
or U8608 (N_8608,N_8590,N_8577);
nand U8609 (N_8609,N_8421,N_8415);
and U8610 (N_8610,N_8438,N_8597);
nand U8611 (N_8611,N_8505,N_8436);
nor U8612 (N_8612,N_8535,N_8448);
nor U8613 (N_8613,N_8403,N_8464);
and U8614 (N_8614,N_8422,N_8442);
nand U8615 (N_8615,N_8585,N_8508);
and U8616 (N_8616,N_8496,N_8480);
or U8617 (N_8617,N_8419,N_8406);
xnor U8618 (N_8618,N_8503,N_8506);
nor U8619 (N_8619,N_8551,N_8450);
or U8620 (N_8620,N_8588,N_8560);
xnor U8621 (N_8621,N_8435,N_8532);
nor U8622 (N_8622,N_8591,N_8434);
nor U8623 (N_8623,N_8437,N_8466);
and U8624 (N_8624,N_8507,N_8525);
nand U8625 (N_8625,N_8424,N_8463);
or U8626 (N_8626,N_8538,N_8524);
xor U8627 (N_8627,N_8510,N_8492);
nor U8628 (N_8628,N_8489,N_8498);
and U8629 (N_8629,N_8493,N_8586);
nor U8630 (N_8630,N_8543,N_8574);
and U8631 (N_8631,N_8520,N_8515);
xor U8632 (N_8632,N_8537,N_8594);
nor U8633 (N_8633,N_8502,N_8474);
or U8634 (N_8634,N_8404,N_8556);
or U8635 (N_8635,N_8485,N_8584);
and U8636 (N_8636,N_8471,N_8553);
nand U8637 (N_8637,N_8456,N_8558);
nand U8638 (N_8638,N_8576,N_8561);
or U8639 (N_8639,N_8495,N_8454);
xnor U8640 (N_8640,N_8418,N_8447);
nor U8641 (N_8641,N_8478,N_8411);
or U8642 (N_8642,N_8444,N_8570);
nor U8643 (N_8643,N_8511,N_8522);
nand U8644 (N_8644,N_8429,N_8530);
nand U8645 (N_8645,N_8539,N_8579);
and U8646 (N_8646,N_8559,N_8548);
and U8647 (N_8647,N_8417,N_8509);
nor U8648 (N_8648,N_8544,N_8428);
xnor U8649 (N_8649,N_8545,N_8483);
xnor U8650 (N_8650,N_8441,N_8516);
nand U8651 (N_8651,N_8512,N_8455);
or U8652 (N_8652,N_8439,N_8410);
nand U8653 (N_8653,N_8491,N_8443);
xor U8654 (N_8654,N_8488,N_8527);
or U8655 (N_8655,N_8465,N_8462);
and U8656 (N_8656,N_8555,N_8523);
xor U8657 (N_8657,N_8592,N_8552);
and U8658 (N_8658,N_8427,N_8533);
nor U8659 (N_8659,N_8446,N_8587);
or U8660 (N_8660,N_8426,N_8568);
nor U8661 (N_8661,N_8598,N_8557);
and U8662 (N_8662,N_8536,N_8534);
xnor U8663 (N_8663,N_8470,N_8497);
xnor U8664 (N_8664,N_8550,N_8423);
xor U8665 (N_8665,N_8432,N_8487);
xnor U8666 (N_8666,N_8514,N_8407);
xor U8667 (N_8667,N_8566,N_8580);
or U8668 (N_8668,N_8440,N_8546);
xor U8669 (N_8669,N_8499,N_8563);
or U8670 (N_8670,N_8569,N_8468);
nor U8671 (N_8671,N_8542,N_8431);
nor U8672 (N_8672,N_8521,N_8461);
or U8673 (N_8673,N_8481,N_8412);
nand U8674 (N_8674,N_8408,N_8564);
or U8675 (N_8675,N_8578,N_8540);
nor U8676 (N_8676,N_8575,N_8565);
and U8677 (N_8677,N_8413,N_8409);
nor U8678 (N_8678,N_8467,N_8596);
or U8679 (N_8679,N_8595,N_8400);
nand U8680 (N_8680,N_8547,N_8541);
xnor U8681 (N_8681,N_8529,N_8453);
nand U8682 (N_8682,N_8519,N_8531);
nand U8683 (N_8683,N_8599,N_8486);
and U8684 (N_8684,N_8458,N_8482);
nor U8685 (N_8685,N_8500,N_8416);
nand U8686 (N_8686,N_8484,N_8460);
or U8687 (N_8687,N_8402,N_8526);
nor U8688 (N_8688,N_8469,N_8589);
and U8689 (N_8689,N_8513,N_8430);
or U8690 (N_8690,N_8401,N_8477);
or U8691 (N_8691,N_8405,N_8562);
and U8692 (N_8692,N_8571,N_8459);
and U8693 (N_8693,N_8528,N_8593);
or U8694 (N_8694,N_8517,N_8549);
or U8695 (N_8695,N_8451,N_8449);
nand U8696 (N_8696,N_8583,N_8473);
nand U8697 (N_8697,N_8452,N_8518);
and U8698 (N_8698,N_8490,N_8501);
xor U8699 (N_8699,N_8572,N_8476);
nor U8700 (N_8700,N_8446,N_8562);
nor U8701 (N_8701,N_8434,N_8459);
and U8702 (N_8702,N_8530,N_8531);
xnor U8703 (N_8703,N_8441,N_8515);
nor U8704 (N_8704,N_8570,N_8578);
or U8705 (N_8705,N_8466,N_8554);
or U8706 (N_8706,N_8462,N_8551);
and U8707 (N_8707,N_8516,N_8445);
nand U8708 (N_8708,N_8414,N_8406);
nor U8709 (N_8709,N_8566,N_8500);
nand U8710 (N_8710,N_8595,N_8474);
nor U8711 (N_8711,N_8558,N_8421);
or U8712 (N_8712,N_8587,N_8530);
xor U8713 (N_8713,N_8416,N_8517);
or U8714 (N_8714,N_8452,N_8538);
nand U8715 (N_8715,N_8482,N_8406);
nand U8716 (N_8716,N_8512,N_8477);
nand U8717 (N_8717,N_8527,N_8443);
and U8718 (N_8718,N_8506,N_8492);
nor U8719 (N_8719,N_8513,N_8539);
or U8720 (N_8720,N_8449,N_8439);
and U8721 (N_8721,N_8437,N_8583);
xnor U8722 (N_8722,N_8521,N_8523);
nand U8723 (N_8723,N_8521,N_8538);
xnor U8724 (N_8724,N_8504,N_8477);
nor U8725 (N_8725,N_8519,N_8408);
and U8726 (N_8726,N_8555,N_8492);
nand U8727 (N_8727,N_8510,N_8431);
nor U8728 (N_8728,N_8420,N_8417);
xor U8729 (N_8729,N_8494,N_8420);
nand U8730 (N_8730,N_8472,N_8474);
xnor U8731 (N_8731,N_8540,N_8589);
and U8732 (N_8732,N_8538,N_8433);
and U8733 (N_8733,N_8428,N_8414);
and U8734 (N_8734,N_8445,N_8466);
or U8735 (N_8735,N_8553,N_8424);
or U8736 (N_8736,N_8499,N_8430);
and U8737 (N_8737,N_8592,N_8493);
nor U8738 (N_8738,N_8520,N_8420);
xnor U8739 (N_8739,N_8591,N_8587);
nand U8740 (N_8740,N_8593,N_8527);
nor U8741 (N_8741,N_8402,N_8531);
or U8742 (N_8742,N_8553,N_8512);
and U8743 (N_8743,N_8419,N_8594);
nor U8744 (N_8744,N_8532,N_8508);
and U8745 (N_8745,N_8485,N_8476);
nor U8746 (N_8746,N_8494,N_8486);
and U8747 (N_8747,N_8514,N_8549);
xor U8748 (N_8748,N_8514,N_8531);
or U8749 (N_8749,N_8572,N_8578);
nand U8750 (N_8750,N_8458,N_8504);
or U8751 (N_8751,N_8422,N_8427);
xnor U8752 (N_8752,N_8421,N_8593);
nor U8753 (N_8753,N_8535,N_8593);
and U8754 (N_8754,N_8472,N_8594);
nor U8755 (N_8755,N_8423,N_8594);
or U8756 (N_8756,N_8500,N_8580);
or U8757 (N_8757,N_8536,N_8496);
and U8758 (N_8758,N_8590,N_8504);
xor U8759 (N_8759,N_8461,N_8442);
nand U8760 (N_8760,N_8584,N_8419);
nor U8761 (N_8761,N_8566,N_8417);
nand U8762 (N_8762,N_8567,N_8480);
nor U8763 (N_8763,N_8558,N_8583);
xnor U8764 (N_8764,N_8470,N_8448);
nor U8765 (N_8765,N_8518,N_8440);
xor U8766 (N_8766,N_8421,N_8436);
xnor U8767 (N_8767,N_8514,N_8576);
nor U8768 (N_8768,N_8446,N_8501);
nand U8769 (N_8769,N_8409,N_8418);
and U8770 (N_8770,N_8423,N_8551);
or U8771 (N_8771,N_8416,N_8550);
nor U8772 (N_8772,N_8561,N_8450);
or U8773 (N_8773,N_8562,N_8597);
and U8774 (N_8774,N_8479,N_8523);
and U8775 (N_8775,N_8557,N_8568);
and U8776 (N_8776,N_8597,N_8491);
and U8777 (N_8777,N_8523,N_8576);
or U8778 (N_8778,N_8460,N_8481);
xor U8779 (N_8779,N_8492,N_8417);
nand U8780 (N_8780,N_8481,N_8506);
nor U8781 (N_8781,N_8456,N_8402);
nand U8782 (N_8782,N_8506,N_8442);
xor U8783 (N_8783,N_8441,N_8574);
nor U8784 (N_8784,N_8443,N_8468);
xnor U8785 (N_8785,N_8591,N_8529);
nand U8786 (N_8786,N_8454,N_8506);
nor U8787 (N_8787,N_8412,N_8500);
and U8788 (N_8788,N_8521,N_8463);
or U8789 (N_8789,N_8456,N_8430);
nor U8790 (N_8790,N_8486,N_8411);
and U8791 (N_8791,N_8508,N_8503);
xor U8792 (N_8792,N_8509,N_8578);
nand U8793 (N_8793,N_8506,N_8551);
or U8794 (N_8794,N_8448,N_8512);
nor U8795 (N_8795,N_8405,N_8456);
and U8796 (N_8796,N_8466,N_8497);
xor U8797 (N_8797,N_8472,N_8548);
and U8798 (N_8798,N_8501,N_8480);
nand U8799 (N_8799,N_8570,N_8562);
nor U8800 (N_8800,N_8797,N_8710);
or U8801 (N_8801,N_8672,N_8759);
or U8802 (N_8802,N_8754,N_8719);
nor U8803 (N_8803,N_8604,N_8784);
or U8804 (N_8804,N_8786,N_8724);
or U8805 (N_8805,N_8678,N_8736);
nor U8806 (N_8806,N_8634,N_8781);
nand U8807 (N_8807,N_8705,N_8645);
nand U8808 (N_8808,N_8639,N_8790);
nand U8809 (N_8809,N_8704,N_8727);
xnor U8810 (N_8810,N_8688,N_8668);
and U8811 (N_8811,N_8624,N_8714);
xor U8812 (N_8812,N_8693,N_8723);
nor U8813 (N_8813,N_8622,N_8715);
nor U8814 (N_8814,N_8737,N_8653);
or U8815 (N_8815,N_8695,N_8751);
nand U8816 (N_8816,N_8654,N_8767);
nand U8817 (N_8817,N_8728,N_8652);
xor U8818 (N_8818,N_8774,N_8713);
nor U8819 (N_8819,N_8756,N_8718);
nand U8820 (N_8820,N_8657,N_8764);
xnor U8821 (N_8821,N_8606,N_8700);
xnor U8822 (N_8822,N_8698,N_8799);
or U8823 (N_8823,N_8721,N_8732);
or U8824 (N_8824,N_8675,N_8619);
and U8825 (N_8825,N_8690,N_8752);
or U8826 (N_8826,N_8703,N_8642);
nor U8827 (N_8827,N_8682,N_8625);
or U8828 (N_8828,N_8745,N_8674);
and U8829 (N_8829,N_8631,N_8646);
nand U8830 (N_8830,N_8649,N_8685);
and U8831 (N_8831,N_8609,N_8670);
nand U8832 (N_8832,N_8716,N_8776);
nor U8833 (N_8833,N_8684,N_8750);
and U8834 (N_8834,N_8779,N_8726);
nor U8835 (N_8835,N_8644,N_8664);
xnor U8836 (N_8836,N_8770,N_8641);
and U8837 (N_8837,N_8738,N_8613);
nand U8838 (N_8838,N_8757,N_8747);
and U8839 (N_8839,N_8697,N_8640);
or U8840 (N_8840,N_8730,N_8782);
xor U8841 (N_8841,N_8771,N_8731);
nand U8842 (N_8842,N_8783,N_8681);
and U8843 (N_8843,N_8761,N_8741);
and U8844 (N_8844,N_8796,N_8701);
nor U8845 (N_8845,N_8614,N_8706);
nand U8846 (N_8846,N_8733,N_8632);
or U8847 (N_8847,N_8659,N_8621);
nand U8848 (N_8848,N_8602,N_8762);
xnor U8849 (N_8849,N_8763,N_8601);
nand U8850 (N_8850,N_8709,N_8671);
nand U8851 (N_8851,N_8648,N_8626);
nand U8852 (N_8852,N_8749,N_8620);
nand U8853 (N_8853,N_8666,N_8734);
nand U8854 (N_8854,N_8708,N_8689);
and U8855 (N_8855,N_8769,N_8742);
nand U8856 (N_8856,N_8760,N_8635);
xnor U8857 (N_8857,N_8777,N_8636);
nand U8858 (N_8858,N_8766,N_8608);
or U8859 (N_8859,N_8679,N_8667);
nand U8860 (N_8860,N_8637,N_8662);
xor U8861 (N_8861,N_8789,N_8661);
nor U8862 (N_8862,N_8699,N_8628);
nand U8863 (N_8863,N_8712,N_8694);
nor U8864 (N_8864,N_8651,N_8618);
nand U8865 (N_8865,N_8656,N_8692);
or U8866 (N_8866,N_8686,N_8753);
nand U8867 (N_8867,N_8629,N_8740);
nor U8868 (N_8868,N_8663,N_8658);
nor U8869 (N_8869,N_8758,N_8735);
nand U8870 (N_8870,N_8650,N_8722);
and U8871 (N_8871,N_8787,N_8788);
nor U8872 (N_8872,N_8603,N_8673);
and U8873 (N_8873,N_8743,N_8611);
or U8874 (N_8874,N_8744,N_8798);
nand U8875 (N_8875,N_8785,N_8739);
nor U8876 (N_8876,N_8775,N_8792);
nor U8877 (N_8877,N_8717,N_8665);
nand U8878 (N_8878,N_8616,N_8725);
xnor U8879 (N_8879,N_8794,N_8702);
and U8880 (N_8880,N_8729,N_8765);
and U8881 (N_8881,N_8772,N_8627);
xor U8882 (N_8882,N_8680,N_8720);
or U8883 (N_8883,N_8617,N_8605);
xor U8884 (N_8884,N_8615,N_8638);
nor U8885 (N_8885,N_8683,N_8791);
nor U8886 (N_8886,N_8607,N_8707);
or U8887 (N_8887,N_8755,N_8711);
nor U8888 (N_8888,N_8623,N_8748);
nor U8889 (N_8889,N_8780,N_8610);
nand U8890 (N_8890,N_8612,N_8660);
nand U8891 (N_8891,N_8773,N_8746);
and U8892 (N_8892,N_8643,N_8696);
nor U8893 (N_8893,N_8647,N_8676);
nor U8894 (N_8894,N_8793,N_8691);
or U8895 (N_8895,N_8768,N_8633);
nand U8896 (N_8896,N_8655,N_8630);
and U8897 (N_8897,N_8600,N_8778);
or U8898 (N_8898,N_8669,N_8687);
nand U8899 (N_8899,N_8677,N_8795);
xor U8900 (N_8900,N_8652,N_8706);
xor U8901 (N_8901,N_8680,N_8609);
and U8902 (N_8902,N_8684,N_8791);
nor U8903 (N_8903,N_8762,N_8679);
and U8904 (N_8904,N_8745,N_8677);
and U8905 (N_8905,N_8614,N_8696);
or U8906 (N_8906,N_8793,N_8634);
or U8907 (N_8907,N_8757,N_8763);
nand U8908 (N_8908,N_8627,N_8712);
nand U8909 (N_8909,N_8631,N_8687);
xor U8910 (N_8910,N_8679,N_8720);
nor U8911 (N_8911,N_8685,N_8607);
or U8912 (N_8912,N_8613,N_8685);
or U8913 (N_8913,N_8678,N_8686);
nand U8914 (N_8914,N_8792,N_8620);
nor U8915 (N_8915,N_8626,N_8664);
nand U8916 (N_8916,N_8779,N_8794);
nor U8917 (N_8917,N_8769,N_8687);
nand U8918 (N_8918,N_8783,N_8735);
xor U8919 (N_8919,N_8736,N_8745);
nand U8920 (N_8920,N_8703,N_8611);
or U8921 (N_8921,N_8753,N_8614);
and U8922 (N_8922,N_8795,N_8614);
xnor U8923 (N_8923,N_8774,N_8683);
or U8924 (N_8924,N_8728,N_8751);
nand U8925 (N_8925,N_8769,N_8696);
or U8926 (N_8926,N_8614,N_8762);
nand U8927 (N_8927,N_8673,N_8605);
nor U8928 (N_8928,N_8688,N_8662);
xor U8929 (N_8929,N_8668,N_8701);
and U8930 (N_8930,N_8730,N_8733);
nand U8931 (N_8931,N_8782,N_8707);
nor U8932 (N_8932,N_8671,N_8766);
or U8933 (N_8933,N_8694,N_8613);
xnor U8934 (N_8934,N_8780,N_8723);
nor U8935 (N_8935,N_8703,N_8767);
nand U8936 (N_8936,N_8685,N_8614);
xor U8937 (N_8937,N_8655,N_8644);
xnor U8938 (N_8938,N_8654,N_8780);
nand U8939 (N_8939,N_8657,N_8726);
nor U8940 (N_8940,N_8609,N_8656);
xnor U8941 (N_8941,N_8780,N_8686);
and U8942 (N_8942,N_8700,N_8658);
nor U8943 (N_8943,N_8765,N_8633);
nor U8944 (N_8944,N_8698,N_8629);
or U8945 (N_8945,N_8783,N_8747);
and U8946 (N_8946,N_8743,N_8634);
and U8947 (N_8947,N_8702,N_8714);
and U8948 (N_8948,N_8708,N_8692);
nor U8949 (N_8949,N_8668,N_8615);
nand U8950 (N_8950,N_8763,N_8625);
nand U8951 (N_8951,N_8701,N_8751);
xnor U8952 (N_8952,N_8668,N_8754);
and U8953 (N_8953,N_8736,N_8775);
and U8954 (N_8954,N_8635,N_8741);
nand U8955 (N_8955,N_8741,N_8720);
nand U8956 (N_8956,N_8650,N_8742);
or U8957 (N_8957,N_8606,N_8719);
xor U8958 (N_8958,N_8665,N_8690);
nor U8959 (N_8959,N_8666,N_8718);
nor U8960 (N_8960,N_8796,N_8629);
and U8961 (N_8961,N_8707,N_8787);
nor U8962 (N_8962,N_8718,N_8699);
and U8963 (N_8963,N_8743,N_8647);
nor U8964 (N_8964,N_8787,N_8694);
xnor U8965 (N_8965,N_8613,N_8661);
nand U8966 (N_8966,N_8632,N_8741);
and U8967 (N_8967,N_8781,N_8700);
xnor U8968 (N_8968,N_8656,N_8705);
or U8969 (N_8969,N_8745,N_8670);
xor U8970 (N_8970,N_8651,N_8707);
nor U8971 (N_8971,N_8746,N_8642);
and U8972 (N_8972,N_8613,N_8710);
and U8973 (N_8973,N_8739,N_8615);
and U8974 (N_8974,N_8691,N_8665);
and U8975 (N_8975,N_8601,N_8622);
nand U8976 (N_8976,N_8787,N_8613);
xnor U8977 (N_8977,N_8705,N_8691);
nor U8978 (N_8978,N_8712,N_8721);
or U8979 (N_8979,N_8758,N_8621);
and U8980 (N_8980,N_8600,N_8722);
nand U8981 (N_8981,N_8615,N_8752);
or U8982 (N_8982,N_8791,N_8609);
xor U8983 (N_8983,N_8678,N_8717);
xor U8984 (N_8984,N_8642,N_8707);
and U8985 (N_8985,N_8612,N_8626);
and U8986 (N_8986,N_8768,N_8720);
xor U8987 (N_8987,N_8749,N_8751);
nand U8988 (N_8988,N_8759,N_8681);
nand U8989 (N_8989,N_8627,N_8707);
nand U8990 (N_8990,N_8675,N_8640);
or U8991 (N_8991,N_8794,N_8678);
xor U8992 (N_8992,N_8734,N_8643);
or U8993 (N_8993,N_8624,N_8651);
or U8994 (N_8994,N_8646,N_8789);
xnor U8995 (N_8995,N_8723,N_8765);
nand U8996 (N_8996,N_8785,N_8684);
nor U8997 (N_8997,N_8769,N_8751);
and U8998 (N_8998,N_8603,N_8672);
or U8999 (N_8999,N_8668,N_8650);
nor U9000 (N_9000,N_8983,N_8823);
nor U9001 (N_9001,N_8998,N_8945);
and U9002 (N_9002,N_8942,N_8965);
and U9003 (N_9003,N_8948,N_8999);
or U9004 (N_9004,N_8938,N_8988);
or U9005 (N_9005,N_8874,N_8892);
nand U9006 (N_9006,N_8963,N_8830);
or U9007 (N_9007,N_8868,N_8814);
xor U9008 (N_9008,N_8884,N_8863);
and U9009 (N_9009,N_8832,N_8978);
nor U9010 (N_9010,N_8807,N_8995);
xor U9011 (N_9011,N_8964,N_8934);
and U9012 (N_9012,N_8960,N_8816);
or U9013 (N_9013,N_8844,N_8831);
and U9014 (N_9014,N_8900,N_8947);
and U9015 (N_9015,N_8801,N_8993);
nand U9016 (N_9016,N_8961,N_8917);
nor U9017 (N_9017,N_8904,N_8856);
or U9018 (N_9018,N_8977,N_8802);
nor U9019 (N_9019,N_8951,N_8922);
or U9020 (N_9020,N_8838,N_8962);
nand U9021 (N_9021,N_8957,N_8845);
and U9022 (N_9022,N_8970,N_8937);
and U9023 (N_9023,N_8818,N_8866);
nor U9024 (N_9024,N_8901,N_8815);
nand U9025 (N_9025,N_8940,N_8827);
xnor U9026 (N_9026,N_8865,N_8852);
xnor U9027 (N_9027,N_8805,N_8822);
or U9028 (N_9028,N_8878,N_8898);
nand U9029 (N_9029,N_8862,N_8897);
and U9030 (N_9030,N_8902,N_8986);
or U9031 (N_9031,N_8987,N_8910);
or U9032 (N_9032,N_8877,N_8976);
xnor U9033 (N_9033,N_8846,N_8925);
or U9034 (N_9034,N_8981,N_8953);
xor U9035 (N_9035,N_8973,N_8817);
nand U9036 (N_9036,N_8843,N_8850);
nand U9037 (N_9037,N_8880,N_8989);
xor U9038 (N_9038,N_8890,N_8848);
and U9039 (N_9039,N_8895,N_8980);
and U9040 (N_9040,N_8870,N_8875);
or U9041 (N_9041,N_8930,N_8984);
xor U9042 (N_9042,N_8835,N_8847);
nand U9043 (N_9043,N_8819,N_8915);
xnor U9044 (N_9044,N_8853,N_8908);
nor U9045 (N_9045,N_8968,N_8979);
and U9046 (N_9046,N_8867,N_8903);
or U9047 (N_9047,N_8972,N_8885);
nor U9048 (N_9048,N_8812,N_8956);
xnor U9049 (N_9049,N_8941,N_8924);
nand U9050 (N_9050,N_8985,N_8912);
or U9051 (N_9051,N_8946,N_8820);
or U9052 (N_9052,N_8899,N_8821);
xnor U9053 (N_9053,N_8907,N_8836);
and U9054 (N_9054,N_8834,N_8881);
nor U9055 (N_9055,N_8905,N_8969);
or U9056 (N_9056,N_8859,N_8994);
xnor U9057 (N_9057,N_8891,N_8921);
and U9058 (N_9058,N_8810,N_8966);
xnor U9059 (N_9059,N_8855,N_8813);
xnor U9060 (N_9060,N_8840,N_8894);
xor U9061 (N_9061,N_8851,N_8974);
and U9062 (N_9062,N_8919,N_8933);
xor U9063 (N_9063,N_8990,N_8871);
or U9064 (N_9064,N_8911,N_8952);
xor U9065 (N_9065,N_8876,N_8918);
or U9066 (N_9066,N_8869,N_8839);
and U9067 (N_9067,N_8975,N_8837);
xnor U9068 (N_9068,N_8829,N_8873);
xor U9069 (N_9069,N_8828,N_8809);
nand U9070 (N_9070,N_8992,N_8889);
and U9071 (N_9071,N_8887,N_8936);
nor U9072 (N_9072,N_8926,N_8800);
and U9073 (N_9073,N_8854,N_8950);
nand U9074 (N_9074,N_8991,N_8833);
nor U9075 (N_9075,N_8872,N_8888);
nor U9076 (N_9076,N_8971,N_8996);
xnor U9077 (N_9077,N_8932,N_8997);
nand U9078 (N_9078,N_8929,N_8955);
and U9079 (N_9079,N_8913,N_8944);
nor U9080 (N_9080,N_8883,N_8982);
xnor U9081 (N_9081,N_8882,N_8824);
nand U9082 (N_9082,N_8808,N_8861);
xor U9083 (N_9083,N_8927,N_8958);
xnor U9084 (N_9084,N_8860,N_8920);
nand U9085 (N_9085,N_8914,N_8949);
xor U9086 (N_9086,N_8825,N_8826);
xnor U9087 (N_9087,N_8909,N_8849);
and U9088 (N_9088,N_8806,N_8906);
and U9089 (N_9089,N_8939,N_8923);
xnor U9090 (N_9090,N_8886,N_8841);
and U9091 (N_9091,N_8857,N_8954);
xnor U9092 (N_9092,N_8879,N_8864);
nor U9093 (N_9093,N_8916,N_8811);
xor U9094 (N_9094,N_8931,N_8842);
nand U9095 (N_9095,N_8967,N_8928);
xor U9096 (N_9096,N_8858,N_8896);
or U9097 (N_9097,N_8893,N_8935);
nor U9098 (N_9098,N_8943,N_8803);
or U9099 (N_9099,N_8959,N_8804);
xnor U9100 (N_9100,N_8914,N_8827);
xnor U9101 (N_9101,N_8972,N_8985);
nor U9102 (N_9102,N_8859,N_8912);
xor U9103 (N_9103,N_8879,N_8811);
and U9104 (N_9104,N_8994,N_8844);
xnor U9105 (N_9105,N_8841,N_8827);
and U9106 (N_9106,N_8824,N_8821);
and U9107 (N_9107,N_8961,N_8971);
and U9108 (N_9108,N_8933,N_8973);
nor U9109 (N_9109,N_8834,N_8869);
or U9110 (N_9110,N_8941,N_8923);
nor U9111 (N_9111,N_8992,N_8913);
nand U9112 (N_9112,N_8944,N_8815);
nand U9113 (N_9113,N_8840,N_8814);
or U9114 (N_9114,N_8802,N_8908);
and U9115 (N_9115,N_8901,N_8909);
or U9116 (N_9116,N_8934,N_8955);
xor U9117 (N_9117,N_8803,N_8805);
nand U9118 (N_9118,N_8885,N_8935);
nor U9119 (N_9119,N_8836,N_8843);
nor U9120 (N_9120,N_8965,N_8901);
or U9121 (N_9121,N_8806,N_8810);
or U9122 (N_9122,N_8928,N_8815);
and U9123 (N_9123,N_8823,N_8878);
nor U9124 (N_9124,N_8926,N_8839);
or U9125 (N_9125,N_8944,N_8905);
and U9126 (N_9126,N_8993,N_8874);
xnor U9127 (N_9127,N_8974,N_8961);
nand U9128 (N_9128,N_8935,N_8924);
nand U9129 (N_9129,N_8927,N_8805);
or U9130 (N_9130,N_8881,N_8904);
and U9131 (N_9131,N_8935,N_8932);
or U9132 (N_9132,N_8843,N_8873);
nand U9133 (N_9133,N_8907,N_8990);
or U9134 (N_9134,N_8908,N_8928);
and U9135 (N_9135,N_8943,N_8976);
or U9136 (N_9136,N_8946,N_8998);
or U9137 (N_9137,N_8960,N_8963);
xor U9138 (N_9138,N_8917,N_8904);
and U9139 (N_9139,N_8911,N_8813);
and U9140 (N_9140,N_8947,N_8906);
or U9141 (N_9141,N_8933,N_8921);
nand U9142 (N_9142,N_8930,N_8843);
or U9143 (N_9143,N_8848,N_8858);
nand U9144 (N_9144,N_8969,N_8801);
nor U9145 (N_9145,N_8980,N_8839);
nor U9146 (N_9146,N_8958,N_8888);
nand U9147 (N_9147,N_8896,N_8861);
and U9148 (N_9148,N_8950,N_8839);
and U9149 (N_9149,N_8988,N_8949);
nor U9150 (N_9150,N_8878,N_8801);
or U9151 (N_9151,N_8833,N_8841);
or U9152 (N_9152,N_8952,N_8977);
or U9153 (N_9153,N_8952,N_8981);
nor U9154 (N_9154,N_8943,N_8914);
nand U9155 (N_9155,N_8961,N_8899);
and U9156 (N_9156,N_8835,N_8927);
nor U9157 (N_9157,N_8863,N_8810);
xor U9158 (N_9158,N_8913,N_8815);
nor U9159 (N_9159,N_8979,N_8995);
xnor U9160 (N_9160,N_8939,N_8958);
or U9161 (N_9161,N_8851,N_8981);
nor U9162 (N_9162,N_8955,N_8809);
xnor U9163 (N_9163,N_8886,N_8898);
nand U9164 (N_9164,N_8870,N_8975);
nor U9165 (N_9165,N_8895,N_8811);
nor U9166 (N_9166,N_8951,N_8924);
and U9167 (N_9167,N_8935,N_8981);
xor U9168 (N_9168,N_8998,N_8865);
nand U9169 (N_9169,N_8993,N_8834);
or U9170 (N_9170,N_8912,N_8956);
nand U9171 (N_9171,N_8818,N_8837);
and U9172 (N_9172,N_8916,N_8951);
nand U9173 (N_9173,N_8877,N_8999);
or U9174 (N_9174,N_8999,N_8814);
or U9175 (N_9175,N_8800,N_8867);
or U9176 (N_9176,N_8938,N_8867);
nor U9177 (N_9177,N_8963,N_8923);
xor U9178 (N_9178,N_8842,N_8858);
nor U9179 (N_9179,N_8966,N_8902);
nand U9180 (N_9180,N_8940,N_8891);
or U9181 (N_9181,N_8837,N_8834);
nand U9182 (N_9182,N_8956,N_8911);
and U9183 (N_9183,N_8999,N_8934);
nor U9184 (N_9184,N_8943,N_8991);
nor U9185 (N_9185,N_8935,N_8864);
or U9186 (N_9186,N_8839,N_8892);
xor U9187 (N_9187,N_8957,N_8888);
nor U9188 (N_9188,N_8916,N_8961);
xnor U9189 (N_9189,N_8814,N_8844);
nor U9190 (N_9190,N_8825,N_8864);
xnor U9191 (N_9191,N_8936,N_8958);
xor U9192 (N_9192,N_8888,N_8823);
and U9193 (N_9193,N_8822,N_8863);
and U9194 (N_9194,N_8922,N_8811);
or U9195 (N_9195,N_8951,N_8848);
or U9196 (N_9196,N_8922,N_8895);
xor U9197 (N_9197,N_8942,N_8841);
xor U9198 (N_9198,N_8960,N_8921);
nand U9199 (N_9199,N_8898,N_8811);
xnor U9200 (N_9200,N_9118,N_9126);
xnor U9201 (N_9201,N_9189,N_9062);
or U9202 (N_9202,N_9150,N_9022);
or U9203 (N_9203,N_9009,N_9198);
or U9204 (N_9204,N_9072,N_9168);
xor U9205 (N_9205,N_9157,N_9160);
nand U9206 (N_9206,N_9130,N_9097);
nand U9207 (N_9207,N_9050,N_9010);
nand U9208 (N_9208,N_9034,N_9045);
nor U9209 (N_9209,N_9170,N_9023);
or U9210 (N_9210,N_9177,N_9102);
nand U9211 (N_9211,N_9103,N_9004);
nor U9212 (N_9212,N_9100,N_9012);
nor U9213 (N_9213,N_9031,N_9145);
nor U9214 (N_9214,N_9019,N_9172);
and U9215 (N_9215,N_9188,N_9075);
nor U9216 (N_9216,N_9042,N_9140);
nand U9217 (N_9217,N_9104,N_9033);
xor U9218 (N_9218,N_9090,N_9053);
nor U9219 (N_9219,N_9190,N_9005);
xor U9220 (N_9220,N_9088,N_9067);
or U9221 (N_9221,N_9182,N_9143);
xor U9222 (N_9222,N_9032,N_9017);
nor U9223 (N_9223,N_9154,N_9052);
nand U9224 (N_9224,N_9132,N_9038);
nor U9225 (N_9225,N_9011,N_9197);
nand U9226 (N_9226,N_9056,N_9024);
and U9227 (N_9227,N_9186,N_9110);
nor U9228 (N_9228,N_9128,N_9036);
nor U9229 (N_9229,N_9046,N_9181);
and U9230 (N_9230,N_9159,N_9028);
and U9231 (N_9231,N_9183,N_9078);
or U9232 (N_9232,N_9002,N_9113);
nor U9233 (N_9233,N_9179,N_9063);
nor U9234 (N_9234,N_9109,N_9173);
nor U9235 (N_9235,N_9124,N_9119);
nand U9236 (N_9236,N_9171,N_9095);
nor U9237 (N_9237,N_9014,N_9057);
xor U9238 (N_9238,N_9089,N_9055);
or U9239 (N_9239,N_9027,N_9060);
and U9240 (N_9240,N_9049,N_9066);
or U9241 (N_9241,N_9117,N_9142);
nand U9242 (N_9242,N_9007,N_9194);
or U9243 (N_9243,N_9184,N_9098);
nor U9244 (N_9244,N_9144,N_9175);
nor U9245 (N_9245,N_9065,N_9092);
xnor U9246 (N_9246,N_9006,N_9137);
nand U9247 (N_9247,N_9085,N_9116);
or U9248 (N_9248,N_9185,N_9153);
nor U9249 (N_9249,N_9058,N_9073);
nor U9250 (N_9250,N_9176,N_9018);
xor U9251 (N_9251,N_9149,N_9030);
or U9252 (N_9252,N_9165,N_9122);
nand U9253 (N_9253,N_9029,N_9141);
nand U9254 (N_9254,N_9147,N_9008);
xor U9255 (N_9255,N_9167,N_9035);
nor U9256 (N_9256,N_9079,N_9081);
nor U9257 (N_9257,N_9086,N_9163);
and U9258 (N_9258,N_9155,N_9051);
and U9259 (N_9259,N_9077,N_9048);
xor U9260 (N_9260,N_9164,N_9064);
nor U9261 (N_9261,N_9121,N_9084);
nand U9262 (N_9262,N_9087,N_9020);
and U9263 (N_9263,N_9151,N_9080);
nor U9264 (N_9264,N_9129,N_9013);
nand U9265 (N_9265,N_9196,N_9021);
xor U9266 (N_9266,N_9091,N_9039);
xor U9267 (N_9267,N_9061,N_9133);
xor U9268 (N_9268,N_9193,N_9037);
nand U9269 (N_9269,N_9094,N_9125);
nand U9270 (N_9270,N_9059,N_9069);
xor U9271 (N_9271,N_9112,N_9099);
nand U9272 (N_9272,N_9044,N_9187);
and U9273 (N_9273,N_9015,N_9076);
nor U9274 (N_9274,N_9123,N_9040);
nor U9275 (N_9275,N_9192,N_9000);
nor U9276 (N_9276,N_9162,N_9139);
and U9277 (N_9277,N_9026,N_9180);
nand U9278 (N_9278,N_9107,N_9174);
or U9279 (N_9279,N_9070,N_9152);
nor U9280 (N_9280,N_9131,N_9111);
nand U9281 (N_9281,N_9146,N_9001);
and U9282 (N_9282,N_9135,N_9161);
and U9283 (N_9283,N_9136,N_9071);
nor U9284 (N_9284,N_9169,N_9105);
nand U9285 (N_9285,N_9083,N_9195);
nor U9286 (N_9286,N_9016,N_9047);
and U9287 (N_9287,N_9158,N_9082);
xor U9288 (N_9288,N_9120,N_9191);
nor U9289 (N_9289,N_9096,N_9041);
nand U9290 (N_9290,N_9114,N_9127);
xnor U9291 (N_9291,N_9003,N_9043);
nand U9292 (N_9292,N_9054,N_9068);
nand U9293 (N_9293,N_9025,N_9156);
or U9294 (N_9294,N_9148,N_9138);
xnor U9295 (N_9295,N_9199,N_9134);
nor U9296 (N_9296,N_9106,N_9074);
or U9297 (N_9297,N_9115,N_9166);
xnor U9298 (N_9298,N_9093,N_9108);
xor U9299 (N_9299,N_9178,N_9101);
nor U9300 (N_9300,N_9145,N_9090);
or U9301 (N_9301,N_9041,N_9164);
or U9302 (N_9302,N_9141,N_9025);
nor U9303 (N_9303,N_9116,N_9181);
nand U9304 (N_9304,N_9181,N_9144);
and U9305 (N_9305,N_9091,N_9016);
or U9306 (N_9306,N_9161,N_9058);
or U9307 (N_9307,N_9011,N_9191);
xor U9308 (N_9308,N_9192,N_9174);
and U9309 (N_9309,N_9192,N_9069);
xnor U9310 (N_9310,N_9118,N_9119);
xnor U9311 (N_9311,N_9053,N_9051);
and U9312 (N_9312,N_9025,N_9042);
xnor U9313 (N_9313,N_9161,N_9173);
or U9314 (N_9314,N_9181,N_9077);
and U9315 (N_9315,N_9189,N_9122);
or U9316 (N_9316,N_9190,N_9164);
nor U9317 (N_9317,N_9142,N_9189);
and U9318 (N_9318,N_9024,N_9191);
nand U9319 (N_9319,N_9078,N_9039);
nand U9320 (N_9320,N_9101,N_9050);
or U9321 (N_9321,N_9013,N_9003);
xor U9322 (N_9322,N_9035,N_9029);
nor U9323 (N_9323,N_9170,N_9019);
or U9324 (N_9324,N_9178,N_9142);
or U9325 (N_9325,N_9099,N_9121);
or U9326 (N_9326,N_9183,N_9011);
nor U9327 (N_9327,N_9194,N_9130);
and U9328 (N_9328,N_9134,N_9138);
nor U9329 (N_9329,N_9121,N_9168);
or U9330 (N_9330,N_9153,N_9163);
nand U9331 (N_9331,N_9110,N_9043);
or U9332 (N_9332,N_9150,N_9009);
nor U9333 (N_9333,N_9005,N_9086);
nor U9334 (N_9334,N_9107,N_9008);
xnor U9335 (N_9335,N_9105,N_9184);
nor U9336 (N_9336,N_9152,N_9082);
nor U9337 (N_9337,N_9122,N_9143);
and U9338 (N_9338,N_9096,N_9130);
nand U9339 (N_9339,N_9162,N_9100);
nor U9340 (N_9340,N_9032,N_9026);
or U9341 (N_9341,N_9179,N_9067);
nor U9342 (N_9342,N_9188,N_9143);
or U9343 (N_9343,N_9114,N_9064);
or U9344 (N_9344,N_9042,N_9067);
nor U9345 (N_9345,N_9119,N_9093);
nand U9346 (N_9346,N_9175,N_9148);
nand U9347 (N_9347,N_9185,N_9158);
and U9348 (N_9348,N_9114,N_9123);
or U9349 (N_9349,N_9108,N_9182);
nand U9350 (N_9350,N_9101,N_9176);
and U9351 (N_9351,N_9037,N_9162);
or U9352 (N_9352,N_9074,N_9066);
nor U9353 (N_9353,N_9137,N_9155);
or U9354 (N_9354,N_9116,N_9013);
and U9355 (N_9355,N_9085,N_9177);
and U9356 (N_9356,N_9180,N_9198);
xor U9357 (N_9357,N_9041,N_9098);
nand U9358 (N_9358,N_9106,N_9048);
nor U9359 (N_9359,N_9007,N_9142);
and U9360 (N_9360,N_9145,N_9003);
xnor U9361 (N_9361,N_9003,N_9072);
or U9362 (N_9362,N_9024,N_9176);
xor U9363 (N_9363,N_9000,N_9004);
or U9364 (N_9364,N_9069,N_9102);
or U9365 (N_9365,N_9103,N_9061);
nor U9366 (N_9366,N_9031,N_9158);
nor U9367 (N_9367,N_9151,N_9167);
and U9368 (N_9368,N_9084,N_9117);
xnor U9369 (N_9369,N_9044,N_9135);
nand U9370 (N_9370,N_9051,N_9149);
or U9371 (N_9371,N_9083,N_9009);
or U9372 (N_9372,N_9030,N_9109);
nand U9373 (N_9373,N_9034,N_9078);
nand U9374 (N_9374,N_9057,N_9112);
and U9375 (N_9375,N_9050,N_9168);
xnor U9376 (N_9376,N_9084,N_9055);
or U9377 (N_9377,N_9011,N_9040);
nor U9378 (N_9378,N_9117,N_9072);
nand U9379 (N_9379,N_9122,N_9183);
xor U9380 (N_9380,N_9110,N_9166);
or U9381 (N_9381,N_9106,N_9139);
or U9382 (N_9382,N_9059,N_9107);
or U9383 (N_9383,N_9053,N_9140);
xnor U9384 (N_9384,N_9068,N_9180);
nand U9385 (N_9385,N_9084,N_9164);
nand U9386 (N_9386,N_9038,N_9076);
and U9387 (N_9387,N_9161,N_9014);
nor U9388 (N_9388,N_9067,N_9175);
or U9389 (N_9389,N_9189,N_9181);
nor U9390 (N_9390,N_9060,N_9172);
or U9391 (N_9391,N_9009,N_9101);
or U9392 (N_9392,N_9194,N_9121);
or U9393 (N_9393,N_9187,N_9021);
xor U9394 (N_9394,N_9108,N_9195);
and U9395 (N_9395,N_9016,N_9188);
nor U9396 (N_9396,N_9187,N_9033);
xnor U9397 (N_9397,N_9167,N_9057);
nor U9398 (N_9398,N_9050,N_9130);
and U9399 (N_9399,N_9076,N_9089);
xor U9400 (N_9400,N_9213,N_9371);
and U9401 (N_9401,N_9307,N_9362);
nand U9402 (N_9402,N_9322,N_9393);
or U9403 (N_9403,N_9334,N_9205);
nand U9404 (N_9404,N_9330,N_9230);
and U9405 (N_9405,N_9285,N_9333);
xnor U9406 (N_9406,N_9346,N_9383);
nor U9407 (N_9407,N_9313,N_9389);
and U9408 (N_9408,N_9271,N_9254);
and U9409 (N_9409,N_9275,N_9258);
xnor U9410 (N_9410,N_9369,N_9326);
and U9411 (N_9411,N_9263,N_9231);
nand U9412 (N_9412,N_9324,N_9204);
or U9413 (N_9413,N_9245,N_9370);
or U9414 (N_9414,N_9239,N_9358);
or U9415 (N_9415,N_9292,N_9257);
xnor U9416 (N_9416,N_9299,N_9396);
nor U9417 (N_9417,N_9363,N_9380);
nor U9418 (N_9418,N_9265,N_9207);
xnor U9419 (N_9419,N_9349,N_9291);
nand U9420 (N_9420,N_9268,N_9248);
nand U9421 (N_9421,N_9323,N_9378);
and U9422 (N_9422,N_9367,N_9214);
or U9423 (N_9423,N_9351,N_9392);
and U9424 (N_9424,N_9296,N_9356);
nor U9425 (N_9425,N_9339,N_9319);
and U9426 (N_9426,N_9293,N_9355);
nand U9427 (N_9427,N_9256,N_9385);
xnor U9428 (N_9428,N_9211,N_9353);
and U9429 (N_9429,N_9295,N_9286);
and U9430 (N_9430,N_9365,N_9298);
or U9431 (N_9431,N_9282,N_9327);
nor U9432 (N_9432,N_9233,N_9395);
nor U9433 (N_9433,N_9225,N_9316);
nor U9434 (N_9434,N_9372,N_9242);
xor U9435 (N_9435,N_9294,N_9218);
nor U9436 (N_9436,N_9272,N_9228);
nor U9437 (N_9437,N_9202,N_9397);
nand U9438 (N_9438,N_9244,N_9366);
xor U9439 (N_9439,N_9344,N_9284);
and U9440 (N_9440,N_9359,N_9252);
or U9441 (N_9441,N_9338,N_9206);
and U9442 (N_9442,N_9278,N_9347);
xor U9443 (N_9443,N_9360,N_9317);
xor U9444 (N_9444,N_9399,N_9279);
and U9445 (N_9445,N_9384,N_9388);
and U9446 (N_9446,N_9283,N_9276);
or U9447 (N_9447,N_9246,N_9303);
and U9448 (N_9448,N_9251,N_9304);
or U9449 (N_9449,N_9273,N_9302);
xor U9450 (N_9450,N_9341,N_9229);
xor U9451 (N_9451,N_9234,N_9364);
nand U9452 (N_9452,N_9373,N_9223);
nor U9453 (N_9453,N_9390,N_9361);
and U9454 (N_9454,N_9217,N_9289);
xnor U9455 (N_9455,N_9287,N_9345);
nor U9456 (N_9456,N_9325,N_9320);
nand U9457 (N_9457,N_9309,N_9288);
or U9458 (N_9458,N_9377,N_9249);
xor U9459 (N_9459,N_9310,N_9306);
or U9460 (N_9460,N_9329,N_9210);
nand U9461 (N_9461,N_9232,N_9352);
and U9462 (N_9462,N_9235,N_9253);
and U9463 (N_9463,N_9220,N_9255);
nor U9464 (N_9464,N_9348,N_9308);
xnor U9465 (N_9465,N_9336,N_9375);
nor U9466 (N_9466,N_9227,N_9398);
xnor U9467 (N_9467,N_9266,N_9269);
nor U9468 (N_9468,N_9222,N_9312);
nand U9469 (N_9469,N_9328,N_9315);
xnor U9470 (N_9470,N_9237,N_9274);
and U9471 (N_9471,N_9219,N_9240);
nand U9472 (N_9472,N_9374,N_9224);
and U9473 (N_9473,N_9368,N_9337);
nand U9474 (N_9474,N_9267,N_9270);
nor U9475 (N_9475,N_9290,N_9354);
and U9476 (N_9476,N_9297,N_9201);
nor U9477 (N_9477,N_9277,N_9357);
or U9478 (N_9478,N_9305,N_9376);
xnor U9479 (N_9479,N_9200,N_9216);
xor U9480 (N_9480,N_9318,N_9387);
xnor U9481 (N_9481,N_9281,N_9241);
nor U9482 (N_9482,N_9247,N_9238);
nand U9483 (N_9483,N_9311,N_9236);
xor U9484 (N_9484,N_9226,N_9335);
or U9485 (N_9485,N_9203,N_9379);
and U9486 (N_9486,N_9314,N_9332);
nand U9487 (N_9487,N_9212,N_9208);
nor U9488 (N_9488,N_9386,N_9261);
nand U9489 (N_9489,N_9340,N_9382);
or U9490 (N_9490,N_9243,N_9259);
nor U9491 (N_9491,N_9342,N_9350);
and U9492 (N_9492,N_9264,N_9262);
nand U9493 (N_9493,N_9381,N_9331);
or U9494 (N_9494,N_9221,N_9394);
xor U9495 (N_9495,N_9321,N_9260);
and U9496 (N_9496,N_9215,N_9391);
xor U9497 (N_9497,N_9280,N_9209);
and U9498 (N_9498,N_9250,N_9343);
nor U9499 (N_9499,N_9300,N_9301);
nand U9500 (N_9500,N_9300,N_9377);
or U9501 (N_9501,N_9274,N_9360);
nand U9502 (N_9502,N_9262,N_9273);
and U9503 (N_9503,N_9363,N_9278);
and U9504 (N_9504,N_9365,N_9354);
xor U9505 (N_9505,N_9281,N_9279);
or U9506 (N_9506,N_9285,N_9357);
nand U9507 (N_9507,N_9231,N_9248);
or U9508 (N_9508,N_9319,N_9352);
nand U9509 (N_9509,N_9372,N_9373);
and U9510 (N_9510,N_9301,N_9298);
or U9511 (N_9511,N_9260,N_9387);
xnor U9512 (N_9512,N_9301,N_9314);
nand U9513 (N_9513,N_9359,N_9206);
and U9514 (N_9514,N_9314,N_9224);
nand U9515 (N_9515,N_9259,N_9317);
nor U9516 (N_9516,N_9342,N_9284);
and U9517 (N_9517,N_9385,N_9392);
xor U9518 (N_9518,N_9246,N_9276);
and U9519 (N_9519,N_9279,N_9387);
nor U9520 (N_9520,N_9357,N_9291);
xnor U9521 (N_9521,N_9333,N_9291);
nand U9522 (N_9522,N_9297,N_9286);
nor U9523 (N_9523,N_9243,N_9348);
nor U9524 (N_9524,N_9211,N_9208);
nor U9525 (N_9525,N_9390,N_9343);
nand U9526 (N_9526,N_9261,N_9225);
and U9527 (N_9527,N_9271,N_9380);
and U9528 (N_9528,N_9269,N_9316);
and U9529 (N_9529,N_9279,N_9215);
xor U9530 (N_9530,N_9244,N_9368);
nor U9531 (N_9531,N_9399,N_9204);
nand U9532 (N_9532,N_9267,N_9204);
or U9533 (N_9533,N_9242,N_9214);
nor U9534 (N_9534,N_9276,N_9273);
nand U9535 (N_9535,N_9271,N_9277);
and U9536 (N_9536,N_9275,N_9371);
and U9537 (N_9537,N_9345,N_9309);
or U9538 (N_9538,N_9355,N_9217);
or U9539 (N_9539,N_9252,N_9275);
nand U9540 (N_9540,N_9223,N_9268);
nand U9541 (N_9541,N_9302,N_9248);
or U9542 (N_9542,N_9253,N_9277);
xor U9543 (N_9543,N_9291,N_9235);
xor U9544 (N_9544,N_9341,N_9280);
nand U9545 (N_9545,N_9294,N_9243);
nand U9546 (N_9546,N_9207,N_9311);
and U9547 (N_9547,N_9205,N_9265);
or U9548 (N_9548,N_9268,N_9257);
nand U9549 (N_9549,N_9251,N_9326);
nand U9550 (N_9550,N_9329,N_9235);
xor U9551 (N_9551,N_9293,N_9202);
nor U9552 (N_9552,N_9299,N_9227);
and U9553 (N_9553,N_9345,N_9377);
nand U9554 (N_9554,N_9387,N_9346);
xnor U9555 (N_9555,N_9256,N_9337);
nand U9556 (N_9556,N_9382,N_9287);
nor U9557 (N_9557,N_9318,N_9240);
or U9558 (N_9558,N_9361,N_9276);
or U9559 (N_9559,N_9395,N_9299);
nor U9560 (N_9560,N_9209,N_9204);
nand U9561 (N_9561,N_9305,N_9278);
xnor U9562 (N_9562,N_9201,N_9324);
and U9563 (N_9563,N_9362,N_9318);
xor U9564 (N_9564,N_9247,N_9269);
nor U9565 (N_9565,N_9232,N_9263);
or U9566 (N_9566,N_9306,N_9369);
xnor U9567 (N_9567,N_9385,N_9228);
nor U9568 (N_9568,N_9377,N_9309);
nor U9569 (N_9569,N_9223,N_9313);
xnor U9570 (N_9570,N_9313,N_9370);
and U9571 (N_9571,N_9286,N_9281);
or U9572 (N_9572,N_9313,N_9240);
nor U9573 (N_9573,N_9297,N_9234);
and U9574 (N_9574,N_9265,N_9377);
or U9575 (N_9575,N_9376,N_9245);
or U9576 (N_9576,N_9371,N_9362);
xor U9577 (N_9577,N_9302,N_9205);
nand U9578 (N_9578,N_9367,N_9270);
or U9579 (N_9579,N_9274,N_9376);
nor U9580 (N_9580,N_9251,N_9346);
or U9581 (N_9581,N_9321,N_9222);
nand U9582 (N_9582,N_9254,N_9253);
or U9583 (N_9583,N_9252,N_9351);
xor U9584 (N_9584,N_9224,N_9202);
nand U9585 (N_9585,N_9217,N_9287);
nor U9586 (N_9586,N_9343,N_9336);
and U9587 (N_9587,N_9334,N_9388);
and U9588 (N_9588,N_9298,N_9342);
and U9589 (N_9589,N_9282,N_9245);
nand U9590 (N_9590,N_9272,N_9220);
or U9591 (N_9591,N_9337,N_9371);
and U9592 (N_9592,N_9398,N_9381);
xor U9593 (N_9593,N_9365,N_9307);
and U9594 (N_9594,N_9221,N_9278);
nor U9595 (N_9595,N_9351,N_9218);
nor U9596 (N_9596,N_9360,N_9205);
and U9597 (N_9597,N_9208,N_9315);
xor U9598 (N_9598,N_9284,N_9231);
nor U9599 (N_9599,N_9226,N_9370);
or U9600 (N_9600,N_9489,N_9550);
nor U9601 (N_9601,N_9521,N_9533);
nand U9602 (N_9602,N_9574,N_9478);
or U9603 (N_9603,N_9530,N_9513);
and U9604 (N_9604,N_9416,N_9594);
or U9605 (N_9605,N_9420,N_9493);
nand U9606 (N_9606,N_9487,N_9418);
and U9607 (N_9607,N_9569,N_9488);
or U9608 (N_9608,N_9525,N_9409);
nand U9609 (N_9609,N_9503,N_9536);
or U9610 (N_9610,N_9452,N_9403);
xnor U9611 (N_9611,N_9494,N_9592);
or U9612 (N_9612,N_9560,N_9504);
nor U9613 (N_9613,N_9573,N_9532);
and U9614 (N_9614,N_9520,N_9438);
nor U9615 (N_9615,N_9408,N_9570);
nand U9616 (N_9616,N_9578,N_9432);
or U9617 (N_9617,N_9528,N_9486);
or U9618 (N_9618,N_9443,N_9511);
nand U9619 (N_9619,N_9501,N_9565);
xnor U9620 (N_9620,N_9453,N_9461);
or U9621 (N_9621,N_9559,N_9546);
nand U9622 (N_9622,N_9545,N_9411);
nand U9623 (N_9623,N_9467,N_9531);
or U9624 (N_9624,N_9466,N_9566);
nand U9625 (N_9625,N_9474,N_9549);
nor U9626 (N_9626,N_9457,N_9459);
nor U9627 (N_9627,N_9534,N_9468);
or U9628 (N_9628,N_9450,N_9480);
nor U9629 (N_9629,N_9458,N_9519);
xor U9630 (N_9630,N_9485,N_9540);
nor U9631 (N_9631,N_9442,N_9568);
or U9632 (N_9632,N_9479,N_9424);
nor U9633 (N_9633,N_9577,N_9596);
and U9634 (N_9634,N_9426,N_9506);
nor U9635 (N_9635,N_9422,N_9512);
xnor U9636 (N_9636,N_9481,N_9529);
or U9637 (N_9637,N_9567,N_9558);
or U9638 (N_9638,N_9412,N_9575);
and U9639 (N_9639,N_9469,N_9579);
xor U9640 (N_9640,N_9456,N_9553);
nor U9641 (N_9641,N_9499,N_9455);
and U9642 (N_9642,N_9510,N_9429);
nand U9643 (N_9643,N_9473,N_9542);
xor U9644 (N_9644,N_9586,N_9509);
nor U9645 (N_9645,N_9562,N_9446);
or U9646 (N_9646,N_9434,N_9564);
xor U9647 (N_9647,N_9597,N_9421);
nand U9648 (N_9648,N_9502,N_9527);
or U9649 (N_9649,N_9537,N_9495);
and U9650 (N_9650,N_9433,N_9507);
and U9651 (N_9651,N_9464,N_9428);
nor U9652 (N_9652,N_9492,N_9599);
nor U9653 (N_9653,N_9516,N_9441);
nor U9654 (N_9654,N_9500,N_9470);
or U9655 (N_9655,N_9535,N_9437);
nor U9656 (N_9656,N_9405,N_9400);
and U9657 (N_9657,N_9454,N_9449);
nor U9658 (N_9658,N_9482,N_9522);
and U9659 (N_9659,N_9517,N_9524);
nor U9660 (N_9660,N_9447,N_9576);
xor U9661 (N_9661,N_9595,N_9491);
or U9662 (N_9662,N_9539,N_9584);
nor U9663 (N_9663,N_9463,N_9490);
nor U9664 (N_9664,N_9430,N_9423);
xnor U9665 (N_9665,N_9483,N_9410);
nand U9666 (N_9666,N_9585,N_9572);
nand U9667 (N_9667,N_9460,N_9498);
nor U9668 (N_9668,N_9414,N_9505);
or U9669 (N_9669,N_9439,N_9419);
xor U9670 (N_9670,N_9514,N_9561);
xor U9671 (N_9671,N_9571,N_9583);
nand U9672 (N_9672,N_9526,N_9598);
nor U9673 (N_9673,N_9477,N_9587);
or U9674 (N_9674,N_9591,N_9465);
or U9675 (N_9675,N_9406,N_9440);
and U9676 (N_9676,N_9552,N_9541);
and U9677 (N_9677,N_9476,N_9462);
or U9678 (N_9678,N_9415,N_9590);
xor U9679 (N_9679,N_9427,N_9548);
or U9680 (N_9680,N_9593,N_9484);
xor U9681 (N_9681,N_9448,N_9589);
or U9682 (N_9682,N_9523,N_9401);
nand U9683 (N_9683,N_9431,N_9547);
nand U9684 (N_9684,N_9402,N_9444);
or U9685 (N_9685,N_9543,N_9556);
and U9686 (N_9686,N_9497,N_9472);
nand U9687 (N_9687,N_9555,N_9407);
xnor U9688 (N_9688,N_9580,N_9417);
nand U9689 (N_9689,N_9551,N_9435);
xnor U9690 (N_9690,N_9515,N_9508);
or U9691 (N_9691,N_9544,N_9581);
nor U9692 (N_9692,N_9451,N_9518);
or U9693 (N_9693,N_9557,N_9471);
or U9694 (N_9694,N_9496,N_9436);
nor U9695 (N_9695,N_9425,N_9404);
xnor U9696 (N_9696,N_9475,N_9588);
xnor U9697 (N_9697,N_9413,N_9554);
nand U9698 (N_9698,N_9445,N_9538);
xnor U9699 (N_9699,N_9563,N_9582);
and U9700 (N_9700,N_9509,N_9591);
or U9701 (N_9701,N_9410,N_9518);
and U9702 (N_9702,N_9518,N_9535);
and U9703 (N_9703,N_9515,N_9544);
nor U9704 (N_9704,N_9461,N_9450);
and U9705 (N_9705,N_9441,N_9515);
or U9706 (N_9706,N_9554,N_9483);
xnor U9707 (N_9707,N_9554,N_9451);
xor U9708 (N_9708,N_9498,N_9473);
or U9709 (N_9709,N_9479,N_9403);
nor U9710 (N_9710,N_9560,N_9462);
nor U9711 (N_9711,N_9556,N_9565);
or U9712 (N_9712,N_9508,N_9479);
and U9713 (N_9713,N_9438,N_9476);
nand U9714 (N_9714,N_9444,N_9484);
nand U9715 (N_9715,N_9521,N_9578);
or U9716 (N_9716,N_9450,N_9577);
nor U9717 (N_9717,N_9597,N_9437);
nor U9718 (N_9718,N_9582,N_9459);
nand U9719 (N_9719,N_9444,N_9556);
and U9720 (N_9720,N_9470,N_9552);
or U9721 (N_9721,N_9533,N_9537);
nand U9722 (N_9722,N_9447,N_9524);
nor U9723 (N_9723,N_9453,N_9481);
nand U9724 (N_9724,N_9521,N_9472);
or U9725 (N_9725,N_9405,N_9527);
nand U9726 (N_9726,N_9503,N_9495);
and U9727 (N_9727,N_9463,N_9416);
or U9728 (N_9728,N_9551,N_9509);
xnor U9729 (N_9729,N_9534,N_9506);
xnor U9730 (N_9730,N_9480,N_9430);
and U9731 (N_9731,N_9417,N_9466);
xnor U9732 (N_9732,N_9440,N_9449);
or U9733 (N_9733,N_9408,N_9520);
nand U9734 (N_9734,N_9549,N_9568);
nor U9735 (N_9735,N_9509,N_9502);
nand U9736 (N_9736,N_9581,N_9435);
nand U9737 (N_9737,N_9533,N_9444);
or U9738 (N_9738,N_9562,N_9458);
or U9739 (N_9739,N_9401,N_9493);
xor U9740 (N_9740,N_9520,N_9589);
nor U9741 (N_9741,N_9589,N_9444);
and U9742 (N_9742,N_9440,N_9412);
nor U9743 (N_9743,N_9564,N_9553);
nand U9744 (N_9744,N_9424,N_9509);
xor U9745 (N_9745,N_9478,N_9493);
nand U9746 (N_9746,N_9468,N_9436);
and U9747 (N_9747,N_9574,N_9511);
nor U9748 (N_9748,N_9592,N_9599);
xnor U9749 (N_9749,N_9573,N_9418);
and U9750 (N_9750,N_9406,N_9457);
nand U9751 (N_9751,N_9491,N_9576);
or U9752 (N_9752,N_9585,N_9514);
xor U9753 (N_9753,N_9407,N_9491);
or U9754 (N_9754,N_9594,N_9417);
nand U9755 (N_9755,N_9591,N_9598);
or U9756 (N_9756,N_9493,N_9507);
nor U9757 (N_9757,N_9409,N_9403);
or U9758 (N_9758,N_9587,N_9424);
or U9759 (N_9759,N_9523,N_9556);
and U9760 (N_9760,N_9440,N_9567);
or U9761 (N_9761,N_9451,N_9460);
and U9762 (N_9762,N_9562,N_9596);
nor U9763 (N_9763,N_9546,N_9544);
and U9764 (N_9764,N_9540,N_9513);
xnor U9765 (N_9765,N_9469,N_9426);
or U9766 (N_9766,N_9543,N_9574);
and U9767 (N_9767,N_9457,N_9532);
nand U9768 (N_9768,N_9519,N_9534);
nand U9769 (N_9769,N_9425,N_9509);
xnor U9770 (N_9770,N_9539,N_9569);
or U9771 (N_9771,N_9523,N_9499);
nand U9772 (N_9772,N_9486,N_9518);
nor U9773 (N_9773,N_9494,N_9448);
and U9774 (N_9774,N_9581,N_9579);
nor U9775 (N_9775,N_9485,N_9498);
xor U9776 (N_9776,N_9594,N_9587);
nand U9777 (N_9777,N_9597,N_9519);
xor U9778 (N_9778,N_9533,N_9590);
or U9779 (N_9779,N_9435,N_9588);
xnor U9780 (N_9780,N_9515,N_9540);
and U9781 (N_9781,N_9486,N_9581);
nor U9782 (N_9782,N_9413,N_9558);
xor U9783 (N_9783,N_9419,N_9491);
nand U9784 (N_9784,N_9481,N_9508);
nor U9785 (N_9785,N_9477,N_9556);
nand U9786 (N_9786,N_9556,N_9535);
nand U9787 (N_9787,N_9516,N_9454);
and U9788 (N_9788,N_9460,N_9446);
and U9789 (N_9789,N_9523,N_9550);
nor U9790 (N_9790,N_9582,N_9513);
nor U9791 (N_9791,N_9418,N_9424);
nand U9792 (N_9792,N_9552,N_9587);
nand U9793 (N_9793,N_9406,N_9548);
nand U9794 (N_9794,N_9578,N_9510);
nor U9795 (N_9795,N_9481,N_9512);
nor U9796 (N_9796,N_9547,N_9494);
and U9797 (N_9797,N_9483,N_9573);
and U9798 (N_9798,N_9443,N_9494);
nand U9799 (N_9799,N_9512,N_9438);
nor U9800 (N_9800,N_9799,N_9606);
xnor U9801 (N_9801,N_9621,N_9673);
nor U9802 (N_9802,N_9603,N_9733);
xnor U9803 (N_9803,N_9792,N_9612);
xor U9804 (N_9804,N_9678,N_9648);
and U9805 (N_9805,N_9778,N_9705);
nor U9806 (N_9806,N_9746,N_9737);
xor U9807 (N_9807,N_9753,N_9661);
and U9808 (N_9808,N_9695,N_9747);
and U9809 (N_9809,N_9738,N_9706);
nand U9810 (N_9810,N_9600,N_9611);
and U9811 (N_9811,N_9759,N_9787);
xnor U9812 (N_9812,N_9666,N_9729);
and U9813 (N_9813,N_9686,N_9779);
xor U9814 (N_9814,N_9632,N_9637);
nand U9815 (N_9815,N_9623,N_9745);
nor U9816 (N_9816,N_9700,N_9780);
and U9817 (N_9817,N_9707,N_9683);
nor U9818 (N_9818,N_9616,N_9735);
xor U9819 (N_9819,N_9667,N_9702);
and U9820 (N_9820,N_9719,N_9676);
nand U9821 (N_9821,N_9766,N_9631);
and U9822 (N_9822,N_9642,N_9756);
and U9823 (N_9823,N_9675,N_9658);
xor U9824 (N_9824,N_9767,N_9730);
or U9825 (N_9825,N_9722,N_9660);
nor U9826 (N_9826,N_9643,N_9717);
nor U9827 (N_9827,N_9723,N_9758);
xor U9828 (N_9828,N_9679,N_9755);
and U9829 (N_9829,N_9699,N_9728);
and U9830 (N_9830,N_9622,N_9605);
nor U9831 (N_9831,N_9774,N_9689);
nand U9832 (N_9832,N_9647,N_9610);
xnor U9833 (N_9833,N_9752,N_9639);
and U9834 (N_9834,N_9732,N_9633);
nor U9835 (N_9835,N_9649,N_9727);
nand U9836 (N_9836,N_9682,N_9688);
nand U9837 (N_9837,N_9736,N_9665);
and U9838 (N_9838,N_9794,N_9762);
or U9839 (N_9839,N_9628,N_9795);
and U9840 (N_9840,N_9760,N_9771);
xnor U9841 (N_9841,N_9655,N_9789);
xor U9842 (N_9842,N_9772,N_9798);
nand U9843 (N_9843,N_9671,N_9783);
and U9844 (N_9844,N_9615,N_9731);
nand U9845 (N_9845,N_9697,N_9634);
nand U9846 (N_9846,N_9650,N_9761);
nor U9847 (N_9847,N_9663,N_9742);
nand U9848 (N_9848,N_9784,N_9711);
nand U9849 (N_9849,N_9716,N_9652);
xnor U9850 (N_9850,N_9629,N_9751);
nor U9851 (N_9851,N_9687,N_9749);
and U9852 (N_9852,N_9786,N_9684);
xnor U9853 (N_9853,N_9659,N_9776);
nor U9854 (N_9854,N_9692,N_9657);
and U9855 (N_9855,N_9651,N_9710);
nor U9856 (N_9856,N_9635,N_9785);
nor U9857 (N_9857,N_9741,N_9703);
nand U9858 (N_9858,N_9626,N_9765);
nand U9859 (N_9859,N_9793,N_9754);
xor U9860 (N_9860,N_9725,N_9768);
nor U9861 (N_9861,N_9654,N_9627);
or U9862 (N_9862,N_9790,N_9644);
nand U9863 (N_9863,N_9690,N_9617);
nand U9864 (N_9864,N_9734,N_9693);
nand U9865 (N_9865,N_9625,N_9618);
or U9866 (N_9866,N_9636,N_9721);
nand U9867 (N_9867,N_9613,N_9630);
and U9868 (N_9868,N_9718,N_9641);
nand U9869 (N_9869,N_9694,N_9638);
xor U9870 (N_9870,N_9724,N_9664);
or U9871 (N_9871,N_9764,N_9775);
or U9872 (N_9872,N_9743,N_9614);
or U9873 (N_9873,N_9669,N_9662);
and U9874 (N_9874,N_9773,N_9796);
xnor U9875 (N_9875,N_9653,N_9791);
nor U9876 (N_9876,N_9640,N_9712);
and U9877 (N_9877,N_9645,N_9704);
nand U9878 (N_9878,N_9701,N_9619);
nor U9879 (N_9879,N_9708,N_9696);
or U9880 (N_9880,N_9750,N_9607);
nor U9881 (N_9881,N_9770,N_9726);
xnor U9882 (N_9882,N_9715,N_9757);
or U9883 (N_9883,N_9601,N_9698);
or U9884 (N_9884,N_9670,N_9685);
xnor U9885 (N_9885,N_9620,N_9624);
and U9886 (N_9886,N_9691,N_9714);
xnor U9887 (N_9887,N_9604,N_9608);
or U9888 (N_9888,N_9781,N_9609);
or U9889 (N_9889,N_9674,N_9677);
or U9890 (N_9890,N_9681,N_9797);
nor U9891 (N_9891,N_9709,N_9713);
and U9892 (N_9892,N_9720,N_9763);
nand U9893 (N_9893,N_9777,N_9672);
nor U9894 (N_9894,N_9646,N_9788);
and U9895 (N_9895,N_9680,N_9782);
nor U9896 (N_9896,N_9739,N_9744);
and U9897 (N_9897,N_9602,N_9668);
or U9898 (N_9898,N_9740,N_9748);
xor U9899 (N_9899,N_9656,N_9769);
and U9900 (N_9900,N_9755,N_9783);
and U9901 (N_9901,N_9777,N_9756);
and U9902 (N_9902,N_9690,N_9607);
xor U9903 (N_9903,N_9799,N_9747);
xor U9904 (N_9904,N_9724,N_9686);
or U9905 (N_9905,N_9776,N_9608);
and U9906 (N_9906,N_9784,N_9626);
nand U9907 (N_9907,N_9751,N_9753);
nand U9908 (N_9908,N_9685,N_9751);
and U9909 (N_9909,N_9778,N_9725);
nor U9910 (N_9910,N_9677,N_9786);
nor U9911 (N_9911,N_9657,N_9636);
and U9912 (N_9912,N_9632,N_9625);
nand U9913 (N_9913,N_9628,N_9622);
xor U9914 (N_9914,N_9684,N_9673);
or U9915 (N_9915,N_9673,N_9755);
or U9916 (N_9916,N_9693,N_9757);
nand U9917 (N_9917,N_9748,N_9755);
and U9918 (N_9918,N_9675,N_9691);
or U9919 (N_9919,N_9655,N_9688);
or U9920 (N_9920,N_9676,N_9786);
nand U9921 (N_9921,N_9657,N_9789);
xnor U9922 (N_9922,N_9772,N_9709);
nand U9923 (N_9923,N_9623,N_9748);
xnor U9924 (N_9924,N_9709,N_9655);
or U9925 (N_9925,N_9748,N_9625);
and U9926 (N_9926,N_9652,N_9677);
or U9927 (N_9927,N_9725,N_9741);
xnor U9928 (N_9928,N_9658,N_9730);
nand U9929 (N_9929,N_9635,N_9654);
xnor U9930 (N_9930,N_9668,N_9719);
and U9931 (N_9931,N_9613,N_9709);
or U9932 (N_9932,N_9734,N_9625);
or U9933 (N_9933,N_9696,N_9772);
nor U9934 (N_9934,N_9630,N_9727);
nand U9935 (N_9935,N_9738,N_9709);
xor U9936 (N_9936,N_9698,N_9795);
or U9937 (N_9937,N_9798,N_9655);
nor U9938 (N_9938,N_9691,N_9696);
xnor U9939 (N_9939,N_9673,N_9789);
xor U9940 (N_9940,N_9698,N_9639);
nand U9941 (N_9941,N_9785,N_9662);
nand U9942 (N_9942,N_9772,N_9766);
nand U9943 (N_9943,N_9627,N_9616);
xnor U9944 (N_9944,N_9720,N_9781);
nand U9945 (N_9945,N_9651,N_9680);
and U9946 (N_9946,N_9760,N_9751);
or U9947 (N_9947,N_9773,N_9705);
or U9948 (N_9948,N_9610,N_9773);
nand U9949 (N_9949,N_9631,N_9692);
nand U9950 (N_9950,N_9772,N_9609);
xnor U9951 (N_9951,N_9661,N_9785);
and U9952 (N_9952,N_9739,N_9603);
nor U9953 (N_9953,N_9760,N_9690);
xnor U9954 (N_9954,N_9612,N_9632);
xnor U9955 (N_9955,N_9713,N_9626);
nor U9956 (N_9956,N_9664,N_9659);
or U9957 (N_9957,N_9722,N_9627);
nand U9958 (N_9958,N_9767,N_9657);
nor U9959 (N_9959,N_9649,N_9713);
and U9960 (N_9960,N_9624,N_9747);
xnor U9961 (N_9961,N_9653,N_9688);
xor U9962 (N_9962,N_9776,N_9619);
and U9963 (N_9963,N_9661,N_9788);
nand U9964 (N_9964,N_9647,N_9672);
and U9965 (N_9965,N_9711,N_9750);
xnor U9966 (N_9966,N_9612,N_9694);
or U9967 (N_9967,N_9778,N_9682);
nand U9968 (N_9968,N_9782,N_9608);
nand U9969 (N_9969,N_9639,N_9732);
and U9970 (N_9970,N_9625,N_9639);
nand U9971 (N_9971,N_9684,N_9628);
and U9972 (N_9972,N_9623,N_9634);
nand U9973 (N_9973,N_9643,N_9793);
and U9974 (N_9974,N_9663,N_9775);
nor U9975 (N_9975,N_9762,N_9659);
nor U9976 (N_9976,N_9705,N_9765);
or U9977 (N_9977,N_9702,N_9759);
nand U9978 (N_9978,N_9752,N_9603);
nand U9979 (N_9979,N_9709,N_9600);
nand U9980 (N_9980,N_9633,N_9798);
xor U9981 (N_9981,N_9797,N_9786);
nor U9982 (N_9982,N_9798,N_9785);
or U9983 (N_9983,N_9658,N_9663);
xor U9984 (N_9984,N_9722,N_9766);
xnor U9985 (N_9985,N_9613,N_9675);
nand U9986 (N_9986,N_9620,N_9645);
nand U9987 (N_9987,N_9773,N_9675);
and U9988 (N_9988,N_9716,N_9784);
nor U9989 (N_9989,N_9715,N_9699);
or U9990 (N_9990,N_9755,N_9627);
or U9991 (N_9991,N_9657,N_9694);
or U9992 (N_9992,N_9685,N_9723);
and U9993 (N_9993,N_9723,N_9647);
xnor U9994 (N_9994,N_9623,N_9687);
xor U9995 (N_9995,N_9616,N_9677);
nand U9996 (N_9996,N_9728,N_9676);
xnor U9997 (N_9997,N_9746,N_9780);
nand U9998 (N_9998,N_9771,N_9725);
nand U9999 (N_9999,N_9738,N_9756);
xnor U10000 (N_10000,N_9844,N_9880);
nand U10001 (N_10001,N_9997,N_9921);
nor U10002 (N_10002,N_9899,N_9900);
nor U10003 (N_10003,N_9989,N_9848);
or U10004 (N_10004,N_9864,N_9819);
nor U10005 (N_10005,N_9872,N_9878);
or U10006 (N_10006,N_9901,N_9926);
xor U10007 (N_10007,N_9811,N_9874);
or U10008 (N_10008,N_9923,N_9852);
nand U10009 (N_10009,N_9807,N_9939);
nor U10010 (N_10010,N_9858,N_9902);
xnor U10011 (N_10011,N_9812,N_9962);
and U10012 (N_10012,N_9938,N_9860);
nand U10013 (N_10013,N_9914,N_9886);
xnor U10014 (N_10014,N_9933,N_9868);
or U10015 (N_10015,N_9907,N_9995);
nor U10016 (N_10016,N_9806,N_9961);
xnor U10017 (N_10017,N_9840,N_9972);
or U10018 (N_10018,N_9959,N_9920);
and U10019 (N_10019,N_9913,N_9835);
nand U10020 (N_10020,N_9814,N_9982);
or U10021 (N_10021,N_9911,N_9969);
nand U10022 (N_10022,N_9897,N_9802);
xnor U10023 (N_10023,N_9871,N_9905);
nand U10024 (N_10024,N_9968,N_9955);
nor U10025 (N_10025,N_9936,N_9849);
and U10026 (N_10026,N_9953,N_9946);
nand U10027 (N_10027,N_9964,N_9949);
and U10028 (N_10028,N_9931,N_9836);
and U10029 (N_10029,N_9838,N_9887);
and U10030 (N_10030,N_9925,N_9956);
or U10031 (N_10031,N_9855,N_9915);
and U10032 (N_10032,N_9842,N_9825);
xnor U10033 (N_10033,N_9948,N_9862);
nor U10034 (N_10034,N_9865,N_9869);
nand U10035 (N_10035,N_9824,N_9859);
or U10036 (N_10036,N_9975,N_9832);
nor U10037 (N_10037,N_9940,N_9996);
nor U10038 (N_10038,N_9892,N_9954);
nor U10039 (N_10039,N_9934,N_9909);
nor U10040 (N_10040,N_9831,N_9922);
and U10041 (N_10041,N_9800,N_9820);
or U10042 (N_10042,N_9957,N_9808);
xor U10043 (N_10043,N_9980,N_9804);
or U10044 (N_10044,N_9993,N_9830);
nand U10045 (N_10045,N_9834,N_9984);
nor U10046 (N_10046,N_9932,N_9809);
and U10047 (N_10047,N_9906,N_9861);
xor U10048 (N_10048,N_9937,N_9942);
nand U10049 (N_10049,N_9882,N_9994);
or U10050 (N_10050,N_9981,N_9884);
xnor U10051 (N_10051,N_9891,N_9875);
and U10052 (N_10052,N_9960,N_9965);
nand U10053 (N_10053,N_9904,N_9847);
xor U10054 (N_10054,N_9898,N_9843);
nand U10055 (N_10055,N_9813,N_9983);
xor U10056 (N_10056,N_9998,N_9851);
nand U10057 (N_10057,N_9927,N_9826);
and U10058 (N_10058,N_9893,N_9990);
or U10059 (N_10059,N_9896,N_9895);
nand U10060 (N_10060,N_9815,N_9818);
and U10061 (N_10061,N_9928,N_9822);
nand U10062 (N_10062,N_9816,N_9857);
nor U10063 (N_10063,N_9979,N_9917);
nand U10064 (N_10064,N_9870,N_9919);
or U10065 (N_10065,N_9973,N_9890);
nor U10066 (N_10066,N_9866,N_9967);
xor U10067 (N_10067,N_9903,N_9951);
nand U10068 (N_10068,N_9889,N_9856);
xor U10069 (N_10069,N_9991,N_9867);
nor U10070 (N_10070,N_9883,N_9810);
and U10071 (N_10071,N_9837,N_9879);
or U10072 (N_10072,N_9978,N_9918);
xnor U10073 (N_10073,N_9801,N_9988);
and U10074 (N_10074,N_9841,N_9952);
xor U10075 (N_10075,N_9924,N_9823);
or U10076 (N_10076,N_9916,N_9910);
or U10077 (N_10077,N_9987,N_9873);
or U10078 (N_10078,N_9929,N_9912);
and U10079 (N_10079,N_9821,N_9992);
or U10080 (N_10080,N_9976,N_9950);
and U10081 (N_10081,N_9963,N_9827);
nor U10082 (N_10082,N_9985,N_9945);
and U10083 (N_10083,N_9894,N_9908);
xnor U10084 (N_10084,N_9947,N_9881);
and U10085 (N_10085,N_9944,N_9888);
nand U10086 (N_10086,N_9941,N_9833);
nand U10087 (N_10087,N_9966,N_9829);
or U10088 (N_10088,N_9828,N_9817);
nand U10089 (N_10089,N_9986,N_9943);
or U10090 (N_10090,N_9850,N_9876);
nor U10091 (N_10091,N_9885,N_9846);
nor U10092 (N_10092,N_9845,N_9958);
and U10093 (N_10093,N_9863,N_9999);
nor U10094 (N_10094,N_9854,N_9803);
nand U10095 (N_10095,N_9877,N_9970);
or U10096 (N_10096,N_9853,N_9935);
nor U10097 (N_10097,N_9930,N_9977);
nor U10098 (N_10098,N_9971,N_9839);
nand U10099 (N_10099,N_9805,N_9974);
nor U10100 (N_10100,N_9984,N_9949);
xnor U10101 (N_10101,N_9946,N_9988);
xor U10102 (N_10102,N_9858,N_9877);
nor U10103 (N_10103,N_9925,N_9941);
or U10104 (N_10104,N_9930,N_9852);
or U10105 (N_10105,N_9893,N_9985);
nand U10106 (N_10106,N_9999,N_9991);
xor U10107 (N_10107,N_9872,N_9963);
and U10108 (N_10108,N_9838,N_9854);
nand U10109 (N_10109,N_9981,N_9808);
nand U10110 (N_10110,N_9883,N_9923);
nor U10111 (N_10111,N_9917,N_9906);
or U10112 (N_10112,N_9938,N_9845);
xnor U10113 (N_10113,N_9837,N_9905);
nor U10114 (N_10114,N_9875,N_9997);
or U10115 (N_10115,N_9891,N_9877);
nor U10116 (N_10116,N_9891,N_9964);
nand U10117 (N_10117,N_9920,N_9845);
or U10118 (N_10118,N_9946,N_9936);
xnor U10119 (N_10119,N_9891,N_9955);
nor U10120 (N_10120,N_9922,N_9941);
nor U10121 (N_10121,N_9825,N_9828);
nor U10122 (N_10122,N_9985,N_9995);
nor U10123 (N_10123,N_9807,N_9947);
nor U10124 (N_10124,N_9870,N_9908);
or U10125 (N_10125,N_9803,N_9914);
nand U10126 (N_10126,N_9990,N_9978);
xnor U10127 (N_10127,N_9901,N_9866);
xnor U10128 (N_10128,N_9814,N_9933);
xor U10129 (N_10129,N_9894,N_9873);
xnor U10130 (N_10130,N_9985,N_9962);
nor U10131 (N_10131,N_9923,N_9880);
nor U10132 (N_10132,N_9995,N_9962);
xnor U10133 (N_10133,N_9845,N_9863);
nand U10134 (N_10134,N_9818,N_9821);
nor U10135 (N_10135,N_9979,N_9895);
xor U10136 (N_10136,N_9962,N_9956);
and U10137 (N_10137,N_9921,N_9949);
xnor U10138 (N_10138,N_9830,N_9961);
xor U10139 (N_10139,N_9808,N_9972);
nor U10140 (N_10140,N_9910,N_9929);
nor U10141 (N_10141,N_9987,N_9975);
and U10142 (N_10142,N_9874,N_9976);
and U10143 (N_10143,N_9937,N_9848);
or U10144 (N_10144,N_9851,N_9873);
nand U10145 (N_10145,N_9885,N_9974);
or U10146 (N_10146,N_9986,N_9952);
xor U10147 (N_10147,N_9804,N_9891);
xor U10148 (N_10148,N_9969,N_9985);
xor U10149 (N_10149,N_9828,N_9957);
and U10150 (N_10150,N_9843,N_9864);
and U10151 (N_10151,N_9838,N_9911);
nor U10152 (N_10152,N_9854,N_9932);
or U10153 (N_10153,N_9838,N_9972);
and U10154 (N_10154,N_9974,N_9963);
xor U10155 (N_10155,N_9923,N_9805);
or U10156 (N_10156,N_9977,N_9984);
or U10157 (N_10157,N_9975,N_9994);
and U10158 (N_10158,N_9987,N_9995);
nand U10159 (N_10159,N_9810,N_9910);
xor U10160 (N_10160,N_9959,N_9853);
nand U10161 (N_10161,N_9890,N_9923);
or U10162 (N_10162,N_9979,N_9835);
and U10163 (N_10163,N_9914,N_9838);
nor U10164 (N_10164,N_9846,N_9872);
nor U10165 (N_10165,N_9862,N_9806);
or U10166 (N_10166,N_9811,N_9944);
xnor U10167 (N_10167,N_9894,N_9863);
and U10168 (N_10168,N_9971,N_9924);
or U10169 (N_10169,N_9926,N_9879);
or U10170 (N_10170,N_9812,N_9898);
nor U10171 (N_10171,N_9909,N_9835);
or U10172 (N_10172,N_9961,N_9933);
and U10173 (N_10173,N_9964,N_9859);
nor U10174 (N_10174,N_9860,N_9820);
nand U10175 (N_10175,N_9965,N_9972);
nand U10176 (N_10176,N_9897,N_9963);
xnor U10177 (N_10177,N_9949,N_9853);
and U10178 (N_10178,N_9918,N_9816);
and U10179 (N_10179,N_9855,N_9806);
nor U10180 (N_10180,N_9850,N_9816);
and U10181 (N_10181,N_9976,N_9841);
nor U10182 (N_10182,N_9836,N_9885);
nand U10183 (N_10183,N_9983,N_9869);
xor U10184 (N_10184,N_9991,N_9938);
nor U10185 (N_10185,N_9918,N_9942);
nor U10186 (N_10186,N_9811,N_9965);
and U10187 (N_10187,N_9977,N_9815);
nor U10188 (N_10188,N_9814,N_9880);
nand U10189 (N_10189,N_9946,N_9808);
nor U10190 (N_10190,N_9917,N_9836);
xnor U10191 (N_10191,N_9993,N_9983);
or U10192 (N_10192,N_9891,N_9862);
and U10193 (N_10193,N_9858,N_9971);
or U10194 (N_10194,N_9855,N_9948);
xnor U10195 (N_10195,N_9888,N_9927);
nor U10196 (N_10196,N_9884,N_9940);
nand U10197 (N_10197,N_9831,N_9880);
or U10198 (N_10198,N_9915,N_9877);
or U10199 (N_10199,N_9870,N_9932);
and U10200 (N_10200,N_10036,N_10144);
or U10201 (N_10201,N_10004,N_10106);
and U10202 (N_10202,N_10085,N_10142);
xor U10203 (N_10203,N_10131,N_10133);
nand U10204 (N_10204,N_10155,N_10068);
and U10205 (N_10205,N_10025,N_10043);
nand U10206 (N_10206,N_10084,N_10054);
or U10207 (N_10207,N_10180,N_10049);
nand U10208 (N_10208,N_10078,N_10058);
nor U10209 (N_10209,N_10127,N_10121);
and U10210 (N_10210,N_10037,N_10104);
nor U10211 (N_10211,N_10022,N_10010);
or U10212 (N_10212,N_10097,N_10169);
and U10213 (N_10213,N_10075,N_10108);
and U10214 (N_10214,N_10184,N_10015);
and U10215 (N_10215,N_10129,N_10044);
nand U10216 (N_10216,N_10113,N_10070);
and U10217 (N_10217,N_10136,N_10159);
nand U10218 (N_10218,N_10164,N_10197);
nor U10219 (N_10219,N_10008,N_10165);
xor U10220 (N_10220,N_10089,N_10107);
nor U10221 (N_10221,N_10065,N_10178);
and U10222 (N_10222,N_10094,N_10125);
or U10223 (N_10223,N_10048,N_10031);
or U10224 (N_10224,N_10013,N_10040);
and U10225 (N_10225,N_10064,N_10011);
and U10226 (N_10226,N_10069,N_10161);
or U10227 (N_10227,N_10172,N_10141);
and U10228 (N_10228,N_10117,N_10122);
nand U10229 (N_10229,N_10187,N_10077);
and U10230 (N_10230,N_10196,N_10096);
or U10231 (N_10231,N_10134,N_10021);
nand U10232 (N_10232,N_10063,N_10111);
and U10233 (N_10233,N_10192,N_10073);
or U10234 (N_10234,N_10060,N_10055);
nor U10235 (N_10235,N_10023,N_10081);
nor U10236 (N_10236,N_10098,N_10140);
nor U10237 (N_10237,N_10170,N_10193);
nand U10238 (N_10238,N_10183,N_10100);
nand U10239 (N_10239,N_10000,N_10088);
nor U10240 (N_10240,N_10188,N_10191);
xor U10241 (N_10241,N_10057,N_10001);
and U10242 (N_10242,N_10119,N_10083);
xnor U10243 (N_10243,N_10150,N_10124);
or U10244 (N_10244,N_10090,N_10130);
xnor U10245 (N_10245,N_10115,N_10110);
xnor U10246 (N_10246,N_10128,N_10116);
or U10247 (N_10247,N_10032,N_10092);
and U10248 (N_10248,N_10093,N_10059);
and U10249 (N_10249,N_10035,N_10042);
or U10250 (N_10250,N_10151,N_10038);
or U10251 (N_10251,N_10074,N_10135);
nand U10252 (N_10252,N_10157,N_10030);
nor U10253 (N_10253,N_10146,N_10095);
nand U10254 (N_10254,N_10179,N_10166);
nand U10255 (N_10255,N_10195,N_10052);
or U10256 (N_10256,N_10174,N_10175);
nor U10257 (N_10257,N_10171,N_10012);
xnor U10258 (N_10258,N_10123,N_10138);
and U10259 (N_10259,N_10027,N_10160);
xor U10260 (N_10260,N_10087,N_10158);
xnor U10261 (N_10261,N_10062,N_10009);
xnor U10262 (N_10262,N_10053,N_10148);
xnor U10263 (N_10263,N_10024,N_10120);
and U10264 (N_10264,N_10041,N_10154);
xnor U10265 (N_10265,N_10047,N_10143);
xnor U10266 (N_10266,N_10051,N_10003);
xnor U10267 (N_10267,N_10002,N_10016);
nor U10268 (N_10268,N_10005,N_10198);
and U10269 (N_10269,N_10071,N_10176);
nand U10270 (N_10270,N_10105,N_10020);
and U10271 (N_10271,N_10039,N_10149);
nand U10272 (N_10272,N_10029,N_10181);
or U10273 (N_10273,N_10173,N_10006);
and U10274 (N_10274,N_10050,N_10018);
nor U10275 (N_10275,N_10079,N_10034);
xor U10276 (N_10276,N_10137,N_10102);
and U10277 (N_10277,N_10182,N_10112);
nor U10278 (N_10278,N_10163,N_10091);
nand U10279 (N_10279,N_10067,N_10177);
and U10280 (N_10280,N_10033,N_10152);
nand U10281 (N_10281,N_10145,N_10019);
nor U10282 (N_10282,N_10118,N_10153);
nand U10283 (N_10283,N_10028,N_10076);
xnor U10284 (N_10284,N_10168,N_10026);
nor U10285 (N_10285,N_10194,N_10156);
nor U10286 (N_10286,N_10086,N_10046);
xor U10287 (N_10287,N_10014,N_10185);
xor U10288 (N_10288,N_10132,N_10056);
xnor U10289 (N_10289,N_10007,N_10189);
or U10290 (N_10290,N_10114,N_10147);
nand U10291 (N_10291,N_10162,N_10072);
and U10292 (N_10292,N_10099,N_10080);
nand U10293 (N_10293,N_10186,N_10199);
nor U10294 (N_10294,N_10190,N_10045);
and U10295 (N_10295,N_10126,N_10139);
and U10296 (N_10296,N_10109,N_10061);
nor U10297 (N_10297,N_10101,N_10017);
xor U10298 (N_10298,N_10103,N_10082);
nand U10299 (N_10299,N_10066,N_10167);
nand U10300 (N_10300,N_10189,N_10137);
or U10301 (N_10301,N_10134,N_10156);
or U10302 (N_10302,N_10005,N_10028);
and U10303 (N_10303,N_10077,N_10090);
or U10304 (N_10304,N_10154,N_10151);
and U10305 (N_10305,N_10083,N_10013);
nand U10306 (N_10306,N_10168,N_10022);
nand U10307 (N_10307,N_10143,N_10157);
nor U10308 (N_10308,N_10054,N_10044);
nor U10309 (N_10309,N_10077,N_10023);
or U10310 (N_10310,N_10098,N_10074);
nor U10311 (N_10311,N_10197,N_10057);
nand U10312 (N_10312,N_10194,N_10115);
or U10313 (N_10313,N_10067,N_10065);
or U10314 (N_10314,N_10146,N_10103);
nand U10315 (N_10315,N_10066,N_10086);
or U10316 (N_10316,N_10111,N_10036);
xnor U10317 (N_10317,N_10006,N_10067);
nor U10318 (N_10318,N_10035,N_10080);
nand U10319 (N_10319,N_10198,N_10116);
or U10320 (N_10320,N_10189,N_10174);
and U10321 (N_10321,N_10130,N_10028);
nor U10322 (N_10322,N_10161,N_10153);
nor U10323 (N_10323,N_10195,N_10162);
xnor U10324 (N_10324,N_10146,N_10108);
xor U10325 (N_10325,N_10168,N_10137);
xor U10326 (N_10326,N_10167,N_10061);
nand U10327 (N_10327,N_10014,N_10123);
xor U10328 (N_10328,N_10001,N_10037);
or U10329 (N_10329,N_10089,N_10035);
nand U10330 (N_10330,N_10118,N_10149);
nand U10331 (N_10331,N_10101,N_10092);
and U10332 (N_10332,N_10163,N_10098);
or U10333 (N_10333,N_10025,N_10189);
or U10334 (N_10334,N_10159,N_10143);
and U10335 (N_10335,N_10143,N_10108);
or U10336 (N_10336,N_10119,N_10130);
xnor U10337 (N_10337,N_10067,N_10196);
nand U10338 (N_10338,N_10010,N_10150);
xor U10339 (N_10339,N_10144,N_10142);
and U10340 (N_10340,N_10060,N_10085);
nand U10341 (N_10341,N_10022,N_10071);
or U10342 (N_10342,N_10193,N_10100);
nor U10343 (N_10343,N_10075,N_10142);
nor U10344 (N_10344,N_10115,N_10111);
xor U10345 (N_10345,N_10078,N_10106);
or U10346 (N_10346,N_10042,N_10120);
or U10347 (N_10347,N_10016,N_10125);
xnor U10348 (N_10348,N_10174,N_10171);
nand U10349 (N_10349,N_10116,N_10090);
or U10350 (N_10350,N_10126,N_10052);
or U10351 (N_10351,N_10046,N_10039);
nand U10352 (N_10352,N_10103,N_10110);
or U10353 (N_10353,N_10163,N_10007);
and U10354 (N_10354,N_10188,N_10143);
nand U10355 (N_10355,N_10153,N_10038);
or U10356 (N_10356,N_10093,N_10058);
xor U10357 (N_10357,N_10146,N_10019);
xnor U10358 (N_10358,N_10034,N_10192);
or U10359 (N_10359,N_10199,N_10079);
or U10360 (N_10360,N_10026,N_10002);
nand U10361 (N_10361,N_10065,N_10169);
nand U10362 (N_10362,N_10123,N_10001);
nand U10363 (N_10363,N_10024,N_10157);
xnor U10364 (N_10364,N_10126,N_10120);
and U10365 (N_10365,N_10062,N_10003);
and U10366 (N_10366,N_10191,N_10155);
nor U10367 (N_10367,N_10165,N_10101);
xnor U10368 (N_10368,N_10077,N_10054);
xor U10369 (N_10369,N_10192,N_10163);
xor U10370 (N_10370,N_10161,N_10059);
nor U10371 (N_10371,N_10083,N_10002);
or U10372 (N_10372,N_10056,N_10094);
xor U10373 (N_10373,N_10048,N_10195);
or U10374 (N_10374,N_10119,N_10163);
nand U10375 (N_10375,N_10101,N_10115);
or U10376 (N_10376,N_10052,N_10136);
xor U10377 (N_10377,N_10116,N_10062);
nor U10378 (N_10378,N_10173,N_10188);
xor U10379 (N_10379,N_10162,N_10179);
and U10380 (N_10380,N_10179,N_10097);
nand U10381 (N_10381,N_10125,N_10165);
nor U10382 (N_10382,N_10045,N_10191);
or U10383 (N_10383,N_10001,N_10016);
nor U10384 (N_10384,N_10180,N_10161);
or U10385 (N_10385,N_10003,N_10034);
xnor U10386 (N_10386,N_10086,N_10103);
nand U10387 (N_10387,N_10134,N_10129);
or U10388 (N_10388,N_10135,N_10017);
and U10389 (N_10389,N_10072,N_10119);
or U10390 (N_10390,N_10128,N_10018);
xnor U10391 (N_10391,N_10137,N_10145);
and U10392 (N_10392,N_10121,N_10007);
or U10393 (N_10393,N_10046,N_10174);
xnor U10394 (N_10394,N_10091,N_10105);
xnor U10395 (N_10395,N_10165,N_10124);
nor U10396 (N_10396,N_10179,N_10016);
xnor U10397 (N_10397,N_10115,N_10124);
or U10398 (N_10398,N_10059,N_10116);
or U10399 (N_10399,N_10133,N_10096);
xor U10400 (N_10400,N_10248,N_10368);
and U10401 (N_10401,N_10317,N_10241);
and U10402 (N_10402,N_10348,N_10207);
nand U10403 (N_10403,N_10389,N_10236);
xor U10404 (N_10404,N_10204,N_10310);
and U10405 (N_10405,N_10315,N_10378);
nand U10406 (N_10406,N_10260,N_10230);
or U10407 (N_10407,N_10321,N_10395);
nor U10408 (N_10408,N_10250,N_10329);
nand U10409 (N_10409,N_10228,N_10373);
nor U10410 (N_10410,N_10278,N_10281);
or U10411 (N_10411,N_10209,N_10353);
nor U10412 (N_10412,N_10382,N_10301);
or U10413 (N_10413,N_10258,N_10326);
xnor U10414 (N_10414,N_10362,N_10202);
nand U10415 (N_10415,N_10351,N_10398);
nor U10416 (N_10416,N_10297,N_10215);
and U10417 (N_10417,N_10303,N_10219);
nor U10418 (N_10418,N_10399,N_10374);
xor U10419 (N_10419,N_10246,N_10232);
or U10420 (N_10420,N_10265,N_10300);
or U10421 (N_10421,N_10269,N_10377);
or U10422 (N_10422,N_10356,N_10305);
and U10423 (N_10423,N_10275,N_10358);
and U10424 (N_10424,N_10213,N_10299);
and U10425 (N_10425,N_10212,N_10397);
or U10426 (N_10426,N_10280,N_10396);
nand U10427 (N_10427,N_10314,N_10330);
and U10428 (N_10428,N_10239,N_10268);
nor U10429 (N_10429,N_10224,N_10355);
nor U10430 (N_10430,N_10393,N_10282);
nand U10431 (N_10431,N_10347,N_10283);
or U10432 (N_10432,N_10243,N_10302);
nand U10433 (N_10433,N_10231,N_10259);
xor U10434 (N_10434,N_10270,N_10341);
or U10435 (N_10435,N_10206,N_10263);
nor U10436 (N_10436,N_10257,N_10276);
and U10437 (N_10437,N_10294,N_10319);
nor U10438 (N_10438,N_10216,N_10376);
nor U10439 (N_10439,N_10237,N_10240);
nand U10440 (N_10440,N_10328,N_10284);
or U10441 (N_10441,N_10298,N_10203);
xor U10442 (N_10442,N_10322,N_10392);
nand U10443 (N_10443,N_10252,N_10244);
xor U10444 (N_10444,N_10226,N_10366);
or U10445 (N_10445,N_10293,N_10372);
xor U10446 (N_10446,N_10323,N_10286);
nor U10447 (N_10447,N_10214,N_10390);
or U10448 (N_10448,N_10221,N_10287);
and U10449 (N_10449,N_10346,N_10251);
xnor U10450 (N_10450,N_10235,N_10253);
nand U10451 (N_10451,N_10267,N_10256);
or U10452 (N_10452,N_10234,N_10318);
xnor U10453 (N_10453,N_10313,N_10340);
or U10454 (N_10454,N_10380,N_10349);
and U10455 (N_10455,N_10332,N_10336);
or U10456 (N_10456,N_10307,N_10290);
and U10457 (N_10457,N_10357,N_10338);
or U10458 (N_10458,N_10249,N_10320);
nand U10459 (N_10459,N_10344,N_10277);
or U10460 (N_10460,N_10364,N_10339);
nand U10461 (N_10461,N_10388,N_10304);
nand U10462 (N_10462,N_10225,N_10296);
or U10463 (N_10463,N_10288,N_10255);
or U10464 (N_10464,N_10291,N_10371);
and U10465 (N_10465,N_10311,N_10279);
nor U10466 (N_10466,N_10201,N_10217);
nand U10467 (N_10467,N_10334,N_10220);
xor U10468 (N_10468,N_10331,N_10261);
nor U10469 (N_10469,N_10208,N_10316);
and U10470 (N_10470,N_10387,N_10327);
nand U10471 (N_10471,N_10271,N_10325);
nor U10472 (N_10472,N_10384,N_10385);
or U10473 (N_10473,N_10292,N_10272);
nand U10474 (N_10474,N_10229,N_10289);
and U10475 (N_10475,N_10274,N_10342);
xnor U10476 (N_10476,N_10354,N_10312);
nand U10477 (N_10477,N_10386,N_10211);
or U10478 (N_10478,N_10266,N_10238);
nor U10479 (N_10479,N_10361,N_10227);
or U10480 (N_10480,N_10222,N_10391);
nor U10481 (N_10481,N_10337,N_10308);
nand U10482 (N_10482,N_10381,N_10394);
xor U10483 (N_10483,N_10352,N_10262);
and U10484 (N_10484,N_10345,N_10383);
and U10485 (N_10485,N_10367,N_10343);
xor U10486 (N_10486,N_10273,N_10324);
nor U10487 (N_10487,N_10295,N_10369);
xnor U10488 (N_10488,N_10245,N_10363);
xnor U10489 (N_10489,N_10350,N_10359);
or U10490 (N_10490,N_10379,N_10285);
or U10491 (N_10491,N_10306,N_10218);
nand U10492 (N_10492,N_10333,N_10264);
xor U10493 (N_10493,N_10233,N_10242);
xnor U10494 (N_10494,N_10375,N_10254);
nor U10495 (N_10495,N_10210,N_10335);
and U10496 (N_10496,N_10360,N_10200);
xor U10497 (N_10497,N_10247,N_10223);
nand U10498 (N_10498,N_10309,N_10205);
nand U10499 (N_10499,N_10365,N_10370);
xor U10500 (N_10500,N_10309,N_10258);
xor U10501 (N_10501,N_10383,N_10338);
nor U10502 (N_10502,N_10347,N_10266);
and U10503 (N_10503,N_10231,N_10351);
nor U10504 (N_10504,N_10381,N_10241);
nor U10505 (N_10505,N_10305,N_10307);
nor U10506 (N_10506,N_10242,N_10206);
xor U10507 (N_10507,N_10354,N_10348);
or U10508 (N_10508,N_10344,N_10205);
nor U10509 (N_10509,N_10265,N_10229);
xor U10510 (N_10510,N_10312,N_10329);
or U10511 (N_10511,N_10319,N_10380);
nor U10512 (N_10512,N_10201,N_10280);
nand U10513 (N_10513,N_10389,N_10243);
and U10514 (N_10514,N_10275,N_10214);
or U10515 (N_10515,N_10207,N_10324);
nor U10516 (N_10516,N_10372,N_10229);
and U10517 (N_10517,N_10227,N_10251);
nor U10518 (N_10518,N_10277,N_10342);
nor U10519 (N_10519,N_10274,N_10219);
nor U10520 (N_10520,N_10322,N_10388);
and U10521 (N_10521,N_10310,N_10248);
and U10522 (N_10522,N_10223,N_10357);
nor U10523 (N_10523,N_10267,N_10309);
or U10524 (N_10524,N_10333,N_10246);
xor U10525 (N_10525,N_10301,N_10380);
nand U10526 (N_10526,N_10354,N_10329);
and U10527 (N_10527,N_10292,N_10363);
xor U10528 (N_10528,N_10332,N_10394);
nor U10529 (N_10529,N_10331,N_10234);
and U10530 (N_10530,N_10387,N_10248);
nand U10531 (N_10531,N_10238,N_10203);
nor U10532 (N_10532,N_10282,N_10205);
or U10533 (N_10533,N_10218,N_10317);
nand U10534 (N_10534,N_10374,N_10275);
and U10535 (N_10535,N_10329,N_10337);
xnor U10536 (N_10536,N_10219,N_10224);
xor U10537 (N_10537,N_10341,N_10232);
nand U10538 (N_10538,N_10225,N_10351);
xnor U10539 (N_10539,N_10233,N_10349);
nor U10540 (N_10540,N_10342,N_10293);
nor U10541 (N_10541,N_10328,N_10378);
nand U10542 (N_10542,N_10332,N_10360);
or U10543 (N_10543,N_10330,N_10380);
xor U10544 (N_10544,N_10213,N_10224);
xnor U10545 (N_10545,N_10347,N_10249);
nand U10546 (N_10546,N_10342,N_10340);
or U10547 (N_10547,N_10216,N_10316);
nor U10548 (N_10548,N_10365,N_10279);
xor U10549 (N_10549,N_10397,N_10234);
nor U10550 (N_10550,N_10301,N_10320);
nand U10551 (N_10551,N_10295,N_10357);
nor U10552 (N_10552,N_10395,N_10248);
nor U10553 (N_10553,N_10393,N_10213);
nor U10554 (N_10554,N_10312,N_10303);
or U10555 (N_10555,N_10306,N_10274);
xor U10556 (N_10556,N_10372,N_10309);
or U10557 (N_10557,N_10318,N_10375);
nor U10558 (N_10558,N_10247,N_10256);
nor U10559 (N_10559,N_10378,N_10332);
and U10560 (N_10560,N_10265,N_10207);
xor U10561 (N_10561,N_10317,N_10388);
or U10562 (N_10562,N_10347,N_10203);
xnor U10563 (N_10563,N_10399,N_10266);
and U10564 (N_10564,N_10234,N_10360);
and U10565 (N_10565,N_10340,N_10215);
nand U10566 (N_10566,N_10360,N_10216);
nand U10567 (N_10567,N_10359,N_10340);
xnor U10568 (N_10568,N_10368,N_10254);
xnor U10569 (N_10569,N_10220,N_10286);
or U10570 (N_10570,N_10274,N_10278);
or U10571 (N_10571,N_10268,N_10316);
or U10572 (N_10572,N_10272,N_10350);
nor U10573 (N_10573,N_10256,N_10223);
nand U10574 (N_10574,N_10349,N_10368);
or U10575 (N_10575,N_10296,N_10281);
and U10576 (N_10576,N_10291,N_10243);
nor U10577 (N_10577,N_10344,N_10202);
or U10578 (N_10578,N_10367,N_10369);
xor U10579 (N_10579,N_10379,N_10289);
or U10580 (N_10580,N_10332,N_10269);
nor U10581 (N_10581,N_10395,N_10380);
nor U10582 (N_10582,N_10331,N_10278);
xnor U10583 (N_10583,N_10233,N_10232);
or U10584 (N_10584,N_10373,N_10218);
nand U10585 (N_10585,N_10221,N_10283);
or U10586 (N_10586,N_10228,N_10375);
xnor U10587 (N_10587,N_10266,N_10201);
nor U10588 (N_10588,N_10345,N_10200);
xnor U10589 (N_10589,N_10297,N_10335);
nand U10590 (N_10590,N_10328,N_10297);
xnor U10591 (N_10591,N_10324,N_10300);
nand U10592 (N_10592,N_10222,N_10277);
xnor U10593 (N_10593,N_10374,N_10350);
nand U10594 (N_10594,N_10320,N_10242);
or U10595 (N_10595,N_10245,N_10235);
or U10596 (N_10596,N_10203,N_10349);
nand U10597 (N_10597,N_10324,N_10377);
and U10598 (N_10598,N_10268,N_10208);
and U10599 (N_10599,N_10234,N_10265);
xor U10600 (N_10600,N_10554,N_10440);
or U10601 (N_10601,N_10536,N_10566);
and U10602 (N_10602,N_10413,N_10533);
xnor U10603 (N_10603,N_10591,N_10436);
and U10604 (N_10604,N_10580,N_10581);
and U10605 (N_10605,N_10483,N_10521);
and U10606 (N_10606,N_10499,N_10504);
or U10607 (N_10607,N_10529,N_10433);
nand U10608 (N_10608,N_10564,N_10401);
or U10609 (N_10609,N_10492,N_10469);
xor U10610 (N_10610,N_10437,N_10471);
and U10611 (N_10611,N_10478,N_10479);
xor U10612 (N_10612,N_10505,N_10474);
nor U10613 (N_10613,N_10527,N_10491);
nand U10614 (N_10614,N_10528,N_10510);
nand U10615 (N_10615,N_10501,N_10463);
xnor U10616 (N_10616,N_10584,N_10578);
and U10617 (N_10617,N_10530,N_10526);
xor U10618 (N_10618,N_10473,N_10408);
nor U10619 (N_10619,N_10496,N_10549);
xnor U10620 (N_10620,N_10590,N_10435);
nor U10621 (N_10621,N_10572,N_10518);
xnor U10622 (N_10622,N_10404,N_10439);
or U10623 (N_10623,N_10438,N_10459);
xnor U10624 (N_10624,N_10506,N_10561);
nand U10625 (N_10625,N_10486,N_10557);
or U10626 (N_10626,N_10507,N_10434);
xnor U10627 (N_10627,N_10538,N_10555);
and U10628 (N_10628,N_10456,N_10570);
nand U10629 (N_10629,N_10500,N_10422);
or U10630 (N_10630,N_10583,N_10517);
xnor U10631 (N_10631,N_10567,N_10443);
or U10632 (N_10632,N_10520,N_10490);
xor U10633 (N_10633,N_10573,N_10462);
or U10634 (N_10634,N_10481,N_10512);
xnor U10635 (N_10635,N_10419,N_10544);
nor U10636 (N_10636,N_10455,N_10460);
nand U10637 (N_10637,N_10508,N_10524);
nor U10638 (N_10638,N_10523,N_10420);
nor U10639 (N_10639,N_10493,N_10596);
or U10640 (N_10640,N_10464,N_10574);
xnor U10641 (N_10641,N_10597,N_10579);
nor U10642 (N_10642,N_10489,N_10402);
xor U10643 (N_10643,N_10430,N_10513);
nand U10644 (N_10644,N_10535,N_10563);
nand U10645 (N_10645,N_10539,N_10550);
xnor U10646 (N_10646,N_10426,N_10458);
and U10647 (N_10647,N_10553,N_10467);
nand U10648 (N_10648,N_10577,N_10444);
nor U10649 (N_10649,N_10448,N_10559);
and U10650 (N_10650,N_10587,N_10470);
nor U10651 (N_10651,N_10441,N_10411);
nand U10652 (N_10652,N_10405,N_10586);
and U10653 (N_10653,N_10475,N_10495);
xnor U10654 (N_10654,N_10525,N_10595);
and U10655 (N_10655,N_10445,N_10542);
and U10656 (N_10656,N_10466,N_10497);
nand U10657 (N_10657,N_10498,N_10477);
or U10658 (N_10658,N_10424,N_10537);
nand U10659 (N_10659,N_10502,N_10418);
nand U10660 (N_10660,N_10482,N_10427);
and U10661 (N_10661,N_10476,N_10576);
or U10662 (N_10662,N_10494,N_10598);
nand U10663 (N_10663,N_10594,N_10589);
nor U10664 (N_10664,N_10565,N_10568);
and U10665 (N_10665,N_10406,N_10534);
nand U10666 (N_10666,N_10472,N_10514);
and U10667 (N_10667,N_10531,N_10503);
nor U10668 (N_10668,N_10516,N_10425);
nor U10669 (N_10669,N_10423,N_10541);
nor U10670 (N_10670,N_10546,N_10453);
nand U10671 (N_10671,N_10571,N_10540);
xor U10672 (N_10672,N_10551,N_10519);
nor U10673 (N_10673,N_10582,N_10522);
and U10674 (N_10674,N_10403,N_10407);
nand U10675 (N_10675,N_10480,N_10446);
and U10676 (N_10676,N_10543,N_10558);
nand U10677 (N_10677,N_10592,N_10447);
xor U10678 (N_10678,N_10585,N_10556);
nor U10679 (N_10679,N_10416,N_10452);
nor U10680 (N_10680,N_10552,N_10417);
and U10681 (N_10681,N_10485,N_10431);
xnor U10682 (N_10682,N_10515,N_10509);
and U10683 (N_10683,N_10412,N_10547);
or U10684 (N_10684,N_10599,N_10429);
and U10685 (N_10685,N_10465,N_10450);
nor U10686 (N_10686,N_10457,N_10442);
and U10687 (N_10687,N_10545,N_10400);
and U10688 (N_10688,N_10560,N_10409);
and U10689 (N_10689,N_10415,N_10532);
nand U10690 (N_10690,N_10575,N_10593);
nand U10691 (N_10691,N_10461,N_10488);
or U10692 (N_10692,N_10410,N_10562);
nand U10693 (N_10693,N_10569,N_10421);
and U10694 (N_10694,N_10487,N_10588);
nor U10695 (N_10695,N_10451,N_10511);
or U10696 (N_10696,N_10414,N_10432);
nand U10697 (N_10697,N_10548,N_10428);
and U10698 (N_10698,N_10484,N_10468);
nand U10699 (N_10699,N_10454,N_10449);
nand U10700 (N_10700,N_10475,N_10497);
nor U10701 (N_10701,N_10506,N_10404);
nand U10702 (N_10702,N_10463,N_10439);
nor U10703 (N_10703,N_10523,N_10418);
nor U10704 (N_10704,N_10431,N_10539);
nand U10705 (N_10705,N_10442,N_10409);
nor U10706 (N_10706,N_10515,N_10545);
nor U10707 (N_10707,N_10456,N_10465);
and U10708 (N_10708,N_10489,N_10549);
nor U10709 (N_10709,N_10526,N_10419);
xnor U10710 (N_10710,N_10424,N_10538);
nand U10711 (N_10711,N_10428,N_10599);
or U10712 (N_10712,N_10597,N_10453);
and U10713 (N_10713,N_10542,N_10400);
or U10714 (N_10714,N_10569,N_10575);
xor U10715 (N_10715,N_10511,N_10418);
nor U10716 (N_10716,N_10474,N_10561);
nand U10717 (N_10717,N_10547,N_10467);
and U10718 (N_10718,N_10448,N_10403);
nand U10719 (N_10719,N_10575,N_10549);
xnor U10720 (N_10720,N_10534,N_10487);
or U10721 (N_10721,N_10483,N_10414);
nand U10722 (N_10722,N_10467,N_10444);
xor U10723 (N_10723,N_10419,N_10580);
or U10724 (N_10724,N_10409,N_10472);
and U10725 (N_10725,N_10451,N_10489);
nand U10726 (N_10726,N_10582,N_10560);
xnor U10727 (N_10727,N_10480,N_10488);
nand U10728 (N_10728,N_10432,N_10508);
or U10729 (N_10729,N_10564,N_10421);
nand U10730 (N_10730,N_10564,N_10496);
and U10731 (N_10731,N_10495,N_10431);
or U10732 (N_10732,N_10509,N_10572);
nand U10733 (N_10733,N_10464,N_10503);
xor U10734 (N_10734,N_10422,N_10438);
nand U10735 (N_10735,N_10482,N_10464);
xor U10736 (N_10736,N_10436,N_10494);
xnor U10737 (N_10737,N_10519,N_10486);
nor U10738 (N_10738,N_10591,N_10519);
nand U10739 (N_10739,N_10467,N_10560);
and U10740 (N_10740,N_10490,N_10480);
xor U10741 (N_10741,N_10582,N_10524);
nand U10742 (N_10742,N_10504,N_10435);
nor U10743 (N_10743,N_10489,N_10514);
or U10744 (N_10744,N_10486,N_10417);
xnor U10745 (N_10745,N_10415,N_10512);
and U10746 (N_10746,N_10588,N_10576);
and U10747 (N_10747,N_10479,N_10512);
nor U10748 (N_10748,N_10540,N_10449);
and U10749 (N_10749,N_10488,N_10402);
nand U10750 (N_10750,N_10544,N_10560);
xnor U10751 (N_10751,N_10589,N_10548);
nor U10752 (N_10752,N_10518,N_10489);
or U10753 (N_10753,N_10437,N_10545);
nor U10754 (N_10754,N_10502,N_10480);
or U10755 (N_10755,N_10443,N_10432);
nor U10756 (N_10756,N_10498,N_10424);
and U10757 (N_10757,N_10480,N_10558);
nand U10758 (N_10758,N_10518,N_10536);
or U10759 (N_10759,N_10585,N_10530);
xnor U10760 (N_10760,N_10444,N_10588);
and U10761 (N_10761,N_10529,N_10459);
or U10762 (N_10762,N_10569,N_10560);
nor U10763 (N_10763,N_10492,N_10512);
nor U10764 (N_10764,N_10531,N_10576);
xor U10765 (N_10765,N_10590,N_10525);
xnor U10766 (N_10766,N_10407,N_10576);
nor U10767 (N_10767,N_10588,N_10566);
and U10768 (N_10768,N_10472,N_10450);
and U10769 (N_10769,N_10569,N_10514);
and U10770 (N_10770,N_10430,N_10509);
nor U10771 (N_10771,N_10457,N_10448);
or U10772 (N_10772,N_10459,N_10518);
xor U10773 (N_10773,N_10417,N_10419);
xor U10774 (N_10774,N_10459,N_10579);
or U10775 (N_10775,N_10507,N_10447);
xor U10776 (N_10776,N_10563,N_10482);
nor U10777 (N_10777,N_10573,N_10590);
nand U10778 (N_10778,N_10583,N_10423);
xnor U10779 (N_10779,N_10598,N_10492);
nand U10780 (N_10780,N_10487,N_10518);
and U10781 (N_10781,N_10439,N_10511);
nand U10782 (N_10782,N_10441,N_10479);
nor U10783 (N_10783,N_10584,N_10507);
xor U10784 (N_10784,N_10486,N_10527);
or U10785 (N_10785,N_10405,N_10537);
and U10786 (N_10786,N_10578,N_10525);
nor U10787 (N_10787,N_10407,N_10400);
or U10788 (N_10788,N_10400,N_10509);
xor U10789 (N_10789,N_10584,N_10597);
nand U10790 (N_10790,N_10465,N_10593);
nand U10791 (N_10791,N_10409,N_10406);
xor U10792 (N_10792,N_10501,N_10573);
or U10793 (N_10793,N_10584,N_10598);
nor U10794 (N_10794,N_10594,N_10456);
or U10795 (N_10795,N_10476,N_10511);
xnor U10796 (N_10796,N_10519,N_10465);
xnor U10797 (N_10797,N_10442,N_10490);
xnor U10798 (N_10798,N_10555,N_10456);
nand U10799 (N_10799,N_10593,N_10524);
xor U10800 (N_10800,N_10748,N_10687);
and U10801 (N_10801,N_10602,N_10605);
or U10802 (N_10802,N_10785,N_10766);
nand U10803 (N_10803,N_10782,N_10610);
nor U10804 (N_10804,N_10781,N_10790);
nand U10805 (N_10805,N_10756,N_10778);
nor U10806 (N_10806,N_10753,N_10788);
and U10807 (N_10807,N_10603,N_10773);
nor U10808 (N_10808,N_10675,N_10656);
and U10809 (N_10809,N_10682,N_10620);
nand U10810 (N_10810,N_10600,N_10689);
xnor U10811 (N_10811,N_10733,N_10613);
nand U10812 (N_10812,N_10601,N_10729);
or U10813 (N_10813,N_10783,N_10767);
and U10814 (N_10814,N_10750,N_10721);
nand U10815 (N_10815,N_10796,N_10726);
nand U10816 (N_10816,N_10761,N_10639);
and U10817 (N_10817,N_10683,N_10702);
nor U10818 (N_10818,N_10752,N_10664);
and U10819 (N_10819,N_10751,N_10673);
nand U10820 (N_10820,N_10650,N_10644);
nor U10821 (N_10821,N_10607,N_10695);
and U10822 (N_10822,N_10626,N_10777);
nand U10823 (N_10823,N_10795,N_10698);
or U10824 (N_10824,N_10658,N_10771);
and U10825 (N_10825,N_10638,N_10780);
and U10826 (N_10826,N_10779,N_10701);
xnor U10827 (N_10827,N_10749,N_10668);
nand U10828 (N_10828,N_10671,N_10714);
and U10829 (N_10829,N_10631,N_10764);
nand U10830 (N_10830,N_10716,N_10768);
xor U10831 (N_10831,N_10792,N_10743);
nor U10832 (N_10832,N_10700,N_10608);
or U10833 (N_10833,N_10623,N_10617);
and U10834 (N_10834,N_10630,N_10797);
nor U10835 (N_10835,N_10635,N_10770);
xnor U10836 (N_10836,N_10677,N_10674);
or U10837 (N_10837,N_10666,N_10662);
nand U10838 (N_10838,N_10755,N_10713);
xor U10839 (N_10839,N_10765,N_10722);
or U10840 (N_10840,N_10669,N_10648);
and U10841 (N_10841,N_10632,N_10615);
nand U10842 (N_10842,N_10734,N_10667);
xor U10843 (N_10843,N_10794,N_10684);
xnor U10844 (N_10844,N_10704,N_10724);
and U10845 (N_10845,N_10690,N_10691);
and U10846 (N_10846,N_10612,N_10637);
nand U10847 (N_10847,N_10665,N_10636);
or U10848 (N_10848,N_10661,N_10705);
nor U10849 (N_10849,N_10679,N_10622);
and U10850 (N_10850,N_10652,N_10659);
and U10851 (N_10851,N_10654,N_10728);
nor U10852 (N_10852,N_10611,N_10757);
xnor U10853 (N_10853,N_10625,N_10686);
nor U10854 (N_10854,N_10774,N_10742);
xnor U10855 (N_10855,N_10629,N_10694);
nand U10856 (N_10856,N_10744,N_10619);
or U10857 (N_10857,N_10719,N_10709);
or U10858 (N_10858,N_10681,N_10618);
nand U10859 (N_10859,N_10799,N_10769);
nor U10860 (N_10860,N_10712,N_10653);
or U10861 (N_10861,N_10786,N_10649);
or U10862 (N_10862,N_10640,N_10663);
and U10863 (N_10863,N_10655,N_10717);
xnor U10864 (N_10864,N_10696,N_10707);
xnor U10865 (N_10865,N_10688,N_10747);
nand U10866 (N_10866,N_10609,N_10685);
nand U10867 (N_10867,N_10754,N_10646);
and U10868 (N_10868,N_10604,N_10736);
xnor U10869 (N_10869,N_10740,N_10624);
nor U10870 (N_10870,N_10730,N_10738);
and U10871 (N_10871,N_10708,N_10657);
nand U10872 (N_10872,N_10776,N_10634);
and U10873 (N_10873,N_10718,N_10614);
and U10874 (N_10874,N_10737,N_10676);
nor U10875 (N_10875,N_10670,N_10772);
and U10876 (N_10876,N_10720,N_10645);
xor U10877 (N_10877,N_10787,N_10745);
or U10878 (N_10878,N_10746,N_10633);
xnor U10879 (N_10879,N_10741,N_10660);
and U10880 (N_10880,N_10735,N_10760);
nand U10881 (N_10881,N_10703,N_10731);
nand U10882 (N_10882,N_10798,N_10789);
or U10883 (N_10883,N_10642,N_10711);
or U10884 (N_10884,N_10759,N_10692);
and U10885 (N_10885,N_10641,N_10758);
or U10886 (N_10886,N_10627,N_10628);
nand U10887 (N_10887,N_10616,N_10775);
xnor U10888 (N_10888,N_10732,N_10643);
and U10889 (N_10889,N_10706,N_10791);
xnor U10890 (N_10890,N_10710,N_10727);
or U10891 (N_10891,N_10784,N_10693);
nor U10892 (N_10892,N_10793,N_10647);
and U10893 (N_10893,N_10621,N_10680);
nand U10894 (N_10894,N_10672,N_10678);
xnor U10895 (N_10895,N_10651,N_10762);
and U10896 (N_10896,N_10697,N_10606);
nor U10897 (N_10897,N_10725,N_10763);
nor U10898 (N_10898,N_10723,N_10715);
or U10899 (N_10899,N_10739,N_10699);
nand U10900 (N_10900,N_10786,N_10799);
or U10901 (N_10901,N_10612,N_10727);
and U10902 (N_10902,N_10695,N_10621);
nand U10903 (N_10903,N_10759,N_10661);
nand U10904 (N_10904,N_10716,N_10747);
and U10905 (N_10905,N_10799,N_10728);
nor U10906 (N_10906,N_10726,N_10607);
nand U10907 (N_10907,N_10613,N_10701);
or U10908 (N_10908,N_10664,N_10728);
xor U10909 (N_10909,N_10611,N_10628);
or U10910 (N_10910,N_10622,N_10793);
or U10911 (N_10911,N_10668,N_10717);
and U10912 (N_10912,N_10736,N_10798);
and U10913 (N_10913,N_10667,N_10753);
and U10914 (N_10914,N_10651,N_10748);
or U10915 (N_10915,N_10698,N_10725);
nor U10916 (N_10916,N_10769,N_10703);
nand U10917 (N_10917,N_10634,N_10658);
nor U10918 (N_10918,N_10798,N_10656);
xnor U10919 (N_10919,N_10783,N_10744);
and U10920 (N_10920,N_10689,N_10634);
nand U10921 (N_10921,N_10791,N_10741);
nand U10922 (N_10922,N_10792,N_10796);
and U10923 (N_10923,N_10700,N_10681);
or U10924 (N_10924,N_10715,N_10781);
and U10925 (N_10925,N_10762,N_10684);
xnor U10926 (N_10926,N_10637,N_10695);
nor U10927 (N_10927,N_10602,N_10633);
nor U10928 (N_10928,N_10761,N_10723);
xnor U10929 (N_10929,N_10728,N_10777);
and U10930 (N_10930,N_10632,N_10742);
xor U10931 (N_10931,N_10722,N_10705);
xor U10932 (N_10932,N_10731,N_10737);
nand U10933 (N_10933,N_10666,N_10703);
or U10934 (N_10934,N_10663,N_10791);
xnor U10935 (N_10935,N_10798,N_10672);
nor U10936 (N_10936,N_10688,N_10643);
and U10937 (N_10937,N_10640,N_10679);
or U10938 (N_10938,N_10608,N_10678);
nor U10939 (N_10939,N_10748,N_10774);
and U10940 (N_10940,N_10755,N_10613);
nor U10941 (N_10941,N_10772,N_10755);
xnor U10942 (N_10942,N_10692,N_10777);
or U10943 (N_10943,N_10741,N_10748);
xor U10944 (N_10944,N_10756,N_10770);
nand U10945 (N_10945,N_10630,N_10781);
nand U10946 (N_10946,N_10728,N_10782);
or U10947 (N_10947,N_10750,N_10637);
nand U10948 (N_10948,N_10773,N_10710);
nor U10949 (N_10949,N_10617,N_10619);
xnor U10950 (N_10950,N_10700,N_10621);
or U10951 (N_10951,N_10749,N_10650);
xnor U10952 (N_10952,N_10720,N_10727);
xor U10953 (N_10953,N_10744,N_10704);
and U10954 (N_10954,N_10711,N_10659);
nor U10955 (N_10955,N_10795,N_10790);
nand U10956 (N_10956,N_10638,N_10722);
nor U10957 (N_10957,N_10794,N_10752);
nand U10958 (N_10958,N_10759,N_10678);
and U10959 (N_10959,N_10642,N_10668);
and U10960 (N_10960,N_10797,N_10728);
nand U10961 (N_10961,N_10787,N_10671);
or U10962 (N_10962,N_10721,N_10710);
nand U10963 (N_10963,N_10675,N_10683);
nor U10964 (N_10964,N_10788,N_10791);
xnor U10965 (N_10965,N_10784,N_10798);
or U10966 (N_10966,N_10711,N_10741);
and U10967 (N_10967,N_10775,N_10637);
and U10968 (N_10968,N_10784,N_10679);
or U10969 (N_10969,N_10799,N_10640);
nand U10970 (N_10970,N_10784,N_10770);
or U10971 (N_10971,N_10613,N_10637);
nor U10972 (N_10972,N_10721,N_10622);
and U10973 (N_10973,N_10634,N_10704);
xor U10974 (N_10974,N_10736,N_10608);
or U10975 (N_10975,N_10724,N_10631);
xnor U10976 (N_10976,N_10656,N_10621);
xnor U10977 (N_10977,N_10646,N_10741);
nand U10978 (N_10978,N_10686,N_10638);
and U10979 (N_10979,N_10655,N_10612);
xor U10980 (N_10980,N_10686,N_10609);
nor U10981 (N_10981,N_10745,N_10672);
nor U10982 (N_10982,N_10762,N_10645);
or U10983 (N_10983,N_10643,N_10703);
and U10984 (N_10984,N_10631,N_10704);
and U10985 (N_10985,N_10763,N_10757);
and U10986 (N_10986,N_10633,N_10783);
xor U10987 (N_10987,N_10617,N_10680);
or U10988 (N_10988,N_10671,N_10640);
xnor U10989 (N_10989,N_10657,N_10707);
nand U10990 (N_10990,N_10655,N_10700);
and U10991 (N_10991,N_10667,N_10756);
nor U10992 (N_10992,N_10638,N_10684);
nand U10993 (N_10993,N_10725,N_10764);
nor U10994 (N_10994,N_10667,N_10759);
nand U10995 (N_10995,N_10716,N_10683);
or U10996 (N_10996,N_10660,N_10654);
nor U10997 (N_10997,N_10676,N_10714);
nor U10998 (N_10998,N_10639,N_10726);
xnor U10999 (N_10999,N_10715,N_10788);
or U11000 (N_11000,N_10997,N_10873);
and U11001 (N_11001,N_10884,N_10810);
and U11002 (N_11002,N_10977,N_10864);
nor U11003 (N_11003,N_10833,N_10968);
and U11004 (N_11004,N_10894,N_10922);
or U11005 (N_11005,N_10842,N_10931);
nor U11006 (N_11006,N_10960,N_10966);
nor U11007 (N_11007,N_10903,N_10988);
nand U11008 (N_11008,N_10885,N_10902);
nand U11009 (N_11009,N_10908,N_10984);
xnor U11010 (N_11010,N_10949,N_10878);
or U11011 (N_11011,N_10897,N_10886);
nand U11012 (N_11012,N_10920,N_10816);
nor U11013 (N_11013,N_10987,N_10856);
nor U11014 (N_11014,N_10893,N_10800);
and U11015 (N_11015,N_10924,N_10803);
or U11016 (N_11016,N_10964,N_10909);
and U11017 (N_11017,N_10995,N_10912);
nand U11018 (N_11018,N_10890,N_10904);
nor U11019 (N_11019,N_10942,N_10828);
xor U11020 (N_11020,N_10906,N_10849);
or U11021 (N_11021,N_10811,N_10944);
or U11022 (N_11022,N_10854,N_10910);
nor U11023 (N_11023,N_10971,N_10870);
and U11024 (N_11024,N_10888,N_10835);
xor U11025 (N_11025,N_10858,N_10972);
and U11026 (N_11026,N_10892,N_10983);
and U11027 (N_11027,N_10999,N_10979);
xor U11028 (N_11028,N_10927,N_10926);
nand U11029 (N_11029,N_10992,N_10941);
nor U11030 (N_11030,N_10895,N_10825);
nand U11031 (N_11031,N_10865,N_10954);
xnor U11032 (N_11032,N_10851,N_10866);
and U11033 (N_11033,N_10883,N_10806);
nor U11034 (N_11034,N_10839,N_10831);
or U11035 (N_11035,N_10932,N_10820);
nor U11036 (N_11036,N_10982,N_10815);
or U11037 (N_11037,N_10925,N_10936);
and U11038 (N_11038,N_10990,N_10808);
nand U11039 (N_11039,N_10996,N_10863);
or U11040 (N_11040,N_10917,N_10834);
xnor U11041 (N_11041,N_10955,N_10846);
or U11042 (N_11042,N_10950,N_10877);
xor U11043 (N_11043,N_10817,N_10953);
and U11044 (N_11044,N_10827,N_10840);
or U11045 (N_11045,N_10847,N_10921);
or U11046 (N_11046,N_10938,N_10887);
nor U11047 (N_11047,N_10930,N_10882);
nand U11048 (N_11048,N_10869,N_10838);
and U11049 (N_11049,N_10812,N_10871);
nand U11050 (N_11050,N_10844,N_10879);
nor U11051 (N_11051,N_10889,N_10937);
nor U11052 (N_11052,N_10829,N_10934);
or U11053 (N_11053,N_10959,N_10807);
and U11054 (N_11054,N_10916,N_10986);
and U11055 (N_11055,N_10980,N_10809);
xnor U11056 (N_11056,N_10928,N_10940);
xor U11057 (N_11057,N_10899,N_10914);
nand U11058 (N_11058,N_10962,N_10985);
and U11059 (N_11059,N_10843,N_10813);
and U11060 (N_11060,N_10989,N_10804);
and U11061 (N_11061,N_10952,N_10969);
nand U11062 (N_11062,N_10961,N_10970);
xnor U11063 (N_11063,N_10876,N_10946);
nor U11064 (N_11064,N_10855,N_10974);
xnor U11065 (N_11065,N_10821,N_10853);
xor U11066 (N_11066,N_10832,N_10905);
or U11067 (N_11067,N_10963,N_10841);
nand U11068 (N_11068,N_10896,N_10836);
or U11069 (N_11069,N_10859,N_10907);
or U11070 (N_11070,N_10824,N_10868);
nand U11071 (N_11071,N_10845,N_10900);
nor U11072 (N_11072,N_10850,N_10981);
nand U11073 (N_11073,N_10978,N_10956);
nor U11074 (N_11074,N_10958,N_10875);
or U11075 (N_11075,N_10998,N_10814);
xnor U11076 (N_11076,N_10881,N_10862);
or U11077 (N_11077,N_10872,N_10852);
nor U11078 (N_11078,N_10973,N_10918);
and U11079 (N_11079,N_10947,N_10919);
and U11080 (N_11080,N_10993,N_10822);
or U11081 (N_11081,N_10965,N_10913);
xnor U11082 (N_11082,N_10975,N_10861);
xnor U11083 (N_11083,N_10911,N_10933);
nor U11084 (N_11084,N_10915,N_10819);
xnor U11085 (N_11085,N_10976,N_10867);
nand U11086 (N_11086,N_10805,N_10874);
or U11087 (N_11087,N_10860,N_10857);
nor U11088 (N_11088,N_10935,N_10802);
nor U11089 (N_11089,N_10898,N_10939);
xnor U11090 (N_11090,N_10891,N_10994);
nand U11091 (N_11091,N_10830,N_10880);
nor U11092 (N_11092,N_10848,N_10945);
nand U11093 (N_11093,N_10837,N_10826);
nand U11094 (N_11094,N_10801,N_10929);
nor U11095 (N_11095,N_10818,N_10943);
nand U11096 (N_11096,N_10923,N_10823);
or U11097 (N_11097,N_10951,N_10957);
xnor U11098 (N_11098,N_10901,N_10967);
and U11099 (N_11099,N_10948,N_10991);
nor U11100 (N_11100,N_10981,N_10949);
nand U11101 (N_11101,N_10998,N_10838);
and U11102 (N_11102,N_10963,N_10943);
xor U11103 (N_11103,N_10838,N_10976);
or U11104 (N_11104,N_10905,N_10873);
nand U11105 (N_11105,N_10804,N_10806);
xor U11106 (N_11106,N_10992,N_10912);
nor U11107 (N_11107,N_10937,N_10857);
nor U11108 (N_11108,N_10839,N_10871);
nor U11109 (N_11109,N_10858,N_10951);
or U11110 (N_11110,N_10816,N_10893);
nand U11111 (N_11111,N_10895,N_10844);
and U11112 (N_11112,N_10953,N_10972);
or U11113 (N_11113,N_10941,N_10801);
nor U11114 (N_11114,N_10943,N_10867);
nand U11115 (N_11115,N_10816,N_10855);
xnor U11116 (N_11116,N_10979,N_10951);
nand U11117 (N_11117,N_10931,N_10818);
nand U11118 (N_11118,N_10935,N_10854);
or U11119 (N_11119,N_10896,N_10865);
and U11120 (N_11120,N_10973,N_10927);
and U11121 (N_11121,N_10919,N_10833);
nand U11122 (N_11122,N_10938,N_10850);
nand U11123 (N_11123,N_10916,N_10801);
xnor U11124 (N_11124,N_10922,N_10877);
nand U11125 (N_11125,N_10846,N_10937);
nor U11126 (N_11126,N_10940,N_10974);
xor U11127 (N_11127,N_10867,N_10941);
xor U11128 (N_11128,N_10830,N_10971);
nor U11129 (N_11129,N_10998,N_10960);
xor U11130 (N_11130,N_10908,N_10811);
and U11131 (N_11131,N_10940,N_10902);
and U11132 (N_11132,N_10919,N_10898);
xnor U11133 (N_11133,N_10969,N_10912);
nor U11134 (N_11134,N_10954,N_10803);
nand U11135 (N_11135,N_10996,N_10895);
nand U11136 (N_11136,N_10819,N_10930);
nand U11137 (N_11137,N_10803,N_10943);
and U11138 (N_11138,N_10979,N_10983);
nand U11139 (N_11139,N_10923,N_10891);
nor U11140 (N_11140,N_10867,N_10869);
and U11141 (N_11141,N_10922,N_10986);
nor U11142 (N_11142,N_10882,N_10909);
nand U11143 (N_11143,N_10863,N_10969);
xor U11144 (N_11144,N_10858,N_10806);
and U11145 (N_11145,N_10897,N_10876);
nor U11146 (N_11146,N_10941,N_10836);
nand U11147 (N_11147,N_10872,N_10876);
nor U11148 (N_11148,N_10909,N_10859);
nor U11149 (N_11149,N_10948,N_10812);
nand U11150 (N_11150,N_10821,N_10989);
xnor U11151 (N_11151,N_10976,N_10989);
nor U11152 (N_11152,N_10884,N_10909);
nor U11153 (N_11153,N_10888,N_10979);
nand U11154 (N_11154,N_10832,N_10897);
and U11155 (N_11155,N_10831,N_10851);
nand U11156 (N_11156,N_10904,N_10801);
xnor U11157 (N_11157,N_10886,N_10998);
and U11158 (N_11158,N_10864,N_10899);
or U11159 (N_11159,N_10810,N_10893);
xor U11160 (N_11160,N_10852,N_10842);
nor U11161 (N_11161,N_10823,N_10810);
nand U11162 (N_11162,N_10859,N_10992);
and U11163 (N_11163,N_10818,N_10808);
xnor U11164 (N_11164,N_10995,N_10936);
xor U11165 (N_11165,N_10965,N_10802);
nand U11166 (N_11166,N_10902,N_10873);
xnor U11167 (N_11167,N_10822,N_10929);
xnor U11168 (N_11168,N_10997,N_10811);
and U11169 (N_11169,N_10854,N_10876);
or U11170 (N_11170,N_10885,N_10828);
nor U11171 (N_11171,N_10863,N_10864);
and U11172 (N_11172,N_10814,N_10966);
and U11173 (N_11173,N_10823,N_10975);
xnor U11174 (N_11174,N_10929,N_10903);
or U11175 (N_11175,N_10913,N_10932);
nor U11176 (N_11176,N_10826,N_10917);
xor U11177 (N_11177,N_10949,N_10947);
or U11178 (N_11178,N_10808,N_10989);
nor U11179 (N_11179,N_10916,N_10914);
nand U11180 (N_11180,N_10878,N_10874);
xor U11181 (N_11181,N_10953,N_10997);
nand U11182 (N_11182,N_10872,N_10809);
nor U11183 (N_11183,N_10889,N_10910);
nor U11184 (N_11184,N_10895,N_10976);
xor U11185 (N_11185,N_10920,N_10985);
xnor U11186 (N_11186,N_10902,N_10802);
nand U11187 (N_11187,N_10808,N_10967);
xnor U11188 (N_11188,N_10894,N_10995);
or U11189 (N_11189,N_10932,N_10919);
nand U11190 (N_11190,N_10905,N_10868);
and U11191 (N_11191,N_10925,N_10954);
or U11192 (N_11192,N_10993,N_10969);
or U11193 (N_11193,N_10981,N_10910);
and U11194 (N_11194,N_10806,N_10980);
nor U11195 (N_11195,N_10807,N_10924);
nand U11196 (N_11196,N_10832,N_10991);
nand U11197 (N_11197,N_10841,N_10927);
nor U11198 (N_11198,N_10958,N_10951);
nor U11199 (N_11199,N_10906,N_10871);
xor U11200 (N_11200,N_11176,N_11167);
nor U11201 (N_11201,N_11095,N_11102);
xnor U11202 (N_11202,N_11074,N_11122);
nor U11203 (N_11203,N_11025,N_11129);
and U11204 (N_11204,N_11022,N_11046);
nor U11205 (N_11205,N_11106,N_11173);
and U11206 (N_11206,N_11030,N_11049);
nand U11207 (N_11207,N_11054,N_11190);
nand U11208 (N_11208,N_11153,N_11137);
and U11209 (N_11209,N_11187,N_11015);
or U11210 (N_11210,N_11115,N_11105);
xnor U11211 (N_11211,N_11011,N_11142);
nor U11212 (N_11212,N_11083,N_11019);
nor U11213 (N_11213,N_11059,N_11112);
nor U11214 (N_11214,N_11077,N_11024);
xor U11215 (N_11215,N_11098,N_11004);
xor U11216 (N_11216,N_11108,N_11027);
or U11217 (N_11217,N_11007,N_11041);
nor U11218 (N_11218,N_11001,N_11010);
nand U11219 (N_11219,N_11076,N_11036);
xor U11220 (N_11220,N_11166,N_11191);
nand U11221 (N_11221,N_11082,N_11174);
and U11222 (N_11222,N_11103,N_11026);
or U11223 (N_11223,N_11151,N_11037);
and U11224 (N_11224,N_11148,N_11075);
xor U11225 (N_11225,N_11078,N_11107);
nand U11226 (N_11226,N_11080,N_11143);
nor U11227 (N_11227,N_11058,N_11051);
xor U11228 (N_11228,N_11017,N_11168);
xnor U11229 (N_11229,N_11152,N_11031);
or U11230 (N_11230,N_11180,N_11057);
and U11231 (N_11231,N_11123,N_11116);
nand U11232 (N_11232,N_11060,N_11088);
and U11233 (N_11233,N_11045,N_11192);
or U11234 (N_11234,N_11120,N_11197);
nand U11235 (N_11235,N_11009,N_11100);
nand U11236 (N_11236,N_11016,N_11195);
xor U11237 (N_11237,N_11172,N_11006);
and U11238 (N_11238,N_11068,N_11136);
nand U11239 (N_11239,N_11056,N_11003);
xnor U11240 (N_11240,N_11144,N_11134);
xor U11241 (N_11241,N_11065,N_11101);
xor U11242 (N_11242,N_11033,N_11114);
nand U11243 (N_11243,N_11038,N_11061);
nor U11244 (N_11244,N_11028,N_11126);
or U11245 (N_11245,N_11050,N_11000);
or U11246 (N_11246,N_11085,N_11042);
nand U11247 (N_11247,N_11196,N_11072);
nand U11248 (N_11248,N_11092,N_11169);
and U11249 (N_11249,N_11145,N_11023);
xnor U11250 (N_11250,N_11018,N_11160);
nand U11251 (N_11251,N_11013,N_11128);
and U11252 (N_11252,N_11014,N_11052);
xor U11253 (N_11253,N_11035,N_11165);
xor U11254 (N_11254,N_11081,N_11139);
or U11255 (N_11255,N_11021,N_11109);
nor U11256 (N_11256,N_11183,N_11154);
xnor U11257 (N_11257,N_11008,N_11161);
nor U11258 (N_11258,N_11094,N_11198);
nand U11259 (N_11259,N_11177,N_11002);
nand U11260 (N_11260,N_11178,N_11199);
xor U11261 (N_11261,N_11097,N_11133);
nand U11262 (N_11262,N_11067,N_11063);
xnor U11263 (N_11263,N_11181,N_11194);
and U11264 (N_11264,N_11053,N_11157);
or U11265 (N_11265,N_11069,N_11182);
or U11266 (N_11266,N_11044,N_11179);
nand U11267 (N_11267,N_11185,N_11090);
or U11268 (N_11268,N_11127,N_11149);
nand U11269 (N_11269,N_11156,N_11189);
or U11270 (N_11270,N_11146,N_11062);
xnor U11271 (N_11271,N_11070,N_11064);
or U11272 (N_11272,N_11073,N_11047);
or U11273 (N_11273,N_11099,N_11093);
and U11274 (N_11274,N_11034,N_11091);
xor U11275 (N_11275,N_11130,N_11117);
nor U11276 (N_11276,N_11096,N_11040);
xor U11277 (N_11277,N_11005,N_11138);
or U11278 (N_11278,N_11079,N_11159);
nor U11279 (N_11279,N_11118,N_11186);
and U11280 (N_11280,N_11131,N_11029);
or U11281 (N_11281,N_11124,N_11104);
nand U11282 (N_11282,N_11039,N_11150);
nor U11283 (N_11283,N_11113,N_11055);
xnor U11284 (N_11284,N_11164,N_11048);
nor U11285 (N_11285,N_11162,N_11089);
nand U11286 (N_11286,N_11066,N_11012);
nand U11287 (N_11287,N_11141,N_11175);
or U11288 (N_11288,N_11121,N_11071);
and U11289 (N_11289,N_11110,N_11125);
nand U11290 (N_11290,N_11163,N_11132);
nand U11291 (N_11291,N_11086,N_11043);
nor U11292 (N_11292,N_11119,N_11140);
nor U11293 (N_11293,N_11147,N_11171);
nor U11294 (N_11294,N_11184,N_11032);
and U11295 (N_11295,N_11087,N_11020);
nor U11296 (N_11296,N_11084,N_11188);
xnor U11297 (N_11297,N_11158,N_11170);
and U11298 (N_11298,N_11111,N_11193);
xor U11299 (N_11299,N_11135,N_11155);
nand U11300 (N_11300,N_11004,N_11176);
nor U11301 (N_11301,N_11180,N_11136);
and U11302 (N_11302,N_11194,N_11077);
xor U11303 (N_11303,N_11027,N_11077);
nor U11304 (N_11304,N_11013,N_11152);
and U11305 (N_11305,N_11092,N_11109);
and U11306 (N_11306,N_11069,N_11144);
nor U11307 (N_11307,N_11189,N_11052);
xor U11308 (N_11308,N_11187,N_11092);
xor U11309 (N_11309,N_11162,N_11141);
xnor U11310 (N_11310,N_11109,N_11152);
or U11311 (N_11311,N_11094,N_11122);
or U11312 (N_11312,N_11071,N_11028);
nand U11313 (N_11313,N_11080,N_11132);
nand U11314 (N_11314,N_11074,N_11052);
nor U11315 (N_11315,N_11026,N_11166);
xnor U11316 (N_11316,N_11146,N_11010);
and U11317 (N_11317,N_11107,N_11191);
nor U11318 (N_11318,N_11071,N_11140);
and U11319 (N_11319,N_11043,N_11064);
xnor U11320 (N_11320,N_11156,N_11108);
nor U11321 (N_11321,N_11131,N_11075);
and U11322 (N_11322,N_11157,N_11064);
nor U11323 (N_11323,N_11010,N_11058);
and U11324 (N_11324,N_11006,N_11113);
xnor U11325 (N_11325,N_11052,N_11163);
and U11326 (N_11326,N_11198,N_11026);
nor U11327 (N_11327,N_11005,N_11091);
or U11328 (N_11328,N_11177,N_11035);
or U11329 (N_11329,N_11198,N_11084);
and U11330 (N_11330,N_11185,N_11048);
and U11331 (N_11331,N_11136,N_11063);
xor U11332 (N_11332,N_11038,N_11041);
nor U11333 (N_11333,N_11186,N_11162);
xnor U11334 (N_11334,N_11007,N_11073);
xnor U11335 (N_11335,N_11025,N_11005);
or U11336 (N_11336,N_11127,N_11059);
nand U11337 (N_11337,N_11054,N_11059);
and U11338 (N_11338,N_11096,N_11058);
or U11339 (N_11339,N_11164,N_11189);
nor U11340 (N_11340,N_11044,N_11005);
and U11341 (N_11341,N_11083,N_11046);
xor U11342 (N_11342,N_11065,N_11123);
nor U11343 (N_11343,N_11002,N_11032);
and U11344 (N_11344,N_11004,N_11045);
xnor U11345 (N_11345,N_11092,N_11002);
nand U11346 (N_11346,N_11083,N_11031);
nor U11347 (N_11347,N_11166,N_11103);
nand U11348 (N_11348,N_11186,N_11071);
xor U11349 (N_11349,N_11037,N_11186);
nand U11350 (N_11350,N_11091,N_11115);
nand U11351 (N_11351,N_11181,N_11038);
nor U11352 (N_11352,N_11183,N_11164);
and U11353 (N_11353,N_11065,N_11194);
xnor U11354 (N_11354,N_11136,N_11012);
and U11355 (N_11355,N_11150,N_11075);
or U11356 (N_11356,N_11127,N_11045);
and U11357 (N_11357,N_11194,N_11021);
nor U11358 (N_11358,N_11072,N_11122);
or U11359 (N_11359,N_11128,N_11071);
nor U11360 (N_11360,N_11188,N_11163);
and U11361 (N_11361,N_11110,N_11107);
nor U11362 (N_11362,N_11094,N_11020);
nor U11363 (N_11363,N_11180,N_11070);
nor U11364 (N_11364,N_11087,N_11004);
xor U11365 (N_11365,N_11165,N_11026);
nor U11366 (N_11366,N_11101,N_11064);
or U11367 (N_11367,N_11195,N_11143);
xnor U11368 (N_11368,N_11155,N_11139);
nor U11369 (N_11369,N_11128,N_11069);
or U11370 (N_11370,N_11193,N_11044);
nand U11371 (N_11371,N_11137,N_11107);
and U11372 (N_11372,N_11129,N_11190);
or U11373 (N_11373,N_11019,N_11114);
or U11374 (N_11374,N_11174,N_11076);
nor U11375 (N_11375,N_11025,N_11093);
or U11376 (N_11376,N_11012,N_11092);
nor U11377 (N_11377,N_11179,N_11080);
nor U11378 (N_11378,N_11119,N_11087);
or U11379 (N_11379,N_11062,N_11021);
xor U11380 (N_11380,N_11073,N_11012);
xor U11381 (N_11381,N_11029,N_11004);
or U11382 (N_11382,N_11049,N_11199);
xnor U11383 (N_11383,N_11074,N_11036);
nor U11384 (N_11384,N_11065,N_11071);
and U11385 (N_11385,N_11151,N_11158);
or U11386 (N_11386,N_11001,N_11134);
and U11387 (N_11387,N_11026,N_11050);
nor U11388 (N_11388,N_11128,N_11054);
nand U11389 (N_11389,N_11181,N_11144);
or U11390 (N_11390,N_11021,N_11026);
xor U11391 (N_11391,N_11198,N_11146);
nor U11392 (N_11392,N_11038,N_11010);
nand U11393 (N_11393,N_11040,N_11095);
nand U11394 (N_11394,N_11189,N_11047);
or U11395 (N_11395,N_11076,N_11010);
nor U11396 (N_11396,N_11065,N_11118);
nor U11397 (N_11397,N_11003,N_11068);
and U11398 (N_11398,N_11045,N_11072);
nand U11399 (N_11399,N_11156,N_11021);
xor U11400 (N_11400,N_11221,N_11364);
nand U11401 (N_11401,N_11272,N_11291);
nor U11402 (N_11402,N_11375,N_11347);
and U11403 (N_11403,N_11337,N_11379);
nand U11404 (N_11404,N_11226,N_11385);
xnor U11405 (N_11405,N_11312,N_11328);
and U11406 (N_11406,N_11296,N_11362);
nand U11407 (N_11407,N_11209,N_11394);
or U11408 (N_11408,N_11270,N_11281);
and U11409 (N_11409,N_11253,N_11338);
or U11410 (N_11410,N_11356,N_11223);
xnor U11411 (N_11411,N_11369,N_11207);
xnor U11412 (N_11412,N_11289,N_11388);
and U11413 (N_11413,N_11395,N_11329);
nand U11414 (N_11414,N_11294,N_11298);
nor U11415 (N_11415,N_11268,N_11236);
nor U11416 (N_11416,N_11214,N_11387);
xnor U11417 (N_11417,N_11286,N_11392);
xor U11418 (N_11418,N_11383,N_11341);
xor U11419 (N_11419,N_11228,N_11215);
and U11420 (N_11420,N_11293,N_11229);
nand U11421 (N_11421,N_11343,N_11244);
and U11422 (N_11422,N_11353,N_11278);
nand U11423 (N_11423,N_11240,N_11288);
xor U11424 (N_11424,N_11201,N_11390);
nor U11425 (N_11425,N_11336,N_11274);
nand U11426 (N_11426,N_11384,N_11299);
nor U11427 (N_11427,N_11357,N_11303);
or U11428 (N_11428,N_11295,N_11378);
or U11429 (N_11429,N_11279,N_11333);
nor U11430 (N_11430,N_11269,N_11249);
or U11431 (N_11431,N_11301,N_11386);
or U11432 (N_11432,N_11350,N_11206);
or U11433 (N_11433,N_11360,N_11399);
nand U11434 (N_11434,N_11212,N_11391);
nand U11435 (N_11435,N_11320,N_11200);
nand U11436 (N_11436,N_11266,N_11211);
or U11437 (N_11437,N_11277,N_11263);
or U11438 (N_11438,N_11305,N_11213);
and U11439 (N_11439,N_11325,N_11344);
xnor U11440 (N_11440,N_11304,N_11242);
nand U11441 (N_11441,N_11275,N_11346);
nand U11442 (N_11442,N_11292,N_11210);
nand U11443 (N_11443,N_11258,N_11372);
or U11444 (N_11444,N_11373,N_11230);
xnor U11445 (N_11445,N_11239,N_11237);
nor U11446 (N_11446,N_11326,N_11246);
or U11447 (N_11447,N_11355,N_11216);
and U11448 (N_11448,N_11302,N_11368);
or U11449 (N_11449,N_11318,N_11339);
nor U11450 (N_11450,N_11248,N_11382);
nand U11451 (N_11451,N_11231,N_11322);
nand U11452 (N_11452,N_11297,N_11280);
and U11453 (N_11453,N_11366,N_11358);
and U11454 (N_11454,N_11363,N_11349);
nor U11455 (N_11455,N_11241,N_11256);
xor U11456 (N_11456,N_11257,N_11306);
xor U11457 (N_11457,N_11290,N_11316);
nor U11458 (N_11458,N_11348,N_11367);
or U11459 (N_11459,N_11398,N_11313);
nand U11460 (N_11460,N_11315,N_11247);
nor U11461 (N_11461,N_11225,N_11202);
and U11462 (N_11462,N_11300,N_11205);
and U11463 (N_11463,N_11307,N_11321);
and U11464 (N_11464,N_11309,N_11352);
nor U11465 (N_11465,N_11351,N_11342);
and U11466 (N_11466,N_11323,N_11265);
and U11467 (N_11467,N_11370,N_11273);
nor U11468 (N_11468,N_11308,N_11245);
or U11469 (N_11469,N_11234,N_11251);
nor U11470 (N_11470,N_11374,N_11262);
nand U11471 (N_11471,N_11377,N_11219);
or U11472 (N_11472,N_11267,N_11361);
xor U11473 (N_11473,N_11243,N_11261);
or U11474 (N_11474,N_11397,N_11319);
xnor U11475 (N_11475,N_11283,N_11396);
nor U11476 (N_11476,N_11220,N_11204);
nor U11477 (N_11477,N_11334,N_11332);
nand U11478 (N_11478,N_11282,N_11381);
or U11479 (N_11479,N_11255,N_11327);
and U11480 (N_11480,N_11380,N_11389);
or U11481 (N_11481,N_11250,N_11287);
and U11482 (N_11482,N_11222,N_11232);
xnor U11483 (N_11483,N_11365,N_11393);
and U11484 (N_11484,N_11354,N_11203);
xor U11485 (N_11485,N_11314,N_11233);
nand U11486 (N_11486,N_11371,N_11331);
nand U11487 (N_11487,N_11252,N_11208);
or U11488 (N_11488,N_11264,N_11238);
xor U11489 (N_11489,N_11317,N_11359);
or U11490 (N_11490,N_11284,N_11254);
nand U11491 (N_11491,N_11271,N_11217);
xor U11492 (N_11492,N_11345,N_11324);
nor U11493 (N_11493,N_11310,N_11218);
or U11494 (N_11494,N_11227,N_11340);
and U11495 (N_11495,N_11260,N_11311);
or U11496 (N_11496,N_11376,N_11285);
or U11497 (N_11497,N_11330,N_11335);
nor U11498 (N_11498,N_11224,N_11276);
nor U11499 (N_11499,N_11235,N_11259);
xnor U11500 (N_11500,N_11362,N_11273);
xor U11501 (N_11501,N_11212,N_11365);
and U11502 (N_11502,N_11256,N_11219);
xor U11503 (N_11503,N_11257,N_11299);
and U11504 (N_11504,N_11214,N_11217);
xor U11505 (N_11505,N_11321,N_11225);
and U11506 (N_11506,N_11321,N_11229);
or U11507 (N_11507,N_11387,N_11309);
xnor U11508 (N_11508,N_11375,N_11274);
xor U11509 (N_11509,N_11373,N_11238);
and U11510 (N_11510,N_11235,N_11269);
xnor U11511 (N_11511,N_11333,N_11388);
nand U11512 (N_11512,N_11229,N_11237);
nand U11513 (N_11513,N_11251,N_11298);
nor U11514 (N_11514,N_11280,N_11251);
nor U11515 (N_11515,N_11370,N_11323);
xor U11516 (N_11516,N_11395,N_11233);
nand U11517 (N_11517,N_11306,N_11278);
or U11518 (N_11518,N_11343,N_11329);
xnor U11519 (N_11519,N_11366,N_11226);
or U11520 (N_11520,N_11342,N_11396);
and U11521 (N_11521,N_11362,N_11257);
and U11522 (N_11522,N_11378,N_11324);
nor U11523 (N_11523,N_11328,N_11285);
or U11524 (N_11524,N_11375,N_11257);
or U11525 (N_11525,N_11355,N_11203);
nor U11526 (N_11526,N_11306,N_11317);
xnor U11527 (N_11527,N_11349,N_11368);
nand U11528 (N_11528,N_11209,N_11333);
nor U11529 (N_11529,N_11287,N_11390);
xnor U11530 (N_11530,N_11301,N_11389);
nor U11531 (N_11531,N_11327,N_11226);
and U11532 (N_11532,N_11388,N_11214);
and U11533 (N_11533,N_11372,N_11249);
nor U11534 (N_11534,N_11374,N_11235);
nor U11535 (N_11535,N_11388,N_11205);
nand U11536 (N_11536,N_11367,N_11390);
and U11537 (N_11537,N_11372,N_11314);
nand U11538 (N_11538,N_11204,N_11398);
and U11539 (N_11539,N_11378,N_11273);
nor U11540 (N_11540,N_11262,N_11235);
nor U11541 (N_11541,N_11211,N_11380);
or U11542 (N_11542,N_11341,N_11388);
or U11543 (N_11543,N_11272,N_11390);
xor U11544 (N_11544,N_11299,N_11212);
nand U11545 (N_11545,N_11348,N_11234);
nor U11546 (N_11546,N_11290,N_11391);
nor U11547 (N_11547,N_11229,N_11256);
xor U11548 (N_11548,N_11392,N_11310);
xnor U11549 (N_11549,N_11351,N_11236);
xor U11550 (N_11550,N_11295,N_11249);
and U11551 (N_11551,N_11292,N_11368);
xor U11552 (N_11552,N_11381,N_11311);
or U11553 (N_11553,N_11234,N_11218);
xnor U11554 (N_11554,N_11361,N_11235);
and U11555 (N_11555,N_11205,N_11250);
nand U11556 (N_11556,N_11368,N_11324);
xnor U11557 (N_11557,N_11337,N_11224);
nor U11558 (N_11558,N_11380,N_11387);
or U11559 (N_11559,N_11317,N_11387);
or U11560 (N_11560,N_11341,N_11214);
and U11561 (N_11561,N_11381,N_11253);
or U11562 (N_11562,N_11353,N_11224);
and U11563 (N_11563,N_11392,N_11267);
or U11564 (N_11564,N_11318,N_11290);
nor U11565 (N_11565,N_11219,N_11209);
and U11566 (N_11566,N_11299,N_11216);
xnor U11567 (N_11567,N_11367,N_11298);
xnor U11568 (N_11568,N_11232,N_11390);
and U11569 (N_11569,N_11249,N_11260);
or U11570 (N_11570,N_11248,N_11276);
nand U11571 (N_11571,N_11364,N_11206);
xor U11572 (N_11572,N_11224,N_11302);
and U11573 (N_11573,N_11359,N_11245);
nor U11574 (N_11574,N_11210,N_11336);
or U11575 (N_11575,N_11266,N_11338);
or U11576 (N_11576,N_11243,N_11231);
and U11577 (N_11577,N_11203,N_11381);
xnor U11578 (N_11578,N_11208,N_11310);
nand U11579 (N_11579,N_11342,N_11340);
nand U11580 (N_11580,N_11247,N_11238);
xnor U11581 (N_11581,N_11263,N_11235);
nand U11582 (N_11582,N_11323,N_11275);
nor U11583 (N_11583,N_11291,N_11372);
nand U11584 (N_11584,N_11300,N_11390);
xnor U11585 (N_11585,N_11393,N_11373);
xor U11586 (N_11586,N_11205,N_11268);
nand U11587 (N_11587,N_11386,N_11365);
or U11588 (N_11588,N_11331,N_11235);
nand U11589 (N_11589,N_11336,N_11347);
nand U11590 (N_11590,N_11218,N_11319);
nor U11591 (N_11591,N_11267,N_11222);
or U11592 (N_11592,N_11249,N_11283);
nor U11593 (N_11593,N_11223,N_11238);
xnor U11594 (N_11594,N_11326,N_11309);
or U11595 (N_11595,N_11310,N_11235);
or U11596 (N_11596,N_11398,N_11229);
xnor U11597 (N_11597,N_11282,N_11286);
nand U11598 (N_11598,N_11360,N_11341);
nand U11599 (N_11599,N_11250,N_11276);
or U11600 (N_11600,N_11594,N_11468);
and U11601 (N_11601,N_11507,N_11589);
or U11602 (N_11602,N_11454,N_11447);
nand U11603 (N_11603,N_11595,N_11596);
and U11604 (N_11604,N_11446,N_11428);
nand U11605 (N_11605,N_11561,N_11484);
and U11606 (N_11606,N_11559,N_11433);
xor U11607 (N_11607,N_11544,N_11469);
xnor U11608 (N_11608,N_11543,N_11542);
or U11609 (N_11609,N_11449,N_11583);
and U11610 (N_11610,N_11475,N_11472);
or U11611 (N_11611,N_11438,N_11523);
nand U11612 (N_11612,N_11509,N_11505);
nand U11613 (N_11613,N_11502,N_11435);
nand U11614 (N_11614,N_11569,N_11577);
nor U11615 (N_11615,N_11551,N_11404);
nand U11616 (N_11616,N_11501,N_11546);
or U11617 (N_11617,N_11578,N_11526);
and U11618 (N_11618,N_11463,N_11567);
and U11619 (N_11619,N_11496,N_11455);
nand U11620 (N_11620,N_11541,N_11481);
nand U11621 (N_11621,N_11512,N_11440);
xor U11622 (N_11622,N_11548,N_11513);
xnor U11623 (N_11623,N_11492,N_11545);
xnor U11624 (N_11624,N_11429,N_11467);
xor U11625 (N_11625,N_11556,N_11464);
xor U11626 (N_11626,N_11430,N_11549);
nand U11627 (N_11627,N_11593,N_11465);
nand U11628 (N_11628,N_11476,N_11439);
and U11629 (N_11629,N_11498,N_11403);
and U11630 (N_11630,N_11407,N_11537);
or U11631 (N_11631,N_11497,N_11565);
xnor U11632 (N_11632,N_11508,N_11487);
xnor U11633 (N_11633,N_11524,N_11584);
nor U11634 (N_11634,N_11431,N_11585);
and U11635 (N_11635,N_11514,N_11536);
nand U11636 (N_11636,N_11448,N_11511);
xor U11637 (N_11637,N_11554,N_11410);
nand U11638 (N_11638,N_11568,N_11528);
nor U11639 (N_11639,N_11444,N_11591);
nor U11640 (N_11640,N_11480,N_11563);
and U11641 (N_11641,N_11408,N_11426);
or U11642 (N_11642,N_11598,N_11470);
nand U11643 (N_11643,N_11510,N_11425);
and U11644 (N_11644,N_11491,N_11570);
xor U11645 (N_11645,N_11489,N_11518);
nand U11646 (N_11646,N_11450,N_11406);
or U11647 (N_11647,N_11499,N_11564);
nor U11648 (N_11648,N_11471,N_11521);
or U11649 (N_11649,N_11416,N_11539);
or U11650 (N_11650,N_11417,N_11495);
or U11651 (N_11651,N_11547,N_11530);
nor U11652 (N_11652,N_11579,N_11405);
or U11653 (N_11653,N_11401,N_11432);
and U11654 (N_11654,N_11478,N_11503);
nor U11655 (N_11655,N_11573,N_11566);
nor U11656 (N_11656,N_11402,N_11400);
nor U11657 (N_11657,N_11443,N_11529);
and U11658 (N_11658,N_11445,N_11456);
nand U11659 (N_11659,N_11562,N_11479);
xnor U11660 (N_11660,N_11553,N_11436);
and U11661 (N_11661,N_11418,N_11415);
and U11662 (N_11662,N_11580,N_11574);
or U11663 (N_11663,N_11571,N_11590);
or U11664 (N_11664,N_11534,N_11540);
nand U11665 (N_11665,N_11588,N_11485);
and U11666 (N_11666,N_11599,N_11576);
and U11667 (N_11667,N_11506,N_11517);
xnor U11668 (N_11668,N_11477,N_11520);
or U11669 (N_11669,N_11460,N_11558);
nor U11670 (N_11670,N_11413,N_11473);
nand U11671 (N_11671,N_11586,N_11519);
or U11672 (N_11672,N_11515,N_11483);
or U11673 (N_11673,N_11424,N_11494);
xnor U11674 (N_11674,N_11592,N_11555);
and U11675 (N_11675,N_11442,N_11525);
nand U11676 (N_11676,N_11532,N_11516);
nand U11677 (N_11677,N_11557,N_11575);
nand U11678 (N_11678,N_11420,N_11482);
nand U11679 (N_11679,N_11422,N_11411);
nor U11680 (N_11680,N_11458,N_11597);
nor U11681 (N_11681,N_11538,N_11437);
or U11682 (N_11682,N_11522,N_11451);
xor U11683 (N_11683,N_11486,N_11504);
or U11684 (N_11684,N_11587,N_11462);
nand U11685 (N_11685,N_11412,N_11434);
or U11686 (N_11686,N_11493,N_11560);
nand U11687 (N_11687,N_11527,N_11427);
nand U11688 (N_11688,N_11459,N_11414);
and U11689 (N_11689,N_11474,N_11490);
nor U11690 (N_11690,N_11457,N_11466);
nand U11691 (N_11691,N_11500,N_11581);
nand U11692 (N_11692,N_11552,N_11572);
or U11693 (N_11693,N_11441,N_11533);
nor U11694 (N_11694,N_11531,N_11419);
xor U11695 (N_11695,N_11488,N_11421);
xnor U11696 (N_11696,N_11535,N_11550);
nand U11697 (N_11697,N_11409,N_11453);
xor U11698 (N_11698,N_11423,N_11582);
nor U11699 (N_11699,N_11452,N_11461);
nor U11700 (N_11700,N_11513,N_11421);
nor U11701 (N_11701,N_11546,N_11418);
or U11702 (N_11702,N_11447,N_11543);
xnor U11703 (N_11703,N_11448,N_11455);
or U11704 (N_11704,N_11493,N_11564);
xnor U11705 (N_11705,N_11542,N_11548);
xnor U11706 (N_11706,N_11569,N_11510);
nand U11707 (N_11707,N_11583,N_11441);
nor U11708 (N_11708,N_11538,N_11586);
or U11709 (N_11709,N_11520,N_11542);
and U11710 (N_11710,N_11489,N_11471);
nand U11711 (N_11711,N_11540,N_11493);
and U11712 (N_11712,N_11501,N_11564);
nand U11713 (N_11713,N_11411,N_11528);
and U11714 (N_11714,N_11520,N_11575);
nor U11715 (N_11715,N_11461,N_11570);
and U11716 (N_11716,N_11454,N_11506);
or U11717 (N_11717,N_11425,N_11513);
or U11718 (N_11718,N_11437,N_11537);
or U11719 (N_11719,N_11498,N_11424);
and U11720 (N_11720,N_11591,N_11548);
and U11721 (N_11721,N_11410,N_11474);
nor U11722 (N_11722,N_11544,N_11466);
and U11723 (N_11723,N_11549,N_11455);
xor U11724 (N_11724,N_11591,N_11462);
nand U11725 (N_11725,N_11480,N_11538);
nand U11726 (N_11726,N_11413,N_11422);
or U11727 (N_11727,N_11426,N_11570);
or U11728 (N_11728,N_11411,N_11489);
nor U11729 (N_11729,N_11511,N_11588);
and U11730 (N_11730,N_11437,N_11555);
nand U11731 (N_11731,N_11595,N_11552);
nand U11732 (N_11732,N_11583,N_11594);
xnor U11733 (N_11733,N_11449,N_11481);
nand U11734 (N_11734,N_11536,N_11422);
xnor U11735 (N_11735,N_11500,N_11448);
xnor U11736 (N_11736,N_11541,N_11437);
and U11737 (N_11737,N_11487,N_11584);
or U11738 (N_11738,N_11488,N_11409);
nand U11739 (N_11739,N_11531,N_11526);
nor U11740 (N_11740,N_11400,N_11547);
xnor U11741 (N_11741,N_11479,N_11519);
and U11742 (N_11742,N_11545,N_11439);
or U11743 (N_11743,N_11521,N_11415);
nor U11744 (N_11744,N_11533,N_11532);
nor U11745 (N_11745,N_11452,N_11470);
and U11746 (N_11746,N_11558,N_11523);
and U11747 (N_11747,N_11431,N_11562);
or U11748 (N_11748,N_11539,N_11535);
or U11749 (N_11749,N_11583,N_11557);
nor U11750 (N_11750,N_11598,N_11472);
nor U11751 (N_11751,N_11560,N_11508);
and U11752 (N_11752,N_11491,N_11454);
and U11753 (N_11753,N_11594,N_11540);
xor U11754 (N_11754,N_11484,N_11415);
xnor U11755 (N_11755,N_11480,N_11477);
nand U11756 (N_11756,N_11546,N_11515);
nand U11757 (N_11757,N_11421,N_11567);
nor U11758 (N_11758,N_11515,N_11502);
nor U11759 (N_11759,N_11588,N_11545);
or U11760 (N_11760,N_11495,N_11487);
nor U11761 (N_11761,N_11420,N_11403);
or U11762 (N_11762,N_11475,N_11536);
nand U11763 (N_11763,N_11554,N_11525);
or U11764 (N_11764,N_11559,N_11443);
nand U11765 (N_11765,N_11489,N_11424);
nor U11766 (N_11766,N_11503,N_11412);
and U11767 (N_11767,N_11557,N_11438);
or U11768 (N_11768,N_11483,N_11599);
or U11769 (N_11769,N_11564,N_11555);
or U11770 (N_11770,N_11531,N_11465);
and U11771 (N_11771,N_11580,N_11442);
nor U11772 (N_11772,N_11510,N_11511);
nor U11773 (N_11773,N_11420,N_11470);
nor U11774 (N_11774,N_11535,N_11549);
nand U11775 (N_11775,N_11516,N_11562);
and U11776 (N_11776,N_11450,N_11519);
nor U11777 (N_11777,N_11419,N_11513);
nor U11778 (N_11778,N_11432,N_11434);
or U11779 (N_11779,N_11435,N_11433);
and U11780 (N_11780,N_11426,N_11421);
and U11781 (N_11781,N_11550,N_11439);
xnor U11782 (N_11782,N_11422,N_11454);
and U11783 (N_11783,N_11524,N_11504);
or U11784 (N_11784,N_11549,N_11500);
or U11785 (N_11785,N_11509,N_11423);
xor U11786 (N_11786,N_11573,N_11527);
xor U11787 (N_11787,N_11480,N_11410);
xnor U11788 (N_11788,N_11409,N_11517);
nand U11789 (N_11789,N_11464,N_11547);
or U11790 (N_11790,N_11477,N_11542);
and U11791 (N_11791,N_11543,N_11424);
or U11792 (N_11792,N_11410,N_11412);
nor U11793 (N_11793,N_11572,N_11472);
and U11794 (N_11794,N_11474,N_11483);
and U11795 (N_11795,N_11488,N_11543);
nand U11796 (N_11796,N_11562,N_11429);
nor U11797 (N_11797,N_11530,N_11431);
xor U11798 (N_11798,N_11496,N_11532);
nor U11799 (N_11799,N_11527,N_11507);
and U11800 (N_11800,N_11694,N_11682);
or U11801 (N_11801,N_11652,N_11797);
or U11802 (N_11802,N_11698,N_11705);
nand U11803 (N_11803,N_11711,N_11741);
and U11804 (N_11804,N_11657,N_11732);
xor U11805 (N_11805,N_11701,N_11615);
xnor U11806 (N_11806,N_11785,N_11750);
nor U11807 (N_11807,N_11727,N_11619);
xor U11808 (N_11808,N_11790,N_11600);
and U11809 (N_11809,N_11607,N_11717);
nand U11810 (N_11810,N_11685,N_11639);
xor U11811 (N_11811,N_11658,N_11742);
and U11812 (N_11812,N_11667,N_11644);
xnor U11813 (N_11813,N_11755,N_11672);
and U11814 (N_11814,N_11788,N_11662);
or U11815 (N_11815,N_11630,N_11798);
nand U11816 (N_11816,N_11631,N_11663);
and U11817 (N_11817,N_11686,N_11641);
nand U11818 (N_11818,N_11603,N_11764);
and U11819 (N_11819,N_11684,N_11771);
nor U11820 (N_11820,N_11642,N_11616);
or U11821 (N_11821,N_11793,N_11775);
xnor U11822 (N_11822,N_11628,N_11740);
or U11823 (N_11823,N_11731,N_11734);
and U11824 (N_11824,N_11736,N_11646);
xnor U11825 (N_11825,N_11670,N_11660);
nor U11826 (N_11826,N_11635,N_11633);
nand U11827 (N_11827,N_11679,N_11689);
nor U11828 (N_11828,N_11782,N_11795);
xnor U11829 (N_11829,N_11620,N_11743);
or U11830 (N_11830,N_11674,N_11638);
nor U11831 (N_11831,N_11604,N_11666);
xnor U11832 (N_11832,N_11703,N_11612);
xnor U11833 (N_11833,N_11766,N_11721);
or U11834 (N_11834,N_11678,N_11702);
or U11835 (N_11835,N_11640,N_11738);
nand U11836 (N_11836,N_11773,N_11709);
and U11837 (N_11837,N_11699,N_11621);
or U11838 (N_11838,N_11602,N_11625);
nor U11839 (N_11839,N_11777,N_11611);
nor U11840 (N_11840,N_11624,N_11763);
xnor U11841 (N_11841,N_11723,N_11760);
or U11842 (N_11842,N_11791,N_11739);
nand U11843 (N_11843,N_11622,N_11735);
nand U11844 (N_11844,N_11729,N_11610);
nor U11845 (N_11845,N_11688,N_11784);
nand U11846 (N_11846,N_11716,N_11707);
nand U11847 (N_11847,N_11737,N_11726);
nand U11848 (N_11848,N_11655,N_11748);
and U11849 (N_11849,N_11697,N_11659);
and U11850 (N_11850,N_11747,N_11783);
or U11851 (N_11851,N_11781,N_11664);
or U11852 (N_11852,N_11643,N_11776);
or U11853 (N_11853,N_11687,N_11745);
or U11854 (N_11854,N_11751,N_11768);
nor U11855 (N_11855,N_11753,N_11700);
or U11856 (N_11856,N_11749,N_11758);
nor U11857 (N_11857,N_11759,N_11634);
and U11858 (N_11858,N_11617,N_11627);
or U11859 (N_11859,N_11724,N_11690);
and U11860 (N_11860,N_11719,N_11668);
or U11861 (N_11861,N_11713,N_11626);
nor U11862 (N_11862,N_11613,N_11681);
and U11863 (N_11863,N_11677,N_11650);
or U11864 (N_11864,N_11706,N_11754);
or U11865 (N_11865,N_11618,N_11714);
or U11866 (N_11866,N_11722,N_11695);
nand U11867 (N_11867,N_11733,N_11704);
nor U11868 (N_11868,N_11730,N_11654);
nand U11869 (N_11869,N_11651,N_11762);
nand U11870 (N_11870,N_11692,N_11669);
nor U11871 (N_11871,N_11725,N_11761);
or U11872 (N_11872,N_11787,N_11718);
nor U11873 (N_11873,N_11765,N_11680);
or U11874 (N_11874,N_11676,N_11614);
nor U11875 (N_11875,N_11696,N_11728);
xnor U11876 (N_11876,N_11712,N_11661);
nor U11877 (N_11877,N_11671,N_11796);
or U11878 (N_11878,N_11608,N_11794);
xnor U11879 (N_11879,N_11789,N_11675);
nor U11880 (N_11880,N_11778,N_11601);
or U11881 (N_11881,N_11780,N_11649);
xnor U11882 (N_11882,N_11767,N_11606);
nand U11883 (N_11883,N_11710,N_11693);
or U11884 (N_11884,N_11632,N_11770);
xor U11885 (N_11885,N_11720,N_11769);
xor U11886 (N_11886,N_11746,N_11708);
or U11887 (N_11887,N_11756,N_11715);
xnor U11888 (N_11888,N_11637,N_11665);
or U11889 (N_11889,N_11774,N_11656);
or U11890 (N_11890,N_11629,N_11744);
nand U11891 (N_11891,N_11799,N_11786);
xor U11892 (N_11892,N_11609,N_11757);
nor U11893 (N_11893,N_11645,N_11623);
and U11894 (N_11894,N_11772,N_11653);
nor U11895 (N_11895,N_11673,N_11752);
nor U11896 (N_11896,N_11636,N_11792);
or U11897 (N_11897,N_11648,N_11605);
xor U11898 (N_11898,N_11683,N_11691);
nor U11899 (N_11899,N_11647,N_11779);
and U11900 (N_11900,N_11612,N_11715);
nor U11901 (N_11901,N_11647,N_11611);
nand U11902 (N_11902,N_11755,N_11788);
xnor U11903 (N_11903,N_11788,N_11750);
nand U11904 (N_11904,N_11653,N_11619);
and U11905 (N_11905,N_11793,N_11633);
or U11906 (N_11906,N_11716,N_11631);
and U11907 (N_11907,N_11718,N_11745);
or U11908 (N_11908,N_11741,N_11653);
nor U11909 (N_11909,N_11629,N_11739);
or U11910 (N_11910,N_11690,N_11617);
nor U11911 (N_11911,N_11690,N_11667);
or U11912 (N_11912,N_11680,N_11647);
xor U11913 (N_11913,N_11724,N_11744);
nor U11914 (N_11914,N_11717,N_11775);
or U11915 (N_11915,N_11777,N_11744);
nor U11916 (N_11916,N_11684,N_11712);
xor U11917 (N_11917,N_11715,N_11607);
nor U11918 (N_11918,N_11659,N_11638);
or U11919 (N_11919,N_11734,N_11674);
xor U11920 (N_11920,N_11776,N_11635);
nor U11921 (N_11921,N_11695,N_11767);
and U11922 (N_11922,N_11646,N_11621);
nor U11923 (N_11923,N_11764,N_11630);
nor U11924 (N_11924,N_11762,N_11652);
nand U11925 (N_11925,N_11717,N_11609);
xnor U11926 (N_11926,N_11708,N_11718);
nand U11927 (N_11927,N_11708,N_11714);
and U11928 (N_11928,N_11616,N_11791);
or U11929 (N_11929,N_11707,N_11640);
or U11930 (N_11930,N_11614,N_11682);
and U11931 (N_11931,N_11791,N_11734);
nor U11932 (N_11932,N_11793,N_11705);
xor U11933 (N_11933,N_11741,N_11641);
and U11934 (N_11934,N_11729,N_11664);
nand U11935 (N_11935,N_11789,N_11781);
or U11936 (N_11936,N_11637,N_11653);
and U11937 (N_11937,N_11704,N_11604);
nand U11938 (N_11938,N_11704,N_11654);
xor U11939 (N_11939,N_11731,N_11641);
nand U11940 (N_11940,N_11665,N_11682);
nand U11941 (N_11941,N_11643,N_11681);
nand U11942 (N_11942,N_11680,N_11791);
and U11943 (N_11943,N_11717,N_11770);
or U11944 (N_11944,N_11706,N_11601);
nand U11945 (N_11945,N_11719,N_11688);
and U11946 (N_11946,N_11716,N_11784);
and U11947 (N_11947,N_11717,N_11783);
nand U11948 (N_11948,N_11709,N_11703);
nor U11949 (N_11949,N_11714,N_11676);
xnor U11950 (N_11950,N_11737,N_11685);
and U11951 (N_11951,N_11610,N_11791);
or U11952 (N_11952,N_11785,N_11760);
nand U11953 (N_11953,N_11693,N_11665);
xnor U11954 (N_11954,N_11631,N_11626);
and U11955 (N_11955,N_11772,N_11705);
and U11956 (N_11956,N_11715,N_11694);
and U11957 (N_11957,N_11605,N_11783);
nand U11958 (N_11958,N_11675,N_11639);
or U11959 (N_11959,N_11772,N_11689);
xnor U11960 (N_11960,N_11761,N_11716);
and U11961 (N_11961,N_11696,N_11698);
or U11962 (N_11962,N_11611,N_11623);
and U11963 (N_11963,N_11609,N_11670);
or U11964 (N_11964,N_11637,N_11767);
or U11965 (N_11965,N_11781,N_11798);
or U11966 (N_11966,N_11663,N_11763);
and U11967 (N_11967,N_11693,N_11688);
xor U11968 (N_11968,N_11612,N_11645);
xnor U11969 (N_11969,N_11696,N_11743);
nand U11970 (N_11970,N_11770,N_11636);
nand U11971 (N_11971,N_11611,N_11732);
nand U11972 (N_11972,N_11661,N_11650);
xor U11973 (N_11973,N_11732,N_11636);
and U11974 (N_11974,N_11788,N_11602);
nor U11975 (N_11975,N_11730,N_11663);
or U11976 (N_11976,N_11766,N_11619);
nor U11977 (N_11977,N_11605,N_11721);
nand U11978 (N_11978,N_11724,N_11685);
and U11979 (N_11979,N_11625,N_11639);
and U11980 (N_11980,N_11697,N_11691);
xor U11981 (N_11981,N_11685,N_11720);
xor U11982 (N_11982,N_11650,N_11672);
xor U11983 (N_11983,N_11636,N_11640);
or U11984 (N_11984,N_11609,N_11716);
nor U11985 (N_11985,N_11753,N_11637);
or U11986 (N_11986,N_11617,N_11721);
and U11987 (N_11987,N_11793,N_11648);
nand U11988 (N_11988,N_11622,N_11676);
nor U11989 (N_11989,N_11679,N_11678);
nand U11990 (N_11990,N_11769,N_11662);
xor U11991 (N_11991,N_11638,N_11616);
and U11992 (N_11992,N_11696,N_11747);
nand U11993 (N_11993,N_11639,N_11638);
nor U11994 (N_11994,N_11695,N_11627);
nor U11995 (N_11995,N_11675,N_11759);
nor U11996 (N_11996,N_11602,N_11624);
or U11997 (N_11997,N_11765,N_11748);
and U11998 (N_11998,N_11794,N_11720);
or U11999 (N_11999,N_11753,N_11790);
and U12000 (N_12000,N_11958,N_11940);
or U12001 (N_12001,N_11852,N_11994);
xnor U12002 (N_12002,N_11986,N_11979);
xor U12003 (N_12003,N_11907,N_11833);
xor U12004 (N_12004,N_11830,N_11855);
nand U12005 (N_12005,N_11921,N_11926);
xor U12006 (N_12006,N_11809,N_11963);
xnor U12007 (N_12007,N_11814,N_11891);
nand U12008 (N_12008,N_11898,N_11983);
nor U12009 (N_12009,N_11853,N_11992);
nor U12010 (N_12010,N_11864,N_11900);
xnor U12011 (N_12011,N_11820,N_11863);
and U12012 (N_12012,N_11970,N_11896);
or U12013 (N_12013,N_11819,N_11893);
nand U12014 (N_12014,N_11959,N_11949);
and U12015 (N_12015,N_11918,N_11845);
xnor U12016 (N_12016,N_11930,N_11905);
nand U12017 (N_12017,N_11812,N_11857);
and U12018 (N_12018,N_11991,N_11880);
or U12019 (N_12019,N_11860,N_11861);
nand U12020 (N_12020,N_11936,N_11965);
or U12021 (N_12021,N_11945,N_11929);
and U12022 (N_12022,N_11976,N_11817);
xor U12023 (N_12023,N_11935,N_11973);
and U12024 (N_12024,N_11876,N_11826);
or U12025 (N_12025,N_11980,N_11834);
nand U12026 (N_12026,N_11866,N_11934);
nor U12027 (N_12027,N_11974,N_11838);
nand U12028 (N_12028,N_11989,N_11953);
nand U12029 (N_12029,N_11908,N_11951);
and U12030 (N_12030,N_11923,N_11913);
or U12031 (N_12031,N_11968,N_11952);
and U12032 (N_12032,N_11844,N_11962);
xnor U12033 (N_12033,N_11858,N_11977);
nor U12034 (N_12034,N_11899,N_11878);
nand U12035 (N_12035,N_11868,N_11933);
nor U12036 (N_12036,N_11990,N_11881);
and U12037 (N_12037,N_11984,N_11993);
or U12038 (N_12038,N_11997,N_11897);
or U12039 (N_12039,N_11960,N_11942);
and U12040 (N_12040,N_11884,N_11919);
nand U12041 (N_12041,N_11943,N_11944);
or U12042 (N_12042,N_11969,N_11922);
nor U12043 (N_12043,N_11810,N_11867);
xnor U12044 (N_12044,N_11800,N_11988);
or U12045 (N_12045,N_11862,N_11957);
nor U12046 (N_12046,N_11815,N_11859);
and U12047 (N_12047,N_11901,N_11879);
and U12048 (N_12048,N_11917,N_11827);
and U12049 (N_12049,N_11840,N_11839);
nand U12050 (N_12050,N_11967,N_11869);
nand U12051 (N_12051,N_11801,N_11854);
or U12052 (N_12052,N_11874,N_11914);
xor U12053 (N_12053,N_11920,N_11909);
nand U12054 (N_12054,N_11882,N_11894);
or U12055 (N_12055,N_11803,N_11831);
or U12056 (N_12056,N_11883,N_11956);
nor U12057 (N_12057,N_11823,N_11811);
nor U12058 (N_12058,N_11902,N_11982);
and U12059 (N_12059,N_11871,N_11821);
nor U12060 (N_12060,N_11938,N_11931);
or U12061 (N_12061,N_11955,N_11837);
or U12062 (N_12062,N_11806,N_11948);
or U12063 (N_12063,N_11996,N_11906);
and U12064 (N_12064,N_11892,N_11822);
nor U12065 (N_12065,N_11824,N_11903);
or U12066 (N_12066,N_11886,N_11865);
nand U12067 (N_12067,N_11964,N_11828);
nor U12068 (N_12068,N_11813,N_11981);
xnor U12069 (N_12069,N_11954,N_11848);
xor U12070 (N_12070,N_11987,N_11999);
nor U12071 (N_12071,N_11829,N_11804);
nand U12072 (N_12072,N_11851,N_11916);
or U12073 (N_12073,N_11932,N_11802);
nand U12074 (N_12074,N_11870,N_11888);
and U12075 (N_12075,N_11808,N_11842);
and U12076 (N_12076,N_11895,N_11873);
or U12077 (N_12077,N_11910,N_11875);
nor U12078 (N_12078,N_11928,N_11805);
nor U12079 (N_12079,N_11978,N_11832);
and U12080 (N_12080,N_11872,N_11847);
nand U12081 (N_12081,N_11966,N_11885);
xnor U12082 (N_12082,N_11915,N_11972);
nor U12083 (N_12083,N_11841,N_11807);
xnor U12084 (N_12084,N_11849,N_11904);
xnor U12085 (N_12085,N_11846,N_11911);
xor U12086 (N_12086,N_11985,N_11939);
and U12087 (N_12087,N_11887,N_11843);
or U12088 (N_12088,N_11924,N_11877);
or U12089 (N_12089,N_11850,N_11950);
nor U12090 (N_12090,N_11927,N_11925);
nand U12091 (N_12091,N_11971,N_11947);
and U12092 (N_12092,N_11961,N_11836);
nand U12093 (N_12093,N_11998,N_11975);
nor U12094 (N_12094,N_11818,N_11890);
nand U12095 (N_12095,N_11889,N_11825);
nand U12096 (N_12096,N_11835,N_11856);
and U12097 (N_12097,N_11816,N_11946);
or U12098 (N_12098,N_11912,N_11937);
xor U12099 (N_12099,N_11941,N_11995);
or U12100 (N_12100,N_11847,N_11875);
nand U12101 (N_12101,N_11969,N_11822);
or U12102 (N_12102,N_11834,N_11811);
and U12103 (N_12103,N_11968,N_11848);
nand U12104 (N_12104,N_11995,N_11873);
xnor U12105 (N_12105,N_11929,N_11915);
and U12106 (N_12106,N_11919,N_11994);
or U12107 (N_12107,N_11942,N_11822);
nand U12108 (N_12108,N_11998,N_11833);
nor U12109 (N_12109,N_11916,N_11855);
nand U12110 (N_12110,N_11968,N_11872);
and U12111 (N_12111,N_11976,N_11900);
and U12112 (N_12112,N_11918,N_11940);
nand U12113 (N_12113,N_11980,N_11847);
nor U12114 (N_12114,N_11957,N_11983);
xnor U12115 (N_12115,N_11816,N_11874);
or U12116 (N_12116,N_11893,N_11807);
xnor U12117 (N_12117,N_11924,N_11911);
nand U12118 (N_12118,N_11914,N_11899);
nand U12119 (N_12119,N_11925,N_11899);
or U12120 (N_12120,N_11981,N_11915);
xor U12121 (N_12121,N_11862,N_11867);
nor U12122 (N_12122,N_11886,N_11984);
or U12123 (N_12123,N_11979,N_11869);
nand U12124 (N_12124,N_11822,N_11963);
nand U12125 (N_12125,N_11993,N_11933);
nor U12126 (N_12126,N_11988,N_11949);
xnor U12127 (N_12127,N_11885,N_11988);
and U12128 (N_12128,N_11842,N_11887);
nand U12129 (N_12129,N_11876,N_11997);
or U12130 (N_12130,N_11879,N_11819);
nand U12131 (N_12131,N_11945,N_11965);
or U12132 (N_12132,N_11868,N_11961);
nor U12133 (N_12133,N_11840,N_11821);
or U12134 (N_12134,N_11925,N_11877);
and U12135 (N_12135,N_11919,N_11856);
nor U12136 (N_12136,N_11917,N_11993);
xor U12137 (N_12137,N_11925,N_11870);
or U12138 (N_12138,N_11835,N_11836);
nor U12139 (N_12139,N_11914,N_11813);
nor U12140 (N_12140,N_11879,N_11964);
nor U12141 (N_12141,N_11861,N_11985);
nand U12142 (N_12142,N_11951,N_11921);
nor U12143 (N_12143,N_11912,N_11952);
xor U12144 (N_12144,N_11838,N_11911);
nand U12145 (N_12145,N_11942,N_11828);
nand U12146 (N_12146,N_11853,N_11873);
and U12147 (N_12147,N_11864,N_11850);
xor U12148 (N_12148,N_11866,N_11988);
nand U12149 (N_12149,N_11921,N_11833);
and U12150 (N_12150,N_11904,N_11894);
or U12151 (N_12151,N_11917,N_11994);
nor U12152 (N_12152,N_11828,N_11869);
and U12153 (N_12153,N_11920,N_11807);
nand U12154 (N_12154,N_11963,N_11966);
or U12155 (N_12155,N_11932,N_11901);
xor U12156 (N_12156,N_11900,N_11837);
nand U12157 (N_12157,N_11972,N_11827);
or U12158 (N_12158,N_11969,N_11811);
and U12159 (N_12159,N_11895,N_11878);
or U12160 (N_12160,N_11925,N_11831);
or U12161 (N_12161,N_11909,N_11999);
xor U12162 (N_12162,N_11904,N_11885);
and U12163 (N_12163,N_11823,N_11851);
and U12164 (N_12164,N_11825,N_11993);
and U12165 (N_12165,N_11990,N_11897);
xnor U12166 (N_12166,N_11977,N_11928);
or U12167 (N_12167,N_11995,N_11992);
nor U12168 (N_12168,N_11870,N_11946);
xnor U12169 (N_12169,N_11961,N_11956);
nor U12170 (N_12170,N_11974,N_11922);
or U12171 (N_12171,N_11971,N_11952);
xnor U12172 (N_12172,N_11987,N_11956);
or U12173 (N_12173,N_11880,N_11852);
nor U12174 (N_12174,N_11884,N_11816);
and U12175 (N_12175,N_11983,N_11819);
xnor U12176 (N_12176,N_11868,N_11948);
and U12177 (N_12177,N_11984,N_11830);
xor U12178 (N_12178,N_11926,N_11826);
nand U12179 (N_12179,N_11810,N_11963);
nand U12180 (N_12180,N_11854,N_11849);
nand U12181 (N_12181,N_11932,N_11819);
or U12182 (N_12182,N_11885,N_11936);
xor U12183 (N_12183,N_11883,N_11821);
or U12184 (N_12184,N_11905,N_11891);
or U12185 (N_12185,N_11856,N_11969);
xor U12186 (N_12186,N_11945,N_11928);
nand U12187 (N_12187,N_11860,N_11873);
nor U12188 (N_12188,N_11909,N_11816);
nand U12189 (N_12189,N_11952,N_11905);
nand U12190 (N_12190,N_11872,N_11991);
xnor U12191 (N_12191,N_11972,N_11880);
xor U12192 (N_12192,N_11997,N_11901);
xnor U12193 (N_12193,N_11924,N_11895);
xor U12194 (N_12194,N_11860,N_11815);
nor U12195 (N_12195,N_11837,N_11932);
xnor U12196 (N_12196,N_11850,N_11966);
xor U12197 (N_12197,N_11953,N_11960);
and U12198 (N_12198,N_11939,N_11952);
xnor U12199 (N_12199,N_11833,N_11817);
xnor U12200 (N_12200,N_12041,N_12025);
xor U12201 (N_12201,N_12143,N_12090);
xor U12202 (N_12202,N_12014,N_12105);
nor U12203 (N_12203,N_12187,N_12083);
and U12204 (N_12204,N_12113,N_12050);
xor U12205 (N_12205,N_12116,N_12075);
nand U12206 (N_12206,N_12148,N_12033);
nor U12207 (N_12207,N_12030,N_12137);
or U12208 (N_12208,N_12173,N_12161);
nand U12209 (N_12209,N_12107,N_12003);
and U12210 (N_12210,N_12051,N_12066);
nand U12211 (N_12211,N_12037,N_12130);
and U12212 (N_12212,N_12154,N_12039);
nand U12213 (N_12213,N_12182,N_12126);
xor U12214 (N_12214,N_12031,N_12132);
or U12215 (N_12215,N_12142,N_12034);
nand U12216 (N_12216,N_12067,N_12035);
nor U12217 (N_12217,N_12159,N_12185);
nor U12218 (N_12218,N_12131,N_12118);
and U12219 (N_12219,N_12189,N_12072);
nand U12220 (N_12220,N_12193,N_12146);
nor U12221 (N_12221,N_12135,N_12099);
nand U12222 (N_12222,N_12054,N_12048);
nand U12223 (N_12223,N_12106,N_12018);
xnor U12224 (N_12224,N_12152,N_12156);
nor U12225 (N_12225,N_12063,N_12027);
or U12226 (N_12226,N_12134,N_12023);
and U12227 (N_12227,N_12078,N_12124);
and U12228 (N_12228,N_12024,N_12017);
and U12229 (N_12229,N_12123,N_12022);
nor U12230 (N_12230,N_12155,N_12028);
xnor U12231 (N_12231,N_12070,N_12056);
nor U12232 (N_12232,N_12151,N_12046);
xnor U12233 (N_12233,N_12176,N_12007);
and U12234 (N_12234,N_12112,N_12086);
or U12235 (N_12235,N_12040,N_12180);
or U12236 (N_12236,N_12062,N_12069);
nor U12237 (N_12237,N_12047,N_12144);
nor U12238 (N_12238,N_12160,N_12188);
and U12239 (N_12239,N_12006,N_12068);
nor U12240 (N_12240,N_12065,N_12094);
and U12241 (N_12241,N_12101,N_12122);
or U12242 (N_12242,N_12038,N_12197);
and U12243 (N_12243,N_12133,N_12195);
and U12244 (N_12244,N_12081,N_12163);
xnor U12245 (N_12245,N_12089,N_12115);
nor U12246 (N_12246,N_12061,N_12000);
xor U12247 (N_12247,N_12172,N_12184);
and U12248 (N_12248,N_12079,N_12042);
nand U12249 (N_12249,N_12002,N_12192);
and U12250 (N_12250,N_12036,N_12170);
nor U12251 (N_12251,N_12167,N_12114);
xor U12252 (N_12252,N_12153,N_12080);
xor U12253 (N_12253,N_12019,N_12026);
xnor U12254 (N_12254,N_12128,N_12129);
nor U12255 (N_12255,N_12140,N_12057);
and U12256 (N_12256,N_12013,N_12104);
nor U12257 (N_12257,N_12071,N_12165);
and U12258 (N_12258,N_12029,N_12044);
nor U12259 (N_12259,N_12136,N_12088);
or U12260 (N_12260,N_12059,N_12150);
or U12261 (N_12261,N_12120,N_12005);
nand U12262 (N_12262,N_12191,N_12084);
or U12263 (N_12263,N_12141,N_12103);
or U12264 (N_12264,N_12181,N_12096);
xor U12265 (N_12265,N_12074,N_12060);
nor U12266 (N_12266,N_12077,N_12053);
xor U12267 (N_12267,N_12064,N_12073);
and U12268 (N_12268,N_12108,N_12093);
xor U12269 (N_12269,N_12009,N_12121);
xnor U12270 (N_12270,N_12032,N_12085);
and U12271 (N_12271,N_12174,N_12102);
or U12272 (N_12272,N_12190,N_12138);
and U12273 (N_12273,N_12171,N_12169);
or U12274 (N_12274,N_12021,N_12175);
nand U12275 (N_12275,N_12194,N_12020);
or U12276 (N_12276,N_12119,N_12091);
xor U12277 (N_12277,N_12095,N_12097);
or U12278 (N_12278,N_12179,N_12186);
nor U12279 (N_12279,N_12058,N_12139);
xor U12280 (N_12280,N_12016,N_12178);
nor U12281 (N_12281,N_12196,N_12109);
nor U12282 (N_12282,N_12012,N_12052);
nor U12283 (N_12283,N_12117,N_12166);
xor U12284 (N_12284,N_12100,N_12145);
or U12285 (N_12285,N_12015,N_12082);
and U12286 (N_12286,N_12049,N_12177);
or U12287 (N_12287,N_12076,N_12111);
nand U12288 (N_12288,N_12004,N_12127);
or U12289 (N_12289,N_12164,N_12043);
nand U12290 (N_12290,N_12092,N_12162);
xor U12291 (N_12291,N_12198,N_12125);
nor U12292 (N_12292,N_12110,N_12199);
xor U12293 (N_12293,N_12010,N_12149);
nand U12294 (N_12294,N_12158,N_12045);
or U12295 (N_12295,N_12008,N_12055);
nand U12296 (N_12296,N_12001,N_12183);
nor U12297 (N_12297,N_12098,N_12147);
xnor U12298 (N_12298,N_12168,N_12011);
nand U12299 (N_12299,N_12087,N_12157);
and U12300 (N_12300,N_12124,N_12145);
and U12301 (N_12301,N_12049,N_12066);
or U12302 (N_12302,N_12159,N_12122);
nor U12303 (N_12303,N_12197,N_12162);
nor U12304 (N_12304,N_12156,N_12137);
nor U12305 (N_12305,N_12062,N_12091);
xnor U12306 (N_12306,N_12149,N_12179);
and U12307 (N_12307,N_12084,N_12142);
nor U12308 (N_12308,N_12004,N_12072);
nor U12309 (N_12309,N_12198,N_12060);
xor U12310 (N_12310,N_12128,N_12034);
nand U12311 (N_12311,N_12043,N_12037);
nor U12312 (N_12312,N_12016,N_12095);
nor U12313 (N_12313,N_12102,N_12025);
xnor U12314 (N_12314,N_12120,N_12088);
nor U12315 (N_12315,N_12135,N_12148);
nand U12316 (N_12316,N_12103,N_12038);
nor U12317 (N_12317,N_12007,N_12048);
or U12318 (N_12318,N_12133,N_12167);
and U12319 (N_12319,N_12081,N_12175);
nand U12320 (N_12320,N_12163,N_12189);
nor U12321 (N_12321,N_12199,N_12135);
nand U12322 (N_12322,N_12021,N_12030);
nand U12323 (N_12323,N_12011,N_12069);
nand U12324 (N_12324,N_12117,N_12103);
xor U12325 (N_12325,N_12125,N_12140);
and U12326 (N_12326,N_12104,N_12053);
nor U12327 (N_12327,N_12173,N_12158);
or U12328 (N_12328,N_12068,N_12069);
or U12329 (N_12329,N_12189,N_12181);
and U12330 (N_12330,N_12153,N_12091);
and U12331 (N_12331,N_12015,N_12196);
or U12332 (N_12332,N_12097,N_12051);
and U12333 (N_12333,N_12049,N_12136);
nand U12334 (N_12334,N_12103,N_12076);
nand U12335 (N_12335,N_12005,N_12040);
and U12336 (N_12336,N_12026,N_12182);
xor U12337 (N_12337,N_12193,N_12112);
xor U12338 (N_12338,N_12015,N_12131);
or U12339 (N_12339,N_12037,N_12006);
nor U12340 (N_12340,N_12064,N_12030);
and U12341 (N_12341,N_12137,N_12006);
nand U12342 (N_12342,N_12025,N_12192);
and U12343 (N_12343,N_12198,N_12170);
xor U12344 (N_12344,N_12107,N_12016);
and U12345 (N_12345,N_12150,N_12168);
nor U12346 (N_12346,N_12164,N_12112);
xnor U12347 (N_12347,N_12074,N_12000);
and U12348 (N_12348,N_12076,N_12190);
nand U12349 (N_12349,N_12143,N_12169);
xnor U12350 (N_12350,N_12075,N_12159);
xor U12351 (N_12351,N_12067,N_12115);
nor U12352 (N_12352,N_12176,N_12000);
or U12353 (N_12353,N_12184,N_12069);
or U12354 (N_12354,N_12009,N_12013);
and U12355 (N_12355,N_12196,N_12123);
or U12356 (N_12356,N_12014,N_12179);
nor U12357 (N_12357,N_12084,N_12094);
xnor U12358 (N_12358,N_12117,N_12168);
or U12359 (N_12359,N_12164,N_12149);
nor U12360 (N_12360,N_12024,N_12158);
xor U12361 (N_12361,N_12012,N_12013);
or U12362 (N_12362,N_12085,N_12103);
xnor U12363 (N_12363,N_12153,N_12112);
nor U12364 (N_12364,N_12109,N_12125);
nor U12365 (N_12365,N_12129,N_12187);
or U12366 (N_12366,N_12176,N_12037);
and U12367 (N_12367,N_12060,N_12046);
xor U12368 (N_12368,N_12013,N_12125);
nor U12369 (N_12369,N_12004,N_12150);
or U12370 (N_12370,N_12163,N_12113);
and U12371 (N_12371,N_12170,N_12143);
and U12372 (N_12372,N_12048,N_12021);
nand U12373 (N_12373,N_12042,N_12106);
xor U12374 (N_12374,N_12062,N_12085);
xnor U12375 (N_12375,N_12057,N_12115);
or U12376 (N_12376,N_12190,N_12139);
nand U12377 (N_12377,N_12082,N_12102);
xnor U12378 (N_12378,N_12015,N_12129);
xnor U12379 (N_12379,N_12121,N_12005);
xor U12380 (N_12380,N_12021,N_12044);
nor U12381 (N_12381,N_12097,N_12165);
xor U12382 (N_12382,N_12123,N_12053);
nand U12383 (N_12383,N_12008,N_12146);
nor U12384 (N_12384,N_12069,N_12111);
and U12385 (N_12385,N_12133,N_12024);
nand U12386 (N_12386,N_12168,N_12008);
and U12387 (N_12387,N_12121,N_12088);
xor U12388 (N_12388,N_12039,N_12120);
xor U12389 (N_12389,N_12027,N_12124);
or U12390 (N_12390,N_12185,N_12042);
nor U12391 (N_12391,N_12038,N_12060);
or U12392 (N_12392,N_12123,N_12173);
and U12393 (N_12393,N_12014,N_12095);
or U12394 (N_12394,N_12069,N_12040);
xnor U12395 (N_12395,N_12143,N_12048);
nand U12396 (N_12396,N_12082,N_12130);
nor U12397 (N_12397,N_12172,N_12000);
or U12398 (N_12398,N_12035,N_12029);
or U12399 (N_12399,N_12191,N_12086);
or U12400 (N_12400,N_12246,N_12243);
or U12401 (N_12401,N_12200,N_12241);
xnor U12402 (N_12402,N_12314,N_12267);
or U12403 (N_12403,N_12342,N_12316);
nor U12404 (N_12404,N_12250,N_12397);
nand U12405 (N_12405,N_12323,N_12318);
and U12406 (N_12406,N_12286,N_12335);
xor U12407 (N_12407,N_12237,N_12333);
or U12408 (N_12408,N_12213,N_12387);
nor U12409 (N_12409,N_12298,N_12370);
and U12410 (N_12410,N_12365,N_12215);
xnor U12411 (N_12411,N_12385,N_12393);
nand U12412 (N_12412,N_12258,N_12339);
nand U12413 (N_12413,N_12277,N_12312);
and U12414 (N_12414,N_12315,N_12260);
and U12415 (N_12415,N_12281,N_12297);
nor U12416 (N_12416,N_12249,N_12271);
and U12417 (N_12417,N_12233,N_12367);
xor U12418 (N_12418,N_12341,N_12372);
nand U12419 (N_12419,N_12302,N_12350);
or U12420 (N_12420,N_12357,N_12324);
xnor U12421 (N_12421,N_12394,N_12236);
nor U12422 (N_12422,N_12280,N_12245);
nor U12423 (N_12423,N_12327,N_12217);
and U12424 (N_12424,N_12306,N_12304);
xnor U12425 (N_12425,N_12309,N_12353);
nor U12426 (N_12426,N_12264,N_12334);
nand U12427 (N_12427,N_12368,N_12235);
nand U12428 (N_12428,N_12225,N_12322);
nand U12429 (N_12429,N_12285,N_12336);
xnor U12430 (N_12430,N_12374,N_12305);
or U12431 (N_12431,N_12279,N_12303);
and U12432 (N_12432,N_12205,N_12240);
xor U12433 (N_12433,N_12253,N_12256);
or U12434 (N_12434,N_12399,N_12263);
or U12435 (N_12435,N_12265,N_12288);
xnor U12436 (N_12436,N_12310,N_12222);
and U12437 (N_12437,N_12278,N_12290);
xnor U12438 (N_12438,N_12344,N_12261);
xnor U12439 (N_12439,N_12377,N_12262);
xnor U12440 (N_12440,N_12358,N_12269);
or U12441 (N_12441,N_12211,N_12202);
xnor U12442 (N_12442,N_12375,N_12380);
nor U12443 (N_12443,N_12234,N_12383);
and U12444 (N_12444,N_12390,N_12227);
nand U12445 (N_12445,N_12294,N_12382);
or U12446 (N_12446,N_12284,N_12347);
nand U12447 (N_12447,N_12376,N_12301);
or U12448 (N_12448,N_12299,N_12228);
xnor U12449 (N_12449,N_12292,N_12275);
and U12450 (N_12450,N_12224,N_12362);
or U12451 (N_12451,N_12360,N_12330);
xnor U12452 (N_12452,N_12254,N_12308);
or U12453 (N_12453,N_12212,N_12274);
nor U12454 (N_12454,N_12244,N_12221);
or U12455 (N_12455,N_12231,N_12238);
nand U12456 (N_12456,N_12338,N_12252);
and U12457 (N_12457,N_12296,N_12201);
and U12458 (N_12458,N_12317,N_12349);
and U12459 (N_12459,N_12326,N_12369);
or U12460 (N_12460,N_12346,N_12251);
and U12461 (N_12461,N_12332,N_12398);
nor U12462 (N_12462,N_12207,N_12340);
and U12463 (N_12463,N_12282,N_12384);
nand U12464 (N_12464,N_12214,N_12355);
and U12465 (N_12465,N_12396,N_12371);
xnor U12466 (N_12466,N_12366,N_12307);
nor U12467 (N_12467,N_12232,N_12361);
xnor U12468 (N_12468,N_12257,N_12255);
xor U12469 (N_12469,N_12389,N_12356);
and U12470 (N_12470,N_12359,N_12378);
or U12471 (N_12471,N_12329,N_12345);
nor U12472 (N_12472,N_12386,N_12352);
or U12473 (N_12473,N_12321,N_12206);
xor U12474 (N_12474,N_12220,N_12328);
or U12475 (N_12475,N_12242,N_12229);
nand U12476 (N_12476,N_12247,N_12319);
xnor U12477 (N_12477,N_12219,N_12295);
nand U12478 (N_12478,N_12320,N_12331);
nor U12479 (N_12479,N_12351,N_12287);
or U12480 (N_12480,N_12239,N_12325);
nor U12481 (N_12481,N_12273,N_12203);
xor U12482 (N_12482,N_12270,N_12266);
or U12483 (N_12483,N_12226,N_12283);
and U12484 (N_12484,N_12364,N_12230);
and U12485 (N_12485,N_12291,N_12204);
or U12486 (N_12486,N_12276,N_12373);
xor U12487 (N_12487,N_12300,N_12272);
and U12488 (N_12488,N_12208,N_12248);
nand U12489 (N_12489,N_12223,N_12311);
nand U12490 (N_12490,N_12289,N_12218);
xor U12491 (N_12491,N_12209,N_12354);
or U12492 (N_12492,N_12343,N_12268);
nor U12493 (N_12493,N_12210,N_12293);
nand U12494 (N_12494,N_12363,N_12348);
or U12495 (N_12495,N_12313,N_12381);
xnor U12496 (N_12496,N_12259,N_12379);
or U12497 (N_12497,N_12395,N_12337);
or U12498 (N_12498,N_12392,N_12388);
nor U12499 (N_12499,N_12391,N_12216);
xnor U12500 (N_12500,N_12222,N_12284);
and U12501 (N_12501,N_12253,N_12334);
xor U12502 (N_12502,N_12332,N_12299);
nand U12503 (N_12503,N_12286,N_12389);
and U12504 (N_12504,N_12220,N_12370);
xnor U12505 (N_12505,N_12384,N_12399);
nor U12506 (N_12506,N_12359,N_12272);
nor U12507 (N_12507,N_12313,N_12320);
or U12508 (N_12508,N_12344,N_12269);
and U12509 (N_12509,N_12357,N_12305);
or U12510 (N_12510,N_12393,N_12327);
nand U12511 (N_12511,N_12248,N_12332);
nor U12512 (N_12512,N_12251,N_12364);
nor U12513 (N_12513,N_12248,N_12272);
or U12514 (N_12514,N_12225,N_12233);
or U12515 (N_12515,N_12360,N_12317);
nor U12516 (N_12516,N_12207,N_12384);
xor U12517 (N_12517,N_12287,N_12271);
nand U12518 (N_12518,N_12326,N_12308);
nand U12519 (N_12519,N_12317,N_12346);
xor U12520 (N_12520,N_12263,N_12381);
nand U12521 (N_12521,N_12386,N_12262);
nor U12522 (N_12522,N_12336,N_12225);
nand U12523 (N_12523,N_12250,N_12302);
nor U12524 (N_12524,N_12358,N_12213);
nor U12525 (N_12525,N_12333,N_12223);
and U12526 (N_12526,N_12297,N_12290);
and U12527 (N_12527,N_12224,N_12353);
xor U12528 (N_12528,N_12328,N_12252);
nor U12529 (N_12529,N_12257,N_12296);
nand U12530 (N_12530,N_12384,N_12220);
or U12531 (N_12531,N_12322,N_12217);
nand U12532 (N_12532,N_12255,N_12303);
xnor U12533 (N_12533,N_12363,N_12310);
and U12534 (N_12534,N_12375,N_12313);
and U12535 (N_12535,N_12379,N_12290);
and U12536 (N_12536,N_12358,N_12228);
nor U12537 (N_12537,N_12366,N_12377);
or U12538 (N_12538,N_12284,N_12387);
and U12539 (N_12539,N_12374,N_12368);
and U12540 (N_12540,N_12215,N_12243);
and U12541 (N_12541,N_12359,N_12315);
or U12542 (N_12542,N_12200,N_12264);
and U12543 (N_12543,N_12263,N_12299);
xnor U12544 (N_12544,N_12354,N_12267);
or U12545 (N_12545,N_12388,N_12311);
nand U12546 (N_12546,N_12355,N_12232);
or U12547 (N_12547,N_12275,N_12215);
and U12548 (N_12548,N_12216,N_12392);
or U12549 (N_12549,N_12276,N_12308);
xor U12550 (N_12550,N_12360,N_12373);
nor U12551 (N_12551,N_12310,N_12321);
or U12552 (N_12552,N_12370,N_12225);
and U12553 (N_12553,N_12328,N_12259);
and U12554 (N_12554,N_12392,N_12361);
and U12555 (N_12555,N_12304,N_12392);
nand U12556 (N_12556,N_12290,N_12218);
or U12557 (N_12557,N_12244,N_12273);
nor U12558 (N_12558,N_12369,N_12284);
or U12559 (N_12559,N_12350,N_12206);
xnor U12560 (N_12560,N_12398,N_12263);
nand U12561 (N_12561,N_12368,N_12349);
nand U12562 (N_12562,N_12365,N_12288);
and U12563 (N_12563,N_12256,N_12227);
nor U12564 (N_12564,N_12201,N_12367);
nor U12565 (N_12565,N_12218,N_12320);
or U12566 (N_12566,N_12206,N_12341);
or U12567 (N_12567,N_12368,N_12245);
nand U12568 (N_12568,N_12244,N_12265);
and U12569 (N_12569,N_12397,N_12291);
xnor U12570 (N_12570,N_12249,N_12327);
or U12571 (N_12571,N_12272,N_12338);
nand U12572 (N_12572,N_12288,N_12359);
nand U12573 (N_12573,N_12312,N_12384);
and U12574 (N_12574,N_12320,N_12397);
xnor U12575 (N_12575,N_12381,N_12355);
xnor U12576 (N_12576,N_12308,N_12283);
or U12577 (N_12577,N_12285,N_12389);
xor U12578 (N_12578,N_12227,N_12234);
xor U12579 (N_12579,N_12306,N_12377);
nor U12580 (N_12580,N_12326,N_12350);
and U12581 (N_12581,N_12356,N_12217);
nor U12582 (N_12582,N_12204,N_12329);
xnor U12583 (N_12583,N_12354,N_12207);
nand U12584 (N_12584,N_12367,N_12284);
nor U12585 (N_12585,N_12253,N_12307);
xor U12586 (N_12586,N_12260,N_12233);
nor U12587 (N_12587,N_12294,N_12301);
and U12588 (N_12588,N_12201,N_12212);
or U12589 (N_12589,N_12237,N_12212);
nand U12590 (N_12590,N_12329,N_12374);
nand U12591 (N_12591,N_12298,N_12351);
nand U12592 (N_12592,N_12223,N_12288);
xor U12593 (N_12593,N_12347,N_12307);
and U12594 (N_12594,N_12323,N_12294);
nor U12595 (N_12595,N_12263,N_12367);
xnor U12596 (N_12596,N_12211,N_12278);
and U12597 (N_12597,N_12210,N_12260);
or U12598 (N_12598,N_12285,N_12294);
nand U12599 (N_12599,N_12316,N_12276);
nand U12600 (N_12600,N_12502,N_12466);
nor U12601 (N_12601,N_12434,N_12490);
nor U12602 (N_12602,N_12593,N_12562);
xor U12603 (N_12603,N_12585,N_12500);
nor U12604 (N_12604,N_12443,N_12408);
and U12605 (N_12605,N_12468,N_12514);
nand U12606 (N_12606,N_12550,N_12507);
nand U12607 (N_12607,N_12565,N_12511);
nor U12608 (N_12608,N_12481,N_12462);
or U12609 (N_12609,N_12575,N_12523);
and U12610 (N_12610,N_12560,N_12469);
xor U12611 (N_12611,N_12584,N_12437);
or U12612 (N_12612,N_12556,N_12431);
and U12613 (N_12613,N_12541,N_12491);
nor U12614 (N_12614,N_12476,N_12577);
xor U12615 (N_12615,N_12455,N_12538);
nor U12616 (N_12616,N_12516,N_12492);
xnor U12617 (N_12617,N_12495,N_12599);
xnor U12618 (N_12618,N_12445,N_12415);
or U12619 (N_12619,N_12578,N_12501);
and U12620 (N_12620,N_12439,N_12519);
nand U12621 (N_12621,N_12489,N_12509);
nor U12622 (N_12622,N_12450,N_12473);
xor U12623 (N_12623,N_12527,N_12539);
nor U12624 (N_12624,N_12428,N_12544);
and U12625 (N_12625,N_12410,N_12569);
xnor U12626 (N_12626,N_12586,N_12447);
xnor U12627 (N_12627,N_12533,N_12432);
or U12628 (N_12628,N_12493,N_12524);
nor U12629 (N_12629,N_12416,N_12441);
nor U12630 (N_12630,N_12554,N_12411);
nand U12631 (N_12631,N_12496,N_12442);
and U12632 (N_12632,N_12594,N_12465);
xor U12633 (N_12633,N_12448,N_12451);
xor U12634 (N_12634,N_12590,N_12477);
nand U12635 (N_12635,N_12400,N_12510);
xnor U12636 (N_12636,N_12535,N_12540);
or U12637 (N_12637,N_12566,N_12504);
or U12638 (N_12638,N_12479,N_12422);
nand U12639 (N_12639,N_12433,N_12409);
nor U12640 (N_12640,N_12574,N_12440);
nor U12641 (N_12641,N_12454,N_12526);
nand U12642 (N_12642,N_12573,N_12478);
and U12643 (N_12643,N_12474,N_12435);
and U12644 (N_12644,N_12436,N_12555);
or U12645 (N_12645,N_12487,N_12446);
nand U12646 (N_12646,N_12583,N_12475);
or U12647 (N_12647,N_12561,N_12460);
or U12648 (N_12648,N_12417,N_12568);
and U12649 (N_12649,N_12518,N_12513);
nand U12650 (N_12650,N_12484,N_12508);
nand U12651 (N_12651,N_12546,N_12595);
nand U12652 (N_12652,N_12459,N_12425);
nor U12653 (N_12653,N_12532,N_12580);
or U12654 (N_12654,N_12559,N_12461);
xnor U12655 (N_12655,N_12529,N_12517);
xor U12656 (N_12656,N_12592,N_12582);
and U12657 (N_12657,N_12452,N_12429);
or U12658 (N_12658,N_12420,N_12551);
nand U12659 (N_12659,N_12503,N_12401);
nor U12660 (N_12660,N_12545,N_12552);
or U12661 (N_12661,N_12421,N_12571);
and U12662 (N_12662,N_12423,N_12467);
or U12663 (N_12663,N_12537,N_12406);
or U12664 (N_12664,N_12444,N_12515);
xnor U12665 (N_12665,N_12482,N_12542);
nor U12666 (N_12666,N_12506,N_12598);
or U12667 (N_12667,N_12525,N_12570);
nand U12668 (N_12668,N_12472,N_12480);
and U12669 (N_12669,N_12404,N_12453);
xor U12670 (N_12670,N_12426,N_12430);
and U12671 (N_12671,N_12485,N_12499);
and U12672 (N_12672,N_12494,N_12438);
and U12673 (N_12673,N_12531,N_12486);
nand U12674 (N_12674,N_12528,N_12596);
nand U12675 (N_12675,N_12483,N_12557);
and U12676 (N_12676,N_12576,N_12418);
xor U12677 (N_12677,N_12588,N_12405);
xor U12678 (N_12678,N_12464,N_12412);
xnor U12679 (N_12679,N_12597,N_12402);
nor U12680 (N_12680,N_12522,N_12581);
nor U12681 (N_12681,N_12549,N_12458);
nor U12682 (N_12682,N_12520,N_12587);
nand U12683 (N_12683,N_12589,N_12564);
nand U12684 (N_12684,N_12498,N_12512);
or U12685 (N_12685,N_12470,N_12534);
and U12686 (N_12686,N_12548,N_12456);
xnor U12687 (N_12687,N_12427,N_12567);
and U12688 (N_12688,N_12563,N_12553);
nor U12689 (N_12689,N_12407,N_12471);
nand U12690 (N_12690,N_12403,N_12543);
or U12691 (N_12691,N_12547,N_12463);
or U12692 (N_12692,N_12424,N_12530);
nor U12693 (N_12693,N_12497,N_12558);
xor U12694 (N_12694,N_12419,N_12449);
nor U12695 (N_12695,N_12413,N_12488);
xnor U12696 (N_12696,N_12579,N_12591);
nand U12697 (N_12697,N_12521,N_12572);
nand U12698 (N_12698,N_12536,N_12505);
nand U12699 (N_12699,N_12457,N_12414);
nor U12700 (N_12700,N_12587,N_12436);
nor U12701 (N_12701,N_12494,N_12420);
and U12702 (N_12702,N_12497,N_12406);
nor U12703 (N_12703,N_12486,N_12521);
xnor U12704 (N_12704,N_12488,N_12473);
nand U12705 (N_12705,N_12461,N_12459);
nand U12706 (N_12706,N_12542,N_12410);
nand U12707 (N_12707,N_12530,N_12515);
nand U12708 (N_12708,N_12451,N_12456);
or U12709 (N_12709,N_12562,N_12568);
nand U12710 (N_12710,N_12433,N_12532);
nor U12711 (N_12711,N_12510,N_12558);
nand U12712 (N_12712,N_12533,N_12596);
xnor U12713 (N_12713,N_12455,N_12475);
or U12714 (N_12714,N_12439,N_12516);
or U12715 (N_12715,N_12534,N_12471);
nand U12716 (N_12716,N_12475,N_12488);
nand U12717 (N_12717,N_12408,N_12470);
nand U12718 (N_12718,N_12426,N_12418);
nor U12719 (N_12719,N_12499,N_12482);
and U12720 (N_12720,N_12464,N_12465);
nor U12721 (N_12721,N_12412,N_12529);
nand U12722 (N_12722,N_12407,N_12532);
or U12723 (N_12723,N_12447,N_12496);
nor U12724 (N_12724,N_12586,N_12400);
and U12725 (N_12725,N_12512,N_12483);
nor U12726 (N_12726,N_12430,N_12503);
and U12727 (N_12727,N_12508,N_12585);
or U12728 (N_12728,N_12538,N_12584);
and U12729 (N_12729,N_12436,N_12553);
xnor U12730 (N_12730,N_12503,N_12587);
nand U12731 (N_12731,N_12586,N_12532);
xor U12732 (N_12732,N_12502,N_12498);
xnor U12733 (N_12733,N_12470,N_12523);
or U12734 (N_12734,N_12501,N_12465);
nor U12735 (N_12735,N_12559,N_12536);
and U12736 (N_12736,N_12565,N_12506);
and U12737 (N_12737,N_12462,N_12483);
and U12738 (N_12738,N_12530,N_12563);
nand U12739 (N_12739,N_12537,N_12485);
and U12740 (N_12740,N_12414,N_12466);
nor U12741 (N_12741,N_12560,N_12442);
and U12742 (N_12742,N_12552,N_12550);
or U12743 (N_12743,N_12577,N_12414);
xnor U12744 (N_12744,N_12438,N_12410);
nor U12745 (N_12745,N_12531,N_12574);
or U12746 (N_12746,N_12552,N_12444);
nor U12747 (N_12747,N_12552,N_12486);
nor U12748 (N_12748,N_12451,N_12598);
nor U12749 (N_12749,N_12524,N_12451);
or U12750 (N_12750,N_12417,N_12413);
and U12751 (N_12751,N_12457,N_12437);
xnor U12752 (N_12752,N_12428,N_12458);
nor U12753 (N_12753,N_12519,N_12583);
nor U12754 (N_12754,N_12552,N_12408);
or U12755 (N_12755,N_12407,N_12437);
xor U12756 (N_12756,N_12527,N_12532);
and U12757 (N_12757,N_12540,N_12590);
and U12758 (N_12758,N_12512,N_12488);
or U12759 (N_12759,N_12450,N_12471);
xnor U12760 (N_12760,N_12477,N_12559);
or U12761 (N_12761,N_12597,N_12536);
nor U12762 (N_12762,N_12424,N_12543);
xor U12763 (N_12763,N_12418,N_12569);
nor U12764 (N_12764,N_12593,N_12423);
nand U12765 (N_12765,N_12405,N_12431);
or U12766 (N_12766,N_12560,N_12483);
or U12767 (N_12767,N_12593,N_12419);
and U12768 (N_12768,N_12418,N_12502);
or U12769 (N_12769,N_12576,N_12569);
or U12770 (N_12770,N_12536,N_12468);
and U12771 (N_12771,N_12510,N_12594);
xnor U12772 (N_12772,N_12569,N_12501);
and U12773 (N_12773,N_12517,N_12597);
nand U12774 (N_12774,N_12420,N_12431);
xor U12775 (N_12775,N_12458,N_12453);
and U12776 (N_12776,N_12437,N_12469);
xnor U12777 (N_12777,N_12551,N_12476);
nor U12778 (N_12778,N_12403,N_12460);
nor U12779 (N_12779,N_12410,N_12551);
and U12780 (N_12780,N_12520,N_12493);
nor U12781 (N_12781,N_12555,N_12462);
and U12782 (N_12782,N_12472,N_12410);
and U12783 (N_12783,N_12519,N_12553);
or U12784 (N_12784,N_12469,N_12575);
nand U12785 (N_12785,N_12594,N_12473);
xnor U12786 (N_12786,N_12400,N_12563);
nor U12787 (N_12787,N_12441,N_12417);
nand U12788 (N_12788,N_12440,N_12451);
nor U12789 (N_12789,N_12557,N_12523);
nor U12790 (N_12790,N_12512,N_12540);
nor U12791 (N_12791,N_12496,N_12429);
or U12792 (N_12792,N_12556,N_12441);
and U12793 (N_12793,N_12519,N_12592);
and U12794 (N_12794,N_12473,N_12504);
or U12795 (N_12795,N_12511,N_12427);
and U12796 (N_12796,N_12523,N_12445);
nor U12797 (N_12797,N_12448,N_12527);
or U12798 (N_12798,N_12588,N_12507);
or U12799 (N_12799,N_12454,N_12551);
nor U12800 (N_12800,N_12743,N_12727);
nand U12801 (N_12801,N_12677,N_12733);
and U12802 (N_12802,N_12652,N_12780);
nor U12803 (N_12803,N_12617,N_12607);
nand U12804 (N_12804,N_12678,N_12672);
nand U12805 (N_12805,N_12693,N_12746);
nand U12806 (N_12806,N_12694,N_12696);
or U12807 (N_12807,N_12615,N_12647);
nand U12808 (N_12808,N_12620,N_12674);
or U12809 (N_12809,N_12793,N_12742);
nand U12810 (N_12810,N_12682,N_12770);
nand U12811 (N_12811,N_12713,N_12728);
nor U12812 (N_12812,N_12619,N_12723);
xor U12813 (N_12813,N_12639,N_12605);
nand U12814 (N_12814,N_12752,N_12760);
xor U12815 (N_12815,N_12698,N_12641);
and U12816 (N_12816,N_12610,N_12786);
or U12817 (N_12817,N_12642,N_12660);
and U12818 (N_12818,N_12799,N_12627);
and U12819 (N_12819,N_12656,N_12625);
xor U12820 (N_12820,N_12691,N_12649);
xor U12821 (N_12821,N_12797,N_12754);
or U12822 (N_12822,N_12753,N_12791);
nand U12823 (N_12823,N_12784,N_12721);
and U12824 (N_12824,N_12734,N_12681);
xor U12825 (N_12825,N_12790,N_12712);
or U12826 (N_12826,N_12767,N_12796);
and U12827 (N_12827,N_12657,N_12795);
and U12828 (N_12828,N_12729,N_12655);
nor U12829 (N_12829,N_12680,N_12749);
or U12830 (N_12830,N_12769,N_12604);
xnor U12831 (N_12831,N_12776,N_12766);
nor U12832 (N_12832,N_12664,N_12716);
xor U12833 (N_12833,N_12745,N_12690);
xnor U12834 (N_12834,N_12777,N_12707);
nor U12835 (N_12835,N_12756,N_12703);
or U12836 (N_12836,N_12683,N_12788);
xor U12837 (N_12837,N_12798,N_12692);
and U12838 (N_12838,N_12640,N_12667);
nand U12839 (N_12839,N_12789,N_12726);
xor U12840 (N_12840,N_12632,N_12714);
or U12841 (N_12841,N_12779,N_12676);
nor U12842 (N_12842,N_12601,N_12787);
nor U12843 (N_12843,N_12759,N_12653);
or U12844 (N_12844,N_12750,N_12751);
or U12845 (N_12845,N_12725,N_12638);
and U12846 (N_12846,N_12700,N_12773);
nor U12847 (N_12847,N_12774,N_12643);
xnor U12848 (N_12848,N_12663,N_12654);
or U12849 (N_12849,N_12628,N_12706);
and U12850 (N_12850,N_12755,N_12741);
and U12851 (N_12851,N_12704,N_12785);
nor U12852 (N_12852,N_12611,N_12722);
nand U12853 (N_12853,N_12781,N_12624);
or U12854 (N_12854,N_12702,N_12646);
nor U12855 (N_12855,N_12668,N_12603);
nand U12856 (N_12856,N_12618,N_12621);
nand U12857 (N_12857,N_12658,N_12671);
nand U12858 (N_12858,N_12709,N_12695);
nand U12859 (N_12859,N_12765,N_12659);
or U12860 (N_12860,N_12730,N_12768);
nor U12861 (N_12861,N_12630,N_12613);
nor U12862 (N_12862,N_12778,N_12736);
xnor U12863 (N_12863,N_12669,N_12708);
nand U12864 (N_12864,N_12724,N_12710);
xor U12865 (N_12865,N_12636,N_12633);
nand U12866 (N_12866,N_12686,N_12718);
and U12867 (N_12867,N_12701,N_12748);
and U12868 (N_12868,N_12747,N_12685);
xor U12869 (N_12869,N_12622,N_12609);
nor U12870 (N_12870,N_12623,N_12740);
or U12871 (N_12871,N_12662,N_12637);
or U12872 (N_12872,N_12792,N_12757);
xor U12873 (N_12873,N_12635,N_12670);
and U12874 (N_12874,N_12616,N_12744);
and U12875 (N_12875,N_12720,N_12600);
nor U12876 (N_12876,N_12731,N_12711);
xor U12877 (N_12877,N_12634,N_12606);
and U12878 (N_12878,N_12735,N_12665);
nor U12879 (N_12879,N_12761,N_12719);
or U12880 (N_12880,N_12715,N_12661);
nor U12881 (N_12881,N_12644,N_12762);
or U12882 (N_12882,N_12631,N_12697);
or U12883 (N_12883,N_12626,N_12783);
nand U12884 (N_12884,N_12614,N_12772);
nor U12885 (N_12885,N_12782,N_12717);
and U12886 (N_12886,N_12794,N_12732);
nand U12887 (N_12887,N_12764,N_12763);
nor U12888 (N_12888,N_12666,N_12684);
nand U12889 (N_12889,N_12648,N_12699);
xor U12890 (N_12890,N_12629,N_12758);
nand U12891 (N_12891,N_12689,N_12602);
or U12892 (N_12892,N_12687,N_12739);
nand U12893 (N_12893,N_12738,N_12645);
nor U12894 (N_12894,N_12673,N_12771);
and U12895 (N_12895,N_12651,N_12608);
and U12896 (N_12896,N_12650,N_12737);
nand U12897 (N_12897,N_12612,N_12688);
nand U12898 (N_12898,N_12775,N_12679);
or U12899 (N_12899,N_12705,N_12675);
or U12900 (N_12900,N_12739,N_12617);
and U12901 (N_12901,N_12634,N_12696);
or U12902 (N_12902,N_12683,N_12741);
or U12903 (N_12903,N_12753,N_12770);
nor U12904 (N_12904,N_12617,N_12667);
xor U12905 (N_12905,N_12726,N_12631);
nand U12906 (N_12906,N_12618,N_12630);
nor U12907 (N_12907,N_12620,N_12682);
and U12908 (N_12908,N_12677,N_12688);
nor U12909 (N_12909,N_12619,N_12792);
xnor U12910 (N_12910,N_12691,N_12694);
xnor U12911 (N_12911,N_12689,N_12660);
or U12912 (N_12912,N_12763,N_12601);
or U12913 (N_12913,N_12722,N_12657);
xnor U12914 (N_12914,N_12620,N_12658);
and U12915 (N_12915,N_12764,N_12629);
xor U12916 (N_12916,N_12755,N_12712);
nand U12917 (N_12917,N_12765,N_12759);
nor U12918 (N_12918,N_12790,N_12676);
or U12919 (N_12919,N_12662,N_12690);
or U12920 (N_12920,N_12618,N_12739);
nor U12921 (N_12921,N_12731,N_12606);
nor U12922 (N_12922,N_12706,N_12780);
nor U12923 (N_12923,N_12737,N_12649);
or U12924 (N_12924,N_12796,N_12690);
and U12925 (N_12925,N_12654,N_12753);
or U12926 (N_12926,N_12646,N_12784);
nand U12927 (N_12927,N_12733,N_12754);
xnor U12928 (N_12928,N_12720,N_12706);
nor U12929 (N_12929,N_12682,N_12799);
and U12930 (N_12930,N_12632,N_12788);
xnor U12931 (N_12931,N_12607,N_12697);
xor U12932 (N_12932,N_12619,N_12718);
nor U12933 (N_12933,N_12761,N_12775);
and U12934 (N_12934,N_12602,N_12756);
and U12935 (N_12935,N_12741,N_12641);
nand U12936 (N_12936,N_12704,N_12629);
or U12937 (N_12937,N_12778,N_12662);
nor U12938 (N_12938,N_12710,N_12632);
nor U12939 (N_12939,N_12681,N_12650);
nor U12940 (N_12940,N_12768,N_12685);
or U12941 (N_12941,N_12789,N_12678);
nand U12942 (N_12942,N_12620,N_12693);
nand U12943 (N_12943,N_12638,N_12751);
nand U12944 (N_12944,N_12653,N_12769);
nand U12945 (N_12945,N_12738,N_12740);
or U12946 (N_12946,N_12620,N_12703);
nand U12947 (N_12947,N_12661,N_12681);
xnor U12948 (N_12948,N_12777,N_12754);
xnor U12949 (N_12949,N_12760,N_12737);
nand U12950 (N_12950,N_12773,N_12620);
nand U12951 (N_12951,N_12776,N_12774);
and U12952 (N_12952,N_12776,N_12762);
xnor U12953 (N_12953,N_12674,N_12747);
and U12954 (N_12954,N_12659,N_12752);
and U12955 (N_12955,N_12655,N_12669);
and U12956 (N_12956,N_12653,N_12740);
or U12957 (N_12957,N_12795,N_12687);
nor U12958 (N_12958,N_12773,N_12705);
nand U12959 (N_12959,N_12745,N_12707);
nand U12960 (N_12960,N_12771,N_12752);
nand U12961 (N_12961,N_12674,N_12758);
xor U12962 (N_12962,N_12795,N_12650);
xnor U12963 (N_12963,N_12725,N_12675);
nor U12964 (N_12964,N_12651,N_12742);
nor U12965 (N_12965,N_12692,N_12716);
and U12966 (N_12966,N_12705,N_12618);
nand U12967 (N_12967,N_12738,N_12654);
and U12968 (N_12968,N_12657,N_12615);
nor U12969 (N_12969,N_12663,N_12790);
xnor U12970 (N_12970,N_12712,N_12774);
or U12971 (N_12971,N_12698,N_12663);
or U12972 (N_12972,N_12640,N_12628);
and U12973 (N_12973,N_12699,N_12620);
or U12974 (N_12974,N_12693,N_12678);
and U12975 (N_12975,N_12612,N_12711);
nand U12976 (N_12976,N_12624,N_12662);
and U12977 (N_12977,N_12728,N_12633);
nand U12978 (N_12978,N_12753,N_12620);
nand U12979 (N_12979,N_12766,N_12691);
or U12980 (N_12980,N_12770,N_12731);
nor U12981 (N_12981,N_12638,N_12710);
nand U12982 (N_12982,N_12681,N_12613);
and U12983 (N_12983,N_12724,N_12622);
and U12984 (N_12984,N_12796,N_12795);
xor U12985 (N_12985,N_12662,N_12666);
nor U12986 (N_12986,N_12619,N_12683);
or U12987 (N_12987,N_12622,N_12747);
xor U12988 (N_12988,N_12722,N_12791);
or U12989 (N_12989,N_12773,N_12668);
or U12990 (N_12990,N_12799,N_12703);
and U12991 (N_12991,N_12673,N_12691);
or U12992 (N_12992,N_12779,N_12687);
nand U12993 (N_12993,N_12660,N_12723);
nand U12994 (N_12994,N_12768,N_12624);
xor U12995 (N_12995,N_12604,N_12760);
and U12996 (N_12996,N_12733,N_12681);
xnor U12997 (N_12997,N_12634,N_12679);
nand U12998 (N_12998,N_12747,N_12675);
nor U12999 (N_12999,N_12687,N_12768);
xor U13000 (N_13000,N_12876,N_12839);
or U13001 (N_13001,N_12980,N_12954);
nand U13002 (N_13002,N_12874,N_12959);
nor U13003 (N_13003,N_12859,N_12873);
nor U13004 (N_13004,N_12907,N_12871);
and U13005 (N_13005,N_12813,N_12815);
and U13006 (N_13006,N_12885,N_12845);
and U13007 (N_13007,N_12913,N_12819);
and U13008 (N_13008,N_12964,N_12951);
and U13009 (N_13009,N_12831,N_12971);
or U13010 (N_13010,N_12965,N_12854);
nor U13011 (N_13011,N_12957,N_12968);
nand U13012 (N_13012,N_12860,N_12979);
nor U13013 (N_13013,N_12838,N_12992);
nor U13014 (N_13014,N_12802,N_12905);
or U13015 (N_13015,N_12982,N_12881);
nor U13016 (N_13016,N_12823,N_12942);
nand U13017 (N_13017,N_12864,N_12840);
nor U13018 (N_13018,N_12941,N_12808);
nor U13019 (N_13019,N_12843,N_12922);
xnor U13020 (N_13020,N_12812,N_12937);
nor U13021 (N_13021,N_12934,N_12896);
and U13022 (N_13022,N_12899,N_12924);
and U13023 (N_13023,N_12927,N_12912);
xor U13024 (N_13024,N_12949,N_12914);
and U13025 (N_13025,N_12870,N_12825);
or U13026 (N_13026,N_12892,N_12966);
nand U13027 (N_13027,N_12879,N_12939);
nor U13028 (N_13028,N_12895,N_12852);
xnor U13029 (N_13029,N_12901,N_12996);
and U13030 (N_13030,N_12990,N_12920);
or U13031 (N_13031,N_12997,N_12950);
nand U13032 (N_13032,N_12917,N_12890);
xnor U13033 (N_13033,N_12875,N_12850);
nand U13034 (N_13034,N_12811,N_12967);
nor U13035 (N_13035,N_12983,N_12827);
and U13036 (N_13036,N_12987,N_12910);
or U13037 (N_13037,N_12940,N_12932);
and U13038 (N_13038,N_12856,N_12805);
nand U13039 (N_13039,N_12902,N_12801);
and U13040 (N_13040,N_12887,N_12989);
nor U13041 (N_13041,N_12826,N_12869);
or U13042 (N_13042,N_12935,N_12849);
xor U13043 (N_13043,N_12824,N_12981);
or U13044 (N_13044,N_12978,N_12842);
or U13045 (N_13045,N_12810,N_12985);
nor U13046 (N_13046,N_12911,N_12848);
xnor U13047 (N_13047,N_12832,N_12923);
and U13048 (N_13048,N_12961,N_12958);
nor U13049 (N_13049,N_12988,N_12906);
nand U13050 (N_13050,N_12821,N_12977);
xnor U13051 (N_13051,N_12948,N_12956);
xor U13052 (N_13052,N_12867,N_12835);
xor U13053 (N_13053,N_12976,N_12915);
nand U13054 (N_13054,N_12804,N_12883);
nand U13055 (N_13055,N_12991,N_12998);
or U13056 (N_13056,N_12947,N_12900);
nor U13057 (N_13057,N_12818,N_12999);
and U13058 (N_13058,N_12898,N_12943);
xor U13059 (N_13059,N_12903,N_12857);
xor U13060 (N_13060,N_12995,N_12847);
or U13061 (N_13061,N_12833,N_12807);
and U13062 (N_13062,N_12861,N_12878);
nand U13063 (N_13063,N_12863,N_12944);
or U13064 (N_13064,N_12925,N_12970);
and U13065 (N_13065,N_12969,N_12938);
and U13066 (N_13066,N_12928,N_12837);
nor U13067 (N_13067,N_12973,N_12884);
nand U13068 (N_13068,N_12889,N_12929);
and U13069 (N_13069,N_12908,N_12865);
nand U13070 (N_13070,N_12877,N_12933);
and U13071 (N_13071,N_12897,N_12962);
or U13072 (N_13072,N_12829,N_12955);
nand U13073 (N_13073,N_12984,N_12853);
nor U13074 (N_13074,N_12834,N_12974);
xor U13075 (N_13075,N_12930,N_12894);
xor U13076 (N_13076,N_12816,N_12936);
nor U13077 (N_13077,N_12886,N_12891);
or U13078 (N_13078,N_12806,N_12960);
and U13079 (N_13079,N_12904,N_12975);
nor U13080 (N_13080,N_12946,N_12953);
xor U13081 (N_13081,N_12830,N_12909);
nand U13082 (N_13082,N_12800,N_12918);
nor U13083 (N_13083,N_12862,N_12814);
and U13084 (N_13084,N_12921,N_12866);
nor U13085 (N_13085,N_12846,N_12963);
nor U13086 (N_13086,N_12822,N_12993);
nor U13087 (N_13087,N_12916,N_12855);
and U13088 (N_13088,N_12820,N_12836);
xor U13089 (N_13089,N_12882,N_12872);
or U13090 (N_13090,N_12926,N_12803);
nor U13091 (N_13091,N_12828,N_12868);
and U13092 (N_13092,N_12893,N_12994);
and U13093 (N_13093,N_12888,N_12919);
nand U13094 (N_13094,N_12972,N_12880);
nor U13095 (N_13095,N_12851,N_12844);
nor U13096 (N_13096,N_12858,N_12817);
xnor U13097 (N_13097,N_12931,N_12986);
nand U13098 (N_13098,N_12952,N_12945);
and U13099 (N_13099,N_12841,N_12809);
nor U13100 (N_13100,N_12887,N_12866);
and U13101 (N_13101,N_12896,N_12840);
xor U13102 (N_13102,N_12879,N_12840);
and U13103 (N_13103,N_12821,N_12895);
nand U13104 (N_13104,N_12871,N_12821);
xnor U13105 (N_13105,N_12837,N_12977);
nand U13106 (N_13106,N_12988,N_12987);
nand U13107 (N_13107,N_12951,N_12896);
or U13108 (N_13108,N_12814,N_12861);
nand U13109 (N_13109,N_12985,N_12828);
or U13110 (N_13110,N_12812,N_12921);
xnor U13111 (N_13111,N_12850,N_12982);
xor U13112 (N_13112,N_12814,N_12975);
or U13113 (N_13113,N_12974,N_12973);
nor U13114 (N_13114,N_12828,N_12800);
nor U13115 (N_13115,N_12976,N_12811);
nand U13116 (N_13116,N_12919,N_12805);
or U13117 (N_13117,N_12893,N_12970);
xnor U13118 (N_13118,N_12912,N_12848);
nor U13119 (N_13119,N_12941,N_12895);
and U13120 (N_13120,N_12807,N_12944);
nor U13121 (N_13121,N_12837,N_12825);
xor U13122 (N_13122,N_12821,N_12854);
xnor U13123 (N_13123,N_12942,N_12958);
nand U13124 (N_13124,N_12825,N_12820);
xnor U13125 (N_13125,N_12969,N_12843);
and U13126 (N_13126,N_12874,N_12925);
and U13127 (N_13127,N_12987,N_12908);
or U13128 (N_13128,N_12946,N_12930);
nor U13129 (N_13129,N_12816,N_12907);
nor U13130 (N_13130,N_12972,N_12816);
or U13131 (N_13131,N_12997,N_12941);
xnor U13132 (N_13132,N_12966,N_12904);
xor U13133 (N_13133,N_12812,N_12831);
xnor U13134 (N_13134,N_12876,N_12896);
and U13135 (N_13135,N_12957,N_12860);
xor U13136 (N_13136,N_12923,N_12843);
xor U13137 (N_13137,N_12879,N_12994);
xnor U13138 (N_13138,N_12853,N_12937);
nand U13139 (N_13139,N_12873,N_12872);
nand U13140 (N_13140,N_12975,N_12934);
and U13141 (N_13141,N_12801,N_12868);
nor U13142 (N_13142,N_12995,N_12834);
nand U13143 (N_13143,N_12957,N_12917);
and U13144 (N_13144,N_12834,N_12862);
nor U13145 (N_13145,N_12975,N_12862);
or U13146 (N_13146,N_12927,N_12853);
xnor U13147 (N_13147,N_12946,N_12917);
xor U13148 (N_13148,N_12930,N_12818);
nor U13149 (N_13149,N_12855,N_12912);
and U13150 (N_13150,N_12921,N_12829);
and U13151 (N_13151,N_12963,N_12985);
xor U13152 (N_13152,N_12967,N_12971);
nor U13153 (N_13153,N_12964,N_12971);
xnor U13154 (N_13154,N_12954,N_12845);
or U13155 (N_13155,N_12928,N_12909);
nand U13156 (N_13156,N_12884,N_12879);
xnor U13157 (N_13157,N_12862,N_12995);
and U13158 (N_13158,N_12890,N_12985);
xnor U13159 (N_13159,N_12821,N_12987);
xor U13160 (N_13160,N_12960,N_12845);
nand U13161 (N_13161,N_12808,N_12975);
and U13162 (N_13162,N_12916,N_12891);
and U13163 (N_13163,N_12803,N_12918);
nor U13164 (N_13164,N_12995,N_12875);
or U13165 (N_13165,N_12808,N_12911);
nor U13166 (N_13166,N_12935,N_12883);
nor U13167 (N_13167,N_12862,N_12924);
nor U13168 (N_13168,N_12964,N_12893);
or U13169 (N_13169,N_12819,N_12975);
xor U13170 (N_13170,N_12960,N_12987);
nor U13171 (N_13171,N_12969,N_12961);
and U13172 (N_13172,N_12914,N_12966);
nand U13173 (N_13173,N_12889,N_12801);
xor U13174 (N_13174,N_12828,N_12990);
xor U13175 (N_13175,N_12838,N_12849);
nor U13176 (N_13176,N_12952,N_12847);
and U13177 (N_13177,N_12922,N_12860);
and U13178 (N_13178,N_12913,N_12992);
and U13179 (N_13179,N_12872,N_12889);
and U13180 (N_13180,N_12975,N_12893);
nor U13181 (N_13181,N_12900,N_12905);
nor U13182 (N_13182,N_12904,N_12832);
or U13183 (N_13183,N_12814,N_12847);
or U13184 (N_13184,N_12823,N_12893);
or U13185 (N_13185,N_12924,N_12984);
and U13186 (N_13186,N_12852,N_12838);
xnor U13187 (N_13187,N_12916,N_12800);
nand U13188 (N_13188,N_12940,N_12893);
nand U13189 (N_13189,N_12930,N_12956);
nand U13190 (N_13190,N_12870,N_12859);
and U13191 (N_13191,N_12818,N_12848);
nor U13192 (N_13192,N_12990,N_12863);
or U13193 (N_13193,N_12958,N_12896);
and U13194 (N_13194,N_12996,N_12868);
or U13195 (N_13195,N_12966,N_12808);
nand U13196 (N_13196,N_12807,N_12823);
and U13197 (N_13197,N_12819,N_12877);
nor U13198 (N_13198,N_12982,N_12916);
nor U13199 (N_13199,N_12884,N_12855);
or U13200 (N_13200,N_13141,N_13010);
nand U13201 (N_13201,N_13103,N_13131);
nor U13202 (N_13202,N_13048,N_13011);
or U13203 (N_13203,N_13008,N_13106);
or U13204 (N_13204,N_13130,N_13060);
xnor U13205 (N_13205,N_13104,N_13109);
and U13206 (N_13206,N_13152,N_13199);
nor U13207 (N_13207,N_13095,N_13001);
nand U13208 (N_13208,N_13022,N_13140);
xnor U13209 (N_13209,N_13111,N_13188);
xnor U13210 (N_13210,N_13115,N_13143);
and U13211 (N_13211,N_13183,N_13003);
xnor U13212 (N_13212,N_13148,N_13053);
nor U13213 (N_13213,N_13161,N_13071);
xor U13214 (N_13214,N_13006,N_13127);
xor U13215 (N_13215,N_13119,N_13047);
or U13216 (N_13216,N_13097,N_13123);
or U13217 (N_13217,N_13050,N_13040);
xor U13218 (N_13218,N_13007,N_13026);
or U13219 (N_13219,N_13159,N_13155);
or U13220 (N_13220,N_13081,N_13124);
nor U13221 (N_13221,N_13023,N_13128);
and U13222 (N_13222,N_13156,N_13142);
and U13223 (N_13223,N_13002,N_13016);
and U13224 (N_13224,N_13158,N_13019);
nor U13225 (N_13225,N_13033,N_13193);
or U13226 (N_13226,N_13056,N_13042);
or U13227 (N_13227,N_13169,N_13195);
nor U13228 (N_13228,N_13151,N_13014);
or U13229 (N_13229,N_13044,N_13046);
xor U13230 (N_13230,N_13105,N_13135);
nand U13231 (N_13231,N_13015,N_13113);
nand U13232 (N_13232,N_13032,N_13174);
nand U13233 (N_13233,N_13004,N_13062);
nor U13234 (N_13234,N_13031,N_13168);
nand U13235 (N_13235,N_13187,N_13117);
or U13236 (N_13236,N_13136,N_13178);
nand U13237 (N_13237,N_13061,N_13120);
and U13238 (N_13238,N_13122,N_13121);
or U13239 (N_13239,N_13133,N_13021);
or U13240 (N_13240,N_13165,N_13180);
nand U13241 (N_13241,N_13146,N_13052);
and U13242 (N_13242,N_13020,N_13126);
nand U13243 (N_13243,N_13179,N_13073);
nor U13244 (N_13244,N_13074,N_13092);
or U13245 (N_13245,N_13157,N_13079);
and U13246 (N_13246,N_13102,N_13110);
nor U13247 (N_13247,N_13041,N_13139);
or U13248 (N_13248,N_13093,N_13112);
nand U13249 (N_13249,N_13163,N_13177);
nand U13250 (N_13250,N_13116,N_13034);
nand U13251 (N_13251,N_13171,N_13114);
nand U13252 (N_13252,N_13125,N_13024);
xor U13253 (N_13253,N_13153,N_13185);
or U13254 (N_13254,N_13076,N_13077);
nand U13255 (N_13255,N_13025,N_13065);
and U13256 (N_13256,N_13108,N_13134);
nand U13257 (N_13257,N_13086,N_13147);
xor U13258 (N_13258,N_13101,N_13162);
or U13259 (N_13259,N_13000,N_13063);
nor U13260 (N_13260,N_13029,N_13045);
nor U13261 (N_13261,N_13039,N_13096);
or U13262 (N_13262,N_13037,N_13196);
nor U13263 (N_13263,N_13057,N_13099);
or U13264 (N_13264,N_13090,N_13059);
nand U13265 (N_13265,N_13181,N_13160);
nand U13266 (N_13266,N_13089,N_13118);
or U13267 (N_13267,N_13064,N_13184);
and U13268 (N_13268,N_13018,N_13068);
or U13269 (N_13269,N_13154,N_13087);
nor U13270 (N_13270,N_13149,N_13189);
nor U13271 (N_13271,N_13085,N_13055);
nand U13272 (N_13272,N_13192,N_13028);
nand U13273 (N_13273,N_13129,N_13166);
or U13274 (N_13274,N_13080,N_13013);
xnor U13275 (N_13275,N_13138,N_13035);
or U13276 (N_13276,N_13078,N_13091);
and U13277 (N_13277,N_13176,N_13194);
nor U13278 (N_13278,N_13038,N_13175);
xor U13279 (N_13279,N_13107,N_13082);
xor U13280 (N_13280,N_13075,N_13030);
xnor U13281 (N_13281,N_13058,N_13172);
nor U13282 (N_13282,N_13144,N_13186);
or U13283 (N_13283,N_13051,N_13049);
nor U13284 (N_13284,N_13167,N_13191);
or U13285 (N_13285,N_13083,N_13070);
nor U13286 (N_13286,N_13084,N_13054);
nand U13287 (N_13287,N_13150,N_13173);
or U13288 (N_13288,N_13027,N_13098);
nor U13289 (N_13289,N_13164,N_13067);
xnor U13290 (N_13290,N_13197,N_13198);
nand U13291 (N_13291,N_13066,N_13094);
or U13292 (N_13292,N_13190,N_13043);
nor U13293 (N_13293,N_13005,N_13069);
nor U13294 (N_13294,N_13088,N_13012);
nor U13295 (N_13295,N_13145,N_13009);
nor U13296 (N_13296,N_13036,N_13132);
xnor U13297 (N_13297,N_13017,N_13137);
or U13298 (N_13298,N_13170,N_13100);
or U13299 (N_13299,N_13072,N_13182);
and U13300 (N_13300,N_13167,N_13049);
xnor U13301 (N_13301,N_13146,N_13007);
nand U13302 (N_13302,N_13038,N_13067);
nand U13303 (N_13303,N_13018,N_13104);
nor U13304 (N_13304,N_13147,N_13062);
and U13305 (N_13305,N_13165,N_13194);
nor U13306 (N_13306,N_13129,N_13194);
or U13307 (N_13307,N_13009,N_13126);
nand U13308 (N_13308,N_13012,N_13071);
nand U13309 (N_13309,N_13075,N_13029);
nor U13310 (N_13310,N_13192,N_13004);
and U13311 (N_13311,N_13018,N_13148);
or U13312 (N_13312,N_13167,N_13108);
and U13313 (N_13313,N_13132,N_13001);
nor U13314 (N_13314,N_13156,N_13089);
nor U13315 (N_13315,N_13090,N_13094);
xnor U13316 (N_13316,N_13183,N_13178);
xor U13317 (N_13317,N_13194,N_13104);
or U13318 (N_13318,N_13194,N_13175);
xnor U13319 (N_13319,N_13072,N_13020);
and U13320 (N_13320,N_13118,N_13040);
and U13321 (N_13321,N_13171,N_13154);
nor U13322 (N_13322,N_13083,N_13181);
xor U13323 (N_13323,N_13039,N_13170);
and U13324 (N_13324,N_13171,N_13071);
or U13325 (N_13325,N_13019,N_13096);
and U13326 (N_13326,N_13146,N_13127);
xor U13327 (N_13327,N_13104,N_13091);
or U13328 (N_13328,N_13129,N_13118);
nor U13329 (N_13329,N_13100,N_13055);
xnor U13330 (N_13330,N_13180,N_13017);
and U13331 (N_13331,N_13122,N_13117);
and U13332 (N_13332,N_13128,N_13188);
and U13333 (N_13333,N_13178,N_13173);
or U13334 (N_13334,N_13122,N_13158);
nand U13335 (N_13335,N_13175,N_13010);
nor U13336 (N_13336,N_13049,N_13070);
nand U13337 (N_13337,N_13056,N_13039);
nor U13338 (N_13338,N_13121,N_13072);
and U13339 (N_13339,N_13119,N_13049);
nand U13340 (N_13340,N_13042,N_13118);
nor U13341 (N_13341,N_13096,N_13125);
nand U13342 (N_13342,N_13175,N_13123);
nor U13343 (N_13343,N_13029,N_13190);
xnor U13344 (N_13344,N_13086,N_13131);
and U13345 (N_13345,N_13083,N_13031);
nand U13346 (N_13346,N_13197,N_13136);
nand U13347 (N_13347,N_13181,N_13132);
nand U13348 (N_13348,N_13072,N_13012);
nor U13349 (N_13349,N_13104,N_13101);
nor U13350 (N_13350,N_13110,N_13075);
and U13351 (N_13351,N_13058,N_13108);
or U13352 (N_13352,N_13143,N_13007);
xnor U13353 (N_13353,N_13141,N_13076);
xor U13354 (N_13354,N_13191,N_13152);
nand U13355 (N_13355,N_13127,N_13155);
xor U13356 (N_13356,N_13007,N_13075);
xor U13357 (N_13357,N_13081,N_13002);
or U13358 (N_13358,N_13148,N_13175);
xor U13359 (N_13359,N_13153,N_13100);
or U13360 (N_13360,N_13097,N_13164);
nor U13361 (N_13361,N_13139,N_13163);
and U13362 (N_13362,N_13188,N_13032);
xor U13363 (N_13363,N_13198,N_13144);
and U13364 (N_13364,N_13046,N_13167);
nor U13365 (N_13365,N_13036,N_13185);
and U13366 (N_13366,N_13121,N_13045);
nor U13367 (N_13367,N_13062,N_13049);
nand U13368 (N_13368,N_13017,N_13116);
or U13369 (N_13369,N_13092,N_13188);
nor U13370 (N_13370,N_13087,N_13195);
nor U13371 (N_13371,N_13075,N_13197);
xnor U13372 (N_13372,N_13028,N_13180);
and U13373 (N_13373,N_13037,N_13150);
nor U13374 (N_13374,N_13056,N_13168);
xnor U13375 (N_13375,N_13028,N_13143);
and U13376 (N_13376,N_13007,N_13006);
and U13377 (N_13377,N_13158,N_13064);
or U13378 (N_13378,N_13105,N_13117);
and U13379 (N_13379,N_13133,N_13035);
xor U13380 (N_13380,N_13008,N_13117);
or U13381 (N_13381,N_13019,N_13012);
nor U13382 (N_13382,N_13103,N_13197);
nor U13383 (N_13383,N_13106,N_13149);
nor U13384 (N_13384,N_13146,N_13149);
xor U13385 (N_13385,N_13175,N_13126);
xor U13386 (N_13386,N_13013,N_13119);
and U13387 (N_13387,N_13008,N_13183);
and U13388 (N_13388,N_13054,N_13087);
and U13389 (N_13389,N_13143,N_13088);
xnor U13390 (N_13390,N_13034,N_13078);
xor U13391 (N_13391,N_13179,N_13064);
or U13392 (N_13392,N_13166,N_13009);
or U13393 (N_13393,N_13050,N_13033);
nand U13394 (N_13394,N_13119,N_13104);
or U13395 (N_13395,N_13041,N_13181);
nor U13396 (N_13396,N_13141,N_13073);
and U13397 (N_13397,N_13106,N_13163);
nand U13398 (N_13398,N_13102,N_13090);
xor U13399 (N_13399,N_13001,N_13045);
nor U13400 (N_13400,N_13224,N_13373);
and U13401 (N_13401,N_13230,N_13304);
and U13402 (N_13402,N_13292,N_13335);
xor U13403 (N_13403,N_13225,N_13353);
nand U13404 (N_13404,N_13347,N_13382);
and U13405 (N_13405,N_13360,N_13247);
or U13406 (N_13406,N_13348,N_13388);
nor U13407 (N_13407,N_13208,N_13262);
xor U13408 (N_13408,N_13368,N_13263);
nor U13409 (N_13409,N_13333,N_13301);
nor U13410 (N_13410,N_13258,N_13370);
nor U13411 (N_13411,N_13234,N_13255);
xor U13412 (N_13412,N_13290,N_13318);
and U13413 (N_13413,N_13351,N_13300);
xnor U13414 (N_13414,N_13244,N_13387);
or U13415 (N_13415,N_13238,N_13286);
or U13416 (N_13416,N_13264,N_13338);
xnor U13417 (N_13417,N_13236,N_13210);
nand U13418 (N_13418,N_13248,N_13352);
nor U13419 (N_13419,N_13294,N_13223);
or U13420 (N_13420,N_13362,N_13345);
or U13421 (N_13421,N_13203,N_13392);
nor U13422 (N_13422,N_13201,N_13291);
and U13423 (N_13423,N_13363,N_13334);
and U13424 (N_13424,N_13349,N_13232);
nor U13425 (N_13425,N_13396,N_13213);
or U13426 (N_13426,N_13252,N_13274);
and U13427 (N_13427,N_13245,N_13293);
nor U13428 (N_13428,N_13273,N_13383);
and U13429 (N_13429,N_13356,N_13280);
nand U13430 (N_13430,N_13271,N_13250);
xor U13431 (N_13431,N_13384,N_13266);
or U13432 (N_13432,N_13342,N_13249);
or U13433 (N_13433,N_13346,N_13319);
xor U13434 (N_13434,N_13235,N_13207);
nor U13435 (N_13435,N_13254,N_13355);
and U13436 (N_13436,N_13251,N_13379);
and U13437 (N_13437,N_13246,N_13243);
or U13438 (N_13438,N_13265,N_13381);
xor U13439 (N_13439,N_13200,N_13276);
nor U13440 (N_13440,N_13378,N_13323);
nor U13441 (N_13441,N_13209,N_13313);
and U13442 (N_13442,N_13284,N_13305);
nor U13443 (N_13443,N_13233,N_13226);
or U13444 (N_13444,N_13214,N_13311);
xnor U13445 (N_13445,N_13205,N_13310);
nand U13446 (N_13446,N_13202,N_13211);
nor U13447 (N_13447,N_13241,N_13339);
nand U13448 (N_13448,N_13315,N_13242);
nor U13449 (N_13449,N_13228,N_13330);
xor U13450 (N_13450,N_13302,N_13324);
or U13451 (N_13451,N_13219,N_13227);
and U13452 (N_13452,N_13393,N_13218);
and U13453 (N_13453,N_13344,N_13260);
nand U13454 (N_13454,N_13328,N_13395);
nor U13455 (N_13455,N_13297,N_13391);
nor U13456 (N_13456,N_13350,N_13336);
nor U13457 (N_13457,N_13231,N_13364);
xnor U13458 (N_13458,N_13303,N_13288);
or U13459 (N_13459,N_13332,N_13341);
nor U13460 (N_13460,N_13340,N_13268);
nor U13461 (N_13461,N_13282,N_13216);
xor U13462 (N_13462,N_13220,N_13212);
and U13463 (N_13463,N_13277,N_13237);
nand U13464 (N_13464,N_13374,N_13257);
xor U13465 (N_13465,N_13390,N_13240);
nor U13466 (N_13466,N_13278,N_13279);
xnor U13467 (N_13467,N_13361,N_13222);
nor U13468 (N_13468,N_13283,N_13397);
or U13469 (N_13469,N_13316,N_13299);
nor U13470 (N_13470,N_13398,N_13357);
nand U13471 (N_13471,N_13317,N_13326);
and U13472 (N_13472,N_13308,N_13371);
xnor U13473 (N_13473,N_13256,N_13285);
and U13474 (N_13474,N_13359,N_13221);
xor U13475 (N_13475,N_13306,N_13259);
or U13476 (N_13476,N_13296,N_13295);
and U13477 (N_13477,N_13327,N_13372);
or U13478 (N_13478,N_13298,N_13272);
nor U13479 (N_13479,N_13369,N_13329);
or U13480 (N_13480,N_13358,N_13386);
xor U13481 (N_13481,N_13399,N_13275);
nand U13482 (N_13482,N_13309,N_13385);
xnor U13483 (N_13483,N_13354,N_13239);
nor U13484 (N_13484,N_13322,N_13267);
nand U13485 (N_13485,N_13376,N_13307);
nand U13486 (N_13486,N_13366,N_13281);
nand U13487 (N_13487,N_13343,N_13380);
nor U13488 (N_13488,N_13289,N_13270);
or U13489 (N_13489,N_13287,N_13206);
nor U13490 (N_13490,N_13337,N_13325);
nor U13491 (N_13491,N_13261,N_13377);
and U13492 (N_13492,N_13269,N_13253);
and U13493 (N_13493,N_13389,N_13320);
and U13494 (N_13494,N_13217,N_13312);
nor U13495 (N_13495,N_13367,N_13365);
nand U13496 (N_13496,N_13375,N_13331);
xnor U13497 (N_13497,N_13204,N_13321);
nor U13498 (N_13498,N_13215,N_13394);
or U13499 (N_13499,N_13314,N_13229);
or U13500 (N_13500,N_13339,N_13279);
xor U13501 (N_13501,N_13206,N_13224);
and U13502 (N_13502,N_13363,N_13378);
nand U13503 (N_13503,N_13251,N_13344);
and U13504 (N_13504,N_13238,N_13330);
or U13505 (N_13505,N_13225,N_13379);
and U13506 (N_13506,N_13249,N_13320);
and U13507 (N_13507,N_13321,N_13226);
xnor U13508 (N_13508,N_13261,N_13307);
nand U13509 (N_13509,N_13397,N_13218);
xor U13510 (N_13510,N_13281,N_13354);
and U13511 (N_13511,N_13218,N_13395);
and U13512 (N_13512,N_13286,N_13314);
nor U13513 (N_13513,N_13233,N_13302);
nor U13514 (N_13514,N_13263,N_13212);
nor U13515 (N_13515,N_13291,N_13380);
nand U13516 (N_13516,N_13237,N_13310);
nand U13517 (N_13517,N_13351,N_13253);
or U13518 (N_13518,N_13347,N_13358);
and U13519 (N_13519,N_13357,N_13337);
nand U13520 (N_13520,N_13266,N_13355);
xnor U13521 (N_13521,N_13344,N_13388);
nand U13522 (N_13522,N_13383,N_13342);
xor U13523 (N_13523,N_13340,N_13377);
or U13524 (N_13524,N_13380,N_13349);
xnor U13525 (N_13525,N_13254,N_13259);
or U13526 (N_13526,N_13209,N_13347);
or U13527 (N_13527,N_13202,N_13361);
xor U13528 (N_13528,N_13372,N_13386);
nand U13529 (N_13529,N_13358,N_13332);
nor U13530 (N_13530,N_13280,N_13271);
nor U13531 (N_13531,N_13201,N_13373);
nor U13532 (N_13532,N_13308,N_13391);
or U13533 (N_13533,N_13306,N_13305);
and U13534 (N_13534,N_13223,N_13261);
nand U13535 (N_13535,N_13202,N_13386);
xor U13536 (N_13536,N_13267,N_13260);
nand U13537 (N_13537,N_13348,N_13363);
or U13538 (N_13538,N_13365,N_13258);
xnor U13539 (N_13539,N_13318,N_13357);
and U13540 (N_13540,N_13331,N_13319);
and U13541 (N_13541,N_13342,N_13293);
and U13542 (N_13542,N_13200,N_13205);
xnor U13543 (N_13543,N_13395,N_13388);
nand U13544 (N_13544,N_13394,N_13201);
nand U13545 (N_13545,N_13327,N_13208);
or U13546 (N_13546,N_13395,N_13217);
xnor U13547 (N_13547,N_13274,N_13325);
or U13548 (N_13548,N_13297,N_13296);
xor U13549 (N_13549,N_13399,N_13308);
and U13550 (N_13550,N_13236,N_13322);
nor U13551 (N_13551,N_13281,N_13217);
and U13552 (N_13552,N_13394,N_13395);
xor U13553 (N_13553,N_13253,N_13358);
or U13554 (N_13554,N_13205,N_13309);
nor U13555 (N_13555,N_13330,N_13203);
or U13556 (N_13556,N_13391,N_13270);
xor U13557 (N_13557,N_13283,N_13336);
or U13558 (N_13558,N_13351,N_13297);
xnor U13559 (N_13559,N_13235,N_13285);
nor U13560 (N_13560,N_13313,N_13282);
nor U13561 (N_13561,N_13392,N_13371);
xnor U13562 (N_13562,N_13297,N_13243);
xnor U13563 (N_13563,N_13301,N_13296);
and U13564 (N_13564,N_13284,N_13299);
nand U13565 (N_13565,N_13360,N_13346);
or U13566 (N_13566,N_13235,N_13292);
and U13567 (N_13567,N_13297,N_13220);
nand U13568 (N_13568,N_13213,N_13399);
and U13569 (N_13569,N_13210,N_13378);
nor U13570 (N_13570,N_13283,N_13398);
xnor U13571 (N_13571,N_13350,N_13243);
and U13572 (N_13572,N_13396,N_13275);
xor U13573 (N_13573,N_13247,N_13202);
nand U13574 (N_13574,N_13212,N_13293);
xor U13575 (N_13575,N_13340,N_13330);
xnor U13576 (N_13576,N_13382,N_13216);
nor U13577 (N_13577,N_13330,N_13229);
xor U13578 (N_13578,N_13316,N_13338);
xnor U13579 (N_13579,N_13310,N_13207);
xnor U13580 (N_13580,N_13252,N_13272);
nand U13581 (N_13581,N_13399,N_13222);
nand U13582 (N_13582,N_13264,N_13306);
nor U13583 (N_13583,N_13267,N_13380);
nor U13584 (N_13584,N_13353,N_13376);
or U13585 (N_13585,N_13299,N_13249);
nor U13586 (N_13586,N_13233,N_13342);
and U13587 (N_13587,N_13255,N_13296);
or U13588 (N_13588,N_13360,N_13236);
or U13589 (N_13589,N_13380,N_13249);
and U13590 (N_13590,N_13232,N_13350);
xnor U13591 (N_13591,N_13376,N_13396);
xor U13592 (N_13592,N_13236,N_13324);
nand U13593 (N_13593,N_13322,N_13283);
xor U13594 (N_13594,N_13201,N_13206);
xnor U13595 (N_13595,N_13216,N_13358);
nand U13596 (N_13596,N_13267,N_13382);
nand U13597 (N_13597,N_13236,N_13356);
or U13598 (N_13598,N_13231,N_13240);
and U13599 (N_13599,N_13201,N_13315);
nor U13600 (N_13600,N_13416,N_13572);
or U13601 (N_13601,N_13408,N_13483);
xor U13602 (N_13602,N_13420,N_13475);
or U13603 (N_13603,N_13595,N_13488);
xor U13604 (N_13604,N_13584,N_13497);
nand U13605 (N_13605,N_13507,N_13557);
nor U13606 (N_13606,N_13533,N_13496);
xnor U13607 (N_13607,N_13444,N_13433);
or U13608 (N_13608,N_13410,N_13553);
and U13609 (N_13609,N_13511,N_13450);
nor U13610 (N_13610,N_13565,N_13413);
nand U13611 (N_13611,N_13494,N_13529);
or U13612 (N_13612,N_13449,N_13447);
or U13613 (N_13613,N_13527,N_13521);
nand U13614 (N_13614,N_13472,N_13574);
nand U13615 (N_13615,N_13436,N_13591);
and U13616 (N_13616,N_13575,N_13482);
and U13617 (N_13617,N_13474,N_13440);
or U13618 (N_13618,N_13461,N_13490);
nor U13619 (N_13619,N_13517,N_13510);
and U13620 (N_13620,N_13592,N_13484);
xnor U13621 (N_13621,N_13438,N_13405);
xnor U13622 (N_13622,N_13593,N_13566);
xnor U13623 (N_13623,N_13470,N_13554);
or U13624 (N_13624,N_13456,N_13513);
xnor U13625 (N_13625,N_13401,N_13495);
nand U13626 (N_13626,N_13538,N_13442);
and U13627 (N_13627,N_13498,N_13535);
or U13628 (N_13628,N_13578,N_13561);
xor U13629 (N_13629,N_13418,N_13515);
nand U13630 (N_13630,N_13589,N_13501);
nor U13631 (N_13631,N_13468,N_13465);
nand U13632 (N_13632,N_13568,N_13471);
or U13633 (N_13633,N_13429,N_13516);
and U13634 (N_13634,N_13500,N_13487);
nand U13635 (N_13635,N_13427,N_13506);
xor U13636 (N_13636,N_13512,N_13426);
nand U13637 (N_13637,N_13469,N_13534);
nor U13638 (N_13638,N_13467,N_13424);
nand U13639 (N_13639,N_13419,N_13505);
and U13640 (N_13640,N_13514,N_13459);
nand U13641 (N_13641,N_13528,N_13588);
xnor U13642 (N_13642,N_13556,N_13551);
nor U13643 (N_13643,N_13422,N_13525);
xnor U13644 (N_13644,N_13569,N_13567);
nand U13645 (N_13645,N_13428,N_13499);
and U13646 (N_13646,N_13432,N_13540);
and U13647 (N_13647,N_13555,N_13594);
nand U13648 (N_13648,N_13587,N_13582);
and U13649 (N_13649,N_13403,N_13570);
nor U13650 (N_13650,N_13400,N_13489);
nor U13651 (N_13651,N_13446,N_13583);
or U13652 (N_13652,N_13542,N_13455);
nand U13653 (N_13653,N_13537,N_13431);
and U13654 (N_13654,N_13562,N_13421);
and U13655 (N_13655,N_13462,N_13573);
nor U13656 (N_13656,N_13434,N_13522);
nand U13657 (N_13657,N_13579,N_13563);
nor U13658 (N_13658,N_13463,N_13406);
nand U13659 (N_13659,N_13597,N_13430);
nor U13660 (N_13660,N_13451,N_13415);
nor U13661 (N_13661,N_13544,N_13473);
xnor U13662 (N_13662,N_13435,N_13523);
or U13663 (N_13663,N_13454,N_13585);
or U13664 (N_13664,N_13576,N_13485);
nor U13665 (N_13665,N_13480,N_13508);
or U13666 (N_13666,N_13407,N_13425);
nor U13667 (N_13667,N_13486,N_13479);
and U13668 (N_13668,N_13504,N_13599);
or U13669 (N_13669,N_13423,N_13560);
and U13670 (N_13670,N_13448,N_13526);
or U13671 (N_13671,N_13550,N_13466);
xor U13672 (N_13672,N_13549,N_13437);
xnor U13673 (N_13673,N_13546,N_13552);
nand U13674 (N_13674,N_13590,N_13477);
nand U13675 (N_13675,N_13414,N_13453);
or U13676 (N_13676,N_13491,N_13586);
nand U13677 (N_13677,N_13458,N_13564);
and U13678 (N_13678,N_13598,N_13492);
nor U13679 (N_13679,N_13404,N_13409);
and U13680 (N_13680,N_13443,N_13417);
nor U13681 (N_13681,N_13532,N_13539);
nand U13682 (N_13682,N_13439,N_13445);
xnor U13683 (N_13683,N_13536,N_13452);
nor U13684 (N_13684,N_13460,N_13411);
or U13685 (N_13685,N_13531,N_13524);
nor U13686 (N_13686,N_13476,N_13559);
and U13687 (N_13687,N_13478,N_13545);
or U13688 (N_13688,N_13518,N_13503);
xor U13689 (N_13689,N_13502,N_13547);
nand U13690 (N_13690,N_13571,N_13493);
xor U13691 (N_13691,N_13581,N_13530);
xnor U13692 (N_13692,N_13519,N_13402);
nor U13693 (N_13693,N_13580,N_13577);
xnor U13694 (N_13694,N_13548,N_13441);
and U13695 (N_13695,N_13457,N_13543);
or U13696 (N_13696,N_13520,N_13464);
or U13697 (N_13697,N_13558,N_13412);
and U13698 (N_13698,N_13481,N_13596);
or U13699 (N_13699,N_13509,N_13541);
and U13700 (N_13700,N_13548,N_13528);
nor U13701 (N_13701,N_13594,N_13540);
and U13702 (N_13702,N_13589,N_13416);
and U13703 (N_13703,N_13589,N_13499);
nor U13704 (N_13704,N_13545,N_13514);
nand U13705 (N_13705,N_13448,N_13589);
nand U13706 (N_13706,N_13418,N_13495);
xnor U13707 (N_13707,N_13447,N_13535);
or U13708 (N_13708,N_13486,N_13445);
and U13709 (N_13709,N_13418,N_13474);
and U13710 (N_13710,N_13586,N_13409);
xor U13711 (N_13711,N_13451,N_13592);
xor U13712 (N_13712,N_13588,N_13510);
xnor U13713 (N_13713,N_13441,N_13532);
or U13714 (N_13714,N_13423,N_13554);
or U13715 (N_13715,N_13459,N_13451);
nand U13716 (N_13716,N_13552,N_13535);
xor U13717 (N_13717,N_13573,N_13444);
or U13718 (N_13718,N_13555,N_13406);
or U13719 (N_13719,N_13499,N_13404);
nand U13720 (N_13720,N_13538,N_13571);
nor U13721 (N_13721,N_13559,N_13512);
xnor U13722 (N_13722,N_13450,N_13401);
nor U13723 (N_13723,N_13525,N_13499);
nand U13724 (N_13724,N_13462,N_13429);
or U13725 (N_13725,N_13438,N_13446);
or U13726 (N_13726,N_13488,N_13518);
nor U13727 (N_13727,N_13403,N_13564);
or U13728 (N_13728,N_13508,N_13587);
and U13729 (N_13729,N_13508,N_13454);
nand U13730 (N_13730,N_13543,N_13429);
and U13731 (N_13731,N_13542,N_13537);
nor U13732 (N_13732,N_13502,N_13486);
and U13733 (N_13733,N_13449,N_13445);
xor U13734 (N_13734,N_13592,N_13431);
or U13735 (N_13735,N_13551,N_13583);
or U13736 (N_13736,N_13444,N_13578);
nand U13737 (N_13737,N_13562,N_13551);
xor U13738 (N_13738,N_13466,N_13591);
xnor U13739 (N_13739,N_13563,N_13491);
and U13740 (N_13740,N_13455,N_13599);
or U13741 (N_13741,N_13540,N_13453);
xnor U13742 (N_13742,N_13518,N_13442);
xor U13743 (N_13743,N_13400,N_13432);
or U13744 (N_13744,N_13577,N_13474);
xnor U13745 (N_13745,N_13467,N_13580);
or U13746 (N_13746,N_13404,N_13541);
xor U13747 (N_13747,N_13535,N_13471);
or U13748 (N_13748,N_13477,N_13512);
xnor U13749 (N_13749,N_13430,N_13421);
and U13750 (N_13750,N_13461,N_13587);
nor U13751 (N_13751,N_13496,N_13551);
nor U13752 (N_13752,N_13520,N_13409);
nand U13753 (N_13753,N_13409,N_13504);
nor U13754 (N_13754,N_13407,N_13520);
nand U13755 (N_13755,N_13454,N_13485);
nand U13756 (N_13756,N_13432,N_13485);
nand U13757 (N_13757,N_13530,N_13491);
and U13758 (N_13758,N_13516,N_13584);
nor U13759 (N_13759,N_13449,N_13502);
nor U13760 (N_13760,N_13514,N_13555);
or U13761 (N_13761,N_13555,N_13567);
or U13762 (N_13762,N_13553,N_13552);
and U13763 (N_13763,N_13599,N_13501);
and U13764 (N_13764,N_13489,N_13542);
xnor U13765 (N_13765,N_13450,N_13552);
nor U13766 (N_13766,N_13468,N_13574);
nor U13767 (N_13767,N_13435,N_13462);
nand U13768 (N_13768,N_13434,N_13500);
nand U13769 (N_13769,N_13403,N_13554);
nand U13770 (N_13770,N_13565,N_13463);
or U13771 (N_13771,N_13447,N_13405);
xnor U13772 (N_13772,N_13508,N_13427);
or U13773 (N_13773,N_13563,N_13452);
nor U13774 (N_13774,N_13552,N_13581);
xor U13775 (N_13775,N_13406,N_13552);
or U13776 (N_13776,N_13428,N_13423);
xnor U13777 (N_13777,N_13475,N_13556);
nor U13778 (N_13778,N_13595,N_13465);
and U13779 (N_13779,N_13461,N_13473);
xor U13780 (N_13780,N_13424,N_13494);
nor U13781 (N_13781,N_13574,N_13579);
or U13782 (N_13782,N_13472,N_13582);
and U13783 (N_13783,N_13555,N_13589);
or U13784 (N_13784,N_13532,N_13586);
nor U13785 (N_13785,N_13541,N_13442);
and U13786 (N_13786,N_13494,N_13428);
xor U13787 (N_13787,N_13551,N_13483);
nor U13788 (N_13788,N_13556,N_13549);
and U13789 (N_13789,N_13449,N_13532);
nor U13790 (N_13790,N_13405,N_13403);
nor U13791 (N_13791,N_13434,N_13431);
nand U13792 (N_13792,N_13580,N_13544);
or U13793 (N_13793,N_13458,N_13584);
or U13794 (N_13794,N_13468,N_13448);
nand U13795 (N_13795,N_13536,N_13455);
or U13796 (N_13796,N_13453,N_13590);
or U13797 (N_13797,N_13566,N_13533);
xor U13798 (N_13798,N_13583,N_13488);
and U13799 (N_13799,N_13551,N_13541);
xnor U13800 (N_13800,N_13794,N_13780);
nand U13801 (N_13801,N_13620,N_13611);
xor U13802 (N_13802,N_13745,N_13621);
and U13803 (N_13803,N_13716,N_13618);
xor U13804 (N_13804,N_13791,N_13732);
and U13805 (N_13805,N_13685,N_13725);
and U13806 (N_13806,N_13761,N_13624);
and U13807 (N_13807,N_13613,N_13634);
and U13808 (N_13808,N_13792,N_13753);
xor U13809 (N_13809,N_13765,N_13667);
nand U13810 (N_13810,N_13734,N_13680);
nand U13811 (N_13811,N_13743,N_13692);
nand U13812 (N_13812,N_13718,N_13741);
xnor U13813 (N_13813,N_13612,N_13642);
nand U13814 (N_13814,N_13783,N_13683);
nand U13815 (N_13815,N_13700,N_13747);
nand U13816 (N_13816,N_13788,N_13755);
or U13817 (N_13817,N_13651,N_13632);
nor U13818 (N_13818,N_13629,N_13724);
nand U13819 (N_13819,N_13695,N_13711);
nor U13820 (N_13820,N_13616,N_13748);
nand U13821 (N_13821,N_13735,N_13701);
nor U13822 (N_13822,N_13602,N_13675);
or U13823 (N_13823,N_13709,N_13609);
and U13824 (N_13824,N_13715,N_13666);
nand U13825 (N_13825,N_13723,N_13657);
and U13826 (N_13826,N_13712,N_13687);
nor U13827 (N_13827,N_13622,N_13610);
nand U13828 (N_13828,N_13654,N_13628);
xor U13829 (N_13829,N_13759,N_13698);
and U13830 (N_13830,N_13647,N_13713);
nor U13831 (N_13831,N_13779,N_13643);
and U13832 (N_13832,N_13708,N_13636);
and U13833 (N_13833,N_13603,N_13659);
nor U13834 (N_13834,N_13789,N_13793);
nand U13835 (N_13835,N_13689,N_13728);
or U13836 (N_13836,N_13742,N_13778);
and U13837 (N_13837,N_13664,N_13645);
or U13838 (N_13838,N_13627,N_13601);
nand U13839 (N_13839,N_13650,N_13691);
and U13840 (N_13840,N_13644,N_13750);
nand U13841 (N_13841,N_13669,N_13688);
nand U13842 (N_13842,N_13782,N_13752);
nand U13843 (N_13843,N_13768,N_13690);
or U13844 (N_13844,N_13606,N_13662);
and U13845 (N_13845,N_13717,N_13762);
and U13846 (N_13846,N_13677,N_13638);
nor U13847 (N_13847,N_13736,N_13703);
nor U13848 (N_13848,N_13721,N_13615);
or U13849 (N_13849,N_13740,N_13770);
xor U13850 (N_13850,N_13674,N_13710);
nand U13851 (N_13851,N_13614,N_13678);
and U13852 (N_13852,N_13658,N_13605);
and U13853 (N_13853,N_13733,N_13769);
nor U13854 (N_13854,N_13767,N_13707);
or U13855 (N_13855,N_13699,N_13705);
or U13856 (N_13856,N_13697,N_13676);
xnor U13857 (N_13857,N_13704,N_13630);
or U13858 (N_13858,N_13639,N_13682);
and U13859 (N_13859,N_13775,N_13652);
nand U13860 (N_13860,N_13608,N_13739);
nor U13861 (N_13861,N_13623,N_13649);
nand U13862 (N_13862,N_13781,N_13702);
xnor U13863 (N_13863,N_13774,N_13773);
nand U13864 (N_13864,N_13787,N_13684);
nor U13865 (N_13865,N_13686,N_13796);
and U13866 (N_13866,N_13681,N_13635);
nor U13867 (N_13867,N_13648,N_13798);
nand U13868 (N_13868,N_13777,N_13668);
nand U13869 (N_13869,N_13729,N_13731);
or U13870 (N_13870,N_13646,N_13764);
nand U13871 (N_13871,N_13637,N_13784);
or U13872 (N_13872,N_13799,N_13633);
and U13873 (N_13873,N_13726,N_13617);
or U13874 (N_13874,N_13757,N_13641);
nor U13875 (N_13875,N_13653,N_13604);
or U13876 (N_13876,N_13673,N_13786);
nand U13877 (N_13877,N_13719,N_13727);
nor U13878 (N_13878,N_13776,N_13640);
and U13879 (N_13879,N_13671,N_13631);
and U13880 (N_13880,N_13760,N_13797);
and U13881 (N_13881,N_13714,N_13720);
nand U13882 (N_13882,N_13607,N_13670);
or U13883 (N_13883,N_13771,N_13672);
or U13884 (N_13884,N_13763,N_13758);
nand U13885 (N_13885,N_13751,N_13694);
nor U13886 (N_13886,N_13600,N_13656);
xnor U13887 (N_13887,N_13679,N_13785);
or U13888 (N_13888,N_13619,N_13756);
or U13889 (N_13889,N_13696,N_13766);
xor U13890 (N_13890,N_13655,N_13663);
xor U13891 (N_13891,N_13738,N_13795);
nor U13892 (N_13892,N_13722,N_13665);
and U13893 (N_13893,N_13706,N_13737);
nand U13894 (N_13894,N_13693,N_13790);
nand U13895 (N_13895,N_13661,N_13772);
nand U13896 (N_13896,N_13626,N_13744);
nand U13897 (N_13897,N_13730,N_13625);
nand U13898 (N_13898,N_13660,N_13754);
and U13899 (N_13899,N_13746,N_13749);
nand U13900 (N_13900,N_13606,N_13677);
nor U13901 (N_13901,N_13643,N_13765);
xnor U13902 (N_13902,N_13602,N_13760);
or U13903 (N_13903,N_13716,N_13723);
xnor U13904 (N_13904,N_13638,N_13715);
nand U13905 (N_13905,N_13691,N_13716);
nand U13906 (N_13906,N_13685,N_13741);
nor U13907 (N_13907,N_13726,N_13716);
nand U13908 (N_13908,N_13724,N_13720);
xnor U13909 (N_13909,N_13657,N_13720);
and U13910 (N_13910,N_13628,N_13610);
nor U13911 (N_13911,N_13682,N_13715);
nor U13912 (N_13912,N_13743,N_13640);
or U13913 (N_13913,N_13689,N_13639);
or U13914 (N_13914,N_13775,N_13641);
and U13915 (N_13915,N_13799,N_13774);
nand U13916 (N_13916,N_13719,N_13791);
and U13917 (N_13917,N_13672,N_13695);
xnor U13918 (N_13918,N_13719,N_13661);
xnor U13919 (N_13919,N_13679,N_13676);
nand U13920 (N_13920,N_13798,N_13692);
xnor U13921 (N_13921,N_13689,N_13675);
xnor U13922 (N_13922,N_13633,N_13674);
xnor U13923 (N_13923,N_13678,N_13717);
nand U13924 (N_13924,N_13777,N_13771);
and U13925 (N_13925,N_13699,N_13608);
xnor U13926 (N_13926,N_13736,N_13618);
nand U13927 (N_13927,N_13754,N_13638);
nor U13928 (N_13928,N_13693,N_13788);
and U13929 (N_13929,N_13709,N_13672);
nor U13930 (N_13930,N_13782,N_13746);
nand U13931 (N_13931,N_13765,N_13700);
xor U13932 (N_13932,N_13734,N_13656);
nand U13933 (N_13933,N_13728,N_13600);
nand U13934 (N_13934,N_13636,N_13707);
nor U13935 (N_13935,N_13652,N_13689);
nand U13936 (N_13936,N_13636,N_13706);
or U13937 (N_13937,N_13719,N_13797);
nor U13938 (N_13938,N_13624,N_13703);
nor U13939 (N_13939,N_13677,N_13666);
nand U13940 (N_13940,N_13789,N_13688);
or U13941 (N_13941,N_13764,N_13769);
xnor U13942 (N_13942,N_13696,N_13754);
xor U13943 (N_13943,N_13658,N_13647);
or U13944 (N_13944,N_13625,N_13691);
xnor U13945 (N_13945,N_13743,N_13624);
and U13946 (N_13946,N_13743,N_13720);
or U13947 (N_13947,N_13623,N_13644);
or U13948 (N_13948,N_13702,N_13727);
xor U13949 (N_13949,N_13735,N_13677);
nand U13950 (N_13950,N_13713,N_13603);
nor U13951 (N_13951,N_13708,N_13682);
nand U13952 (N_13952,N_13715,N_13620);
or U13953 (N_13953,N_13754,N_13618);
nand U13954 (N_13954,N_13604,N_13623);
and U13955 (N_13955,N_13725,N_13681);
nand U13956 (N_13956,N_13604,N_13703);
and U13957 (N_13957,N_13705,N_13694);
or U13958 (N_13958,N_13745,N_13770);
nand U13959 (N_13959,N_13669,N_13782);
xor U13960 (N_13960,N_13722,N_13600);
nor U13961 (N_13961,N_13666,N_13686);
xnor U13962 (N_13962,N_13645,N_13792);
or U13963 (N_13963,N_13653,N_13630);
xor U13964 (N_13964,N_13716,N_13735);
or U13965 (N_13965,N_13764,N_13658);
nand U13966 (N_13966,N_13737,N_13634);
or U13967 (N_13967,N_13711,N_13688);
nor U13968 (N_13968,N_13624,N_13641);
or U13969 (N_13969,N_13691,N_13743);
nand U13970 (N_13970,N_13705,N_13686);
or U13971 (N_13971,N_13624,N_13681);
or U13972 (N_13972,N_13751,N_13737);
nand U13973 (N_13973,N_13617,N_13787);
and U13974 (N_13974,N_13667,N_13779);
nand U13975 (N_13975,N_13703,N_13615);
nor U13976 (N_13976,N_13653,N_13721);
nand U13977 (N_13977,N_13653,N_13795);
nand U13978 (N_13978,N_13689,N_13765);
or U13979 (N_13979,N_13694,N_13636);
nand U13980 (N_13980,N_13651,N_13628);
or U13981 (N_13981,N_13648,N_13695);
and U13982 (N_13982,N_13698,N_13678);
and U13983 (N_13983,N_13655,N_13727);
xor U13984 (N_13984,N_13763,N_13749);
or U13985 (N_13985,N_13738,N_13787);
xnor U13986 (N_13986,N_13729,N_13631);
nor U13987 (N_13987,N_13655,N_13642);
nand U13988 (N_13988,N_13603,N_13614);
xor U13989 (N_13989,N_13603,N_13766);
nor U13990 (N_13990,N_13683,N_13706);
xnor U13991 (N_13991,N_13782,N_13713);
nand U13992 (N_13992,N_13713,N_13609);
or U13993 (N_13993,N_13643,N_13727);
xnor U13994 (N_13994,N_13719,N_13790);
nor U13995 (N_13995,N_13697,N_13641);
or U13996 (N_13996,N_13722,N_13658);
xor U13997 (N_13997,N_13734,N_13622);
nor U13998 (N_13998,N_13654,N_13637);
and U13999 (N_13999,N_13601,N_13618);
xor U14000 (N_14000,N_13964,N_13879);
xor U14001 (N_14001,N_13908,N_13862);
nand U14002 (N_14002,N_13940,N_13913);
and U14003 (N_14003,N_13969,N_13825);
xnor U14004 (N_14004,N_13980,N_13943);
nor U14005 (N_14005,N_13998,N_13993);
and U14006 (N_14006,N_13840,N_13925);
nand U14007 (N_14007,N_13972,N_13977);
or U14008 (N_14008,N_13822,N_13893);
and U14009 (N_14009,N_13952,N_13990);
xor U14010 (N_14010,N_13898,N_13882);
or U14011 (N_14011,N_13987,N_13911);
nand U14012 (N_14012,N_13803,N_13880);
and U14013 (N_14013,N_13931,N_13810);
and U14014 (N_14014,N_13957,N_13890);
or U14015 (N_14015,N_13858,N_13863);
nor U14016 (N_14016,N_13874,N_13923);
xor U14017 (N_14017,N_13839,N_13995);
xnor U14018 (N_14018,N_13820,N_13988);
or U14019 (N_14019,N_13849,N_13801);
nand U14020 (N_14020,N_13836,N_13832);
nand U14021 (N_14021,N_13846,N_13919);
and U14022 (N_14022,N_13864,N_13888);
nor U14023 (N_14023,N_13920,N_13973);
xor U14024 (N_14024,N_13907,N_13866);
and U14025 (N_14025,N_13837,N_13905);
nor U14026 (N_14026,N_13891,N_13806);
nor U14027 (N_14027,N_13855,N_13968);
nor U14028 (N_14028,N_13851,N_13966);
nor U14029 (N_14029,N_13805,N_13902);
nand U14030 (N_14030,N_13928,N_13946);
nand U14031 (N_14031,N_13815,N_13814);
and U14032 (N_14032,N_13953,N_13934);
nor U14033 (N_14033,N_13950,N_13848);
or U14034 (N_14034,N_13826,N_13892);
or U14035 (N_14035,N_13812,N_13813);
nor U14036 (N_14036,N_13816,N_13944);
nor U14037 (N_14037,N_13949,N_13999);
nor U14038 (N_14038,N_13835,N_13938);
nand U14039 (N_14039,N_13854,N_13906);
nor U14040 (N_14040,N_13904,N_13819);
and U14041 (N_14041,N_13917,N_13914);
xnor U14042 (N_14042,N_13942,N_13915);
nand U14043 (N_14043,N_13982,N_13885);
nor U14044 (N_14044,N_13827,N_13965);
or U14045 (N_14045,N_13833,N_13881);
and U14046 (N_14046,N_13896,N_13901);
xnor U14047 (N_14047,N_13875,N_13900);
nor U14048 (N_14048,N_13985,N_13852);
and U14049 (N_14049,N_13870,N_13824);
or U14050 (N_14050,N_13984,N_13847);
or U14051 (N_14051,N_13935,N_13918);
and U14052 (N_14052,N_13960,N_13959);
xor U14053 (N_14053,N_13830,N_13996);
and U14054 (N_14054,N_13844,N_13926);
xnor U14055 (N_14055,N_13948,N_13976);
nand U14056 (N_14056,N_13922,N_13994);
nand U14057 (N_14057,N_13916,N_13842);
nand U14058 (N_14058,N_13967,N_13895);
nand U14059 (N_14059,N_13981,N_13989);
nand U14060 (N_14060,N_13997,N_13877);
nand U14061 (N_14061,N_13829,N_13886);
or U14062 (N_14062,N_13856,N_13838);
xor U14063 (N_14063,N_13834,N_13868);
or U14064 (N_14064,N_13889,N_13903);
nand U14065 (N_14065,N_13894,N_13831);
or U14066 (N_14066,N_13921,N_13865);
xnor U14067 (N_14067,N_13927,N_13954);
nand U14068 (N_14068,N_13843,N_13991);
or U14069 (N_14069,N_13850,N_13929);
or U14070 (N_14070,N_13817,N_13800);
or U14071 (N_14071,N_13932,N_13802);
xor U14072 (N_14072,N_13956,N_13986);
nand U14073 (N_14073,N_13930,N_13808);
nor U14074 (N_14074,N_13878,N_13978);
nor U14075 (N_14075,N_13897,N_13962);
nor U14076 (N_14076,N_13909,N_13945);
and U14077 (N_14077,N_13807,N_13947);
or U14078 (N_14078,N_13818,N_13869);
nor U14079 (N_14079,N_13961,N_13955);
xor U14080 (N_14080,N_13939,N_13859);
or U14081 (N_14081,N_13867,N_13887);
or U14082 (N_14082,N_13883,N_13963);
and U14083 (N_14083,N_13884,N_13841);
nand U14084 (N_14084,N_13958,N_13861);
nor U14085 (N_14085,N_13936,N_13974);
and U14086 (N_14086,N_13971,N_13857);
and U14087 (N_14087,N_13809,N_13823);
or U14088 (N_14088,N_13811,N_13992);
and U14089 (N_14089,N_13983,N_13845);
and U14090 (N_14090,N_13873,N_13860);
nor U14091 (N_14091,N_13951,N_13912);
nor U14092 (N_14092,N_13828,N_13871);
or U14093 (N_14093,N_13970,N_13924);
or U14094 (N_14094,N_13804,N_13910);
xor U14095 (N_14095,N_13975,N_13876);
nor U14096 (N_14096,N_13979,N_13853);
xor U14097 (N_14097,N_13937,N_13941);
nand U14098 (N_14098,N_13899,N_13872);
nor U14099 (N_14099,N_13933,N_13821);
nand U14100 (N_14100,N_13952,N_13992);
and U14101 (N_14101,N_13830,N_13849);
and U14102 (N_14102,N_13833,N_13944);
and U14103 (N_14103,N_13846,N_13982);
nand U14104 (N_14104,N_13919,N_13850);
and U14105 (N_14105,N_13812,N_13895);
nor U14106 (N_14106,N_13896,N_13866);
and U14107 (N_14107,N_13981,N_13957);
and U14108 (N_14108,N_13801,N_13871);
or U14109 (N_14109,N_13975,N_13801);
xnor U14110 (N_14110,N_13842,N_13972);
or U14111 (N_14111,N_13837,N_13937);
nand U14112 (N_14112,N_13966,N_13898);
and U14113 (N_14113,N_13887,N_13840);
nand U14114 (N_14114,N_13959,N_13908);
or U14115 (N_14115,N_13878,N_13811);
or U14116 (N_14116,N_13880,N_13926);
and U14117 (N_14117,N_13917,N_13865);
and U14118 (N_14118,N_13858,N_13987);
nor U14119 (N_14119,N_13983,N_13812);
nor U14120 (N_14120,N_13862,N_13953);
or U14121 (N_14121,N_13953,N_13809);
nor U14122 (N_14122,N_13985,N_13899);
or U14123 (N_14123,N_13835,N_13870);
and U14124 (N_14124,N_13811,N_13909);
or U14125 (N_14125,N_13878,N_13868);
nand U14126 (N_14126,N_13984,N_13863);
nand U14127 (N_14127,N_13933,N_13819);
or U14128 (N_14128,N_13836,N_13962);
nand U14129 (N_14129,N_13923,N_13820);
xor U14130 (N_14130,N_13853,N_13877);
and U14131 (N_14131,N_13852,N_13973);
or U14132 (N_14132,N_13850,N_13827);
nand U14133 (N_14133,N_13951,N_13880);
or U14134 (N_14134,N_13976,N_13978);
and U14135 (N_14135,N_13969,N_13837);
and U14136 (N_14136,N_13919,N_13924);
nor U14137 (N_14137,N_13906,N_13951);
xor U14138 (N_14138,N_13803,N_13996);
nor U14139 (N_14139,N_13854,N_13929);
xnor U14140 (N_14140,N_13884,N_13966);
and U14141 (N_14141,N_13860,N_13997);
nand U14142 (N_14142,N_13888,N_13973);
nand U14143 (N_14143,N_13951,N_13839);
or U14144 (N_14144,N_13851,N_13879);
nor U14145 (N_14145,N_13943,N_13858);
nor U14146 (N_14146,N_13901,N_13894);
or U14147 (N_14147,N_13972,N_13872);
and U14148 (N_14148,N_13922,N_13871);
or U14149 (N_14149,N_13811,N_13957);
nor U14150 (N_14150,N_13820,N_13885);
or U14151 (N_14151,N_13921,N_13935);
xor U14152 (N_14152,N_13882,N_13965);
nor U14153 (N_14153,N_13940,N_13829);
and U14154 (N_14154,N_13940,N_13883);
nand U14155 (N_14155,N_13998,N_13930);
xor U14156 (N_14156,N_13924,N_13949);
nand U14157 (N_14157,N_13825,N_13868);
nor U14158 (N_14158,N_13801,N_13878);
xnor U14159 (N_14159,N_13918,N_13801);
nand U14160 (N_14160,N_13997,N_13951);
or U14161 (N_14161,N_13806,N_13863);
and U14162 (N_14162,N_13884,N_13941);
xor U14163 (N_14163,N_13994,N_13928);
nor U14164 (N_14164,N_13988,N_13807);
nor U14165 (N_14165,N_13937,N_13844);
or U14166 (N_14166,N_13854,N_13998);
nand U14167 (N_14167,N_13947,N_13906);
and U14168 (N_14168,N_13843,N_13850);
nand U14169 (N_14169,N_13815,N_13840);
nor U14170 (N_14170,N_13915,N_13931);
nor U14171 (N_14171,N_13830,N_13840);
nor U14172 (N_14172,N_13959,N_13969);
nor U14173 (N_14173,N_13928,N_13903);
nor U14174 (N_14174,N_13829,N_13916);
or U14175 (N_14175,N_13962,N_13881);
xnor U14176 (N_14176,N_13890,N_13944);
and U14177 (N_14177,N_13928,N_13965);
nor U14178 (N_14178,N_13867,N_13847);
xor U14179 (N_14179,N_13834,N_13996);
or U14180 (N_14180,N_13968,N_13942);
nand U14181 (N_14181,N_13840,N_13875);
and U14182 (N_14182,N_13819,N_13804);
nand U14183 (N_14183,N_13863,N_13895);
or U14184 (N_14184,N_13972,N_13840);
xor U14185 (N_14185,N_13958,N_13952);
and U14186 (N_14186,N_13818,N_13912);
xor U14187 (N_14187,N_13954,N_13994);
nor U14188 (N_14188,N_13841,N_13891);
nor U14189 (N_14189,N_13908,N_13899);
nand U14190 (N_14190,N_13884,N_13991);
and U14191 (N_14191,N_13816,N_13803);
nand U14192 (N_14192,N_13884,N_13800);
xnor U14193 (N_14193,N_13916,N_13806);
xnor U14194 (N_14194,N_13820,N_13927);
and U14195 (N_14195,N_13881,N_13874);
nand U14196 (N_14196,N_13838,N_13893);
and U14197 (N_14197,N_13945,N_13830);
and U14198 (N_14198,N_13855,N_13854);
nand U14199 (N_14199,N_13963,N_13860);
or U14200 (N_14200,N_14100,N_14170);
and U14201 (N_14201,N_14037,N_14092);
or U14202 (N_14202,N_14117,N_14042);
nor U14203 (N_14203,N_14013,N_14127);
and U14204 (N_14204,N_14122,N_14104);
nand U14205 (N_14205,N_14128,N_14192);
or U14206 (N_14206,N_14019,N_14008);
and U14207 (N_14207,N_14103,N_14082);
xnor U14208 (N_14208,N_14155,N_14083);
or U14209 (N_14209,N_14084,N_14167);
xnor U14210 (N_14210,N_14041,N_14156);
nor U14211 (N_14211,N_14190,N_14069);
nor U14212 (N_14212,N_14081,N_14057);
or U14213 (N_14213,N_14040,N_14126);
and U14214 (N_14214,N_14185,N_14134);
xnor U14215 (N_14215,N_14178,N_14006);
and U14216 (N_14216,N_14036,N_14067);
or U14217 (N_14217,N_14063,N_14091);
or U14218 (N_14218,N_14166,N_14053);
nor U14219 (N_14219,N_14137,N_14193);
nand U14220 (N_14220,N_14133,N_14094);
nand U14221 (N_14221,N_14175,N_14055);
or U14222 (N_14222,N_14197,N_14097);
or U14223 (N_14223,N_14050,N_14187);
xor U14224 (N_14224,N_14182,N_14096);
xnor U14225 (N_14225,N_14088,N_14076);
nand U14226 (N_14226,N_14020,N_14003);
xor U14227 (N_14227,N_14065,N_14043);
xor U14228 (N_14228,N_14184,N_14132);
nor U14229 (N_14229,N_14007,N_14147);
nor U14230 (N_14230,N_14004,N_14143);
or U14231 (N_14231,N_14047,N_14110);
nor U14232 (N_14232,N_14161,N_14164);
xor U14233 (N_14233,N_14171,N_14017);
or U14234 (N_14234,N_14108,N_14099);
or U14235 (N_14235,N_14179,N_14168);
nor U14236 (N_14236,N_14027,N_14044);
nor U14237 (N_14237,N_14048,N_14118);
nor U14238 (N_14238,N_14089,N_14148);
nor U14239 (N_14239,N_14086,N_14066);
and U14240 (N_14240,N_14150,N_14105);
nand U14241 (N_14241,N_14123,N_14060);
and U14242 (N_14242,N_14079,N_14174);
xor U14243 (N_14243,N_14029,N_14199);
nor U14244 (N_14244,N_14090,N_14030);
nor U14245 (N_14245,N_14095,N_14068);
and U14246 (N_14246,N_14102,N_14162);
nand U14247 (N_14247,N_14176,N_14141);
and U14248 (N_14248,N_14074,N_14101);
nand U14249 (N_14249,N_14125,N_14151);
and U14250 (N_14250,N_14183,N_14152);
nor U14251 (N_14251,N_14106,N_14080);
nand U14252 (N_14252,N_14158,N_14181);
or U14253 (N_14253,N_14034,N_14028);
nand U14254 (N_14254,N_14139,N_14136);
xor U14255 (N_14255,N_14111,N_14109);
nand U14256 (N_14256,N_14116,N_14075);
or U14257 (N_14257,N_14054,N_14191);
nor U14258 (N_14258,N_14130,N_14014);
nor U14259 (N_14259,N_14023,N_14138);
nand U14260 (N_14260,N_14188,N_14159);
nor U14261 (N_14261,N_14085,N_14169);
or U14262 (N_14262,N_14153,N_14021);
and U14263 (N_14263,N_14000,N_14035);
xnor U14264 (N_14264,N_14015,N_14002);
and U14265 (N_14265,N_14196,N_14010);
xnor U14266 (N_14266,N_14038,N_14142);
xor U14267 (N_14267,N_14011,N_14033);
xnor U14268 (N_14268,N_14064,N_14098);
or U14269 (N_14269,N_14077,N_14059);
nor U14270 (N_14270,N_14012,N_14195);
and U14271 (N_14271,N_14049,N_14058);
and U14272 (N_14272,N_14124,N_14112);
or U14273 (N_14273,N_14121,N_14018);
and U14274 (N_14274,N_14045,N_14039);
or U14275 (N_14275,N_14157,N_14165);
xnor U14276 (N_14276,N_14071,N_14078);
xor U14277 (N_14277,N_14072,N_14131);
xnor U14278 (N_14278,N_14189,N_14140);
nand U14279 (N_14279,N_14149,N_14144);
and U14280 (N_14280,N_14146,N_14070);
nor U14281 (N_14281,N_14001,N_14186);
nand U14282 (N_14282,N_14135,N_14032);
and U14283 (N_14283,N_14107,N_14163);
nand U14284 (N_14284,N_14160,N_14087);
or U14285 (N_14285,N_14114,N_14026);
nand U14286 (N_14286,N_14145,N_14052);
or U14287 (N_14287,N_14073,N_14046);
or U14288 (N_14288,N_14056,N_14198);
nor U14289 (N_14289,N_14129,N_14051);
nor U14290 (N_14290,N_14120,N_14113);
nand U14291 (N_14291,N_14024,N_14173);
nor U14292 (N_14292,N_14031,N_14061);
or U14293 (N_14293,N_14180,N_14115);
nand U14294 (N_14294,N_14154,N_14062);
and U14295 (N_14295,N_14093,N_14022);
nand U14296 (N_14296,N_14005,N_14194);
or U14297 (N_14297,N_14172,N_14016);
xor U14298 (N_14298,N_14119,N_14009);
and U14299 (N_14299,N_14025,N_14177);
nand U14300 (N_14300,N_14085,N_14048);
xnor U14301 (N_14301,N_14081,N_14103);
nand U14302 (N_14302,N_14098,N_14074);
and U14303 (N_14303,N_14002,N_14058);
nor U14304 (N_14304,N_14029,N_14154);
nor U14305 (N_14305,N_14094,N_14002);
or U14306 (N_14306,N_14108,N_14127);
nand U14307 (N_14307,N_14164,N_14037);
nor U14308 (N_14308,N_14021,N_14147);
xor U14309 (N_14309,N_14172,N_14199);
and U14310 (N_14310,N_14092,N_14022);
nand U14311 (N_14311,N_14102,N_14087);
and U14312 (N_14312,N_14198,N_14087);
or U14313 (N_14313,N_14106,N_14190);
nor U14314 (N_14314,N_14088,N_14121);
nand U14315 (N_14315,N_14127,N_14085);
or U14316 (N_14316,N_14107,N_14036);
xnor U14317 (N_14317,N_14177,N_14084);
nor U14318 (N_14318,N_14005,N_14041);
xnor U14319 (N_14319,N_14026,N_14087);
nand U14320 (N_14320,N_14113,N_14013);
xnor U14321 (N_14321,N_14149,N_14034);
xor U14322 (N_14322,N_14131,N_14182);
or U14323 (N_14323,N_14115,N_14121);
nor U14324 (N_14324,N_14106,N_14052);
nor U14325 (N_14325,N_14017,N_14198);
or U14326 (N_14326,N_14004,N_14044);
and U14327 (N_14327,N_14135,N_14004);
or U14328 (N_14328,N_14165,N_14024);
nand U14329 (N_14329,N_14191,N_14154);
or U14330 (N_14330,N_14189,N_14149);
or U14331 (N_14331,N_14124,N_14061);
nor U14332 (N_14332,N_14121,N_14180);
and U14333 (N_14333,N_14139,N_14170);
nor U14334 (N_14334,N_14014,N_14069);
xnor U14335 (N_14335,N_14175,N_14047);
nand U14336 (N_14336,N_14146,N_14199);
or U14337 (N_14337,N_14004,N_14028);
nor U14338 (N_14338,N_14061,N_14043);
nor U14339 (N_14339,N_14076,N_14171);
or U14340 (N_14340,N_14138,N_14180);
nand U14341 (N_14341,N_14095,N_14115);
and U14342 (N_14342,N_14040,N_14117);
nor U14343 (N_14343,N_14158,N_14045);
and U14344 (N_14344,N_14153,N_14147);
or U14345 (N_14345,N_14023,N_14038);
nor U14346 (N_14346,N_14150,N_14163);
nand U14347 (N_14347,N_14187,N_14139);
nand U14348 (N_14348,N_14007,N_14088);
or U14349 (N_14349,N_14041,N_14148);
and U14350 (N_14350,N_14062,N_14145);
xnor U14351 (N_14351,N_14198,N_14140);
nand U14352 (N_14352,N_14015,N_14018);
nor U14353 (N_14353,N_14150,N_14115);
or U14354 (N_14354,N_14139,N_14134);
nand U14355 (N_14355,N_14089,N_14171);
or U14356 (N_14356,N_14147,N_14027);
and U14357 (N_14357,N_14187,N_14096);
nor U14358 (N_14358,N_14024,N_14169);
or U14359 (N_14359,N_14064,N_14198);
and U14360 (N_14360,N_14007,N_14048);
or U14361 (N_14361,N_14195,N_14091);
nand U14362 (N_14362,N_14063,N_14067);
nand U14363 (N_14363,N_14145,N_14106);
and U14364 (N_14364,N_14144,N_14100);
nand U14365 (N_14365,N_14168,N_14196);
and U14366 (N_14366,N_14197,N_14154);
or U14367 (N_14367,N_14184,N_14143);
nor U14368 (N_14368,N_14135,N_14015);
nor U14369 (N_14369,N_14022,N_14041);
and U14370 (N_14370,N_14156,N_14166);
nand U14371 (N_14371,N_14161,N_14095);
nand U14372 (N_14372,N_14025,N_14061);
xor U14373 (N_14373,N_14031,N_14092);
or U14374 (N_14374,N_14102,N_14050);
or U14375 (N_14375,N_14145,N_14070);
and U14376 (N_14376,N_14007,N_14036);
nand U14377 (N_14377,N_14181,N_14030);
nor U14378 (N_14378,N_14059,N_14115);
or U14379 (N_14379,N_14108,N_14146);
xor U14380 (N_14380,N_14017,N_14196);
nor U14381 (N_14381,N_14019,N_14012);
xnor U14382 (N_14382,N_14135,N_14055);
nand U14383 (N_14383,N_14105,N_14148);
xnor U14384 (N_14384,N_14055,N_14179);
or U14385 (N_14385,N_14061,N_14004);
and U14386 (N_14386,N_14134,N_14081);
or U14387 (N_14387,N_14063,N_14116);
or U14388 (N_14388,N_14006,N_14175);
nand U14389 (N_14389,N_14124,N_14069);
nor U14390 (N_14390,N_14068,N_14182);
nor U14391 (N_14391,N_14009,N_14160);
nand U14392 (N_14392,N_14128,N_14014);
and U14393 (N_14393,N_14083,N_14041);
and U14394 (N_14394,N_14153,N_14125);
nor U14395 (N_14395,N_14143,N_14181);
xor U14396 (N_14396,N_14015,N_14055);
xor U14397 (N_14397,N_14158,N_14006);
and U14398 (N_14398,N_14064,N_14061);
nor U14399 (N_14399,N_14166,N_14133);
nand U14400 (N_14400,N_14228,N_14285);
xor U14401 (N_14401,N_14377,N_14303);
and U14402 (N_14402,N_14233,N_14288);
and U14403 (N_14403,N_14304,N_14336);
and U14404 (N_14404,N_14300,N_14396);
nor U14405 (N_14405,N_14337,N_14324);
nor U14406 (N_14406,N_14229,N_14232);
xor U14407 (N_14407,N_14399,N_14217);
nand U14408 (N_14408,N_14338,N_14390);
or U14409 (N_14409,N_14247,N_14392);
nor U14410 (N_14410,N_14287,N_14207);
xor U14411 (N_14411,N_14249,N_14383);
and U14412 (N_14412,N_14208,N_14226);
or U14413 (N_14413,N_14279,N_14277);
or U14414 (N_14414,N_14298,N_14393);
or U14415 (N_14415,N_14345,N_14366);
and U14416 (N_14416,N_14314,N_14294);
or U14417 (N_14417,N_14375,N_14351);
nor U14418 (N_14418,N_14237,N_14251);
nor U14419 (N_14419,N_14268,N_14267);
or U14420 (N_14420,N_14310,N_14344);
nor U14421 (N_14421,N_14335,N_14203);
or U14422 (N_14422,N_14348,N_14382);
or U14423 (N_14423,N_14308,N_14329);
xor U14424 (N_14424,N_14376,N_14224);
nor U14425 (N_14425,N_14302,N_14241);
xnor U14426 (N_14426,N_14385,N_14256);
xor U14427 (N_14427,N_14284,N_14215);
xor U14428 (N_14428,N_14397,N_14373);
or U14429 (N_14429,N_14391,N_14363);
or U14430 (N_14430,N_14331,N_14272);
nand U14431 (N_14431,N_14210,N_14227);
xnor U14432 (N_14432,N_14225,N_14289);
nand U14433 (N_14433,N_14269,N_14212);
and U14434 (N_14434,N_14368,N_14263);
xnor U14435 (N_14435,N_14386,N_14291);
or U14436 (N_14436,N_14326,N_14311);
xnor U14437 (N_14437,N_14305,N_14301);
and U14438 (N_14438,N_14262,N_14250);
xor U14439 (N_14439,N_14221,N_14293);
nor U14440 (N_14440,N_14266,N_14299);
nor U14441 (N_14441,N_14209,N_14222);
nor U14442 (N_14442,N_14248,N_14264);
nor U14443 (N_14443,N_14357,N_14352);
or U14444 (N_14444,N_14290,N_14327);
or U14445 (N_14445,N_14297,N_14276);
and U14446 (N_14446,N_14309,N_14218);
nor U14447 (N_14447,N_14394,N_14312);
nand U14448 (N_14448,N_14253,N_14339);
nor U14449 (N_14449,N_14332,N_14204);
and U14450 (N_14450,N_14260,N_14340);
nor U14451 (N_14451,N_14246,N_14216);
nand U14452 (N_14452,N_14349,N_14273);
and U14453 (N_14453,N_14346,N_14259);
xor U14454 (N_14454,N_14236,N_14343);
and U14455 (N_14455,N_14323,N_14231);
xor U14456 (N_14456,N_14261,N_14234);
and U14457 (N_14457,N_14270,N_14361);
and U14458 (N_14458,N_14370,N_14325);
nand U14459 (N_14459,N_14313,N_14318);
xor U14460 (N_14460,N_14358,N_14282);
nor U14461 (N_14461,N_14239,N_14374);
and U14462 (N_14462,N_14200,N_14362);
nand U14463 (N_14463,N_14317,N_14372);
and U14464 (N_14464,N_14205,N_14381);
nor U14465 (N_14465,N_14350,N_14320);
nand U14466 (N_14466,N_14292,N_14342);
nor U14467 (N_14467,N_14354,N_14254);
nor U14468 (N_14468,N_14322,N_14258);
xnor U14469 (N_14469,N_14265,N_14388);
xnor U14470 (N_14470,N_14206,N_14295);
nor U14471 (N_14471,N_14243,N_14379);
and U14472 (N_14472,N_14334,N_14235);
nor U14473 (N_14473,N_14306,N_14271);
nor U14474 (N_14474,N_14353,N_14389);
or U14475 (N_14475,N_14307,N_14380);
or U14476 (N_14476,N_14367,N_14280);
or U14477 (N_14477,N_14201,N_14378);
nor U14478 (N_14478,N_14330,N_14321);
and U14479 (N_14479,N_14283,N_14355);
xnor U14480 (N_14480,N_14245,N_14213);
or U14481 (N_14481,N_14341,N_14274);
nor U14482 (N_14482,N_14316,N_14364);
nand U14483 (N_14483,N_14244,N_14238);
nor U14484 (N_14484,N_14333,N_14359);
and U14485 (N_14485,N_14219,N_14369);
and U14486 (N_14486,N_14275,N_14387);
and U14487 (N_14487,N_14356,N_14257);
and U14488 (N_14488,N_14252,N_14319);
or U14489 (N_14489,N_14371,N_14384);
xor U14490 (N_14490,N_14296,N_14230);
nor U14491 (N_14491,N_14347,N_14202);
xor U14492 (N_14492,N_14242,N_14220);
and U14493 (N_14493,N_14240,N_14315);
nand U14494 (N_14494,N_14395,N_14278);
or U14495 (N_14495,N_14214,N_14398);
and U14496 (N_14496,N_14328,N_14286);
nand U14497 (N_14497,N_14281,N_14255);
and U14498 (N_14498,N_14365,N_14360);
nand U14499 (N_14499,N_14211,N_14223);
and U14500 (N_14500,N_14291,N_14233);
or U14501 (N_14501,N_14311,N_14254);
or U14502 (N_14502,N_14313,N_14347);
and U14503 (N_14503,N_14316,N_14349);
nand U14504 (N_14504,N_14315,N_14335);
nor U14505 (N_14505,N_14333,N_14346);
nand U14506 (N_14506,N_14286,N_14237);
and U14507 (N_14507,N_14357,N_14267);
nand U14508 (N_14508,N_14360,N_14203);
nor U14509 (N_14509,N_14202,N_14283);
and U14510 (N_14510,N_14280,N_14357);
and U14511 (N_14511,N_14366,N_14378);
nand U14512 (N_14512,N_14339,N_14231);
nand U14513 (N_14513,N_14381,N_14225);
nand U14514 (N_14514,N_14334,N_14268);
nand U14515 (N_14515,N_14203,N_14316);
and U14516 (N_14516,N_14323,N_14253);
nor U14517 (N_14517,N_14289,N_14221);
and U14518 (N_14518,N_14214,N_14284);
xor U14519 (N_14519,N_14268,N_14395);
or U14520 (N_14520,N_14255,N_14320);
nor U14521 (N_14521,N_14352,N_14202);
nand U14522 (N_14522,N_14204,N_14355);
nor U14523 (N_14523,N_14294,N_14302);
or U14524 (N_14524,N_14394,N_14380);
nand U14525 (N_14525,N_14385,N_14328);
nand U14526 (N_14526,N_14320,N_14285);
or U14527 (N_14527,N_14205,N_14217);
or U14528 (N_14528,N_14384,N_14327);
nand U14529 (N_14529,N_14233,N_14201);
nor U14530 (N_14530,N_14304,N_14286);
or U14531 (N_14531,N_14308,N_14241);
nor U14532 (N_14532,N_14382,N_14313);
xnor U14533 (N_14533,N_14279,N_14263);
nor U14534 (N_14534,N_14297,N_14225);
xnor U14535 (N_14535,N_14256,N_14304);
xor U14536 (N_14536,N_14208,N_14337);
xnor U14537 (N_14537,N_14354,N_14245);
nand U14538 (N_14538,N_14315,N_14239);
nand U14539 (N_14539,N_14363,N_14378);
or U14540 (N_14540,N_14256,N_14353);
and U14541 (N_14541,N_14362,N_14232);
nand U14542 (N_14542,N_14347,N_14260);
or U14543 (N_14543,N_14225,N_14356);
or U14544 (N_14544,N_14244,N_14348);
nor U14545 (N_14545,N_14206,N_14286);
and U14546 (N_14546,N_14280,N_14305);
xor U14547 (N_14547,N_14217,N_14379);
xor U14548 (N_14548,N_14209,N_14306);
and U14549 (N_14549,N_14310,N_14309);
or U14550 (N_14550,N_14381,N_14253);
and U14551 (N_14551,N_14388,N_14353);
nor U14552 (N_14552,N_14240,N_14325);
xor U14553 (N_14553,N_14316,N_14245);
nor U14554 (N_14554,N_14331,N_14399);
xnor U14555 (N_14555,N_14273,N_14310);
or U14556 (N_14556,N_14307,N_14356);
xor U14557 (N_14557,N_14274,N_14293);
nor U14558 (N_14558,N_14387,N_14223);
nand U14559 (N_14559,N_14214,N_14286);
and U14560 (N_14560,N_14298,N_14288);
xnor U14561 (N_14561,N_14258,N_14396);
and U14562 (N_14562,N_14243,N_14245);
nand U14563 (N_14563,N_14226,N_14333);
or U14564 (N_14564,N_14293,N_14240);
nor U14565 (N_14565,N_14217,N_14339);
nand U14566 (N_14566,N_14304,N_14357);
or U14567 (N_14567,N_14247,N_14281);
nand U14568 (N_14568,N_14256,N_14230);
or U14569 (N_14569,N_14231,N_14213);
xnor U14570 (N_14570,N_14379,N_14359);
or U14571 (N_14571,N_14227,N_14223);
xor U14572 (N_14572,N_14288,N_14286);
or U14573 (N_14573,N_14227,N_14233);
xnor U14574 (N_14574,N_14299,N_14324);
or U14575 (N_14575,N_14222,N_14390);
nand U14576 (N_14576,N_14373,N_14368);
nand U14577 (N_14577,N_14214,N_14219);
xor U14578 (N_14578,N_14338,N_14222);
xor U14579 (N_14579,N_14275,N_14337);
or U14580 (N_14580,N_14216,N_14352);
xor U14581 (N_14581,N_14293,N_14364);
nand U14582 (N_14582,N_14262,N_14329);
and U14583 (N_14583,N_14297,N_14254);
nor U14584 (N_14584,N_14302,N_14356);
nor U14585 (N_14585,N_14344,N_14268);
or U14586 (N_14586,N_14345,N_14380);
xnor U14587 (N_14587,N_14293,N_14324);
nor U14588 (N_14588,N_14282,N_14220);
nand U14589 (N_14589,N_14368,N_14398);
and U14590 (N_14590,N_14355,N_14364);
xnor U14591 (N_14591,N_14354,N_14262);
or U14592 (N_14592,N_14219,N_14323);
nand U14593 (N_14593,N_14252,N_14315);
nor U14594 (N_14594,N_14263,N_14326);
or U14595 (N_14595,N_14319,N_14284);
or U14596 (N_14596,N_14223,N_14305);
or U14597 (N_14597,N_14258,N_14354);
nand U14598 (N_14598,N_14382,N_14355);
nor U14599 (N_14599,N_14249,N_14385);
and U14600 (N_14600,N_14459,N_14472);
or U14601 (N_14601,N_14435,N_14524);
nand U14602 (N_14602,N_14579,N_14411);
and U14603 (N_14603,N_14549,N_14504);
or U14604 (N_14604,N_14457,N_14410);
or U14605 (N_14605,N_14422,N_14434);
nor U14606 (N_14606,N_14546,N_14482);
or U14607 (N_14607,N_14574,N_14441);
nand U14608 (N_14608,N_14424,N_14429);
nor U14609 (N_14609,N_14570,N_14406);
and U14610 (N_14610,N_14499,N_14597);
nand U14611 (N_14611,N_14454,N_14523);
or U14612 (N_14612,N_14505,N_14465);
and U14613 (N_14613,N_14554,N_14517);
or U14614 (N_14614,N_14527,N_14427);
nor U14615 (N_14615,N_14593,N_14537);
nand U14616 (N_14616,N_14532,N_14521);
xor U14617 (N_14617,N_14552,N_14589);
nor U14618 (N_14618,N_14415,N_14467);
xnor U14619 (N_14619,N_14433,N_14571);
and U14620 (N_14620,N_14413,N_14449);
nand U14621 (N_14621,N_14494,N_14536);
or U14622 (N_14622,N_14451,N_14453);
nor U14623 (N_14623,N_14520,N_14588);
and U14624 (N_14624,N_14471,N_14509);
or U14625 (N_14625,N_14529,N_14428);
or U14626 (N_14626,N_14475,N_14445);
xor U14627 (N_14627,N_14559,N_14567);
xnor U14628 (N_14628,N_14468,N_14414);
nand U14629 (N_14629,N_14511,N_14486);
nor U14630 (N_14630,N_14452,N_14572);
nor U14631 (N_14631,N_14558,N_14405);
xor U14632 (N_14632,N_14569,N_14587);
nor U14633 (N_14633,N_14501,N_14513);
nand U14634 (N_14634,N_14561,N_14566);
nand U14635 (N_14635,N_14481,N_14512);
nor U14636 (N_14636,N_14470,N_14510);
nor U14637 (N_14637,N_14476,N_14599);
and U14638 (N_14638,N_14477,N_14514);
nand U14639 (N_14639,N_14403,N_14490);
and U14640 (N_14640,N_14551,N_14506);
or U14641 (N_14641,N_14489,N_14446);
or U14642 (N_14642,N_14444,N_14448);
nand U14643 (N_14643,N_14580,N_14430);
nand U14644 (N_14644,N_14522,N_14450);
nand U14645 (N_14645,N_14479,N_14423);
and U14646 (N_14646,N_14436,N_14402);
and U14647 (N_14647,N_14496,N_14582);
nor U14648 (N_14648,N_14495,N_14417);
or U14649 (N_14649,N_14548,N_14426);
xor U14650 (N_14650,N_14575,N_14466);
or U14651 (N_14651,N_14455,N_14592);
or U14652 (N_14652,N_14584,N_14456);
xor U14653 (N_14653,N_14576,N_14563);
nor U14654 (N_14654,N_14556,N_14526);
or U14655 (N_14655,N_14591,N_14595);
xor U14656 (N_14656,N_14550,N_14507);
nand U14657 (N_14657,N_14491,N_14531);
or U14658 (N_14658,N_14508,N_14578);
xor U14659 (N_14659,N_14420,N_14525);
or U14660 (N_14660,N_14502,N_14503);
or U14661 (N_14661,N_14432,N_14542);
xor U14662 (N_14662,N_14461,N_14442);
xor U14663 (N_14663,N_14439,N_14401);
nand U14664 (N_14664,N_14586,N_14443);
xnor U14665 (N_14665,N_14598,N_14573);
nand U14666 (N_14666,N_14437,N_14545);
and U14667 (N_14667,N_14590,N_14585);
xor U14668 (N_14668,N_14487,N_14462);
and U14669 (N_14669,N_14485,N_14412);
and U14670 (N_14670,N_14583,N_14409);
nand U14671 (N_14671,N_14530,N_14493);
xor U14672 (N_14672,N_14419,N_14538);
xor U14673 (N_14673,N_14483,N_14594);
nand U14674 (N_14674,N_14543,N_14539);
and U14675 (N_14675,N_14440,N_14474);
and U14676 (N_14676,N_14421,N_14418);
nand U14677 (N_14677,N_14535,N_14540);
xor U14678 (N_14678,N_14407,N_14464);
and U14679 (N_14679,N_14519,N_14425);
xor U14680 (N_14680,N_14564,N_14562);
and U14681 (N_14681,N_14544,N_14469);
and U14682 (N_14682,N_14577,N_14438);
nor U14683 (N_14683,N_14463,N_14460);
or U14684 (N_14684,N_14447,N_14416);
nand U14685 (N_14685,N_14404,N_14488);
xor U14686 (N_14686,N_14528,N_14500);
xor U14687 (N_14687,N_14518,N_14547);
and U14688 (N_14688,N_14560,N_14568);
or U14689 (N_14689,N_14492,N_14533);
and U14690 (N_14690,N_14458,N_14581);
xnor U14691 (N_14691,N_14516,N_14408);
nor U14692 (N_14692,N_14555,N_14565);
nor U14693 (N_14693,N_14484,N_14541);
nor U14694 (N_14694,N_14498,N_14480);
or U14695 (N_14695,N_14400,N_14515);
xor U14696 (N_14696,N_14473,N_14497);
nand U14697 (N_14697,N_14596,N_14478);
and U14698 (N_14698,N_14553,N_14534);
or U14699 (N_14699,N_14557,N_14431);
nand U14700 (N_14700,N_14511,N_14530);
nand U14701 (N_14701,N_14596,N_14590);
and U14702 (N_14702,N_14599,N_14439);
nor U14703 (N_14703,N_14522,N_14566);
and U14704 (N_14704,N_14464,N_14438);
nor U14705 (N_14705,N_14454,N_14480);
and U14706 (N_14706,N_14482,N_14538);
nand U14707 (N_14707,N_14450,N_14416);
or U14708 (N_14708,N_14430,N_14512);
nand U14709 (N_14709,N_14486,N_14431);
nand U14710 (N_14710,N_14407,N_14546);
and U14711 (N_14711,N_14437,N_14539);
or U14712 (N_14712,N_14440,N_14511);
and U14713 (N_14713,N_14490,N_14506);
and U14714 (N_14714,N_14589,N_14402);
or U14715 (N_14715,N_14491,N_14557);
and U14716 (N_14716,N_14438,N_14459);
xnor U14717 (N_14717,N_14425,N_14468);
and U14718 (N_14718,N_14456,N_14482);
nand U14719 (N_14719,N_14428,N_14477);
nor U14720 (N_14720,N_14449,N_14502);
nand U14721 (N_14721,N_14484,N_14589);
nand U14722 (N_14722,N_14461,N_14553);
xnor U14723 (N_14723,N_14530,N_14469);
nor U14724 (N_14724,N_14524,N_14441);
nand U14725 (N_14725,N_14537,N_14559);
nor U14726 (N_14726,N_14431,N_14483);
nand U14727 (N_14727,N_14467,N_14488);
and U14728 (N_14728,N_14542,N_14544);
nor U14729 (N_14729,N_14482,N_14404);
or U14730 (N_14730,N_14596,N_14580);
nand U14731 (N_14731,N_14520,N_14571);
or U14732 (N_14732,N_14415,N_14441);
or U14733 (N_14733,N_14590,N_14540);
nand U14734 (N_14734,N_14530,N_14591);
or U14735 (N_14735,N_14499,N_14489);
or U14736 (N_14736,N_14410,N_14592);
and U14737 (N_14737,N_14543,N_14447);
nand U14738 (N_14738,N_14492,N_14536);
and U14739 (N_14739,N_14440,N_14540);
and U14740 (N_14740,N_14455,N_14440);
or U14741 (N_14741,N_14549,N_14487);
nand U14742 (N_14742,N_14404,N_14531);
nor U14743 (N_14743,N_14472,N_14528);
or U14744 (N_14744,N_14422,N_14497);
xor U14745 (N_14745,N_14556,N_14452);
nand U14746 (N_14746,N_14561,N_14480);
nand U14747 (N_14747,N_14537,N_14454);
nor U14748 (N_14748,N_14553,N_14446);
nand U14749 (N_14749,N_14436,N_14595);
nand U14750 (N_14750,N_14464,N_14525);
nand U14751 (N_14751,N_14521,N_14528);
xor U14752 (N_14752,N_14459,N_14408);
nor U14753 (N_14753,N_14532,N_14539);
nor U14754 (N_14754,N_14431,N_14504);
nor U14755 (N_14755,N_14518,N_14404);
nand U14756 (N_14756,N_14423,N_14459);
xor U14757 (N_14757,N_14550,N_14429);
and U14758 (N_14758,N_14519,N_14444);
or U14759 (N_14759,N_14467,N_14598);
nand U14760 (N_14760,N_14565,N_14465);
or U14761 (N_14761,N_14582,N_14549);
nor U14762 (N_14762,N_14437,N_14442);
nand U14763 (N_14763,N_14499,N_14456);
or U14764 (N_14764,N_14597,N_14535);
nand U14765 (N_14765,N_14488,N_14537);
and U14766 (N_14766,N_14510,N_14587);
and U14767 (N_14767,N_14480,N_14523);
xnor U14768 (N_14768,N_14447,N_14429);
nor U14769 (N_14769,N_14553,N_14503);
nand U14770 (N_14770,N_14406,N_14403);
nor U14771 (N_14771,N_14412,N_14408);
or U14772 (N_14772,N_14551,N_14586);
or U14773 (N_14773,N_14435,N_14473);
or U14774 (N_14774,N_14430,N_14409);
nor U14775 (N_14775,N_14490,N_14411);
xnor U14776 (N_14776,N_14425,N_14511);
nand U14777 (N_14777,N_14528,N_14587);
xnor U14778 (N_14778,N_14401,N_14597);
xor U14779 (N_14779,N_14492,N_14409);
nor U14780 (N_14780,N_14443,N_14437);
nor U14781 (N_14781,N_14449,N_14591);
nand U14782 (N_14782,N_14524,N_14541);
nand U14783 (N_14783,N_14409,N_14481);
and U14784 (N_14784,N_14459,N_14410);
or U14785 (N_14785,N_14518,N_14442);
or U14786 (N_14786,N_14579,N_14461);
or U14787 (N_14787,N_14545,N_14468);
nor U14788 (N_14788,N_14481,N_14499);
and U14789 (N_14789,N_14585,N_14461);
xor U14790 (N_14790,N_14540,N_14437);
nor U14791 (N_14791,N_14413,N_14403);
or U14792 (N_14792,N_14579,N_14473);
xor U14793 (N_14793,N_14586,N_14424);
or U14794 (N_14794,N_14582,N_14528);
xnor U14795 (N_14795,N_14532,N_14522);
and U14796 (N_14796,N_14450,N_14492);
and U14797 (N_14797,N_14539,N_14501);
and U14798 (N_14798,N_14571,N_14418);
nor U14799 (N_14799,N_14442,N_14547);
nor U14800 (N_14800,N_14772,N_14650);
and U14801 (N_14801,N_14744,N_14605);
nor U14802 (N_14802,N_14642,N_14667);
xnor U14803 (N_14803,N_14665,N_14763);
xnor U14804 (N_14804,N_14627,N_14733);
xor U14805 (N_14805,N_14643,N_14698);
and U14806 (N_14806,N_14678,N_14654);
xor U14807 (N_14807,N_14797,N_14616);
nand U14808 (N_14808,N_14610,N_14641);
nand U14809 (N_14809,N_14769,N_14789);
xor U14810 (N_14810,N_14609,N_14708);
xnor U14811 (N_14811,N_14685,N_14786);
nand U14812 (N_14812,N_14730,N_14765);
or U14813 (N_14813,N_14745,N_14779);
nand U14814 (N_14814,N_14635,N_14751);
or U14815 (N_14815,N_14639,N_14660);
and U14816 (N_14816,N_14787,N_14696);
nand U14817 (N_14817,N_14777,N_14647);
xnor U14818 (N_14818,N_14653,N_14792);
and U14819 (N_14819,N_14659,N_14675);
nand U14820 (N_14820,N_14798,N_14759);
nor U14821 (N_14821,N_14767,N_14640);
nor U14822 (N_14822,N_14741,N_14790);
xnor U14823 (N_14823,N_14711,N_14607);
xor U14824 (N_14824,N_14718,N_14634);
nor U14825 (N_14825,N_14602,N_14783);
or U14826 (N_14826,N_14756,N_14734);
xor U14827 (N_14827,N_14713,N_14776);
and U14828 (N_14828,N_14753,N_14699);
and U14829 (N_14829,N_14621,N_14773);
nand U14830 (N_14830,N_14742,N_14766);
nand U14831 (N_14831,N_14752,N_14714);
xnor U14832 (N_14832,N_14774,N_14788);
or U14833 (N_14833,N_14796,N_14760);
or U14834 (N_14834,N_14666,N_14604);
nand U14835 (N_14835,N_14630,N_14780);
nor U14836 (N_14836,N_14732,N_14695);
nand U14837 (N_14837,N_14704,N_14631);
or U14838 (N_14838,N_14663,N_14683);
xnor U14839 (N_14839,N_14706,N_14617);
nor U14840 (N_14840,N_14717,N_14775);
and U14841 (N_14841,N_14727,N_14613);
nand U14842 (N_14842,N_14646,N_14747);
and U14843 (N_14843,N_14748,N_14655);
nand U14844 (N_14844,N_14652,N_14636);
and U14845 (N_14845,N_14686,N_14782);
and U14846 (N_14846,N_14672,N_14677);
xor U14847 (N_14847,N_14720,N_14632);
and U14848 (N_14848,N_14676,N_14633);
or U14849 (N_14849,N_14735,N_14731);
nand U14850 (N_14850,N_14618,N_14791);
xnor U14851 (N_14851,N_14669,N_14619);
or U14852 (N_14852,N_14721,N_14690);
or U14853 (N_14853,N_14680,N_14674);
nand U14854 (N_14854,N_14729,N_14645);
and U14855 (N_14855,N_14625,N_14637);
and U14856 (N_14856,N_14601,N_14784);
nor U14857 (N_14857,N_14719,N_14755);
nor U14858 (N_14858,N_14606,N_14628);
or U14859 (N_14859,N_14638,N_14707);
and U14860 (N_14860,N_14673,N_14768);
nor U14861 (N_14861,N_14770,N_14691);
or U14862 (N_14862,N_14629,N_14795);
nand U14863 (N_14863,N_14716,N_14725);
nand U14864 (N_14864,N_14703,N_14692);
and U14865 (N_14865,N_14608,N_14681);
xnor U14866 (N_14866,N_14778,N_14657);
nand U14867 (N_14867,N_14710,N_14709);
or U14868 (N_14868,N_14722,N_14738);
nand U14869 (N_14869,N_14702,N_14656);
nor U14870 (N_14870,N_14705,N_14712);
nand U14871 (N_14871,N_14689,N_14758);
nor U14872 (N_14872,N_14694,N_14794);
nor U14873 (N_14873,N_14737,N_14603);
nand U14874 (N_14874,N_14764,N_14740);
xnor U14875 (N_14875,N_14700,N_14600);
or U14876 (N_14876,N_14693,N_14623);
or U14877 (N_14877,N_14743,N_14668);
and U14878 (N_14878,N_14622,N_14754);
nor U14879 (N_14879,N_14761,N_14762);
nor U14880 (N_14880,N_14658,N_14726);
nor U14881 (N_14881,N_14771,N_14626);
nand U14882 (N_14882,N_14662,N_14781);
nand U14883 (N_14883,N_14749,N_14620);
xor U14884 (N_14884,N_14785,N_14661);
or U14885 (N_14885,N_14644,N_14757);
xnor U14886 (N_14886,N_14664,N_14614);
and U14887 (N_14887,N_14651,N_14611);
nor U14888 (N_14888,N_14746,N_14688);
or U14889 (N_14889,N_14697,N_14687);
xor U14890 (N_14890,N_14684,N_14648);
xor U14891 (N_14891,N_14723,N_14671);
xor U14892 (N_14892,N_14736,N_14724);
nand U14893 (N_14893,N_14799,N_14728);
xor U14894 (N_14894,N_14649,N_14701);
xor U14895 (N_14895,N_14715,N_14670);
xor U14896 (N_14896,N_14682,N_14739);
nor U14897 (N_14897,N_14624,N_14793);
nor U14898 (N_14898,N_14679,N_14750);
xnor U14899 (N_14899,N_14615,N_14612);
nand U14900 (N_14900,N_14742,N_14794);
and U14901 (N_14901,N_14717,N_14606);
nor U14902 (N_14902,N_14605,N_14752);
xor U14903 (N_14903,N_14782,N_14752);
or U14904 (N_14904,N_14688,N_14694);
nand U14905 (N_14905,N_14609,N_14784);
nand U14906 (N_14906,N_14607,N_14660);
nor U14907 (N_14907,N_14738,N_14780);
or U14908 (N_14908,N_14660,N_14781);
nor U14909 (N_14909,N_14744,N_14742);
or U14910 (N_14910,N_14697,N_14780);
nor U14911 (N_14911,N_14685,N_14730);
and U14912 (N_14912,N_14658,N_14746);
and U14913 (N_14913,N_14662,N_14665);
xor U14914 (N_14914,N_14702,N_14749);
xnor U14915 (N_14915,N_14630,N_14754);
or U14916 (N_14916,N_14661,N_14635);
nand U14917 (N_14917,N_14690,N_14652);
nor U14918 (N_14918,N_14622,N_14628);
xor U14919 (N_14919,N_14706,N_14751);
nand U14920 (N_14920,N_14769,N_14721);
or U14921 (N_14921,N_14694,N_14701);
and U14922 (N_14922,N_14608,N_14623);
or U14923 (N_14923,N_14645,N_14702);
nand U14924 (N_14924,N_14602,N_14732);
and U14925 (N_14925,N_14731,N_14747);
and U14926 (N_14926,N_14616,N_14618);
and U14927 (N_14927,N_14626,N_14702);
and U14928 (N_14928,N_14675,N_14786);
or U14929 (N_14929,N_14733,N_14657);
nor U14930 (N_14930,N_14694,N_14730);
or U14931 (N_14931,N_14750,N_14716);
or U14932 (N_14932,N_14766,N_14664);
and U14933 (N_14933,N_14695,N_14661);
and U14934 (N_14934,N_14786,N_14604);
and U14935 (N_14935,N_14740,N_14700);
nor U14936 (N_14936,N_14783,N_14784);
or U14937 (N_14937,N_14704,N_14698);
nand U14938 (N_14938,N_14674,N_14605);
or U14939 (N_14939,N_14656,N_14659);
nor U14940 (N_14940,N_14627,N_14651);
xnor U14941 (N_14941,N_14737,N_14675);
nor U14942 (N_14942,N_14676,N_14636);
xor U14943 (N_14943,N_14706,N_14658);
and U14944 (N_14944,N_14675,N_14706);
nor U14945 (N_14945,N_14671,N_14711);
or U14946 (N_14946,N_14748,N_14678);
xor U14947 (N_14947,N_14704,N_14721);
nand U14948 (N_14948,N_14681,N_14755);
nor U14949 (N_14949,N_14740,N_14775);
xor U14950 (N_14950,N_14607,N_14606);
and U14951 (N_14951,N_14729,N_14777);
nor U14952 (N_14952,N_14767,N_14650);
nand U14953 (N_14953,N_14778,N_14673);
nand U14954 (N_14954,N_14722,N_14615);
nand U14955 (N_14955,N_14664,N_14794);
or U14956 (N_14956,N_14794,N_14780);
and U14957 (N_14957,N_14654,N_14772);
or U14958 (N_14958,N_14672,N_14743);
and U14959 (N_14959,N_14760,N_14792);
and U14960 (N_14960,N_14779,N_14608);
nor U14961 (N_14961,N_14623,N_14643);
and U14962 (N_14962,N_14791,N_14664);
nor U14963 (N_14963,N_14770,N_14690);
xor U14964 (N_14964,N_14734,N_14675);
or U14965 (N_14965,N_14643,N_14744);
or U14966 (N_14966,N_14689,N_14686);
or U14967 (N_14967,N_14759,N_14693);
nor U14968 (N_14968,N_14786,N_14616);
or U14969 (N_14969,N_14786,N_14600);
nand U14970 (N_14970,N_14715,N_14606);
nand U14971 (N_14971,N_14605,N_14749);
nor U14972 (N_14972,N_14627,N_14684);
and U14973 (N_14973,N_14771,N_14677);
nand U14974 (N_14974,N_14634,N_14661);
and U14975 (N_14975,N_14704,N_14628);
and U14976 (N_14976,N_14621,N_14731);
xnor U14977 (N_14977,N_14619,N_14709);
or U14978 (N_14978,N_14667,N_14649);
nand U14979 (N_14979,N_14622,N_14683);
nor U14980 (N_14980,N_14719,N_14647);
and U14981 (N_14981,N_14650,N_14719);
nor U14982 (N_14982,N_14690,N_14635);
xor U14983 (N_14983,N_14607,N_14760);
nand U14984 (N_14984,N_14625,N_14705);
xnor U14985 (N_14985,N_14657,N_14633);
and U14986 (N_14986,N_14649,N_14645);
nand U14987 (N_14987,N_14615,N_14743);
or U14988 (N_14988,N_14681,N_14739);
and U14989 (N_14989,N_14792,N_14659);
nand U14990 (N_14990,N_14619,N_14717);
nor U14991 (N_14991,N_14697,N_14700);
or U14992 (N_14992,N_14719,N_14686);
xor U14993 (N_14993,N_14798,N_14730);
and U14994 (N_14994,N_14616,N_14619);
nand U14995 (N_14995,N_14618,N_14700);
xor U14996 (N_14996,N_14752,N_14727);
or U14997 (N_14997,N_14739,N_14795);
and U14998 (N_14998,N_14686,N_14691);
nand U14999 (N_14999,N_14788,N_14707);
xnor U15000 (N_15000,N_14864,N_14871);
or U15001 (N_15001,N_14845,N_14972);
or U15002 (N_15002,N_14925,N_14839);
xnor U15003 (N_15003,N_14975,N_14825);
nand U15004 (N_15004,N_14982,N_14811);
nor U15005 (N_15005,N_14977,N_14922);
nand U15006 (N_15006,N_14892,N_14911);
xnor U15007 (N_15007,N_14955,N_14857);
and U15008 (N_15008,N_14807,N_14872);
and U15009 (N_15009,N_14859,N_14906);
nand U15010 (N_15010,N_14909,N_14919);
xnor U15011 (N_15011,N_14868,N_14969);
and U15012 (N_15012,N_14855,N_14877);
xnor U15013 (N_15013,N_14945,N_14820);
or U15014 (N_15014,N_14953,N_14921);
nand U15015 (N_15015,N_14970,N_14880);
and U15016 (N_15016,N_14998,N_14973);
xnor U15017 (N_15017,N_14850,N_14858);
nand U15018 (N_15018,N_14822,N_14810);
and U15019 (N_15019,N_14938,N_14804);
nor U15020 (N_15020,N_14971,N_14918);
nand U15021 (N_15021,N_14933,N_14950);
and U15022 (N_15022,N_14937,N_14849);
nand U15023 (N_15023,N_14819,N_14979);
nor U15024 (N_15024,N_14854,N_14996);
or U15025 (N_15025,N_14896,N_14876);
nor U15026 (N_15026,N_14885,N_14856);
nor U15027 (N_15027,N_14917,N_14823);
or U15028 (N_15028,N_14986,N_14948);
nor U15029 (N_15029,N_14983,N_14842);
xnor U15030 (N_15030,N_14992,N_14828);
and U15031 (N_15031,N_14994,N_14812);
or U15032 (N_15032,N_14987,N_14847);
or U15033 (N_15033,N_14974,N_14827);
and U15034 (N_15034,N_14824,N_14960);
and U15035 (N_15035,N_14836,N_14862);
or U15036 (N_15036,N_14863,N_14866);
and U15037 (N_15037,N_14988,N_14878);
nand U15038 (N_15038,N_14894,N_14879);
nand U15039 (N_15039,N_14914,N_14813);
and U15040 (N_15040,N_14958,N_14883);
or U15041 (N_15041,N_14818,N_14908);
xor U15042 (N_15042,N_14840,N_14816);
nor U15043 (N_15043,N_14852,N_14904);
and U15044 (N_15044,N_14841,N_14947);
or U15045 (N_15045,N_14999,N_14803);
and U15046 (N_15046,N_14890,N_14993);
and U15047 (N_15047,N_14949,N_14805);
nand U15048 (N_15048,N_14932,N_14963);
nor U15049 (N_15049,N_14800,N_14965);
xnor U15050 (N_15050,N_14814,N_14899);
nor U15051 (N_15051,N_14838,N_14957);
or U15052 (N_15052,N_14935,N_14926);
or U15053 (N_15053,N_14873,N_14954);
nand U15054 (N_15054,N_14830,N_14942);
xor U15055 (N_15055,N_14889,N_14920);
xor U15056 (N_15056,N_14821,N_14980);
xor U15057 (N_15057,N_14956,N_14978);
xor U15058 (N_15058,N_14888,N_14981);
nor U15059 (N_15059,N_14934,N_14865);
or U15060 (N_15060,N_14834,N_14989);
and U15061 (N_15061,N_14815,N_14843);
and U15062 (N_15062,N_14829,N_14928);
nor U15063 (N_15063,N_14936,N_14910);
nand U15064 (N_15064,N_14844,N_14806);
xnor U15065 (N_15065,N_14923,N_14968);
and U15066 (N_15066,N_14808,N_14991);
or U15067 (N_15067,N_14916,N_14881);
or U15068 (N_15068,N_14902,N_14875);
nor U15069 (N_15069,N_14801,N_14995);
nand U15070 (N_15070,N_14985,N_14901);
nand U15071 (N_15071,N_14826,N_14915);
nor U15072 (N_15072,N_14861,N_14853);
nor U15073 (N_15073,N_14860,N_14900);
or U15074 (N_15074,N_14831,N_14967);
nand U15075 (N_15075,N_14893,N_14837);
xnor U15076 (N_15076,N_14886,N_14930);
or U15077 (N_15077,N_14943,N_14951);
or U15078 (N_15078,N_14833,N_14898);
xor U15079 (N_15079,N_14882,N_14964);
xnor U15080 (N_15080,N_14846,N_14962);
and U15081 (N_15081,N_14912,N_14997);
and U15082 (N_15082,N_14941,N_14905);
or U15083 (N_15083,N_14874,N_14887);
nand U15084 (N_15084,N_14939,N_14895);
nor U15085 (N_15085,N_14851,N_14891);
or U15086 (N_15086,N_14867,N_14884);
nand U15087 (N_15087,N_14870,N_14931);
and U15088 (N_15088,N_14848,N_14952);
nor U15089 (N_15089,N_14940,N_14966);
or U15090 (N_15090,N_14897,N_14976);
xnor U15091 (N_15091,N_14809,N_14927);
or U15092 (N_15092,N_14959,N_14832);
nor U15093 (N_15093,N_14913,N_14907);
or U15094 (N_15094,N_14817,N_14903);
xnor U15095 (N_15095,N_14929,N_14869);
and U15096 (N_15096,N_14984,N_14944);
and U15097 (N_15097,N_14802,N_14835);
nand U15098 (N_15098,N_14961,N_14924);
nor U15099 (N_15099,N_14946,N_14990);
or U15100 (N_15100,N_14935,N_14909);
and U15101 (N_15101,N_14848,N_14925);
and U15102 (N_15102,N_14996,N_14855);
nor U15103 (N_15103,N_14822,N_14817);
xor U15104 (N_15104,N_14847,N_14985);
and U15105 (N_15105,N_14930,N_14957);
xor U15106 (N_15106,N_14890,N_14963);
nor U15107 (N_15107,N_14811,N_14972);
nand U15108 (N_15108,N_14952,N_14802);
and U15109 (N_15109,N_14940,N_14856);
xnor U15110 (N_15110,N_14958,N_14999);
nor U15111 (N_15111,N_14824,N_14942);
nand U15112 (N_15112,N_14926,N_14991);
and U15113 (N_15113,N_14819,N_14926);
xnor U15114 (N_15114,N_14912,N_14965);
nand U15115 (N_15115,N_14932,N_14873);
or U15116 (N_15116,N_14926,N_14917);
nor U15117 (N_15117,N_14843,N_14948);
nand U15118 (N_15118,N_14839,N_14945);
or U15119 (N_15119,N_14928,N_14805);
nor U15120 (N_15120,N_14818,N_14902);
nand U15121 (N_15121,N_14850,N_14968);
and U15122 (N_15122,N_14891,N_14963);
or U15123 (N_15123,N_14891,N_14915);
nor U15124 (N_15124,N_14940,N_14887);
or U15125 (N_15125,N_14979,N_14971);
nand U15126 (N_15126,N_14803,N_14980);
or U15127 (N_15127,N_14984,N_14900);
xnor U15128 (N_15128,N_14941,N_14930);
nor U15129 (N_15129,N_14935,N_14898);
and U15130 (N_15130,N_14845,N_14809);
nand U15131 (N_15131,N_14995,N_14980);
or U15132 (N_15132,N_14934,N_14910);
and U15133 (N_15133,N_14959,N_14864);
nor U15134 (N_15134,N_14938,N_14930);
xnor U15135 (N_15135,N_14972,N_14863);
nor U15136 (N_15136,N_14904,N_14958);
or U15137 (N_15137,N_14873,N_14957);
and U15138 (N_15138,N_14821,N_14967);
or U15139 (N_15139,N_14887,N_14886);
nand U15140 (N_15140,N_14901,N_14914);
xor U15141 (N_15141,N_14947,N_14875);
or U15142 (N_15142,N_14881,N_14952);
xor U15143 (N_15143,N_14936,N_14853);
nand U15144 (N_15144,N_14898,N_14970);
and U15145 (N_15145,N_14928,N_14879);
xnor U15146 (N_15146,N_14986,N_14820);
or U15147 (N_15147,N_14935,N_14983);
or U15148 (N_15148,N_14925,N_14987);
nand U15149 (N_15149,N_14876,N_14843);
or U15150 (N_15150,N_14993,N_14869);
and U15151 (N_15151,N_14957,N_14918);
xor U15152 (N_15152,N_14877,N_14852);
and U15153 (N_15153,N_14861,N_14815);
nand U15154 (N_15154,N_14814,N_14975);
xor U15155 (N_15155,N_14903,N_14960);
and U15156 (N_15156,N_14981,N_14946);
or U15157 (N_15157,N_14841,N_14949);
nand U15158 (N_15158,N_14998,N_14864);
nor U15159 (N_15159,N_14945,N_14904);
or U15160 (N_15160,N_14820,N_14993);
nand U15161 (N_15161,N_14903,N_14943);
nand U15162 (N_15162,N_14808,N_14930);
nor U15163 (N_15163,N_14945,N_14862);
nand U15164 (N_15164,N_14970,N_14992);
nor U15165 (N_15165,N_14906,N_14923);
and U15166 (N_15166,N_14858,N_14901);
nand U15167 (N_15167,N_14822,N_14919);
nand U15168 (N_15168,N_14855,N_14906);
or U15169 (N_15169,N_14978,N_14829);
and U15170 (N_15170,N_14872,N_14912);
or U15171 (N_15171,N_14843,N_14914);
or U15172 (N_15172,N_14855,N_14927);
or U15173 (N_15173,N_14975,N_14851);
or U15174 (N_15174,N_14921,N_14856);
or U15175 (N_15175,N_14929,N_14959);
or U15176 (N_15176,N_14895,N_14843);
nand U15177 (N_15177,N_14803,N_14915);
xnor U15178 (N_15178,N_14919,N_14991);
and U15179 (N_15179,N_14810,N_14803);
nand U15180 (N_15180,N_14925,N_14822);
nor U15181 (N_15181,N_14848,N_14961);
nand U15182 (N_15182,N_14824,N_14841);
nor U15183 (N_15183,N_14839,N_14869);
nor U15184 (N_15184,N_14954,N_14984);
and U15185 (N_15185,N_14972,N_14830);
or U15186 (N_15186,N_14912,N_14957);
nand U15187 (N_15187,N_14862,N_14979);
xor U15188 (N_15188,N_14987,N_14941);
or U15189 (N_15189,N_14821,N_14820);
nand U15190 (N_15190,N_14957,N_14910);
and U15191 (N_15191,N_14995,N_14978);
nor U15192 (N_15192,N_14878,N_14802);
or U15193 (N_15193,N_14925,N_14974);
nand U15194 (N_15194,N_14954,N_14971);
nor U15195 (N_15195,N_14871,N_14993);
nor U15196 (N_15196,N_14819,N_14822);
nor U15197 (N_15197,N_14968,N_14800);
or U15198 (N_15198,N_14830,N_14916);
nand U15199 (N_15199,N_14817,N_14984);
and U15200 (N_15200,N_15063,N_15164);
or U15201 (N_15201,N_15088,N_15123);
xor U15202 (N_15202,N_15058,N_15178);
and U15203 (N_15203,N_15101,N_15004);
xnor U15204 (N_15204,N_15054,N_15079);
and U15205 (N_15205,N_15048,N_15107);
xor U15206 (N_15206,N_15174,N_15171);
and U15207 (N_15207,N_15185,N_15018);
nor U15208 (N_15208,N_15147,N_15096);
xor U15209 (N_15209,N_15023,N_15150);
nand U15210 (N_15210,N_15127,N_15108);
nand U15211 (N_15211,N_15102,N_15074);
or U15212 (N_15212,N_15175,N_15124);
nor U15213 (N_15213,N_15151,N_15037);
nor U15214 (N_15214,N_15136,N_15009);
xor U15215 (N_15215,N_15053,N_15126);
nand U15216 (N_15216,N_15194,N_15033);
nor U15217 (N_15217,N_15121,N_15120);
xor U15218 (N_15218,N_15133,N_15131);
and U15219 (N_15219,N_15105,N_15049);
and U15220 (N_15220,N_15183,N_15104);
or U15221 (N_15221,N_15060,N_15006);
nand U15222 (N_15222,N_15122,N_15115);
nand U15223 (N_15223,N_15027,N_15180);
nand U15224 (N_15224,N_15062,N_15137);
and U15225 (N_15225,N_15197,N_15003);
nand U15226 (N_15226,N_15119,N_15128);
nand U15227 (N_15227,N_15116,N_15158);
or U15228 (N_15228,N_15140,N_15153);
nand U15229 (N_15229,N_15012,N_15092);
and U15230 (N_15230,N_15052,N_15129);
xnor U15231 (N_15231,N_15076,N_15106);
and U15232 (N_15232,N_15082,N_15013);
and U15233 (N_15233,N_15125,N_15103);
xnor U15234 (N_15234,N_15169,N_15196);
nor U15235 (N_15235,N_15142,N_15064);
xnor U15236 (N_15236,N_15149,N_15166);
xor U15237 (N_15237,N_15177,N_15040);
xnor U15238 (N_15238,N_15181,N_15067);
or U15239 (N_15239,N_15110,N_15090);
xor U15240 (N_15240,N_15000,N_15097);
or U15241 (N_15241,N_15039,N_15160);
nand U15242 (N_15242,N_15043,N_15186);
or U15243 (N_15243,N_15077,N_15051);
or U15244 (N_15244,N_15024,N_15044);
and U15245 (N_15245,N_15146,N_15007);
nor U15246 (N_15246,N_15193,N_15112);
or U15247 (N_15247,N_15032,N_15179);
xor U15248 (N_15248,N_15008,N_15173);
and U15249 (N_15249,N_15144,N_15176);
xor U15250 (N_15250,N_15162,N_15065);
or U15251 (N_15251,N_15189,N_15005);
or U15252 (N_15252,N_15159,N_15094);
nand U15253 (N_15253,N_15168,N_15055);
nor U15254 (N_15254,N_15010,N_15152);
nor U15255 (N_15255,N_15098,N_15117);
xnor U15256 (N_15256,N_15187,N_15093);
xor U15257 (N_15257,N_15070,N_15130);
or U15258 (N_15258,N_15069,N_15132);
and U15259 (N_15259,N_15199,N_15167);
or U15260 (N_15260,N_15085,N_15025);
or U15261 (N_15261,N_15163,N_15056);
xor U15262 (N_15262,N_15157,N_15099);
nand U15263 (N_15263,N_15072,N_15172);
xnor U15264 (N_15264,N_15091,N_15138);
and U15265 (N_15265,N_15141,N_15081);
xnor U15266 (N_15266,N_15030,N_15087);
xor U15267 (N_15267,N_15182,N_15190);
nand U15268 (N_15268,N_15073,N_15028);
or U15269 (N_15269,N_15059,N_15148);
nor U15270 (N_15270,N_15002,N_15078);
nor U15271 (N_15271,N_15041,N_15042);
nand U15272 (N_15272,N_15089,N_15165);
nand U15273 (N_15273,N_15035,N_15170);
nor U15274 (N_15274,N_15071,N_15014);
or U15275 (N_15275,N_15047,N_15020);
nor U15276 (N_15276,N_15083,N_15111);
nand U15277 (N_15277,N_15019,N_15075);
xnor U15278 (N_15278,N_15038,N_15046);
nand U15279 (N_15279,N_15135,N_15026);
and U15280 (N_15280,N_15015,N_15068);
nor U15281 (N_15281,N_15192,N_15114);
and U15282 (N_15282,N_15095,N_15066);
nor U15283 (N_15283,N_15084,N_15045);
and U15284 (N_15284,N_15134,N_15154);
and U15285 (N_15285,N_15021,N_15188);
or U15286 (N_15286,N_15016,N_15057);
xor U15287 (N_15287,N_15100,N_15195);
nor U15288 (N_15288,N_15143,N_15191);
nor U15289 (N_15289,N_15029,N_15080);
nor U15290 (N_15290,N_15139,N_15155);
xor U15291 (N_15291,N_15011,N_15036);
or U15292 (N_15292,N_15086,N_15050);
nor U15293 (N_15293,N_15001,N_15156);
or U15294 (N_15294,N_15184,N_15113);
xor U15295 (N_15295,N_15145,N_15118);
and U15296 (N_15296,N_15198,N_15061);
or U15297 (N_15297,N_15017,N_15031);
or U15298 (N_15298,N_15109,N_15034);
or U15299 (N_15299,N_15022,N_15161);
or U15300 (N_15300,N_15069,N_15163);
and U15301 (N_15301,N_15144,N_15026);
and U15302 (N_15302,N_15184,N_15047);
and U15303 (N_15303,N_15183,N_15169);
or U15304 (N_15304,N_15004,N_15031);
nand U15305 (N_15305,N_15156,N_15136);
nor U15306 (N_15306,N_15143,N_15146);
and U15307 (N_15307,N_15036,N_15059);
nand U15308 (N_15308,N_15102,N_15163);
xor U15309 (N_15309,N_15132,N_15011);
xor U15310 (N_15310,N_15029,N_15098);
nand U15311 (N_15311,N_15094,N_15059);
xor U15312 (N_15312,N_15051,N_15152);
or U15313 (N_15313,N_15179,N_15100);
nand U15314 (N_15314,N_15090,N_15029);
nor U15315 (N_15315,N_15194,N_15034);
nand U15316 (N_15316,N_15181,N_15166);
or U15317 (N_15317,N_15158,N_15177);
xor U15318 (N_15318,N_15082,N_15042);
nand U15319 (N_15319,N_15011,N_15120);
nor U15320 (N_15320,N_15163,N_15132);
and U15321 (N_15321,N_15153,N_15078);
xnor U15322 (N_15322,N_15096,N_15004);
or U15323 (N_15323,N_15127,N_15000);
nor U15324 (N_15324,N_15115,N_15064);
xnor U15325 (N_15325,N_15199,N_15074);
nand U15326 (N_15326,N_15002,N_15180);
and U15327 (N_15327,N_15016,N_15006);
nand U15328 (N_15328,N_15132,N_15084);
and U15329 (N_15329,N_15163,N_15038);
nor U15330 (N_15330,N_15062,N_15056);
or U15331 (N_15331,N_15102,N_15177);
nand U15332 (N_15332,N_15137,N_15080);
or U15333 (N_15333,N_15068,N_15131);
nand U15334 (N_15334,N_15109,N_15164);
nand U15335 (N_15335,N_15064,N_15103);
xor U15336 (N_15336,N_15007,N_15028);
and U15337 (N_15337,N_15169,N_15097);
or U15338 (N_15338,N_15189,N_15104);
nor U15339 (N_15339,N_15092,N_15019);
and U15340 (N_15340,N_15029,N_15112);
xnor U15341 (N_15341,N_15185,N_15084);
xnor U15342 (N_15342,N_15000,N_15174);
nand U15343 (N_15343,N_15023,N_15009);
nor U15344 (N_15344,N_15156,N_15008);
xnor U15345 (N_15345,N_15164,N_15135);
or U15346 (N_15346,N_15118,N_15039);
xor U15347 (N_15347,N_15042,N_15084);
or U15348 (N_15348,N_15043,N_15007);
xor U15349 (N_15349,N_15062,N_15135);
and U15350 (N_15350,N_15079,N_15041);
nand U15351 (N_15351,N_15009,N_15108);
xnor U15352 (N_15352,N_15123,N_15007);
xor U15353 (N_15353,N_15060,N_15029);
xnor U15354 (N_15354,N_15035,N_15017);
or U15355 (N_15355,N_15032,N_15017);
nand U15356 (N_15356,N_15190,N_15173);
xnor U15357 (N_15357,N_15145,N_15037);
nor U15358 (N_15358,N_15135,N_15127);
nand U15359 (N_15359,N_15017,N_15053);
xor U15360 (N_15360,N_15005,N_15061);
xor U15361 (N_15361,N_15103,N_15084);
and U15362 (N_15362,N_15165,N_15112);
and U15363 (N_15363,N_15100,N_15005);
xnor U15364 (N_15364,N_15119,N_15089);
xor U15365 (N_15365,N_15128,N_15044);
nand U15366 (N_15366,N_15004,N_15006);
or U15367 (N_15367,N_15104,N_15030);
or U15368 (N_15368,N_15007,N_15086);
and U15369 (N_15369,N_15010,N_15183);
and U15370 (N_15370,N_15167,N_15006);
and U15371 (N_15371,N_15185,N_15183);
xnor U15372 (N_15372,N_15006,N_15087);
and U15373 (N_15373,N_15083,N_15140);
and U15374 (N_15374,N_15013,N_15111);
nor U15375 (N_15375,N_15181,N_15138);
or U15376 (N_15376,N_15020,N_15140);
xnor U15377 (N_15377,N_15002,N_15169);
or U15378 (N_15378,N_15094,N_15100);
xor U15379 (N_15379,N_15157,N_15031);
xor U15380 (N_15380,N_15110,N_15173);
or U15381 (N_15381,N_15156,N_15172);
and U15382 (N_15382,N_15170,N_15167);
xnor U15383 (N_15383,N_15004,N_15069);
nor U15384 (N_15384,N_15066,N_15034);
or U15385 (N_15385,N_15098,N_15146);
xor U15386 (N_15386,N_15049,N_15166);
and U15387 (N_15387,N_15147,N_15171);
nand U15388 (N_15388,N_15151,N_15106);
and U15389 (N_15389,N_15173,N_15021);
xor U15390 (N_15390,N_15094,N_15024);
nand U15391 (N_15391,N_15021,N_15091);
nand U15392 (N_15392,N_15035,N_15019);
xor U15393 (N_15393,N_15197,N_15009);
xor U15394 (N_15394,N_15010,N_15050);
nand U15395 (N_15395,N_15171,N_15194);
nor U15396 (N_15396,N_15159,N_15143);
nand U15397 (N_15397,N_15001,N_15179);
and U15398 (N_15398,N_15140,N_15067);
or U15399 (N_15399,N_15135,N_15159);
nand U15400 (N_15400,N_15398,N_15358);
and U15401 (N_15401,N_15213,N_15389);
nor U15402 (N_15402,N_15261,N_15320);
or U15403 (N_15403,N_15317,N_15267);
or U15404 (N_15404,N_15342,N_15349);
nand U15405 (N_15405,N_15322,N_15390);
xor U15406 (N_15406,N_15260,N_15396);
and U15407 (N_15407,N_15232,N_15345);
and U15408 (N_15408,N_15235,N_15397);
and U15409 (N_15409,N_15370,N_15343);
nor U15410 (N_15410,N_15333,N_15284);
and U15411 (N_15411,N_15387,N_15354);
and U15412 (N_15412,N_15233,N_15250);
and U15413 (N_15413,N_15236,N_15371);
nor U15414 (N_15414,N_15326,N_15243);
or U15415 (N_15415,N_15339,N_15381);
xnor U15416 (N_15416,N_15265,N_15307);
nand U15417 (N_15417,N_15348,N_15297);
nor U15418 (N_15418,N_15360,N_15292);
or U15419 (N_15419,N_15368,N_15201);
nor U15420 (N_15420,N_15319,N_15399);
and U15421 (N_15421,N_15378,N_15242);
nand U15422 (N_15422,N_15221,N_15227);
nor U15423 (N_15423,N_15309,N_15251);
nor U15424 (N_15424,N_15214,N_15329);
nor U15425 (N_15425,N_15341,N_15335);
nand U15426 (N_15426,N_15324,N_15253);
or U15427 (N_15427,N_15323,N_15287);
xor U15428 (N_15428,N_15388,N_15269);
xor U15429 (N_15429,N_15316,N_15218);
nand U15430 (N_15430,N_15364,N_15392);
and U15431 (N_15431,N_15255,N_15264);
nor U15432 (N_15432,N_15330,N_15222);
or U15433 (N_15433,N_15229,N_15271);
nand U15434 (N_15434,N_15332,N_15248);
and U15435 (N_15435,N_15303,N_15262);
and U15436 (N_15436,N_15268,N_15254);
xor U15437 (N_15437,N_15241,N_15350);
nor U15438 (N_15438,N_15346,N_15247);
or U15439 (N_15439,N_15220,N_15362);
and U15440 (N_15440,N_15312,N_15209);
and U15441 (N_15441,N_15263,N_15270);
xnor U15442 (N_15442,N_15373,N_15274);
nor U15443 (N_15443,N_15304,N_15299);
or U15444 (N_15444,N_15256,N_15377);
xnor U15445 (N_15445,N_15206,N_15257);
xor U15446 (N_15446,N_15286,N_15200);
or U15447 (N_15447,N_15318,N_15234);
and U15448 (N_15448,N_15310,N_15275);
nor U15449 (N_15449,N_15369,N_15203);
nor U15450 (N_15450,N_15308,N_15386);
xor U15451 (N_15451,N_15353,N_15288);
nor U15452 (N_15452,N_15301,N_15283);
nor U15453 (N_15453,N_15336,N_15219);
or U15454 (N_15454,N_15207,N_15295);
and U15455 (N_15455,N_15300,N_15311);
or U15456 (N_15456,N_15212,N_15258);
xnor U15457 (N_15457,N_15216,N_15215);
or U15458 (N_15458,N_15293,N_15249);
nand U15459 (N_15459,N_15372,N_15290);
and U15460 (N_15460,N_15211,N_15347);
xnor U15461 (N_15461,N_15328,N_15305);
and U15462 (N_15462,N_15334,N_15384);
xnor U15463 (N_15463,N_15223,N_15355);
and U15464 (N_15464,N_15266,N_15210);
or U15465 (N_15465,N_15202,N_15325);
xnor U15466 (N_15466,N_15383,N_15224);
nand U15467 (N_15467,N_15291,N_15337);
nor U15468 (N_15468,N_15230,N_15302);
xor U15469 (N_15469,N_15367,N_15273);
or U15470 (N_15470,N_15280,N_15361);
xnor U15471 (N_15471,N_15205,N_15228);
nand U15472 (N_15472,N_15237,N_15289);
or U15473 (N_15473,N_15217,N_15294);
or U15474 (N_15474,N_15357,N_15285);
nor U15475 (N_15475,N_15277,N_15238);
nand U15476 (N_15476,N_15244,N_15296);
xnor U15477 (N_15477,N_15385,N_15239);
nor U15478 (N_15478,N_15315,N_15380);
nand U15479 (N_15479,N_15379,N_15281);
or U15480 (N_15480,N_15225,N_15240);
and U15481 (N_15481,N_15282,N_15204);
xnor U15482 (N_15482,N_15331,N_15338);
nor U15483 (N_15483,N_15344,N_15394);
or U15484 (N_15484,N_15395,N_15382);
nor U15485 (N_15485,N_15252,N_15272);
or U15486 (N_15486,N_15356,N_15391);
or U15487 (N_15487,N_15226,N_15245);
nor U15488 (N_15488,N_15313,N_15321);
nor U15489 (N_15489,N_15375,N_15208);
and U15490 (N_15490,N_15306,N_15246);
nand U15491 (N_15491,N_15352,N_15231);
nand U15492 (N_15492,N_15374,N_15363);
nand U15493 (N_15493,N_15298,N_15259);
nand U15494 (N_15494,N_15359,N_15393);
nand U15495 (N_15495,N_15314,N_15327);
and U15496 (N_15496,N_15376,N_15365);
nor U15497 (N_15497,N_15276,N_15278);
nand U15498 (N_15498,N_15351,N_15366);
or U15499 (N_15499,N_15340,N_15279);
nand U15500 (N_15500,N_15270,N_15352);
xnor U15501 (N_15501,N_15226,N_15270);
and U15502 (N_15502,N_15357,N_15280);
and U15503 (N_15503,N_15320,N_15339);
xnor U15504 (N_15504,N_15309,N_15218);
and U15505 (N_15505,N_15347,N_15350);
or U15506 (N_15506,N_15331,N_15397);
or U15507 (N_15507,N_15258,N_15253);
nor U15508 (N_15508,N_15269,N_15339);
xor U15509 (N_15509,N_15361,N_15383);
or U15510 (N_15510,N_15383,N_15279);
xnor U15511 (N_15511,N_15256,N_15363);
xnor U15512 (N_15512,N_15328,N_15304);
and U15513 (N_15513,N_15329,N_15391);
and U15514 (N_15514,N_15297,N_15386);
and U15515 (N_15515,N_15366,N_15354);
nor U15516 (N_15516,N_15326,N_15351);
xnor U15517 (N_15517,N_15304,N_15247);
and U15518 (N_15518,N_15395,N_15223);
or U15519 (N_15519,N_15243,N_15372);
xor U15520 (N_15520,N_15376,N_15360);
or U15521 (N_15521,N_15248,N_15214);
and U15522 (N_15522,N_15243,N_15271);
or U15523 (N_15523,N_15232,N_15293);
nor U15524 (N_15524,N_15233,N_15372);
or U15525 (N_15525,N_15367,N_15298);
nor U15526 (N_15526,N_15272,N_15331);
xnor U15527 (N_15527,N_15289,N_15219);
and U15528 (N_15528,N_15360,N_15280);
xnor U15529 (N_15529,N_15259,N_15271);
xnor U15530 (N_15530,N_15241,N_15297);
nor U15531 (N_15531,N_15377,N_15305);
xor U15532 (N_15532,N_15287,N_15326);
xnor U15533 (N_15533,N_15255,N_15377);
nor U15534 (N_15534,N_15209,N_15283);
nor U15535 (N_15535,N_15393,N_15368);
xor U15536 (N_15536,N_15332,N_15262);
nor U15537 (N_15537,N_15212,N_15257);
and U15538 (N_15538,N_15259,N_15344);
and U15539 (N_15539,N_15229,N_15200);
xor U15540 (N_15540,N_15342,N_15228);
xor U15541 (N_15541,N_15213,N_15394);
xor U15542 (N_15542,N_15219,N_15392);
and U15543 (N_15543,N_15252,N_15367);
nor U15544 (N_15544,N_15261,N_15311);
or U15545 (N_15545,N_15342,N_15394);
and U15546 (N_15546,N_15321,N_15292);
or U15547 (N_15547,N_15255,N_15252);
and U15548 (N_15548,N_15263,N_15271);
nand U15549 (N_15549,N_15341,N_15249);
and U15550 (N_15550,N_15287,N_15232);
nand U15551 (N_15551,N_15241,N_15335);
nand U15552 (N_15552,N_15393,N_15224);
nand U15553 (N_15553,N_15216,N_15258);
nand U15554 (N_15554,N_15392,N_15333);
or U15555 (N_15555,N_15271,N_15230);
nor U15556 (N_15556,N_15308,N_15292);
or U15557 (N_15557,N_15305,N_15218);
and U15558 (N_15558,N_15215,N_15307);
xor U15559 (N_15559,N_15352,N_15224);
and U15560 (N_15560,N_15386,N_15376);
nand U15561 (N_15561,N_15316,N_15216);
and U15562 (N_15562,N_15212,N_15250);
and U15563 (N_15563,N_15324,N_15243);
or U15564 (N_15564,N_15272,N_15245);
and U15565 (N_15565,N_15263,N_15219);
nor U15566 (N_15566,N_15322,N_15240);
nand U15567 (N_15567,N_15362,N_15372);
nand U15568 (N_15568,N_15214,N_15306);
nand U15569 (N_15569,N_15286,N_15336);
xor U15570 (N_15570,N_15369,N_15370);
nand U15571 (N_15571,N_15303,N_15268);
nand U15572 (N_15572,N_15322,N_15388);
nand U15573 (N_15573,N_15256,N_15388);
xor U15574 (N_15574,N_15361,N_15397);
xor U15575 (N_15575,N_15215,N_15360);
nor U15576 (N_15576,N_15204,N_15315);
nor U15577 (N_15577,N_15313,N_15246);
nor U15578 (N_15578,N_15392,N_15358);
nor U15579 (N_15579,N_15219,N_15300);
nand U15580 (N_15580,N_15215,N_15284);
nor U15581 (N_15581,N_15261,N_15395);
nor U15582 (N_15582,N_15281,N_15269);
and U15583 (N_15583,N_15209,N_15301);
xor U15584 (N_15584,N_15286,N_15334);
nor U15585 (N_15585,N_15236,N_15338);
xnor U15586 (N_15586,N_15205,N_15355);
xnor U15587 (N_15587,N_15388,N_15303);
nand U15588 (N_15588,N_15243,N_15240);
nand U15589 (N_15589,N_15229,N_15316);
nor U15590 (N_15590,N_15392,N_15342);
xnor U15591 (N_15591,N_15272,N_15367);
nand U15592 (N_15592,N_15375,N_15331);
nor U15593 (N_15593,N_15204,N_15347);
nand U15594 (N_15594,N_15325,N_15382);
and U15595 (N_15595,N_15259,N_15289);
or U15596 (N_15596,N_15295,N_15307);
nor U15597 (N_15597,N_15230,N_15322);
and U15598 (N_15598,N_15376,N_15236);
xnor U15599 (N_15599,N_15312,N_15249);
or U15600 (N_15600,N_15447,N_15597);
or U15601 (N_15601,N_15434,N_15472);
nand U15602 (N_15602,N_15431,N_15422);
or U15603 (N_15603,N_15419,N_15408);
nand U15604 (N_15604,N_15494,N_15556);
or U15605 (N_15605,N_15577,N_15443);
or U15606 (N_15606,N_15518,N_15468);
nand U15607 (N_15607,N_15595,N_15473);
nor U15608 (N_15608,N_15437,N_15416);
or U15609 (N_15609,N_15582,N_15414);
or U15610 (N_15610,N_15497,N_15528);
or U15611 (N_15611,N_15533,N_15527);
nand U15612 (N_15612,N_15507,N_15530);
or U15613 (N_15613,N_15482,N_15540);
or U15614 (N_15614,N_15498,N_15409);
nand U15615 (N_15615,N_15546,N_15535);
or U15616 (N_15616,N_15478,N_15561);
xor U15617 (N_15617,N_15519,N_15536);
xor U15618 (N_15618,N_15517,N_15584);
nand U15619 (N_15619,N_15491,N_15513);
xor U15620 (N_15620,N_15407,N_15523);
xnor U15621 (N_15621,N_15558,N_15501);
nand U15622 (N_15622,N_15543,N_15598);
or U15623 (N_15623,N_15538,N_15585);
and U15624 (N_15624,N_15442,N_15544);
or U15625 (N_15625,N_15406,N_15521);
nand U15626 (N_15626,N_15565,N_15547);
nand U15627 (N_15627,N_15426,N_15573);
or U15628 (N_15628,N_15432,N_15554);
and U15629 (N_15629,N_15457,N_15485);
or U15630 (N_15630,N_15508,N_15516);
or U15631 (N_15631,N_15462,N_15435);
xor U15632 (N_15632,N_15571,N_15417);
and U15633 (N_15633,N_15480,N_15496);
or U15634 (N_15634,N_15549,N_15539);
nor U15635 (N_15635,N_15579,N_15487);
nand U15636 (N_15636,N_15504,N_15511);
or U15637 (N_15637,N_15502,N_15402);
nand U15638 (N_15638,N_15476,N_15455);
xnor U15639 (N_15639,N_15505,N_15404);
and U15640 (N_15640,N_15524,N_15529);
and U15641 (N_15641,N_15557,N_15514);
xor U15642 (N_15642,N_15566,N_15492);
xnor U15643 (N_15643,N_15415,N_15403);
and U15644 (N_15644,N_15541,N_15532);
and U15645 (N_15645,N_15474,N_15596);
nor U15646 (N_15646,N_15405,N_15486);
and U15647 (N_15647,N_15465,N_15593);
xnor U15648 (N_15648,N_15428,N_15470);
nand U15649 (N_15649,N_15429,N_15522);
xor U15650 (N_15650,N_15481,N_15545);
xor U15651 (N_15651,N_15548,N_15510);
nor U15652 (N_15652,N_15412,N_15526);
and U15653 (N_15653,N_15564,N_15594);
nand U15654 (N_15654,N_15588,N_15427);
nor U15655 (N_15655,N_15424,N_15423);
nor U15656 (N_15656,N_15438,N_15551);
nor U15657 (N_15657,N_15479,N_15459);
nand U15658 (N_15658,N_15441,N_15440);
nand U15659 (N_15659,N_15568,N_15534);
and U15660 (N_15660,N_15449,N_15591);
and U15661 (N_15661,N_15413,N_15483);
nand U15662 (N_15662,N_15581,N_15460);
xor U15663 (N_15663,N_15587,N_15461);
nor U15664 (N_15664,N_15425,N_15500);
nor U15665 (N_15665,N_15531,N_15467);
and U15666 (N_15666,N_15537,N_15562);
nand U15667 (N_15667,N_15503,N_15477);
and U15668 (N_15668,N_15489,N_15563);
nand U15669 (N_15669,N_15555,N_15574);
nand U15670 (N_15670,N_15401,N_15488);
and U15671 (N_15671,N_15575,N_15410);
nand U15672 (N_15672,N_15430,N_15444);
nor U15673 (N_15673,N_15493,N_15553);
xnor U15674 (N_15674,N_15570,N_15436);
nor U15675 (N_15675,N_15560,N_15475);
or U15676 (N_15676,N_15433,N_15454);
or U15677 (N_15677,N_15506,N_15569);
or U15678 (N_15678,N_15445,N_15471);
and U15679 (N_15679,N_15420,N_15451);
nor U15680 (N_15680,N_15450,N_15515);
or U15681 (N_15681,N_15464,N_15509);
nor U15682 (N_15682,N_15484,N_15463);
nand U15683 (N_15683,N_15439,N_15411);
and U15684 (N_15684,N_15452,N_15499);
xor U15685 (N_15685,N_15495,N_15583);
nand U15686 (N_15686,N_15466,N_15580);
and U15687 (N_15687,N_15458,N_15559);
and U15688 (N_15688,N_15448,N_15421);
nor U15689 (N_15689,N_15446,N_15469);
and U15690 (N_15690,N_15542,N_15578);
xor U15691 (N_15691,N_15453,N_15576);
nor U15692 (N_15692,N_15592,N_15599);
and U15693 (N_15693,N_15550,N_15400);
and U15694 (N_15694,N_15552,N_15456);
nand U15695 (N_15695,N_15520,N_15572);
xor U15696 (N_15696,N_15589,N_15590);
nand U15697 (N_15697,N_15512,N_15490);
and U15698 (N_15698,N_15567,N_15418);
and U15699 (N_15699,N_15525,N_15586);
and U15700 (N_15700,N_15530,N_15451);
and U15701 (N_15701,N_15593,N_15432);
xnor U15702 (N_15702,N_15457,N_15501);
and U15703 (N_15703,N_15537,N_15432);
nor U15704 (N_15704,N_15540,N_15546);
nor U15705 (N_15705,N_15416,N_15433);
xor U15706 (N_15706,N_15546,N_15512);
xnor U15707 (N_15707,N_15468,N_15596);
nand U15708 (N_15708,N_15518,N_15437);
and U15709 (N_15709,N_15521,N_15585);
and U15710 (N_15710,N_15433,N_15599);
or U15711 (N_15711,N_15540,N_15533);
nand U15712 (N_15712,N_15401,N_15570);
nor U15713 (N_15713,N_15540,N_15470);
or U15714 (N_15714,N_15595,N_15520);
and U15715 (N_15715,N_15546,N_15584);
and U15716 (N_15716,N_15532,N_15422);
nand U15717 (N_15717,N_15492,N_15466);
or U15718 (N_15718,N_15563,N_15508);
xor U15719 (N_15719,N_15573,N_15434);
xor U15720 (N_15720,N_15432,N_15431);
or U15721 (N_15721,N_15593,N_15421);
and U15722 (N_15722,N_15480,N_15526);
nand U15723 (N_15723,N_15406,N_15437);
xnor U15724 (N_15724,N_15424,N_15493);
or U15725 (N_15725,N_15520,N_15492);
xor U15726 (N_15726,N_15455,N_15532);
and U15727 (N_15727,N_15431,N_15414);
and U15728 (N_15728,N_15546,N_15530);
xnor U15729 (N_15729,N_15427,N_15469);
nor U15730 (N_15730,N_15545,N_15527);
xnor U15731 (N_15731,N_15443,N_15524);
nand U15732 (N_15732,N_15577,N_15479);
nor U15733 (N_15733,N_15504,N_15456);
and U15734 (N_15734,N_15571,N_15457);
nor U15735 (N_15735,N_15447,N_15587);
nor U15736 (N_15736,N_15565,N_15505);
or U15737 (N_15737,N_15539,N_15491);
nand U15738 (N_15738,N_15536,N_15478);
nor U15739 (N_15739,N_15413,N_15510);
nor U15740 (N_15740,N_15586,N_15500);
xor U15741 (N_15741,N_15595,N_15528);
nand U15742 (N_15742,N_15498,N_15447);
or U15743 (N_15743,N_15575,N_15488);
xnor U15744 (N_15744,N_15429,N_15414);
or U15745 (N_15745,N_15536,N_15550);
nand U15746 (N_15746,N_15441,N_15514);
or U15747 (N_15747,N_15591,N_15467);
nor U15748 (N_15748,N_15503,N_15561);
nand U15749 (N_15749,N_15548,N_15516);
nor U15750 (N_15750,N_15521,N_15477);
xor U15751 (N_15751,N_15568,N_15535);
nor U15752 (N_15752,N_15406,N_15578);
or U15753 (N_15753,N_15420,N_15578);
nand U15754 (N_15754,N_15486,N_15400);
nand U15755 (N_15755,N_15429,N_15496);
xnor U15756 (N_15756,N_15533,N_15460);
nor U15757 (N_15757,N_15495,N_15558);
and U15758 (N_15758,N_15443,N_15547);
nand U15759 (N_15759,N_15433,N_15438);
nor U15760 (N_15760,N_15432,N_15477);
nor U15761 (N_15761,N_15486,N_15437);
nor U15762 (N_15762,N_15412,N_15488);
and U15763 (N_15763,N_15538,N_15473);
xor U15764 (N_15764,N_15427,N_15580);
and U15765 (N_15765,N_15401,N_15499);
xor U15766 (N_15766,N_15462,N_15508);
nor U15767 (N_15767,N_15565,N_15446);
nand U15768 (N_15768,N_15572,N_15560);
nand U15769 (N_15769,N_15411,N_15557);
or U15770 (N_15770,N_15517,N_15480);
and U15771 (N_15771,N_15580,N_15419);
nand U15772 (N_15772,N_15429,N_15471);
or U15773 (N_15773,N_15535,N_15429);
nor U15774 (N_15774,N_15577,N_15533);
nand U15775 (N_15775,N_15525,N_15584);
nand U15776 (N_15776,N_15528,N_15413);
and U15777 (N_15777,N_15418,N_15474);
or U15778 (N_15778,N_15523,N_15471);
nand U15779 (N_15779,N_15403,N_15452);
nor U15780 (N_15780,N_15439,N_15446);
or U15781 (N_15781,N_15591,N_15404);
nor U15782 (N_15782,N_15529,N_15495);
or U15783 (N_15783,N_15523,N_15541);
and U15784 (N_15784,N_15491,N_15403);
nand U15785 (N_15785,N_15514,N_15488);
and U15786 (N_15786,N_15551,N_15452);
or U15787 (N_15787,N_15582,N_15563);
and U15788 (N_15788,N_15576,N_15594);
nor U15789 (N_15789,N_15405,N_15465);
nand U15790 (N_15790,N_15417,N_15481);
and U15791 (N_15791,N_15403,N_15542);
and U15792 (N_15792,N_15587,N_15474);
or U15793 (N_15793,N_15512,N_15554);
or U15794 (N_15794,N_15527,N_15554);
nor U15795 (N_15795,N_15588,N_15574);
nor U15796 (N_15796,N_15496,N_15481);
and U15797 (N_15797,N_15592,N_15490);
nor U15798 (N_15798,N_15519,N_15573);
xor U15799 (N_15799,N_15555,N_15444);
nand U15800 (N_15800,N_15743,N_15733);
xnor U15801 (N_15801,N_15674,N_15642);
nor U15802 (N_15802,N_15604,N_15671);
and U15803 (N_15803,N_15727,N_15770);
nor U15804 (N_15804,N_15600,N_15618);
nand U15805 (N_15805,N_15632,N_15644);
nand U15806 (N_15806,N_15658,N_15657);
and U15807 (N_15807,N_15752,N_15746);
and U15808 (N_15808,N_15608,N_15641);
nand U15809 (N_15809,N_15755,N_15653);
nand U15810 (N_15810,N_15615,N_15664);
xor U15811 (N_15811,N_15612,N_15738);
and U15812 (N_15812,N_15617,N_15648);
and U15813 (N_15813,N_15799,N_15702);
xnor U15814 (N_15814,N_15790,N_15669);
or U15815 (N_15815,N_15601,N_15781);
nor U15816 (N_15816,N_15668,N_15689);
and U15817 (N_15817,N_15791,N_15663);
xor U15818 (N_15818,N_15767,N_15715);
or U15819 (N_15819,N_15602,N_15623);
nor U15820 (N_15820,N_15643,N_15740);
xor U15821 (N_15821,N_15724,N_15704);
or U15822 (N_15822,N_15652,N_15798);
and U15823 (N_15823,N_15741,N_15666);
nand U15824 (N_15824,N_15645,N_15751);
and U15825 (N_15825,N_15711,N_15782);
nor U15826 (N_15826,N_15695,N_15766);
xnor U15827 (N_15827,N_15759,N_15661);
or U15828 (N_15828,N_15678,N_15605);
nor U15829 (N_15829,N_15705,N_15613);
nor U15830 (N_15830,N_15684,N_15688);
nor U15831 (N_15831,N_15628,N_15655);
nor U15832 (N_15832,N_15725,N_15774);
or U15833 (N_15833,N_15780,N_15750);
nand U15834 (N_15834,N_15619,N_15764);
and U15835 (N_15835,N_15636,N_15673);
or U15836 (N_15836,N_15679,N_15776);
and U15837 (N_15837,N_15614,N_15718);
nand U15838 (N_15838,N_15756,N_15685);
nor U15839 (N_15839,N_15789,N_15795);
or U15840 (N_15840,N_15620,N_15728);
and U15841 (N_15841,N_15659,N_15682);
nor U15842 (N_15842,N_15754,N_15701);
and U15843 (N_15843,N_15749,N_15650);
nor U15844 (N_15844,N_15649,N_15792);
xnor U15845 (N_15845,N_15730,N_15622);
xor U15846 (N_15846,N_15700,N_15630);
and U15847 (N_15847,N_15680,N_15626);
nand U15848 (N_15848,N_15635,N_15773);
or U15849 (N_15849,N_15771,N_15697);
nand U15850 (N_15850,N_15670,N_15777);
or U15851 (N_15851,N_15775,N_15656);
xnor U15852 (N_15852,N_15772,N_15762);
or U15853 (N_15853,N_15698,N_15717);
nor U15854 (N_15854,N_15735,N_15758);
and U15855 (N_15855,N_15634,N_15676);
nand U15856 (N_15856,N_15760,N_15786);
xor U15857 (N_15857,N_15721,N_15651);
xnor U15858 (N_15858,N_15763,N_15631);
xor U15859 (N_15859,N_15796,N_15637);
and U15860 (N_15860,N_15753,N_15744);
nor U15861 (N_15861,N_15709,N_15739);
xnor U15862 (N_15862,N_15687,N_15625);
and U15863 (N_15863,N_15660,N_15633);
or U15864 (N_15864,N_15616,N_15765);
xor U15865 (N_15865,N_15640,N_15693);
xnor U15866 (N_15866,N_15797,N_15779);
or U15867 (N_15867,N_15610,N_15794);
or U15868 (N_15868,N_15785,N_15624);
nor U15869 (N_15869,N_15742,N_15707);
nand U15870 (N_15870,N_15647,N_15665);
nor U15871 (N_15871,N_15731,N_15722);
or U15872 (N_15872,N_15716,N_15606);
and U15873 (N_15873,N_15694,N_15607);
xnor U15874 (N_15874,N_15603,N_15748);
nand U15875 (N_15875,N_15706,N_15691);
and U15876 (N_15876,N_15736,N_15646);
nand U15877 (N_15877,N_15783,N_15690);
xnor U15878 (N_15878,N_15611,N_15708);
or U15879 (N_15879,N_15692,N_15720);
nand U15880 (N_15880,N_15769,N_15788);
nor U15881 (N_15881,N_15714,N_15703);
and U15882 (N_15882,N_15729,N_15726);
or U15883 (N_15883,N_15757,N_15677);
nor U15884 (N_15884,N_15638,N_15745);
xor U15885 (N_15885,N_15732,N_15734);
nand U15886 (N_15886,N_15654,N_15683);
xor U15887 (N_15887,N_15662,N_15787);
nand U15888 (N_15888,N_15667,N_15621);
xor U15889 (N_15889,N_15629,N_15719);
and U15890 (N_15890,N_15609,N_15784);
nor U15891 (N_15891,N_15686,N_15672);
xor U15892 (N_15892,N_15699,N_15713);
or U15893 (N_15893,N_15723,N_15712);
and U15894 (N_15894,N_15793,N_15675);
xor U15895 (N_15895,N_15696,N_15681);
and U15896 (N_15896,N_15627,N_15747);
and U15897 (N_15897,N_15737,N_15639);
nand U15898 (N_15898,N_15761,N_15710);
nor U15899 (N_15899,N_15778,N_15768);
xnor U15900 (N_15900,N_15768,N_15647);
or U15901 (N_15901,N_15704,N_15661);
and U15902 (N_15902,N_15669,N_15763);
nand U15903 (N_15903,N_15682,N_15683);
nor U15904 (N_15904,N_15704,N_15677);
and U15905 (N_15905,N_15744,N_15724);
nor U15906 (N_15906,N_15785,N_15648);
xor U15907 (N_15907,N_15741,N_15705);
or U15908 (N_15908,N_15624,N_15737);
nor U15909 (N_15909,N_15750,N_15623);
nand U15910 (N_15910,N_15780,N_15733);
xor U15911 (N_15911,N_15781,N_15610);
or U15912 (N_15912,N_15793,N_15703);
nor U15913 (N_15913,N_15714,N_15610);
nand U15914 (N_15914,N_15746,N_15609);
and U15915 (N_15915,N_15747,N_15601);
or U15916 (N_15916,N_15762,N_15799);
nand U15917 (N_15917,N_15779,N_15722);
nor U15918 (N_15918,N_15635,N_15616);
nor U15919 (N_15919,N_15717,N_15641);
and U15920 (N_15920,N_15772,N_15620);
nor U15921 (N_15921,N_15641,N_15776);
or U15922 (N_15922,N_15663,N_15692);
and U15923 (N_15923,N_15666,N_15638);
or U15924 (N_15924,N_15690,N_15781);
or U15925 (N_15925,N_15707,N_15660);
and U15926 (N_15926,N_15661,N_15794);
xnor U15927 (N_15927,N_15655,N_15672);
and U15928 (N_15928,N_15663,N_15615);
or U15929 (N_15929,N_15679,N_15613);
xnor U15930 (N_15930,N_15607,N_15618);
nand U15931 (N_15931,N_15689,N_15612);
xnor U15932 (N_15932,N_15798,N_15662);
nor U15933 (N_15933,N_15624,N_15714);
xnor U15934 (N_15934,N_15662,N_15648);
or U15935 (N_15935,N_15721,N_15657);
xnor U15936 (N_15936,N_15698,N_15607);
and U15937 (N_15937,N_15760,N_15750);
xnor U15938 (N_15938,N_15733,N_15761);
xor U15939 (N_15939,N_15702,N_15766);
nand U15940 (N_15940,N_15715,N_15693);
nand U15941 (N_15941,N_15620,N_15747);
nand U15942 (N_15942,N_15771,N_15628);
xor U15943 (N_15943,N_15633,N_15609);
nor U15944 (N_15944,N_15720,N_15611);
xnor U15945 (N_15945,N_15719,N_15756);
and U15946 (N_15946,N_15657,N_15743);
nand U15947 (N_15947,N_15710,N_15648);
nand U15948 (N_15948,N_15681,N_15742);
xnor U15949 (N_15949,N_15635,N_15644);
xnor U15950 (N_15950,N_15794,N_15703);
and U15951 (N_15951,N_15709,N_15681);
nand U15952 (N_15952,N_15675,N_15612);
nor U15953 (N_15953,N_15654,N_15632);
and U15954 (N_15954,N_15695,N_15739);
nand U15955 (N_15955,N_15722,N_15729);
nand U15956 (N_15956,N_15789,N_15622);
and U15957 (N_15957,N_15697,N_15729);
xor U15958 (N_15958,N_15688,N_15627);
xnor U15959 (N_15959,N_15736,N_15645);
xnor U15960 (N_15960,N_15726,N_15663);
nor U15961 (N_15961,N_15660,N_15790);
nor U15962 (N_15962,N_15655,N_15747);
and U15963 (N_15963,N_15788,N_15732);
and U15964 (N_15964,N_15666,N_15703);
nor U15965 (N_15965,N_15626,N_15772);
xor U15966 (N_15966,N_15640,N_15742);
nand U15967 (N_15967,N_15784,N_15620);
or U15968 (N_15968,N_15674,N_15614);
nand U15969 (N_15969,N_15769,N_15669);
or U15970 (N_15970,N_15729,N_15629);
nor U15971 (N_15971,N_15724,N_15665);
or U15972 (N_15972,N_15608,N_15703);
nor U15973 (N_15973,N_15717,N_15728);
nor U15974 (N_15974,N_15640,N_15653);
or U15975 (N_15975,N_15606,N_15787);
or U15976 (N_15976,N_15666,N_15671);
and U15977 (N_15977,N_15752,N_15767);
and U15978 (N_15978,N_15656,N_15689);
nand U15979 (N_15979,N_15775,N_15791);
and U15980 (N_15980,N_15641,N_15761);
or U15981 (N_15981,N_15729,N_15673);
or U15982 (N_15982,N_15655,N_15754);
xor U15983 (N_15983,N_15770,N_15787);
and U15984 (N_15984,N_15634,N_15621);
and U15985 (N_15985,N_15608,N_15638);
or U15986 (N_15986,N_15706,N_15683);
nand U15987 (N_15987,N_15693,N_15775);
and U15988 (N_15988,N_15796,N_15625);
nand U15989 (N_15989,N_15617,N_15694);
xnor U15990 (N_15990,N_15717,N_15776);
nand U15991 (N_15991,N_15681,N_15741);
xor U15992 (N_15992,N_15650,N_15634);
nand U15993 (N_15993,N_15768,N_15601);
nand U15994 (N_15994,N_15730,N_15715);
nor U15995 (N_15995,N_15770,N_15719);
or U15996 (N_15996,N_15629,N_15787);
and U15997 (N_15997,N_15686,N_15677);
xnor U15998 (N_15998,N_15667,N_15616);
nor U15999 (N_15999,N_15749,N_15743);
xnor U16000 (N_16000,N_15938,N_15978);
xnor U16001 (N_16001,N_15895,N_15896);
or U16002 (N_16002,N_15839,N_15875);
nor U16003 (N_16003,N_15937,N_15921);
or U16004 (N_16004,N_15997,N_15821);
nand U16005 (N_16005,N_15856,N_15946);
nor U16006 (N_16006,N_15909,N_15907);
nor U16007 (N_16007,N_15905,N_15925);
xor U16008 (N_16008,N_15805,N_15927);
or U16009 (N_16009,N_15986,N_15918);
xor U16010 (N_16010,N_15928,N_15852);
or U16011 (N_16011,N_15824,N_15913);
or U16012 (N_16012,N_15923,N_15823);
and U16013 (N_16013,N_15877,N_15902);
or U16014 (N_16014,N_15843,N_15813);
xor U16015 (N_16015,N_15848,N_15984);
nor U16016 (N_16016,N_15903,N_15936);
xnor U16017 (N_16017,N_15939,N_15948);
nand U16018 (N_16018,N_15947,N_15945);
xnor U16019 (N_16019,N_15959,N_15952);
and U16020 (N_16020,N_15870,N_15956);
nor U16021 (N_16021,N_15942,N_15960);
nor U16022 (N_16022,N_15804,N_15838);
and U16023 (N_16023,N_15811,N_15842);
or U16024 (N_16024,N_15964,N_15957);
nand U16025 (N_16025,N_15915,N_15916);
or U16026 (N_16026,N_15985,N_15990);
nand U16027 (N_16027,N_15841,N_15994);
nand U16028 (N_16028,N_15965,N_15963);
nand U16029 (N_16029,N_15887,N_15967);
xnor U16030 (N_16030,N_15835,N_15966);
or U16031 (N_16031,N_15800,N_15981);
nor U16032 (N_16032,N_15815,N_15836);
and U16033 (N_16033,N_15934,N_15866);
nand U16034 (N_16034,N_15961,N_15943);
or U16035 (N_16035,N_15980,N_15874);
or U16036 (N_16036,N_15944,N_15847);
nand U16037 (N_16037,N_15924,N_15975);
nand U16038 (N_16038,N_15954,N_15914);
or U16039 (N_16039,N_15894,N_15880);
or U16040 (N_16040,N_15970,N_15968);
nor U16041 (N_16041,N_15814,N_15910);
xor U16042 (N_16042,N_15816,N_15817);
or U16043 (N_16043,N_15865,N_15859);
nand U16044 (N_16044,N_15897,N_15893);
and U16045 (N_16045,N_15806,N_15993);
nor U16046 (N_16046,N_15983,N_15830);
and U16047 (N_16047,N_15818,N_15969);
xnor U16048 (N_16048,N_15860,N_15809);
xnor U16049 (N_16049,N_15955,N_15958);
nand U16050 (N_16050,N_15920,N_15857);
xor U16051 (N_16051,N_15844,N_15876);
nand U16052 (N_16052,N_15881,N_15884);
xor U16053 (N_16053,N_15826,N_15855);
nor U16054 (N_16054,N_15850,N_15917);
and U16055 (N_16055,N_15930,N_15892);
xnor U16056 (N_16056,N_15845,N_15971);
and U16057 (N_16057,N_15995,N_15974);
or U16058 (N_16058,N_15831,N_15940);
xnor U16059 (N_16059,N_15950,N_15822);
nand U16060 (N_16060,N_15911,N_15849);
or U16061 (N_16061,N_15863,N_15882);
nor U16062 (N_16062,N_15941,N_15825);
and U16063 (N_16063,N_15977,N_15899);
xnor U16064 (N_16064,N_15868,N_15901);
or U16065 (N_16065,N_15982,N_15932);
xnor U16066 (N_16066,N_15992,N_15854);
nand U16067 (N_16067,N_15951,N_15929);
or U16068 (N_16068,N_15987,N_15908);
or U16069 (N_16069,N_15931,N_15890);
and U16070 (N_16070,N_15869,N_15837);
xnor U16071 (N_16071,N_15953,N_15832);
xor U16072 (N_16072,N_15834,N_15900);
nor U16073 (N_16073,N_15829,N_15888);
and U16074 (N_16074,N_15996,N_15807);
and U16075 (N_16075,N_15889,N_15879);
xnor U16076 (N_16076,N_15808,N_15933);
and U16077 (N_16077,N_15904,N_15926);
nor U16078 (N_16078,N_15872,N_15853);
xor U16079 (N_16079,N_15801,N_15886);
or U16080 (N_16080,N_15802,N_15828);
xor U16081 (N_16081,N_15988,N_15864);
nor U16082 (N_16082,N_15867,N_15906);
or U16083 (N_16083,N_15871,N_15810);
or U16084 (N_16084,N_15861,N_15919);
nand U16085 (N_16085,N_15812,N_15922);
xnor U16086 (N_16086,N_15885,N_15803);
or U16087 (N_16087,N_15998,N_15827);
xor U16088 (N_16088,N_15989,N_15846);
or U16089 (N_16089,N_15972,N_15878);
nor U16090 (N_16090,N_15883,N_15840);
nor U16091 (N_16091,N_15891,N_15912);
xor U16092 (N_16092,N_15976,N_15949);
xnor U16093 (N_16093,N_15873,N_15973);
or U16094 (N_16094,N_15991,N_15858);
nand U16095 (N_16095,N_15819,N_15935);
xor U16096 (N_16096,N_15833,N_15962);
and U16097 (N_16097,N_15979,N_15898);
or U16098 (N_16098,N_15999,N_15851);
nor U16099 (N_16099,N_15862,N_15820);
nand U16100 (N_16100,N_15881,N_15905);
nor U16101 (N_16101,N_15857,N_15867);
or U16102 (N_16102,N_15902,N_15813);
nand U16103 (N_16103,N_15996,N_15925);
and U16104 (N_16104,N_15984,N_15859);
nor U16105 (N_16105,N_15862,N_15821);
xnor U16106 (N_16106,N_15884,N_15994);
nand U16107 (N_16107,N_15853,N_15930);
and U16108 (N_16108,N_15820,N_15993);
nor U16109 (N_16109,N_15904,N_15934);
and U16110 (N_16110,N_15841,N_15892);
xor U16111 (N_16111,N_15806,N_15824);
and U16112 (N_16112,N_15831,N_15893);
nand U16113 (N_16113,N_15909,N_15826);
nand U16114 (N_16114,N_15909,N_15980);
and U16115 (N_16115,N_15993,N_15827);
or U16116 (N_16116,N_15998,N_15938);
xnor U16117 (N_16117,N_15831,N_15858);
xnor U16118 (N_16118,N_15991,N_15838);
xnor U16119 (N_16119,N_15953,N_15906);
nand U16120 (N_16120,N_15922,N_15800);
nor U16121 (N_16121,N_15851,N_15905);
nand U16122 (N_16122,N_15912,N_15875);
xor U16123 (N_16123,N_15980,N_15822);
or U16124 (N_16124,N_15904,N_15930);
and U16125 (N_16125,N_15881,N_15917);
or U16126 (N_16126,N_15959,N_15909);
nor U16127 (N_16127,N_15897,N_15877);
nor U16128 (N_16128,N_15916,N_15842);
or U16129 (N_16129,N_15976,N_15812);
nor U16130 (N_16130,N_15915,N_15974);
nand U16131 (N_16131,N_15814,N_15811);
or U16132 (N_16132,N_15892,N_15980);
and U16133 (N_16133,N_15832,N_15985);
nand U16134 (N_16134,N_15893,N_15946);
and U16135 (N_16135,N_15868,N_15811);
and U16136 (N_16136,N_15856,N_15884);
and U16137 (N_16137,N_15832,N_15840);
and U16138 (N_16138,N_15872,N_15823);
nand U16139 (N_16139,N_15816,N_15981);
nor U16140 (N_16140,N_15802,N_15854);
nand U16141 (N_16141,N_15827,N_15912);
xor U16142 (N_16142,N_15838,N_15980);
xor U16143 (N_16143,N_15855,N_15907);
nor U16144 (N_16144,N_15837,N_15812);
nor U16145 (N_16145,N_15873,N_15879);
and U16146 (N_16146,N_15836,N_15933);
xnor U16147 (N_16147,N_15836,N_15928);
and U16148 (N_16148,N_15983,N_15809);
xor U16149 (N_16149,N_15807,N_15999);
xor U16150 (N_16150,N_15998,N_15926);
or U16151 (N_16151,N_15869,N_15828);
nand U16152 (N_16152,N_15805,N_15847);
or U16153 (N_16153,N_15866,N_15912);
nand U16154 (N_16154,N_15986,N_15847);
nand U16155 (N_16155,N_15922,N_15976);
nand U16156 (N_16156,N_15980,N_15829);
nor U16157 (N_16157,N_15819,N_15967);
xor U16158 (N_16158,N_15811,N_15805);
nor U16159 (N_16159,N_15938,N_15844);
nand U16160 (N_16160,N_15815,N_15801);
or U16161 (N_16161,N_15806,N_15877);
xor U16162 (N_16162,N_15849,N_15860);
nand U16163 (N_16163,N_15877,N_15903);
nand U16164 (N_16164,N_15913,N_15838);
or U16165 (N_16165,N_15928,N_15946);
and U16166 (N_16166,N_15881,N_15940);
xnor U16167 (N_16167,N_15811,N_15844);
nand U16168 (N_16168,N_15824,N_15846);
and U16169 (N_16169,N_15938,N_15889);
xnor U16170 (N_16170,N_15991,N_15845);
xor U16171 (N_16171,N_15840,N_15868);
nor U16172 (N_16172,N_15844,N_15872);
nor U16173 (N_16173,N_15951,N_15932);
nor U16174 (N_16174,N_15878,N_15871);
nor U16175 (N_16175,N_15962,N_15984);
and U16176 (N_16176,N_15927,N_15988);
nor U16177 (N_16177,N_15809,N_15869);
xnor U16178 (N_16178,N_15873,N_15823);
nand U16179 (N_16179,N_15944,N_15870);
or U16180 (N_16180,N_15856,N_15952);
nor U16181 (N_16181,N_15853,N_15999);
xor U16182 (N_16182,N_15810,N_15962);
and U16183 (N_16183,N_15915,N_15999);
nand U16184 (N_16184,N_15950,N_15804);
xor U16185 (N_16185,N_15851,N_15979);
xor U16186 (N_16186,N_15808,N_15923);
or U16187 (N_16187,N_15950,N_15905);
and U16188 (N_16188,N_15886,N_15831);
and U16189 (N_16189,N_15910,N_15895);
nor U16190 (N_16190,N_15900,N_15925);
or U16191 (N_16191,N_15885,N_15953);
nand U16192 (N_16192,N_15803,N_15988);
xnor U16193 (N_16193,N_15956,N_15884);
nand U16194 (N_16194,N_15935,N_15920);
or U16195 (N_16195,N_15803,N_15903);
xnor U16196 (N_16196,N_15852,N_15821);
nand U16197 (N_16197,N_15946,N_15802);
nor U16198 (N_16198,N_15804,N_15883);
xnor U16199 (N_16199,N_15886,N_15978);
nor U16200 (N_16200,N_16084,N_16105);
xor U16201 (N_16201,N_16082,N_16020);
nor U16202 (N_16202,N_16063,N_16030);
or U16203 (N_16203,N_16095,N_16035);
nand U16204 (N_16204,N_16191,N_16012);
or U16205 (N_16205,N_16056,N_16041);
or U16206 (N_16206,N_16036,N_16042);
nand U16207 (N_16207,N_16178,N_16026);
and U16208 (N_16208,N_16138,N_16183);
or U16209 (N_16209,N_16137,N_16145);
and U16210 (N_16210,N_16007,N_16108);
or U16211 (N_16211,N_16112,N_16081);
or U16212 (N_16212,N_16061,N_16047);
nand U16213 (N_16213,N_16045,N_16064);
nand U16214 (N_16214,N_16051,N_16163);
and U16215 (N_16215,N_16087,N_16156);
nand U16216 (N_16216,N_16185,N_16129);
nand U16217 (N_16217,N_16008,N_16148);
nor U16218 (N_16218,N_16066,N_16161);
nor U16219 (N_16219,N_16104,N_16194);
xnor U16220 (N_16220,N_16062,N_16180);
nor U16221 (N_16221,N_16027,N_16141);
or U16222 (N_16222,N_16155,N_16109);
nand U16223 (N_16223,N_16015,N_16044);
nor U16224 (N_16224,N_16014,N_16039);
or U16225 (N_16225,N_16181,N_16147);
and U16226 (N_16226,N_16009,N_16059);
xnor U16227 (N_16227,N_16174,N_16072);
nor U16228 (N_16228,N_16043,N_16170);
nor U16229 (N_16229,N_16077,N_16005);
nor U16230 (N_16230,N_16193,N_16037);
xor U16231 (N_16231,N_16158,N_16190);
nor U16232 (N_16232,N_16151,N_16143);
xnor U16233 (N_16233,N_16118,N_16052);
and U16234 (N_16234,N_16177,N_16149);
nor U16235 (N_16235,N_16090,N_16013);
nand U16236 (N_16236,N_16079,N_16127);
nand U16237 (N_16237,N_16176,N_16167);
and U16238 (N_16238,N_16164,N_16093);
nor U16239 (N_16239,N_16102,N_16006);
nand U16240 (N_16240,N_16186,N_16133);
or U16241 (N_16241,N_16154,N_16004);
nor U16242 (N_16242,N_16049,N_16113);
or U16243 (N_16243,N_16131,N_16182);
and U16244 (N_16244,N_16083,N_16116);
and U16245 (N_16245,N_16085,N_16075);
or U16246 (N_16246,N_16139,N_16175);
xnor U16247 (N_16247,N_16057,N_16073);
nor U16248 (N_16248,N_16126,N_16123);
or U16249 (N_16249,N_16146,N_16196);
or U16250 (N_16250,N_16120,N_16136);
or U16251 (N_16251,N_16162,N_16103);
xor U16252 (N_16252,N_16010,N_16157);
nor U16253 (N_16253,N_16099,N_16018);
xor U16254 (N_16254,N_16048,N_16021);
or U16255 (N_16255,N_16184,N_16098);
xnor U16256 (N_16256,N_16001,N_16074);
and U16257 (N_16257,N_16058,N_16144);
and U16258 (N_16258,N_16195,N_16140);
and U16259 (N_16259,N_16187,N_16189);
nand U16260 (N_16260,N_16171,N_16069);
and U16261 (N_16261,N_16038,N_16022);
nor U16262 (N_16262,N_16115,N_16086);
or U16263 (N_16263,N_16053,N_16122);
or U16264 (N_16264,N_16078,N_16111);
xnor U16265 (N_16265,N_16179,N_16097);
nor U16266 (N_16266,N_16152,N_16169);
or U16267 (N_16267,N_16031,N_16130);
or U16268 (N_16268,N_16166,N_16100);
nand U16269 (N_16269,N_16150,N_16165);
and U16270 (N_16270,N_16071,N_16132);
nor U16271 (N_16271,N_16067,N_16055);
xnor U16272 (N_16272,N_16068,N_16024);
and U16273 (N_16273,N_16107,N_16076);
and U16274 (N_16274,N_16199,N_16094);
xor U16275 (N_16275,N_16125,N_16114);
xnor U16276 (N_16276,N_16160,N_16159);
nand U16277 (N_16277,N_16070,N_16142);
nand U16278 (N_16278,N_16032,N_16197);
and U16279 (N_16279,N_16054,N_16119);
and U16280 (N_16280,N_16023,N_16106);
xnor U16281 (N_16281,N_16019,N_16025);
or U16282 (N_16282,N_16117,N_16168);
xnor U16283 (N_16283,N_16080,N_16065);
nor U16284 (N_16284,N_16017,N_16016);
and U16285 (N_16285,N_16034,N_16003);
nor U16286 (N_16286,N_16198,N_16046);
nor U16287 (N_16287,N_16096,N_16124);
or U16288 (N_16288,N_16121,N_16029);
nor U16289 (N_16289,N_16060,N_16101);
or U16290 (N_16290,N_16135,N_16040);
nand U16291 (N_16291,N_16011,N_16088);
nand U16292 (N_16292,N_16089,N_16188);
and U16293 (N_16293,N_16000,N_16153);
xor U16294 (N_16294,N_16173,N_16110);
nand U16295 (N_16295,N_16092,N_16134);
nor U16296 (N_16296,N_16033,N_16091);
xnor U16297 (N_16297,N_16128,N_16172);
and U16298 (N_16298,N_16050,N_16028);
nand U16299 (N_16299,N_16002,N_16192);
xor U16300 (N_16300,N_16145,N_16010);
or U16301 (N_16301,N_16132,N_16036);
nor U16302 (N_16302,N_16103,N_16046);
or U16303 (N_16303,N_16182,N_16020);
nand U16304 (N_16304,N_16196,N_16093);
nor U16305 (N_16305,N_16019,N_16013);
nor U16306 (N_16306,N_16138,N_16186);
and U16307 (N_16307,N_16063,N_16077);
or U16308 (N_16308,N_16192,N_16067);
and U16309 (N_16309,N_16156,N_16095);
or U16310 (N_16310,N_16065,N_16111);
nand U16311 (N_16311,N_16040,N_16154);
nor U16312 (N_16312,N_16159,N_16136);
and U16313 (N_16313,N_16176,N_16194);
or U16314 (N_16314,N_16051,N_16084);
or U16315 (N_16315,N_16177,N_16140);
xor U16316 (N_16316,N_16143,N_16145);
nand U16317 (N_16317,N_16154,N_16092);
nor U16318 (N_16318,N_16109,N_16153);
nor U16319 (N_16319,N_16056,N_16034);
nor U16320 (N_16320,N_16049,N_16027);
xor U16321 (N_16321,N_16021,N_16009);
and U16322 (N_16322,N_16067,N_16111);
nor U16323 (N_16323,N_16112,N_16197);
and U16324 (N_16324,N_16166,N_16142);
and U16325 (N_16325,N_16160,N_16194);
or U16326 (N_16326,N_16023,N_16140);
and U16327 (N_16327,N_16045,N_16047);
nand U16328 (N_16328,N_16061,N_16074);
or U16329 (N_16329,N_16108,N_16190);
or U16330 (N_16330,N_16039,N_16023);
xor U16331 (N_16331,N_16042,N_16103);
nor U16332 (N_16332,N_16175,N_16183);
nor U16333 (N_16333,N_16134,N_16013);
nor U16334 (N_16334,N_16086,N_16018);
or U16335 (N_16335,N_16190,N_16077);
nand U16336 (N_16336,N_16078,N_16023);
nand U16337 (N_16337,N_16098,N_16162);
xnor U16338 (N_16338,N_16187,N_16030);
nand U16339 (N_16339,N_16110,N_16192);
xnor U16340 (N_16340,N_16074,N_16186);
or U16341 (N_16341,N_16199,N_16132);
nor U16342 (N_16342,N_16070,N_16066);
or U16343 (N_16343,N_16115,N_16199);
and U16344 (N_16344,N_16032,N_16042);
xnor U16345 (N_16345,N_16002,N_16000);
xor U16346 (N_16346,N_16113,N_16136);
nand U16347 (N_16347,N_16004,N_16119);
xor U16348 (N_16348,N_16116,N_16154);
and U16349 (N_16349,N_16184,N_16165);
xor U16350 (N_16350,N_16190,N_16023);
and U16351 (N_16351,N_16081,N_16079);
and U16352 (N_16352,N_16158,N_16063);
nand U16353 (N_16353,N_16170,N_16180);
xnor U16354 (N_16354,N_16105,N_16110);
and U16355 (N_16355,N_16159,N_16172);
nand U16356 (N_16356,N_16005,N_16083);
and U16357 (N_16357,N_16054,N_16160);
or U16358 (N_16358,N_16004,N_16112);
xor U16359 (N_16359,N_16198,N_16150);
and U16360 (N_16360,N_16022,N_16092);
and U16361 (N_16361,N_16098,N_16136);
or U16362 (N_16362,N_16058,N_16097);
and U16363 (N_16363,N_16102,N_16061);
xor U16364 (N_16364,N_16110,N_16030);
nand U16365 (N_16365,N_16008,N_16093);
nor U16366 (N_16366,N_16120,N_16002);
nand U16367 (N_16367,N_16103,N_16149);
xor U16368 (N_16368,N_16026,N_16153);
nor U16369 (N_16369,N_16070,N_16030);
nand U16370 (N_16370,N_16178,N_16185);
xor U16371 (N_16371,N_16031,N_16040);
and U16372 (N_16372,N_16192,N_16196);
or U16373 (N_16373,N_16018,N_16075);
xor U16374 (N_16374,N_16006,N_16111);
nor U16375 (N_16375,N_16065,N_16009);
xnor U16376 (N_16376,N_16074,N_16133);
nor U16377 (N_16377,N_16062,N_16032);
and U16378 (N_16378,N_16163,N_16059);
nor U16379 (N_16379,N_16002,N_16060);
nand U16380 (N_16380,N_16181,N_16033);
nor U16381 (N_16381,N_16115,N_16082);
or U16382 (N_16382,N_16079,N_16140);
nand U16383 (N_16383,N_16050,N_16166);
nor U16384 (N_16384,N_16043,N_16068);
and U16385 (N_16385,N_16107,N_16173);
nand U16386 (N_16386,N_16126,N_16145);
nand U16387 (N_16387,N_16066,N_16168);
and U16388 (N_16388,N_16139,N_16046);
or U16389 (N_16389,N_16114,N_16048);
nor U16390 (N_16390,N_16097,N_16007);
and U16391 (N_16391,N_16150,N_16121);
and U16392 (N_16392,N_16147,N_16104);
xnor U16393 (N_16393,N_16007,N_16080);
nand U16394 (N_16394,N_16026,N_16125);
xnor U16395 (N_16395,N_16089,N_16101);
nand U16396 (N_16396,N_16008,N_16014);
xor U16397 (N_16397,N_16024,N_16118);
nor U16398 (N_16398,N_16044,N_16196);
nand U16399 (N_16399,N_16164,N_16127);
and U16400 (N_16400,N_16354,N_16349);
and U16401 (N_16401,N_16376,N_16267);
nand U16402 (N_16402,N_16230,N_16283);
and U16403 (N_16403,N_16325,N_16280);
nor U16404 (N_16404,N_16229,N_16355);
xnor U16405 (N_16405,N_16323,N_16331);
or U16406 (N_16406,N_16210,N_16217);
or U16407 (N_16407,N_16255,N_16377);
and U16408 (N_16408,N_16251,N_16307);
nor U16409 (N_16409,N_16254,N_16305);
and U16410 (N_16410,N_16277,N_16272);
nor U16411 (N_16411,N_16322,N_16279);
nor U16412 (N_16412,N_16339,N_16208);
or U16413 (N_16413,N_16232,N_16231);
and U16414 (N_16414,N_16356,N_16304);
and U16415 (N_16415,N_16236,N_16319);
nor U16416 (N_16416,N_16380,N_16292);
nand U16417 (N_16417,N_16332,N_16249);
or U16418 (N_16418,N_16389,N_16333);
and U16419 (N_16419,N_16214,N_16371);
or U16420 (N_16420,N_16264,N_16365);
nand U16421 (N_16421,N_16291,N_16224);
or U16422 (N_16422,N_16341,N_16212);
nand U16423 (N_16423,N_16266,N_16282);
xor U16424 (N_16424,N_16330,N_16218);
or U16425 (N_16425,N_16386,N_16387);
nand U16426 (N_16426,N_16335,N_16316);
nand U16427 (N_16427,N_16343,N_16309);
or U16428 (N_16428,N_16327,N_16385);
xor U16429 (N_16429,N_16259,N_16394);
nand U16430 (N_16430,N_16326,N_16329);
and U16431 (N_16431,N_16225,N_16248);
and U16432 (N_16432,N_16368,N_16374);
nand U16433 (N_16433,N_16346,N_16347);
nor U16434 (N_16434,N_16258,N_16297);
nand U16435 (N_16435,N_16233,N_16301);
xnor U16436 (N_16436,N_16362,N_16300);
nor U16437 (N_16437,N_16364,N_16234);
nor U16438 (N_16438,N_16281,N_16393);
nand U16439 (N_16439,N_16201,N_16289);
nor U16440 (N_16440,N_16246,N_16392);
and U16441 (N_16441,N_16285,N_16382);
xor U16442 (N_16442,N_16293,N_16314);
and U16443 (N_16443,N_16378,N_16398);
nor U16444 (N_16444,N_16381,N_16286);
nand U16445 (N_16445,N_16317,N_16227);
or U16446 (N_16446,N_16342,N_16265);
xnor U16447 (N_16447,N_16357,N_16296);
nor U16448 (N_16448,N_16253,N_16351);
or U16449 (N_16449,N_16226,N_16216);
nand U16450 (N_16450,N_16337,N_16245);
or U16451 (N_16451,N_16324,N_16370);
nor U16452 (N_16452,N_16363,N_16271);
xnor U16453 (N_16453,N_16353,N_16284);
and U16454 (N_16454,N_16369,N_16261);
and U16455 (N_16455,N_16312,N_16373);
or U16456 (N_16456,N_16313,N_16310);
nor U16457 (N_16457,N_16311,N_16207);
or U16458 (N_16458,N_16256,N_16344);
xor U16459 (N_16459,N_16205,N_16270);
nor U16460 (N_16460,N_16395,N_16384);
and U16461 (N_16461,N_16320,N_16388);
and U16462 (N_16462,N_16383,N_16367);
and U16463 (N_16463,N_16278,N_16321);
nand U16464 (N_16464,N_16390,N_16243);
or U16465 (N_16465,N_16223,N_16338);
nand U16466 (N_16466,N_16274,N_16200);
and U16467 (N_16467,N_16379,N_16399);
nor U16468 (N_16468,N_16220,N_16275);
and U16469 (N_16469,N_16352,N_16299);
and U16470 (N_16470,N_16302,N_16268);
and U16471 (N_16471,N_16202,N_16209);
and U16472 (N_16472,N_16361,N_16318);
nor U16473 (N_16473,N_16391,N_16219);
xnor U16474 (N_16474,N_16239,N_16345);
nand U16475 (N_16475,N_16396,N_16228);
or U16476 (N_16476,N_16288,N_16269);
and U16477 (N_16477,N_16241,N_16360);
xnor U16478 (N_16478,N_16372,N_16303);
nand U16479 (N_16479,N_16375,N_16237);
xnor U16480 (N_16480,N_16244,N_16306);
or U16481 (N_16481,N_16235,N_16262);
and U16482 (N_16482,N_16221,N_16203);
nor U16483 (N_16483,N_16250,N_16328);
and U16484 (N_16484,N_16257,N_16215);
or U16485 (N_16485,N_16276,N_16242);
nor U16486 (N_16486,N_16295,N_16213);
nand U16487 (N_16487,N_16260,N_16348);
xor U16488 (N_16488,N_16206,N_16366);
xnor U16489 (N_16489,N_16290,N_16240);
nor U16490 (N_16490,N_16287,N_16359);
nand U16491 (N_16491,N_16350,N_16222);
and U16492 (N_16492,N_16294,N_16238);
or U16493 (N_16493,N_16273,N_16211);
or U16494 (N_16494,N_16308,N_16315);
nor U16495 (N_16495,N_16358,N_16334);
xnor U16496 (N_16496,N_16247,N_16340);
nand U16497 (N_16497,N_16336,N_16397);
and U16498 (N_16498,N_16252,N_16263);
and U16499 (N_16499,N_16298,N_16204);
nor U16500 (N_16500,N_16286,N_16301);
or U16501 (N_16501,N_16345,N_16251);
nor U16502 (N_16502,N_16384,N_16315);
nor U16503 (N_16503,N_16383,N_16205);
nor U16504 (N_16504,N_16347,N_16390);
xnor U16505 (N_16505,N_16272,N_16243);
or U16506 (N_16506,N_16277,N_16204);
and U16507 (N_16507,N_16275,N_16225);
xor U16508 (N_16508,N_16302,N_16378);
nor U16509 (N_16509,N_16206,N_16219);
nor U16510 (N_16510,N_16254,N_16275);
xnor U16511 (N_16511,N_16297,N_16265);
and U16512 (N_16512,N_16389,N_16282);
xor U16513 (N_16513,N_16200,N_16320);
nand U16514 (N_16514,N_16239,N_16397);
xor U16515 (N_16515,N_16324,N_16383);
and U16516 (N_16516,N_16366,N_16227);
xnor U16517 (N_16517,N_16225,N_16357);
and U16518 (N_16518,N_16241,N_16369);
or U16519 (N_16519,N_16236,N_16291);
and U16520 (N_16520,N_16373,N_16342);
nor U16521 (N_16521,N_16276,N_16323);
nor U16522 (N_16522,N_16363,N_16387);
xor U16523 (N_16523,N_16332,N_16251);
xnor U16524 (N_16524,N_16342,N_16243);
nor U16525 (N_16525,N_16326,N_16207);
nor U16526 (N_16526,N_16203,N_16340);
or U16527 (N_16527,N_16399,N_16314);
xnor U16528 (N_16528,N_16200,N_16201);
nor U16529 (N_16529,N_16382,N_16200);
nor U16530 (N_16530,N_16322,N_16333);
or U16531 (N_16531,N_16356,N_16239);
or U16532 (N_16532,N_16340,N_16284);
nand U16533 (N_16533,N_16243,N_16227);
or U16534 (N_16534,N_16260,N_16216);
xor U16535 (N_16535,N_16251,N_16258);
xnor U16536 (N_16536,N_16250,N_16276);
xor U16537 (N_16537,N_16327,N_16238);
nor U16538 (N_16538,N_16221,N_16303);
or U16539 (N_16539,N_16227,N_16228);
nand U16540 (N_16540,N_16268,N_16275);
nand U16541 (N_16541,N_16277,N_16314);
nand U16542 (N_16542,N_16320,N_16326);
and U16543 (N_16543,N_16205,N_16374);
xor U16544 (N_16544,N_16248,N_16373);
and U16545 (N_16545,N_16252,N_16247);
or U16546 (N_16546,N_16225,N_16378);
nand U16547 (N_16547,N_16357,N_16270);
xnor U16548 (N_16548,N_16279,N_16345);
nor U16549 (N_16549,N_16295,N_16339);
and U16550 (N_16550,N_16238,N_16380);
and U16551 (N_16551,N_16384,N_16218);
or U16552 (N_16552,N_16333,N_16392);
and U16553 (N_16553,N_16314,N_16214);
or U16554 (N_16554,N_16299,N_16263);
xnor U16555 (N_16555,N_16286,N_16316);
xnor U16556 (N_16556,N_16246,N_16330);
nand U16557 (N_16557,N_16385,N_16391);
and U16558 (N_16558,N_16243,N_16386);
and U16559 (N_16559,N_16269,N_16245);
and U16560 (N_16560,N_16293,N_16290);
xor U16561 (N_16561,N_16394,N_16398);
and U16562 (N_16562,N_16388,N_16299);
or U16563 (N_16563,N_16210,N_16342);
nand U16564 (N_16564,N_16384,N_16262);
nand U16565 (N_16565,N_16350,N_16223);
xor U16566 (N_16566,N_16373,N_16365);
or U16567 (N_16567,N_16204,N_16369);
xor U16568 (N_16568,N_16271,N_16281);
and U16569 (N_16569,N_16390,N_16380);
nor U16570 (N_16570,N_16391,N_16399);
or U16571 (N_16571,N_16229,N_16224);
nor U16572 (N_16572,N_16251,N_16394);
and U16573 (N_16573,N_16295,N_16227);
nand U16574 (N_16574,N_16388,N_16214);
and U16575 (N_16575,N_16342,N_16242);
and U16576 (N_16576,N_16224,N_16227);
nor U16577 (N_16577,N_16393,N_16337);
nor U16578 (N_16578,N_16344,N_16335);
nor U16579 (N_16579,N_16309,N_16353);
and U16580 (N_16580,N_16306,N_16220);
and U16581 (N_16581,N_16368,N_16335);
xnor U16582 (N_16582,N_16243,N_16297);
or U16583 (N_16583,N_16215,N_16306);
nor U16584 (N_16584,N_16268,N_16221);
or U16585 (N_16585,N_16392,N_16307);
nor U16586 (N_16586,N_16247,N_16342);
nor U16587 (N_16587,N_16200,N_16258);
nor U16588 (N_16588,N_16325,N_16214);
xor U16589 (N_16589,N_16260,N_16322);
nand U16590 (N_16590,N_16298,N_16361);
or U16591 (N_16591,N_16213,N_16293);
or U16592 (N_16592,N_16299,N_16360);
nor U16593 (N_16593,N_16346,N_16334);
xnor U16594 (N_16594,N_16341,N_16359);
nor U16595 (N_16595,N_16224,N_16218);
xnor U16596 (N_16596,N_16323,N_16356);
nor U16597 (N_16597,N_16305,N_16286);
and U16598 (N_16598,N_16242,N_16258);
xor U16599 (N_16599,N_16251,N_16370);
nand U16600 (N_16600,N_16414,N_16487);
nand U16601 (N_16601,N_16485,N_16444);
and U16602 (N_16602,N_16461,N_16580);
xor U16603 (N_16603,N_16413,N_16501);
xor U16604 (N_16604,N_16525,N_16590);
and U16605 (N_16605,N_16405,N_16498);
nor U16606 (N_16606,N_16472,N_16446);
nor U16607 (N_16607,N_16576,N_16522);
nand U16608 (N_16608,N_16436,N_16479);
nand U16609 (N_16609,N_16513,N_16482);
nor U16610 (N_16610,N_16528,N_16567);
and U16611 (N_16611,N_16551,N_16497);
and U16612 (N_16612,N_16570,N_16494);
or U16613 (N_16613,N_16425,N_16592);
nor U16614 (N_16614,N_16424,N_16583);
nor U16615 (N_16615,N_16532,N_16599);
or U16616 (N_16616,N_16421,N_16574);
nor U16617 (N_16617,N_16471,N_16523);
or U16618 (N_16618,N_16554,N_16489);
or U16619 (N_16619,N_16556,N_16437);
and U16620 (N_16620,N_16406,N_16573);
xor U16621 (N_16621,N_16582,N_16459);
nand U16622 (N_16622,N_16597,N_16533);
and U16623 (N_16623,N_16475,N_16465);
nor U16624 (N_16624,N_16428,N_16577);
nor U16625 (N_16625,N_16499,N_16466);
or U16626 (N_16626,N_16433,N_16504);
and U16627 (N_16627,N_16568,N_16490);
nor U16628 (N_16628,N_16547,N_16470);
or U16629 (N_16629,N_16564,N_16429);
or U16630 (N_16630,N_16520,N_16559);
nor U16631 (N_16631,N_16516,N_16594);
nand U16632 (N_16632,N_16541,N_16578);
and U16633 (N_16633,N_16557,N_16512);
nor U16634 (N_16634,N_16515,N_16514);
and U16635 (N_16635,N_16527,N_16431);
xor U16636 (N_16636,N_16500,N_16550);
nand U16637 (N_16637,N_16565,N_16535);
xor U16638 (N_16638,N_16521,N_16450);
nor U16639 (N_16639,N_16588,N_16548);
or U16640 (N_16640,N_16427,N_16447);
nor U16641 (N_16641,N_16455,N_16418);
and U16642 (N_16642,N_16566,N_16561);
nand U16643 (N_16643,N_16430,N_16488);
or U16644 (N_16644,N_16453,N_16586);
and U16645 (N_16645,N_16549,N_16503);
and U16646 (N_16646,N_16416,N_16439);
and U16647 (N_16647,N_16589,N_16519);
xor U16648 (N_16648,N_16442,N_16462);
xor U16649 (N_16649,N_16478,N_16420);
xnor U16650 (N_16650,N_16432,N_16440);
xnor U16651 (N_16651,N_16451,N_16545);
or U16652 (N_16652,N_16401,N_16587);
nor U16653 (N_16653,N_16441,N_16408);
nand U16654 (N_16654,N_16474,N_16595);
xnor U16655 (N_16655,N_16508,N_16419);
or U16656 (N_16656,N_16569,N_16558);
or U16657 (N_16657,N_16581,N_16445);
or U16658 (N_16658,N_16552,N_16495);
or U16659 (N_16659,N_16435,N_16524);
nand U16660 (N_16660,N_16518,N_16491);
nor U16661 (N_16661,N_16531,N_16449);
or U16662 (N_16662,N_16536,N_16448);
or U16663 (N_16663,N_16506,N_16526);
nand U16664 (N_16664,N_16477,N_16510);
or U16665 (N_16665,N_16596,N_16534);
xor U16666 (N_16666,N_16409,N_16404);
nand U16667 (N_16667,N_16509,N_16412);
and U16668 (N_16668,N_16537,N_16400);
xnor U16669 (N_16669,N_16434,N_16460);
nor U16670 (N_16670,N_16492,N_16572);
nor U16671 (N_16671,N_16458,N_16483);
xor U16672 (N_16672,N_16542,N_16563);
nand U16673 (N_16673,N_16407,N_16463);
nand U16674 (N_16674,N_16598,N_16546);
nand U16675 (N_16675,N_16452,N_16467);
nand U16676 (N_16676,N_16454,N_16538);
and U16677 (N_16677,N_16496,N_16464);
or U16678 (N_16678,N_16553,N_16502);
or U16679 (N_16679,N_16505,N_16543);
nor U16680 (N_16680,N_16585,N_16457);
nand U16681 (N_16681,N_16529,N_16539);
nor U16682 (N_16682,N_16402,N_16484);
nor U16683 (N_16683,N_16540,N_16417);
xor U16684 (N_16684,N_16481,N_16426);
nor U16685 (N_16685,N_16530,N_16456);
or U16686 (N_16686,N_16410,N_16443);
nor U16687 (N_16687,N_16411,N_16544);
nand U16688 (N_16688,N_16438,N_16468);
or U16689 (N_16689,N_16555,N_16480);
or U16690 (N_16690,N_16584,N_16507);
nand U16691 (N_16691,N_16423,N_16517);
or U16692 (N_16692,N_16415,N_16486);
nand U16693 (N_16693,N_16562,N_16575);
nand U16694 (N_16694,N_16511,N_16593);
nand U16695 (N_16695,N_16571,N_16493);
nor U16696 (N_16696,N_16476,N_16469);
and U16697 (N_16697,N_16422,N_16473);
nand U16698 (N_16698,N_16403,N_16579);
nor U16699 (N_16699,N_16591,N_16560);
nand U16700 (N_16700,N_16460,N_16515);
or U16701 (N_16701,N_16512,N_16513);
xnor U16702 (N_16702,N_16525,N_16447);
and U16703 (N_16703,N_16492,N_16412);
xnor U16704 (N_16704,N_16542,N_16567);
xnor U16705 (N_16705,N_16422,N_16415);
nor U16706 (N_16706,N_16562,N_16475);
xor U16707 (N_16707,N_16446,N_16540);
and U16708 (N_16708,N_16572,N_16403);
xor U16709 (N_16709,N_16483,N_16506);
nand U16710 (N_16710,N_16478,N_16528);
nor U16711 (N_16711,N_16519,N_16561);
and U16712 (N_16712,N_16449,N_16509);
and U16713 (N_16713,N_16556,N_16460);
nor U16714 (N_16714,N_16410,N_16532);
nor U16715 (N_16715,N_16537,N_16535);
nand U16716 (N_16716,N_16433,N_16424);
and U16717 (N_16717,N_16575,N_16438);
nand U16718 (N_16718,N_16466,N_16582);
nor U16719 (N_16719,N_16481,N_16525);
and U16720 (N_16720,N_16595,N_16445);
and U16721 (N_16721,N_16516,N_16472);
xor U16722 (N_16722,N_16579,N_16490);
nor U16723 (N_16723,N_16481,N_16528);
and U16724 (N_16724,N_16422,N_16596);
xnor U16725 (N_16725,N_16575,N_16598);
or U16726 (N_16726,N_16519,N_16424);
xor U16727 (N_16727,N_16517,N_16492);
or U16728 (N_16728,N_16537,N_16511);
xnor U16729 (N_16729,N_16426,N_16458);
xor U16730 (N_16730,N_16574,N_16460);
and U16731 (N_16731,N_16468,N_16527);
or U16732 (N_16732,N_16472,N_16585);
nand U16733 (N_16733,N_16534,N_16443);
and U16734 (N_16734,N_16543,N_16450);
nor U16735 (N_16735,N_16465,N_16549);
and U16736 (N_16736,N_16544,N_16514);
nor U16737 (N_16737,N_16420,N_16598);
nand U16738 (N_16738,N_16443,N_16424);
or U16739 (N_16739,N_16468,N_16577);
and U16740 (N_16740,N_16510,N_16474);
nor U16741 (N_16741,N_16560,N_16579);
xor U16742 (N_16742,N_16450,N_16556);
nor U16743 (N_16743,N_16471,N_16484);
xnor U16744 (N_16744,N_16570,N_16586);
xor U16745 (N_16745,N_16528,N_16487);
nor U16746 (N_16746,N_16455,N_16421);
and U16747 (N_16747,N_16542,N_16580);
nor U16748 (N_16748,N_16500,N_16539);
or U16749 (N_16749,N_16406,N_16485);
or U16750 (N_16750,N_16572,N_16508);
xnor U16751 (N_16751,N_16415,N_16446);
nor U16752 (N_16752,N_16485,N_16577);
or U16753 (N_16753,N_16420,N_16536);
and U16754 (N_16754,N_16548,N_16408);
and U16755 (N_16755,N_16430,N_16555);
nand U16756 (N_16756,N_16497,N_16520);
or U16757 (N_16757,N_16540,N_16574);
or U16758 (N_16758,N_16585,N_16445);
and U16759 (N_16759,N_16471,N_16568);
and U16760 (N_16760,N_16520,N_16455);
xor U16761 (N_16761,N_16476,N_16453);
nand U16762 (N_16762,N_16541,N_16447);
xnor U16763 (N_16763,N_16543,N_16539);
nor U16764 (N_16764,N_16541,N_16539);
or U16765 (N_16765,N_16484,N_16575);
nand U16766 (N_16766,N_16458,N_16448);
xnor U16767 (N_16767,N_16564,N_16474);
and U16768 (N_16768,N_16570,N_16510);
nor U16769 (N_16769,N_16503,N_16596);
nor U16770 (N_16770,N_16438,N_16526);
and U16771 (N_16771,N_16512,N_16520);
xor U16772 (N_16772,N_16518,N_16425);
xnor U16773 (N_16773,N_16472,N_16450);
and U16774 (N_16774,N_16496,N_16441);
nor U16775 (N_16775,N_16451,N_16549);
nor U16776 (N_16776,N_16459,N_16490);
or U16777 (N_16777,N_16516,N_16485);
nand U16778 (N_16778,N_16538,N_16573);
nor U16779 (N_16779,N_16444,N_16403);
or U16780 (N_16780,N_16502,N_16555);
nor U16781 (N_16781,N_16571,N_16546);
nand U16782 (N_16782,N_16548,N_16561);
nand U16783 (N_16783,N_16576,N_16541);
nand U16784 (N_16784,N_16445,N_16575);
or U16785 (N_16785,N_16403,N_16495);
and U16786 (N_16786,N_16507,N_16544);
nor U16787 (N_16787,N_16572,N_16466);
nand U16788 (N_16788,N_16569,N_16576);
and U16789 (N_16789,N_16563,N_16521);
xnor U16790 (N_16790,N_16591,N_16491);
or U16791 (N_16791,N_16508,N_16571);
nor U16792 (N_16792,N_16597,N_16549);
or U16793 (N_16793,N_16475,N_16495);
and U16794 (N_16794,N_16400,N_16475);
nor U16795 (N_16795,N_16506,N_16458);
and U16796 (N_16796,N_16581,N_16517);
xnor U16797 (N_16797,N_16401,N_16527);
nand U16798 (N_16798,N_16450,N_16498);
or U16799 (N_16799,N_16478,N_16588);
or U16800 (N_16800,N_16610,N_16659);
nand U16801 (N_16801,N_16661,N_16627);
xnor U16802 (N_16802,N_16635,N_16769);
or U16803 (N_16803,N_16788,N_16752);
nor U16804 (N_16804,N_16740,N_16742);
and U16805 (N_16805,N_16653,N_16671);
xnor U16806 (N_16806,N_16674,N_16728);
or U16807 (N_16807,N_16628,N_16605);
nand U16808 (N_16808,N_16690,N_16637);
or U16809 (N_16809,N_16639,N_16640);
xor U16810 (N_16810,N_16600,N_16729);
nor U16811 (N_16811,N_16603,N_16669);
nor U16812 (N_16812,N_16623,N_16702);
xnor U16813 (N_16813,N_16749,N_16707);
or U16814 (N_16814,N_16775,N_16730);
xnor U16815 (N_16815,N_16648,N_16761);
or U16816 (N_16816,N_16753,N_16660);
nand U16817 (N_16817,N_16708,N_16695);
and U16818 (N_16818,N_16774,N_16617);
or U16819 (N_16819,N_16703,N_16783);
xnor U16820 (N_16820,N_16691,N_16747);
nand U16821 (N_16821,N_16687,N_16667);
and U16822 (N_16822,N_16737,N_16722);
nand U16823 (N_16823,N_16762,N_16765);
xnor U16824 (N_16824,N_16607,N_16676);
xnor U16825 (N_16825,N_16625,N_16631);
nand U16826 (N_16826,N_16777,N_16698);
nor U16827 (N_16827,N_16618,N_16719);
nor U16828 (N_16828,N_16681,N_16606);
nand U16829 (N_16829,N_16644,N_16656);
or U16830 (N_16830,N_16650,N_16620);
nand U16831 (N_16831,N_16647,N_16713);
nor U16832 (N_16832,N_16732,N_16643);
nor U16833 (N_16833,N_16645,N_16649);
nor U16834 (N_16834,N_16770,N_16616);
nand U16835 (N_16835,N_16701,N_16678);
and U16836 (N_16836,N_16633,N_16683);
nand U16837 (N_16837,N_16685,N_16652);
or U16838 (N_16838,N_16725,N_16654);
or U16839 (N_16839,N_16721,N_16791);
nor U16840 (N_16840,N_16748,N_16686);
or U16841 (N_16841,N_16641,N_16798);
and U16842 (N_16842,N_16682,N_16630);
and U16843 (N_16843,N_16621,N_16709);
nand U16844 (N_16844,N_16779,N_16608);
xnor U16845 (N_16845,N_16785,N_16796);
and U16846 (N_16846,N_16771,N_16634);
nor U16847 (N_16847,N_16750,N_16781);
and U16848 (N_16848,N_16756,N_16764);
nor U16849 (N_16849,N_16733,N_16795);
and U16850 (N_16850,N_16755,N_16738);
nand U16851 (N_16851,N_16772,N_16697);
or U16852 (N_16852,N_16664,N_16699);
or U16853 (N_16853,N_16613,N_16794);
nor U16854 (N_16854,N_16763,N_16670);
or U16855 (N_16855,N_16679,N_16780);
and U16856 (N_16856,N_16773,N_16723);
or U16857 (N_16857,N_16636,N_16693);
xnor U16858 (N_16858,N_16714,N_16776);
nor U16859 (N_16859,N_16767,N_16799);
nor U16860 (N_16860,N_16716,N_16632);
and U16861 (N_16861,N_16758,N_16673);
xor U16862 (N_16862,N_16662,N_16768);
nor U16863 (N_16863,N_16668,N_16651);
nor U16864 (N_16864,N_16622,N_16629);
nand U16865 (N_16865,N_16757,N_16754);
or U16866 (N_16866,N_16744,N_16615);
and U16867 (N_16867,N_16666,N_16789);
nor U16868 (N_16868,N_16745,N_16705);
or U16869 (N_16869,N_16680,N_16684);
xor U16870 (N_16870,N_16797,N_16782);
or U16871 (N_16871,N_16766,N_16751);
and U16872 (N_16872,N_16675,N_16646);
and U16873 (N_16873,N_16715,N_16727);
or U16874 (N_16874,N_16759,N_16692);
xor U16875 (N_16875,N_16711,N_16609);
nor U16876 (N_16876,N_16663,N_16694);
nand U16877 (N_16877,N_16688,N_16619);
nand U16878 (N_16878,N_16743,N_16658);
nand U16879 (N_16879,N_16706,N_16793);
xor U16880 (N_16880,N_16624,N_16735);
and U16881 (N_16881,N_16790,N_16677);
xnor U16882 (N_16882,N_16604,N_16720);
nor U16883 (N_16883,N_16786,N_16704);
and U16884 (N_16884,N_16792,N_16778);
xor U16885 (N_16885,N_16726,N_16700);
and U16886 (N_16886,N_16657,N_16731);
nor U16887 (N_16887,N_16626,N_16710);
and U16888 (N_16888,N_16689,N_16734);
nor U16889 (N_16889,N_16601,N_16787);
nor U16890 (N_16890,N_16611,N_16712);
and U16891 (N_16891,N_16741,N_16718);
nor U16892 (N_16892,N_16655,N_16614);
or U16893 (N_16893,N_16696,N_16760);
nor U16894 (N_16894,N_16717,N_16665);
and U16895 (N_16895,N_16672,N_16739);
and U16896 (N_16896,N_16638,N_16784);
nor U16897 (N_16897,N_16736,N_16642);
xnor U16898 (N_16898,N_16724,N_16612);
and U16899 (N_16899,N_16746,N_16602);
and U16900 (N_16900,N_16601,N_16783);
nor U16901 (N_16901,N_16795,N_16605);
nor U16902 (N_16902,N_16789,N_16737);
and U16903 (N_16903,N_16748,N_16605);
nor U16904 (N_16904,N_16646,N_16679);
or U16905 (N_16905,N_16615,N_16747);
and U16906 (N_16906,N_16624,N_16626);
and U16907 (N_16907,N_16741,N_16640);
xnor U16908 (N_16908,N_16707,N_16742);
nand U16909 (N_16909,N_16770,N_16678);
or U16910 (N_16910,N_16623,N_16712);
xnor U16911 (N_16911,N_16792,N_16604);
or U16912 (N_16912,N_16675,N_16695);
nand U16913 (N_16913,N_16625,N_16735);
or U16914 (N_16914,N_16696,N_16798);
or U16915 (N_16915,N_16774,N_16754);
and U16916 (N_16916,N_16733,N_16637);
and U16917 (N_16917,N_16787,N_16773);
or U16918 (N_16918,N_16768,N_16729);
and U16919 (N_16919,N_16649,N_16653);
nor U16920 (N_16920,N_16652,N_16679);
and U16921 (N_16921,N_16656,N_16772);
nor U16922 (N_16922,N_16695,N_16698);
and U16923 (N_16923,N_16761,N_16770);
and U16924 (N_16924,N_16604,N_16782);
and U16925 (N_16925,N_16747,N_16754);
or U16926 (N_16926,N_16699,N_16638);
nor U16927 (N_16927,N_16763,N_16637);
nor U16928 (N_16928,N_16611,N_16757);
xor U16929 (N_16929,N_16774,N_16779);
xnor U16930 (N_16930,N_16759,N_16625);
or U16931 (N_16931,N_16601,N_16731);
nand U16932 (N_16932,N_16618,N_16688);
nand U16933 (N_16933,N_16625,N_16799);
nand U16934 (N_16934,N_16666,N_16693);
or U16935 (N_16935,N_16702,N_16670);
nand U16936 (N_16936,N_16614,N_16625);
or U16937 (N_16937,N_16752,N_16694);
nor U16938 (N_16938,N_16659,N_16749);
or U16939 (N_16939,N_16776,N_16726);
and U16940 (N_16940,N_16608,N_16630);
or U16941 (N_16941,N_16652,N_16737);
and U16942 (N_16942,N_16714,N_16767);
and U16943 (N_16943,N_16712,N_16741);
nand U16944 (N_16944,N_16695,N_16719);
nand U16945 (N_16945,N_16694,N_16638);
xnor U16946 (N_16946,N_16730,N_16612);
or U16947 (N_16947,N_16759,N_16638);
and U16948 (N_16948,N_16798,N_16737);
xnor U16949 (N_16949,N_16766,N_16621);
nand U16950 (N_16950,N_16612,N_16726);
or U16951 (N_16951,N_16782,N_16763);
nor U16952 (N_16952,N_16662,N_16787);
or U16953 (N_16953,N_16606,N_16751);
nand U16954 (N_16954,N_16698,N_16748);
nor U16955 (N_16955,N_16656,N_16614);
nor U16956 (N_16956,N_16633,N_16790);
and U16957 (N_16957,N_16762,N_16662);
and U16958 (N_16958,N_16758,N_16660);
and U16959 (N_16959,N_16767,N_16762);
or U16960 (N_16960,N_16694,N_16640);
and U16961 (N_16961,N_16727,N_16770);
and U16962 (N_16962,N_16709,N_16782);
and U16963 (N_16963,N_16765,N_16797);
xor U16964 (N_16964,N_16780,N_16724);
and U16965 (N_16965,N_16748,N_16741);
xor U16966 (N_16966,N_16757,N_16766);
and U16967 (N_16967,N_16663,N_16676);
xor U16968 (N_16968,N_16674,N_16773);
nor U16969 (N_16969,N_16719,N_16797);
or U16970 (N_16970,N_16639,N_16633);
nand U16971 (N_16971,N_16633,N_16708);
xor U16972 (N_16972,N_16694,N_16730);
and U16973 (N_16973,N_16656,N_16730);
and U16974 (N_16974,N_16642,N_16604);
or U16975 (N_16975,N_16721,N_16666);
or U16976 (N_16976,N_16631,N_16713);
nand U16977 (N_16977,N_16741,N_16654);
nor U16978 (N_16978,N_16625,N_16641);
xor U16979 (N_16979,N_16614,N_16759);
and U16980 (N_16980,N_16669,N_16708);
xor U16981 (N_16981,N_16742,N_16772);
and U16982 (N_16982,N_16737,N_16689);
xor U16983 (N_16983,N_16700,N_16717);
and U16984 (N_16984,N_16780,N_16789);
nor U16985 (N_16985,N_16749,N_16651);
nor U16986 (N_16986,N_16601,N_16778);
and U16987 (N_16987,N_16738,N_16730);
and U16988 (N_16988,N_16649,N_16728);
nor U16989 (N_16989,N_16705,N_16695);
or U16990 (N_16990,N_16649,N_16689);
or U16991 (N_16991,N_16769,N_16735);
and U16992 (N_16992,N_16699,N_16797);
or U16993 (N_16993,N_16667,N_16763);
nand U16994 (N_16994,N_16759,N_16699);
nor U16995 (N_16995,N_16607,N_16624);
and U16996 (N_16996,N_16734,N_16719);
or U16997 (N_16997,N_16706,N_16653);
and U16998 (N_16998,N_16665,N_16708);
nand U16999 (N_16999,N_16745,N_16777);
nor U17000 (N_17000,N_16841,N_16957);
or U17001 (N_17001,N_16831,N_16999);
nand U17002 (N_17002,N_16806,N_16908);
xor U17003 (N_17003,N_16919,N_16853);
nand U17004 (N_17004,N_16829,N_16873);
nand U17005 (N_17005,N_16929,N_16949);
nor U17006 (N_17006,N_16954,N_16973);
nand U17007 (N_17007,N_16932,N_16802);
and U17008 (N_17008,N_16903,N_16801);
nand U17009 (N_17009,N_16983,N_16901);
or U17010 (N_17010,N_16905,N_16852);
or U17011 (N_17011,N_16924,N_16984);
nor U17012 (N_17012,N_16943,N_16878);
nand U17013 (N_17013,N_16930,N_16914);
or U17014 (N_17014,N_16987,N_16972);
or U17015 (N_17015,N_16915,N_16800);
xor U17016 (N_17016,N_16911,N_16961);
or U17017 (N_17017,N_16870,N_16855);
or U17018 (N_17018,N_16836,N_16886);
or U17019 (N_17019,N_16958,N_16996);
and U17020 (N_17020,N_16995,N_16854);
or U17021 (N_17021,N_16944,N_16940);
nand U17022 (N_17022,N_16969,N_16970);
and U17023 (N_17023,N_16814,N_16893);
or U17024 (N_17024,N_16845,N_16861);
nor U17025 (N_17025,N_16840,N_16827);
xor U17026 (N_17026,N_16869,N_16980);
nor U17027 (N_17027,N_16913,N_16826);
nor U17028 (N_17028,N_16993,N_16948);
xor U17029 (N_17029,N_16860,N_16867);
nand U17030 (N_17030,N_16927,N_16894);
xor U17031 (N_17031,N_16876,N_16979);
or U17032 (N_17032,N_16823,N_16967);
nor U17033 (N_17033,N_16921,N_16912);
nor U17034 (N_17034,N_16922,N_16889);
xnor U17035 (N_17035,N_16879,N_16994);
nand U17036 (N_17036,N_16891,N_16935);
xor U17037 (N_17037,N_16892,N_16842);
and U17038 (N_17038,N_16926,N_16896);
xnor U17039 (N_17039,N_16863,N_16988);
nand U17040 (N_17040,N_16849,N_16821);
and U17041 (N_17041,N_16865,N_16884);
nand U17042 (N_17042,N_16937,N_16968);
or U17043 (N_17043,N_16824,N_16925);
and U17044 (N_17044,N_16811,N_16907);
nor U17045 (N_17045,N_16991,N_16837);
xor U17046 (N_17046,N_16898,N_16864);
or U17047 (N_17047,N_16882,N_16981);
nor U17048 (N_17048,N_16830,N_16890);
and U17049 (N_17049,N_16868,N_16885);
or U17050 (N_17050,N_16866,N_16959);
and U17051 (N_17051,N_16945,N_16874);
or U17052 (N_17052,N_16978,N_16939);
xor U17053 (N_17053,N_16818,N_16875);
nor U17054 (N_17054,N_16812,N_16900);
nor U17055 (N_17055,N_16834,N_16971);
nand U17056 (N_17056,N_16858,N_16871);
nor U17057 (N_17057,N_16833,N_16904);
and U17058 (N_17058,N_16817,N_16955);
xnor U17059 (N_17059,N_16951,N_16966);
nand U17060 (N_17060,N_16974,N_16942);
nor U17061 (N_17061,N_16928,N_16920);
or U17062 (N_17062,N_16810,N_16976);
nand U17063 (N_17063,N_16828,N_16846);
nor U17064 (N_17064,N_16963,N_16918);
nand U17065 (N_17065,N_16883,N_16964);
nor U17066 (N_17066,N_16986,N_16950);
nand U17067 (N_17067,N_16997,N_16897);
nand U17068 (N_17068,N_16805,N_16902);
nand U17069 (N_17069,N_16835,N_16888);
nand U17070 (N_17070,N_16909,N_16856);
and U17071 (N_17071,N_16803,N_16838);
xor U17072 (N_17072,N_16804,N_16936);
and U17073 (N_17073,N_16880,N_16808);
and U17074 (N_17074,N_16872,N_16887);
nor U17075 (N_17075,N_16895,N_16960);
nand U17076 (N_17076,N_16839,N_16975);
nor U17077 (N_17077,N_16815,N_16946);
or U17078 (N_17078,N_16998,N_16938);
xor U17079 (N_17079,N_16947,N_16807);
nor U17080 (N_17080,N_16899,N_16931);
or U17081 (N_17081,N_16989,N_16813);
nor U17082 (N_17082,N_16933,N_16847);
nand U17083 (N_17083,N_16844,N_16952);
and U17084 (N_17084,N_16862,N_16962);
nor U17085 (N_17085,N_16877,N_16819);
nor U17086 (N_17086,N_16916,N_16990);
and U17087 (N_17087,N_16917,N_16906);
or U17088 (N_17088,N_16857,N_16816);
nand U17089 (N_17089,N_16977,N_16992);
nor U17090 (N_17090,N_16843,N_16982);
and U17091 (N_17091,N_16934,N_16820);
and U17092 (N_17092,N_16848,N_16953);
and U17093 (N_17093,N_16859,N_16923);
and U17094 (N_17094,N_16850,N_16809);
nand U17095 (N_17095,N_16941,N_16822);
nor U17096 (N_17096,N_16825,N_16832);
and U17097 (N_17097,N_16985,N_16851);
nand U17098 (N_17098,N_16956,N_16881);
or U17099 (N_17099,N_16910,N_16965);
nand U17100 (N_17100,N_16902,N_16985);
xor U17101 (N_17101,N_16903,N_16965);
xnor U17102 (N_17102,N_16854,N_16966);
and U17103 (N_17103,N_16999,N_16868);
or U17104 (N_17104,N_16971,N_16911);
xnor U17105 (N_17105,N_16910,N_16824);
nor U17106 (N_17106,N_16870,N_16812);
nor U17107 (N_17107,N_16924,N_16845);
nor U17108 (N_17108,N_16963,N_16934);
or U17109 (N_17109,N_16977,N_16804);
nor U17110 (N_17110,N_16995,N_16841);
nand U17111 (N_17111,N_16826,N_16899);
nor U17112 (N_17112,N_16931,N_16871);
or U17113 (N_17113,N_16901,N_16834);
and U17114 (N_17114,N_16835,N_16803);
nand U17115 (N_17115,N_16910,N_16862);
nand U17116 (N_17116,N_16892,N_16913);
and U17117 (N_17117,N_16928,N_16827);
nand U17118 (N_17118,N_16930,N_16836);
and U17119 (N_17119,N_16882,N_16832);
and U17120 (N_17120,N_16969,N_16883);
or U17121 (N_17121,N_16986,N_16882);
nand U17122 (N_17122,N_16888,N_16854);
nand U17123 (N_17123,N_16925,N_16830);
or U17124 (N_17124,N_16854,N_16904);
and U17125 (N_17125,N_16874,N_16810);
xor U17126 (N_17126,N_16922,N_16865);
xor U17127 (N_17127,N_16862,N_16900);
nand U17128 (N_17128,N_16882,N_16979);
and U17129 (N_17129,N_16989,N_16974);
or U17130 (N_17130,N_16822,N_16876);
nand U17131 (N_17131,N_16815,N_16845);
nor U17132 (N_17132,N_16836,N_16961);
or U17133 (N_17133,N_16988,N_16860);
xor U17134 (N_17134,N_16882,N_16968);
xnor U17135 (N_17135,N_16917,N_16832);
or U17136 (N_17136,N_16966,N_16822);
nor U17137 (N_17137,N_16961,N_16906);
or U17138 (N_17138,N_16883,N_16959);
xor U17139 (N_17139,N_16888,N_16844);
nand U17140 (N_17140,N_16819,N_16962);
xor U17141 (N_17141,N_16906,N_16862);
nand U17142 (N_17142,N_16981,N_16812);
or U17143 (N_17143,N_16951,N_16882);
or U17144 (N_17144,N_16827,N_16955);
xor U17145 (N_17145,N_16962,N_16945);
nor U17146 (N_17146,N_16930,N_16829);
or U17147 (N_17147,N_16888,N_16996);
nand U17148 (N_17148,N_16833,N_16902);
or U17149 (N_17149,N_16948,N_16973);
nand U17150 (N_17150,N_16924,N_16983);
or U17151 (N_17151,N_16939,N_16959);
and U17152 (N_17152,N_16809,N_16973);
or U17153 (N_17153,N_16816,N_16937);
or U17154 (N_17154,N_16831,N_16841);
nand U17155 (N_17155,N_16917,N_16854);
xor U17156 (N_17156,N_16827,N_16960);
nand U17157 (N_17157,N_16959,N_16899);
nand U17158 (N_17158,N_16985,N_16888);
nor U17159 (N_17159,N_16938,N_16970);
and U17160 (N_17160,N_16918,N_16913);
or U17161 (N_17161,N_16915,N_16876);
or U17162 (N_17162,N_16982,N_16827);
nor U17163 (N_17163,N_16970,N_16874);
and U17164 (N_17164,N_16864,N_16810);
and U17165 (N_17165,N_16802,N_16827);
and U17166 (N_17166,N_16870,N_16936);
or U17167 (N_17167,N_16978,N_16877);
or U17168 (N_17168,N_16918,N_16863);
and U17169 (N_17169,N_16892,N_16914);
or U17170 (N_17170,N_16805,N_16848);
or U17171 (N_17171,N_16808,N_16846);
or U17172 (N_17172,N_16998,N_16869);
and U17173 (N_17173,N_16841,N_16999);
and U17174 (N_17174,N_16850,N_16962);
xnor U17175 (N_17175,N_16800,N_16846);
or U17176 (N_17176,N_16835,N_16809);
or U17177 (N_17177,N_16988,N_16807);
nand U17178 (N_17178,N_16962,N_16874);
xnor U17179 (N_17179,N_16885,N_16987);
nand U17180 (N_17180,N_16917,N_16834);
and U17181 (N_17181,N_16910,N_16925);
nand U17182 (N_17182,N_16840,N_16885);
nand U17183 (N_17183,N_16864,N_16988);
xor U17184 (N_17184,N_16829,N_16835);
xnor U17185 (N_17185,N_16849,N_16887);
xor U17186 (N_17186,N_16885,N_16923);
or U17187 (N_17187,N_16840,N_16923);
or U17188 (N_17188,N_16859,N_16885);
and U17189 (N_17189,N_16810,N_16968);
nor U17190 (N_17190,N_16854,N_16979);
nor U17191 (N_17191,N_16996,N_16810);
and U17192 (N_17192,N_16924,N_16936);
or U17193 (N_17193,N_16827,N_16823);
and U17194 (N_17194,N_16992,N_16911);
xnor U17195 (N_17195,N_16909,N_16967);
and U17196 (N_17196,N_16951,N_16833);
xor U17197 (N_17197,N_16951,N_16842);
and U17198 (N_17198,N_16889,N_16898);
xor U17199 (N_17199,N_16864,N_16859);
and U17200 (N_17200,N_17163,N_17113);
or U17201 (N_17201,N_17042,N_17178);
and U17202 (N_17202,N_17162,N_17085);
nand U17203 (N_17203,N_17084,N_17112);
nand U17204 (N_17204,N_17010,N_17058);
or U17205 (N_17205,N_17027,N_17095);
or U17206 (N_17206,N_17199,N_17141);
or U17207 (N_17207,N_17136,N_17089);
xor U17208 (N_17208,N_17183,N_17166);
and U17209 (N_17209,N_17186,N_17195);
nand U17210 (N_17210,N_17043,N_17131);
nor U17211 (N_17211,N_17132,N_17160);
nor U17212 (N_17212,N_17031,N_17137);
nand U17213 (N_17213,N_17127,N_17119);
xnor U17214 (N_17214,N_17152,N_17125);
and U17215 (N_17215,N_17017,N_17111);
nand U17216 (N_17216,N_17075,N_17139);
or U17217 (N_17217,N_17123,N_17090);
nor U17218 (N_17218,N_17102,N_17138);
nand U17219 (N_17219,N_17192,N_17171);
nand U17220 (N_17220,N_17002,N_17001);
and U17221 (N_17221,N_17045,N_17145);
xor U17222 (N_17222,N_17114,N_17173);
and U17223 (N_17223,N_17037,N_17154);
nand U17224 (N_17224,N_17153,N_17074);
nor U17225 (N_17225,N_17087,N_17105);
and U17226 (N_17226,N_17038,N_17046);
nand U17227 (N_17227,N_17184,N_17118);
and U17228 (N_17228,N_17078,N_17073);
nor U17229 (N_17229,N_17011,N_17181);
xnor U17230 (N_17230,N_17099,N_17096);
xnor U17231 (N_17231,N_17142,N_17097);
nor U17232 (N_17232,N_17187,N_17028);
or U17233 (N_17233,N_17040,N_17080);
nor U17234 (N_17234,N_17059,N_17103);
nor U17235 (N_17235,N_17077,N_17168);
xnor U17236 (N_17236,N_17193,N_17176);
nand U17237 (N_17237,N_17051,N_17021);
and U17238 (N_17238,N_17106,N_17120);
and U17239 (N_17239,N_17128,N_17052);
nand U17240 (N_17240,N_17057,N_17025);
nor U17241 (N_17241,N_17047,N_17065);
or U17242 (N_17242,N_17140,N_17034);
xor U17243 (N_17243,N_17061,N_17134);
nand U17244 (N_17244,N_17069,N_17158);
or U17245 (N_17245,N_17117,N_17100);
nand U17246 (N_17246,N_17003,N_17126);
and U17247 (N_17247,N_17086,N_17108);
or U17248 (N_17248,N_17161,N_17135);
nor U17249 (N_17249,N_17129,N_17014);
xor U17250 (N_17250,N_17004,N_17169);
nor U17251 (N_17251,N_17091,N_17109);
xor U17252 (N_17252,N_17094,N_17185);
or U17253 (N_17253,N_17013,N_17008);
xor U17254 (N_17254,N_17067,N_17194);
xor U17255 (N_17255,N_17143,N_17180);
xor U17256 (N_17256,N_17019,N_17115);
or U17257 (N_17257,N_17079,N_17036);
xor U17258 (N_17258,N_17083,N_17093);
or U17259 (N_17259,N_17060,N_17012);
xnor U17260 (N_17260,N_17006,N_17054);
or U17261 (N_17261,N_17015,N_17072);
or U17262 (N_17262,N_17023,N_17053);
nand U17263 (N_17263,N_17104,N_17035);
and U17264 (N_17264,N_17039,N_17020);
nor U17265 (N_17265,N_17157,N_17167);
xor U17266 (N_17266,N_17101,N_17197);
xnor U17267 (N_17267,N_17107,N_17070);
nor U17268 (N_17268,N_17055,N_17190);
nor U17269 (N_17269,N_17066,N_17018);
nor U17270 (N_17270,N_17076,N_17068);
and U17271 (N_17271,N_17170,N_17164);
nand U17272 (N_17272,N_17177,N_17148);
and U17273 (N_17273,N_17005,N_17081);
or U17274 (N_17274,N_17071,N_17029);
xor U17275 (N_17275,N_17174,N_17048);
and U17276 (N_17276,N_17150,N_17124);
nor U17277 (N_17277,N_17026,N_17044);
and U17278 (N_17278,N_17041,N_17182);
and U17279 (N_17279,N_17024,N_17189);
and U17280 (N_17280,N_17121,N_17030);
nor U17281 (N_17281,N_17151,N_17092);
nand U17282 (N_17282,N_17196,N_17188);
nand U17283 (N_17283,N_17191,N_17049);
or U17284 (N_17284,N_17050,N_17064);
xnor U17285 (N_17285,N_17149,N_17172);
or U17286 (N_17286,N_17063,N_17144);
and U17287 (N_17287,N_17198,N_17116);
or U17288 (N_17288,N_17098,N_17155);
nand U17289 (N_17289,N_17156,N_17130);
xor U17290 (N_17290,N_17062,N_17175);
nor U17291 (N_17291,N_17122,N_17146);
xor U17292 (N_17292,N_17009,N_17033);
or U17293 (N_17293,N_17088,N_17147);
or U17294 (N_17294,N_17110,N_17159);
nand U17295 (N_17295,N_17165,N_17082);
and U17296 (N_17296,N_17000,N_17179);
xnor U17297 (N_17297,N_17133,N_17032);
nand U17298 (N_17298,N_17016,N_17007);
and U17299 (N_17299,N_17056,N_17022);
or U17300 (N_17300,N_17046,N_17083);
xor U17301 (N_17301,N_17002,N_17078);
nor U17302 (N_17302,N_17162,N_17196);
and U17303 (N_17303,N_17191,N_17175);
or U17304 (N_17304,N_17182,N_17072);
and U17305 (N_17305,N_17066,N_17135);
and U17306 (N_17306,N_17028,N_17020);
nor U17307 (N_17307,N_17122,N_17195);
or U17308 (N_17308,N_17081,N_17006);
or U17309 (N_17309,N_17085,N_17080);
xnor U17310 (N_17310,N_17000,N_17128);
or U17311 (N_17311,N_17061,N_17001);
or U17312 (N_17312,N_17005,N_17042);
and U17313 (N_17313,N_17128,N_17044);
xor U17314 (N_17314,N_17186,N_17180);
and U17315 (N_17315,N_17057,N_17054);
or U17316 (N_17316,N_17006,N_17077);
nand U17317 (N_17317,N_17085,N_17079);
nor U17318 (N_17318,N_17136,N_17023);
or U17319 (N_17319,N_17071,N_17165);
nor U17320 (N_17320,N_17023,N_17110);
xor U17321 (N_17321,N_17031,N_17003);
xor U17322 (N_17322,N_17194,N_17037);
or U17323 (N_17323,N_17104,N_17057);
nor U17324 (N_17324,N_17053,N_17196);
nor U17325 (N_17325,N_17043,N_17081);
xnor U17326 (N_17326,N_17029,N_17135);
or U17327 (N_17327,N_17000,N_17101);
xnor U17328 (N_17328,N_17067,N_17172);
nand U17329 (N_17329,N_17144,N_17158);
xnor U17330 (N_17330,N_17020,N_17057);
xnor U17331 (N_17331,N_17135,N_17071);
or U17332 (N_17332,N_17187,N_17144);
xnor U17333 (N_17333,N_17056,N_17045);
xnor U17334 (N_17334,N_17150,N_17005);
nand U17335 (N_17335,N_17061,N_17139);
nor U17336 (N_17336,N_17000,N_17196);
and U17337 (N_17337,N_17109,N_17132);
nand U17338 (N_17338,N_17176,N_17140);
and U17339 (N_17339,N_17143,N_17127);
nor U17340 (N_17340,N_17128,N_17039);
and U17341 (N_17341,N_17175,N_17010);
and U17342 (N_17342,N_17163,N_17095);
or U17343 (N_17343,N_17179,N_17082);
nand U17344 (N_17344,N_17130,N_17190);
or U17345 (N_17345,N_17018,N_17137);
nand U17346 (N_17346,N_17154,N_17160);
or U17347 (N_17347,N_17149,N_17085);
nor U17348 (N_17348,N_17134,N_17000);
nand U17349 (N_17349,N_17128,N_17048);
nor U17350 (N_17350,N_17017,N_17175);
nor U17351 (N_17351,N_17000,N_17178);
or U17352 (N_17352,N_17019,N_17098);
nand U17353 (N_17353,N_17091,N_17077);
xnor U17354 (N_17354,N_17195,N_17182);
nor U17355 (N_17355,N_17017,N_17145);
xor U17356 (N_17356,N_17100,N_17167);
nand U17357 (N_17357,N_17083,N_17174);
xor U17358 (N_17358,N_17185,N_17036);
or U17359 (N_17359,N_17034,N_17049);
or U17360 (N_17360,N_17162,N_17069);
nand U17361 (N_17361,N_17199,N_17019);
nand U17362 (N_17362,N_17150,N_17138);
nor U17363 (N_17363,N_17127,N_17008);
nand U17364 (N_17364,N_17025,N_17022);
or U17365 (N_17365,N_17135,N_17010);
nor U17366 (N_17366,N_17112,N_17013);
xor U17367 (N_17367,N_17079,N_17119);
nand U17368 (N_17368,N_17176,N_17117);
or U17369 (N_17369,N_17186,N_17171);
nor U17370 (N_17370,N_17087,N_17164);
or U17371 (N_17371,N_17193,N_17157);
or U17372 (N_17372,N_17082,N_17005);
nand U17373 (N_17373,N_17075,N_17129);
xnor U17374 (N_17374,N_17016,N_17071);
xnor U17375 (N_17375,N_17178,N_17080);
nand U17376 (N_17376,N_17133,N_17007);
and U17377 (N_17377,N_17021,N_17150);
nor U17378 (N_17378,N_17064,N_17163);
or U17379 (N_17379,N_17116,N_17167);
or U17380 (N_17380,N_17085,N_17150);
nand U17381 (N_17381,N_17074,N_17011);
xor U17382 (N_17382,N_17082,N_17037);
nor U17383 (N_17383,N_17011,N_17174);
nor U17384 (N_17384,N_17166,N_17076);
and U17385 (N_17385,N_17129,N_17085);
nor U17386 (N_17386,N_17102,N_17183);
nand U17387 (N_17387,N_17101,N_17071);
and U17388 (N_17388,N_17056,N_17069);
and U17389 (N_17389,N_17121,N_17199);
nand U17390 (N_17390,N_17083,N_17065);
nand U17391 (N_17391,N_17047,N_17129);
nor U17392 (N_17392,N_17105,N_17113);
nor U17393 (N_17393,N_17018,N_17010);
xnor U17394 (N_17394,N_17068,N_17074);
nor U17395 (N_17395,N_17183,N_17055);
nor U17396 (N_17396,N_17140,N_17068);
or U17397 (N_17397,N_17175,N_17182);
xor U17398 (N_17398,N_17050,N_17157);
or U17399 (N_17399,N_17162,N_17019);
xnor U17400 (N_17400,N_17343,N_17296);
nand U17401 (N_17401,N_17306,N_17240);
xor U17402 (N_17402,N_17214,N_17337);
nand U17403 (N_17403,N_17212,N_17218);
nand U17404 (N_17404,N_17208,N_17287);
nor U17405 (N_17405,N_17352,N_17265);
and U17406 (N_17406,N_17272,N_17248);
or U17407 (N_17407,N_17327,N_17295);
nor U17408 (N_17408,N_17275,N_17252);
nand U17409 (N_17409,N_17390,N_17294);
nor U17410 (N_17410,N_17396,N_17378);
nand U17411 (N_17411,N_17215,N_17235);
or U17412 (N_17412,N_17326,N_17388);
xor U17413 (N_17413,N_17342,N_17331);
xor U17414 (N_17414,N_17260,N_17340);
nand U17415 (N_17415,N_17268,N_17317);
and U17416 (N_17416,N_17348,N_17321);
and U17417 (N_17417,N_17316,N_17264);
nand U17418 (N_17418,N_17257,N_17332);
nand U17419 (N_17419,N_17293,N_17262);
or U17420 (N_17420,N_17357,N_17242);
nor U17421 (N_17421,N_17395,N_17291);
or U17422 (N_17422,N_17339,N_17376);
nor U17423 (N_17423,N_17303,N_17251);
and U17424 (N_17424,N_17325,N_17322);
xor U17425 (N_17425,N_17206,N_17282);
and U17426 (N_17426,N_17372,N_17399);
and U17427 (N_17427,N_17209,N_17245);
nand U17428 (N_17428,N_17261,N_17213);
nor U17429 (N_17429,N_17375,N_17389);
and U17430 (N_17430,N_17356,N_17284);
and U17431 (N_17431,N_17380,N_17216);
and U17432 (N_17432,N_17315,N_17397);
xnor U17433 (N_17433,N_17207,N_17387);
or U17434 (N_17434,N_17367,N_17308);
xnor U17435 (N_17435,N_17362,N_17392);
nor U17436 (N_17436,N_17220,N_17297);
nand U17437 (N_17437,N_17274,N_17283);
or U17438 (N_17438,N_17219,N_17353);
nor U17439 (N_17439,N_17255,N_17358);
nor U17440 (N_17440,N_17278,N_17314);
xor U17441 (N_17441,N_17319,N_17254);
and U17442 (N_17442,N_17224,N_17301);
or U17443 (N_17443,N_17323,N_17328);
or U17444 (N_17444,N_17365,N_17217);
nor U17445 (N_17445,N_17205,N_17344);
and U17446 (N_17446,N_17288,N_17229);
xor U17447 (N_17447,N_17371,N_17318);
xnor U17448 (N_17448,N_17253,N_17230);
and U17449 (N_17449,N_17335,N_17292);
and U17450 (N_17450,N_17241,N_17305);
nand U17451 (N_17451,N_17223,N_17243);
or U17452 (N_17452,N_17202,N_17310);
xor U17453 (N_17453,N_17354,N_17382);
nand U17454 (N_17454,N_17329,N_17290);
nor U17455 (N_17455,N_17263,N_17232);
nand U17456 (N_17456,N_17204,N_17200);
or U17457 (N_17457,N_17302,N_17393);
xor U17458 (N_17458,N_17313,N_17211);
xor U17459 (N_17459,N_17298,N_17304);
xor U17460 (N_17460,N_17234,N_17269);
or U17461 (N_17461,N_17355,N_17227);
nand U17462 (N_17462,N_17320,N_17270);
nand U17463 (N_17463,N_17256,N_17300);
nor U17464 (N_17464,N_17345,N_17259);
nor U17465 (N_17465,N_17276,N_17277);
or U17466 (N_17466,N_17346,N_17394);
nor U17467 (N_17467,N_17379,N_17370);
nor U17468 (N_17468,N_17384,N_17368);
and U17469 (N_17469,N_17398,N_17312);
nand U17470 (N_17470,N_17360,N_17299);
nand U17471 (N_17471,N_17369,N_17289);
nor U17472 (N_17472,N_17273,N_17203);
and U17473 (N_17473,N_17201,N_17381);
xnor U17474 (N_17474,N_17373,N_17333);
and U17475 (N_17475,N_17236,N_17351);
nand U17476 (N_17476,N_17350,N_17285);
nor U17477 (N_17477,N_17233,N_17341);
nand U17478 (N_17478,N_17249,N_17246);
and U17479 (N_17479,N_17386,N_17377);
nand U17480 (N_17480,N_17334,N_17391);
or U17481 (N_17481,N_17324,N_17266);
xnor U17482 (N_17482,N_17349,N_17239);
xor U17483 (N_17483,N_17311,N_17286);
nor U17484 (N_17484,N_17231,N_17363);
nand U17485 (N_17485,N_17244,N_17336);
or U17486 (N_17486,N_17226,N_17364);
and U17487 (N_17487,N_17330,N_17338);
nand U17488 (N_17488,N_17366,N_17238);
or U17489 (N_17489,N_17361,N_17271);
nor U17490 (N_17490,N_17307,N_17210);
nor U17491 (N_17491,N_17250,N_17281);
nor U17492 (N_17492,N_17385,N_17247);
and U17493 (N_17493,N_17222,N_17258);
nor U17494 (N_17494,N_17347,N_17383);
nor U17495 (N_17495,N_17374,N_17225);
or U17496 (N_17496,N_17267,N_17309);
xnor U17497 (N_17497,N_17280,N_17359);
xnor U17498 (N_17498,N_17237,N_17228);
or U17499 (N_17499,N_17279,N_17221);
and U17500 (N_17500,N_17243,N_17212);
nor U17501 (N_17501,N_17346,N_17290);
and U17502 (N_17502,N_17326,N_17324);
and U17503 (N_17503,N_17358,N_17310);
nor U17504 (N_17504,N_17368,N_17314);
nor U17505 (N_17505,N_17300,N_17387);
or U17506 (N_17506,N_17287,N_17309);
or U17507 (N_17507,N_17337,N_17209);
xor U17508 (N_17508,N_17259,N_17374);
nand U17509 (N_17509,N_17365,N_17385);
and U17510 (N_17510,N_17392,N_17384);
nor U17511 (N_17511,N_17389,N_17209);
xor U17512 (N_17512,N_17360,N_17242);
nand U17513 (N_17513,N_17390,N_17279);
and U17514 (N_17514,N_17208,N_17379);
or U17515 (N_17515,N_17398,N_17385);
or U17516 (N_17516,N_17226,N_17248);
nand U17517 (N_17517,N_17334,N_17204);
nor U17518 (N_17518,N_17240,N_17269);
or U17519 (N_17519,N_17302,N_17215);
nor U17520 (N_17520,N_17219,N_17222);
or U17521 (N_17521,N_17263,N_17227);
nand U17522 (N_17522,N_17295,N_17368);
nor U17523 (N_17523,N_17297,N_17240);
and U17524 (N_17524,N_17385,N_17283);
nor U17525 (N_17525,N_17257,N_17269);
xnor U17526 (N_17526,N_17336,N_17329);
nor U17527 (N_17527,N_17209,N_17376);
or U17528 (N_17528,N_17339,N_17392);
or U17529 (N_17529,N_17395,N_17269);
and U17530 (N_17530,N_17304,N_17327);
xor U17531 (N_17531,N_17276,N_17361);
and U17532 (N_17532,N_17382,N_17286);
or U17533 (N_17533,N_17342,N_17350);
and U17534 (N_17534,N_17281,N_17334);
xor U17535 (N_17535,N_17256,N_17252);
xor U17536 (N_17536,N_17207,N_17209);
xnor U17537 (N_17537,N_17328,N_17204);
nor U17538 (N_17538,N_17212,N_17309);
nor U17539 (N_17539,N_17332,N_17395);
nand U17540 (N_17540,N_17385,N_17246);
nor U17541 (N_17541,N_17385,N_17294);
nand U17542 (N_17542,N_17296,N_17353);
nor U17543 (N_17543,N_17331,N_17290);
or U17544 (N_17544,N_17256,N_17307);
and U17545 (N_17545,N_17287,N_17315);
nor U17546 (N_17546,N_17254,N_17346);
or U17547 (N_17547,N_17306,N_17239);
nor U17548 (N_17548,N_17203,N_17359);
nand U17549 (N_17549,N_17207,N_17366);
nor U17550 (N_17550,N_17325,N_17371);
and U17551 (N_17551,N_17261,N_17269);
nor U17552 (N_17552,N_17268,N_17300);
nor U17553 (N_17553,N_17238,N_17358);
nor U17554 (N_17554,N_17270,N_17326);
or U17555 (N_17555,N_17277,N_17223);
or U17556 (N_17556,N_17222,N_17243);
nand U17557 (N_17557,N_17347,N_17251);
or U17558 (N_17558,N_17398,N_17244);
and U17559 (N_17559,N_17203,N_17279);
xnor U17560 (N_17560,N_17316,N_17330);
nor U17561 (N_17561,N_17386,N_17363);
or U17562 (N_17562,N_17312,N_17309);
and U17563 (N_17563,N_17260,N_17203);
or U17564 (N_17564,N_17265,N_17371);
and U17565 (N_17565,N_17299,N_17242);
and U17566 (N_17566,N_17383,N_17329);
xnor U17567 (N_17567,N_17379,N_17309);
or U17568 (N_17568,N_17215,N_17399);
and U17569 (N_17569,N_17347,N_17218);
xor U17570 (N_17570,N_17367,N_17337);
nand U17571 (N_17571,N_17280,N_17361);
xor U17572 (N_17572,N_17331,N_17234);
nand U17573 (N_17573,N_17367,N_17216);
nand U17574 (N_17574,N_17257,N_17268);
and U17575 (N_17575,N_17354,N_17301);
nand U17576 (N_17576,N_17394,N_17239);
xnor U17577 (N_17577,N_17316,N_17275);
or U17578 (N_17578,N_17311,N_17384);
nand U17579 (N_17579,N_17270,N_17253);
nand U17580 (N_17580,N_17250,N_17384);
xnor U17581 (N_17581,N_17328,N_17368);
and U17582 (N_17582,N_17266,N_17364);
or U17583 (N_17583,N_17390,N_17211);
or U17584 (N_17584,N_17357,N_17279);
and U17585 (N_17585,N_17377,N_17253);
xor U17586 (N_17586,N_17305,N_17264);
nand U17587 (N_17587,N_17246,N_17391);
and U17588 (N_17588,N_17352,N_17396);
nor U17589 (N_17589,N_17203,N_17277);
nand U17590 (N_17590,N_17354,N_17309);
and U17591 (N_17591,N_17372,N_17242);
or U17592 (N_17592,N_17202,N_17349);
nor U17593 (N_17593,N_17351,N_17231);
and U17594 (N_17594,N_17335,N_17390);
nor U17595 (N_17595,N_17381,N_17220);
nor U17596 (N_17596,N_17388,N_17281);
xor U17597 (N_17597,N_17214,N_17308);
or U17598 (N_17598,N_17279,N_17231);
and U17599 (N_17599,N_17216,N_17361);
and U17600 (N_17600,N_17551,N_17486);
nor U17601 (N_17601,N_17539,N_17590);
and U17602 (N_17602,N_17589,N_17520);
or U17603 (N_17603,N_17555,N_17548);
and U17604 (N_17604,N_17402,N_17403);
xnor U17605 (N_17605,N_17412,N_17511);
xor U17606 (N_17606,N_17411,N_17429);
xor U17607 (N_17607,N_17423,N_17501);
and U17608 (N_17608,N_17512,N_17453);
and U17609 (N_17609,N_17416,N_17533);
nor U17610 (N_17610,N_17503,N_17461);
nor U17611 (N_17611,N_17581,N_17517);
nand U17612 (N_17612,N_17466,N_17424);
or U17613 (N_17613,N_17550,N_17583);
xor U17614 (N_17614,N_17495,N_17440);
and U17615 (N_17615,N_17490,N_17471);
nand U17616 (N_17616,N_17454,N_17469);
or U17617 (N_17617,N_17561,N_17530);
and U17618 (N_17618,N_17518,N_17436);
or U17619 (N_17619,N_17558,N_17541);
and U17620 (N_17620,N_17527,N_17578);
nor U17621 (N_17621,N_17542,N_17462);
and U17622 (N_17622,N_17475,N_17405);
and U17623 (N_17623,N_17445,N_17477);
xor U17624 (N_17624,N_17594,N_17598);
or U17625 (N_17625,N_17443,N_17513);
nand U17626 (N_17626,N_17549,N_17450);
xor U17627 (N_17627,N_17498,N_17409);
nor U17628 (N_17628,N_17444,N_17468);
xnor U17629 (N_17629,N_17597,N_17474);
or U17630 (N_17630,N_17588,N_17400);
nand U17631 (N_17631,N_17569,N_17538);
and U17632 (N_17632,N_17565,N_17419);
nor U17633 (N_17633,N_17582,N_17510);
nand U17634 (N_17634,N_17413,N_17570);
or U17635 (N_17635,N_17430,N_17485);
nand U17636 (N_17636,N_17425,N_17407);
or U17637 (N_17637,N_17532,N_17516);
and U17638 (N_17638,N_17492,N_17448);
or U17639 (N_17639,N_17568,N_17553);
xor U17640 (N_17640,N_17526,N_17507);
or U17641 (N_17641,N_17540,N_17500);
nor U17642 (N_17642,N_17427,N_17567);
nand U17643 (N_17643,N_17459,N_17487);
or U17644 (N_17644,N_17547,N_17483);
xnor U17645 (N_17645,N_17446,N_17408);
nand U17646 (N_17646,N_17438,N_17496);
nand U17647 (N_17647,N_17531,N_17580);
and U17648 (N_17648,N_17599,N_17519);
and U17649 (N_17649,N_17481,N_17447);
nor U17650 (N_17650,N_17441,N_17595);
nand U17651 (N_17651,N_17417,N_17451);
nor U17652 (N_17652,N_17428,N_17418);
nor U17653 (N_17653,N_17470,N_17457);
xnor U17654 (N_17654,N_17494,N_17421);
nand U17655 (N_17655,N_17571,N_17489);
or U17656 (N_17656,N_17509,N_17562);
and U17657 (N_17657,N_17563,N_17442);
or U17658 (N_17658,N_17506,N_17593);
nor U17659 (N_17659,N_17596,N_17502);
nor U17660 (N_17660,N_17406,N_17434);
and U17661 (N_17661,N_17410,N_17432);
nor U17662 (N_17662,N_17585,N_17437);
and U17663 (N_17663,N_17505,N_17479);
nor U17664 (N_17664,N_17433,N_17404);
or U17665 (N_17665,N_17534,N_17439);
xor U17666 (N_17666,N_17420,N_17452);
and U17667 (N_17667,N_17573,N_17545);
nor U17668 (N_17668,N_17480,N_17478);
xnor U17669 (N_17669,N_17491,N_17586);
nand U17670 (N_17670,N_17525,N_17514);
or U17671 (N_17671,N_17576,N_17546);
or U17672 (N_17672,N_17463,N_17464);
xnor U17673 (N_17673,N_17499,N_17488);
nand U17674 (N_17674,N_17473,N_17587);
xnor U17675 (N_17675,N_17435,N_17415);
or U17676 (N_17676,N_17557,N_17426);
nand U17677 (N_17677,N_17536,N_17401);
nand U17678 (N_17678,N_17508,N_17472);
nor U17679 (N_17679,N_17560,N_17535);
or U17680 (N_17680,N_17566,N_17572);
nor U17681 (N_17681,N_17543,N_17592);
xor U17682 (N_17682,N_17515,N_17449);
or U17683 (N_17683,N_17552,N_17537);
xnor U17684 (N_17684,N_17524,N_17456);
nand U17685 (N_17685,N_17431,N_17554);
xor U17686 (N_17686,N_17497,N_17584);
xor U17687 (N_17687,N_17579,N_17493);
or U17688 (N_17688,N_17504,N_17529);
nand U17689 (N_17689,N_17523,N_17564);
nor U17690 (N_17690,N_17544,N_17522);
xor U17691 (N_17691,N_17476,N_17575);
or U17692 (N_17692,N_17521,N_17414);
nand U17693 (N_17693,N_17528,N_17465);
or U17694 (N_17694,N_17422,N_17556);
and U17695 (N_17695,N_17577,N_17455);
nor U17696 (N_17696,N_17574,N_17482);
or U17697 (N_17697,N_17559,N_17460);
nand U17698 (N_17698,N_17467,N_17458);
nand U17699 (N_17699,N_17484,N_17591);
xor U17700 (N_17700,N_17542,N_17506);
nand U17701 (N_17701,N_17527,N_17589);
and U17702 (N_17702,N_17523,N_17449);
nand U17703 (N_17703,N_17506,N_17409);
nand U17704 (N_17704,N_17528,N_17537);
nand U17705 (N_17705,N_17420,N_17485);
nor U17706 (N_17706,N_17452,N_17431);
xnor U17707 (N_17707,N_17560,N_17447);
or U17708 (N_17708,N_17535,N_17506);
nor U17709 (N_17709,N_17417,N_17547);
and U17710 (N_17710,N_17545,N_17596);
or U17711 (N_17711,N_17478,N_17425);
xor U17712 (N_17712,N_17431,N_17504);
nand U17713 (N_17713,N_17415,N_17463);
nand U17714 (N_17714,N_17478,N_17599);
and U17715 (N_17715,N_17584,N_17531);
xnor U17716 (N_17716,N_17480,N_17425);
or U17717 (N_17717,N_17490,N_17501);
nor U17718 (N_17718,N_17576,N_17504);
and U17719 (N_17719,N_17481,N_17478);
nand U17720 (N_17720,N_17548,N_17545);
or U17721 (N_17721,N_17541,N_17403);
or U17722 (N_17722,N_17590,N_17538);
xnor U17723 (N_17723,N_17523,N_17574);
nor U17724 (N_17724,N_17479,N_17564);
and U17725 (N_17725,N_17414,N_17406);
and U17726 (N_17726,N_17558,N_17475);
and U17727 (N_17727,N_17594,N_17473);
nor U17728 (N_17728,N_17530,N_17577);
nor U17729 (N_17729,N_17459,N_17539);
and U17730 (N_17730,N_17539,N_17581);
xnor U17731 (N_17731,N_17532,N_17473);
nand U17732 (N_17732,N_17464,N_17544);
or U17733 (N_17733,N_17503,N_17535);
nor U17734 (N_17734,N_17519,N_17551);
or U17735 (N_17735,N_17485,N_17521);
and U17736 (N_17736,N_17567,N_17583);
nor U17737 (N_17737,N_17457,N_17569);
nor U17738 (N_17738,N_17532,N_17586);
and U17739 (N_17739,N_17577,N_17511);
nand U17740 (N_17740,N_17513,N_17589);
nor U17741 (N_17741,N_17527,N_17565);
or U17742 (N_17742,N_17491,N_17402);
nor U17743 (N_17743,N_17510,N_17490);
xnor U17744 (N_17744,N_17516,N_17545);
nand U17745 (N_17745,N_17549,N_17589);
nand U17746 (N_17746,N_17413,N_17524);
nand U17747 (N_17747,N_17479,N_17463);
xor U17748 (N_17748,N_17549,N_17418);
or U17749 (N_17749,N_17480,N_17566);
or U17750 (N_17750,N_17551,N_17453);
xor U17751 (N_17751,N_17427,N_17491);
nor U17752 (N_17752,N_17558,N_17587);
xnor U17753 (N_17753,N_17546,N_17513);
or U17754 (N_17754,N_17457,N_17448);
nor U17755 (N_17755,N_17526,N_17547);
nand U17756 (N_17756,N_17501,N_17459);
or U17757 (N_17757,N_17492,N_17403);
xnor U17758 (N_17758,N_17479,N_17518);
nor U17759 (N_17759,N_17550,N_17548);
nand U17760 (N_17760,N_17526,N_17559);
nor U17761 (N_17761,N_17488,N_17507);
nand U17762 (N_17762,N_17479,N_17551);
or U17763 (N_17763,N_17451,N_17425);
or U17764 (N_17764,N_17569,N_17523);
and U17765 (N_17765,N_17556,N_17528);
xor U17766 (N_17766,N_17533,N_17555);
xor U17767 (N_17767,N_17459,N_17502);
xnor U17768 (N_17768,N_17581,N_17576);
nor U17769 (N_17769,N_17420,N_17491);
xor U17770 (N_17770,N_17539,N_17503);
and U17771 (N_17771,N_17464,N_17426);
xnor U17772 (N_17772,N_17533,N_17500);
or U17773 (N_17773,N_17483,N_17472);
or U17774 (N_17774,N_17563,N_17476);
and U17775 (N_17775,N_17415,N_17462);
and U17776 (N_17776,N_17506,N_17591);
and U17777 (N_17777,N_17475,N_17492);
or U17778 (N_17778,N_17401,N_17549);
xor U17779 (N_17779,N_17488,N_17562);
and U17780 (N_17780,N_17574,N_17554);
nor U17781 (N_17781,N_17563,N_17474);
nor U17782 (N_17782,N_17515,N_17507);
nor U17783 (N_17783,N_17492,N_17478);
nand U17784 (N_17784,N_17542,N_17437);
xnor U17785 (N_17785,N_17536,N_17581);
and U17786 (N_17786,N_17427,N_17499);
nand U17787 (N_17787,N_17547,N_17572);
nand U17788 (N_17788,N_17553,N_17564);
or U17789 (N_17789,N_17532,N_17411);
or U17790 (N_17790,N_17408,N_17427);
nor U17791 (N_17791,N_17454,N_17533);
or U17792 (N_17792,N_17422,N_17589);
nand U17793 (N_17793,N_17517,N_17455);
and U17794 (N_17794,N_17509,N_17550);
or U17795 (N_17795,N_17405,N_17562);
nand U17796 (N_17796,N_17413,N_17542);
or U17797 (N_17797,N_17426,N_17417);
or U17798 (N_17798,N_17586,N_17523);
nor U17799 (N_17799,N_17444,N_17501);
nand U17800 (N_17800,N_17621,N_17667);
nand U17801 (N_17801,N_17654,N_17758);
or U17802 (N_17802,N_17774,N_17742);
or U17803 (N_17803,N_17727,N_17629);
or U17804 (N_17804,N_17648,N_17757);
or U17805 (N_17805,N_17668,N_17689);
nor U17806 (N_17806,N_17790,N_17762);
and U17807 (N_17807,N_17747,N_17679);
xor U17808 (N_17808,N_17680,N_17616);
nor U17809 (N_17809,N_17661,N_17746);
xnor U17810 (N_17810,N_17653,N_17763);
or U17811 (N_17811,N_17701,N_17752);
xor U17812 (N_17812,N_17784,N_17641);
xor U17813 (N_17813,N_17755,N_17799);
nor U17814 (N_17814,N_17764,N_17712);
xnor U17815 (N_17815,N_17726,N_17602);
xor U17816 (N_17816,N_17776,N_17778);
or U17817 (N_17817,N_17618,N_17798);
or U17818 (N_17818,N_17739,N_17636);
xor U17819 (N_17819,N_17625,N_17714);
or U17820 (N_17820,N_17611,N_17786);
nor U17821 (N_17821,N_17657,N_17613);
or U17822 (N_17822,N_17633,N_17745);
nand U17823 (N_17823,N_17743,N_17619);
xor U17824 (N_17824,N_17687,N_17785);
xor U17825 (N_17825,N_17777,N_17637);
xor U17826 (N_17826,N_17646,N_17794);
or U17827 (N_17827,N_17631,N_17634);
nand U17828 (N_17828,N_17605,N_17649);
nand U17829 (N_17829,N_17644,N_17737);
nor U17830 (N_17830,N_17734,N_17783);
or U17831 (N_17831,N_17789,N_17676);
or U17832 (N_17832,N_17732,N_17688);
and U17833 (N_17833,N_17779,N_17756);
nor U17834 (N_17834,N_17738,N_17693);
or U17835 (N_17835,N_17719,N_17640);
xor U17836 (N_17836,N_17761,N_17682);
or U17837 (N_17837,N_17673,N_17768);
and U17838 (N_17838,N_17706,N_17659);
nand U17839 (N_17839,N_17665,N_17696);
nor U17840 (N_17840,N_17617,N_17697);
or U17841 (N_17841,N_17788,N_17632);
or U17842 (N_17842,N_17702,N_17751);
nand U17843 (N_17843,N_17769,N_17700);
nand U17844 (N_17844,N_17626,N_17715);
and U17845 (N_17845,N_17683,N_17759);
and U17846 (N_17846,N_17627,N_17717);
and U17847 (N_17847,N_17698,N_17670);
or U17848 (N_17848,N_17731,N_17672);
and U17849 (N_17849,N_17730,N_17674);
or U17850 (N_17850,N_17782,N_17638);
nor U17851 (N_17851,N_17750,N_17623);
nand U17852 (N_17852,N_17787,N_17615);
xnor U17853 (N_17853,N_17710,N_17694);
or U17854 (N_17854,N_17797,N_17642);
or U17855 (N_17855,N_17766,N_17760);
nor U17856 (N_17856,N_17610,N_17724);
nor U17857 (N_17857,N_17614,N_17684);
nor U17858 (N_17858,N_17728,N_17772);
nor U17859 (N_17859,N_17666,N_17681);
nand U17860 (N_17860,N_17663,N_17690);
and U17861 (N_17861,N_17765,N_17624);
nand U17862 (N_17862,N_17645,N_17740);
and U17863 (N_17863,N_17741,N_17716);
and U17864 (N_17864,N_17600,N_17733);
nand U17865 (N_17865,N_17604,N_17669);
xor U17866 (N_17866,N_17647,N_17664);
nor U17867 (N_17867,N_17713,N_17792);
xor U17868 (N_17868,N_17748,N_17795);
or U17869 (N_17869,N_17707,N_17630);
nand U17870 (N_17870,N_17705,N_17695);
or U17871 (N_17871,N_17671,N_17767);
xnor U17872 (N_17872,N_17791,N_17651);
nand U17873 (N_17873,N_17662,N_17639);
or U17874 (N_17874,N_17780,N_17607);
or U17875 (N_17875,N_17675,N_17796);
nor U17876 (N_17876,N_17773,N_17704);
nor U17877 (N_17877,N_17685,N_17736);
nor U17878 (N_17878,N_17708,N_17793);
nor U17879 (N_17879,N_17606,N_17622);
xor U17880 (N_17880,N_17753,N_17729);
nand U17881 (N_17881,N_17749,N_17620);
nand U17882 (N_17882,N_17628,N_17658);
xor U17883 (N_17883,N_17711,N_17735);
nand U17884 (N_17884,N_17723,N_17775);
or U17885 (N_17885,N_17678,N_17643);
or U17886 (N_17886,N_17703,N_17601);
and U17887 (N_17887,N_17652,N_17692);
nand U17888 (N_17888,N_17709,N_17603);
nand U17889 (N_17889,N_17770,N_17699);
nand U17890 (N_17890,N_17660,N_17771);
nand U17891 (N_17891,N_17720,N_17612);
or U17892 (N_17892,N_17635,N_17608);
nand U17893 (N_17893,N_17650,N_17718);
and U17894 (N_17894,N_17754,N_17725);
and U17895 (N_17895,N_17655,N_17722);
xnor U17896 (N_17896,N_17721,N_17744);
nand U17897 (N_17897,N_17781,N_17686);
and U17898 (N_17898,N_17656,N_17609);
xnor U17899 (N_17899,N_17677,N_17691);
or U17900 (N_17900,N_17698,N_17661);
nand U17901 (N_17901,N_17774,N_17665);
xor U17902 (N_17902,N_17733,N_17758);
or U17903 (N_17903,N_17728,N_17705);
xnor U17904 (N_17904,N_17710,N_17685);
nor U17905 (N_17905,N_17709,N_17602);
or U17906 (N_17906,N_17721,N_17675);
or U17907 (N_17907,N_17609,N_17761);
and U17908 (N_17908,N_17695,N_17693);
xor U17909 (N_17909,N_17683,N_17675);
xor U17910 (N_17910,N_17616,N_17791);
and U17911 (N_17911,N_17658,N_17610);
nand U17912 (N_17912,N_17712,N_17762);
nor U17913 (N_17913,N_17614,N_17750);
nand U17914 (N_17914,N_17655,N_17624);
xnor U17915 (N_17915,N_17654,N_17669);
or U17916 (N_17916,N_17689,N_17649);
nand U17917 (N_17917,N_17647,N_17615);
xnor U17918 (N_17918,N_17730,N_17768);
and U17919 (N_17919,N_17732,N_17637);
nor U17920 (N_17920,N_17697,N_17797);
xnor U17921 (N_17921,N_17717,N_17715);
nand U17922 (N_17922,N_17705,N_17799);
nor U17923 (N_17923,N_17688,N_17779);
nor U17924 (N_17924,N_17676,N_17660);
or U17925 (N_17925,N_17613,N_17649);
or U17926 (N_17926,N_17697,N_17785);
and U17927 (N_17927,N_17758,N_17773);
nand U17928 (N_17928,N_17614,N_17799);
xor U17929 (N_17929,N_17795,N_17714);
xor U17930 (N_17930,N_17624,N_17676);
or U17931 (N_17931,N_17643,N_17685);
or U17932 (N_17932,N_17708,N_17734);
nor U17933 (N_17933,N_17757,N_17643);
xnor U17934 (N_17934,N_17735,N_17621);
or U17935 (N_17935,N_17632,N_17722);
xnor U17936 (N_17936,N_17647,N_17665);
xor U17937 (N_17937,N_17678,N_17687);
xnor U17938 (N_17938,N_17634,N_17628);
and U17939 (N_17939,N_17766,N_17662);
and U17940 (N_17940,N_17734,N_17774);
nand U17941 (N_17941,N_17706,N_17756);
and U17942 (N_17942,N_17750,N_17682);
nand U17943 (N_17943,N_17707,N_17600);
and U17944 (N_17944,N_17612,N_17704);
or U17945 (N_17945,N_17735,N_17609);
nor U17946 (N_17946,N_17722,N_17788);
or U17947 (N_17947,N_17781,N_17703);
xor U17948 (N_17948,N_17723,N_17670);
and U17949 (N_17949,N_17653,N_17764);
or U17950 (N_17950,N_17610,N_17653);
or U17951 (N_17951,N_17691,N_17615);
nor U17952 (N_17952,N_17777,N_17796);
nor U17953 (N_17953,N_17654,N_17730);
and U17954 (N_17954,N_17746,N_17775);
xor U17955 (N_17955,N_17650,N_17692);
and U17956 (N_17956,N_17750,N_17764);
nor U17957 (N_17957,N_17722,N_17643);
and U17958 (N_17958,N_17716,N_17691);
or U17959 (N_17959,N_17650,N_17706);
and U17960 (N_17960,N_17683,N_17684);
xor U17961 (N_17961,N_17756,N_17602);
nand U17962 (N_17962,N_17734,N_17772);
and U17963 (N_17963,N_17706,N_17779);
nor U17964 (N_17964,N_17735,N_17782);
nor U17965 (N_17965,N_17736,N_17678);
nand U17966 (N_17966,N_17789,N_17771);
nand U17967 (N_17967,N_17718,N_17793);
nor U17968 (N_17968,N_17617,N_17791);
nor U17969 (N_17969,N_17797,N_17738);
nand U17970 (N_17970,N_17663,N_17640);
xor U17971 (N_17971,N_17721,N_17726);
and U17972 (N_17972,N_17758,N_17761);
and U17973 (N_17973,N_17717,N_17691);
or U17974 (N_17974,N_17787,N_17608);
nand U17975 (N_17975,N_17732,N_17613);
or U17976 (N_17976,N_17661,N_17672);
nand U17977 (N_17977,N_17761,N_17605);
and U17978 (N_17978,N_17648,N_17698);
or U17979 (N_17979,N_17715,N_17712);
and U17980 (N_17980,N_17727,N_17721);
and U17981 (N_17981,N_17798,N_17704);
nand U17982 (N_17982,N_17652,N_17725);
xor U17983 (N_17983,N_17661,N_17683);
nand U17984 (N_17984,N_17753,N_17637);
nor U17985 (N_17985,N_17679,N_17717);
xor U17986 (N_17986,N_17652,N_17743);
nand U17987 (N_17987,N_17733,N_17791);
or U17988 (N_17988,N_17743,N_17765);
nand U17989 (N_17989,N_17781,N_17788);
or U17990 (N_17990,N_17635,N_17798);
nor U17991 (N_17991,N_17777,N_17769);
xnor U17992 (N_17992,N_17672,N_17651);
or U17993 (N_17993,N_17744,N_17691);
nor U17994 (N_17994,N_17774,N_17670);
nor U17995 (N_17995,N_17648,N_17730);
nor U17996 (N_17996,N_17719,N_17714);
or U17997 (N_17997,N_17771,N_17601);
nor U17998 (N_17998,N_17783,N_17741);
nand U17999 (N_17999,N_17790,N_17600);
nand U18000 (N_18000,N_17823,N_17873);
nand U18001 (N_18001,N_17901,N_17822);
nor U18002 (N_18002,N_17881,N_17907);
nand U18003 (N_18003,N_17933,N_17999);
xnor U18004 (N_18004,N_17997,N_17819);
or U18005 (N_18005,N_17812,N_17824);
nand U18006 (N_18006,N_17930,N_17856);
or U18007 (N_18007,N_17820,N_17831);
nand U18008 (N_18008,N_17804,N_17991);
and U18009 (N_18009,N_17803,N_17946);
xnor U18010 (N_18010,N_17979,N_17854);
and U18011 (N_18011,N_17852,N_17877);
nor U18012 (N_18012,N_17943,N_17821);
nor U18013 (N_18013,N_17968,N_17818);
xnor U18014 (N_18014,N_17983,N_17861);
nand U18015 (N_18015,N_17964,N_17934);
xor U18016 (N_18016,N_17848,N_17838);
or U18017 (N_18017,N_17816,N_17894);
nor U18018 (N_18018,N_17951,N_17844);
nand U18019 (N_18019,N_17898,N_17817);
xor U18020 (N_18020,N_17839,N_17875);
or U18021 (N_18021,N_17961,N_17887);
nand U18022 (N_18022,N_17928,N_17906);
xor U18023 (N_18023,N_17802,N_17940);
or U18024 (N_18024,N_17919,N_17902);
and U18025 (N_18025,N_17895,N_17865);
and U18026 (N_18026,N_17850,N_17973);
or U18027 (N_18027,N_17886,N_17927);
nand U18028 (N_18028,N_17845,N_17932);
nand U18029 (N_18029,N_17834,N_17897);
and U18030 (N_18030,N_17936,N_17876);
xor U18031 (N_18031,N_17862,N_17908);
and U18032 (N_18032,N_17892,N_17958);
xor U18033 (N_18033,N_17985,N_17893);
and U18034 (N_18034,N_17939,N_17984);
nor U18035 (N_18035,N_17801,N_17885);
or U18036 (N_18036,N_17829,N_17814);
nor U18037 (N_18037,N_17981,N_17912);
xnor U18038 (N_18038,N_17995,N_17855);
nor U18039 (N_18039,N_17952,N_17948);
and U18040 (N_18040,N_17996,N_17921);
nor U18041 (N_18041,N_17903,N_17994);
and U18042 (N_18042,N_17860,N_17840);
nor U18043 (N_18043,N_17828,N_17851);
xor U18044 (N_18044,N_17805,N_17953);
nor U18045 (N_18045,N_17896,N_17858);
and U18046 (N_18046,N_17917,N_17808);
nand U18047 (N_18047,N_17807,N_17972);
nor U18048 (N_18048,N_17969,N_17869);
nand U18049 (N_18049,N_17947,N_17986);
nor U18050 (N_18050,N_17910,N_17827);
or U18051 (N_18051,N_17931,N_17900);
nand U18052 (N_18052,N_17954,N_17843);
or U18053 (N_18053,N_17905,N_17925);
or U18054 (N_18054,N_17920,N_17945);
or U18055 (N_18055,N_17915,N_17842);
or U18056 (N_18056,N_17941,N_17809);
nand U18057 (N_18057,N_17811,N_17864);
xor U18058 (N_18058,N_17857,N_17863);
and U18059 (N_18059,N_17955,N_17993);
nand U18060 (N_18060,N_17882,N_17975);
or U18061 (N_18061,N_17835,N_17880);
or U18062 (N_18062,N_17868,N_17833);
or U18063 (N_18063,N_17935,N_17988);
or U18064 (N_18064,N_17942,N_17825);
nand U18065 (N_18065,N_17890,N_17916);
nand U18066 (N_18066,N_17978,N_17965);
and U18067 (N_18067,N_17909,N_17974);
xor U18068 (N_18068,N_17982,N_17963);
nand U18069 (N_18069,N_17967,N_17923);
and U18070 (N_18070,N_17966,N_17846);
xnor U18071 (N_18071,N_17976,N_17980);
or U18072 (N_18072,N_17841,N_17849);
nand U18073 (N_18073,N_17938,N_17911);
or U18074 (N_18074,N_17957,N_17806);
xnor U18075 (N_18075,N_17826,N_17918);
xnor U18076 (N_18076,N_17870,N_17949);
nor U18077 (N_18077,N_17832,N_17971);
and U18078 (N_18078,N_17891,N_17914);
and U18079 (N_18079,N_17924,N_17960);
nand U18080 (N_18080,N_17987,N_17853);
nor U18081 (N_18081,N_17889,N_17970);
xnor U18082 (N_18082,N_17883,N_17859);
and U18083 (N_18083,N_17837,N_17810);
nor U18084 (N_18084,N_17815,N_17962);
xor U18085 (N_18085,N_17888,N_17878);
xnor U18086 (N_18086,N_17904,N_17989);
nand U18087 (N_18087,N_17836,N_17871);
nor U18088 (N_18088,N_17992,N_17959);
nand U18089 (N_18089,N_17872,N_17884);
nand U18090 (N_18090,N_17899,N_17977);
and U18091 (N_18091,N_17830,N_17937);
or U18092 (N_18092,N_17998,N_17800);
or U18093 (N_18093,N_17956,N_17944);
xnor U18094 (N_18094,N_17847,N_17813);
or U18095 (N_18095,N_17867,N_17922);
xor U18096 (N_18096,N_17866,N_17879);
xor U18097 (N_18097,N_17874,N_17950);
nand U18098 (N_18098,N_17990,N_17929);
or U18099 (N_18099,N_17926,N_17913);
nor U18100 (N_18100,N_17843,N_17858);
or U18101 (N_18101,N_17907,N_17801);
or U18102 (N_18102,N_17859,N_17868);
nor U18103 (N_18103,N_17847,N_17855);
nor U18104 (N_18104,N_17914,N_17916);
nor U18105 (N_18105,N_17997,N_17855);
xor U18106 (N_18106,N_17825,N_17930);
nand U18107 (N_18107,N_17833,N_17924);
nor U18108 (N_18108,N_17920,N_17852);
xor U18109 (N_18109,N_17915,N_17909);
xor U18110 (N_18110,N_17822,N_17860);
and U18111 (N_18111,N_17803,N_17888);
and U18112 (N_18112,N_17863,N_17906);
and U18113 (N_18113,N_17860,N_17990);
nand U18114 (N_18114,N_17923,N_17993);
nand U18115 (N_18115,N_17865,N_17806);
nand U18116 (N_18116,N_17924,N_17923);
or U18117 (N_18117,N_17900,N_17886);
or U18118 (N_18118,N_17898,N_17805);
nand U18119 (N_18119,N_17881,N_17932);
xnor U18120 (N_18120,N_17999,N_17837);
nor U18121 (N_18121,N_17820,N_17852);
nand U18122 (N_18122,N_17951,N_17935);
nor U18123 (N_18123,N_17806,N_17886);
xor U18124 (N_18124,N_17933,N_17885);
nor U18125 (N_18125,N_17882,N_17950);
nand U18126 (N_18126,N_17926,N_17841);
xnor U18127 (N_18127,N_17936,N_17962);
xor U18128 (N_18128,N_17949,N_17974);
xnor U18129 (N_18129,N_17929,N_17914);
xnor U18130 (N_18130,N_17959,N_17877);
and U18131 (N_18131,N_17887,N_17837);
xnor U18132 (N_18132,N_17885,N_17805);
xor U18133 (N_18133,N_17830,N_17804);
xor U18134 (N_18134,N_17929,N_17948);
nand U18135 (N_18135,N_17849,N_17838);
xor U18136 (N_18136,N_17956,N_17805);
and U18137 (N_18137,N_17930,N_17803);
nor U18138 (N_18138,N_17807,N_17889);
nand U18139 (N_18139,N_17920,N_17815);
nand U18140 (N_18140,N_17924,N_17952);
nor U18141 (N_18141,N_17876,N_17976);
nand U18142 (N_18142,N_17860,N_17874);
xnor U18143 (N_18143,N_17998,N_17824);
nand U18144 (N_18144,N_17859,N_17827);
or U18145 (N_18145,N_17998,N_17924);
xor U18146 (N_18146,N_17804,N_17995);
nor U18147 (N_18147,N_17984,N_17805);
xor U18148 (N_18148,N_17855,N_17982);
xnor U18149 (N_18149,N_17802,N_17835);
nand U18150 (N_18150,N_17984,N_17835);
xnor U18151 (N_18151,N_17950,N_17989);
nor U18152 (N_18152,N_17868,N_17805);
nor U18153 (N_18153,N_17877,N_17969);
nand U18154 (N_18154,N_17877,N_17961);
xnor U18155 (N_18155,N_17842,N_17880);
or U18156 (N_18156,N_17894,N_17972);
or U18157 (N_18157,N_17866,N_17970);
nor U18158 (N_18158,N_17846,N_17986);
or U18159 (N_18159,N_17959,N_17987);
xor U18160 (N_18160,N_17959,N_17931);
xor U18161 (N_18161,N_17979,N_17917);
nand U18162 (N_18162,N_17841,N_17814);
and U18163 (N_18163,N_17909,N_17815);
and U18164 (N_18164,N_17864,N_17827);
nand U18165 (N_18165,N_17878,N_17938);
nand U18166 (N_18166,N_17988,N_17883);
nor U18167 (N_18167,N_17929,N_17979);
and U18168 (N_18168,N_17817,N_17806);
or U18169 (N_18169,N_17850,N_17936);
xor U18170 (N_18170,N_17916,N_17822);
or U18171 (N_18171,N_17950,N_17856);
xor U18172 (N_18172,N_17953,N_17922);
nor U18173 (N_18173,N_17962,N_17836);
and U18174 (N_18174,N_17975,N_17957);
nand U18175 (N_18175,N_17929,N_17830);
xnor U18176 (N_18176,N_17975,N_17891);
or U18177 (N_18177,N_17978,N_17963);
nand U18178 (N_18178,N_17849,N_17810);
xor U18179 (N_18179,N_17954,N_17810);
nor U18180 (N_18180,N_17847,N_17862);
and U18181 (N_18181,N_17947,N_17834);
nor U18182 (N_18182,N_17876,N_17853);
nand U18183 (N_18183,N_17826,N_17907);
and U18184 (N_18184,N_17942,N_17973);
xor U18185 (N_18185,N_17931,N_17956);
nor U18186 (N_18186,N_17827,N_17877);
or U18187 (N_18187,N_17855,N_17974);
xor U18188 (N_18188,N_17988,N_17903);
or U18189 (N_18189,N_17818,N_17999);
nand U18190 (N_18190,N_17965,N_17993);
nor U18191 (N_18191,N_17996,N_17948);
and U18192 (N_18192,N_17895,N_17823);
or U18193 (N_18193,N_17948,N_17967);
and U18194 (N_18194,N_17947,N_17874);
and U18195 (N_18195,N_17888,N_17853);
nand U18196 (N_18196,N_17957,N_17938);
nor U18197 (N_18197,N_17950,N_17879);
or U18198 (N_18198,N_17952,N_17839);
or U18199 (N_18199,N_17898,N_17992);
xor U18200 (N_18200,N_18160,N_18020);
nor U18201 (N_18201,N_18129,N_18078);
and U18202 (N_18202,N_18192,N_18029);
and U18203 (N_18203,N_18105,N_18171);
and U18204 (N_18204,N_18038,N_18065);
nand U18205 (N_18205,N_18079,N_18043);
nand U18206 (N_18206,N_18115,N_18170);
and U18207 (N_18207,N_18062,N_18163);
nand U18208 (N_18208,N_18000,N_18179);
and U18209 (N_18209,N_18198,N_18197);
or U18210 (N_18210,N_18025,N_18026);
nor U18211 (N_18211,N_18044,N_18128);
nand U18212 (N_18212,N_18089,N_18074);
or U18213 (N_18213,N_18070,N_18094);
or U18214 (N_18214,N_18085,N_18185);
or U18215 (N_18215,N_18072,N_18154);
or U18216 (N_18216,N_18075,N_18058);
nor U18217 (N_18217,N_18112,N_18022);
nor U18218 (N_18218,N_18139,N_18186);
nor U18219 (N_18219,N_18162,N_18141);
and U18220 (N_18220,N_18104,N_18155);
nor U18221 (N_18221,N_18190,N_18123);
and U18222 (N_18222,N_18042,N_18133);
nor U18223 (N_18223,N_18030,N_18173);
nor U18224 (N_18224,N_18084,N_18066);
nor U18225 (N_18225,N_18068,N_18165);
nand U18226 (N_18226,N_18087,N_18049);
xnor U18227 (N_18227,N_18125,N_18191);
and U18228 (N_18228,N_18111,N_18081);
xor U18229 (N_18229,N_18161,N_18177);
or U18230 (N_18230,N_18059,N_18151);
nand U18231 (N_18231,N_18187,N_18095);
nor U18232 (N_18232,N_18109,N_18144);
nand U18233 (N_18233,N_18126,N_18047);
nand U18234 (N_18234,N_18060,N_18182);
and U18235 (N_18235,N_18132,N_18031);
or U18236 (N_18236,N_18122,N_18184);
or U18237 (N_18237,N_18120,N_18054);
xor U18238 (N_18238,N_18166,N_18008);
xor U18239 (N_18239,N_18015,N_18053);
nor U18240 (N_18240,N_18093,N_18032);
nand U18241 (N_18241,N_18052,N_18037);
xnor U18242 (N_18242,N_18056,N_18013);
xnor U18243 (N_18243,N_18168,N_18157);
and U18244 (N_18244,N_18117,N_18045);
and U18245 (N_18245,N_18135,N_18082);
nor U18246 (N_18246,N_18012,N_18131);
xor U18247 (N_18247,N_18021,N_18127);
nor U18248 (N_18248,N_18167,N_18050);
and U18249 (N_18249,N_18034,N_18090);
nand U18250 (N_18250,N_18069,N_18039);
nand U18251 (N_18251,N_18083,N_18147);
and U18252 (N_18252,N_18103,N_18033);
or U18253 (N_18253,N_18016,N_18011);
xor U18254 (N_18254,N_18143,N_18027);
and U18255 (N_18255,N_18193,N_18055);
nor U18256 (N_18256,N_18181,N_18010);
nor U18257 (N_18257,N_18051,N_18017);
nand U18258 (N_18258,N_18110,N_18116);
or U18259 (N_18259,N_18099,N_18091);
xor U18260 (N_18260,N_18114,N_18001);
nand U18261 (N_18261,N_18145,N_18118);
xnor U18262 (N_18262,N_18063,N_18149);
and U18263 (N_18263,N_18180,N_18005);
and U18264 (N_18264,N_18014,N_18004);
or U18265 (N_18265,N_18088,N_18189);
xnor U18266 (N_18266,N_18048,N_18137);
xor U18267 (N_18267,N_18130,N_18156);
nand U18268 (N_18268,N_18196,N_18086);
xnor U18269 (N_18269,N_18077,N_18152);
or U18270 (N_18270,N_18002,N_18134);
xor U18271 (N_18271,N_18100,N_18019);
nor U18272 (N_18272,N_18153,N_18124);
nand U18273 (N_18273,N_18057,N_18023);
nand U18274 (N_18274,N_18178,N_18041);
nor U18275 (N_18275,N_18195,N_18106);
and U18276 (N_18276,N_18024,N_18183);
xnor U18277 (N_18277,N_18148,N_18092);
xor U18278 (N_18278,N_18175,N_18146);
or U18279 (N_18279,N_18073,N_18028);
nand U18280 (N_18280,N_18119,N_18009);
xnor U18281 (N_18281,N_18046,N_18061);
nor U18282 (N_18282,N_18101,N_18006);
xnor U18283 (N_18283,N_18113,N_18199);
and U18284 (N_18284,N_18188,N_18142);
nand U18285 (N_18285,N_18140,N_18067);
nor U18286 (N_18286,N_18003,N_18040);
or U18287 (N_18287,N_18071,N_18007);
or U18288 (N_18288,N_18018,N_18194);
xnor U18289 (N_18289,N_18172,N_18064);
nor U18290 (N_18290,N_18107,N_18108);
xor U18291 (N_18291,N_18158,N_18164);
nor U18292 (N_18292,N_18150,N_18098);
xnor U18293 (N_18293,N_18121,N_18136);
or U18294 (N_18294,N_18036,N_18035);
or U18295 (N_18295,N_18096,N_18174);
nand U18296 (N_18296,N_18169,N_18076);
xor U18297 (N_18297,N_18097,N_18080);
or U18298 (N_18298,N_18159,N_18138);
or U18299 (N_18299,N_18176,N_18102);
nand U18300 (N_18300,N_18081,N_18189);
nand U18301 (N_18301,N_18076,N_18182);
nand U18302 (N_18302,N_18175,N_18102);
and U18303 (N_18303,N_18033,N_18023);
or U18304 (N_18304,N_18109,N_18115);
xnor U18305 (N_18305,N_18142,N_18084);
nand U18306 (N_18306,N_18179,N_18015);
or U18307 (N_18307,N_18022,N_18015);
nor U18308 (N_18308,N_18022,N_18023);
nand U18309 (N_18309,N_18138,N_18180);
or U18310 (N_18310,N_18109,N_18040);
or U18311 (N_18311,N_18015,N_18116);
and U18312 (N_18312,N_18056,N_18179);
nand U18313 (N_18313,N_18096,N_18112);
or U18314 (N_18314,N_18002,N_18014);
nand U18315 (N_18315,N_18038,N_18193);
nand U18316 (N_18316,N_18047,N_18128);
xnor U18317 (N_18317,N_18191,N_18070);
or U18318 (N_18318,N_18043,N_18120);
or U18319 (N_18319,N_18083,N_18066);
nand U18320 (N_18320,N_18118,N_18152);
nand U18321 (N_18321,N_18006,N_18068);
nor U18322 (N_18322,N_18115,N_18188);
nand U18323 (N_18323,N_18164,N_18193);
xor U18324 (N_18324,N_18148,N_18042);
nand U18325 (N_18325,N_18138,N_18081);
xnor U18326 (N_18326,N_18179,N_18100);
or U18327 (N_18327,N_18127,N_18068);
or U18328 (N_18328,N_18013,N_18154);
xnor U18329 (N_18329,N_18058,N_18004);
nand U18330 (N_18330,N_18139,N_18120);
nand U18331 (N_18331,N_18115,N_18151);
and U18332 (N_18332,N_18158,N_18083);
and U18333 (N_18333,N_18038,N_18115);
nand U18334 (N_18334,N_18106,N_18008);
nand U18335 (N_18335,N_18152,N_18159);
or U18336 (N_18336,N_18069,N_18193);
xor U18337 (N_18337,N_18132,N_18059);
nor U18338 (N_18338,N_18175,N_18193);
nand U18339 (N_18339,N_18006,N_18123);
xnor U18340 (N_18340,N_18004,N_18088);
or U18341 (N_18341,N_18172,N_18127);
nand U18342 (N_18342,N_18167,N_18006);
nand U18343 (N_18343,N_18099,N_18148);
xor U18344 (N_18344,N_18198,N_18173);
nor U18345 (N_18345,N_18139,N_18168);
xnor U18346 (N_18346,N_18100,N_18025);
or U18347 (N_18347,N_18096,N_18185);
nor U18348 (N_18348,N_18127,N_18175);
nand U18349 (N_18349,N_18131,N_18098);
xnor U18350 (N_18350,N_18061,N_18045);
nand U18351 (N_18351,N_18028,N_18130);
or U18352 (N_18352,N_18037,N_18101);
nand U18353 (N_18353,N_18077,N_18099);
xnor U18354 (N_18354,N_18101,N_18111);
and U18355 (N_18355,N_18192,N_18058);
xor U18356 (N_18356,N_18192,N_18036);
nor U18357 (N_18357,N_18120,N_18049);
xor U18358 (N_18358,N_18191,N_18124);
and U18359 (N_18359,N_18152,N_18012);
or U18360 (N_18360,N_18027,N_18165);
xor U18361 (N_18361,N_18196,N_18183);
xnor U18362 (N_18362,N_18007,N_18181);
and U18363 (N_18363,N_18039,N_18055);
nor U18364 (N_18364,N_18045,N_18179);
nand U18365 (N_18365,N_18105,N_18051);
and U18366 (N_18366,N_18109,N_18026);
nor U18367 (N_18367,N_18035,N_18140);
or U18368 (N_18368,N_18168,N_18051);
xnor U18369 (N_18369,N_18097,N_18015);
or U18370 (N_18370,N_18050,N_18149);
xor U18371 (N_18371,N_18070,N_18151);
xor U18372 (N_18372,N_18170,N_18083);
nand U18373 (N_18373,N_18050,N_18027);
nand U18374 (N_18374,N_18094,N_18065);
xor U18375 (N_18375,N_18084,N_18192);
nand U18376 (N_18376,N_18011,N_18084);
or U18377 (N_18377,N_18129,N_18087);
xnor U18378 (N_18378,N_18132,N_18164);
nand U18379 (N_18379,N_18152,N_18117);
nor U18380 (N_18380,N_18104,N_18122);
or U18381 (N_18381,N_18063,N_18075);
and U18382 (N_18382,N_18113,N_18097);
nand U18383 (N_18383,N_18092,N_18145);
and U18384 (N_18384,N_18056,N_18027);
xnor U18385 (N_18385,N_18009,N_18115);
or U18386 (N_18386,N_18028,N_18157);
or U18387 (N_18387,N_18058,N_18098);
xor U18388 (N_18388,N_18088,N_18116);
xor U18389 (N_18389,N_18199,N_18030);
nand U18390 (N_18390,N_18094,N_18182);
nand U18391 (N_18391,N_18111,N_18109);
and U18392 (N_18392,N_18133,N_18114);
xor U18393 (N_18393,N_18080,N_18177);
xnor U18394 (N_18394,N_18020,N_18154);
nor U18395 (N_18395,N_18043,N_18110);
nand U18396 (N_18396,N_18002,N_18040);
and U18397 (N_18397,N_18048,N_18186);
xor U18398 (N_18398,N_18180,N_18171);
nor U18399 (N_18399,N_18194,N_18108);
xor U18400 (N_18400,N_18355,N_18341);
nand U18401 (N_18401,N_18327,N_18264);
nor U18402 (N_18402,N_18257,N_18283);
nand U18403 (N_18403,N_18316,N_18242);
nand U18404 (N_18404,N_18352,N_18362);
xnor U18405 (N_18405,N_18351,N_18328);
and U18406 (N_18406,N_18388,N_18346);
xnor U18407 (N_18407,N_18286,N_18349);
nand U18408 (N_18408,N_18322,N_18337);
nand U18409 (N_18409,N_18291,N_18356);
xor U18410 (N_18410,N_18266,N_18376);
and U18411 (N_18411,N_18292,N_18323);
nand U18412 (N_18412,N_18299,N_18224);
nor U18413 (N_18413,N_18281,N_18294);
and U18414 (N_18414,N_18343,N_18329);
xnor U18415 (N_18415,N_18339,N_18354);
or U18416 (N_18416,N_18201,N_18295);
xor U18417 (N_18417,N_18317,N_18319);
nor U18418 (N_18418,N_18280,N_18331);
xor U18419 (N_18419,N_18208,N_18240);
or U18420 (N_18420,N_18261,N_18296);
nor U18421 (N_18421,N_18209,N_18350);
nand U18422 (N_18422,N_18321,N_18369);
and U18423 (N_18423,N_18333,N_18393);
nand U18424 (N_18424,N_18255,N_18210);
or U18425 (N_18425,N_18342,N_18326);
nand U18426 (N_18426,N_18310,N_18397);
nor U18427 (N_18427,N_18315,N_18392);
or U18428 (N_18428,N_18248,N_18269);
and U18429 (N_18429,N_18290,N_18345);
and U18430 (N_18430,N_18277,N_18385);
or U18431 (N_18431,N_18231,N_18366);
and U18432 (N_18432,N_18271,N_18212);
nor U18433 (N_18433,N_18359,N_18372);
or U18434 (N_18434,N_18398,N_18311);
nor U18435 (N_18435,N_18222,N_18370);
nor U18436 (N_18436,N_18371,N_18272);
or U18437 (N_18437,N_18226,N_18396);
or U18438 (N_18438,N_18288,N_18206);
nand U18439 (N_18439,N_18344,N_18236);
and U18440 (N_18440,N_18218,N_18249);
nor U18441 (N_18441,N_18330,N_18252);
xor U18442 (N_18442,N_18263,N_18347);
nand U18443 (N_18443,N_18217,N_18304);
nand U18444 (N_18444,N_18320,N_18273);
or U18445 (N_18445,N_18207,N_18293);
nor U18446 (N_18446,N_18307,N_18223);
and U18447 (N_18447,N_18214,N_18363);
nand U18448 (N_18448,N_18309,N_18358);
nand U18449 (N_18449,N_18360,N_18233);
nor U18450 (N_18450,N_18395,N_18379);
xor U18451 (N_18451,N_18243,N_18361);
xor U18452 (N_18452,N_18336,N_18238);
nor U18453 (N_18453,N_18237,N_18260);
or U18454 (N_18454,N_18232,N_18225);
nor U18455 (N_18455,N_18303,N_18332);
xnor U18456 (N_18456,N_18306,N_18340);
nor U18457 (N_18457,N_18205,N_18284);
xnor U18458 (N_18458,N_18251,N_18268);
and U18459 (N_18459,N_18334,N_18270);
or U18460 (N_18460,N_18312,N_18227);
xor U18461 (N_18461,N_18245,N_18386);
and U18462 (N_18462,N_18384,N_18382);
xor U18463 (N_18463,N_18374,N_18367);
xnor U18464 (N_18464,N_18211,N_18200);
xnor U18465 (N_18465,N_18348,N_18254);
and U18466 (N_18466,N_18308,N_18282);
nor U18467 (N_18467,N_18318,N_18324);
or U18468 (N_18468,N_18364,N_18373);
nand U18469 (N_18469,N_18219,N_18338);
xor U18470 (N_18470,N_18241,N_18313);
nor U18471 (N_18471,N_18215,N_18378);
or U18472 (N_18472,N_18297,N_18262);
and U18473 (N_18473,N_18353,N_18253);
nand U18474 (N_18474,N_18213,N_18394);
nand U18475 (N_18475,N_18380,N_18228);
nor U18476 (N_18476,N_18300,N_18368);
nand U18477 (N_18477,N_18305,N_18377);
or U18478 (N_18478,N_18221,N_18234);
nor U18479 (N_18479,N_18230,N_18250);
nand U18480 (N_18480,N_18259,N_18391);
nand U18481 (N_18481,N_18387,N_18229);
or U18482 (N_18482,N_18390,N_18365);
xor U18483 (N_18483,N_18389,N_18239);
xnor U18484 (N_18484,N_18314,N_18375);
nand U18485 (N_18485,N_18202,N_18216);
or U18486 (N_18486,N_18325,N_18246);
nand U18487 (N_18487,N_18285,N_18256);
xor U18488 (N_18488,N_18258,N_18399);
nand U18489 (N_18489,N_18267,N_18275);
xor U18490 (N_18490,N_18289,N_18279);
or U18491 (N_18491,N_18203,N_18302);
nand U18492 (N_18492,N_18265,N_18244);
nand U18493 (N_18493,N_18278,N_18274);
nand U18494 (N_18494,N_18276,N_18204);
nand U18495 (N_18495,N_18235,N_18301);
nand U18496 (N_18496,N_18298,N_18383);
xor U18497 (N_18497,N_18247,N_18381);
xor U18498 (N_18498,N_18220,N_18335);
nand U18499 (N_18499,N_18287,N_18357);
xor U18500 (N_18500,N_18265,N_18329);
xor U18501 (N_18501,N_18275,N_18336);
nand U18502 (N_18502,N_18202,N_18358);
xnor U18503 (N_18503,N_18397,N_18202);
nor U18504 (N_18504,N_18238,N_18347);
and U18505 (N_18505,N_18229,N_18270);
and U18506 (N_18506,N_18217,N_18222);
nand U18507 (N_18507,N_18202,N_18211);
and U18508 (N_18508,N_18224,N_18389);
and U18509 (N_18509,N_18278,N_18236);
and U18510 (N_18510,N_18226,N_18296);
nor U18511 (N_18511,N_18391,N_18280);
nand U18512 (N_18512,N_18374,N_18331);
and U18513 (N_18513,N_18221,N_18360);
nor U18514 (N_18514,N_18200,N_18381);
or U18515 (N_18515,N_18267,N_18356);
nor U18516 (N_18516,N_18308,N_18270);
nand U18517 (N_18517,N_18316,N_18235);
and U18518 (N_18518,N_18222,N_18279);
nor U18519 (N_18519,N_18234,N_18204);
or U18520 (N_18520,N_18343,N_18202);
xnor U18521 (N_18521,N_18348,N_18352);
nor U18522 (N_18522,N_18388,N_18300);
nor U18523 (N_18523,N_18303,N_18354);
nand U18524 (N_18524,N_18260,N_18204);
nand U18525 (N_18525,N_18392,N_18294);
nor U18526 (N_18526,N_18375,N_18346);
nand U18527 (N_18527,N_18336,N_18350);
nor U18528 (N_18528,N_18360,N_18312);
nand U18529 (N_18529,N_18226,N_18366);
and U18530 (N_18530,N_18269,N_18200);
nor U18531 (N_18531,N_18381,N_18223);
and U18532 (N_18532,N_18311,N_18222);
xnor U18533 (N_18533,N_18305,N_18394);
xnor U18534 (N_18534,N_18373,N_18249);
nor U18535 (N_18535,N_18291,N_18226);
nor U18536 (N_18536,N_18284,N_18391);
xor U18537 (N_18537,N_18341,N_18349);
nand U18538 (N_18538,N_18295,N_18215);
and U18539 (N_18539,N_18249,N_18342);
nand U18540 (N_18540,N_18374,N_18354);
xor U18541 (N_18541,N_18320,N_18361);
xor U18542 (N_18542,N_18372,N_18238);
or U18543 (N_18543,N_18206,N_18247);
xor U18544 (N_18544,N_18333,N_18367);
xor U18545 (N_18545,N_18292,N_18299);
nor U18546 (N_18546,N_18354,N_18253);
nand U18547 (N_18547,N_18325,N_18214);
and U18548 (N_18548,N_18282,N_18314);
nand U18549 (N_18549,N_18333,N_18211);
or U18550 (N_18550,N_18281,N_18391);
xnor U18551 (N_18551,N_18320,N_18284);
and U18552 (N_18552,N_18363,N_18370);
or U18553 (N_18553,N_18348,N_18392);
nor U18554 (N_18554,N_18244,N_18288);
nor U18555 (N_18555,N_18291,N_18321);
and U18556 (N_18556,N_18228,N_18254);
and U18557 (N_18557,N_18260,N_18353);
nand U18558 (N_18558,N_18215,N_18318);
or U18559 (N_18559,N_18310,N_18261);
xnor U18560 (N_18560,N_18375,N_18342);
nand U18561 (N_18561,N_18324,N_18396);
nand U18562 (N_18562,N_18344,N_18363);
or U18563 (N_18563,N_18236,N_18283);
nor U18564 (N_18564,N_18277,N_18285);
and U18565 (N_18565,N_18240,N_18223);
and U18566 (N_18566,N_18331,N_18212);
xnor U18567 (N_18567,N_18217,N_18226);
nand U18568 (N_18568,N_18384,N_18310);
or U18569 (N_18569,N_18219,N_18262);
and U18570 (N_18570,N_18206,N_18227);
or U18571 (N_18571,N_18312,N_18310);
and U18572 (N_18572,N_18337,N_18266);
and U18573 (N_18573,N_18223,N_18355);
nand U18574 (N_18574,N_18326,N_18302);
nor U18575 (N_18575,N_18368,N_18321);
and U18576 (N_18576,N_18237,N_18347);
or U18577 (N_18577,N_18208,N_18289);
nor U18578 (N_18578,N_18340,N_18270);
xor U18579 (N_18579,N_18338,N_18293);
and U18580 (N_18580,N_18359,N_18321);
xnor U18581 (N_18581,N_18376,N_18244);
xor U18582 (N_18582,N_18385,N_18218);
or U18583 (N_18583,N_18364,N_18225);
nand U18584 (N_18584,N_18264,N_18284);
or U18585 (N_18585,N_18392,N_18318);
or U18586 (N_18586,N_18397,N_18327);
or U18587 (N_18587,N_18248,N_18381);
nor U18588 (N_18588,N_18286,N_18361);
or U18589 (N_18589,N_18362,N_18247);
xnor U18590 (N_18590,N_18245,N_18334);
or U18591 (N_18591,N_18223,N_18204);
xor U18592 (N_18592,N_18295,N_18291);
or U18593 (N_18593,N_18306,N_18229);
or U18594 (N_18594,N_18239,N_18351);
nand U18595 (N_18595,N_18215,N_18264);
nor U18596 (N_18596,N_18341,N_18346);
and U18597 (N_18597,N_18240,N_18306);
nand U18598 (N_18598,N_18291,N_18399);
nor U18599 (N_18599,N_18346,N_18266);
or U18600 (N_18600,N_18522,N_18518);
nor U18601 (N_18601,N_18593,N_18556);
xnor U18602 (N_18602,N_18525,N_18511);
nor U18603 (N_18603,N_18452,N_18542);
or U18604 (N_18604,N_18442,N_18594);
nor U18605 (N_18605,N_18595,N_18496);
and U18606 (N_18606,N_18422,N_18480);
and U18607 (N_18607,N_18517,N_18408);
xor U18608 (N_18608,N_18471,N_18481);
nand U18609 (N_18609,N_18513,N_18538);
or U18610 (N_18610,N_18430,N_18548);
or U18611 (N_18611,N_18571,N_18494);
xor U18612 (N_18612,N_18493,N_18532);
nand U18613 (N_18613,N_18404,N_18465);
or U18614 (N_18614,N_18438,N_18443);
nor U18615 (N_18615,N_18516,N_18403);
nor U18616 (N_18616,N_18464,N_18551);
nor U18617 (N_18617,N_18509,N_18570);
xnor U18618 (N_18618,N_18425,N_18544);
or U18619 (N_18619,N_18470,N_18417);
nand U18620 (N_18620,N_18599,N_18439);
or U18621 (N_18621,N_18447,N_18483);
nor U18622 (N_18622,N_18562,N_18445);
or U18623 (N_18623,N_18536,N_18486);
and U18624 (N_18624,N_18402,N_18547);
xor U18625 (N_18625,N_18434,N_18411);
xnor U18626 (N_18626,N_18590,N_18441);
xor U18627 (N_18627,N_18416,N_18540);
nor U18628 (N_18628,N_18506,N_18533);
nor U18629 (N_18629,N_18484,N_18576);
xnor U18630 (N_18630,N_18567,N_18529);
xor U18631 (N_18631,N_18444,N_18499);
nand U18632 (N_18632,N_18453,N_18539);
or U18633 (N_18633,N_18462,N_18450);
nand U18634 (N_18634,N_18437,N_18427);
and U18635 (N_18635,N_18466,N_18420);
nor U18636 (N_18636,N_18467,N_18561);
or U18637 (N_18637,N_18537,N_18559);
nor U18638 (N_18638,N_18456,N_18419);
nand U18639 (N_18639,N_18498,N_18526);
and U18640 (N_18640,N_18401,N_18565);
nand U18641 (N_18641,N_18508,N_18545);
and U18642 (N_18642,N_18431,N_18578);
nand U18643 (N_18643,N_18541,N_18472);
and U18644 (N_18644,N_18485,N_18409);
or U18645 (N_18645,N_18504,N_18554);
xor U18646 (N_18646,N_18591,N_18586);
nand U18647 (N_18647,N_18503,N_18455);
nand U18648 (N_18648,N_18569,N_18407);
nand U18649 (N_18649,N_18563,N_18560);
xor U18650 (N_18650,N_18458,N_18495);
nand U18651 (N_18651,N_18473,N_18478);
and U18652 (N_18652,N_18491,N_18476);
xnor U18653 (N_18653,N_18580,N_18482);
xnor U18654 (N_18654,N_18568,N_18423);
xnor U18655 (N_18655,N_18415,N_18585);
nor U18656 (N_18656,N_18449,N_18448);
and U18657 (N_18657,N_18512,N_18553);
nand U18658 (N_18658,N_18421,N_18461);
nor U18659 (N_18659,N_18557,N_18474);
and U18660 (N_18660,N_18429,N_18405);
nand U18661 (N_18661,N_18400,N_18497);
or U18662 (N_18662,N_18468,N_18460);
xnor U18663 (N_18663,N_18477,N_18435);
and U18664 (N_18664,N_18574,N_18535);
nor U18665 (N_18665,N_18433,N_18523);
or U18666 (N_18666,N_18579,N_18558);
nand U18667 (N_18667,N_18475,N_18589);
xnor U18668 (N_18668,N_18413,N_18410);
or U18669 (N_18669,N_18488,N_18550);
nand U18670 (N_18670,N_18446,N_18534);
and U18671 (N_18671,N_18436,N_18524);
nand U18672 (N_18672,N_18502,N_18577);
and U18673 (N_18673,N_18501,N_18587);
or U18674 (N_18674,N_18469,N_18597);
nor U18675 (N_18675,N_18418,N_18521);
and U18676 (N_18676,N_18515,N_18479);
and U18677 (N_18677,N_18457,N_18514);
nand U18678 (N_18678,N_18566,N_18459);
or U18679 (N_18679,N_18546,N_18412);
xnor U18680 (N_18680,N_18490,N_18500);
nand U18681 (N_18681,N_18582,N_18424);
nor U18682 (N_18682,N_18451,N_18564);
xnor U18683 (N_18683,N_18489,N_18432);
nand U18684 (N_18684,N_18575,N_18531);
nand U18685 (N_18685,N_18492,N_18463);
and U18686 (N_18686,N_18440,N_18555);
nand U18687 (N_18687,N_18406,N_18583);
nand U18688 (N_18688,N_18428,N_18454);
and U18689 (N_18689,N_18520,N_18510);
nand U18690 (N_18690,N_18549,N_18426);
nand U18691 (N_18691,N_18414,N_18596);
xnor U18692 (N_18692,N_18573,N_18507);
and U18693 (N_18693,N_18572,N_18487);
nand U18694 (N_18694,N_18505,N_18527);
xor U18695 (N_18695,N_18588,N_18552);
nand U18696 (N_18696,N_18530,N_18598);
nand U18697 (N_18697,N_18543,N_18528);
or U18698 (N_18698,N_18584,N_18592);
and U18699 (N_18699,N_18581,N_18519);
or U18700 (N_18700,N_18532,N_18496);
xor U18701 (N_18701,N_18540,N_18573);
or U18702 (N_18702,N_18440,N_18562);
xnor U18703 (N_18703,N_18588,N_18539);
nand U18704 (N_18704,N_18586,N_18517);
xor U18705 (N_18705,N_18540,N_18550);
or U18706 (N_18706,N_18532,N_18583);
and U18707 (N_18707,N_18500,N_18543);
and U18708 (N_18708,N_18509,N_18540);
and U18709 (N_18709,N_18477,N_18524);
and U18710 (N_18710,N_18577,N_18478);
or U18711 (N_18711,N_18446,N_18564);
or U18712 (N_18712,N_18465,N_18412);
and U18713 (N_18713,N_18413,N_18438);
xnor U18714 (N_18714,N_18483,N_18467);
nor U18715 (N_18715,N_18537,N_18489);
or U18716 (N_18716,N_18599,N_18570);
xnor U18717 (N_18717,N_18496,N_18423);
xnor U18718 (N_18718,N_18509,N_18493);
or U18719 (N_18719,N_18531,N_18530);
nand U18720 (N_18720,N_18577,N_18451);
and U18721 (N_18721,N_18437,N_18523);
xor U18722 (N_18722,N_18414,N_18535);
nand U18723 (N_18723,N_18533,N_18438);
nand U18724 (N_18724,N_18501,N_18439);
and U18725 (N_18725,N_18493,N_18516);
and U18726 (N_18726,N_18520,N_18549);
xnor U18727 (N_18727,N_18591,N_18472);
nand U18728 (N_18728,N_18443,N_18405);
and U18729 (N_18729,N_18595,N_18572);
nor U18730 (N_18730,N_18463,N_18472);
nor U18731 (N_18731,N_18467,N_18400);
nor U18732 (N_18732,N_18427,N_18497);
nand U18733 (N_18733,N_18540,N_18419);
xnor U18734 (N_18734,N_18552,N_18506);
xor U18735 (N_18735,N_18531,N_18556);
xnor U18736 (N_18736,N_18504,N_18568);
or U18737 (N_18737,N_18503,N_18558);
nand U18738 (N_18738,N_18501,N_18444);
and U18739 (N_18739,N_18536,N_18437);
nor U18740 (N_18740,N_18476,N_18544);
and U18741 (N_18741,N_18418,N_18500);
or U18742 (N_18742,N_18446,N_18427);
xor U18743 (N_18743,N_18489,N_18414);
xor U18744 (N_18744,N_18530,N_18446);
nor U18745 (N_18745,N_18453,N_18414);
and U18746 (N_18746,N_18576,N_18508);
xnor U18747 (N_18747,N_18499,N_18551);
nor U18748 (N_18748,N_18462,N_18457);
xor U18749 (N_18749,N_18596,N_18586);
and U18750 (N_18750,N_18503,N_18438);
xnor U18751 (N_18751,N_18491,N_18421);
nand U18752 (N_18752,N_18476,N_18527);
xor U18753 (N_18753,N_18431,N_18484);
xnor U18754 (N_18754,N_18503,N_18597);
or U18755 (N_18755,N_18583,N_18490);
nand U18756 (N_18756,N_18541,N_18528);
nand U18757 (N_18757,N_18501,N_18482);
and U18758 (N_18758,N_18548,N_18414);
xor U18759 (N_18759,N_18527,N_18543);
nor U18760 (N_18760,N_18492,N_18576);
nand U18761 (N_18761,N_18428,N_18498);
nand U18762 (N_18762,N_18402,N_18497);
nand U18763 (N_18763,N_18535,N_18482);
xnor U18764 (N_18764,N_18547,N_18537);
nor U18765 (N_18765,N_18427,N_18490);
xnor U18766 (N_18766,N_18447,N_18401);
and U18767 (N_18767,N_18417,N_18430);
or U18768 (N_18768,N_18577,N_18434);
nand U18769 (N_18769,N_18537,N_18589);
xor U18770 (N_18770,N_18417,N_18412);
or U18771 (N_18771,N_18529,N_18427);
nand U18772 (N_18772,N_18426,N_18433);
nor U18773 (N_18773,N_18578,N_18465);
or U18774 (N_18774,N_18554,N_18446);
and U18775 (N_18775,N_18567,N_18576);
or U18776 (N_18776,N_18530,N_18412);
nand U18777 (N_18777,N_18532,N_18436);
and U18778 (N_18778,N_18523,N_18494);
nor U18779 (N_18779,N_18451,N_18587);
xor U18780 (N_18780,N_18449,N_18465);
nand U18781 (N_18781,N_18470,N_18517);
nand U18782 (N_18782,N_18589,N_18492);
xor U18783 (N_18783,N_18436,N_18541);
xor U18784 (N_18784,N_18545,N_18482);
nand U18785 (N_18785,N_18473,N_18484);
xnor U18786 (N_18786,N_18417,N_18531);
or U18787 (N_18787,N_18496,N_18569);
xor U18788 (N_18788,N_18599,N_18536);
nor U18789 (N_18789,N_18527,N_18447);
or U18790 (N_18790,N_18581,N_18555);
or U18791 (N_18791,N_18453,N_18569);
and U18792 (N_18792,N_18527,N_18568);
nand U18793 (N_18793,N_18411,N_18565);
or U18794 (N_18794,N_18585,N_18531);
or U18795 (N_18795,N_18466,N_18529);
nand U18796 (N_18796,N_18514,N_18538);
nand U18797 (N_18797,N_18573,N_18484);
xnor U18798 (N_18798,N_18517,N_18555);
nor U18799 (N_18799,N_18428,N_18438);
nor U18800 (N_18800,N_18732,N_18616);
nor U18801 (N_18801,N_18753,N_18751);
nand U18802 (N_18802,N_18643,N_18782);
nor U18803 (N_18803,N_18705,N_18772);
nor U18804 (N_18804,N_18778,N_18637);
or U18805 (N_18805,N_18608,N_18748);
or U18806 (N_18806,N_18755,N_18634);
xnor U18807 (N_18807,N_18600,N_18791);
or U18808 (N_18808,N_18707,N_18777);
or U18809 (N_18809,N_18613,N_18630);
xor U18810 (N_18810,N_18728,N_18695);
nand U18811 (N_18811,N_18680,N_18696);
and U18812 (N_18812,N_18700,N_18736);
nand U18813 (N_18813,N_18744,N_18617);
nor U18814 (N_18814,N_18684,N_18750);
or U18815 (N_18815,N_18688,N_18653);
xor U18816 (N_18816,N_18789,N_18687);
or U18817 (N_18817,N_18759,N_18620);
and U18818 (N_18818,N_18741,N_18745);
or U18819 (N_18819,N_18636,N_18783);
or U18820 (N_18820,N_18793,N_18664);
and U18821 (N_18821,N_18735,N_18763);
xor U18822 (N_18822,N_18709,N_18683);
nand U18823 (N_18823,N_18762,N_18788);
or U18824 (N_18824,N_18767,N_18747);
nor U18825 (N_18825,N_18639,N_18731);
or U18826 (N_18826,N_18646,N_18628);
xor U18827 (N_18827,N_18773,N_18678);
nor U18828 (N_18828,N_18659,N_18652);
or U18829 (N_18829,N_18623,N_18648);
nor U18830 (N_18830,N_18645,N_18784);
and U18831 (N_18831,N_18656,N_18609);
nor U18832 (N_18832,N_18698,N_18670);
or U18833 (N_18833,N_18692,N_18757);
nor U18834 (N_18834,N_18758,N_18672);
or U18835 (N_18835,N_18701,N_18682);
nor U18836 (N_18836,N_18733,N_18712);
nor U18837 (N_18837,N_18734,N_18714);
and U18838 (N_18838,N_18756,N_18655);
xor U18839 (N_18839,N_18699,N_18702);
nor U18840 (N_18840,N_18726,N_18729);
and U18841 (N_18841,N_18677,N_18671);
and U18842 (N_18842,N_18711,N_18657);
and U18843 (N_18843,N_18704,N_18641);
xor U18844 (N_18844,N_18665,N_18694);
nor U18845 (N_18845,N_18632,N_18681);
nand U18846 (N_18846,N_18754,N_18689);
and U18847 (N_18847,N_18651,N_18764);
nand U18848 (N_18848,N_18765,N_18622);
nor U18849 (N_18849,N_18794,N_18661);
or U18850 (N_18850,N_18724,N_18710);
or U18851 (N_18851,N_18770,N_18673);
or U18852 (N_18852,N_18780,N_18706);
nand U18853 (N_18853,N_18676,N_18727);
xor U18854 (N_18854,N_18739,N_18752);
nor U18855 (N_18855,N_18660,N_18796);
or U18856 (N_18856,N_18766,N_18760);
or U18857 (N_18857,N_18790,N_18693);
nor U18858 (N_18858,N_18740,N_18647);
xor U18859 (N_18859,N_18743,N_18618);
nor U18860 (N_18860,N_18602,N_18685);
xnor U18861 (N_18861,N_18721,N_18662);
xor U18862 (N_18862,N_18742,N_18723);
nand U18863 (N_18863,N_18635,N_18633);
and U18864 (N_18864,N_18638,N_18674);
or U18865 (N_18865,N_18615,N_18654);
or U18866 (N_18866,N_18667,N_18621);
nand U18867 (N_18867,N_18626,N_18775);
and U18868 (N_18868,N_18614,N_18776);
and U18869 (N_18869,N_18658,N_18730);
nor U18870 (N_18870,N_18774,N_18691);
xnor U18871 (N_18871,N_18779,N_18675);
or U18872 (N_18872,N_18605,N_18603);
and U18873 (N_18873,N_18715,N_18619);
or U18874 (N_18874,N_18611,N_18792);
nand U18875 (N_18875,N_18798,N_18781);
or U18876 (N_18876,N_18668,N_18717);
and U18877 (N_18877,N_18703,N_18612);
xnor U18878 (N_18878,N_18746,N_18697);
and U18879 (N_18879,N_18787,N_18624);
and U18880 (N_18880,N_18669,N_18631);
xor U18881 (N_18881,N_18771,N_18690);
nand U18882 (N_18882,N_18708,N_18769);
xnor U18883 (N_18883,N_18761,N_18720);
nand U18884 (N_18884,N_18718,N_18650);
nand U18885 (N_18885,N_18722,N_18716);
and U18886 (N_18886,N_18642,N_18786);
nor U18887 (N_18887,N_18713,N_18640);
nand U18888 (N_18888,N_18644,N_18663);
and U18889 (N_18889,N_18737,N_18749);
nor U18890 (N_18890,N_18629,N_18719);
nand U18891 (N_18891,N_18666,N_18768);
nand U18892 (N_18892,N_18725,N_18797);
or U18893 (N_18893,N_18606,N_18738);
nand U18894 (N_18894,N_18607,N_18610);
nor U18895 (N_18895,N_18686,N_18649);
nand U18896 (N_18896,N_18785,N_18679);
xor U18897 (N_18897,N_18601,N_18799);
nand U18898 (N_18898,N_18604,N_18627);
nor U18899 (N_18899,N_18625,N_18795);
nor U18900 (N_18900,N_18758,N_18743);
and U18901 (N_18901,N_18775,N_18740);
or U18902 (N_18902,N_18607,N_18741);
or U18903 (N_18903,N_18760,N_18795);
nor U18904 (N_18904,N_18675,N_18775);
or U18905 (N_18905,N_18796,N_18619);
nor U18906 (N_18906,N_18689,N_18611);
and U18907 (N_18907,N_18746,N_18757);
or U18908 (N_18908,N_18781,N_18650);
nor U18909 (N_18909,N_18707,N_18608);
and U18910 (N_18910,N_18681,N_18624);
nor U18911 (N_18911,N_18693,N_18670);
nor U18912 (N_18912,N_18626,N_18644);
and U18913 (N_18913,N_18602,N_18670);
xor U18914 (N_18914,N_18762,N_18750);
and U18915 (N_18915,N_18704,N_18749);
or U18916 (N_18916,N_18643,N_18607);
nand U18917 (N_18917,N_18641,N_18735);
nand U18918 (N_18918,N_18760,N_18638);
nand U18919 (N_18919,N_18643,N_18669);
and U18920 (N_18920,N_18672,N_18791);
or U18921 (N_18921,N_18674,N_18637);
xor U18922 (N_18922,N_18689,N_18732);
nand U18923 (N_18923,N_18620,N_18612);
nor U18924 (N_18924,N_18659,N_18775);
xor U18925 (N_18925,N_18671,N_18645);
and U18926 (N_18926,N_18695,N_18735);
nor U18927 (N_18927,N_18644,N_18784);
nand U18928 (N_18928,N_18613,N_18629);
nor U18929 (N_18929,N_18768,N_18758);
xnor U18930 (N_18930,N_18640,N_18754);
and U18931 (N_18931,N_18633,N_18743);
xor U18932 (N_18932,N_18631,N_18693);
xor U18933 (N_18933,N_18771,N_18777);
nor U18934 (N_18934,N_18708,N_18750);
and U18935 (N_18935,N_18609,N_18607);
xnor U18936 (N_18936,N_18649,N_18746);
and U18937 (N_18937,N_18636,N_18685);
nand U18938 (N_18938,N_18721,N_18749);
and U18939 (N_18939,N_18739,N_18612);
nand U18940 (N_18940,N_18657,N_18622);
xnor U18941 (N_18941,N_18687,N_18607);
nand U18942 (N_18942,N_18751,N_18666);
nor U18943 (N_18943,N_18749,N_18621);
nand U18944 (N_18944,N_18702,N_18657);
nand U18945 (N_18945,N_18794,N_18650);
or U18946 (N_18946,N_18784,N_18693);
nand U18947 (N_18947,N_18607,N_18756);
and U18948 (N_18948,N_18717,N_18770);
nand U18949 (N_18949,N_18601,N_18635);
nand U18950 (N_18950,N_18632,N_18721);
nand U18951 (N_18951,N_18636,N_18749);
and U18952 (N_18952,N_18658,N_18755);
or U18953 (N_18953,N_18741,N_18730);
or U18954 (N_18954,N_18727,N_18764);
nand U18955 (N_18955,N_18730,N_18617);
or U18956 (N_18956,N_18668,N_18797);
and U18957 (N_18957,N_18622,N_18757);
and U18958 (N_18958,N_18731,N_18680);
xnor U18959 (N_18959,N_18623,N_18644);
and U18960 (N_18960,N_18744,N_18739);
nand U18961 (N_18961,N_18693,N_18645);
nor U18962 (N_18962,N_18705,N_18652);
xor U18963 (N_18963,N_18777,N_18772);
nor U18964 (N_18964,N_18794,N_18771);
nor U18965 (N_18965,N_18632,N_18658);
xnor U18966 (N_18966,N_18733,N_18675);
and U18967 (N_18967,N_18633,N_18657);
nor U18968 (N_18968,N_18650,N_18761);
or U18969 (N_18969,N_18701,N_18663);
or U18970 (N_18970,N_18748,N_18744);
or U18971 (N_18971,N_18636,N_18673);
nand U18972 (N_18972,N_18752,N_18704);
xor U18973 (N_18973,N_18757,N_18603);
or U18974 (N_18974,N_18750,N_18788);
or U18975 (N_18975,N_18749,N_18603);
nand U18976 (N_18976,N_18607,N_18795);
or U18977 (N_18977,N_18729,N_18755);
nor U18978 (N_18978,N_18630,N_18650);
and U18979 (N_18979,N_18703,N_18765);
xor U18980 (N_18980,N_18667,N_18643);
nor U18981 (N_18981,N_18712,N_18746);
nand U18982 (N_18982,N_18622,N_18646);
nand U18983 (N_18983,N_18624,N_18613);
or U18984 (N_18984,N_18758,N_18696);
and U18985 (N_18985,N_18664,N_18696);
xor U18986 (N_18986,N_18708,N_18747);
and U18987 (N_18987,N_18735,N_18642);
or U18988 (N_18988,N_18765,N_18627);
and U18989 (N_18989,N_18663,N_18607);
or U18990 (N_18990,N_18727,N_18630);
xor U18991 (N_18991,N_18686,N_18622);
or U18992 (N_18992,N_18784,N_18777);
nand U18993 (N_18993,N_18799,N_18618);
nand U18994 (N_18994,N_18703,N_18655);
or U18995 (N_18995,N_18773,N_18748);
nor U18996 (N_18996,N_18796,N_18643);
nand U18997 (N_18997,N_18620,N_18780);
or U18998 (N_18998,N_18704,N_18645);
nand U18999 (N_18999,N_18705,N_18640);
xor U19000 (N_19000,N_18832,N_18869);
and U19001 (N_19001,N_18851,N_18893);
and U19002 (N_19002,N_18899,N_18971);
nor U19003 (N_19003,N_18822,N_18951);
nand U19004 (N_19004,N_18993,N_18942);
xnor U19005 (N_19005,N_18863,N_18818);
or U19006 (N_19006,N_18875,N_18906);
xnor U19007 (N_19007,N_18902,N_18895);
and U19008 (N_19008,N_18932,N_18955);
or U19009 (N_19009,N_18909,N_18918);
nor U19010 (N_19010,N_18961,N_18824);
nand U19011 (N_19011,N_18810,N_18852);
nor U19012 (N_19012,N_18867,N_18920);
nor U19013 (N_19013,N_18897,N_18996);
and U19014 (N_19014,N_18966,N_18845);
nor U19015 (N_19015,N_18854,N_18905);
or U19016 (N_19016,N_18928,N_18913);
nor U19017 (N_19017,N_18935,N_18853);
nor U19018 (N_19018,N_18860,N_18990);
nor U19019 (N_19019,N_18894,N_18983);
nor U19020 (N_19020,N_18844,N_18938);
xnor U19021 (N_19021,N_18956,N_18960);
or U19022 (N_19022,N_18807,N_18915);
nor U19023 (N_19023,N_18922,N_18891);
xnor U19024 (N_19024,N_18884,N_18847);
nand U19025 (N_19025,N_18934,N_18917);
xnor U19026 (N_19026,N_18923,N_18883);
xor U19027 (N_19027,N_18873,N_18911);
nand U19028 (N_19028,N_18892,N_18819);
or U19029 (N_19029,N_18858,N_18953);
nor U19030 (N_19030,N_18820,N_18840);
or U19031 (N_19031,N_18944,N_18937);
nand U19032 (N_19032,N_18825,N_18912);
nor U19033 (N_19033,N_18806,N_18963);
xnor U19034 (N_19034,N_18994,N_18921);
and U19035 (N_19035,N_18805,N_18919);
and U19036 (N_19036,N_18855,N_18871);
nand U19037 (N_19037,N_18866,N_18817);
nor U19038 (N_19038,N_18856,N_18811);
nand U19039 (N_19039,N_18801,N_18927);
or U19040 (N_19040,N_18815,N_18870);
or U19041 (N_19041,N_18859,N_18988);
or U19042 (N_19042,N_18992,N_18826);
and U19043 (N_19043,N_18835,N_18833);
or U19044 (N_19044,N_18984,N_18809);
xnor U19045 (N_19045,N_18903,N_18967);
and U19046 (N_19046,N_18802,N_18874);
or U19047 (N_19047,N_18837,N_18940);
nand U19048 (N_19048,N_18986,N_18958);
or U19049 (N_19049,N_18916,N_18901);
nand U19050 (N_19050,N_18885,N_18970);
nand U19051 (N_19051,N_18933,N_18957);
nor U19052 (N_19052,N_18804,N_18925);
xnor U19053 (N_19053,N_18991,N_18949);
or U19054 (N_19054,N_18989,N_18943);
and U19055 (N_19055,N_18841,N_18827);
and U19056 (N_19056,N_18836,N_18800);
and U19057 (N_19057,N_18981,N_18979);
xor U19058 (N_19058,N_18864,N_18877);
xor U19059 (N_19059,N_18982,N_18872);
or U19060 (N_19060,N_18977,N_18904);
xor U19061 (N_19061,N_18931,N_18812);
nand U19062 (N_19062,N_18946,N_18985);
xor U19063 (N_19063,N_18881,N_18876);
xor U19064 (N_19064,N_18834,N_18887);
xnor U19065 (N_19065,N_18980,N_18965);
nand U19066 (N_19066,N_18936,N_18898);
xor U19067 (N_19067,N_18964,N_18974);
or U19068 (N_19068,N_18839,N_18828);
nor U19069 (N_19069,N_18850,N_18830);
xor U19070 (N_19070,N_18908,N_18890);
nand U19071 (N_19071,N_18880,N_18808);
nand U19072 (N_19072,N_18952,N_18846);
xnor U19073 (N_19073,N_18865,N_18862);
nor U19074 (N_19074,N_18997,N_18995);
or U19075 (N_19075,N_18941,N_18914);
nand U19076 (N_19076,N_18842,N_18907);
nor U19077 (N_19077,N_18930,N_18948);
and U19078 (N_19078,N_18816,N_18972);
xnor U19079 (N_19079,N_18987,N_18889);
nor U19080 (N_19080,N_18803,N_18947);
or U19081 (N_19081,N_18962,N_18831);
and U19082 (N_19082,N_18857,N_18813);
and U19083 (N_19083,N_18969,N_18926);
nand U19084 (N_19084,N_18945,N_18882);
nand U19085 (N_19085,N_18878,N_18968);
nand U19086 (N_19086,N_18924,N_18896);
nand U19087 (N_19087,N_18848,N_18849);
nor U19088 (N_19088,N_18999,N_18959);
and U19089 (N_19089,N_18829,N_18823);
nor U19090 (N_19090,N_18843,N_18998);
or U19091 (N_19091,N_18978,N_18975);
and U19092 (N_19092,N_18886,N_18868);
nand U19093 (N_19093,N_18973,N_18888);
nand U19094 (N_19094,N_18954,N_18838);
xor U19095 (N_19095,N_18900,N_18879);
or U19096 (N_19096,N_18910,N_18929);
or U19097 (N_19097,N_18861,N_18950);
or U19098 (N_19098,N_18821,N_18939);
or U19099 (N_19099,N_18976,N_18814);
and U19100 (N_19100,N_18956,N_18935);
and U19101 (N_19101,N_18861,N_18976);
xnor U19102 (N_19102,N_18831,N_18855);
and U19103 (N_19103,N_18847,N_18987);
or U19104 (N_19104,N_18861,N_18866);
nand U19105 (N_19105,N_18969,N_18877);
nand U19106 (N_19106,N_18813,N_18923);
nor U19107 (N_19107,N_18895,N_18986);
nand U19108 (N_19108,N_18838,N_18817);
xor U19109 (N_19109,N_18888,N_18813);
and U19110 (N_19110,N_18972,N_18822);
or U19111 (N_19111,N_18928,N_18924);
nor U19112 (N_19112,N_18943,N_18962);
nand U19113 (N_19113,N_18825,N_18965);
nand U19114 (N_19114,N_18972,N_18940);
or U19115 (N_19115,N_18903,N_18955);
nor U19116 (N_19116,N_18888,N_18876);
and U19117 (N_19117,N_18967,N_18961);
xor U19118 (N_19118,N_18855,N_18927);
nand U19119 (N_19119,N_18900,N_18856);
and U19120 (N_19120,N_18811,N_18940);
and U19121 (N_19121,N_18870,N_18915);
xor U19122 (N_19122,N_18851,N_18875);
nor U19123 (N_19123,N_18875,N_18959);
nor U19124 (N_19124,N_18970,N_18977);
or U19125 (N_19125,N_18862,N_18883);
or U19126 (N_19126,N_18847,N_18994);
nand U19127 (N_19127,N_18930,N_18860);
and U19128 (N_19128,N_18900,N_18907);
xnor U19129 (N_19129,N_18892,N_18953);
xor U19130 (N_19130,N_18840,N_18898);
and U19131 (N_19131,N_18933,N_18804);
nor U19132 (N_19132,N_18957,N_18802);
nand U19133 (N_19133,N_18916,N_18841);
nor U19134 (N_19134,N_18940,N_18899);
and U19135 (N_19135,N_18996,N_18953);
nand U19136 (N_19136,N_18817,N_18991);
xnor U19137 (N_19137,N_18959,N_18939);
and U19138 (N_19138,N_18861,N_18911);
nor U19139 (N_19139,N_18960,N_18921);
xnor U19140 (N_19140,N_18816,N_18903);
or U19141 (N_19141,N_18936,N_18924);
and U19142 (N_19142,N_18813,N_18802);
nand U19143 (N_19143,N_18950,N_18966);
nor U19144 (N_19144,N_18948,N_18831);
nor U19145 (N_19145,N_18865,N_18890);
xnor U19146 (N_19146,N_18949,N_18854);
nand U19147 (N_19147,N_18914,N_18915);
xnor U19148 (N_19148,N_18817,N_18855);
nand U19149 (N_19149,N_18980,N_18974);
xnor U19150 (N_19150,N_18838,N_18952);
and U19151 (N_19151,N_18893,N_18889);
nand U19152 (N_19152,N_18847,N_18861);
or U19153 (N_19153,N_18828,N_18859);
xor U19154 (N_19154,N_18966,N_18941);
nor U19155 (N_19155,N_18991,N_18935);
nand U19156 (N_19156,N_18807,N_18902);
nand U19157 (N_19157,N_18953,N_18844);
and U19158 (N_19158,N_18893,N_18844);
and U19159 (N_19159,N_18888,N_18804);
or U19160 (N_19160,N_18929,N_18942);
or U19161 (N_19161,N_18928,N_18863);
xor U19162 (N_19162,N_18997,N_18834);
xnor U19163 (N_19163,N_18925,N_18984);
xor U19164 (N_19164,N_18840,N_18905);
and U19165 (N_19165,N_18950,N_18959);
or U19166 (N_19166,N_18929,N_18919);
and U19167 (N_19167,N_18886,N_18888);
xor U19168 (N_19168,N_18850,N_18973);
and U19169 (N_19169,N_18827,N_18839);
nor U19170 (N_19170,N_18908,N_18877);
nor U19171 (N_19171,N_18965,N_18848);
or U19172 (N_19172,N_18819,N_18810);
xnor U19173 (N_19173,N_18959,N_18809);
nor U19174 (N_19174,N_18886,N_18883);
xnor U19175 (N_19175,N_18934,N_18986);
xnor U19176 (N_19176,N_18870,N_18806);
xor U19177 (N_19177,N_18892,N_18960);
nand U19178 (N_19178,N_18871,N_18877);
nand U19179 (N_19179,N_18933,N_18888);
nor U19180 (N_19180,N_18940,N_18948);
xor U19181 (N_19181,N_18843,N_18932);
nor U19182 (N_19182,N_18965,N_18838);
nand U19183 (N_19183,N_18860,N_18931);
and U19184 (N_19184,N_18897,N_18802);
nand U19185 (N_19185,N_18976,N_18995);
or U19186 (N_19186,N_18857,N_18896);
nor U19187 (N_19187,N_18939,N_18998);
xnor U19188 (N_19188,N_18918,N_18944);
nor U19189 (N_19189,N_18853,N_18868);
xnor U19190 (N_19190,N_18930,N_18896);
nand U19191 (N_19191,N_18896,N_18964);
nand U19192 (N_19192,N_18925,N_18975);
xor U19193 (N_19193,N_18919,N_18822);
or U19194 (N_19194,N_18884,N_18915);
nor U19195 (N_19195,N_18883,N_18967);
xnor U19196 (N_19196,N_18837,N_18927);
and U19197 (N_19197,N_18965,N_18992);
xnor U19198 (N_19198,N_18897,N_18857);
nor U19199 (N_19199,N_18875,N_18957);
and U19200 (N_19200,N_19084,N_19137);
nor U19201 (N_19201,N_19007,N_19072);
nor U19202 (N_19202,N_19033,N_19188);
xnor U19203 (N_19203,N_19161,N_19189);
or U19204 (N_19204,N_19143,N_19014);
nand U19205 (N_19205,N_19070,N_19095);
nor U19206 (N_19206,N_19107,N_19015);
nor U19207 (N_19207,N_19063,N_19067);
nand U19208 (N_19208,N_19083,N_19085);
or U19209 (N_19209,N_19100,N_19048);
nand U19210 (N_19210,N_19088,N_19090);
and U19211 (N_19211,N_19196,N_19087);
and U19212 (N_19212,N_19195,N_19108);
xnor U19213 (N_19213,N_19191,N_19180);
and U19214 (N_19214,N_19086,N_19153);
and U19215 (N_19215,N_19016,N_19022);
nor U19216 (N_19216,N_19064,N_19120);
or U19217 (N_19217,N_19165,N_19110);
or U19218 (N_19218,N_19045,N_19093);
nor U19219 (N_19219,N_19124,N_19020);
or U19220 (N_19220,N_19010,N_19071);
nor U19221 (N_19221,N_19183,N_19027);
nand U19222 (N_19222,N_19044,N_19170);
xnor U19223 (N_19223,N_19029,N_19163);
and U19224 (N_19224,N_19035,N_19121);
or U19225 (N_19225,N_19198,N_19006);
nand U19226 (N_19226,N_19129,N_19103);
nand U19227 (N_19227,N_19102,N_19004);
xnor U19228 (N_19228,N_19173,N_19075);
nor U19229 (N_19229,N_19089,N_19178);
and U19230 (N_19230,N_19054,N_19190);
xnor U19231 (N_19231,N_19098,N_19028);
or U19232 (N_19232,N_19078,N_19026);
nand U19233 (N_19233,N_19032,N_19148);
xnor U19234 (N_19234,N_19140,N_19001);
and U19235 (N_19235,N_19167,N_19128);
or U19236 (N_19236,N_19145,N_19080);
or U19237 (N_19237,N_19159,N_19142);
nor U19238 (N_19238,N_19116,N_19122);
nor U19239 (N_19239,N_19031,N_19117);
xnor U19240 (N_19240,N_19123,N_19050);
nor U19241 (N_19241,N_19130,N_19105);
xnor U19242 (N_19242,N_19176,N_19036);
nor U19243 (N_19243,N_19009,N_19127);
nor U19244 (N_19244,N_19179,N_19030);
and U19245 (N_19245,N_19039,N_19019);
nand U19246 (N_19246,N_19096,N_19109);
nand U19247 (N_19247,N_19082,N_19000);
or U19248 (N_19248,N_19125,N_19194);
or U19249 (N_19249,N_19181,N_19150);
and U19250 (N_19250,N_19040,N_19059);
and U19251 (N_19251,N_19113,N_19132);
or U19252 (N_19252,N_19034,N_19172);
and U19253 (N_19253,N_19185,N_19136);
xor U19254 (N_19254,N_19043,N_19164);
nand U19255 (N_19255,N_19073,N_19002);
nor U19256 (N_19256,N_19152,N_19154);
xor U19257 (N_19257,N_19158,N_19079);
xor U19258 (N_19258,N_19193,N_19101);
and U19259 (N_19259,N_19046,N_19023);
or U19260 (N_19260,N_19038,N_19119);
nor U19261 (N_19261,N_19091,N_19138);
and U19262 (N_19262,N_19062,N_19131);
nor U19263 (N_19263,N_19133,N_19174);
and U19264 (N_19264,N_19012,N_19135);
or U19265 (N_19265,N_19076,N_19057);
nand U19266 (N_19266,N_19011,N_19114);
or U19267 (N_19267,N_19017,N_19134);
nor U19268 (N_19268,N_19092,N_19041);
nand U19269 (N_19269,N_19005,N_19175);
or U19270 (N_19270,N_19097,N_19192);
or U19271 (N_19271,N_19171,N_19018);
and U19272 (N_19272,N_19066,N_19106);
nor U19273 (N_19273,N_19169,N_19042);
nor U19274 (N_19274,N_19149,N_19141);
nor U19275 (N_19275,N_19187,N_19024);
nor U19276 (N_19276,N_19013,N_19157);
or U19277 (N_19277,N_19168,N_19146);
and U19278 (N_19278,N_19126,N_19025);
and U19279 (N_19279,N_19051,N_19037);
nand U19280 (N_19280,N_19052,N_19094);
nand U19281 (N_19281,N_19184,N_19155);
nand U19282 (N_19282,N_19104,N_19053);
xor U19283 (N_19283,N_19160,N_19177);
and U19284 (N_19284,N_19021,N_19112);
xnor U19285 (N_19285,N_19069,N_19139);
and U19286 (N_19286,N_19055,N_19162);
or U19287 (N_19287,N_19074,N_19197);
nor U19288 (N_19288,N_19199,N_19060);
and U19289 (N_19289,N_19008,N_19056);
xnor U19290 (N_19290,N_19099,N_19077);
and U19291 (N_19291,N_19049,N_19156);
nand U19292 (N_19292,N_19111,N_19166);
nor U19293 (N_19293,N_19151,N_19003);
xor U19294 (N_19294,N_19144,N_19182);
and U19295 (N_19295,N_19047,N_19147);
nand U19296 (N_19296,N_19115,N_19058);
nor U19297 (N_19297,N_19065,N_19068);
nor U19298 (N_19298,N_19081,N_19118);
or U19299 (N_19299,N_19186,N_19061);
nand U19300 (N_19300,N_19076,N_19188);
or U19301 (N_19301,N_19188,N_19065);
nor U19302 (N_19302,N_19032,N_19070);
nand U19303 (N_19303,N_19045,N_19100);
or U19304 (N_19304,N_19010,N_19021);
and U19305 (N_19305,N_19015,N_19066);
nand U19306 (N_19306,N_19040,N_19099);
or U19307 (N_19307,N_19122,N_19123);
nor U19308 (N_19308,N_19123,N_19000);
xnor U19309 (N_19309,N_19101,N_19097);
xor U19310 (N_19310,N_19065,N_19005);
nand U19311 (N_19311,N_19171,N_19060);
and U19312 (N_19312,N_19013,N_19155);
nand U19313 (N_19313,N_19037,N_19077);
and U19314 (N_19314,N_19039,N_19122);
and U19315 (N_19315,N_19108,N_19192);
xor U19316 (N_19316,N_19008,N_19078);
xor U19317 (N_19317,N_19194,N_19067);
or U19318 (N_19318,N_19114,N_19041);
and U19319 (N_19319,N_19006,N_19109);
nor U19320 (N_19320,N_19094,N_19167);
xnor U19321 (N_19321,N_19197,N_19130);
and U19322 (N_19322,N_19162,N_19097);
or U19323 (N_19323,N_19082,N_19027);
nor U19324 (N_19324,N_19199,N_19147);
nand U19325 (N_19325,N_19007,N_19129);
or U19326 (N_19326,N_19052,N_19179);
nor U19327 (N_19327,N_19098,N_19113);
nand U19328 (N_19328,N_19057,N_19158);
or U19329 (N_19329,N_19016,N_19127);
xor U19330 (N_19330,N_19086,N_19191);
nor U19331 (N_19331,N_19088,N_19009);
nor U19332 (N_19332,N_19188,N_19167);
xor U19333 (N_19333,N_19071,N_19150);
nor U19334 (N_19334,N_19006,N_19038);
or U19335 (N_19335,N_19033,N_19030);
and U19336 (N_19336,N_19132,N_19126);
xor U19337 (N_19337,N_19070,N_19015);
xnor U19338 (N_19338,N_19179,N_19071);
and U19339 (N_19339,N_19102,N_19021);
and U19340 (N_19340,N_19072,N_19039);
nor U19341 (N_19341,N_19092,N_19194);
nor U19342 (N_19342,N_19018,N_19065);
and U19343 (N_19343,N_19087,N_19190);
xor U19344 (N_19344,N_19137,N_19181);
or U19345 (N_19345,N_19187,N_19137);
or U19346 (N_19346,N_19021,N_19030);
xor U19347 (N_19347,N_19129,N_19060);
nand U19348 (N_19348,N_19056,N_19045);
and U19349 (N_19349,N_19057,N_19154);
nor U19350 (N_19350,N_19078,N_19151);
and U19351 (N_19351,N_19090,N_19054);
and U19352 (N_19352,N_19027,N_19004);
or U19353 (N_19353,N_19154,N_19096);
nand U19354 (N_19354,N_19086,N_19116);
or U19355 (N_19355,N_19028,N_19123);
xor U19356 (N_19356,N_19061,N_19131);
nor U19357 (N_19357,N_19004,N_19091);
xor U19358 (N_19358,N_19021,N_19065);
nor U19359 (N_19359,N_19129,N_19119);
and U19360 (N_19360,N_19057,N_19172);
nand U19361 (N_19361,N_19054,N_19115);
and U19362 (N_19362,N_19007,N_19021);
nand U19363 (N_19363,N_19127,N_19110);
nand U19364 (N_19364,N_19061,N_19005);
xnor U19365 (N_19365,N_19012,N_19118);
nand U19366 (N_19366,N_19096,N_19075);
and U19367 (N_19367,N_19162,N_19124);
or U19368 (N_19368,N_19129,N_19123);
nor U19369 (N_19369,N_19115,N_19128);
nand U19370 (N_19370,N_19115,N_19031);
xnor U19371 (N_19371,N_19035,N_19075);
or U19372 (N_19372,N_19092,N_19170);
or U19373 (N_19373,N_19102,N_19180);
xnor U19374 (N_19374,N_19129,N_19145);
xor U19375 (N_19375,N_19162,N_19175);
and U19376 (N_19376,N_19056,N_19070);
nand U19377 (N_19377,N_19183,N_19157);
nand U19378 (N_19378,N_19100,N_19022);
nor U19379 (N_19379,N_19195,N_19098);
and U19380 (N_19380,N_19122,N_19194);
xor U19381 (N_19381,N_19060,N_19066);
and U19382 (N_19382,N_19086,N_19105);
and U19383 (N_19383,N_19010,N_19120);
nand U19384 (N_19384,N_19168,N_19135);
and U19385 (N_19385,N_19134,N_19158);
nor U19386 (N_19386,N_19087,N_19070);
nand U19387 (N_19387,N_19154,N_19108);
nor U19388 (N_19388,N_19184,N_19000);
nor U19389 (N_19389,N_19054,N_19163);
xnor U19390 (N_19390,N_19037,N_19078);
and U19391 (N_19391,N_19154,N_19053);
nor U19392 (N_19392,N_19033,N_19090);
nor U19393 (N_19393,N_19081,N_19151);
nand U19394 (N_19394,N_19073,N_19045);
and U19395 (N_19395,N_19104,N_19045);
nand U19396 (N_19396,N_19057,N_19128);
nand U19397 (N_19397,N_19067,N_19172);
nor U19398 (N_19398,N_19115,N_19139);
nor U19399 (N_19399,N_19088,N_19033);
or U19400 (N_19400,N_19384,N_19237);
and U19401 (N_19401,N_19214,N_19376);
nor U19402 (N_19402,N_19238,N_19329);
xor U19403 (N_19403,N_19322,N_19358);
xor U19404 (N_19404,N_19388,N_19389);
nand U19405 (N_19405,N_19328,N_19293);
and U19406 (N_19406,N_19263,N_19259);
nand U19407 (N_19407,N_19352,N_19220);
xnor U19408 (N_19408,N_19399,N_19209);
nand U19409 (N_19409,N_19251,N_19223);
and U19410 (N_19410,N_19337,N_19225);
nor U19411 (N_19411,N_19202,N_19260);
or U19412 (N_19412,N_19262,N_19326);
and U19413 (N_19413,N_19341,N_19249);
nor U19414 (N_19414,N_19299,N_19362);
or U19415 (N_19415,N_19386,N_19394);
xor U19416 (N_19416,N_19374,N_19216);
and U19417 (N_19417,N_19321,N_19372);
or U19418 (N_19418,N_19242,N_19219);
nand U19419 (N_19419,N_19235,N_19305);
or U19420 (N_19420,N_19272,N_19343);
or U19421 (N_19421,N_19391,N_19256);
xnor U19422 (N_19422,N_19271,N_19266);
and U19423 (N_19423,N_19356,N_19330);
nor U19424 (N_19424,N_19303,N_19261);
and U19425 (N_19425,N_19312,N_19240);
and U19426 (N_19426,N_19387,N_19208);
or U19427 (N_19427,N_19215,N_19311);
or U19428 (N_19428,N_19254,N_19340);
and U19429 (N_19429,N_19335,N_19276);
xor U19430 (N_19430,N_19331,N_19232);
and U19431 (N_19431,N_19357,N_19230);
and U19432 (N_19432,N_19281,N_19346);
and U19433 (N_19433,N_19309,N_19245);
nand U19434 (N_19434,N_19284,N_19307);
nand U19435 (N_19435,N_19333,N_19236);
nor U19436 (N_19436,N_19393,N_19224);
xnor U19437 (N_19437,N_19353,N_19246);
nor U19438 (N_19438,N_19258,N_19205);
or U19439 (N_19439,N_19213,N_19228);
and U19440 (N_19440,N_19318,N_19222);
nor U19441 (N_19441,N_19257,N_19278);
and U19442 (N_19442,N_19368,N_19392);
and U19443 (N_19443,N_19347,N_19348);
xnor U19444 (N_19444,N_19227,N_19378);
nor U19445 (N_19445,N_19339,N_19306);
xor U19446 (N_19446,N_19390,N_19360);
xor U19447 (N_19447,N_19325,N_19320);
and U19448 (N_19448,N_19231,N_19200);
nand U19449 (N_19449,N_19201,N_19300);
nor U19450 (N_19450,N_19323,N_19267);
nor U19451 (N_19451,N_19313,N_19302);
xnor U19452 (N_19452,N_19233,N_19319);
nor U19453 (N_19453,N_19212,N_19285);
and U19454 (N_19454,N_19297,N_19204);
nor U19455 (N_19455,N_19274,N_19275);
xor U19456 (N_19456,N_19317,N_19345);
and U19457 (N_19457,N_19277,N_19290);
and U19458 (N_19458,N_19367,N_19255);
and U19459 (N_19459,N_19273,N_19316);
xnor U19460 (N_19460,N_19369,N_19379);
nor U19461 (N_19461,N_19380,N_19396);
or U19462 (N_19462,N_19289,N_19286);
or U19463 (N_19463,N_19265,N_19247);
nor U19464 (N_19464,N_19203,N_19253);
or U19465 (N_19465,N_19308,N_19243);
and U19466 (N_19466,N_19366,N_19226);
xor U19467 (N_19467,N_19398,N_19363);
nor U19468 (N_19468,N_19383,N_19332);
or U19469 (N_19469,N_19234,N_19291);
or U19470 (N_19470,N_19295,N_19324);
nor U19471 (N_19471,N_19351,N_19244);
nor U19472 (N_19472,N_19395,N_19211);
or U19473 (N_19473,N_19252,N_19314);
nand U19474 (N_19474,N_19248,N_19221);
nor U19475 (N_19475,N_19250,N_19292);
xnor U19476 (N_19476,N_19382,N_19371);
nor U19477 (N_19477,N_19349,N_19241);
and U19478 (N_19478,N_19282,N_19218);
xnor U19479 (N_19479,N_19361,N_19350);
nor U19480 (N_19480,N_19355,N_19359);
and U19481 (N_19481,N_19397,N_19210);
xor U19482 (N_19482,N_19229,N_19375);
or U19483 (N_19483,N_19294,N_19364);
nor U19484 (N_19484,N_19370,N_19298);
nor U19485 (N_19485,N_19365,N_19310);
and U19486 (N_19486,N_19338,N_19334);
and U19487 (N_19487,N_19279,N_19207);
nand U19488 (N_19488,N_19296,N_19385);
nand U19489 (N_19489,N_19264,N_19288);
or U19490 (N_19490,N_19217,N_19344);
nor U19491 (N_19491,N_19287,N_19280);
xor U19492 (N_19492,N_19336,N_19304);
nor U19493 (N_19493,N_19283,N_19381);
and U19494 (N_19494,N_19377,N_19269);
nand U19495 (N_19495,N_19268,N_19354);
and U19496 (N_19496,N_19342,N_19315);
xnor U19497 (N_19497,N_19270,N_19327);
nand U19498 (N_19498,N_19301,N_19239);
and U19499 (N_19499,N_19206,N_19373);
or U19500 (N_19500,N_19273,N_19208);
and U19501 (N_19501,N_19355,N_19327);
nand U19502 (N_19502,N_19274,N_19231);
nand U19503 (N_19503,N_19236,N_19312);
and U19504 (N_19504,N_19254,N_19266);
nand U19505 (N_19505,N_19290,N_19322);
or U19506 (N_19506,N_19313,N_19319);
and U19507 (N_19507,N_19252,N_19379);
xnor U19508 (N_19508,N_19334,N_19272);
and U19509 (N_19509,N_19282,N_19328);
nand U19510 (N_19510,N_19238,N_19213);
nor U19511 (N_19511,N_19283,N_19212);
xor U19512 (N_19512,N_19259,N_19273);
or U19513 (N_19513,N_19283,N_19282);
nand U19514 (N_19514,N_19261,N_19243);
nor U19515 (N_19515,N_19200,N_19320);
or U19516 (N_19516,N_19259,N_19213);
or U19517 (N_19517,N_19369,N_19316);
or U19518 (N_19518,N_19384,N_19286);
or U19519 (N_19519,N_19352,N_19362);
and U19520 (N_19520,N_19315,N_19216);
nor U19521 (N_19521,N_19297,N_19313);
nor U19522 (N_19522,N_19350,N_19280);
nand U19523 (N_19523,N_19318,N_19352);
xor U19524 (N_19524,N_19211,N_19355);
or U19525 (N_19525,N_19236,N_19269);
nor U19526 (N_19526,N_19211,N_19307);
or U19527 (N_19527,N_19275,N_19278);
xor U19528 (N_19528,N_19346,N_19387);
nand U19529 (N_19529,N_19229,N_19238);
nor U19530 (N_19530,N_19310,N_19312);
and U19531 (N_19531,N_19321,N_19229);
and U19532 (N_19532,N_19252,N_19241);
nand U19533 (N_19533,N_19299,N_19336);
nor U19534 (N_19534,N_19313,N_19353);
or U19535 (N_19535,N_19248,N_19272);
or U19536 (N_19536,N_19376,N_19318);
xnor U19537 (N_19537,N_19352,N_19382);
nand U19538 (N_19538,N_19363,N_19242);
or U19539 (N_19539,N_19348,N_19224);
nand U19540 (N_19540,N_19240,N_19394);
xnor U19541 (N_19541,N_19376,N_19252);
and U19542 (N_19542,N_19236,N_19314);
xnor U19543 (N_19543,N_19276,N_19256);
and U19544 (N_19544,N_19324,N_19391);
xnor U19545 (N_19545,N_19360,N_19200);
xor U19546 (N_19546,N_19254,N_19358);
or U19547 (N_19547,N_19224,N_19342);
xnor U19548 (N_19548,N_19395,N_19345);
or U19549 (N_19549,N_19238,N_19325);
and U19550 (N_19550,N_19201,N_19253);
xnor U19551 (N_19551,N_19279,N_19301);
nor U19552 (N_19552,N_19294,N_19277);
and U19553 (N_19553,N_19348,N_19304);
and U19554 (N_19554,N_19289,N_19353);
xor U19555 (N_19555,N_19359,N_19285);
nor U19556 (N_19556,N_19331,N_19236);
nand U19557 (N_19557,N_19385,N_19212);
nand U19558 (N_19558,N_19270,N_19396);
and U19559 (N_19559,N_19287,N_19300);
and U19560 (N_19560,N_19380,N_19388);
nor U19561 (N_19561,N_19368,N_19285);
nand U19562 (N_19562,N_19228,N_19381);
nand U19563 (N_19563,N_19327,N_19295);
nand U19564 (N_19564,N_19385,N_19285);
xnor U19565 (N_19565,N_19289,N_19347);
or U19566 (N_19566,N_19296,N_19300);
and U19567 (N_19567,N_19288,N_19306);
and U19568 (N_19568,N_19228,N_19254);
xnor U19569 (N_19569,N_19349,N_19314);
nor U19570 (N_19570,N_19267,N_19284);
or U19571 (N_19571,N_19371,N_19396);
and U19572 (N_19572,N_19306,N_19284);
xor U19573 (N_19573,N_19365,N_19260);
nand U19574 (N_19574,N_19219,N_19203);
nand U19575 (N_19575,N_19331,N_19229);
xor U19576 (N_19576,N_19333,N_19277);
xnor U19577 (N_19577,N_19357,N_19309);
xnor U19578 (N_19578,N_19390,N_19309);
nand U19579 (N_19579,N_19338,N_19275);
and U19580 (N_19580,N_19248,N_19349);
xor U19581 (N_19581,N_19335,N_19212);
or U19582 (N_19582,N_19392,N_19247);
nand U19583 (N_19583,N_19340,N_19258);
nor U19584 (N_19584,N_19250,N_19269);
xnor U19585 (N_19585,N_19221,N_19293);
xnor U19586 (N_19586,N_19355,N_19292);
nand U19587 (N_19587,N_19396,N_19334);
or U19588 (N_19588,N_19301,N_19247);
xor U19589 (N_19589,N_19381,N_19394);
nor U19590 (N_19590,N_19377,N_19320);
or U19591 (N_19591,N_19245,N_19217);
xor U19592 (N_19592,N_19313,N_19383);
and U19593 (N_19593,N_19367,N_19394);
nand U19594 (N_19594,N_19209,N_19245);
xor U19595 (N_19595,N_19251,N_19379);
nor U19596 (N_19596,N_19322,N_19361);
nor U19597 (N_19597,N_19228,N_19210);
or U19598 (N_19598,N_19327,N_19308);
nor U19599 (N_19599,N_19352,N_19296);
or U19600 (N_19600,N_19419,N_19460);
nand U19601 (N_19601,N_19503,N_19550);
or U19602 (N_19602,N_19484,N_19496);
xnor U19603 (N_19603,N_19507,N_19546);
nor U19604 (N_19604,N_19434,N_19429);
nor U19605 (N_19605,N_19476,N_19539);
nand U19606 (N_19606,N_19424,N_19598);
and U19607 (N_19607,N_19459,N_19464);
nor U19608 (N_19608,N_19401,N_19482);
nand U19609 (N_19609,N_19443,N_19588);
xnor U19610 (N_19610,N_19495,N_19566);
nor U19611 (N_19611,N_19409,N_19447);
nand U19612 (N_19612,N_19491,N_19540);
or U19613 (N_19613,N_19557,N_19551);
and U19614 (N_19614,N_19508,N_19417);
nand U19615 (N_19615,N_19572,N_19514);
nor U19616 (N_19616,N_19414,N_19579);
and U19617 (N_19617,N_19560,N_19400);
xnor U19618 (N_19618,N_19524,N_19472);
nand U19619 (N_19619,N_19585,N_19559);
and U19620 (N_19620,N_19450,N_19488);
nand U19621 (N_19621,N_19578,N_19543);
nand U19622 (N_19622,N_19549,N_19473);
xor U19623 (N_19623,N_19413,N_19519);
xor U19624 (N_19624,N_19527,N_19467);
and U19625 (N_19625,N_19465,N_19510);
or U19626 (N_19626,N_19475,N_19437);
nand U19627 (N_19627,N_19581,N_19574);
or U19628 (N_19628,N_19497,N_19517);
nand U19629 (N_19629,N_19405,N_19421);
nand U19630 (N_19630,N_19536,N_19534);
nand U19631 (N_19631,N_19458,N_19478);
and U19632 (N_19632,N_19480,N_19509);
or U19633 (N_19633,N_19529,N_19569);
and U19634 (N_19634,N_19556,N_19580);
and U19635 (N_19635,N_19532,N_19483);
nor U19636 (N_19636,N_19455,N_19403);
nand U19637 (N_19637,N_19561,N_19404);
nand U19638 (N_19638,N_19470,N_19412);
and U19639 (N_19639,N_19541,N_19555);
nand U19640 (N_19640,N_19592,N_19521);
and U19641 (N_19641,N_19596,N_19451);
nor U19642 (N_19642,N_19554,N_19594);
xor U19643 (N_19643,N_19542,N_19586);
or U19644 (N_19644,N_19501,N_19474);
and U19645 (N_19645,N_19548,N_19446);
xor U19646 (N_19646,N_19430,N_19498);
xnor U19647 (N_19647,N_19492,N_19528);
nor U19648 (N_19648,N_19454,N_19530);
or U19649 (N_19649,N_19444,N_19456);
or U19650 (N_19650,N_19563,N_19570);
and U19651 (N_19651,N_19442,N_19425);
or U19652 (N_19652,N_19547,N_19573);
or U19653 (N_19653,N_19471,N_19537);
and U19654 (N_19654,N_19564,N_19433);
xnor U19655 (N_19655,N_19562,N_19558);
nand U19656 (N_19656,N_19411,N_19408);
and U19657 (N_19657,N_19435,N_19533);
xnor U19658 (N_19658,N_19552,N_19591);
and U19659 (N_19659,N_19597,N_19441);
xnor U19660 (N_19660,N_19577,N_19440);
nor U19661 (N_19661,N_19506,N_19479);
or U19662 (N_19662,N_19439,N_19595);
xnor U19663 (N_19663,N_19576,N_19553);
and U19664 (N_19664,N_19448,N_19516);
and U19665 (N_19665,N_19410,N_19452);
xor U19666 (N_19666,N_19599,N_19489);
xnor U19667 (N_19667,N_19449,N_19583);
nand U19668 (N_19668,N_19406,N_19518);
nor U19669 (N_19669,N_19526,N_19582);
and U19670 (N_19670,N_19571,N_19453);
and U19671 (N_19671,N_19587,N_19584);
nand U19672 (N_19672,N_19502,N_19485);
nor U19673 (N_19673,N_19462,N_19477);
or U19674 (N_19674,N_19565,N_19481);
and U19675 (N_19675,N_19538,N_19487);
nand U19676 (N_19676,N_19522,N_19428);
xor U19677 (N_19677,N_19545,N_19494);
nor U19678 (N_19678,N_19525,N_19515);
nand U19679 (N_19679,N_19589,N_19427);
nor U19680 (N_19680,N_19513,N_19415);
xor U19681 (N_19681,N_19422,N_19457);
xor U19682 (N_19682,N_19407,N_19436);
nor U19683 (N_19683,N_19493,N_19431);
or U19684 (N_19684,N_19432,N_19511);
and U19685 (N_19685,N_19531,N_19568);
xnor U19686 (N_19686,N_19490,N_19523);
nor U19687 (N_19687,N_19504,N_19499);
or U19688 (N_19688,N_19520,N_19468);
xnor U19689 (N_19689,N_19423,N_19590);
or U19690 (N_19690,N_19445,N_19463);
or U19691 (N_19691,N_19402,N_19575);
and U19692 (N_19692,N_19486,N_19500);
nand U19693 (N_19693,N_19593,N_19469);
nand U19694 (N_19694,N_19416,N_19426);
or U19695 (N_19695,N_19535,N_19438);
nand U19696 (N_19696,N_19466,N_19418);
nand U19697 (N_19697,N_19461,N_19567);
or U19698 (N_19698,N_19544,N_19512);
and U19699 (N_19699,N_19420,N_19505);
xor U19700 (N_19700,N_19409,N_19557);
nor U19701 (N_19701,N_19526,N_19422);
and U19702 (N_19702,N_19552,N_19509);
or U19703 (N_19703,N_19512,N_19418);
or U19704 (N_19704,N_19463,N_19414);
and U19705 (N_19705,N_19401,N_19582);
xor U19706 (N_19706,N_19599,N_19466);
or U19707 (N_19707,N_19451,N_19473);
xnor U19708 (N_19708,N_19457,N_19445);
xnor U19709 (N_19709,N_19443,N_19422);
or U19710 (N_19710,N_19427,N_19445);
nor U19711 (N_19711,N_19550,N_19542);
xor U19712 (N_19712,N_19474,N_19417);
or U19713 (N_19713,N_19592,N_19472);
or U19714 (N_19714,N_19425,N_19534);
or U19715 (N_19715,N_19583,N_19498);
nand U19716 (N_19716,N_19442,N_19519);
xnor U19717 (N_19717,N_19442,N_19508);
or U19718 (N_19718,N_19594,N_19480);
or U19719 (N_19719,N_19420,N_19519);
nor U19720 (N_19720,N_19495,N_19558);
and U19721 (N_19721,N_19458,N_19400);
and U19722 (N_19722,N_19484,N_19425);
nor U19723 (N_19723,N_19521,N_19535);
and U19724 (N_19724,N_19540,N_19488);
nand U19725 (N_19725,N_19485,N_19557);
nand U19726 (N_19726,N_19430,N_19563);
nor U19727 (N_19727,N_19484,N_19422);
nand U19728 (N_19728,N_19519,N_19563);
nand U19729 (N_19729,N_19447,N_19505);
nor U19730 (N_19730,N_19429,N_19532);
and U19731 (N_19731,N_19412,N_19593);
or U19732 (N_19732,N_19487,N_19445);
nor U19733 (N_19733,N_19521,N_19476);
nand U19734 (N_19734,N_19492,N_19427);
nand U19735 (N_19735,N_19513,N_19467);
and U19736 (N_19736,N_19426,N_19566);
or U19737 (N_19737,N_19427,N_19586);
nor U19738 (N_19738,N_19432,N_19452);
nand U19739 (N_19739,N_19599,N_19528);
nor U19740 (N_19740,N_19444,N_19434);
nor U19741 (N_19741,N_19425,N_19515);
and U19742 (N_19742,N_19512,N_19554);
xor U19743 (N_19743,N_19426,N_19432);
nand U19744 (N_19744,N_19534,N_19412);
nor U19745 (N_19745,N_19477,N_19520);
or U19746 (N_19746,N_19410,N_19507);
and U19747 (N_19747,N_19516,N_19582);
xnor U19748 (N_19748,N_19580,N_19430);
nand U19749 (N_19749,N_19421,N_19529);
nand U19750 (N_19750,N_19425,N_19575);
or U19751 (N_19751,N_19408,N_19558);
xor U19752 (N_19752,N_19581,N_19584);
and U19753 (N_19753,N_19462,N_19502);
or U19754 (N_19754,N_19563,N_19447);
or U19755 (N_19755,N_19554,N_19497);
xnor U19756 (N_19756,N_19498,N_19573);
nand U19757 (N_19757,N_19562,N_19477);
and U19758 (N_19758,N_19568,N_19447);
nand U19759 (N_19759,N_19535,N_19478);
nand U19760 (N_19760,N_19587,N_19402);
and U19761 (N_19761,N_19478,N_19475);
nor U19762 (N_19762,N_19468,N_19472);
or U19763 (N_19763,N_19436,N_19533);
nand U19764 (N_19764,N_19477,N_19429);
xor U19765 (N_19765,N_19528,N_19478);
nor U19766 (N_19766,N_19580,N_19509);
nand U19767 (N_19767,N_19589,N_19457);
nand U19768 (N_19768,N_19584,N_19563);
and U19769 (N_19769,N_19497,N_19544);
nor U19770 (N_19770,N_19574,N_19465);
and U19771 (N_19771,N_19519,N_19515);
and U19772 (N_19772,N_19483,N_19469);
and U19773 (N_19773,N_19486,N_19467);
or U19774 (N_19774,N_19465,N_19496);
or U19775 (N_19775,N_19503,N_19463);
or U19776 (N_19776,N_19414,N_19475);
or U19777 (N_19777,N_19430,N_19581);
nor U19778 (N_19778,N_19593,N_19547);
xor U19779 (N_19779,N_19415,N_19478);
or U19780 (N_19780,N_19552,N_19482);
xnor U19781 (N_19781,N_19448,N_19561);
and U19782 (N_19782,N_19457,N_19425);
nand U19783 (N_19783,N_19455,N_19513);
xor U19784 (N_19784,N_19431,N_19416);
nand U19785 (N_19785,N_19562,N_19533);
or U19786 (N_19786,N_19585,N_19508);
and U19787 (N_19787,N_19552,N_19548);
or U19788 (N_19788,N_19577,N_19548);
nor U19789 (N_19789,N_19486,N_19436);
xnor U19790 (N_19790,N_19459,N_19466);
nor U19791 (N_19791,N_19522,N_19448);
nor U19792 (N_19792,N_19470,N_19530);
and U19793 (N_19793,N_19527,N_19440);
nand U19794 (N_19794,N_19484,N_19469);
nor U19795 (N_19795,N_19568,N_19413);
and U19796 (N_19796,N_19575,N_19488);
and U19797 (N_19797,N_19570,N_19509);
xnor U19798 (N_19798,N_19492,N_19474);
or U19799 (N_19799,N_19433,N_19421);
nand U19800 (N_19800,N_19679,N_19754);
nor U19801 (N_19801,N_19678,N_19694);
xor U19802 (N_19802,N_19723,N_19671);
nor U19803 (N_19803,N_19649,N_19607);
nor U19804 (N_19804,N_19625,N_19670);
nor U19805 (N_19805,N_19601,N_19697);
nor U19806 (N_19806,N_19627,N_19646);
nor U19807 (N_19807,N_19763,N_19779);
and U19808 (N_19808,N_19735,N_19715);
and U19809 (N_19809,N_19668,N_19630);
or U19810 (N_19810,N_19682,N_19609);
or U19811 (N_19811,N_19772,N_19714);
nor U19812 (N_19812,N_19762,N_19767);
nor U19813 (N_19813,N_19796,N_19699);
xor U19814 (N_19814,N_19680,N_19764);
nor U19815 (N_19815,N_19747,N_19766);
xor U19816 (N_19816,N_19736,N_19613);
nand U19817 (N_19817,N_19626,N_19750);
nor U19818 (N_19818,N_19794,N_19786);
or U19819 (N_19819,N_19732,N_19744);
nor U19820 (N_19820,N_19693,N_19645);
xnor U19821 (N_19821,N_19666,N_19662);
nand U19822 (N_19822,N_19780,N_19711);
or U19823 (N_19823,N_19660,N_19741);
and U19824 (N_19824,N_19717,N_19621);
nand U19825 (N_19825,N_19742,N_19651);
nand U19826 (N_19826,N_19691,N_19791);
nor U19827 (N_19827,N_19781,N_19797);
nor U19828 (N_19828,N_19698,N_19727);
or U19829 (N_19829,N_19792,N_19657);
nor U19830 (N_19830,N_19604,N_19676);
or U19831 (N_19831,N_19718,N_19749);
and U19832 (N_19832,N_19673,N_19640);
nor U19833 (N_19833,N_19739,N_19789);
or U19834 (N_19834,N_19667,N_19659);
nor U19835 (N_19835,N_19624,N_19687);
and U19836 (N_19836,N_19684,N_19755);
nand U19837 (N_19837,N_19610,N_19600);
xnor U19838 (N_19838,N_19740,N_19690);
xnor U19839 (N_19839,N_19704,N_19703);
or U19840 (N_19840,N_19701,N_19709);
nand U19841 (N_19841,N_19720,N_19719);
nand U19842 (N_19842,N_19793,N_19706);
and U19843 (N_19843,N_19643,N_19669);
nand U19844 (N_19844,N_19707,N_19788);
nand U19845 (N_19845,N_19637,N_19746);
nand U19846 (N_19846,N_19724,N_19716);
and U19847 (N_19847,N_19631,N_19665);
nor U19848 (N_19848,N_19777,N_19773);
xor U19849 (N_19849,N_19795,N_19710);
nand U19850 (N_19850,N_19708,N_19644);
or U19851 (N_19851,N_19752,N_19784);
nor U19852 (N_19852,N_19785,N_19765);
or U19853 (N_19853,N_19688,N_19775);
xor U19854 (N_19854,N_19738,N_19638);
and U19855 (N_19855,N_19743,N_19683);
xnor U19856 (N_19856,N_19611,N_19712);
nand U19857 (N_19857,N_19686,N_19639);
nand U19858 (N_19858,N_19648,N_19705);
or U19859 (N_19859,N_19776,N_19692);
xor U19860 (N_19860,N_19672,N_19636);
nor U19861 (N_19861,N_19725,N_19615);
nand U19862 (N_19862,N_19761,N_19658);
xnor U19863 (N_19863,N_19619,N_19602);
nand U19864 (N_19864,N_19632,N_19647);
xnor U19865 (N_19865,N_19650,N_19674);
xnor U19866 (N_19866,N_19799,N_19713);
and U19867 (N_19867,N_19603,N_19753);
and U19868 (N_19868,N_19617,N_19729);
xor U19869 (N_19869,N_19663,N_19737);
or U19870 (N_19870,N_19721,N_19722);
or U19871 (N_19871,N_19790,N_19745);
nand U19872 (N_19872,N_19677,N_19614);
nand U19873 (N_19873,N_19634,N_19618);
nand U19874 (N_19874,N_19778,N_19702);
xor U19875 (N_19875,N_19756,N_19655);
and U19876 (N_19876,N_19608,N_19748);
xnor U19877 (N_19877,N_19734,N_19787);
or U19878 (N_19878,N_19757,N_19652);
xnor U19879 (N_19879,N_19689,N_19760);
or U19880 (N_19880,N_19774,N_19782);
nand U19881 (N_19881,N_19642,N_19759);
and U19882 (N_19882,N_19623,N_19622);
nand U19883 (N_19883,N_19769,N_19770);
xnor U19884 (N_19884,N_19606,N_19664);
and U19885 (N_19885,N_19675,N_19696);
or U19886 (N_19886,N_19612,N_19620);
and U19887 (N_19887,N_19681,N_19635);
nor U19888 (N_19888,N_19728,N_19695);
and U19889 (N_19889,N_19726,N_19768);
xnor U19890 (N_19890,N_19798,N_19730);
nand U19891 (N_19891,N_19605,N_19685);
nand U19892 (N_19892,N_19731,N_19700);
nand U19893 (N_19893,N_19661,N_19783);
xnor U19894 (N_19894,N_19616,N_19771);
or U19895 (N_19895,N_19633,N_19629);
nor U19896 (N_19896,N_19641,N_19653);
and U19897 (N_19897,N_19751,N_19656);
xor U19898 (N_19898,N_19654,N_19733);
or U19899 (N_19899,N_19628,N_19758);
and U19900 (N_19900,N_19695,N_19654);
nor U19901 (N_19901,N_19623,N_19619);
xnor U19902 (N_19902,N_19680,N_19709);
xor U19903 (N_19903,N_19729,N_19650);
or U19904 (N_19904,N_19734,N_19694);
or U19905 (N_19905,N_19797,N_19752);
nor U19906 (N_19906,N_19630,N_19643);
nand U19907 (N_19907,N_19677,N_19773);
xnor U19908 (N_19908,N_19753,N_19621);
nor U19909 (N_19909,N_19798,N_19601);
nor U19910 (N_19910,N_19695,N_19726);
and U19911 (N_19911,N_19687,N_19788);
xor U19912 (N_19912,N_19601,N_19793);
nand U19913 (N_19913,N_19733,N_19775);
nand U19914 (N_19914,N_19747,N_19690);
and U19915 (N_19915,N_19610,N_19626);
and U19916 (N_19916,N_19751,N_19715);
and U19917 (N_19917,N_19790,N_19791);
and U19918 (N_19918,N_19642,N_19673);
nor U19919 (N_19919,N_19669,N_19756);
nand U19920 (N_19920,N_19797,N_19635);
nor U19921 (N_19921,N_19675,N_19639);
and U19922 (N_19922,N_19778,N_19696);
or U19923 (N_19923,N_19629,N_19718);
nand U19924 (N_19924,N_19786,N_19628);
nor U19925 (N_19925,N_19603,N_19705);
and U19926 (N_19926,N_19778,N_19724);
nand U19927 (N_19927,N_19753,N_19733);
nand U19928 (N_19928,N_19622,N_19707);
nand U19929 (N_19929,N_19633,N_19703);
nor U19930 (N_19930,N_19785,N_19725);
nor U19931 (N_19931,N_19687,N_19634);
and U19932 (N_19932,N_19789,N_19737);
nand U19933 (N_19933,N_19638,N_19602);
nand U19934 (N_19934,N_19638,N_19692);
or U19935 (N_19935,N_19705,N_19747);
or U19936 (N_19936,N_19620,N_19756);
and U19937 (N_19937,N_19641,N_19615);
xor U19938 (N_19938,N_19781,N_19626);
and U19939 (N_19939,N_19753,N_19784);
and U19940 (N_19940,N_19674,N_19720);
nand U19941 (N_19941,N_19786,N_19680);
nor U19942 (N_19942,N_19670,N_19657);
xor U19943 (N_19943,N_19767,N_19651);
or U19944 (N_19944,N_19623,N_19675);
nand U19945 (N_19945,N_19638,N_19726);
xor U19946 (N_19946,N_19651,N_19699);
and U19947 (N_19947,N_19738,N_19617);
or U19948 (N_19948,N_19671,N_19792);
and U19949 (N_19949,N_19744,N_19621);
nor U19950 (N_19950,N_19613,N_19769);
nand U19951 (N_19951,N_19658,N_19747);
nor U19952 (N_19952,N_19747,N_19773);
nor U19953 (N_19953,N_19765,N_19743);
or U19954 (N_19954,N_19725,N_19672);
or U19955 (N_19955,N_19724,N_19726);
nor U19956 (N_19956,N_19796,N_19754);
or U19957 (N_19957,N_19706,N_19750);
and U19958 (N_19958,N_19644,N_19631);
nand U19959 (N_19959,N_19619,N_19787);
nor U19960 (N_19960,N_19625,N_19799);
xor U19961 (N_19961,N_19646,N_19765);
nand U19962 (N_19962,N_19745,N_19615);
nand U19963 (N_19963,N_19717,N_19782);
and U19964 (N_19964,N_19697,N_19785);
nand U19965 (N_19965,N_19775,N_19612);
or U19966 (N_19966,N_19621,N_19684);
or U19967 (N_19967,N_19603,N_19606);
xor U19968 (N_19968,N_19684,N_19731);
xor U19969 (N_19969,N_19791,N_19780);
nand U19970 (N_19970,N_19642,N_19760);
xor U19971 (N_19971,N_19749,N_19796);
or U19972 (N_19972,N_19724,N_19648);
xor U19973 (N_19973,N_19711,N_19622);
nand U19974 (N_19974,N_19688,N_19746);
xor U19975 (N_19975,N_19780,N_19712);
nand U19976 (N_19976,N_19656,N_19601);
nor U19977 (N_19977,N_19730,N_19620);
xor U19978 (N_19978,N_19639,N_19685);
or U19979 (N_19979,N_19634,N_19792);
nor U19980 (N_19980,N_19647,N_19625);
and U19981 (N_19981,N_19625,N_19674);
nand U19982 (N_19982,N_19735,N_19609);
xor U19983 (N_19983,N_19767,N_19790);
nand U19984 (N_19984,N_19774,N_19663);
nor U19985 (N_19985,N_19743,N_19608);
nand U19986 (N_19986,N_19644,N_19794);
nor U19987 (N_19987,N_19667,N_19775);
and U19988 (N_19988,N_19693,N_19652);
nor U19989 (N_19989,N_19659,N_19712);
xnor U19990 (N_19990,N_19728,N_19689);
xnor U19991 (N_19991,N_19642,N_19683);
nor U19992 (N_19992,N_19613,N_19783);
nand U19993 (N_19993,N_19658,N_19609);
xor U19994 (N_19994,N_19629,N_19738);
nand U19995 (N_19995,N_19653,N_19782);
nand U19996 (N_19996,N_19798,N_19687);
xnor U19997 (N_19997,N_19694,N_19617);
and U19998 (N_19998,N_19785,N_19653);
xor U19999 (N_19999,N_19701,N_19657);
and UO_0 (O_0,N_19885,N_19959);
nand UO_1 (O_1,N_19891,N_19962);
or UO_2 (O_2,N_19915,N_19889);
nand UO_3 (O_3,N_19957,N_19807);
and UO_4 (O_4,N_19861,N_19966);
nand UO_5 (O_5,N_19803,N_19883);
or UO_6 (O_6,N_19832,N_19984);
nand UO_7 (O_7,N_19894,N_19995);
and UO_8 (O_8,N_19846,N_19872);
or UO_9 (O_9,N_19992,N_19963);
nand UO_10 (O_10,N_19802,N_19845);
or UO_11 (O_11,N_19912,N_19982);
and UO_12 (O_12,N_19970,N_19818);
and UO_13 (O_13,N_19882,N_19838);
nor UO_14 (O_14,N_19911,N_19909);
and UO_15 (O_15,N_19814,N_19965);
xor UO_16 (O_16,N_19948,N_19858);
and UO_17 (O_17,N_19835,N_19870);
or UO_18 (O_18,N_19997,N_19810);
xor UO_19 (O_19,N_19955,N_19827);
or UO_20 (O_20,N_19923,N_19864);
or UO_21 (O_21,N_19983,N_19991);
nand UO_22 (O_22,N_19905,N_19893);
and UO_23 (O_23,N_19886,N_19951);
nor UO_24 (O_24,N_19877,N_19918);
nor UO_25 (O_25,N_19840,N_19985);
or UO_26 (O_26,N_19956,N_19800);
nand UO_27 (O_27,N_19866,N_19859);
or UO_28 (O_28,N_19841,N_19852);
and UO_29 (O_29,N_19953,N_19935);
and UO_30 (O_30,N_19813,N_19968);
and UO_31 (O_31,N_19952,N_19820);
xor UO_32 (O_32,N_19898,N_19831);
nand UO_33 (O_33,N_19837,N_19920);
and UO_34 (O_34,N_19849,N_19925);
nor UO_35 (O_35,N_19843,N_19830);
xnor UO_36 (O_36,N_19922,N_19809);
or UO_37 (O_37,N_19977,N_19884);
or UO_38 (O_38,N_19943,N_19961);
xnor UO_39 (O_39,N_19853,N_19890);
nor UO_40 (O_40,N_19805,N_19811);
and UO_41 (O_41,N_19910,N_19914);
nor UO_42 (O_42,N_19850,N_19931);
xnor UO_43 (O_43,N_19823,N_19851);
nor UO_44 (O_44,N_19919,N_19871);
or UO_45 (O_45,N_19806,N_19828);
xor UO_46 (O_46,N_19873,N_19964);
nand UO_47 (O_47,N_19990,N_19825);
xnor UO_48 (O_48,N_19987,N_19979);
or UO_49 (O_49,N_19801,N_19933);
or UO_50 (O_50,N_19892,N_19836);
xor UO_51 (O_51,N_19904,N_19865);
nand UO_52 (O_52,N_19895,N_19969);
nor UO_53 (O_53,N_19896,N_19868);
and UO_54 (O_54,N_19842,N_19958);
nor UO_55 (O_55,N_19942,N_19917);
or UO_56 (O_56,N_19879,N_19834);
or UO_57 (O_57,N_19869,N_19934);
and UO_58 (O_58,N_19973,N_19875);
nand UO_59 (O_59,N_19899,N_19876);
or UO_60 (O_60,N_19857,N_19817);
and UO_61 (O_61,N_19862,N_19816);
nand UO_62 (O_62,N_19902,N_19900);
or UO_63 (O_63,N_19906,N_19901);
and UO_64 (O_64,N_19939,N_19867);
xor UO_65 (O_65,N_19921,N_19822);
nor UO_66 (O_66,N_19993,N_19996);
nand UO_67 (O_67,N_19897,N_19854);
nand UO_68 (O_68,N_19887,N_19916);
nand UO_69 (O_69,N_19998,N_19888);
nor UO_70 (O_70,N_19978,N_19949);
or UO_71 (O_71,N_19945,N_19860);
or UO_72 (O_72,N_19960,N_19981);
xor UO_73 (O_73,N_19954,N_19881);
nand UO_74 (O_74,N_19847,N_19880);
xnor UO_75 (O_75,N_19839,N_19930);
nor UO_76 (O_76,N_19994,N_19974);
xor UO_77 (O_77,N_19913,N_19844);
and UO_78 (O_78,N_19826,N_19928);
xnor UO_79 (O_79,N_19936,N_19819);
nor UO_80 (O_80,N_19808,N_19947);
xor UO_81 (O_81,N_19856,N_19967);
or UO_82 (O_82,N_19824,N_19940);
xnor UO_83 (O_83,N_19821,N_19907);
and UO_84 (O_84,N_19924,N_19975);
nor UO_85 (O_85,N_19855,N_19833);
xor UO_86 (O_86,N_19999,N_19946);
xor UO_87 (O_87,N_19863,N_19932);
nor UO_88 (O_88,N_19988,N_19941);
and UO_89 (O_89,N_19938,N_19976);
or UO_90 (O_90,N_19950,N_19815);
nand UO_91 (O_91,N_19986,N_19829);
nor UO_92 (O_92,N_19926,N_19903);
or UO_93 (O_93,N_19937,N_19972);
and UO_94 (O_94,N_19804,N_19812);
nand UO_95 (O_95,N_19848,N_19980);
nand UO_96 (O_96,N_19878,N_19927);
xor UO_97 (O_97,N_19908,N_19944);
xor UO_98 (O_98,N_19874,N_19929);
nand UO_99 (O_99,N_19971,N_19989);
and UO_100 (O_100,N_19804,N_19900);
nor UO_101 (O_101,N_19996,N_19970);
nand UO_102 (O_102,N_19874,N_19879);
and UO_103 (O_103,N_19829,N_19980);
xor UO_104 (O_104,N_19862,N_19808);
and UO_105 (O_105,N_19943,N_19889);
nor UO_106 (O_106,N_19864,N_19952);
nand UO_107 (O_107,N_19833,N_19901);
and UO_108 (O_108,N_19880,N_19961);
or UO_109 (O_109,N_19904,N_19859);
nor UO_110 (O_110,N_19982,N_19971);
and UO_111 (O_111,N_19837,N_19820);
nor UO_112 (O_112,N_19854,N_19973);
or UO_113 (O_113,N_19910,N_19919);
nand UO_114 (O_114,N_19938,N_19893);
or UO_115 (O_115,N_19858,N_19877);
or UO_116 (O_116,N_19897,N_19921);
nand UO_117 (O_117,N_19910,N_19903);
nand UO_118 (O_118,N_19819,N_19857);
nor UO_119 (O_119,N_19971,N_19891);
and UO_120 (O_120,N_19804,N_19947);
or UO_121 (O_121,N_19826,N_19898);
or UO_122 (O_122,N_19825,N_19813);
xnor UO_123 (O_123,N_19938,N_19939);
or UO_124 (O_124,N_19952,N_19973);
nor UO_125 (O_125,N_19988,N_19876);
nand UO_126 (O_126,N_19924,N_19855);
xnor UO_127 (O_127,N_19959,N_19902);
and UO_128 (O_128,N_19867,N_19802);
xnor UO_129 (O_129,N_19852,N_19910);
or UO_130 (O_130,N_19997,N_19896);
xnor UO_131 (O_131,N_19994,N_19975);
nand UO_132 (O_132,N_19801,N_19805);
and UO_133 (O_133,N_19982,N_19887);
xor UO_134 (O_134,N_19964,N_19950);
xor UO_135 (O_135,N_19824,N_19972);
nand UO_136 (O_136,N_19921,N_19905);
nand UO_137 (O_137,N_19806,N_19864);
xnor UO_138 (O_138,N_19907,N_19858);
nor UO_139 (O_139,N_19966,N_19950);
nand UO_140 (O_140,N_19939,N_19813);
nor UO_141 (O_141,N_19812,N_19872);
xnor UO_142 (O_142,N_19983,N_19845);
or UO_143 (O_143,N_19852,N_19897);
nor UO_144 (O_144,N_19883,N_19902);
or UO_145 (O_145,N_19903,N_19944);
xnor UO_146 (O_146,N_19815,N_19824);
or UO_147 (O_147,N_19999,N_19956);
xor UO_148 (O_148,N_19904,N_19850);
and UO_149 (O_149,N_19928,N_19804);
nand UO_150 (O_150,N_19912,N_19860);
nor UO_151 (O_151,N_19880,N_19956);
nand UO_152 (O_152,N_19853,N_19858);
and UO_153 (O_153,N_19962,N_19835);
nand UO_154 (O_154,N_19948,N_19982);
nand UO_155 (O_155,N_19982,N_19803);
nor UO_156 (O_156,N_19991,N_19801);
and UO_157 (O_157,N_19896,N_19938);
nand UO_158 (O_158,N_19966,N_19830);
nand UO_159 (O_159,N_19936,N_19853);
or UO_160 (O_160,N_19980,N_19883);
or UO_161 (O_161,N_19873,N_19917);
xor UO_162 (O_162,N_19870,N_19889);
nor UO_163 (O_163,N_19877,N_19965);
nor UO_164 (O_164,N_19976,N_19982);
nand UO_165 (O_165,N_19943,N_19810);
and UO_166 (O_166,N_19874,N_19983);
or UO_167 (O_167,N_19939,N_19869);
or UO_168 (O_168,N_19928,N_19880);
and UO_169 (O_169,N_19911,N_19846);
and UO_170 (O_170,N_19901,N_19915);
or UO_171 (O_171,N_19808,N_19888);
xnor UO_172 (O_172,N_19889,N_19919);
and UO_173 (O_173,N_19989,N_19940);
xnor UO_174 (O_174,N_19809,N_19872);
and UO_175 (O_175,N_19917,N_19863);
nand UO_176 (O_176,N_19877,N_19823);
nand UO_177 (O_177,N_19810,N_19820);
xnor UO_178 (O_178,N_19936,N_19971);
nand UO_179 (O_179,N_19889,N_19802);
or UO_180 (O_180,N_19959,N_19942);
or UO_181 (O_181,N_19839,N_19953);
or UO_182 (O_182,N_19826,N_19912);
or UO_183 (O_183,N_19978,N_19970);
nand UO_184 (O_184,N_19960,N_19832);
nor UO_185 (O_185,N_19895,N_19937);
or UO_186 (O_186,N_19919,N_19986);
and UO_187 (O_187,N_19998,N_19910);
nand UO_188 (O_188,N_19997,N_19959);
nand UO_189 (O_189,N_19808,N_19965);
and UO_190 (O_190,N_19869,N_19966);
and UO_191 (O_191,N_19902,N_19865);
xor UO_192 (O_192,N_19890,N_19858);
or UO_193 (O_193,N_19940,N_19844);
nand UO_194 (O_194,N_19884,N_19866);
and UO_195 (O_195,N_19877,N_19924);
xnor UO_196 (O_196,N_19899,N_19800);
nor UO_197 (O_197,N_19871,N_19953);
nor UO_198 (O_198,N_19983,N_19942);
or UO_199 (O_199,N_19941,N_19898);
nor UO_200 (O_200,N_19852,N_19834);
and UO_201 (O_201,N_19956,N_19859);
and UO_202 (O_202,N_19847,N_19991);
nor UO_203 (O_203,N_19972,N_19985);
xnor UO_204 (O_204,N_19929,N_19813);
or UO_205 (O_205,N_19977,N_19969);
xor UO_206 (O_206,N_19931,N_19889);
nand UO_207 (O_207,N_19825,N_19849);
nand UO_208 (O_208,N_19937,N_19824);
nor UO_209 (O_209,N_19861,N_19915);
or UO_210 (O_210,N_19955,N_19979);
nand UO_211 (O_211,N_19993,N_19827);
nor UO_212 (O_212,N_19821,N_19916);
nand UO_213 (O_213,N_19989,N_19951);
and UO_214 (O_214,N_19953,N_19835);
nand UO_215 (O_215,N_19940,N_19929);
nor UO_216 (O_216,N_19821,N_19997);
nand UO_217 (O_217,N_19917,N_19980);
nand UO_218 (O_218,N_19814,N_19933);
xnor UO_219 (O_219,N_19901,N_19800);
and UO_220 (O_220,N_19908,N_19920);
and UO_221 (O_221,N_19934,N_19808);
nand UO_222 (O_222,N_19977,N_19853);
nand UO_223 (O_223,N_19886,N_19905);
and UO_224 (O_224,N_19909,N_19836);
nand UO_225 (O_225,N_19878,N_19984);
xnor UO_226 (O_226,N_19886,N_19974);
and UO_227 (O_227,N_19964,N_19920);
xor UO_228 (O_228,N_19873,N_19878);
nand UO_229 (O_229,N_19840,N_19987);
nand UO_230 (O_230,N_19853,N_19941);
nor UO_231 (O_231,N_19898,N_19870);
nor UO_232 (O_232,N_19848,N_19817);
or UO_233 (O_233,N_19853,N_19940);
nand UO_234 (O_234,N_19814,N_19971);
or UO_235 (O_235,N_19870,N_19844);
xor UO_236 (O_236,N_19886,N_19980);
and UO_237 (O_237,N_19854,N_19986);
and UO_238 (O_238,N_19938,N_19852);
or UO_239 (O_239,N_19809,N_19819);
or UO_240 (O_240,N_19870,N_19911);
nand UO_241 (O_241,N_19904,N_19975);
nand UO_242 (O_242,N_19976,N_19857);
xor UO_243 (O_243,N_19997,N_19940);
xnor UO_244 (O_244,N_19882,N_19935);
xor UO_245 (O_245,N_19934,N_19891);
nor UO_246 (O_246,N_19874,N_19894);
or UO_247 (O_247,N_19847,N_19972);
xnor UO_248 (O_248,N_19829,N_19820);
or UO_249 (O_249,N_19898,N_19841);
or UO_250 (O_250,N_19947,N_19857);
and UO_251 (O_251,N_19919,N_19959);
and UO_252 (O_252,N_19982,N_19923);
or UO_253 (O_253,N_19889,N_19906);
or UO_254 (O_254,N_19991,N_19863);
nand UO_255 (O_255,N_19988,N_19998);
and UO_256 (O_256,N_19956,N_19855);
and UO_257 (O_257,N_19914,N_19868);
or UO_258 (O_258,N_19806,N_19964);
nand UO_259 (O_259,N_19988,N_19987);
or UO_260 (O_260,N_19823,N_19970);
xnor UO_261 (O_261,N_19828,N_19891);
nand UO_262 (O_262,N_19971,N_19830);
xnor UO_263 (O_263,N_19899,N_19820);
nor UO_264 (O_264,N_19817,N_19872);
xnor UO_265 (O_265,N_19907,N_19896);
nand UO_266 (O_266,N_19915,N_19906);
and UO_267 (O_267,N_19978,N_19910);
nand UO_268 (O_268,N_19841,N_19914);
or UO_269 (O_269,N_19826,N_19965);
nand UO_270 (O_270,N_19880,N_19809);
nand UO_271 (O_271,N_19902,N_19970);
or UO_272 (O_272,N_19994,N_19925);
and UO_273 (O_273,N_19893,N_19874);
nor UO_274 (O_274,N_19935,N_19803);
and UO_275 (O_275,N_19816,N_19921);
nand UO_276 (O_276,N_19872,N_19947);
nor UO_277 (O_277,N_19862,N_19877);
nand UO_278 (O_278,N_19948,N_19959);
and UO_279 (O_279,N_19917,N_19811);
and UO_280 (O_280,N_19912,N_19960);
and UO_281 (O_281,N_19808,N_19833);
nor UO_282 (O_282,N_19936,N_19889);
nor UO_283 (O_283,N_19993,N_19970);
or UO_284 (O_284,N_19922,N_19999);
nand UO_285 (O_285,N_19899,N_19941);
nand UO_286 (O_286,N_19908,N_19911);
xnor UO_287 (O_287,N_19966,N_19842);
nand UO_288 (O_288,N_19875,N_19847);
or UO_289 (O_289,N_19873,N_19887);
xnor UO_290 (O_290,N_19978,N_19836);
and UO_291 (O_291,N_19821,N_19901);
xor UO_292 (O_292,N_19836,N_19950);
and UO_293 (O_293,N_19812,N_19929);
or UO_294 (O_294,N_19939,N_19891);
and UO_295 (O_295,N_19929,N_19912);
xnor UO_296 (O_296,N_19844,N_19850);
nor UO_297 (O_297,N_19857,N_19884);
xor UO_298 (O_298,N_19975,N_19990);
nor UO_299 (O_299,N_19840,N_19895);
nor UO_300 (O_300,N_19992,N_19999);
or UO_301 (O_301,N_19932,N_19835);
or UO_302 (O_302,N_19978,N_19880);
xnor UO_303 (O_303,N_19811,N_19931);
and UO_304 (O_304,N_19917,N_19993);
nand UO_305 (O_305,N_19972,N_19918);
nor UO_306 (O_306,N_19822,N_19848);
xor UO_307 (O_307,N_19931,N_19817);
nand UO_308 (O_308,N_19969,N_19952);
nor UO_309 (O_309,N_19866,N_19870);
or UO_310 (O_310,N_19899,N_19888);
nand UO_311 (O_311,N_19963,N_19816);
or UO_312 (O_312,N_19960,N_19828);
xnor UO_313 (O_313,N_19808,N_19967);
and UO_314 (O_314,N_19892,N_19837);
xnor UO_315 (O_315,N_19864,N_19986);
nor UO_316 (O_316,N_19815,N_19975);
or UO_317 (O_317,N_19908,N_19919);
and UO_318 (O_318,N_19916,N_19912);
and UO_319 (O_319,N_19811,N_19926);
nor UO_320 (O_320,N_19987,N_19875);
or UO_321 (O_321,N_19811,N_19858);
xnor UO_322 (O_322,N_19813,N_19904);
nand UO_323 (O_323,N_19815,N_19853);
nor UO_324 (O_324,N_19836,N_19855);
or UO_325 (O_325,N_19835,N_19867);
nand UO_326 (O_326,N_19959,N_19994);
and UO_327 (O_327,N_19943,N_19904);
and UO_328 (O_328,N_19964,N_19827);
nand UO_329 (O_329,N_19835,N_19989);
nor UO_330 (O_330,N_19970,N_19831);
or UO_331 (O_331,N_19952,N_19857);
and UO_332 (O_332,N_19939,N_19916);
nor UO_333 (O_333,N_19970,N_19982);
or UO_334 (O_334,N_19832,N_19891);
or UO_335 (O_335,N_19989,N_19845);
nand UO_336 (O_336,N_19925,N_19920);
and UO_337 (O_337,N_19845,N_19817);
nor UO_338 (O_338,N_19992,N_19868);
and UO_339 (O_339,N_19820,N_19812);
and UO_340 (O_340,N_19982,N_19990);
nor UO_341 (O_341,N_19895,N_19908);
nor UO_342 (O_342,N_19812,N_19845);
or UO_343 (O_343,N_19964,N_19955);
nor UO_344 (O_344,N_19813,N_19937);
or UO_345 (O_345,N_19928,N_19961);
nand UO_346 (O_346,N_19871,N_19878);
nor UO_347 (O_347,N_19950,N_19954);
nor UO_348 (O_348,N_19888,N_19849);
nor UO_349 (O_349,N_19808,N_19917);
nand UO_350 (O_350,N_19850,N_19807);
or UO_351 (O_351,N_19960,N_19990);
and UO_352 (O_352,N_19993,N_19966);
and UO_353 (O_353,N_19857,N_19888);
xnor UO_354 (O_354,N_19925,N_19949);
xnor UO_355 (O_355,N_19863,N_19998);
nor UO_356 (O_356,N_19949,N_19819);
nor UO_357 (O_357,N_19800,N_19945);
xor UO_358 (O_358,N_19896,N_19853);
or UO_359 (O_359,N_19980,N_19909);
nor UO_360 (O_360,N_19837,N_19995);
and UO_361 (O_361,N_19843,N_19861);
or UO_362 (O_362,N_19873,N_19857);
and UO_363 (O_363,N_19960,N_19904);
or UO_364 (O_364,N_19970,N_19928);
or UO_365 (O_365,N_19873,N_19816);
and UO_366 (O_366,N_19915,N_19975);
nor UO_367 (O_367,N_19926,N_19870);
or UO_368 (O_368,N_19835,N_19991);
and UO_369 (O_369,N_19839,N_19971);
nor UO_370 (O_370,N_19971,N_19974);
xor UO_371 (O_371,N_19843,N_19887);
xor UO_372 (O_372,N_19927,N_19921);
and UO_373 (O_373,N_19894,N_19970);
and UO_374 (O_374,N_19942,N_19990);
nand UO_375 (O_375,N_19954,N_19946);
nand UO_376 (O_376,N_19802,N_19941);
xnor UO_377 (O_377,N_19824,N_19812);
nand UO_378 (O_378,N_19890,N_19902);
nor UO_379 (O_379,N_19975,N_19823);
nand UO_380 (O_380,N_19947,N_19852);
nand UO_381 (O_381,N_19827,N_19895);
nor UO_382 (O_382,N_19829,N_19915);
or UO_383 (O_383,N_19827,N_19900);
nand UO_384 (O_384,N_19941,N_19969);
and UO_385 (O_385,N_19914,N_19973);
nand UO_386 (O_386,N_19824,N_19854);
or UO_387 (O_387,N_19845,N_19835);
and UO_388 (O_388,N_19818,N_19877);
or UO_389 (O_389,N_19837,N_19957);
and UO_390 (O_390,N_19960,N_19853);
or UO_391 (O_391,N_19863,N_19984);
xor UO_392 (O_392,N_19869,N_19901);
or UO_393 (O_393,N_19808,N_19889);
and UO_394 (O_394,N_19997,N_19978);
nand UO_395 (O_395,N_19943,N_19995);
nor UO_396 (O_396,N_19864,N_19820);
and UO_397 (O_397,N_19935,N_19892);
nor UO_398 (O_398,N_19982,N_19992);
nand UO_399 (O_399,N_19925,N_19928);
and UO_400 (O_400,N_19983,N_19841);
and UO_401 (O_401,N_19913,N_19912);
or UO_402 (O_402,N_19867,N_19936);
nand UO_403 (O_403,N_19900,N_19925);
and UO_404 (O_404,N_19947,N_19858);
or UO_405 (O_405,N_19863,N_19927);
nand UO_406 (O_406,N_19843,N_19829);
or UO_407 (O_407,N_19966,N_19982);
and UO_408 (O_408,N_19942,N_19919);
nand UO_409 (O_409,N_19825,N_19920);
nor UO_410 (O_410,N_19820,N_19986);
nor UO_411 (O_411,N_19980,N_19965);
nand UO_412 (O_412,N_19977,N_19915);
xor UO_413 (O_413,N_19851,N_19955);
nor UO_414 (O_414,N_19860,N_19870);
or UO_415 (O_415,N_19835,N_19946);
or UO_416 (O_416,N_19857,N_19978);
xnor UO_417 (O_417,N_19835,N_19971);
nand UO_418 (O_418,N_19987,N_19926);
nor UO_419 (O_419,N_19910,N_19987);
nor UO_420 (O_420,N_19973,N_19953);
nand UO_421 (O_421,N_19867,N_19908);
nor UO_422 (O_422,N_19890,N_19889);
nor UO_423 (O_423,N_19994,N_19936);
xor UO_424 (O_424,N_19928,N_19995);
and UO_425 (O_425,N_19903,N_19954);
nor UO_426 (O_426,N_19941,N_19800);
xnor UO_427 (O_427,N_19997,N_19891);
and UO_428 (O_428,N_19879,N_19990);
nand UO_429 (O_429,N_19975,N_19814);
nor UO_430 (O_430,N_19803,N_19991);
xnor UO_431 (O_431,N_19913,N_19933);
xor UO_432 (O_432,N_19845,N_19841);
or UO_433 (O_433,N_19940,N_19829);
nor UO_434 (O_434,N_19936,N_19944);
and UO_435 (O_435,N_19922,N_19937);
nand UO_436 (O_436,N_19884,N_19990);
or UO_437 (O_437,N_19833,N_19960);
or UO_438 (O_438,N_19916,N_19925);
nor UO_439 (O_439,N_19918,N_19984);
nor UO_440 (O_440,N_19838,N_19892);
or UO_441 (O_441,N_19814,N_19877);
and UO_442 (O_442,N_19932,N_19807);
nand UO_443 (O_443,N_19811,N_19839);
and UO_444 (O_444,N_19999,N_19813);
xor UO_445 (O_445,N_19919,N_19876);
or UO_446 (O_446,N_19993,N_19820);
nor UO_447 (O_447,N_19876,N_19811);
nand UO_448 (O_448,N_19993,N_19903);
or UO_449 (O_449,N_19836,N_19803);
xnor UO_450 (O_450,N_19917,N_19825);
and UO_451 (O_451,N_19947,N_19987);
nand UO_452 (O_452,N_19936,N_19800);
or UO_453 (O_453,N_19841,N_19947);
nor UO_454 (O_454,N_19850,N_19840);
xor UO_455 (O_455,N_19951,N_19884);
xor UO_456 (O_456,N_19991,N_19842);
xor UO_457 (O_457,N_19810,N_19846);
nor UO_458 (O_458,N_19809,N_19861);
nor UO_459 (O_459,N_19908,N_19970);
nand UO_460 (O_460,N_19817,N_19916);
or UO_461 (O_461,N_19953,N_19951);
nor UO_462 (O_462,N_19905,N_19972);
and UO_463 (O_463,N_19923,N_19854);
nor UO_464 (O_464,N_19931,N_19942);
nand UO_465 (O_465,N_19953,N_19802);
nand UO_466 (O_466,N_19901,N_19832);
nor UO_467 (O_467,N_19999,N_19995);
xnor UO_468 (O_468,N_19811,N_19889);
nor UO_469 (O_469,N_19959,N_19802);
and UO_470 (O_470,N_19817,N_19830);
nor UO_471 (O_471,N_19958,N_19973);
nand UO_472 (O_472,N_19951,N_19917);
nand UO_473 (O_473,N_19810,N_19909);
xor UO_474 (O_474,N_19964,N_19947);
nor UO_475 (O_475,N_19959,N_19950);
and UO_476 (O_476,N_19805,N_19833);
or UO_477 (O_477,N_19912,N_19925);
nand UO_478 (O_478,N_19859,N_19858);
and UO_479 (O_479,N_19952,N_19876);
and UO_480 (O_480,N_19853,N_19814);
and UO_481 (O_481,N_19838,N_19880);
nor UO_482 (O_482,N_19832,N_19865);
xnor UO_483 (O_483,N_19918,N_19988);
xor UO_484 (O_484,N_19808,N_19926);
xor UO_485 (O_485,N_19825,N_19985);
nand UO_486 (O_486,N_19834,N_19994);
and UO_487 (O_487,N_19849,N_19976);
nand UO_488 (O_488,N_19920,N_19872);
or UO_489 (O_489,N_19917,N_19814);
nand UO_490 (O_490,N_19989,N_19810);
or UO_491 (O_491,N_19967,N_19899);
and UO_492 (O_492,N_19944,N_19912);
nor UO_493 (O_493,N_19917,N_19906);
xor UO_494 (O_494,N_19906,N_19902);
or UO_495 (O_495,N_19883,N_19916);
nand UO_496 (O_496,N_19817,N_19849);
nor UO_497 (O_497,N_19969,N_19982);
nand UO_498 (O_498,N_19899,N_19992);
nor UO_499 (O_499,N_19836,N_19974);
or UO_500 (O_500,N_19925,N_19803);
xor UO_501 (O_501,N_19805,N_19816);
xnor UO_502 (O_502,N_19822,N_19906);
xnor UO_503 (O_503,N_19860,N_19913);
nand UO_504 (O_504,N_19977,N_19843);
or UO_505 (O_505,N_19874,N_19978);
and UO_506 (O_506,N_19855,N_19823);
and UO_507 (O_507,N_19800,N_19867);
nand UO_508 (O_508,N_19935,N_19888);
nand UO_509 (O_509,N_19909,N_19887);
and UO_510 (O_510,N_19807,N_19937);
nor UO_511 (O_511,N_19944,N_19857);
and UO_512 (O_512,N_19890,N_19941);
or UO_513 (O_513,N_19935,N_19895);
nand UO_514 (O_514,N_19995,N_19897);
and UO_515 (O_515,N_19920,N_19855);
nand UO_516 (O_516,N_19904,N_19902);
xor UO_517 (O_517,N_19896,N_19986);
nand UO_518 (O_518,N_19852,N_19990);
nor UO_519 (O_519,N_19967,N_19800);
xnor UO_520 (O_520,N_19804,N_19873);
nand UO_521 (O_521,N_19990,N_19851);
and UO_522 (O_522,N_19866,N_19868);
nor UO_523 (O_523,N_19867,N_19989);
xor UO_524 (O_524,N_19962,N_19992);
nor UO_525 (O_525,N_19818,N_19979);
nor UO_526 (O_526,N_19810,N_19801);
xor UO_527 (O_527,N_19815,N_19917);
nand UO_528 (O_528,N_19986,N_19893);
and UO_529 (O_529,N_19891,N_19834);
or UO_530 (O_530,N_19827,N_19965);
xor UO_531 (O_531,N_19987,N_19862);
nand UO_532 (O_532,N_19841,N_19839);
nand UO_533 (O_533,N_19848,N_19958);
nor UO_534 (O_534,N_19934,N_19990);
xor UO_535 (O_535,N_19810,N_19867);
or UO_536 (O_536,N_19957,N_19952);
nand UO_537 (O_537,N_19814,N_19839);
xor UO_538 (O_538,N_19947,N_19867);
nand UO_539 (O_539,N_19803,N_19840);
nand UO_540 (O_540,N_19923,N_19939);
nor UO_541 (O_541,N_19843,N_19996);
nor UO_542 (O_542,N_19808,N_19817);
and UO_543 (O_543,N_19935,N_19889);
nor UO_544 (O_544,N_19864,N_19880);
and UO_545 (O_545,N_19951,N_19859);
and UO_546 (O_546,N_19803,N_19952);
nor UO_547 (O_547,N_19966,N_19880);
or UO_548 (O_548,N_19923,N_19913);
nand UO_549 (O_549,N_19836,N_19955);
nor UO_550 (O_550,N_19991,N_19980);
xor UO_551 (O_551,N_19957,N_19855);
xnor UO_552 (O_552,N_19852,N_19944);
or UO_553 (O_553,N_19973,N_19999);
nor UO_554 (O_554,N_19882,N_19896);
nor UO_555 (O_555,N_19847,N_19944);
nor UO_556 (O_556,N_19920,N_19853);
or UO_557 (O_557,N_19912,N_19881);
or UO_558 (O_558,N_19914,N_19932);
and UO_559 (O_559,N_19950,N_19807);
and UO_560 (O_560,N_19855,N_19970);
nor UO_561 (O_561,N_19830,N_19998);
and UO_562 (O_562,N_19802,N_19824);
xnor UO_563 (O_563,N_19883,N_19912);
nor UO_564 (O_564,N_19961,N_19870);
or UO_565 (O_565,N_19865,N_19953);
xor UO_566 (O_566,N_19947,N_19934);
nand UO_567 (O_567,N_19966,N_19836);
nor UO_568 (O_568,N_19835,N_19957);
and UO_569 (O_569,N_19895,N_19832);
or UO_570 (O_570,N_19997,N_19853);
nor UO_571 (O_571,N_19929,N_19942);
nor UO_572 (O_572,N_19880,N_19827);
xor UO_573 (O_573,N_19862,N_19933);
nand UO_574 (O_574,N_19872,N_19829);
xor UO_575 (O_575,N_19957,N_19843);
xnor UO_576 (O_576,N_19801,N_19978);
or UO_577 (O_577,N_19961,N_19906);
nor UO_578 (O_578,N_19958,N_19945);
nor UO_579 (O_579,N_19831,N_19887);
nor UO_580 (O_580,N_19941,N_19896);
nand UO_581 (O_581,N_19813,N_19801);
nand UO_582 (O_582,N_19883,N_19847);
nand UO_583 (O_583,N_19875,N_19992);
xor UO_584 (O_584,N_19938,N_19943);
nand UO_585 (O_585,N_19960,N_19957);
nor UO_586 (O_586,N_19827,N_19963);
nand UO_587 (O_587,N_19874,N_19835);
or UO_588 (O_588,N_19829,N_19822);
xor UO_589 (O_589,N_19945,N_19828);
or UO_590 (O_590,N_19843,N_19967);
nor UO_591 (O_591,N_19922,N_19926);
nand UO_592 (O_592,N_19847,N_19864);
nor UO_593 (O_593,N_19801,N_19828);
or UO_594 (O_594,N_19812,N_19936);
or UO_595 (O_595,N_19879,N_19885);
nand UO_596 (O_596,N_19922,N_19803);
nand UO_597 (O_597,N_19939,N_19843);
and UO_598 (O_598,N_19901,N_19873);
and UO_599 (O_599,N_19900,N_19857);
or UO_600 (O_600,N_19808,N_19876);
or UO_601 (O_601,N_19883,N_19893);
or UO_602 (O_602,N_19947,N_19860);
nor UO_603 (O_603,N_19883,N_19855);
nor UO_604 (O_604,N_19827,N_19989);
nor UO_605 (O_605,N_19996,N_19870);
xor UO_606 (O_606,N_19823,N_19943);
nand UO_607 (O_607,N_19854,N_19865);
nor UO_608 (O_608,N_19991,N_19994);
nor UO_609 (O_609,N_19845,N_19964);
nor UO_610 (O_610,N_19811,N_19976);
nor UO_611 (O_611,N_19848,N_19900);
and UO_612 (O_612,N_19945,N_19812);
xor UO_613 (O_613,N_19974,N_19821);
nor UO_614 (O_614,N_19910,N_19948);
and UO_615 (O_615,N_19832,N_19873);
nor UO_616 (O_616,N_19827,N_19866);
xnor UO_617 (O_617,N_19827,N_19953);
xor UO_618 (O_618,N_19848,N_19991);
nand UO_619 (O_619,N_19919,N_19852);
nor UO_620 (O_620,N_19907,N_19874);
xnor UO_621 (O_621,N_19962,N_19928);
and UO_622 (O_622,N_19956,N_19945);
xor UO_623 (O_623,N_19981,N_19950);
xor UO_624 (O_624,N_19840,N_19923);
nor UO_625 (O_625,N_19877,N_19802);
xor UO_626 (O_626,N_19984,N_19855);
nand UO_627 (O_627,N_19830,N_19984);
xnor UO_628 (O_628,N_19911,N_19976);
nand UO_629 (O_629,N_19965,N_19832);
and UO_630 (O_630,N_19866,N_19837);
xor UO_631 (O_631,N_19858,N_19895);
or UO_632 (O_632,N_19874,N_19876);
nand UO_633 (O_633,N_19820,N_19828);
xnor UO_634 (O_634,N_19972,N_19872);
or UO_635 (O_635,N_19856,N_19862);
nand UO_636 (O_636,N_19820,N_19832);
nand UO_637 (O_637,N_19958,N_19911);
and UO_638 (O_638,N_19983,N_19923);
nand UO_639 (O_639,N_19885,N_19973);
or UO_640 (O_640,N_19904,N_19830);
nor UO_641 (O_641,N_19907,N_19963);
nand UO_642 (O_642,N_19806,N_19933);
nor UO_643 (O_643,N_19939,N_19851);
and UO_644 (O_644,N_19960,N_19845);
xnor UO_645 (O_645,N_19875,N_19865);
xor UO_646 (O_646,N_19958,N_19886);
nand UO_647 (O_647,N_19920,N_19935);
or UO_648 (O_648,N_19827,N_19876);
or UO_649 (O_649,N_19866,N_19968);
and UO_650 (O_650,N_19876,N_19801);
xor UO_651 (O_651,N_19961,N_19923);
and UO_652 (O_652,N_19898,N_19863);
nor UO_653 (O_653,N_19915,N_19830);
xnor UO_654 (O_654,N_19838,N_19906);
nand UO_655 (O_655,N_19908,N_19996);
and UO_656 (O_656,N_19979,N_19880);
nand UO_657 (O_657,N_19803,N_19930);
nor UO_658 (O_658,N_19989,N_19998);
xnor UO_659 (O_659,N_19994,N_19870);
nor UO_660 (O_660,N_19890,N_19968);
nand UO_661 (O_661,N_19948,N_19932);
nand UO_662 (O_662,N_19980,N_19900);
xor UO_663 (O_663,N_19972,N_19823);
or UO_664 (O_664,N_19881,N_19968);
nor UO_665 (O_665,N_19960,N_19949);
xor UO_666 (O_666,N_19928,N_19923);
or UO_667 (O_667,N_19942,N_19803);
and UO_668 (O_668,N_19975,N_19878);
xnor UO_669 (O_669,N_19849,N_19964);
and UO_670 (O_670,N_19821,N_19817);
xor UO_671 (O_671,N_19897,N_19983);
or UO_672 (O_672,N_19910,N_19924);
nand UO_673 (O_673,N_19918,N_19944);
xor UO_674 (O_674,N_19909,N_19882);
nor UO_675 (O_675,N_19992,N_19970);
and UO_676 (O_676,N_19873,N_19865);
nand UO_677 (O_677,N_19932,N_19999);
xnor UO_678 (O_678,N_19950,N_19909);
or UO_679 (O_679,N_19918,N_19913);
or UO_680 (O_680,N_19983,N_19959);
and UO_681 (O_681,N_19947,N_19990);
nor UO_682 (O_682,N_19882,N_19831);
nor UO_683 (O_683,N_19978,N_19804);
and UO_684 (O_684,N_19891,N_19987);
and UO_685 (O_685,N_19950,N_19948);
and UO_686 (O_686,N_19941,N_19966);
nand UO_687 (O_687,N_19869,N_19857);
or UO_688 (O_688,N_19926,N_19857);
xor UO_689 (O_689,N_19910,N_19832);
nand UO_690 (O_690,N_19826,N_19863);
or UO_691 (O_691,N_19894,N_19882);
and UO_692 (O_692,N_19932,N_19905);
nand UO_693 (O_693,N_19829,N_19909);
nand UO_694 (O_694,N_19801,N_19981);
or UO_695 (O_695,N_19833,N_19877);
nor UO_696 (O_696,N_19987,N_19822);
or UO_697 (O_697,N_19876,N_19894);
nand UO_698 (O_698,N_19881,N_19839);
nor UO_699 (O_699,N_19823,N_19982);
nand UO_700 (O_700,N_19999,N_19939);
and UO_701 (O_701,N_19803,N_19969);
xnor UO_702 (O_702,N_19816,N_19838);
or UO_703 (O_703,N_19882,N_19854);
xnor UO_704 (O_704,N_19975,N_19889);
or UO_705 (O_705,N_19897,N_19887);
xor UO_706 (O_706,N_19977,N_19870);
nand UO_707 (O_707,N_19933,N_19950);
xnor UO_708 (O_708,N_19849,N_19895);
nand UO_709 (O_709,N_19895,N_19802);
xnor UO_710 (O_710,N_19952,N_19825);
xor UO_711 (O_711,N_19841,N_19974);
xor UO_712 (O_712,N_19837,N_19952);
xor UO_713 (O_713,N_19857,N_19852);
xor UO_714 (O_714,N_19952,N_19902);
or UO_715 (O_715,N_19875,N_19948);
or UO_716 (O_716,N_19822,N_19959);
nor UO_717 (O_717,N_19888,N_19956);
nor UO_718 (O_718,N_19874,N_19853);
nor UO_719 (O_719,N_19847,N_19828);
and UO_720 (O_720,N_19869,N_19964);
and UO_721 (O_721,N_19997,N_19888);
nand UO_722 (O_722,N_19841,N_19955);
nand UO_723 (O_723,N_19954,N_19909);
and UO_724 (O_724,N_19931,N_19915);
nor UO_725 (O_725,N_19947,N_19938);
or UO_726 (O_726,N_19940,N_19833);
or UO_727 (O_727,N_19826,N_19934);
nor UO_728 (O_728,N_19987,N_19961);
or UO_729 (O_729,N_19905,N_19846);
nand UO_730 (O_730,N_19942,N_19810);
nor UO_731 (O_731,N_19924,N_19869);
xnor UO_732 (O_732,N_19982,N_19849);
xor UO_733 (O_733,N_19945,N_19920);
xor UO_734 (O_734,N_19867,N_19972);
nor UO_735 (O_735,N_19973,N_19940);
xnor UO_736 (O_736,N_19888,N_19975);
xor UO_737 (O_737,N_19873,N_19925);
and UO_738 (O_738,N_19893,N_19999);
nand UO_739 (O_739,N_19853,N_19913);
and UO_740 (O_740,N_19914,N_19840);
and UO_741 (O_741,N_19886,N_19981);
nor UO_742 (O_742,N_19952,N_19836);
xor UO_743 (O_743,N_19874,N_19892);
xor UO_744 (O_744,N_19897,N_19813);
or UO_745 (O_745,N_19823,N_19951);
nand UO_746 (O_746,N_19868,N_19860);
and UO_747 (O_747,N_19948,N_19920);
or UO_748 (O_748,N_19812,N_19828);
or UO_749 (O_749,N_19950,N_19852);
and UO_750 (O_750,N_19891,N_19874);
and UO_751 (O_751,N_19885,N_19834);
nor UO_752 (O_752,N_19875,N_19826);
nand UO_753 (O_753,N_19833,N_19842);
xor UO_754 (O_754,N_19830,N_19827);
and UO_755 (O_755,N_19886,N_19858);
nor UO_756 (O_756,N_19989,N_19991);
xor UO_757 (O_757,N_19943,N_19835);
nor UO_758 (O_758,N_19847,N_19802);
or UO_759 (O_759,N_19974,N_19923);
nor UO_760 (O_760,N_19941,N_19880);
xor UO_761 (O_761,N_19920,N_19900);
nor UO_762 (O_762,N_19857,N_19970);
nand UO_763 (O_763,N_19923,N_19966);
nor UO_764 (O_764,N_19993,N_19999);
nand UO_765 (O_765,N_19982,N_19826);
nand UO_766 (O_766,N_19882,N_19906);
nor UO_767 (O_767,N_19809,N_19926);
or UO_768 (O_768,N_19806,N_19950);
nor UO_769 (O_769,N_19929,N_19830);
xor UO_770 (O_770,N_19851,N_19809);
nand UO_771 (O_771,N_19842,N_19967);
nor UO_772 (O_772,N_19804,N_19860);
xnor UO_773 (O_773,N_19962,N_19849);
or UO_774 (O_774,N_19910,N_19891);
or UO_775 (O_775,N_19977,N_19909);
and UO_776 (O_776,N_19844,N_19834);
or UO_777 (O_777,N_19980,N_19887);
and UO_778 (O_778,N_19911,N_19984);
nand UO_779 (O_779,N_19807,N_19951);
nor UO_780 (O_780,N_19820,N_19821);
and UO_781 (O_781,N_19958,N_19954);
and UO_782 (O_782,N_19926,N_19996);
nand UO_783 (O_783,N_19904,N_19901);
xor UO_784 (O_784,N_19863,N_19825);
nor UO_785 (O_785,N_19890,N_19843);
nand UO_786 (O_786,N_19831,N_19896);
or UO_787 (O_787,N_19936,N_19904);
xor UO_788 (O_788,N_19870,N_19927);
nand UO_789 (O_789,N_19894,N_19962);
xor UO_790 (O_790,N_19841,N_19888);
nor UO_791 (O_791,N_19937,N_19959);
and UO_792 (O_792,N_19822,N_19967);
nand UO_793 (O_793,N_19806,N_19837);
nor UO_794 (O_794,N_19956,N_19996);
or UO_795 (O_795,N_19862,N_19962);
xor UO_796 (O_796,N_19971,N_19961);
and UO_797 (O_797,N_19827,N_19938);
nand UO_798 (O_798,N_19893,N_19933);
nor UO_799 (O_799,N_19876,N_19859);
or UO_800 (O_800,N_19843,N_19948);
or UO_801 (O_801,N_19821,N_19853);
and UO_802 (O_802,N_19922,N_19965);
or UO_803 (O_803,N_19835,N_19954);
or UO_804 (O_804,N_19982,N_19846);
nor UO_805 (O_805,N_19863,N_19996);
xnor UO_806 (O_806,N_19928,N_19869);
or UO_807 (O_807,N_19869,N_19881);
nor UO_808 (O_808,N_19812,N_19925);
nor UO_809 (O_809,N_19972,N_19852);
xor UO_810 (O_810,N_19942,N_19887);
nand UO_811 (O_811,N_19808,N_19971);
or UO_812 (O_812,N_19994,N_19976);
xnor UO_813 (O_813,N_19916,N_19846);
nor UO_814 (O_814,N_19833,N_19926);
nor UO_815 (O_815,N_19864,N_19902);
or UO_816 (O_816,N_19803,N_19824);
or UO_817 (O_817,N_19902,N_19876);
or UO_818 (O_818,N_19897,N_19975);
nand UO_819 (O_819,N_19822,N_19907);
nand UO_820 (O_820,N_19837,N_19958);
or UO_821 (O_821,N_19802,N_19842);
nand UO_822 (O_822,N_19980,N_19898);
nand UO_823 (O_823,N_19916,N_19800);
nor UO_824 (O_824,N_19867,N_19997);
xor UO_825 (O_825,N_19966,N_19980);
xor UO_826 (O_826,N_19944,N_19969);
nand UO_827 (O_827,N_19978,N_19863);
nand UO_828 (O_828,N_19815,N_19947);
or UO_829 (O_829,N_19982,N_19868);
nor UO_830 (O_830,N_19844,N_19946);
nor UO_831 (O_831,N_19898,N_19930);
xnor UO_832 (O_832,N_19949,N_19859);
xor UO_833 (O_833,N_19925,N_19952);
and UO_834 (O_834,N_19862,N_19905);
and UO_835 (O_835,N_19895,N_19837);
nand UO_836 (O_836,N_19859,N_19968);
and UO_837 (O_837,N_19918,N_19997);
or UO_838 (O_838,N_19987,N_19904);
nor UO_839 (O_839,N_19907,N_19802);
nor UO_840 (O_840,N_19898,N_19884);
nor UO_841 (O_841,N_19836,N_19953);
nor UO_842 (O_842,N_19855,N_19860);
or UO_843 (O_843,N_19964,N_19930);
nor UO_844 (O_844,N_19856,N_19888);
and UO_845 (O_845,N_19844,N_19959);
or UO_846 (O_846,N_19866,N_19944);
and UO_847 (O_847,N_19974,N_19804);
xor UO_848 (O_848,N_19897,N_19965);
nand UO_849 (O_849,N_19960,N_19829);
or UO_850 (O_850,N_19850,N_19895);
xnor UO_851 (O_851,N_19998,N_19957);
or UO_852 (O_852,N_19881,N_19800);
and UO_853 (O_853,N_19894,N_19866);
and UO_854 (O_854,N_19823,N_19818);
nor UO_855 (O_855,N_19828,N_19884);
and UO_856 (O_856,N_19864,N_19982);
and UO_857 (O_857,N_19846,N_19973);
nand UO_858 (O_858,N_19809,N_19991);
xnor UO_859 (O_859,N_19971,N_19932);
nand UO_860 (O_860,N_19806,N_19815);
xor UO_861 (O_861,N_19948,N_19952);
nand UO_862 (O_862,N_19969,N_19800);
and UO_863 (O_863,N_19961,N_19947);
and UO_864 (O_864,N_19975,N_19992);
or UO_865 (O_865,N_19937,N_19893);
or UO_866 (O_866,N_19929,N_19811);
or UO_867 (O_867,N_19830,N_19848);
and UO_868 (O_868,N_19826,N_19808);
nand UO_869 (O_869,N_19961,N_19970);
nand UO_870 (O_870,N_19985,N_19971);
or UO_871 (O_871,N_19921,N_19815);
nand UO_872 (O_872,N_19882,N_19965);
nor UO_873 (O_873,N_19980,N_19942);
and UO_874 (O_874,N_19873,N_19902);
xor UO_875 (O_875,N_19914,N_19925);
nor UO_876 (O_876,N_19888,N_19905);
nor UO_877 (O_877,N_19834,N_19883);
and UO_878 (O_878,N_19940,N_19969);
and UO_879 (O_879,N_19818,N_19916);
and UO_880 (O_880,N_19912,N_19873);
nor UO_881 (O_881,N_19965,N_19836);
or UO_882 (O_882,N_19982,N_19818);
and UO_883 (O_883,N_19888,N_19973);
nand UO_884 (O_884,N_19992,N_19989);
or UO_885 (O_885,N_19801,N_19990);
and UO_886 (O_886,N_19816,N_19847);
and UO_887 (O_887,N_19843,N_19904);
xor UO_888 (O_888,N_19935,N_19963);
xnor UO_889 (O_889,N_19989,N_19913);
and UO_890 (O_890,N_19999,N_19984);
xor UO_891 (O_891,N_19874,N_19919);
or UO_892 (O_892,N_19893,N_19815);
nand UO_893 (O_893,N_19824,N_19856);
or UO_894 (O_894,N_19947,N_19978);
nor UO_895 (O_895,N_19904,N_19816);
nand UO_896 (O_896,N_19983,N_19990);
and UO_897 (O_897,N_19846,N_19909);
nor UO_898 (O_898,N_19984,N_19915);
or UO_899 (O_899,N_19927,N_19866);
nor UO_900 (O_900,N_19874,N_19831);
or UO_901 (O_901,N_19857,N_19989);
nand UO_902 (O_902,N_19830,N_19997);
nand UO_903 (O_903,N_19930,N_19957);
nor UO_904 (O_904,N_19856,N_19829);
nor UO_905 (O_905,N_19979,N_19925);
nand UO_906 (O_906,N_19915,N_19869);
or UO_907 (O_907,N_19895,N_19916);
nor UO_908 (O_908,N_19978,N_19995);
or UO_909 (O_909,N_19890,N_19879);
nor UO_910 (O_910,N_19858,N_19898);
or UO_911 (O_911,N_19948,N_19958);
xnor UO_912 (O_912,N_19899,N_19893);
nand UO_913 (O_913,N_19986,N_19808);
and UO_914 (O_914,N_19913,N_19968);
nor UO_915 (O_915,N_19868,N_19941);
nand UO_916 (O_916,N_19875,N_19850);
xor UO_917 (O_917,N_19885,N_19856);
xnor UO_918 (O_918,N_19950,N_19949);
or UO_919 (O_919,N_19991,N_19877);
and UO_920 (O_920,N_19800,N_19960);
nor UO_921 (O_921,N_19976,N_19832);
nor UO_922 (O_922,N_19992,N_19872);
nand UO_923 (O_923,N_19877,N_19914);
nand UO_924 (O_924,N_19937,N_19866);
xnor UO_925 (O_925,N_19809,N_19869);
or UO_926 (O_926,N_19994,N_19886);
nand UO_927 (O_927,N_19995,N_19971);
nand UO_928 (O_928,N_19952,N_19817);
and UO_929 (O_929,N_19911,N_19879);
nor UO_930 (O_930,N_19937,N_19855);
xnor UO_931 (O_931,N_19981,N_19952);
and UO_932 (O_932,N_19874,N_19950);
nand UO_933 (O_933,N_19858,N_19892);
xnor UO_934 (O_934,N_19943,N_19870);
or UO_935 (O_935,N_19908,N_19807);
or UO_936 (O_936,N_19965,N_19847);
or UO_937 (O_937,N_19943,N_19928);
and UO_938 (O_938,N_19903,N_19831);
and UO_939 (O_939,N_19950,N_19958);
or UO_940 (O_940,N_19849,N_19942);
nand UO_941 (O_941,N_19938,N_19940);
nand UO_942 (O_942,N_19967,N_19958);
and UO_943 (O_943,N_19996,N_19838);
nand UO_944 (O_944,N_19958,N_19878);
and UO_945 (O_945,N_19996,N_19856);
nand UO_946 (O_946,N_19952,N_19845);
xor UO_947 (O_947,N_19920,N_19878);
or UO_948 (O_948,N_19955,N_19821);
and UO_949 (O_949,N_19995,N_19857);
or UO_950 (O_950,N_19846,N_19825);
nand UO_951 (O_951,N_19997,N_19850);
or UO_952 (O_952,N_19884,N_19890);
or UO_953 (O_953,N_19930,N_19888);
nand UO_954 (O_954,N_19874,N_19936);
or UO_955 (O_955,N_19862,N_19809);
and UO_956 (O_956,N_19957,N_19910);
or UO_957 (O_957,N_19919,N_19855);
or UO_958 (O_958,N_19940,N_19870);
or UO_959 (O_959,N_19986,N_19944);
xor UO_960 (O_960,N_19891,N_19819);
nand UO_961 (O_961,N_19942,N_19976);
nor UO_962 (O_962,N_19951,N_19972);
and UO_963 (O_963,N_19924,N_19828);
or UO_964 (O_964,N_19863,N_19955);
and UO_965 (O_965,N_19942,N_19884);
nand UO_966 (O_966,N_19992,N_19843);
xnor UO_967 (O_967,N_19939,N_19919);
nand UO_968 (O_968,N_19803,N_19960);
nand UO_969 (O_969,N_19875,N_19986);
nand UO_970 (O_970,N_19967,N_19891);
xor UO_971 (O_971,N_19997,N_19892);
xnor UO_972 (O_972,N_19811,N_19818);
nand UO_973 (O_973,N_19942,N_19970);
nor UO_974 (O_974,N_19974,N_19846);
and UO_975 (O_975,N_19915,N_19919);
nor UO_976 (O_976,N_19817,N_19980);
nor UO_977 (O_977,N_19903,N_19833);
nand UO_978 (O_978,N_19992,N_19956);
nand UO_979 (O_979,N_19924,N_19843);
xor UO_980 (O_980,N_19974,N_19922);
nor UO_981 (O_981,N_19977,N_19950);
nand UO_982 (O_982,N_19996,N_19959);
xor UO_983 (O_983,N_19933,N_19890);
and UO_984 (O_984,N_19811,N_19820);
xnor UO_985 (O_985,N_19924,N_19949);
nand UO_986 (O_986,N_19876,N_19916);
nor UO_987 (O_987,N_19942,N_19908);
xnor UO_988 (O_988,N_19937,N_19993);
xor UO_989 (O_989,N_19998,N_19954);
nor UO_990 (O_990,N_19875,N_19914);
or UO_991 (O_991,N_19929,N_19939);
or UO_992 (O_992,N_19978,N_19891);
nor UO_993 (O_993,N_19914,N_19906);
nor UO_994 (O_994,N_19890,N_19995);
or UO_995 (O_995,N_19950,N_19916);
or UO_996 (O_996,N_19976,N_19845);
xnor UO_997 (O_997,N_19940,N_19945);
xnor UO_998 (O_998,N_19897,N_19918);
or UO_999 (O_999,N_19871,N_19816);
nor UO_1000 (O_1000,N_19933,N_19981);
xnor UO_1001 (O_1001,N_19998,N_19854);
nor UO_1002 (O_1002,N_19970,N_19989);
nand UO_1003 (O_1003,N_19901,N_19877);
xor UO_1004 (O_1004,N_19816,N_19859);
nor UO_1005 (O_1005,N_19926,N_19925);
or UO_1006 (O_1006,N_19990,N_19991);
or UO_1007 (O_1007,N_19950,N_19920);
xor UO_1008 (O_1008,N_19981,N_19804);
and UO_1009 (O_1009,N_19945,N_19908);
and UO_1010 (O_1010,N_19809,N_19942);
nand UO_1011 (O_1011,N_19886,N_19868);
xor UO_1012 (O_1012,N_19972,N_19893);
or UO_1013 (O_1013,N_19929,N_19842);
xnor UO_1014 (O_1014,N_19839,N_19989);
nand UO_1015 (O_1015,N_19973,N_19906);
or UO_1016 (O_1016,N_19968,N_19905);
and UO_1017 (O_1017,N_19889,N_19902);
or UO_1018 (O_1018,N_19916,N_19967);
nand UO_1019 (O_1019,N_19892,N_19982);
nor UO_1020 (O_1020,N_19860,N_19905);
nand UO_1021 (O_1021,N_19913,N_19969);
nor UO_1022 (O_1022,N_19968,N_19897);
and UO_1023 (O_1023,N_19934,N_19999);
xnor UO_1024 (O_1024,N_19879,N_19883);
xnor UO_1025 (O_1025,N_19904,N_19892);
xnor UO_1026 (O_1026,N_19940,N_19977);
xnor UO_1027 (O_1027,N_19896,N_19964);
nand UO_1028 (O_1028,N_19818,N_19887);
xor UO_1029 (O_1029,N_19877,N_19955);
and UO_1030 (O_1030,N_19895,N_19871);
or UO_1031 (O_1031,N_19841,N_19883);
or UO_1032 (O_1032,N_19921,N_19879);
nor UO_1033 (O_1033,N_19999,N_19898);
nor UO_1034 (O_1034,N_19831,N_19814);
nor UO_1035 (O_1035,N_19845,N_19840);
or UO_1036 (O_1036,N_19959,N_19816);
xnor UO_1037 (O_1037,N_19895,N_19879);
and UO_1038 (O_1038,N_19982,N_19874);
nor UO_1039 (O_1039,N_19908,N_19926);
or UO_1040 (O_1040,N_19932,N_19936);
and UO_1041 (O_1041,N_19986,N_19976);
nor UO_1042 (O_1042,N_19853,N_19942);
nand UO_1043 (O_1043,N_19800,N_19875);
and UO_1044 (O_1044,N_19825,N_19982);
nand UO_1045 (O_1045,N_19979,N_19900);
nor UO_1046 (O_1046,N_19993,N_19883);
xor UO_1047 (O_1047,N_19986,N_19853);
or UO_1048 (O_1048,N_19863,N_19959);
nor UO_1049 (O_1049,N_19983,N_19882);
xor UO_1050 (O_1050,N_19889,N_19856);
xor UO_1051 (O_1051,N_19995,N_19951);
and UO_1052 (O_1052,N_19884,N_19955);
xor UO_1053 (O_1053,N_19872,N_19937);
nand UO_1054 (O_1054,N_19834,N_19856);
or UO_1055 (O_1055,N_19840,N_19992);
xnor UO_1056 (O_1056,N_19913,N_19864);
nand UO_1057 (O_1057,N_19843,N_19968);
and UO_1058 (O_1058,N_19834,N_19912);
nand UO_1059 (O_1059,N_19833,N_19880);
xnor UO_1060 (O_1060,N_19940,N_19898);
nor UO_1061 (O_1061,N_19805,N_19917);
xor UO_1062 (O_1062,N_19884,N_19810);
nand UO_1063 (O_1063,N_19929,N_19949);
xnor UO_1064 (O_1064,N_19867,N_19981);
nand UO_1065 (O_1065,N_19883,N_19973);
or UO_1066 (O_1066,N_19894,N_19936);
and UO_1067 (O_1067,N_19827,N_19803);
xnor UO_1068 (O_1068,N_19951,N_19897);
nand UO_1069 (O_1069,N_19994,N_19917);
xor UO_1070 (O_1070,N_19861,N_19908);
xnor UO_1071 (O_1071,N_19864,N_19825);
nand UO_1072 (O_1072,N_19819,N_19847);
xnor UO_1073 (O_1073,N_19865,N_19989);
and UO_1074 (O_1074,N_19905,N_19845);
nand UO_1075 (O_1075,N_19924,N_19926);
or UO_1076 (O_1076,N_19893,N_19801);
and UO_1077 (O_1077,N_19891,N_19928);
nand UO_1078 (O_1078,N_19996,N_19907);
or UO_1079 (O_1079,N_19962,N_19948);
nor UO_1080 (O_1080,N_19825,N_19958);
or UO_1081 (O_1081,N_19871,N_19802);
and UO_1082 (O_1082,N_19801,N_19925);
nor UO_1083 (O_1083,N_19957,N_19862);
nor UO_1084 (O_1084,N_19930,N_19842);
nand UO_1085 (O_1085,N_19883,N_19994);
xor UO_1086 (O_1086,N_19972,N_19895);
or UO_1087 (O_1087,N_19941,N_19861);
and UO_1088 (O_1088,N_19814,N_19837);
nor UO_1089 (O_1089,N_19943,N_19967);
xor UO_1090 (O_1090,N_19946,N_19846);
nor UO_1091 (O_1091,N_19812,N_19821);
nand UO_1092 (O_1092,N_19908,N_19803);
nor UO_1093 (O_1093,N_19826,N_19879);
nand UO_1094 (O_1094,N_19837,N_19823);
nor UO_1095 (O_1095,N_19925,N_19981);
and UO_1096 (O_1096,N_19868,N_19931);
xnor UO_1097 (O_1097,N_19856,N_19960);
nor UO_1098 (O_1098,N_19900,N_19833);
nor UO_1099 (O_1099,N_19959,N_19951);
and UO_1100 (O_1100,N_19801,N_19888);
nand UO_1101 (O_1101,N_19950,N_19878);
xor UO_1102 (O_1102,N_19848,N_19888);
or UO_1103 (O_1103,N_19960,N_19917);
nand UO_1104 (O_1104,N_19866,N_19959);
and UO_1105 (O_1105,N_19973,N_19842);
nor UO_1106 (O_1106,N_19858,N_19830);
or UO_1107 (O_1107,N_19873,N_19893);
or UO_1108 (O_1108,N_19953,N_19943);
and UO_1109 (O_1109,N_19864,N_19917);
nand UO_1110 (O_1110,N_19804,N_19910);
or UO_1111 (O_1111,N_19910,N_19929);
or UO_1112 (O_1112,N_19879,N_19967);
nand UO_1113 (O_1113,N_19830,N_19861);
xor UO_1114 (O_1114,N_19863,N_19870);
nand UO_1115 (O_1115,N_19918,N_19952);
or UO_1116 (O_1116,N_19984,N_19868);
xnor UO_1117 (O_1117,N_19983,N_19849);
nand UO_1118 (O_1118,N_19992,N_19991);
xnor UO_1119 (O_1119,N_19880,N_19858);
xor UO_1120 (O_1120,N_19975,N_19905);
and UO_1121 (O_1121,N_19877,N_19852);
and UO_1122 (O_1122,N_19852,N_19853);
xnor UO_1123 (O_1123,N_19826,N_19938);
xor UO_1124 (O_1124,N_19864,N_19827);
and UO_1125 (O_1125,N_19882,N_19988);
or UO_1126 (O_1126,N_19901,N_19820);
or UO_1127 (O_1127,N_19863,N_19916);
nand UO_1128 (O_1128,N_19968,N_19999);
and UO_1129 (O_1129,N_19823,N_19980);
and UO_1130 (O_1130,N_19946,N_19937);
nor UO_1131 (O_1131,N_19967,N_19830);
xor UO_1132 (O_1132,N_19913,N_19862);
or UO_1133 (O_1133,N_19994,N_19937);
nor UO_1134 (O_1134,N_19892,N_19912);
xnor UO_1135 (O_1135,N_19968,N_19834);
and UO_1136 (O_1136,N_19870,N_19938);
xnor UO_1137 (O_1137,N_19844,N_19929);
or UO_1138 (O_1138,N_19898,N_19827);
or UO_1139 (O_1139,N_19901,N_19825);
nor UO_1140 (O_1140,N_19862,N_19992);
and UO_1141 (O_1141,N_19828,N_19949);
and UO_1142 (O_1142,N_19846,N_19945);
and UO_1143 (O_1143,N_19911,N_19828);
or UO_1144 (O_1144,N_19971,N_19978);
nand UO_1145 (O_1145,N_19977,N_19813);
nor UO_1146 (O_1146,N_19989,N_19804);
and UO_1147 (O_1147,N_19875,N_19808);
and UO_1148 (O_1148,N_19826,N_19957);
xor UO_1149 (O_1149,N_19877,N_19936);
or UO_1150 (O_1150,N_19899,N_19929);
nor UO_1151 (O_1151,N_19963,N_19906);
xor UO_1152 (O_1152,N_19912,N_19876);
or UO_1153 (O_1153,N_19933,N_19984);
xor UO_1154 (O_1154,N_19913,N_19994);
and UO_1155 (O_1155,N_19838,N_19860);
nor UO_1156 (O_1156,N_19975,N_19942);
xor UO_1157 (O_1157,N_19897,N_19960);
nand UO_1158 (O_1158,N_19987,N_19844);
or UO_1159 (O_1159,N_19836,N_19998);
xnor UO_1160 (O_1160,N_19969,N_19921);
and UO_1161 (O_1161,N_19800,N_19913);
xor UO_1162 (O_1162,N_19965,N_19991);
xnor UO_1163 (O_1163,N_19805,N_19997);
nand UO_1164 (O_1164,N_19871,N_19927);
nor UO_1165 (O_1165,N_19986,N_19991);
nor UO_1166 (O_1166,N_19883,N_19997);
nor UO_1167 (O_1167,N_19987,N_19927);
or UO_1168 (O_1168,N_19826,N_19832);
nor UO_1169 (O_1169,N_19873,N_19907);
nand UO_1170 (O_1170,N_19806,N_19875);
nand UO_1171 (O_1171,N_19857,N_19820);
and UO_1172 (O_1172,N_19899,N_19831);
or UO_1173 (O_1173,N_19812,N_19871);
or UO_1174 (O_1174,N_19968,N_19891);
nand UO_1175 (O_1175,N_19900,N_19964);
or UO_1176 (O_1176,N_19968,N_19857);
xnor UO_1177 (O_1177,N_19816,N_19802);
nand UO_1178 (O_1178,N_19964,N_19898);
xnor UO_1179 (O_1179,N_19945,N_19892);
xnor UO_1180 (O_1180,N_19929,N_19859);
nor UO_1181 (O_1181,N_19826,N_19873);
xor UO_1182 (O_1182,N_19953,N_19873);
and UO_1183 (O_1183,N_19810,N_19902);
or UO_1184 (O_1184,N_19826,N_19853);
nand UO_1185 (O_1185,N_19946,N_19932);
and UO_1186 (O_1186,N_19926,N_19800);
and UO_1187 (O_1187,N_19847,N_19893);
or UO_1188 (O_1188,N_19896,N_19951);
nor UO_1189 (O_1189,N_19997,N_19885);
or UO_1190 (O_1190,N_19979,N_19968);
and UO_1191 (O_1191,N_19819,N_19937);
xor UO_1192 (O_1192,N_19841,N_19806);
and UO_1193 (O_1193,N_19992,N_19922);
and UO_1194 (O_1194,N_19975,N_19901);
nor UO_1195 (O_1195,N_19866,N_19863);
xnor UO_1196 (O_1196,N_19990,N_19913);
nand UO_1197 (O_1197,N_19815,N_19967);
or UO_1198 (O_1198,N_19950,N_19893);
xnor UO_1199 (O_1199,N_19901,N_19882);
xor UO_1200 (O_1200,N_19927,N_19832);
and UO_1201 (O_1201,N_19914,N_19874);
nand UO_1202 (O_1202,N_19803,N_19818);
and UO_1203 (O_1203,N_19961,N_19807);
and UO_1204 (O_1204,N_19985,N_19833);
nand UO_1205 (O_1205,N_19847,N_19848);
nand UO_1206 (O_1206,N_19859,N_19918);
nand UO_1207 (O_1207,N_19961,N_19829);
or UO_1208 (O_1208,N_19884,N_19853);
nand UO_1209 (O_1209,N_19861,N_19968);
nor UO_1210 (O_1210,N_19850,N_19897);
or UO_1211 (O_1211,N_19984,N_19847);
nand UO_1212 (O_1212,N_19962,N_19877);
or UO_1213 (O_1213,N_19814,N_19970);
nand UO_1214 (O_1214,N_19805,N_19896);
nand UO_1215 (O_1215,N_19833,N_19947);
nand UO_1216 (O_1216,N_19962,N_19899);
nand UO_1217 (O_1217,N_19808,N_19824);
xor UO_1218 (O_1218,N_19929,N_19884);
nand UO_1219 (O_1219,N_19890,N_19974);
or UO_1220 (O_1220,N_19986,N_19950);
nand UO_1221 (O_1221,N_19803,N_19919);
nand UO_1222 (O_1222,N_19831,N_19961);
nand UO_1223 (O_1223,N_19844,N_19982);
xor UO_1224 (O_1224,N_19970,N_19835);
nand UO_1225 (O_1225,N_19911,N_19900);
xor UO_1226 (O_1226,N_19890,N_19887);
or UO_1227 (O_1227,N_19919,N_19931);
nand UO_1228 (O_1228,N_19973,N_19818);
xor UO_1229 (O_1229,N_19847,N_19869);
and UO_1230 (O_1230,N_19838,N_19971);
and UO_1231 (O_1231,N_19852,N_19933);
xor UO_1232 (O_1232,N_19937,N_19815);
or UO_1233 (O_1233,N_19813,N_19802);
or UO_1234 (O_1234,N_19976,N_19837);
or UO_1235 (O_1235,N_19956,N_19931);
nand UO_1236 (O_1236,N_19925,N_19842);
and UO_1237 (O_1237,N_19943,N_19897);
nor UO_1238 (O_1238,N_19908,N_19912);
nand UO_1239 (O_1239,N_19842,N_19836);
or UO_1240 (O_1240,N_19950,N_19834);
or UO_1241 (O_1241,N_19992,N_19867);
and UO_1242 (O_1242,N_19850,N_19970);
and UO_1243 (O_1243,N_19976,N_19945);
and UO_1244 (O_1244,N_19990,N_19988);
and UO_1245 (O_1245,N_19903,N_19951);
nand UO_1246 (O_1246,N_19970,N_19858);
nand UO_1247 (O_1247,N_19924,N_19868);
nor UO_1248 (O_1248,N_19948,N_19916);
nand UO_1249 (O_1249,N_19835,N_19960);
xnor UO_1250 (O_1250,N_19957,N_19831);
or UO_1251 (O_1251,N_19931,N_19854);
and UO_1252 (O_1252,N_19940,N_19876);
xnor UO_1253 (O_1253,N_19844,N_19839);
xnor UO_1254 (O_1254,N_19978,N_19830);
nand UO_1255 (O_1255,N_19892,N_19802);
nand UO_1256 (O_1256,N_19854,N_19859);
and UO_1257 (O_1257,N_19871,N_19830);
or UO_1258 (O_1258,N_19969,N_19942);
or UO_1259 (O_1259,N_19937,N_19991);
nor UO_1260 (O_1260,N_19873,N_19994);
xor UO_1261 (O_1261,N_19842,N_19878);
nor UO_1262 (O_1262,N_19901,N_19878);
and UO_1263 (O_1263,N_19874,N_19823);
and UO_1264 (O_1264,N_19977,N_19941);
or UO_1265 (O_1265,N_19874,N_19992);
or UO_1266 (O_1266,N_19912,N_19801);
xor UO_1267 (O_1267,N_19996,N_19979);
nand UO_1268 (O_1268,N_19979,N_19876);
nor UO_1269 (O_1269,N_19807,N_19952);
nand UO_1270 (O_1270,N_19838,N_19899);
xnor UO_1271 (O_1271,N_19805,N_19941);
and UO_1272 (O_1272,N_19928,N_19807);
nand UO_1273 (O_1273,N_19943,N_19896);
and UO_1274 (O_1274,N_19910,N_19927);
nor UO_1275 (O_1275,N_19888,N_19916);
and UO_1276 (O_1276,N_19804,N_19850);
and UO_1277 (O_1277,N_19858,N_19855);
xor UO_1278 (O_1278,N_19883,N_19813);
or UO_1279 (O_1279,N_19932,N_19881);
and UO_1280 (O_1280,N_19902,N_19985);
xor UO_1281 (O_1281,N_19908,N_19983);
and UO_1282 (O_1282,N_19921,N_19895);
or UO_1283 (O_1283,N_19812,N_19985);
nor UO_1284 (O_1284,N_19906,N_19832);
xor UO_1285 (O_1285,N_19885,N_19913);
nor UO_1286 (O_1286,N_19952,N_19889);
nand UO_1287 (O_1287,N_19984,N_19998);
nor UO_1288 (O_1288,N_19835,N_19988);
nor UO_1289 (O_1289,N_19937,N_19878);
or UO_1290 (O_1290,N_19942,N_19918);
nand UO_1291 (O_1291,N_19989,N_19864);
and UO_1292 (O_1292,N_19866,N_19931);
nor UO_1293 (O_1293,N_19911,N_19808);
xnor UO_1294 (O_1294,N_19919,N_19963);
and UO_1295 (O_1295,N_19830,N_19981);
xnor UO_1296 (O_1296,N_19897,N_19898);
xor UO_1297 (O_1297,N_19962,N_19918);
and UO_1298 (O_1298,N_19978,N_19904);
nor UO_1299 (O_1299,N_19837,N_19876);
nand UO_1300 (O_1300,N_19878,N_19823);
nor UO_1301 (O_1301,N_19970,N_19822);
nand UO_1302 (O_1302,N_19910,N_19920);
nand UO_1303 (O_1303,N_19981,N_19993);
xor UO_1304 (O_1304,N_19856,N_19920);
nor UO_1305 (O_1305,N_19948,N_19805);
nand UO_1306 (O_1306,N_19863,N_19874);
nor UO_1307 (O_1307,N_19955,N_19934);
xnor UO_1308 (O_1308,N_19835,N_19884);
xnor UO_1309 (O_1309,N_19906,N_19934);
or UO_1310 (O_1310,N_19872,N_19977);
and UO_1311 (O_1311,N_19947,N_19930);
or UO_1312 (O_1312,N_19893,N_19870);
nand UO_1313 (O_1313,N_19814,N_19816);
and UO_1314 (O_1314,N_19931,N_19821);
xnor UO_1315 (O_1315,N_19863,N_19940);
nor UO_1316 (O_1316,N_19842,N_19916);
or UO_1317 (O_1317,N_19844,N_19824);
and UO_1318 (O_1318,N_19965,N_19946);
xor UO_1319 (O_1319,N_19862,N_19830);
or UO_1320 (O_1320,N_19908,N_19864);
nor UO_1321 (O_1321,N_19949,N_19809);
nor UO_1322 (O_1322,N_19816,N_19880);
xor UO_1323 (O_1323,N_19963,N_19800);
nor UO_1324 (O_1324,N_19847,N_19952);
nor UO_1325 (O_1325,N_19977,N_19857);
and UO_1326 (O_1326,N_19962,N_19940);
or UO_1327 (O_1327,N_19912,N_19956);
nor UO_1328 (O_1328,N_19929,N_19927);
nand UO_1329 (O_1329,N_19892,N_19827);
and UO_1330 (O_1330,N_19862,N_19951);
or UO_1331 (O_1331,N_19939,N_19893);
nor UO_1332 (O_1332,N_19933,N_19886);
or UO_1333 (O_1333,N_19993,N_19885);
nor UO_1334 (O_1334,N_19824,N_19931);
nand UO_1335 (O_1335,N_19984,N_19914);
xor UO_1336 (O_1336,N_19965,N_19853);
and UO_1337 (O_1337,N_19855,N_19989);
xor UO_1338 (O_1338,N_19993,N_19987);
xor UO_1339 (O_1339,N_19895,N_19833);
nand UO_1340 (O_1340,N_19815,N_19909);
xor UO_1341 (O_1341,N_19880,N_19831);
nor UO_1342 (O_1342,N_19891,N_19979);
nand UO_1343 (O_1343,N_19919,N_19971);
xnor UO_1344 (O_1344,N_19914,N_19975);
nor UO_1345 (O_1345,N_19986,N_19901);
and UO_1346 (O_1346,N_19850,N_19868);
nor UO_1347 (O_1347,N_19904,N_19992);
nor UO_1348 (O_1348,N_19923,N_19986);
nor UO_1349 (O_1349,N_19914,N_19960);
or UO_1350 (O_1350,N_19958,N_19876);
nand UO_1351 (O_1351,N_19978,N_19950);
nor UO_1352 (O_1352,N_19897,N_19982);
xnor UO_1353 (O_1353,N_19881,N_19885);
nand UO_1354 (O_1354,N_19832,N_19988);
nand UO_1355 (O_1355,N_19865,N_19905);
xnor UO_1356 (O_1356,N_19892,N_19833);
and UO_1357 (O_1357,N_19870,N_19905);
or UO_1358 (O_1358,N_19951,N_19871);
nand UO_1359 (O_1359,N_19928,N_19940);
xnor UO_1360 (O_1360,N_19902,N_19931);
xnor UO_1361 (O_1361,N_19925,N_19936);
and UO_1362 (O_1362,N_19944,N_19924);
xor UO_1363 (O_1363,N_19859,N_19917);
xnor UO_1364 (O_1364,N_19819,N_19920);
and UO_1365 (O_1365,N_19924,N_19821);
nand UO_1366 (O_1366,N_19972,N_19936);
xnor UO_1367 (O_1367,N_19978,N_19817);
xor UO_1368 (O_1368,N_19839,N_19820);
nor UO_1369 (O_1369,N_19983,N_19986);
xor UO_1370 (O_1370,N_19834,N_19855);
or UO_1371 (O_1371,N_19836,N_19814);
and UO_1372 (O_1372,N_19954,N_19846);
nand UO_1373 (O_1373,N_19812,N_19907);
nand UO_1374 (O_1374,N_19855,N_19890);
xnor UO_1375 (O_1375,N_19945,N_19901);
and UO_1376 (O_1376,N_19921,N_19926);
and UO_1377 (O_1377,N_19920,N_19880);
nor UO_1378 (O_1378,N_19980,N_19935);
and UO_1379 (O_1379,N_19985,N_19835);
nand UO_1380 (O_1380,N_19971,N_19937);
or UO_1381 (O_1381,N_19934,N_19914);
nand UO_1382 (O_1382,N_19994,N_19918);
or UO_1383 (O_1383,N_19909,N_19843);
nor UO_1384 (O_1384,N_19937,N_19883);
xnor UO_1385 (O_1385,N_19860,N_19951);
and UO_1386 (O_1386,N_19887,N_19845);
xnor UO_1387 (O_1387,N_19931,N_19888);
nand UO_1388 (O_1388,N_19990,N_19848);
or UO_1389 (O_1389,N_19867,N_19832);
xnor UO_1390 (O_1390,N_19871,N_19809);
xor UO_1391 (O_1391,N_19977,N_19874);
and UO_1392 (O_1392,N_19992,N_19949);
nor UO_1393 (O_1393,N_19964,N_19815);
and UO_1394 (O_1394,N_19921,N_19909);
nor UO_1395 (O_1395,N_19924,N_19922);
nor UO_1396 (O_1396,N_19943,N_19882);
nor UO_1397 (O_1397,N_19948,N_19989);
nor UO_1398 (O_1398,N_19820,N_19892);
nand UO_1399 (O_1399,N_19889,N_19949);
nand UO_1400 (O_1400,N_19849,N_19845);
nand UO_1401 (O_1401,N_19946,N_19980);
xnor UO_1402 (O_1402,N_19848,N_19853);
xnor UO_1403 (O_1403,N_19859,N_19955);
and UO_1404 (O_1404,N_19954,N_19947);
or UO_1405 (O_1405,N_19831,N_19883);
nor UO_1406 (O_1406,N_19974,N_19956);
nand UO_1407 (O_1407,N_19854,N_19871);
nor UO_1408 (O_1408,N_19928,N_19811);
or UO_1409 (O_1409,N_19868,N_19990);
or UO_1410 (O_1410,N_19893,N_19814);
xnor UO_1411 (O_1411,N_19967,N_19801);
xor UO_1412 (O_1412,N_19821,N_19937);
and UO_1413 (O_1413,N_19886,N_19845);
or UO_1414 (O_1414,N_19806,N_19843);
xnor UO_1415 (O_1415,N_19917,N_19895);
nand UO_1416 (O_1416,N_19984,N_19949);
nand UO_1417 (O_1417,N_19991,N_19806);
xnor UO_1418 (O_1418,N_19806,N_19819);
nand UO_1419 (O_1419,N_19816,N_19984);
nor UO_1420 (O_1420,N_19838,N_19803);
nor UO_1421 (O_1421,N_19971,N_19939);
nor UO_1422 (O_1422,N_19909,N_19842);
and UO_1423 (O_1423,N_19932,N_19817);
or UO_1424 (O_1424,N_19886,N_19969);
or UO_1425 (O_1425,N_19858,N_19807);
and UO_1426 (O_1426,N_19953,N_19946);
nand UO_1427 (O_1427,N_19993,N_19909);
or UO_1428 (O_1428,N_19870,N_19823);
nor UO_1429 (O_1429,N_19847,N_19829);
xnor UO_1430 (O_1430,N_19804,N_19904);
or UO_1431 (O_1431,N_19800,N_19948);
nor UO_1432 (O_1432,N_19841,N_19801);
and UO_1433 (O_1433,N_19909,N_19861);
and UO_1434 (O_1434,N_19891,N_19888);
nand UO_1435 (O_1435,N_19843,N_19944);
nand UO_1436 (O_1436,N_19914,N_19921);
nor UO_1437 (O_1437,N_19857,N_19901);
nand UO_1438 (O_1438,N_19977,N_19906);
nand UO_1439 (O_1439,N_19988,N_19923);
xnor UO_1440 (O_1440,N_19841,N_19824);
nand UO_1441 (O_1441,N_19881,N_19904);
xnor UO_1442 (O_1442,N_19873,N_19936);
nor UO_1443 (O_1443,N_19893,N_19856);
or UO_1444 (O_1444,N_19861,N_19900);
or UO_1445 (O_1445,N_19817,N_19967);
xnor UO_1446 (O_1446,N_19967,N_19912);
nand UO_1447 (O_1447,N_19842,N_19807);
nand UO_1448 (O_1448,N_19883,N_19809);
or UO_1449 (O_1449,N_19910,N_19907);
nand UO_1450 (O_1450,N_19924,N_19816);
xor UO_1451 (O_1451,N_19822,N_19838);
xnor UO_1452 (O_1452,N_19945,N_19883);
or UO_1453 (O_1453,N_19807,N_19840);
nand UO_1454 (O_1454,N_19899,N_19854);
xor UO_1455 (O_1455,N_19885,N_19860);
or UO_1456 (O_1456,N_19862,N_19929);
nand UO_1457 (O_1457,N_19842,N_19934);
or UO_1458 (O_1458,N_19820,N_19924);
or UO_1459 (O_1459,N_19970,N_19810);
xnor UO_1460 (O_1460,N_19901,N_19938);
nand UO_1461 (O_1461,N_19975,N_19916);
or UO_1462 (O_1462,N_19888,N_19870);
and UO_1463 (O_1463,N_19965,N_19909);
and UO_1464 (O_1464,N_19920,N_19965);
and UO_1465 (O_1465,N_19966,N_19807);
and UO_1466 (O_1466,N_19869,N_19842);
or UO_1467 (O_1467,N_19923,N_19898);
or UO_1468 (O_1468,N_19990,N_19936);
and UO_1469 (O_1469,N_19901,N_19897);
and UO_1470 (O_1470,N_19862,N_19834);
or UO_1471 (O_1471,N_19819,N_19898);
nor UO_1472 (O_1472,N_19886,N_19819);
nand UO_1473 (O_1473,N_19911,N_19805);
nor UO_1474 (O_1474,N_19929,N_19835);
or UO_1475 (O_1475,N_19920,N_19991);
nand UO_1476 (O_1476,N_19937,N_19931);
and UO_1477 (O_1477,N_19837,N_19803);
or UO_1478 (O_1478,N_19878,N_19815);
nor UO_1479 (O_1479,N_19855,N_19817);
xnor UO_1480 (O_1480,N_19957,N_19948);
or UO_1481 (O_1481,N_19805,N_19842);
xor UO_1482 (O_1482,N_19819,N_19868);
nor UO_1483 (O_1483,N_19901,N_19898);
xor UO_1484 (O_1484,N_19830,N_19867);
nand UO_1485 (O_1485,N_19863,N_19903);
and UO_1486 (O_1486,N_19946,N_19899);
and UO_1487 (O_1487,N_19869,N_19980);
and UO_1488 (O_1488,N_19906,N_19989);
nor UO_1489 (O_1489,N_19873,N_19858);
nand UO_1490 (O_1490,N_19847,N_19937);
nor UO_1491 (O_1491,N_19866,N_19836);
and UO_1492 (O_1492,N_19867,N_19929);
or UO_1493 (O_1493,N_19918,N_19839);
nand UO_1494 (O_1494,N_19842,N_19921);
nand UO_1495 (O_1495,N_19814,N_19862);
nand UO_1496 (O_1496,N_19840,N_19882);
and UO_1497 (O_1497,N_19903,N_19959);
xnor UO_1498 (O_1498,N_19956,N_19930);
or UO_1499 (O_1499,N_19956,N_19921);
nor UO_1500 (O_1500,N_19974,N_19966);
nand UO_1501 (O_1501,N_19856,N_19850);
xor UO_1502 (O_1502,N_19957,N_19877);
or UO_1503 (O_1503,N_19964,N_19979);
nand UO_1504 (O_1504,N_19866,N_19822);
and UO_1505 (O_1505,N_19896,N_19819);
nor UO_1506 (O_1506,N_19852,N_19855);
nand UO_1507 (O_1507,N_19906,N_19875);
and UO_1508 (O_1508,N_19935,N_19834);
nand UO_1509 (O_1509,N_19853,N_19878);
xor UO_1510 (O_1510,N_19985,N_19931);
nand UO_1511 (O_1511,N_19866,N_19844);
nor UO_1512 (O_1512,N_19829,N_19963);
nor UO_1513 (O_1513,N_19851,N_19967);
nand UO_1514 (O_1514,N_19931,N_19961);
or UO_1515 (O_1515,N_19894,N_19833);
nor UO_1516 (O_1516,N_19882,N_19811);
or UO_1517 (O_1517,N_19975,N_19940);
xnor UO_1518 (O_1518,N_19901,N_19844);
or UO_1519 (O_1519,N_19942,N_19933);
and UO_1520 (O_1520,N_19948,N_19983);
and UO_1521 (O_1521,N_19862,N_19938);
xor UO_1522 (O_1522,N_19814,N_19846);
and UO_1523 (O_1523,N_19801,N_19881);
or UO_1524 (O_1524,N_19984,N_19905);
and UO_1525 (O_1525,N_19952,N_19950);
and UO_1526 (O_1526,N_19955,N_19970);
and UO_1527 (O_1527,N_19869,N_19873);
xnor UO_1528 (O_1528,N_19985,N_19995);
xnor UO_1529 (O_1529,N_19923,N_19863);
nor UO_1530 (O_1530,N_19880,N_19997);
xnor UO_1531 (O_1531,N_19816,N_19834);
xor UO_1532 (O_1532,N_19906,N_19859);
xnor UO_1533 (O_1533,N_19861,N_19967);
and UO_1534 (O_1534,N_19928,N_19958);
xnor UO_1535 (O_1535,N_19825,N_19899);
and UO_1536 (O_1536,N_19935,N_19913);
and UO_1537 (O_1537,N_19874,N_19937);
nand UO_1538 (O_1538,N_19918,N_19981);
nand UO_1539 (O_1539,N_19930,N_19862);
and UO_1540 (O_1540,N_19968,N_19888);
xnor UO_1541 (O_1541,N_19802,N_19976);
xnor UO_1542 (O_1542,N_19958,N_19815);
or UO_1543 (O_1543,N_19985,N_19987);
nor UO_1544 (O_1544,N_19933,N_19830);
xnor UO_1545 (O_1545,N_19890,N_19897);
nor UO_1546 (O_1546,N_19931,N_19903);
xor UO_1547 (O_1547,N_19808,N_19908);
and UO_1548 (O_1548,N_19977,N_19833);
or UO_1549 (O_1549,N_19828,N_19825);
xor UO_1550 (O_1550,N_19933,N_19979);
xor UO_1551 (O_1551,N_19973,N_19894);
nand UO_1552 (O_1552,N_19884,N_19904);
nor UO_1553 (O_1553,N_19815,N_19927);
nor UO_1554 (O_1554,N_19925,N_19855);
xor UO_1555 (O_1555,N_19825,N_19870);
xor UO_1556 (O_1556,N_19887,N_19996);
nor UO_1557 (O_1557,N_19876,N_19986);
xnor UO_1558 (O_1558,N_19964,N_19931);
nand UO_1559 (O_1559,N_19850,N_19975);
nand UO_1560 (O_1560,N_19814,N_19930);
xnor UO_1561 (O_1561,N_19856,N_19800);
nor UO_1562 (O_1562,N_19983,N_19999);
or UO_1563 (O_1563,N_19940,N_19850);
and UO_1564 (O_1564,N_19839,N_19902);
and UO_1565 (O_1565,N_19800,N_19850);
nand UO_1566 (O_1566,N_19991,N_19802);
xnor UO_1567 (O_1567,N_19974,N_19871);
nor UO_1568 (O_1568,N_19885,N_19833);
or UO_1569 (O_1569,N_19851,N_19921);
nand UO_1570 (O_1570,N_19977,N_19963);
or UO_1571 (O_1571,N_19973,N_19878);
or UO_1572 (O_1572,N_19997,N_19917);
nor UO_1573 (O_1573,N_19881,N_19845);
and UO_1574 (O_1574,N_19865,N_19958);
nand UO_1575 (O_1575,N_19806,N_19814);
xnor UO_1576 (O_1576,N_19873,N_19899);
xor UO_1577 (O_1577,N_19823,N_19959);
nand UO_1578 (O_1578,N_19846,N_19860);
and UO_1579 (O_1579,N_19884,N_19805);
nor UO_1580 (O_1580,N_19923,N_19832);
nor UO_1581 (O_1581,N_19929,N_19850);
xnor UO_1582 (O_1582,N_19928,N_19935);
and UO_1583 (O_1583,N_19818,N_19870);
and UO_1584 (O_1584,N_19812,N_19949);
nand UO_1585 (O_1585,N_19950,N_19867);
xor UO_1586 (O_1586,N_19933,N_19904);
and UO_1587 (O_1587,N_19930,N_19922);
xnor UO_1588 (O_1588,N_19959,N_19826);
and UO_1589 (O_1589,N_19954,N_19966);
xnor UO_1590 (O_1590,N_19983,N_19964);
nor UO_1591 (O_1591,N_19958,N_19881);
xnor UO_1592 (O_1592,N_19802,N_19884);
nor UO_1593 (O_1593,N_19834,N_19874);
xnor UO_1594 (O_1594,N_19926,N_19810);
nor UO_1595 (O_1595,N_19873,N_19918);
and UO_1596 (O_1596,N_19987,N_19815);
nor UO_1597 (O_1597,N_19857,N_19863);
and UO_1598 (O_1598,N_19803,N_19909);
xor UO_1599 (O_1599,N_19998,N_19892);
nor UO_1600 (O_1600,N_19812,N_19902);
or UO_1601 (O_1601,N_19823,N_19814);
nand UO_1602 (O_1602,N_19844,N_19851);
nor UO_1603 (O_1603,N_19960,N_19933);
nand UO_1604 (O_1604,N_19812,N_19951);
and UO_1605 (O_1605,N_19852,N_19849);
xor UO_1606 (O_1606,N_19859,N_19948);
nand UO_1607 (O_1607,N_19852,N_19854);
nand UO_1608 (O_1608,N_19804,N_19806);
nor UO_1609 (O_1609,N_19819,N_19911);
or UO_1610 (O_1610,N_19846,N_19842);
xor UO_1611 (O_1611,N_19893,N_19896);
nor UO_1612 (O_1612,N_19902,N_19868);
or UO_1613 (O_1613,N_19909,N_19889);
xnor UO_1614 (O_1614,N_19808,N_19981);
nor UO_1615 (O_1615,N_19907,N_19941);
and UO_1616 (O_1616,N_19849,N_19975);
nand UO_1617 (O_1617,N_19892,N_19987);
or UO_1618 (O_1618,N_19974,N_19908);
or UO_1619 (O_1619,N_19966,N_19907);
nor UO_1620 (O_1620,N_19942,N_19939);
nor UO_1621 (O_1621,N_19964,N_19888);
xor UO_1622 (O_1622,N_19871,N_19967);
xnor UO_1623 (O_1623,N_19910,N_19896);
nor UO_1624 (O_1624,N_19928,N_19976);
and UO_1625 (O_1625,N_19940,N_19925);
or UO_1626 (O_1626,N_19849,N_19831);
nor UO_1627 (O_1627,N_19831,N_19816);
or UO_1628 (O_1628,N_19829,N_19995);
nand UO_1629 (O_1629,N_19844,N_19878);
nor UO_1630 (O_1630,N_19892,N_19939);
xnor UO_1631 (O_1631,N_19841,N_19926);
and UO_1632 (O_1632,N_19916,N_19961);
and UO_1633 (O_1633,N_19983,N_19810);
and UO_1634 (O_1634,N_19954,N_19866);
nand UO_1635 (O_1635,N_19812,N_19957);
xnor UO_1636 (O_1636,N_19863,N_19967);
nor UO_1637 (O_1637,N_19807,N_19996);
nor UO_1638 (O_1638,N_19880,N_19931);
and UO_1639 (O_1639,N_19891,N_19894);
xnor UO_1640 (O_1640,N_19885,N_19940);
xor UO_1641 (O_1641,N_19816,N_19967);
xnor UO_1642 (O_1642,N_19901,N_19829);
and UO_1643 (O_1643,N_19996,N_19852);
nor UO_1644 (O_1644,N_19961,N_19908);
nor UO_1645 (O_1645,N_19816,N_19875);
nand UO_1646 (O_1646,N_19961,N_19950);
and UO_1647 (O_1647,N_19842,N_19896);
or UO_1648 (O_1648,N_19810,N_19924);
nand UO_1649 (O_1649,N_19805,N_19874);
or UO_1650 (O_1650,N_19932,N_19995);
nor UO_1651 (O_1651,N_19925,N_19963);
xnor UO_1652 (O_1652,N_19850,N_19954);
xor UO_1653 (O_1653,N_19983,N_19924);
nand UO_1654 (O_1654,N_19846,N_19913);
or UO_1655 (O_1655,N_19847,N_19863);
and UO_1656 (O_1656,N_19817,N_19992);
or UO_1657 (O_1657,N_19927,N_19996);
xnor UO_1658 (O_1658,N_19913,N_19857);
nor UO_1659 (O_1659,N_19897,N_19970);
and UO_1660 (O_1660,N_19843,N_19801);
nor UO_1661 (O_1661,N_19853,N_19866);
and UO_1662 (O_1662,N_19812,N_19980);
nand UO_1663 (O_1663,N_19989,N_19952);
nor UO_1664 (O_1664,N_19813,N_19893);
or UO_1665 (O_1665,N_19827,N_19987);
nand UO_1666 (O_1666,N_19835,N_19910);
xnor UO_1667 (O_1667,N_19991,N_19869);
xor UO_1668 (O_1668,N_19855,N_19888);
nor UO_1669 (O_1669,N_19899,N_19862);
nand UO_1670 (O_1670,N_19982,N_19888);
xor UO_1671 (O_1671,N_19970,N_19865);
and UO_1672 (O_1672,N_19902,N_19894);
and UO_1673 (O_1673,N_19962,N_19949);
or UO_1674 (O_1674,N_19905,N_19927);
nor UO_1675 (O_1675,N_19999,N_19817);
xor UO_1676 (O_1676,N_19893,N_19858);
nor UO_1677 (O_1677,N_19974,N_19926);
xor UO_1678 (O_1678,N_19902,N_19939);
or UO_1679 (O_1679,N_19825,N_19866);
xor UO_1680 (O_1680,N_19841,N_19820);
xnor UO_1681 (O_1681,N_19800,N_19888);
or UO_1682 (O_1682,N_19876,N_19943);
nand UO_1683 (O_1683,N_19922,N_19918);
xnor UO_1684 (O_1684,N_19866,N_19817);
and UO_1685 (O_1685,N_19885,N_19903);
nand UO_1686 (O_1686,N_19932,N_19960);
or UO_1687 (O_1687,N_19861,N_19888);
nor UO_1688 (O_1688,N_19868,N_19839);
and UO_1689 (O_1689,N_19842,N_19999);
xor UO_1690 (O_1690,N_19809,N_19848);
xor UO_1691 (O_1691,N_19872,N_19957);
xor UO_1692 (O_1692,N_19940,N_19936);
or UO_1693 (O_1693,N_19853,N_19859);
nand UO_1694 (O_1694,N_19962,N_19950);
or UO_1695 (O_1695,N_19877,N_19972);
or UO_1696 (O_1696,N_19925,N_19885);
nor UO_1697 (O_1697,N_19971,N_19809);
and UO_1698 (O_1698,N_19880,N_19846);
xor UO_1699 (O_1699,N_19822,N_19864);
or UO_1700 (O_1700,N_19872,N_19935);
nand UO_1701 (O_1701,N_19935,N_19800);
nor UO_1702 (O_1702,N_19954,N_19814);
and UO_1703 (O_1703,N_19901,N_19983);
nor UO_1704 (O_1704,N_19854,N_19917);
nor UO_1705 (O_1705,N_19975,N_19867);
nand UO_1706 (O_1706,N_19803,N_19861);
or UO_1707 (O_1707,N_19984,N_19923);
and UO_1708 (O_1708,N_19871,N_19855);
and UO_1709 (O_1709,N_19843,N_19922);
nor UO_1710 (O_1710,N_19950,N_19881);
or UO_1711 (O_1711,N_19837,N_19910);
xnor UO_1712 (O_1712,N_19986,N_19817);
nor UO_1713 (O_1713,N_19970,N_19963);
or UO_1714 (O_1714,N_19970,N_19935);
nor UO_1715 (O_1715,N_19861,N_19902);
nand UO_1716 (O_1716,N_19851,N_19832);
xnor UO_1717 (O_1717,N_19969,N_19930);
or UO_1718 (O_1718,N_19849,N_19823);
nor UO_1719 (O_1719,N_19943,N_19843);
nand UO_1720 (O_1720,N_19827,N_19838);
or UO_1721 (O_1721,N_19869,N_19975);
nand UO_1722 (O_1722,N_19865,N_19984);
and UO_1723 (O_1723,N_19827,N_19923);
or UO_1724 (O_1724,N_19829,N_19837);
nor UO_1725 (O_1725,N_19849,N_19866);
nand UO_1726 (O_1726,N_19902,N_19851);
or UO_1727 (O_1727,N_19927,N_19918);
xor UO_1728 (O_1728,N_19879,N_19962);
and UO_1729 (O_1729,N_19995,N_19809);
nor UO_1730 (O_1730,N_19862,N_19828);
nand UO_1731 (O_1731,N_19843,N_19930);
or UO_1732 (O_1732,N_19801,N_19974);
or UO_1733 (O_1733,N_19941,N_19874);
nand UO_1734 (O_1734,N_19888,N_19925);
or UO_1735 (O_1735,N_19816,N_19982);
xnor UO_1736 (O_1736,N_19873,N_19849);
and UO_1737 (O_1737,N_19879,N_19861);
xor UO_1738 (O_1738,N_19979,N_19831);
and UO_1739 (O_1739,N_19801,N_19951);
xor UO_1740 (O_1740,N_19987,N_19983);
nand UO_1741 (O_1741,N_19901,N_19917);
nand UO_1742 (O_1742,N_19860,N_19895);
and UO_1743 (O_1743,N_19819,N_19984);
xor UO_1744 (O_1744,N_19873,N_19937);
xor UO_1745 (O_1745,N_19966,N_19864);
and UO_1746 (O_1746,N_19869,N_19977);
nor UO_1747 (O_1747,N_19853,N_19809);
nand UO_1748 (O_1748,N_19900,N_19929);
xnor UO_1749 (O_1749,N_19959,N_19851);
xnor UO_1750 (O_1750,N_19888,N_19853);
nor UO_1751 (O_1751,N_19915,N_19902);
xnor UO_1752 (O_1752,N_19921,N_19875);
xor UO_1753 (O_1753,N_19932,N_19888);
xnor UO_1754 (O_1754,N_19806,N_19844);
nor UO_1755 (O_1755,N_19914,N_19842);
or UO_1756 (O_1756,N_19929,N_19852);
or UO_1757 (O_1757,N_19975,N_19986);
or UO_1758 (O_1758,N_19990,N_19920);
xor UO_1759 (O_1759,N_19875,N_19951);
or UO_1760 (O_1760,N_19927,N_19820);
or UO_1761 (O_1761,N_19905,N_19879);
or UO_1762 (O_1762,N_19801,N_19875);
or UO_1763 (O_1763,N_19893,N_19943);
nor UO_1764 (O_1764,N_19876,N_19968);
or UO_1765 (O_1765,N_19887,N_19911);
nor UO_1766 (O_1766,N_19812,N_19842);
and UO_1767 (O_1767,N_19861,N_19845);
nor UO_1768 (O_1768,N_19995,N_19986);
xor UO_1769 (O_1769,N_19914,N_19928);
xnor UO_1770 (O_1770,N_19945,N_19925);
xnor UO_1771 (O_1771,N_19839,N_19904);
nor UO_1772 (O_1772,N_19994,N_19951);
or UO_1773 (O_1773,N_19855,N_19991);
nand UO_1774 (O_1774,N_19863,N_19987);
xor UO_1775 (O_1775,N_19879,N_19969);
or UO_1776 (O_1776,N_19811,N_19971);
or UO_1777 (O_1777,N_19854,N_19835);
nor UO_1778 (O_1778,N_19831,N_19891);
nand UO_1779 (O_1779,N_19884,N_19814);
nand UO_1780 (O_1780,N_19840,N_19831);
or UO_1781 (O_1781,N_19864,N_19805);
nor UO_1782 (O_1782,N_19846,N_19907);
nor UO_1783 (O_1783,N_19817,N_19875);
and UO_1784 (O_1784,N_19868,N_19905);
or UO_1785 (O_1785,N_19870,N_19947);
and UO_1786 (O_1786,N_19910,N_19986);
or UO_1787 (O_1787,N_19978,N_19854);
xor UO_1788 (O_1788,N_19866,N_19854);
xor UO_1789 (O_1789,N_19907,N_19837);
nand UO_1790 (O_1790,N_19810,N_19822);
nand UO_1791 (O_1791,N_19941,N_19809);
nor UO_1792 (O_1792,N_19903,N_19801);
xnor UO_1793 (O_1793,N_19866,N_19873);
nor UO_1794 (O_1794,N_19822,N_19905);
nand UO_1795 (O_1795,N_19866,N_19867);
or UO_1796 (O_1796,N_19921,N_19818);
nand UO_1797 (O_1797,N_19989,N_19946);
nand UO_1798 (O_1798,N_19940,N_19953);
or UO_1799 (O_1799,N_19892,N_19841);
xnor UO_1800 (O_1800,N_19944,N_19956);
nand UO_1801 (O_1801,N_19912,N_19850);
or UO_1802 (O_1802,N_19905,N_19914);
nand UO_1803 (O_1803,N_19823,N_19873);
xnor UO_1804 (O_1804,N_19815,N_19962);
xor UO_1805 (O_1805,N_19918,N_19974);
or UO_1806 (O_1806,N_19879,N_19979);
nand UO_1807 (O_1807,N_19887,N_19802);
nor UO_1808 (O_1808,N_19942,N_19886);
or UO_1809 (O_1809,N_19989,N_19975);
xor UO_1810 (O_1810,N_19839,N_19921);
and UO_1811 (O_1811,N_19912,N_19909);
nor UO_1812 (O_1812,N_19857,N_19935);
xnor UO_1813 (O_1813,N_19993,N_19948);
or UO_1814 (O_1814,N_19953,N_19868);
or UO_1815 (O_1815,N_19800,N_19857);
or UO_1816 (O_1816,N_19829,N_19833);
nand UO_1817 (O_1817,N_19850,N_19968);
and UO_1818 (O_1818,N_19942,N_19877);
xor UO_1819 (O_1819,N_19944,N_19820);
or UO_1820 (O_1820,N_19944,N_19888);
xnor UO_1821 (O_1821,N_19862,N_19965);
nor UO_1822 (O_1822,N_19896,N_19802);
or UO_1823 (O_1823,N_19868,N_19895);
and UO_1824 (O_1824,N_19984,N_19840);
or UO_1825 (O_1825,N_19922,N_19882);
nor UO_1826 (O_1826,N_19987,N_19968);
nand UO_1827 (O_1827,N_19862,N_19924);
xnor UO_1828 (O_1828,N_19972,N_19817);
nor UO_1829 (O_1829,N_19976,N_19853);
nor UO_1830 (O_1830,N_19949,N_19987);
and UO_1831 (O_1831,N_19870,N_19966);
xnor UO_1832 (O_1832,N_19937,N_19912);
xor UO_1833 (O_1833,N_19944,N_19906);
and UO_1834 (O_1834,N_19845,N_19936);
and UO_1835 (O_1835,N_19998,N_19808);
nand UO_1836 (O_1836,N_19813,N_19886);
and UO_1837 (O_1837,N_19981,N_19812);
nor UO_1838 (O_1838,N_19903,N_19946);
or UO_1839 (O_1839,N_19928,N_19893);
xor UO_1840 (O_1840,N_19825,N_19925);
nand UO_1841 (O_1841,N_19846,N_19921);
or UO_1842 (O_1842,N_19869,N_19814);
nand UO_1843 (O_1843,N_19969,N_19962);
or UO_1844 (O_1844,N_19964,N_19953);
nor UO_1845 (O_1845,N_19868,N_19821);
nor UO_1846 (O_1846,N_19896,N_19895);
nand UO_1847 (O_1847,N_19984,N_19972);
xor UO_1848 (O_1848,N_19881,N_19930);
xor UO_1849 (O_1849,N_19989,N_19929);
and UO_1850 (O_1850,N_19997,N_19834);
nand UO_1851 (O_1851,N_19825,N_19977);
nand UO_1852 (O_1852,N_19913,N_19805);
xnor UO_1853 (O_1853,N_19864,N_19963);
or UO_1854 (O_1854,N_19872,N_19816);
and UO_1855 (O_1855,N_19839,N_19879);
nand UO_1856 (O_1856,N_19983,N_19825);
nor UO_1857 (O_1857,N_19950,N_19918);
xnor UO_1858 (O_1858,N_19931,N_19816);
and UO_1859 (O_1859,N_19954,N_19925);
or UO_1860 (O_1860,N_19926,N_19913);
or UO_1861 (O_1861,N_19890,N_19977);
nor UO_1862 (O_1862,N_19954,N_19993);
nand UO_1863 (O_1863,N_19932,N_19869);
and UO_1864 (O_1864,N_19861,N_19974);
nor UO_1865 (O_1865,N_19864,N_19960);
xnor UO_1866 (O_1866,N_19908,N_19989);
or UO_1867 (O_1867,N_19824,N_19928);
and UO_1868 (O_1868,N_19996,N_19890);
or UO_1869 (O_1869,N_19912,N_19984);
nor UO_1870 (O_1870,N_19923,N_19902);
and UO_1871 (O_1871,N_19956,N_19914);
nor UO_1872 (O_1872,N_19909,N_19863);
or UO_1873 (O_1873,N_19955,N_19976);
nand UO_1874 (O_1874,N_19945,N_19879);
and UO_1875 (O_1875,N_19981,N_19901);
xnor UO_1876 (O_1876,N_19823,N_19893);
and UO_1877 (O_1877,N_19817,N_19883);
xor UO_1878 (O_1878,N_19949,N_19821);
nand UO_1879 (O_1879,N_19963,N_19852);
nor UO_1880 (O_1880,N_19802,N_19831);
and UO_1881 (O_1881,N_19913,N_19810);
nor UO_1882 (O_1882,N_19935,N_19912);
and UO_1883 (O_1883,N_19992,N_19976);
nand UO_1884 (O_1884,N_19834,N_19955);
nand UO_1885 (O_1885,N_19843,N_19984);
nand UO_1886 (O_1886,N_19984,N_19941);
and UO_1887 (O_1887,N_19993,N_19836);
or UO_1888 (O_1888,N_19818,N_19926);
xor UO_1889 (O_1889,N_19815,N_19861);
and UO_1890 (O_1890,N_19824,N_19806);
nor UO_1891 (O_1891,N_19806,N_19909);
nor UO_1892 (O_1892,N_19837,N_19825);
nor UO_1893 (O_1893,N_19941,N_19997);
or UO_1894 (O_1894,N_19859,N_19941);
nor UO_1895 (O_1895,N_19820,N_19919);
nor UO_1896 (O_1896,N_19836,N_19911);
or UO_1897 (O_1897,N_19820,N_19902);
nor UO_1898 (O_1898,N_19835,N_19875);
and UO_1899 (O_1899,N_19829,N_19888);
and UO_1900 (O_1900,N_19992,N_19938);
or UO_1901 (O_1901,N_19945,N_19898);
xnor UO_1902 (O_1902,N_19926,N_19868);
nand UO_1903 (O_1903,N_19990,N_19830);
nor UO_1904 (O_1904,N_19860,N_19965);
nand UO_1905 (O_1905,N_19987,N_19960);
nor UO_1906 (O_1906,N_19803,N_19873);
nand UO_1907 (O_1907,N_19940,N_19971);
nor UO_1908 (O_1908,N_19895,N_19823);
or UO_1909 (O_1909,N_19835,N_19930);
and UO_1910 (O_1910,N_19868,N_19890);
nor UO_1911 (O_1911,N_19933,N_19819);
and UO_1912 (O_1912,N_19903,N_19856);
or UO_1913 (O_1913,N_19928,N_19966);
xnor UO_1914 (O_1914,N_19836,N_19926);
nand UO_1915 (O_1915,N_19834,N_19892);
nor UO_1916 (O_1916,N_19803,N_19934);
nor UO_1917 (O_1917,N_19828,N_19921);
nor UO_1918 (O_1918,N_19861,N_19959);
nor UO_1919 (O_1919,N_19800,N_19822);
nor UO_1920 (O_1920,N_19958,N_19863);
nand UO_1921 (O_1921,N_19937,N_19860);
nand UO_1922 (O_1922,N_19923,N_19934);
and UO_1923 (O_1923,N_19815,N_19980);
nor UO_1924 (O_1924,N_19885,N_19984);
and UO_1925 (O_1925,N_19814,N_19946);
xnor UO_1926 (O_1926,N_19909,N_19931);
or UO_1927 (O_1927,N_19800,N_19943);
and UO_1928 (O_1928,N_19934,N_19859);
nand UO_1929 (O_1929,N_19939,N_19807);
nor UO_1930 (O_1930,N_19863,N_19982);
xnor UO_1931 (O_1931,N_19864,N_19954);
nor UO_1932 (O_1932,N_19958,N_19839);
nand UO_1933 (O_1933,N_19839,N_19823);
xor UO_1934 (O_1934,N_19910,N_19888);
and UO_1935 (O_1935,N_19836,N_19890);
and UO_1936 (O_1936,N_19927,N_19995);
or UO_1937 (O_1937,N_19931,N_19862);
nand UO_1938 (O_1938,N_19801,N_19998);
nand UO_1939 (O_1939,N_19835,N_19973);
and UO_1940 (O_1940,N_19910,N_19931);
xor UO_1941 (O_1941,N_19978,N_19998);
nand UO_1942 (O_1942,N_19994,N_19996);
nand UO_1943 (O_1943,N_19840,N_19804);
and UO_1944 (O_1944,N_19887,N_19880);
nand UO_1945 (O_1945,N_19943,N_19880);
nand UO_1946 (O_1946,N_19901,N_19834);
xnor UO_1947 (O_1947,N_19890,N_19854);
nand UO_1948 (O_1948,N_19850,N_19845);
nor UO_1949 (O_1949,N_19807,N_19913);
xnor UO_1950 (O_1950,N_19824,N_19835);
xor UO_1951 (O_1951,N_19907,N_19977);
or UO_1952 (O_1952,N_19908,N_19946);
or UO_1953 (O_1953,N_19963,N_19879);
nor UO_1954 (O_1954,N_19930,N_19910);
nand UO_1955 (O_1955,N_19895,N_19978);
nor UO_1956 (O_1956,N_19968,N_19852);
and UO_1957 (O_1957,N_19866,N_19881);
nor UO_1958 (O_1958,N_19935,N_19942);
nand UO_1959 (O_1959,N_19826,N_19951);
xor UO_1960 (O_1960,N_19844,N_19859);
nand UO_1961 (O_1961,N_19802,N_19827);
xnor UO_1962 (O_1962,N_19954,N_19878);
and UO_1963 (O_1963,N_19865,N_19917);
nand UO_1964 (O_1964,N_19851,N_19989);
and UO_1965 (O_1965,N_19861,N_19997);
nor UO_1966 (O_1966,N_19923,N_19899);
nand UO_1967 (O_1967,N_19955,N_19911);
or UO_1968 (O_1968,N_19914,N_19829);
xnor UO_1969 (O_1969,N_19800,N_19898);
or UO_1970 (O_1970,N_19984,N_19953);
and UO_1971 (O_1971,N_19808,N_19944);
and UO_1972 (O_1972,N_19903,N_19919);
and UO_1973 (O_1973,N_19926,N_19846);
or UO_1974 (O_1974,N_19926,N_19928);
and UO_1975 (O_1975,N_19943,N_19988);
and UO_1976 (O_1976,N_19962,N_19957);
nor UO_1977 (O_1977,N_19911,N_19848);
nor UO_1978 (O_1978,N_19893,N_19957);
nor UO_1979 (O_1979,N_19861,N_19884);
nand UO_1980 (O_1980,N_19932,N_19846);
or UO_1981 (O_1981,N_19843,N_19933);
xor UO_1982 (O_1982,N_19822,N_19844);
or UO_1983 (O_1983,N_19970,N_19811);
nand UO_1984 (O_1984,N_19912,N_19855);
or UO_1985 (O_1985,N_19841,N_19890);
or UO_1986 (O_1986,N_19834,N_19931);
xnor UO_1987 (O_1987,N_19911,N_19842);
nor UO_1988 (O_1988,N_19890,N_19803);
xnor UO_1989 (O_1989,N_19987,N_19861);
or UO_1990 (O_1990,N_19870,N_19879);
and UO_1991 (O_1991,N_19882,N_19944);
nand UO_1992 (O_1992,N_19969,N_19902);
xnor UO_1993 (O_1993,N_19953,N_19949);
or UO_1994 (O_1994,N_19843,N_19958);
and UO_1995 (O_1995,N_19867,N_19960);
or UO_1996 (O_1996,N_19835,N_19816);
or UO_1997 (O_1997,N_19987,N_19957);
nand UO_1998 (O_1998,N_19811,N_19938);
nor UO_1999 (O_1999,N_19906,N_19938);
xnor UO_2000 (O_2000,N_19998,N_19804);
nand UO_2001 (O_2001,N_19814,N_19926);
nand UO_2002 (O_2002,N_19835,N_19982);
nand UO_2003 (O_2003,N_19901,N_19944);
nor UO_2004 (O_2004,N_19966,N_19801);
xnor UO_2005 (O_2005,N_19953,N_19956);
or UO_2006 (O_2006,N_19899,N_19988);
nand UO_2007 (O_2007,N_19850,N_19823);
nand UO_2008 (O_2008,N_19803,N_19914);
xor UO_2009 (O_2009,N_19875,N_19848);
xor UO_2010 (O_2010,N_19871,N_19981);
nand UO_2011 (O_2011,N_19990,N_19815);
xnor UO_2012 (O_2012,N_19816,N_19955);
nand UO_2013 (O_2013,N_19865,N_19921);
and UO_2014 (O_2014,N_19904,N_19860);
xor UO_2015 (O_2015,N_19905,N_19873);
or UO_2016 (O_2016,N_19813,N_19946);
or UO_2017 (O_2017,N_19966,N_19968);
and UO_2018 (O_2018,N_19867,N_19996);
or UO_2019 (O_2019,N_19968,N_19973);
nand UO_2020 (O_2020,N_19888,N_19906);
nand UO_2021 (O_2021,N_19956,N_19903);
xnor UO_2022 (O_2022,N_19944,N_19919);
or UO_2023 (O_2023,N_19853,N_19894);
or UO_2024 (O_2024,N_19872,N_19940);
and UO_2025 (O_2025,N_19857,N_19886);
and UO_2026 (O_2026,N_19823,N_19826);
and UO_2027 (O_2027,N_19882,N_19904);
xor UO_2028 (O_2028,N_19806,N_19925);
and UO_2029 (O_2029,N_19925,N_19841);
xnor UO_2030 (O_2030,N_19806,N_19854);
and UO_2031 (O_2031,N_19832,N_19997);
xnor UO_2032 (O_2032,N_19811,N_19855);
xor UO_2033 (O_2033,N_19942,N_19965);
nor UO_2034 (O_2034,N_19891,N_19879);
and UO_2035 (O_2035,N_19887,N_19928);
nand UO_2036 (O_2036,N_19824,N_19896);
nor UO_2037 (O_2037,N_19954,N_19869);
nor UO_2038 (O_2038,N_19965,N_19878);
nand UO_2039 (O_2039,N_19868,N_19802);
or UO_2040 (O_2040,N_19872,N_19848);
nand UO_2041 (O_2041,N_19974,N_19930);
nor UO_2042 (O_2042,N_19823,N_19876);
and UO_2043 (O_2043,N_19872,N_19902);
xnor UO_2044 (O_2044,N_19964,N_19982);
nand UO_2045 (O_2045,N_19898,N_19921);
and UO_2046 (O_2046,N_19830,N_19906);
and UO_2047 (O_2047,N_19819,N_19931);
nand UO_2048 (O_2048,N_19996,N_19865);
nor UO_2049 (O_2049,N_19870,N_19839);
or UO_2050 (O_2050,N_19944,N_19894);
and UO_2051 (O_2051,N_19804,N_19943);
nand UO_2052 (O_2052,N_19999,N_19866);
xnor UO_2053 (O_2053,N_19981,N_19884);
xor UO_2054 (O_2054,N_19859,N_19907);
and UO_2055 (O_2055,N_19916,N_19905);
nand UO_2056 (O_2056,N_19834,N_19865);
xor UO_2057 (O_2057,N_19874,N_19872);
xor UO_2058 (O_2058,N_19923,N_19846);
nand UO_2059 (O_2059,N_19878,N_19969);
or UO_2060 (O_2060,N_19918,N_19954);
or UO_2061 (O_2061,N_19846,N_19823);
xnor UO_2062 (O_2062,N_19850,N_19937);
xnor UO_2063 (O_2063,N_19828,N_19915);
nand UO_2064 (O_2064,N_19923,N_19912);
and UO_2065 (O_2065,N_19896,N_19920);
nor UO_2066 (O_2066,N_19858,N_19934);
xnor UO_2067 (O_2067,N_19938,N_19872);
and UO_2068 (O_2068,N_19966,N_19825);
and UO_2069 (O_2069,N_19926,N_19946);
nor UO_2070 (O_2070,N_19817,N_19965);
xnor UO_2071 (O_2071,N_19944,N_19851);
nor UO_2072 (O_2072,N_19832,N_19893);
or UO_2073 (O_2073,N_19852,N_19833);
xor UO_2074 (O_2074,N_19879,N_19954);
or UO_2075 (O_2075,N_19809,N_19992);
or UO_2076 (O_2076,N_19825,N_19935);
and UO_2077 (O_2077,N_19953,N_19970);
and UO_2078 (O_2078,N_19895,N_19857);
nor UO_2079 (O_2079,N_19801,N_19862);
or UO_2080 (O_2080,N_19975,N_19956);
nand UO_2081 (O_2081,N_19983,N_19994);
nor UO_2082 (O_2082,N_19942,N_19819);
or UO_2083 (O_2083,N_19863,N_19949);
or UO_2084 (O_2084,N_19876,N_19854);
nor UO_2085 (O_2085,N_19816,N_19966);
nor UO_2086 (O_2086,N_19986,N_19926);
xor UO_2087 (O_2087,N_19892,N_19940);
nor UO_2088 (O_2088,N_19970,N_19872);
nand UO_2089 (O_2089,N_19992,N_19933);
and UO_2090 (O_2090,N_19942,N_19968);
xor UO_2091 (O_2091,N_19801,N_19988);
and UO_2092 (O_2092,N_19981,N_19809);
nor UO_2093 (O_2093,N_19922,N_19881);
xor UO_2094 (O_2094,N_19904,N_19991);
and UO_2095 (O_2095,N_19869,N_19972);
or UO_2096 (O_2096,N_19990,N_19817);
and UO_2097 (O_2097,N_19823,N_19857);
nor UO_2098 (O_2098,N_19877,N_19897);
xor UO_2099 (O_2099,N_19846,N_19894);
nand UO_2100 (O_2100,N_19965,N_19819);
or UO_2101 (O_2101,N_19921,N_19860);
and UO_2102 (O_2102,N_19933,N_19832);
and UO_2103 (O_2103,N_19897,N_19801);
nor UO_2104 (O_2104,N_19804,N_19911);
nor UO_2105 (O_2105,N_19932,N_19822);
and UO_2106 (O_2106,N_19915,N_19936);
and UO_2107 (O_2107,N_19962,N_19974);
xnor UO_2108 (O_2108,N_19850,N_19974);
and UO_2109 (O_2109,N_19885,N_19847);
xor UO_2110 (O_2110,N_19954,N_19943);
nor UO_2111 (O_2111,N_19870,N_19836);
nor UO_2112 (O_2112,N_19934,N_19807);
xor UO_2113 (O_2113,N_19903,N_19969);
xor UO_2114 (O_2114,N_19898,N_19825);
nand UO_2115 (O_2115,N_19969,N_19901);
or UO_2116 (O_2116,N_19801,N_19921);
nand UO_2117 (O_2117,N_19933,N_19856);
nand UO_2118 (O_2118,N_19974,N_19997);
xnor UO_2119 (O_2119,N_19879,N_19854);
xor UO_2120 (O_2120,N_19812,N_19930);
nand UO_2121 (O_2121,N_19940,N_19905);
nor UO_2122 (O_2122,N_19912,N_19864);
xor UO_2123 (O_2123,N_19998,N_19964);
xnor UO_2124 (O_2124,N_19861,N_19834);
nand UO_2125 (O_2125,N_19999,N_19989);
or UO_2126 (O_2126,N_19817,N_19804);
xor UO_2127 (O_2127,N_19962,N_19850);
or UO_2128 (O_2128,N_19966,N_19990);
nor UO_2129 (O_2129,N_19875,N_19931);
nor UO_2130 (O_2130,N_19962,N_19963);
nor UO_2131 (O_2131,N_19813,N_19823);
nor UO_2132 (O_2132,N_19836,N_19830);
xnor UO_2133 (O_2133,N_19906,N_19809);
nor UO_2134 (O_2134,N_19945,N_19952);
or UO_2135 (O_2135,N_19808,N_19871);
nor UO_2136 (O_2136,N_19934,N_19954);
xnor UO_2137 (O_2137,N_19973,N_19904);
nand UO_2138 (O_2138,N_19991,N_19981);
and UO_2139 (O_2139,N_19973,N_19992);
and UO_2140 (O_2140,N_19846,N_19807);
or UO_2141 (O_2141,N_19969,N_19867);
nand UO_2142 (O_2142,N_19963,N_19847);
or UO_2143 (O_2143,N_19878,N_19935);
or UO_2144 (O_2144,N_19887,N_19896);
and UO_2145 (O_2145,N_19990,N_19923);
nand UO_2146 (O_2146,N_19848,N_19950);
or UO_2147 (O_2147,N_19842,N_19917);
nand UO_2148 (O_2148,N_19884,N_19975);
xnor UO_2149 (O_2149,N_19902,N_19829);
xnor UO_2150 (O_2150,N_19962,N_19972);
and UO_2151 (O_2151,N_19973,N_19870);
and UO_2152 (O_2152,N_19887,N_19852);
xnor UO_2153 (O_2153,N_19827,N_19997);
or UO_2154 (O_2154,N_19880,N_19863);
nand UO_2155 (O_2155,N_19831,N_19846);
and UO_2156 (O_2156,N_19860,N_19812);
xnor UO_2157 (O_2157,N_19979,N_19823);
and UO_2158 (O_2158,N_19903,N_19813);
nor UO_2159 (O_2159,N_19851,N_19886);
nor UO_2160 (O_2160,N_19885,N_19889);
and UO_2161 (O_2161,N_19895,N_19824);
or UO_2162 (O_2162,N_19866,N_19920);
or UO_2163 (O_2163,N_19874,N_19800);
nand UO_2164 (O_2164,N_19993,N_19851);
xor UO_2165 (O_2165,N_19973,N_19868);
nand UO_2166 (O_2166,N_19896,N_19892);
or UO_2167 (O_2167,N_19806,N_19987);
xor UO_2168 (O_2168,N_19823,N_19925);
nor UO_2169 (O_2169,N_19981,N_19865);
nand UO_2170 (O_2170,N_19856,N_19836);
xnor UO_2171 (O_2171,N_19981,N_19902);
nand UO_2172 (O_2172,N_19833,N_19811);
or UO_2173 (O_2173,N_19829,N_19896);
and UO_2174 (O_2174,N_19872,N_19832);
nand UO_2175 (O_2175,N_19859,N_19885);
or UO_2176 (O_2176,N_19848,N_19916);
nor UO_2177 (O_2177,N_19851,N_19999);
or UO_2178 (O_2178,N_19846,N_19891);
xnor UO_2179 (O_2179,N_19958,N_19893);
or UO_2180 (O_2180,N_19885,N_19862);
or UO_2181 (O_2181,N_19975,N_19966);
nand UO_2182 (O_2182,N_19982,N_19894);
nand UO_2183 (O_2183,N_19825,N_19963);
and UO_2184 (O_2184,N_19940,N_19800);
and UO_2185 (O_2185,N_19999,N_19913);
or UO_2186 (O_2186,N_19805,N_19981);
xor UO_2187 (O_2187,N_19968,N_19832);
or UO_2188 (O_2188,N_19805,N_19869);
nor UO_2189 (O_2189,N_19898,N_19933);
nand UO_2190 (O_2190,N_19894,N_19959);
nand UO_2191 (O_2191,N_19870,N_19930);
nor UO_2192 (O_2192,N_19965,N_19972);
or UO_2193 (O_2193,N_19960,N_19863);
and UO_2194 (O_2194,N_19944,N_19998);
and UO_2195 (O_2195,N_19975,N_19987);
or UO_2196 (O_2196,N_19825,N_19809);
xor UO_2197 (O_2197,N_19917,N_19818);
nand UO_2198 (O_2198,N_19892,N_19825);
nand UO_2199 (O_2199,N_19941,N_19810);
and UO_2200 (O_2200,N_19853,N_19988);
nand UO_2201 (O_2201,N_19854,N_19954);
nor UO_2202 (O_2202,N_19965,N_19928);
or UO_2203 (O_2203,N_19827,N_19857);
nand UO_2204 (O_2204,N_19920,N_19835);
xnor UO_2205 (O_2205,N_19994,N_19891);
nand UO_2206 (O_2206,N_19807,N_19918);
nand UO_2207 (O_2207,N_19807,N_19991);
and UO_2208 (O_2208,N_19904,N_19866);
and UO_2209 (O_2209,N_19940,N_19960);
xor UO_2210 (O_2210,N_19952,N_19882);
or UO_2211 (O_2211,N_19921,N_19949);
and UO_2212 (O_2212,N_19919,N_19965);
nand UO_2213 (O_2213,N_19953,N_19811);
xor UO_2214 (O_2214,N_19966,N_19804);
nor UO_2215 (O_2215,N_19819,N_19860);
or UO_2216 (O_2216,N_19826,N_19907);
nor UO_2217 (O_2217,N_19916,N_19921);
xnor UO_2218 (O_2218,N_19889,N_19837);
nand UO_2219 (O_2219,N_19865,N_19820);
nand UO_2220 (O_2220,N_19853,N_19903);
xnor UO_2221 (O_2221,N_19971,N_19977);
nand UO_2222 (O_2222,N_19916,N_19867);
and UO_2223 (O_2223,N_19801,N_19928);
xor UO_2224 (O_2224,N_19958,N_19808);
nand UO_2225 (O_2225,N_19917,N_19974);
and UO_2226 (O_2226,N_19973,N_19994);
xor UO_2227 (O_2227,N_19826,N_19935);
or UO_2228 (O_2228,N_19865,N_19869);
or UO_2229 (O_2229,N_19994,N_19807);
nand UO_2230 (O_2230,N_19867,N_19860);
and UO_2231 (O_2231,N_19849,N_19909);
or UO_2232 (O_2232,N_19965,N_19885);
xnor UO_2233 (O_2233,N_19896,N_19871);
xor UO_2234 (O_2234,N_19969,N_19953);
xor UO_2235 (O_2235,N_19806,N_19865);
and UO_2236 (O_2236,N_19894,N_19989);
nor UO_2237 (O_2237,N_19953,N_19859);
xnor UO_2238 (O_2238,N_19812,N_19895);
nand UO_2239 (O_2239,N_19974,N_19985);
nand UO_2240 (O_2240,N_19915,N_19868);
and UO_2241 (O_2241,N_19888,N_19966);
nor UO_2242 (O_2242,N_19802,N_19893);
or UO_2243 (O_2243,N_19919,N_19800);
nor UO_2244 (O_2244,N_19850,N_19842);
xnor UO_2245 (O_2245,N_19869,N_19832);
nor UO_2246 (O_2246,N_19923,N_19920);
xnor UO_2247 (O_2247,N_19892,N_19900);
nand UO_2248 (O_2248,N_19803,N_19989);
nand UO_2249 (O_2249,N_19981,N_19947);
nor UO_2250 (O_2250,N_19875,N_19884);
or UO_2251 (O_2251,N_19938,N_19849);
nand UO_2252 (O_2252,N_19817,N_19800);
or UO_2253 (O_2253,N_19833,N_19888);
nand UO_2254 (O_2254,N_19866,N_19979);
or UO_2255 (O_2255,N_19883,N_19921);
nand UO_2256 (O_2256,N_19987,N_19982);
or UO_2257 (O_2257,N_19900,N_19871);
nor UO_2258 (O_2258,N_19950,N_19936);
xor UO_2259 (O_2259,N_19934,N_19839);
xor UO_2260 (O_2260,N_19969,N_19974);
xnor UO_2261 (O_2261,N_19939,N_19990);
nor UO_2262 (O_2262,N_19811,N_19867);
nand UO_2263 (O_2263,N_19862,N_19944);
nand UO_2264 (O_2264,N_19917,N_19996);
nand UO_2265 (O_2265,N_19936,N_19934);
xor UO_2266 (O_2266,N_19978,N_19924);
and UO_2267 (O_2267,N_19889,N_19842);
or UO_2268 (O_2268,N_19810,N_19988);
and UO_2269 (O_2269,N_19885,N_19933);
nand UO_2270 (O_2270,N_19895,N_19839);
or UO_2271 (O_2271,N_19868,N_19873);
nor UO_2272 (O_2272,N_19989,N_19805);
nor UO_2273 (O_2273,N_19814,N_19830);
or UO_2274 (O_2274,N_19834,N_19921);
xor UO_2275 (O_2275,N_19934,N_19950);
nor UO_2276 (O_2276,N_19878,N_19825);
or UO_2277 (O_2277,N_19870,N_19840);
or UO_2278 (O_2278,N_19862,N_19998);
and UO_2279 (O_2279,N_19826,N_19983);
or UO_2280 (O_2280,N_19811,N_19902);
xor UO_2281 (O_2281,N_19991,N_19875);
nand UO_2282 (O_2282,N_19860,N_19828);
and UO_2283 (O_2283,N_19867,N_19859);
nand UO_2284 (O_2284,N_19982,N_19839);
nand UO_2285 (O_2285,N_19974,N_19832);
nand UO_2286 (O_2286,N_19825,N_19851);
nand UO_2287 (O_2287,N_19864,N_19996);
and UO_2288 (O_2288,N_19887,N_19836);
and UO_2289 (O_2289,N_19891,N_19969);
or UO_2290 (O_2290,N_19815,N_19920);
nand UO_2291 (O_2291,N_19862,N_19803);
nor UO_2292 (O_2292,N_19841,N_19909);
nor UO_2293 (O_2293,N_19947,N_19822);
or UO_2294 (O_2294,N_19848,N_19852);
nor UO_2295 (O_2295,N_19893,N_19850);
nor UO_2296 (O_2296,N_19835,N_19890);
nor UO_2297 (O_2297,N_19979,N_19846);
xnor UO_2298 (O_2298,N_19958,N_19853);
nor UO_2299 (O_2299,N_19867,N_19878);
or UO_2300 (O_2300,N_19810,N_19910);
or UO_2301 (O_2301,N_19926,N_19995);
nand UO_2302 (O_2302,N_19927,N_19816);
nand UO_2303 (O_2303,N_19991,N_19969);
nand UO_2304 (O_2304,N_19999,N_19927);
xor UO_2305 (O_2305,N_19858,N_19828);
nand UO_2306 (O_2306,N_19991,N_19957);
and UO_2307 (O_2307,N_19965,N_19881);
nand UO_2308 (O_2308,N_19966,N_19994);
or UO_2309 (O_2309,N_19922,N_19813);
nor UO_2310 (O_2310,N_19942,N_19888);
nand UO_2311 (O_2311,N_19936,N_19835);
xnor UO_2312 (O_2312,N_19903,N_19921);
and UO_2313 (O_2313,N_19989,N_19925);
nor UO_2314 (O_2314,N_19898,N_19850);
nor UO_2315 (O_2315,N_19820,N_19975);
or UO_2316 (O_2316,N_19801,N_19846);
nor UO_2317 (O_2317,N_19802,N_19978);
nand UO_2318 (O_2318,N_19927,N_19873);
nand UO_2319 (O_2319,N_19963,N_19846);
and UO_2320 (O_2320,N_19974,N_19983);
or UO_2321 (O_2321,N_19972,N_19988);
nand UO_2322 (O_2322,N_19936,N_19997);
nor UO_2323 (O_2323,N_19810,N_19874);
nand UO_2324 (O_2324,N_19940,N_19812);
or UO_2325 (O_2325,N_19834,N_19887);
and UO_2326 (O_2326,N_19999,N_19966);
nand UO_2327 (O_2327,N_19830,N_19851);
or UO_2328 (O_2328,N_19952,N_19974);
or UO_2329 (O_2329,N_19999,N_19883);
or UO_2330 (O_2330,N_19948,N_19967);
nand UO_2331 (O_2331,N_19969,N_19997);
or UO_2332 (O_2332,N_19877,N_19875);
and UO_2333 (O_2333,N_19866,N_19879);
or UO_2334 (O_2334,N_19993,N_19850);
and UO_2335 (O_2335,N_19953,N_19934);
or UO_2336 (O_2336,N_19877,N_19920);
xnor UO_2337 (O_2337,N_19937,N_19949);
or UO_2338 (O_2338,N_19995,N_19919);
nor UO_2339 (O_2339,N_19892,N_19960);
xor UO_2340 (O_2340,N_19862,N_19852);
or UO_2341 (O_2341,N_19855,N_19847);
nand UO_2342 (O_2342,N_19848,N_19957);
and UO_2343 (O_2343,N_19933,N_19841);
nor UO_2344 (O_2344,N_19995,N_19974);
nor UO_2345 (O_2345,N_19834,N_19801);
nand UO_2346 (O_2346,N_19880,N_19930);
or UO_2347 (O_2347,N_19940,N_19805);
xnor UO_2348 (O_2348,N_19838,N_19819);
and UO_2349 (O_2349,N_19899,N_19925);
nand UO_2350 (O_2350,N_19879,N_19928);
and UO_2351 (O_2351,N_19938,N_19954);
nand UO_2352 (O_2352,N_19919,N_19907);
nand UO_2353 (O_2353,N_19914,N_19891);
and UO_2354 (O_2354,N_19901,N_19886);
nand UO_2355 (O_2355,N_19926,N_19966);
or UO_2356 (O_2356,N_19840,N_19871);
or UO_2357 (O_2357,N_19878,N_19866);
nor UO_2358 (O_2358,N_19949,N_19986);
nand UO_2359 (O_2359,N_19866,N_19974);
and UO_2360 (O_2360,N_19814,N_19821);
xor UO_2361 (O_2361,N_19850,N_19918);
or UO_2362 (O_2362,N_19963,N_19901);
and UO_2363 (O_2363,N_19999,N_19909);
and UO_2364 (O_2364,N_19877,N_19941);
or UO_2365 (O_2365,N_19981,N_19978);
nand UO_2366 (O_2366,N_19960,N_19814);
or UO_2367 (O_2367,N_19973,N_19832);
and UO_2368 (O_2368,N_19986,N_19892);
xnor UO_2369 (O_2369,N_19866,N_19949);
and UO_2370 (O_2370,N_19803,N_19804);
and UO_2371 (O_2371,N_19883,N_19878);
or UO_2372 (O_2372,N_19839,N_19894);
xor UO_2373 (O_2373,N_19984,N_19899);
and UO_2374 (O_2374,N_19898,N_19839);
xnor UO_2375 (O_2375,N_19825,N_19800);
nor UO_2376 (O_2376,N_19810,N_19851);
nor UO_2377 (O_2377,N_19870,N_19971);
nand UO_2378 (O_2378,N_19993,N_19941);
or UO_2379 (O_2379,N_19935,N_19887);
nand UO_2380 (O_2380,N_19803,N_19896);
nand UO_2381 (O_2381,N_19832,N_19874);
and UO_2382 (O_2382,N_19838,N_19901);
nor UO_2383 (O_2383,N_19806,N_19850);
nor UO_2384 (O_2384,N_19871,N_19937);
and UO_2385 (O_2385,N_19804,N_19996);
or UO_2386 (O_2386,N_19920,N_19811);
and UO_2387 (O_2387,N_19967,N_19947);
or UO_2388 (O_2388,N_19901,N_19868);
or UO_2389 (O_2389,N_19821,N_19846);
and UO_2390 (O_2390,N_19813,N_19936);
nand UO_2391 (O_2391,N_19909,N_19990);
xor UO_2392 (O_2392,N_19804,N_19859);
and UO_2393 (O_2393,N_19998,N_19856);
and UO_2394 (O_2394,N_19837,N_19821);
or UO_2395 (O_2395,N_19868,N_19887);
nor UO_2396 (O_2396,N_19877,N_19921);
nor UO_2397 (O_2397,N_19910,N_19966);
xor UO_2398 (O_2398,N_19970,N_19813);
nor UO_2399 (O_2399,N_19987,N_19930);
or UO_2400 (O_2400,N_19916,N_19879);
nor UO_2401 (O_2401,N_19937,N_19928);
and UO_2402 (O_2402,N_19870,N_19987);
or UO_2403 (O_2403,N_19932,N_19800);
nor UO_2404 (O_2404,N_19800,N_19865);
nor UO_2405 (O_2405,N_19879,N_19955);
nand UO_2406 (O_2406,N_19998,N_19900);
or UO_2407 (O_2407,N_19856,N_19879);
and UO_2408 (O_2408,N_19893,N_19863);
xor UO_2409 (O_2409,N_19915,N_19916);
nand UO_2410 (O_2410,N_19896,N_19911);
or UO_2411 (O_2411,N_19856,N_19852);
nand UO_2412 (O_2412,N_19903,N_19898);
nor UO_2413 (O_2413,N_19944,N_19989);
or UO_2414 (O_2414,N_19984,N_19821);
nand UO_2415 (O_2415,N_19802,N_19971);
xnor UO_2416 (O_2416,N_19805,N_19950);
and UO_2417 (O_2417,N_19858,N_19857);
nand UO_2418 (O_2418,N_19810,N_19993);
nand UO_2419 (O_2419,N_19906,N_19868);
or UO_2420 (O_2420,N_19828,N_19982);
xnor UO_2421 (O_2421,N_19986,N_19890);
xnor UO_2422 (O_2422,N_19920,N_19979);
or UO_2423 (O_2423,N_19901,N_19920);
or UO_2424 (O_2424,N_19957,N_19922);
nand UO_2425 (O_2425,N_19836,N_19882);
and UO_2426 (O_2426,N_19843,N_19850);
nand UO_2427 (O_2427,N_19858,N_19933);
and UO_2428 (O_2428,N_19853,N_19957);
nand UO_2429 (O_2429,N_19974,N_19810);
xnor UO_2430 (O_2430,N_19956,N_19840);
nor UO_2431 (O_2431,N_19928,N_19910);
nand UO_2432 (O_2432,N_19957,N_19980);
nor UO_2433 (O_2433,N_19867,N_19982);
xnor UO_2434 (O_2434,N_19921,N_19939);
xnor UO_2435 (O_2435,N_19945,N_19890);
nand UO_2436 (O_2436,N_19803,N_19839);
xor UO_2437 (O_2437,N_19842,N_19980);
xnor UO_2438 (O_2438,N_19919,N_19825);
or UO_2439 (O_2439,N_19929,N_19941);
or UO_2440 (O_2440,N_19941,N_19902);
nor UO_2441 (O_2441,N_19982,N_19994);
nor UO_2442 (O_2442,N_19866,N_19923);
and UO_2443 (O_2443,N_19908,N_19950);
and UO_2444 (O_2444,N_19824,N_19915);
xnor UO_2445 (O_2445,N_19802,N_19801);
and UO_2446 (O_2446,N_19867,N_19893);
xor UO_2447 (O_2447,N_19862,N_19811);
or UO_2448 (O_2448,N_19913,N_19949);
nand UO_2449 (O_2449,N_19888,N_19804);
nand UO_2450 (O_2450,N_19911,N_19916);
nor UO_2451 (O_2451,N_19979,N_19950);
and UO_2452 (O_2452,N_19835,N_19825);
nand UO_2453 (O_2453,N_19838,N_19963);
nor UO_2454 (O_2454,N_19915,N_19934);
nand UO_2455 (O_2455,N_19899,N_19865);
or UO_2456 (O_2456,N_19910,N_19824);
xnor UO_2457 (O_2457,N_19856,N_19832);
nor UO_2458 (O_2458,N_19927,N_19922);
nor UO_2459 (O_2459,N_19812,N_19891);
and UO_2460 (O_2460,N_19865,N_19867);
nor UO_2461 (O_2461,N_19905,N_19899);
or UO_2462 (O_2462,N_19878,N_19813);
nand UO_2463 (O_2463,N_19985,N_19982);
xor UO_2464 (O_2464,N_19833,N_19963);
xnor UO_2465 (O_2465,N_19858,N_19917);
and UO_2466 (O_2466,N_19920,N_19865);
nand UO_2467 (O_2467,N_19977,N_19875);
nor UO_2468 (O_2468,N_19808,N_19970);
nand UO_2469 (O_2469,N_19911,N_19968);
xnor UO_2470 (O_2470,N_19833,N_19967);
nor UO_2471 (O_2471,N_19855,N_19832);
or UO_2472 (O_2472,N_19903,N_19948);
xor UO_2473 (O_2473,N_19837,N_19904);
xor UO_2474 (O_2474,N_19996,N_19886);
and UO_2475 (O_2475,N_19878,N_19964);
and UO_2476 (O_2476,N_19927,N_19994);
nor UO_2477 (O_2477,N_19891,N_19996);
nor UO_2478 (O_2478,N_19829,N_19925);
xnor UO_2479 (O_2479,N_19817,N_19816);
nand UO_2480 (O_2480,N_19990,N_19945);
xor UO_2481 (O_2481,N_19967,N_19853);
xor UO_2482 (O_2482,N_19940,N_19904);
or UO_2483 (O_2483,N_19864,N_19980);
xnor UO_2484 (O_2484,N_19849,N_19901);
and UO_2485 (O_2485,N_19943,N_19926);
nand UO_2486 (O_2486,N_19837,N_19878);
xor UO_2487 (O_2487,N_19993,N_19933);
nor UO_2488 (O_2488,N_19871,N_19933);
or UO_2489 (O_2489,N_19855,N_19990);
and UO_2490 (O_2490,N_19818,N_19906);
nor UO_2491 (O_2491,N_19898,N_19842);
or UO_2492 (O_2492,N_19934,N_19860);
nand UO_2493 (O_2493,N_19876,N_19835);
and UO_2494 (O_2494,N_19937,N_19995);
nor UO_2495 (O_2495,N_19861,N_19813);
xnor UO_2496 (O_2496,N_19930,N_19878);
or UO_2497 (O_2497,N_19909,N_19938);
nor UO_2498 (O_2498,N_19963,N_19865);
and UO_2499 (O_2499,N_19845,N_19984);
endmodule