module basic_2000_20000_2500_125_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1517,In_1312);
nor U1 (N_1,In_108,In_1398);
nor U2 (N_2,In_1725,In_1974);
nor U3 (N_3,In_1032,In_997);
xnor U4 (N_4,In_1946,In_344);
or U5 (N_5,In_748,In_1018);
nor U6 (N_6,In_1419,In_3);
nor U7 (N_7,In_1898,In_1785);
nor U8 (N_8,In_1798,In_1962);
nand U9 (N_9,In_361,In_903);
nor U10 (N_10,In_1320,In_1815);
nor U11 (N_11,In_1707,In_1452);
or U12 (N_12,In_1835,In_276);
nand U13 (N_13,In_787,In_137);
and U14 (N_14,In_1972,In_1739);
or U15 (N_15,In_463,In_662);
xor U16 (N_16,In_798,In_1742);
nand U17 (N_17,In_135,In_1729);
nor U18 (N_18,In_1367,In_822);
xnor U19 (N_19,In_1358,In_687);
nor U20 (N_20,In_1324,In_1316);
nand U21 (N_21,In_1651,In_597);
and U22 (N_22,In_471,In_175);
xnor U23 (N_23,In_384,In_1361);
or U24 (N_24,In_1404,In_701);
nand U25 (N_25,In_582,In_1861);
xnor U26 (N_26,In_1541,In_1087);
or U27 (N_27,In_185,In_412);
or U28 (N_28,In_1104,In_692);
xor U29 (N_29,In_333,In_844);
or U30 (N_30,In_1304,In_1240);
nand U31 (N_31,In_1108,In_1003);
nand U32 (N_32,In_1378,In_159);
and U33 (N_33,In_1136,In_489);
or U34 (N_34,In_335,In_200);
and U35 (N_35,In_1868,In_677);
or U36 (N_36,In_1716,In_60);
or U37 (N_37,In_1603,In_648);
nor U38 (N_38,In_1330,In_814);
or U39 (N_39,In_1471,In_1035);
nor U40 (N_40,In_581,In_1678);
or U41 (N_41,In_771,In_1746);
xor U42 (N_42,In_1368,In_1797);
or U43 (N_43,In_759,In_317);
or U44 (N_44,In_1019,In_1227);
nor U45 (N_45,In_1990,In_1880);
and U46 (N_46,In_1936,In_741);
xor U47 (N_47,In_1736,In_70);
or U48 (N_48,In_181,In_1261);
or U49 (N_49,In_1406,In_297);
nand U50 (N_50,In_1924,In_826);
nand U51 (N_51,In_1433,In_1874);
or U52 (N_52,In_1468,In_248);
and U53 (N_53,In_31,In_643);
or U54 (N_54,In_513,In_583);
nor U55 (N_55,In_265,In_1635);
nand U56 (N_56,In_948,In_1583);
or U57 (N_57,In_1431,In_1409);
or U58 (N_58,In_1676,In_1191);
or U59 (N_59,In_1885,In_993);
or U60 (N_60,In_724,In_48);
nand U61 (N_61,In_1935,In_1429);
nand U62 (N_62,In_174,In_32);
xnor U63 (N_63,In_1118,In_1645);
nor U64 (N_64,In_1672,In_202);
nand U65 (N_65,In_1024,In_1335);
nor U66 (N_66,In_1668,In_1343);
nand U67 (N_67,In_213,In_49);
and U68 (N_68,In_1437,In_1389);
nand U69 (N_69,In_481,In_682);
and U70 (N_70,In_1467,In_473);
nand U71 (N_71,In_1410,In_1278);
nor U72 (N_72,In_1959,In_829);
and U73 (N_73,In_1669,In_1573);
and U74 (N_74,In_633,In_1511);
nand U75 (N_75,In_1077,In_1545);
xnor U76 (N_76,In_890,In_1047);
and U77 (N_77,In_622,In_1288);
and U78 (N_78,In_1253,In_732);
nand U79 (N_79,In_1753,In_504);
and U80 (N_80,In_756,In_492);
nand U81 (N_81,In_1658,In_968);
nand U82 (N_82,In_1040,In_270);
and U83 (N_83,In_495,In_1955);
nand U84 (N_84,In_877,In_305);
nand U85 (N_85,In_1366,In_994);
nor U86 (N_86,In_467,In_1958);
or U87 (N_87,In_910,In_1988);
and U88 (N_88,In_1177,In_1916);
xor U89 (N_89,In_847,In_1061);
and U90 (N_90,In_430,In_1385);
nor U91 (N_91,In_1840,In_1085);
and U92 (N_92,In_133,In_1664);
or U93 (N_93,In_414,In_1649);
xor U94 (N_94,In_201,In_1347);
xnor U95 (N_95,In_74,In_387);
nand U96 (N_96,In_1162,In_164);
xnor U97 (N_97,In_1071,In_1720);
xnor U98 (N_98,In_1355,In_1801);
nand U99 (N_99,In_1580,In_862);
or U100 (N_100,In_1770,In_1257);
or U101 (N_101,In_1620,In_239);
nand U102 (N_102,In_1397,In_1561);
and U103 (N_103,In_337,In_864);
or U104 (N_104,In_725,In_22);
or U105 (N_105,In_792,In_243);
or U106 (N_106,In_1263,In_1457);
or U107 (N_107,In_965,In_71);
or U108 (N_108,In_589,In_1439);
xor U109 (N_109,In_300,In_1910);
and U110 (N_110,In_1284,In_571);
xnor U111 (N_111,In_702,In_925);
nand U112 (N_112,In_331,In_620);
nand U113 (N_113,In_1585,In_1799);
nor U114 (N_114,In_720,In_1233);
and U115 (N_115,In_519,In_617);
or U116 (N_116,In_416,In_1554);
and U117 (N_117,In_982,In_5);
nor U118 (N_118,In_221,In_686);
nor U119 (N_119,In_1947,In_1841);
nor U120 (N_120,In_1758,In_256);
xor U121 (N_121,In_418,In_894);
or U122 (N_122,In_1391,In_1349);
and U123 (N_123,In_1838,In_809);
or U124 (N_124,In_1154,In_1530);
xor U125 (N_125,In_611,In_1734);
nand U126 (N_126,In_751,In_38);
xnor U127 (N_127,In_421,In_143);
xor U128 (N_128,In_1951,In_1460);
xor U129 (N_129,In_909,In_1048);
and U130 (N_130,In_56,In_99);
or U131 (N_131,In_605,In_619);
nor U132 (N_132,In_1377,In_1986);
nor U133 (N_133,In_1379,In_775);
nor U134 (N_134,In_1522,In_296);
xor U135 (N_135,In_314,In_1172);
nand U136 (N_136,In_721,In_247);
and U137 (N_137,In_2,In_1265);
nand U138 (N_138,In_111,In_394);
nor U139 (N_139,In_1748,In_1450);
nand U140 (N_140,In_1703,In_584);
nand U141 (N_141,In_911,In_1081);
and U142 (N_142,In_98,In_816);
nor U143 (N_143,In_642,In_293);
xnor U144 (N_144,In_1507,In_550);
xnor U145 (N_145,In_180,In_570);
or U146 (N_146,In_1917,In_1111);
or U147 (N_147,In_112,In_943);
or U148 (N_148,In_1991,In_674);
xnor U149 (N_149,In_1808,In_183);
or U150 (N_150,In_229,In_1211);
and U151 (N_151,In_1694,In_469);
nand U152 (N_152,In_1934,In_659);
nand U153 (N_153,In_374,In_93);
nand U154 (N_154,In_1667,In_241);
nand U155 (N_155,In_291,In_884);
nor U156 (N_156,In_845,In_288);
nand U157 (N_157,In_1440,In_260);
xor U158 (N_158,In_1836,In_1247);
nand U159 (N_159,In_553,In_419);
nor U160 (N_160,In_426,In_1380);
xor U161 (N_161,In_197,In_1960);
or U162 (N_162,In_743,In_1228);
or U163 (N_163,In_271,In_710);
xnor U164 (N_164,In_472,In_969);
xor U165 (N_165,In_1775,In_476);
nand U166 (N_166,In_290,In_783);
xnor U167 (N_167,In_433,In_1351);
xnor U168 (N_168,In_371,In_1607);
nor U169 (N_169,In_1093,In_134);
and U170 (N_170,In_514,In_1096);
xnor U171 (N_171,In_744,In_992);
and U172 (N_172,In_530,In_1549);
or U173 (N_173,In_1559,In_1867);
xor U174 (N_174,In_364,In_1403);
xnor U175 (N_175,N_92,In_1090);
and U176 (N_176,N_48,In_577);
and U177 (N_177,In_1560,In_634);
or U178 (N_178,In_409,In_1188);
nor U179 (N_179,In_1921,In_540);
xor U180 (N_180,In_964,In_306);
or U181 (N_181,In_1839,In_1014);
and U182 (N_182,In_1639,In_304);
or U183 (N_183,In_1383,In_977);
or U184 (N_184,In_1183,In_1809);
and U185 (N_185,In_781,In_1943);
nor U186 (N_186,In_151,In_474);
xor U187 (N_187,In_36,In_1225);
or U188 (N_188,In_155,In_389);
xor U189 (N_189,In_1857,N_115);
and U190 (N_190,In_1870,In_1715);
and U191 (N_191,In_630,In_1072);
nor U192 (N_192,In_1570,In_1526);
nand U193 (N_193,In_1311,In_897);
nor U194 (N_194,In_1689,In_1806);
and U195 (N_195,N_17,In_208);
nand U196 (N_196,In_1337,In_1903);
nand U197 (N_197,In_753,In_1594);
xor U198 (N_198,In_1661,In_1466);
or U199 (N_199,N_145,In_493);
nand U200 (N_200,In_113,In_1193);
nand U201 (N_201,In_1281,In_1473);
and U202 (N_202,In_1376,In_315);
nor U203 (N_203,In_1074,In_1558);
and U204 (N_204,In_295,In_233);
nor U205 (N_205,N_85,In_1137);
or U206 (N_206,In_652,In_1474);
nor U207 (N_207,In_908,In_560);
nand U208 (N_208,In_1975,In_33);
or U209 (N_209,In_178,In_244);
xnor U210 (N_210,In_848,In_654);
nand U211 (N_211,In_1904,In_951);
and U212 (N_212,In_850,In_1387);
xnor U213 (N_213,In_1519,In_486);
nor U214 (N_214,In_507,In_1322);
nor U215 (N_215,In_1723,In_1502);
or U216 (N_216,N_112,In_1218);
nand U217 (N_217,In_1480,In_670);
nor U218 (N_218,In_334,In_719);
nor U219 (N_219,In_127,In_945);
xnor U220 (N_220,In_1789,N_127);
xnor U221 (N_221,In_1185,In_1568);
or U222 (N_222,In_576,In_1267);
or U223 (N_223,In_1527,In_891);
or U224 (N_224,In_711,In_480);
nor U225 (N_225,In_776,In_1037);
xor U226 (N_226,In_1538,In_1360);
nor U227 (N_227,In_813,In_1976);
xnor U228 (N_228,In_1684,N_140);
or U229 (N_229,In_203,N_121);
nand U230 (N_230,In_539,In_382);
nor U231 (N_231,In_920,In_846);
nor U232 (N_232,In_1636,In_1339);
or U233 (N_233,In_146,In_1971);
nor U234 (N_234,In_673,In_534);
and U235 (N_235,In_252,In_100);
nor U236 (N_236,In_1083,In_1245);
or U237 (N_237,In_1407,In_1189);
or U238 (N_238,In_1279,In_1053);
nor U239 (N_239,In_967,In_258);
xor U240 (N_240,In_1015,In_407);
nand U241 (N_241,In_1531,In_57);
or U242 (N_242,In_896,In_1750);
xor U243 (N_243,N_44,In_1685);
xnor U244 (N_244,In_1057,In_986);
and U245 (N_245,In_50,In_696);
xnor U246 (N_246,In_1925,In_54);
nor U247 (N_247,In_1630,In_470);
nor U248 (N_248,In_1158,In_957);
nand U249 (N_249,In_1484,N_50);
or U250 (N_250,N_41,In_666);
nor U251 (N_251,In_1747,In_512);
or U252 (N_252,In_1028,In_215);
nand U253 (N_253,In_918,In_212);
nand U254 (N_254,In_1408,In_90);
nor U255 (N_255,In_1855,In_1321);
xor U256 (N_256,In_1130,In_429);
and U257 (N_257,In_1565,In_851);
nor U258 (N_258,In_780,In_704);
and U259 (N_259,In_1231,In_1049);
and U260 (N_260,In_1039,In_614);
nand U261 (N_261,In_515,N_133);
nor U262 (N_262,In_52,In_447);
nand U263 (N_263,In_1906,In_1209);
nand U264 (N_264,In_1851,In_1660);
or U265 (N_265,N_79,N_64);
and U266 (N_266,In_689,In_811);
or U267 (N_267,In_1127,In_464);
nand U268 (N_268,In_1881,In_1613);
and U269 (N_269,In_795,In_511);
nor U270 (N_270,N_9,In_591);
xnor U271 (N_271,In_703,In_912);
nand U272 (N_272,In_535,In_1411);
or U273 (N_273,In_1886,In_259);
nor U274 (N_274,N_114,In_1082);
and U275 (N_275,In_313,In_556);
or U276 (N_276,In_1598,In_217);
and U277 (N_277,In_349,In_1301);
xnor U278 (N_278,In_1864,In_681);
nand U279 (N_279,In_1950,In_938);
nand U280 (N_280,In_655,In_263);
nor U281 (N_281,In_179,In_1606);
nand U282 (N_282,In_1711,In_638);
nand U283 (N_283,In_1068,In_1291);
and U284 (N_284,N_28,N_35);
nand U285 (N_285,In_508,In_1126);
or U286 (N_286,In_541,In_210);
nor U287 (N_287,In_1800,In_1241);
nand U288 (N_288,In_1547,In_559);
xor U289 (N_289,In_301,In_1119);
xor U290 (N_290,In_207,In_1728);
or U291 (N_291,In_1315,In_1016);
nand U292 (N_292,N_36,In_927);
xnor U293 (N_293,In_1712,In_1425);
xor U294 (N_294,In_1171,In_1303);
nand U295 (N_295,In_1372,In_144);
and U296 (N_296,In_1120,In_859);
xnor U297 (N_297,In_947,In_251);
nor U298 (N_298,In_479,In_1940);
nand U299 (N_299,In_747,In_697);
or U300 (N_300,In_1076,In_1997);
nand U301 (N_301,In_698,In_1138);
and U302 (N_302,N_77,N_5);
and U303 (N_303,In_237,In_328);
or U304 (N_304,In_1751,In_405);
and U305 (N_305,N_60,In_799);
nor U306 (N_306,In_445,In_1113);
xor U307 (N_307,In_356,In_145);
nor U308 (N_308,In_1441,In_1807);
xor U309 (N_309,In_600,In_1198);
nor U310 (N_310,In_1160,N_99);
and U311 (N_311,In_932,In_841);
nand U312 (N_312,In_522,In_316);
and U313 (N_313,In_922,In_1948);
and U314 (N_314,In_1516,In_773);
nor U315 (N_315,In_1783,In_941);
or U316 (N_316,In_726,In_462);
xnor U317 (N_317,In_205,In_294);
or U318 (N_318,In_122,In_461);
xnor U319 (N_319,In_285,In_1978);
xor U320 (N_320,In_1447,In_1796);
nand U321 (N_321,In_119,In_1994);
and U322 (N_322,In_76,In_272);
xor U323 (N_323,In_1006,In_1067);
or U324 (N_324,In_1289,N_275);
or U325 (N_325,In_339,In_959);
or U326 (N_326,In_1030,In_746);
nor U327 (N_327,In_61,In_765);
nor U328 (N_328,In_1611,N_131);
or U329 (N_329,In_1930,In_1213);
xnor U330 (N_330,N_82,N_113);
or U331 (N_331,In_1744,In_1495);
xnor U332 (N_332,In_1812,In_46);
nor U333 (N_333,In_53,In_1862);
and U334 (N_334,In_393,In_1998);
and U335 (N_335,In_1095,In_456);
and U336 (N_336,In_284,In_1226);
and U337 (N_337,N_201,In_1369);
nand U338 (N_338,In_1135,In_1069);
nand U339 (N_339,In_1010,N_153);
xor U340 (N_340,In_678,In_160);
nand U341 (N_341,In_1766,In_41);
nor U342 (N_342,In_1309,In_824);
xor U343 (N_343,In_1833,In_656);
and U344 (N_344,N_63,In_273);
nand U345 (N_345,In_401,In_955);
xnor U346 (N_346,In_1614,In_1764);
or U347 (N_347,In_353,In_105);
nor U348 (N_348,In_234,In_1727);
xor U349 (N_349,In_1816,In_101);
or U350 (N_350,In_970,In_1989);
or U351 (N_351,In_1422,In_1179);
or U352 (N_352,In_1506,In_11);
and U353 (N_353,In_590,In_173);
and U354 (N_354,In_1164,In_936);
or U355 (N_355,In_1326,In_1187);
nand U356 (N_356,In_510,In_245);
and U357 (N_357,In_902,N_255);
and U358 (N_358,In_1207,In_691);
and U359 (N_359,In_1724,In_1600);
xnor U360 (N_360,In_1416,In_132);
nand U361 (N_361,In_1325,N_307);
xor U362 (N_362,In_1999,In_341);
xor U363 (N_363,In_1283,N_154);
xnor U364 (N_364,N_88,In_1737);
nor U365 (N_365,In_1754,In_1306);
or U366 (N_366,In_1681,N_190);
nand U367 (N_367,In_729,In_1670);
and U368 (N_368,In_1626,N_24);
nor U369 (N_369,In_365,N_176);
xor U370 (N_370,In_230,In_114);
xnor U371 (N_371,In_1967,In_1979);
nor U372 (N_372,In_1033,In_1299);
nand U373 (N_373,In_96,In_1749);
or U374 (N_374,In_1772,In_1515);
xor U375 (N_375,In_1503,In_924);
xnor U376 (N_376,In_601,In_867);
xnor U377 (N_377,In_1790,In_1501);
and U378 (N_378,In_806,In_665);
nor U379 (N_379,In_1273,In_264);
and U380 (N_380,In_299,N_18);
nand U381 (N_381,In_713,In_1638);
or U382 (N_382,N_149,In_618);
nand U383 (N_383,In_1248,In_423);
or U384 (N_384,In_901,In_1157);
nor U385 (N_385,In_1810,In_563);
xnor U386 (N_386,In_27,N_199);
or U387 (N_387,N_216,In_573);
nand U388 (N_388,In_1755,In_1025);
nand U389 (N_389,In_989,In_1919);
or U390 (N_390,In_1295,N_30);
or U391 (N_391,N_266,In_1652);
and U392 (N_392,In_1091,In_1846);
nand U393 (N_393,In_63,In_1964);
nor U394 (N_394,In_336,In_1827);
nand U395 (N_395,In_383,In_303);
nor U396 (N_396,In_1463,In_836);
or U397 (N_397,In_1202,In_1182);
or U398 (N_398,In_152,In_685);
nor U399 (N_399,In_1918,In_87);
or U400 (N_400,In_1644,In_40);
or U401 (N_401,In_1390,In_631);
nor U402 (N_402,In_1788,In_913);
nand U403 (N_403,In_855,In_565);
and U404 (N_404,In_1292,In_1493);
nor U405 (N_405,N_134,In_1535);
or U406 (N_406,In_422,In_167);
and U407 (N_407,In_608,In_424);
nor U408 (N_408,N_252,In_899);
xnor U409 (N_409,N_135,N_251);
nand U410 (N_410,In_1144,In_868);
nand U411 (N_411,In_973,In_1174);
nand U412 (N_412,In_502,In_453);
or U413 (N_413,In_588,N_284);
nor U414 (N_414,In_1587,In_398);
xnor U415 (N_415,In_1084,In_1927);
xor U416 (N_416,In_1201,N_297);
nand U417 (N_417,In_359,N_246);
or U418 (N_418,N_236,In_794);
and U419 (N_419,In_983,In_1062);
and U420 (N_420,In_219,In_1696);
nor U421 (N_421,N_47,In_518);
and U422 (N_422,In_1622,In_1740);
nor U423 (N_423,In_1317,In_1872);
and U424 (N_424,In_649,In_1181);
or U425 (N_425,N_7,In_465);
xor U426 (N_426,In_446,N_299);
nand U427 (N_427,N_119,N_301);
xnor U428 (N_428,In_1963,N_312);
and U429 (N_429,In_1856,In_420);
xor U430 (N_430,In_278,In_820);
and U431 (N_431,In_1610,In_1743);
nand U432 (N_432,In_193,In_1627);
nand U433 (N_433,In_1131,In_1066);
and U434 (N_434,In_1145,In_1784);
nor U435 (N_435,In_8,In_839);
xnor U436 (N_436,N_150,In_980);
or U437 (N_437,N_293,N_291);
nor U438 (N_438,In_1534,In_190);
and U439 (N_439,N_211,In_1509);
nand U440 (N_440,N_230,In_1643);
and U441 (N_441,In_255,In_999);
nor U442 (N_442,In_1052,N_142);
and U443 (N_443,In_1887,N_217);
and U444 (N_444,N_295,In_1352);
nand U445 (N_445,N_270,N_62);
and U446 (N_446,In_575,In_808);
nand U447 (N_447,In_1341,N_225);
and U448 (N_448,N_90,In_1246);
and U449 (N_449,In_517,In_123);
or U450 (N_450,N_292,In_157);
or U451 (N_451,N_12,In_1548);
nor U452 (N_452,In_934,In_138);
or U453 (N_453,In_1498,In_72);
xnor U454 (N_454,In_1114,N_179);
nor U455 (N_455,In_1673,In_604);
or U456 (N_456,In_1953,In_330);
and U457 (N_457,In_683,In_1605);
nand U458 (N_458,N_38,In_843);
or U459 (N_459,In_397,In_1254);
and U460 (N_460,In_222,In_529);
xor U461 (N_461,N_314,In_236);
nor U462 (N_462,In_366,In_13);
and U463 (N_463,In_1128,In_158);
xor U464 (N_464,In_802,In_253);
or U465 (N_465,In_1562,In_1448);
nand U466 (N_466,In_1161,In_1704);
xnor U467 (N_467,In_1877,N_203);
xnor U468 (N_468,N_296,In_694);
or U469 (N_469,In_893,In_417);
and U470 (N_470,In_17,In_521);
xnor U471 (N_471,In_385,N_287);
and U472 (N_472,In_1826,In_857);
and U473 (N_473,In_1250,In_1031);
nor U474 (N_474,In_1995,In_1539);
xor U475 (N_475,N_243,In_214);
xor U476 (N_476,N_78,N_202);
and U477 (N_477,In_0,In_7);
or U478 (N_478,In_231,N_194);
and U479 (N_479,In_1259,In_1396);
and U480 (N_480,In_579,In_1017);
nand U481 (N_481,In_196,N_249);
nand U482 (N_482,In_1821,In_572);
or U483 (N_483,In_1532,In_926);
nor U484 (N_484,N_477,N_185);
xor U485 (N_485,In_1794,In_156);
and U486 (N_486,In_1888,In_378);
and U487 (N_487,N_231,In_1370);
or U488 (N_488,N_374,In_546);
xnor U489 (N_489,In_232,N_22);
xnor U490 (N_490,In_1640,In_1494);
and U491 (N_491,N_120,In_764);
nand U492 (N_492,N_256,In_990);
and U493 (N_493,In_532,In_1103);
and U494 (N_494,In_1593,In_668);
xor U495 (N_495,In_131,In_1388);
nand U496 (N_496,N_55,In_1345);
or U497 (N_497,N_300,In_380);
or U498 (N_498,N_180,In_223);
nor U499 (N_499,N_136,In_533);
or U500 (N_500,In_292,In_77);
nor U501 (N_501,In_1581,In_399);
and U502 (N_502,N_171,N_37);
xnor U503 (N_503,In_1615,N_89);
nor U504 (N_504,In_568,In_501);
nor U505 (N_505,In_1665,In_369);
or U506 (N_506,In_483,In_1086);
nor U507 (N_507,In_1708,In_162);
nor U508 (N_508,In_825,N_110);
xor U509 (N_509,In_88,In_1782);
nor U510 (N_510,N_161,N_43);
and U511 (N_511,In_147,N_338);
nor U512 (N_512,In_796,N_101);
xor U513 (N_513,In_628,N_274);
xnor U514 (N_514,In_1344,In_396);
nand U515 (N_515,In_1786,N_466);
or U516 (N_516,In_391,N_80);
and U517 (N_517,In_931,In_1869);
nor U518 (N_518,In_834,N_235);
nand U519 (N_519,In_738,In_1346);
and U520 (N_520,In_199,In_632);
nor U521 (N_521,In_705,In_449);
nor U522 (N_522,In_693,N_168);
nor U523 (N_523,In_1243,In_593);
and U524 (N_524,N_67,In_1599);
nor U525 (N_525,N_322,In_1500);
nand U526 (N_526,N_118,N_162);
and U527 (N_527,In_154,In_351);
xnor U528 (N_528,In_623,In_1980);
or U529 (N_529,In_1269,N_364);
nand U530 (N_530,In_1075,N_264);
nand U531 (N_531,N_206,In_195);
and U532 (N_532,In_1297,N_159);
and U533 (N_533,N_424,In_370);
nand U534 (N_534,N_105,N_347);
xor U535 (N_535,In_805,In_404);
and U536 (N_536,In_606,In_500);
nand U537 (N_537,N_265,In_1146);
and U538 (N_538,In_684,In_1204);
or U539 (N_539,In_372,In_1834);
and U540 (N_540,In_224,In_1180);
nor U541 (N_541,In_345,In_1757);
or U542 (N_542,In_66,In_832);
and U543 (N_543,In_1543,In_1588);
and U544 (N_544,In_283,In_254);
or U545 (N_545,In_1491,In_1470);
or U546 (N_546,In_1675,N_366);
nand U547 (N_547,In_165,N_315);
nor U548 (N_548,In_1731,In_1569);
xor U549 (N_549,In_1000,In_59);
nand U550 (N_550,N_317,In_695);
xor U551 (N_551,In_1151,In_438);
nand U552 (N_552,In_1464,N_373);
or U553 (N_553,N_289,N_237);
xor U554 (N_554,In_346,In_586);
nand U555 (N_555,In_170,N_220);
nor U556 (N_556,In_1551,N_467);
and U557 (N_557,In_1307,N_124);
nor U558 (N_558,In_1483,In_332);
nor U559 (N_559,In_1893,N_412);
and U560 (N_560,In_1909,In_1595);
or U561 (N_561,In_1098,N_31);
xor U562 (N_562,In_488,In_413);
xnor U563 (N_563,In_1051,In_789);
nand U564 (N_564,In_1780,In_1700);
nor U565 (N_565,In_368,In_406);
or U566 (N_566,In_837,In_878);
xor U567 (N_567,In_906,In_1891);
and U568 (N_568,In_706,In_117);
xor U569 (N_569,In_1106,In_774);
xnor U570 (N_570,In_1741,In_1894);
nand U571 (N_571,N_298,In_1695);
and U572 (N_572,In_1628,In_1333);
and U573 (N_573,In_779,N_81);
nand U574 (N_574,In_815,N_33);
or U575 (N_575,N_406,In_527);
nor U576 (N_576,In_885,In_621);
xnor U577 (N_577,In_1064,In_1271);
and U578 (N_578,In_1802,In_1913);
or U579 (N_579,In_1592,In_452);
or U580 (N_580,N_416,N_87);
or U581 (N_581,In_1621,N_15);
nor U582 (N_582,In_1186,N_248);
or U583 (N_583,In_1987,In_1659);
or U584 (N_584,N_97,In_1196);
nor U585 (N_585,N_458,In_95);
or U586 (N_586,In_1818,N_263);
nor U587 (N_587,N_109,In_946);
xor U588 (N_588,In_707,In_64);
or U589 (N_589,In_1080,In_436);
xor U590 (N_590,N_473,N_268);
nand U591 (N_591,In_1625,In_1199);
nor U592 (N_592,In_42,In_1314);
or U593 (N_593,In_1911,In_1134);
and U594 (N_594,In_1323,In_1602);
nand U595 (N_595,In_950,In_1022);
nor U596 (N_596,In_1451,N_376);
and U597 (N_597,In_1327,In_1901);
nand U598 (N_598,In_1928,In_1476);
nor U599 (N_599,In_1216,In_1996);
xor U600 (N_600,In_444,In_1843);
nand U601 (N_601,In_1336,In_103);
nand U602 (N_602,In_599,N_65);
and U603 (N_603,In_1567,N_215);
nor U604 (N_604,In_325,N_382);
xnor U605 (N_605,In_400,In_1497);
or U606 (N_606,In_1873,N_448);
nor U607 (N_607,In_496,In_737);
nor U608 (N_608,In_250,In_1969);
xnor U609 (N_609,In_937,In_307);
nand U610 (N_610,In_933,In_1733);
and U611 (N_611,In_1296,In_875);
nor U612 (N_612,N_93,In_731);
xor U613 (N_613,In_1932,In_1683);
and U614 (N_614,In_835,In_440);
or U615 (N_615,N_423,In_1722);
nor U616 (N_616,In_431,N_344);
or U617 (N_617,In_1642,In_876);
nor U618 (N_618,N_333,In_730);
xor U619 (N_619,In_68,In_1884);
nor U620 (N_620,In_1590,In_435);
nand U621 (N_621,N_102,In_1102);
and U622 (N_622,In_1706,In_1426);
or U623 (N_623,In_1272,In_1771);
and U624 (N_624,In_381,In_39);
xor U625 (N_625,In_1584,In_1435);
and U626 (N_626,In_246,In_1637);
nand U627 (N_627,N_413,N_74);
or U628 (N_628,N_447,N_1);
nor U629 (N_629,In_110,In_942);
or U630 (N_630,N_422,In_425);
or U631 (N_631,In_958,N_470);
xor U632 (N_632,In_30,In_840);
and U633 (N_633,In_83,In_51);
and U634 (N_634,In_1957,In_1858);
nand U635 (N_635,N_455,N_151);
and U636 (N_636,N_371,In_1036);
xor U637 (N_637,In_82,In_1359);
nand U638 (N_638,N_173,In_1300);
and U639 (N_639,In_1005,In_1671);
nand U640 (N_640,In_1155,In_1449);
or U641 (N_641,In_1779,N_362);
nand U642 (N_642,In_358,In_1277);
or U643 (N_643,In_1690,In_1482);
nand U644 (N_644,In_679,In_1804);
xnor U645 (N_645,N_407,In_557);
or U646 (N_646,In_1899,N_582);
xor U647 (N_647,In_242,In_140);
or U648 (N_648,In_1550,N_303);
nor U649 (N_649,In_1041,In_1523);
xnor U650 (N_650,In_1462,In_1973);
or U651 (N_651,In_347,N_69);
nand U652 (N_652,In_1148,In_1831);
and U653 (N_653,In_1329,In_972);
nor U654 (N_654,N_245,In_739);
xnor U655 (N_655,N_386,In_1674);
and U656 (N_656,In_1229,N_95);
xor U657 (N_657,N_508,In_189);
or U658 (N_658,In_1401,In_1260);
nand U659 (N_659,In_240,In_1465);
and U660 (N_660,N_355,In_1354);
and U661 (N_661,N_613,In_1662);
nand U662 (N_662,N_535,In_1860);
nand U663 (N_663,In_1822,In_1115);
or U664 (N_664,In_1849,In_1063);
nor U665 (N_665,N_599,In_900);
and U666 (N_666,N_392,In_1097);
and U667 (N_667,In_1150,In_717);
xor U668 (N_668,N_6,N_241);
xor U669 (N_669,N_184,In_1778);
or U670 (N_670,In_1163,N_148);
and U671 (N_671,In_1692,In_1124);
xor U672 (N_672,In_79,In_1865);
nand U673 (N_673,In_544,In_1769);
or U674 (N_674,N_327,In_238);
and U675 (N_675,In_410,N_116);
xnor U676 (N_676,N_579,In_1184);
nor U677 (N_677,In_1079,In_321);
nand U678 (N_678,In_1170,In_1985);
nor U679 (N_679,N_369,N_603);
xnor U680 (N_680,In_612,In_858);
xnor U681 (N_681,N_581,In_1752);
nor U682 (N_682,N_61,N_519);
nand U683 (N_683,N_638,In_1045);
and U684 (N_684,N_546,In_1828);
and U685 (N_685,In_24,In_120);
nor U686 (N_686,In_1572,In_657);
xor U687 (N_687,N_21,In_257);
nor U688 (N_688,N_523,In_791);
nand U689 (N_689,In_803,In_1208);
nor U690 (N_690,In_1803,In_1952);
nor U691 (N_691,In_1302,N_612);
or U692 (N_692,N_342,In_1011);
and U693 (N_693,In_979,N_637);
and U694 (N_694,In_852,In_1166);
xor U695 (N_695,In_1481,N_586);
or U696 (N_696,In_1854,In_833);
xor U697 (N_697,In_1001,N_469);
xor U698 (N_698,In_1489,In_1399);
nor U699 (N_699,In_29,In_1415);
and U700 (N_700,In_784,N_26);
and U701 (N_701,In_261,N_106);
nor U702 (N_702,In_62,In_377);
nor U703 (N_703,N_528,N_506);
xnor U704 (N_704,In_1105,In_1374);
xnor U705 (N_705,In_1402,In_733);
or U706 (N_706,In_1656,N_427);
nor U707 (N_707,N_486,N_221);
xnor U708 (N_708,In_1938,N_304);
nand U709 (N_709,In_661,N_187);
xor U710 (N_710,In_963,In_498);
nor U711 (N_711,In_1109,In_1478);
nand U712 (N_712,In_1552,N_415);
or U713 (N_713,N_379,In_1863);
and U714 (N_714,In_506,N_381);
xor U715 (N_715,In_1206,In_749);
nor U716 (N_716,In_1176,In_1249);
nand U717 (N_717,N_489,N_429);
nor U718 (N_718,In_863,In_129);
nand U719 (N_719,In_326,In_375);
xor U720 (N_720,In_520,In_136);
or U721 (N_721,N_491,In_499);
nor U722 (N_722,N_476,N_547);
nor U723 (N_723,In_1900,N_308);
xor U724 (N_724,N_192,N_388);
nor U725 (N_725,In_402,N_417);
nand U726 (N_726,In_1054,N_498);
xor U727 (N_727,In_728,N_224);
nand U728 (N_728,N_590,In_1939);
or U729 (N_729,In_960,In_1937);
nand U730 (N_730,N_393,In_763);
nor U731 (N_731,In_1905,N_479);
or U732 (N_732,N_593,In_477);
and U733 (N_733,In_1424,In_130);
and U734 (N_734,In_308,In_1143);
or U735 (N_735,In_4,In_128);
or U736 (N_736,In_355,N_279);
nor U737 (N_737,N_269,In_1612);
nand U738 (N_738,N_580,N_2);
or U739 (N_739,In_785,N_98);
xnor U740 (N_740,In_777,N_219);
nor U741 (N_741,In_949,N_227);
and U742 (N_742,N_513,In_1009);
or U743 (N_743,In_1023,In_817);
xnor U744 (N_744,In_1167,In_675);
nand U745 (N_745,In_1871,N_282);
xnor U746 (N_746,In_1485,In_1853);
and U747 (N_747,In_1710,N_551);
and U748 (N_748,N_499,In_1713);
xnor U749 (N_749,In_1702,N_32);
nor U750 (N_750,In_1825,N_343);
xor U751 (N_751,N_401,N_45);
nand U752 (N_752,N_618,In_1697);
nor U753 (N_753,In_558,In_923);
nor U754 (N_754,In_625,N_167);
xor U755 (N_755,In_548,In_842);
or U756 (N_756,In_889,In_466);
or U757 (N_757,In_818,In_1837);
nand U758 (N_758,In_1443,In_991);
nor U759 (N_759,In_536,In_650);
and U760 (N_760,In_1056,N_639);
or U761 (N_761,In_865,In_43);
nand U762 (N_762,N_398,N_285);
nor U763 (N_763,In_329,N_370);
nor U764 (N_764,In_459,In_757);
and U765 (N_765,In_121,In_18);
nor U766 (N_766,In_1629,In_281);
xnor U767 (N_767,N_213,In_286);
and U768 (N_768,N_400,In_1721);
and U769 (N_769,In_227,N_205);
nor U770 (N_770,N_563,In_287);
and U771 (N_771,In_85,In_1647);
nor U772 (N_772,In_1197,In_549);
and U773 (N_773,In_646,N_250);
xor U774 (N_774,In_1002,In_1895);
and U775 (N_775,In_194,In_944);
or U776 (N_776,In_1342,In_1381);
or U777 (N_777,In_566,In_153);
and U778 (N_778,N_441,In_1586);
nor U779 (N_779,N_390,In_1153);
and U780 (N_780,In_641,N_143);
or U781 (N_781,In_266,In_1305);
nor U782 (N_782,In_1528,In_124);
or U783 (N_783,In_554,In_1933);
or U784 (N_784,In_1582,In_669);
nand U785 (N_785,In_770,In_1405);
nand U786 (N_786,N_434,N_40);
xor U787 (N_787,N_170,In_1842);
and U788 (N_788,In_1576,In_874);
or U789 (N_789,In_1892,In_503);
nor U790 (N_790,N_411,N_571);
nor U791 (N_791,N_404,In_1116);
or U792 (N_792,In_1107,In_984);
or U793 (N_793,N_261,In_561);
or U794 (N_794,In_598,N_541);
nand U795 (N_795,In_1472,N_527);
or U796 (N_796,N_622,In_531);
xor U797 (N_797,In_228,In_1577);
and U798 (N_798,N_286,In_390);
nand U799 (N_799,In_1357,In_1824);
nand U800 (N_800,In_109,N_737);
nor U801 (N_801,N_643,N_776);
xnor U802 (N_802,In_367,N_218);
or U803 (N_803,N_329,In_1121);
xnor U804 (N_804,In_302,N_544);
or U805 (N_805,In_1112,In_1508);
xnor U806 (N_806,N_208,In_1915);
xor U807 (N_807,N_346,In_1286);
and U808 (N_808,N_52,N_352);
or U809 (N_809,N_550,In_595);
or U810 (N_810,In_542,In_1793);
xor U811 (N_811,N_664,N_280);
nor U812 (N_812,In_277,In_974);
and U813 (N_813,N_389,In_1945);
and U814 (N_814,In_663,In_25);
nand U815 (N_815,In_1845,N_538);
xor U816 (N_816,N_70,In_1275);
nand U817 (N_817,N_126,N_620);
xnor U818 (N_818,In_860,N_679);
and U819 (N_819,N_59,In_115);
nand U820 (N_820,N_799,In_988);
or U821 (N_821,In_1129,In_21);
and U822 (N_822,In_340,In_1663);
and U823 (N_823,N_34,In_1393);
or U824 (N_824,In_709,N_751);
and U825 (N_825,In_75,In_1691);
nor U826 (N_826,In_1012,In_1088);
or U827 (N_827,N_27,N_531);
nor U828 (N_828,N_648,N_661);
or U829 (N_829,N_645,In_1469);
or U830 (N_830,In_443,In_1709);
or U831 (N_831,In_150,N_597);
and U832 (N_832,N_439,In_279);
and U833 (N_833,N_774,N_450);
xnor U834 (N_834,In_1459,N_768);
or U835 (N_835,In_343,In_1596);
or U836 (N_836,N_340,In_1008);
xor U837 (N_837,In_1256,In_1026);
nand U838 (N_838,N_653,N_226);
and U839 (N_839,N_516,N_775);
and U840 (N_840,N_330,In_1505);
nor U841 (N_841,In_626,In_1220);
nor U842 (N_842,In_690,In_742);
and U843 (N_843,In_1479,N_475);
nand U844 (N_844,In_34,In_441);
and U845 (N_845,In_745,N_743);
xnor U846 (N_846,In_1897,In_879);
and U847 (N_847,In_1859,N_591);
xnor U848 (N_848,N_572,N_526);
or U849 (N_849,In_274,In_939);
or U850 (N_850,N_695,In_1252);
nor U851 (N_851,In_455,N_445);
xor U852 (N_852,In_672,In_551);
nand U853 (N_853,N_565,N_144);
and U854 (N_854,In_1878,N_607);
or U855 (N_855,In_562,In_1941);
and U856 (N_856,In_1537,N_693);
nor U857 (N_857,In_1092,In_1236);
nor U858 (N_858,In_1499,In_1239);
or U859 (N_859,N_460,In_1169);
or U860 (N_860,In_1616,N_524);
and U861 (N_861,In_768,In_1641);
nand U862 (N_862,N_56,N_644);
xor U863 (N_863,N_501,In_1194);
nor U864 (N_864,In_1089,N_186);
nand U865 (N_865,N_574,In_1875);
xor U866 (N_866,N_358,N_332);
nand U867 (N_867,N_178,In_211);
xor U868 (N_868,N_487,In_1929);
nor U869 (N_869,In_1421,In_182);
and U870 (N_870,N_86,In_1823);
and U871 (N_871,N_662,N_738);
nand U872 (N_872,In_880,N_503);
or U873 (N_873,N_481,N_354);
and U874 (N_874,In_1065,In_1428);
or U875 (N_875,In_1332,In_482);
nor U876 (N_876,In_607,N_686);
nand U877 (N_877,In_904,N_474);
nor U878 (N_878,In_104,N_708);
nand U879 (N_879,N_552,N_71);
xnor U880 (N_880,In_450,N_387);
or U881 (N_881,N_517,N_172);
nand U882 (N_882,In_1830,N_583);
nor U883 (N_883,In_1525,N_309);
and U884 (N_884,In_676,In_1414);
nand U885 (N_885,N_518,In_395);
nor U886 (N_886,N_537,N_363);
nand U887 (N_887,In_1717,In_1190);
xor U888 (N_888,N_646,In_790);
nand U889 (N_889,N_57,In_1544);
and U890 (N_890,N_244,In_1215);
xnor U891 (N_891,In_935,In_226);
xnor U892 (N_892,In_1688,In_1285);
nor U893 (N_893,N_740,In_1234);
nor U894 (N_894,In_176,N_709);
nand U895 (N_895,In_289,In_1759);
nand U896 (N_896,In_1004,In_1222);
nand U897 (N_897,N_356,In_1968);
nor U898 (N_898,N_677,In_1266);
or U899 (N_899,In_338,N_534);
and U900 (N_900,In_1242,In_1034);
nand U901 (N_901,In_107,N_197);
nand U902 (N_902,In_1230,N_747);
nor U903 (N_903,N_426,In_1382);
and U904 (N_904,In_357,In_1591);
or U905 (N_905,In_962,N_430);
and U906 (N_906,N_259,In_930);
nor U907 (N_907,In_762,In_1262);
and U908 (N_908,In_1632,In_491);
nor U909 (N_909,In_636,In_1657);
or U910 (N_910,In_1781,N_310);
nor U911 (N_911,N_396,In_1773);
nor U912 (N_912,In_324,N_598);
xnor U913 (N_913,N_391,In_1646);
nor U914 (N_914,In_1122,N_763);
and U915 (N_915,N_688,In_1791);
or U916 (N_916,In_1504,In_1094);
or U917 (N_917,In_198,In_1223);
nand U918 (N_918,N_754,N_23);
or U919 (N_919,N_683,In_1384);
nand U920 (N_920,In_1847,N_609);
or U921 (N_921,N_335,In_475);
nand U922 (N_922,N_605,N_108);
or U923 (N_923,In_1029,N_758);
xor U924 (N_924,In_580,In_1282);
or U925 (N_925,In_1436,In_1981);
and U926 (N_926,In_886,N_351);
or U927 (N_927,In_873,In_1334);
and U928 (N_928,N_687,N_789);
or U929 (N_929,In_1521,N_626);
or U930 (N_930,In_1578,In_658);
and U931 (N_931,In_298,In_1123);
nand U932 (N_932,N_446,In_1811);
nor U933 (N_933,N_438,In_432);
nor U934 (N_934,In_1147,In_587);
or U935 (N_935,In_856,N_200);
nand U936 (N_936,In_1310,In_1255);
nand U937 (N_937,In_1922,In_187);
xnor U938 (N_938,In_1042,In_149);
and U939 (N_939,In_602,In_543);
nand U940 (N_940,In_1977,In_1070);
xor U941 (N_941,In_1574,N_242);
nand U942 (N_942,In_1908,In_1966);
nand U943 (N_943,In_142,In_172);
nor U944 (N_944,N_510,In_92);
xnor U945 (N_945,In_1876,In_1338);
nor U946 (N_946,N_785,N_4);
nor U947 (N_947,N_568,In_976);
nor U948 (N_948,N_188,In_35);
or U949 (N_949,In_1984,In_1777);
xnor U950 (N_950,In_1557,In_388);
nand U951 (N_951,In_97,In_1617);
or U952 (N_952,N_158,N_752);
or U953 (N_953,In_1013,In_940);
xor U954 (N_954,In_1513,N_659);
or U955 (N_955,In_1942,In_929);
or U956 (N_956,In_1110,N_324);
xnor U957 (N_957,N_750,N_11);
and U958 (N_958,N_104,In_1520);
nor U959 (N_959,N_339,In_1763);
and U960 (N_960,N_437,N_557);
xnor U961 (N_961,N_838,N_278);
or U962 (N_962,In_907,N_895);
and U963 (N_963,N_453,In_869);
and U964 (N_964,In_58,N_357);
xnor U965 (N_965,N_616,N_608);
or U966 (N_966,N_780,N_174);
nand U967 (N_967,N_896,In_1430);
nor U968 (N_968,N_953,N_569);
or U969 (N_969,In_1563,In_1251);
or U970 (N_970,In_769,In_1648);
xor U971 (N_971,N_20,N_919);
nand U972 (N_972,In_1510,N_228);
and U973 (N_973,N_685,In_1073);
or U974 (N_974,In_1038,N_260);
nand U975 (N_975,In_1564,N_689);
or U976 (N_976,In_1308,N_846);
xnor U977 (N_977,N_617,In_1879);
xnor U978 (N_978,N_640,N_817);
nor U979 (N_979,N_808,N_764);
or U980 (N_980,In_1152,In_592);
or U981 (N_981,N_858,In_1101);
xor U982 (N_982,In_1375,N_8);
nand U983 (N_983,In_1487,N_887);
xnor U984 (N_984,In_596,In_921);
or U985 (N_985,In_460,In_1623);
nand U986 (N_986,In_1687,In_352);
xnor U987 (N_987,N_156,N_420);
and U988 (N_988,In_1058,N_777);
xnor U989 (N_989,N_484,In_1624);
and U990 (N_990,In_786,N_769);
xnor U991 (N_991,N_111,In_699);
or U992 (N_992,In_1956,In_644);
nand U993 (N_993,In_1392,N_377);
nand U994 (N_994,N_832,N_497);
xnor U995 (N_995,N_647,In_1738);
nand U996 (N_996,N_652,N_463);
nor U997 (N_997,In_1293,N_913);
nor U998 (N_998,In_671,In_350);
or U999 (N_999,N_732,In_1417);
nor U1000 (N_1000,N_916,N_556);
or U1001 (N_1001,N_520,N_163);
nand U1002 (N_1002,N_13,In_1701);
xor U1003 (N_1003,In_249,In_1);
xor U1004 (N_1004,N_701,In_1214);
xor U1005 (N_1005,In_1258,N_103);
xnor U1006 (N_1006,N_921,In_629);
or U1007 (N_1007,N_670,In_594);
and U1008 (N_1008,In_700,N_543);
and U1009 (N_1009,In_161,In_1400);
nor U1010 (N_1010,In_1205,In_723);
nor U1011 (N_1011,N_676,In_1453);
and U1012 (N_1012,N_829,N_635);
nor U1013 (N_1013,N_191,N_421);
or U1014 (N_1014,N_806,In_603);
xnor U1015 (N_1015,N_525,In_1496);
nor U1016 (N_1016,N_691,In_1461);
nor U1017 (N_1017,N_480,In_1203);
xor U1018 (N_1018,N_828,N_319);
xor U1019 (N_1019,N_147,N_502);
xnor U1020 (N_1020,In_1666,N_650);
xnor U1021 (N_1021,In_1445,N_843);
or U1022 (N_1022,In_1395,N_428);
xor U1023 (N_1023,In_1514,In_280);
and U1024 (N_1024,N_870,N_573);
or U1025 (N_1025,N_859,N_642);
or U1026 (N_1026,N_783,N_132);
nand U1027 (N_1027,N_238,N_696);
and U1028 (N_1028,N_712,N_820);
nor U1029 (N_1029,In_65,N_958);
nand U1030 (N_1030,N_611,N_772);
or U1031 (N_1031,N_222,In_1579);
or U1032 (N_1032,In_437,N_924);
or U1033 (N_1033,N_53,In_637);
nor U1034 (N_1034,N_930,In_342);
nand U1035 (N_1035,N_901,In_1813);
and U1036 (N_1036,In_171,N_472);
xor U1037 (N_1037,In_454,N_365);
nand U1038 (N_1038,In_1931,N_871);
or U1039 (N_1039,N_629,N_883);
nand U1040 (N_1040,In_807,In_118);
and U1041 (N_1041,N_562,In_1486);
or U1042 (N_1042,In_1883,In_1597);
or U1043 (N_1043,N_578,N_10);
xor U1044 (N_1044,N_152,In_434);
xor U1045 (N_1045,N_452,In_1442);
nand U1046 (N_1046,N_779,N_853);
nand U1047 (N_1047,N_164,N_726);
xnor U1048 (N_1048,In_141,N_146);
or U1049 (N_1049,N_815,In_45);
or U1050 (N_1050,In_866,N_673);
or U1051 (N_1051,In_1961,N_936);
nand U1052 (N_1052,N_866,N_383);
nor U1053 (N_1053,In_615,N_950);
xor U1054 (N_1054,N_850,In_73);
xnor U1055 (N_1055,N_39,In_1714);
xnor U1056 (N_1056,N_567,N_731);
xor U1057 (N_1057,In_647,N_633);
or U1058 (N_1058,In_716,In_564);
nor U1059 (N_1059,In_1475,N_610);
nor U1060 (N_1060,N_440,In_478);
nor U1061 (N_1061,N_824,N_727);
or U1062 (N_1062,In_376,N_885);
or U1063 (N_1063,In_1328,N_49);
nor U1064 (N_1064,N_681,N_100);
nand U1065 (N_1065,N_781,N_394);
nor U1066 (N_1066,N_254,In_191);
nor U1067 (N_1067,In_1200,N_803);
nor U1068 (N_1068,N_945,N_770);
and U1069 (N_1069,In_1765,In_715);
nor U1070 (N_1070,In_1432,N_302);
nand U1071 (N_1071,In_1698,N_797);
nand U1072 (N_1072,In_793,In_585);
nor U1073 (N_1073,N_917,In_1235);
nor U1074 (N_1074,N_76,In_1546);
nand U1075 (N_1075,In_1682,In_1619);
nor U1076 (N_1076,N_914,In_184);
and U1077 (N_1077,N_925,In_640);
xnor U1078 (N_1078,N_418,In_269);
nand U1079 (N_1079,N_884,N_794);
and U1080 (N_1080,N_800,In_928);
or U1081 (N_1081,In_497,In_1575);
nor U1082 (N_1082,In_1745,In_1178);
nor U1083 (N_1083,In_1902,N_810);
and U1084 (N_1084,N_881,N_336);
and U1085 (N_1085,N_840,In_1244);
nor U1086 (N_1086,In_225,In_1566);
nand U1087 (N_1087,In_1168,In_1232);
and U1088 (N_1088,N_947,In_12);
nor U1089 (N_1089,N_536,N_665);
and U1090 (N_1090,N_94,In_354);
nor U1091 (N_1091,N_699,N_229);
and U1092 (N_1092,In_755,In_1007);
and U1093 (N_1093,In_1149,In_28);
nor U1094 (N_1094,In_1132,In_362);
and U1095 (N_1095,In_1173,In_1529);
and U1096 (N_1096,In_714,N_666);
and U1097 (N_1097,N_873,N_348);
nand U1098 (N_1098,N_744,In_1264);
or U1099 (N_1099,In_1444,N_29);
or U1100 (N_1100,N_504,N_325);
nor U1101 (N_1101,In_1420,In_1907);
xnor U1102 (N_1102,In_1365,In_1618);
or U1103 (N_1103,In_905,N_735);
xnor U1104 (N_1104,N_807,N_922);
nor U1105 (N_1105,N_625,N_444);
xnor U1106 (N_1106,N_657,N_353);
nand U1107 (N_1107,In_1634,In_1756);
nor U1108 (N_1108,In_915,N_223);
nand U1109 (N_1109,N_848,N_867);
nor U1110 (N_1110,N_619,In_1434);
nand U1111 (N_1111,In_801,In_526);
or U1112 (N_1112,N_630,N_514);
or U1113 (N_1113,In_1556,N_464);
or U1114 (N_1114,In_712,N_575);
xnor U1115 (N_1115,N_212,N_753);
nand U1116 (N_1116,In_888,N_14);
nor U1117 (N_1117,N_952,In_892);
and U1118 (N_1118,N_765,N_125);
and U1119 (N_1119,N_833,In_996);
and U1120 (N_1120,In_1413,In_882);
or U1121 (N_1121,N_902,N_1045);
xor U1122 (N_1122,In_1456,N_288);
xnor U1123 (N_1123,N_375,N_459);
and U1124 (N_1124,N_239,N_1052);
nand U1125 (N_1125,N_904,In_651);
and U1126 (N_1126,N_831,N_1034);
or U1127 (N_1127,N_155,In_538);
xor U1128 (N_1128,In_1604,N_385);
and U1129 (N_1129,In_1792,In_1319);
xnor U1130 (N_1130,N_733,N_694);
nand U1131 (N_1131,N_966,In_6);
nor U1132 (N_1132,N_1005,N_1016);
nand U1133 (N_1133,N_814,In_1492);
nor U1134 (N_1134,In_1850,In_788);
and U1135 (N_1135,N_548,In_505);
xnor U1136 (N_1136,In_1992,In_1195);
nor U1137 (N_1137,N_232,N_522);
nor U1138 (N_1138,N_589,N_461);
nor U1139 (N_1139,N_860,In_192);
nor U1140 (N_1140,N_857,N_706);
nand U1141 (N_1141,N_918,N_323);
and U1142 (N_1142,N_311,In_282);
nor U1143 (N_1143,N_318,In_1536);
xor U1144 (N_1144,N_1107,N_948);
nand U1145 (N_1145,N_397,N_926);
nand U1146 (N_1146,N_558,N_842);
and U1147 (N_1147,In_1060,N_1035);
or U1148 (N_1148,In_1455,N_628);
nor U1149 (N_1149,N_454,In_828);
nand U1150 (N_1150,N_849,In_1719);
or U1151 (N_1151,N_1084,N_756);
and U1152 (N_1152,In_821,N_993);
and U1153 (N_1153,N_1055,In_823);
xor U1154 (N_1154,N_992,N_977);
or U1155 (N_1155,N_1073,N_660);
xor U1156 (N_1156,In_760,N_1097);
or U1157 (N_1157,In_734,N_972);
xor U1158 (N_1158,N_564,In_1192);
nand U1159 (N_1159,N_405,N_724);
or U1160 (N_1160,N_122,In_1553);
or U1161 (N_1161,N_91,In_971);
and U1162 (N_1162,In_1889,In_1954);
or U1163 (N_1163,In_552,N_710);
and U1164 (N_1164,N_897,N_1048);
xor U1165 (N_1165,N_723,N_1027);
nor U1166 (N_1166,N_1026,N_500);
nand U1167 (N_1167,N_1032,N_830);
xor U1168 (N_1168,N_507,In_186);
nand U1169 (N_1169,N_903,N_349);
nand U1170 (N_1170,N_939,N_271);
nor U1171 (N_1171,In_20,N_821);
xor U1172 (N_1172,N_889,N_395);
nand U1173 (N_1173,N_816,In_1268);
nand U1174 (N_1174,N_963,N_755);
nand U1175 (N_1175,N_431,In_310);
nor U1176 (N_1176,N_985,In_1760);
xnor U1177 (N_1177,In_311,In_966);
xor U1178 (N_1178,N_942,In_169);
nand U1179 (N_1179,N_1008,N_667);
and U1180 (N_1180,In_881,In_1923);
or U1181 (N_1181,N_839,N_847);
xor U1182 (N_1182,N_802,N_1115);
or U1183 (N_1183,N_615,N_601);
and U1184 (N_1184,In_403,In_78);
or U1185 (N_1185,In_1165,N_964);
nand U1186 (N_1186,N_851,In_722);
nor U1187 (N_1187,N_410,N_204);
nor U1188 (N_1188,N_784,N_425);
nor U1189 (N_1189,N_361,N_96);
nor U1190 (N_1190,In_831,N_1100);
or U1191 (N_1191,In_523,N_345);
xnor U1192 (N_1192,In_487,N_975);
xnor U1193 (N_1193,In_1217,N_462);
and U1194 (N_1194,In_830,In_1270);
nand U1195 (N_1195,In_1540,N_707);
nor U1196 (N_1196,N_878,N_465);
nor U1197 (N_1197,N_967,N_1085);
and U1198 (N_1198,In_1512,N_674);
and U1199 (N_1199,In_516,In_1650);
and U1200 (N_1200,In_919,N_604);
nand U1201 (N_1201,N_711,N_990);
nor U1202 (N_1202,In_1787,N_576);
and U1203 (N_1203,N_414,N_1051);
nor U1204 (N_1204,In_386,In_1477);
xnor U1205 (N_1205,In_363,In_635);
nand U1206 (N_1206,N_559,In_1795);
xnor U1207 (N_1207,N_1063,N_128);
and U1208 (N_1208,N_1012,N_561);
or U1209 (N_1209,N_214,In_978);
nand U1210 (N_1210,N_725,N_66);
nor U1211 (N_1211,In_139,N_521);
and U1212 (N_1212,In_987,N_1113);
xnor U1213 (N_1213,In_660,In_1446);
and U1214 (N_1214,In_616,In_1142);
nand U1215 (N_1215,N_969,N_636);
and U1216 (N_1216,N_631,N_1119);
nand U1217 (N_1217,In_639,In_1735);
nand U1218 (N_1218,In_708,N_1007);
xor U1219 (N_1219,N_1040,N_529);
or U1220 (N_1220,In_917,N_1103);
nand U1221 (N_1221,In_1438,In_1212);
or U1222 (N_1222,N_334,N_978);
nand U1223 (N_1223,In_218,N_1047);
nor U1224 (N_1224,In_37,N_313);
nand U1225 (N_1225,N_350,N_443);
or U1226 (N_1226,N_734,In_268);
xnor U1227 (N_1227,In_323,N_545);
and U1228 (N_1228,In_415,N_941);
and U1229 (N_1229,N_720,In_1608);
or U1230 (N_1230,N_854,In_688);
or U1231 (N_1231,In_718,N_762);
and U1232 (N_1232,In_427,N_3);
nand U1233 (N_1233,In_1693,N_253);
or U1234 (N_1234,In_81,In_509);
and U1235 (N_1235,In_800,In_1418);
and U1236 (N_1236,N_1004,N_570);
and U1237 (N_1237,N_909,N_195);
nor U1238 (N_1238,N_981,N_402);
nand U1239 (N_1239,N_984,In_275);
and U1240 (N_1240,In_578,In_1356);
nor U1241 (N_1241,In_537,N_654);
or U1242 (N_1242,N_721,N_378);
nor U1243 (N_1243,In_319,N_372);
or U1244 (N_1244,N_915,N_1019);
or U1245 (N_1245,N_1087,N_533);
nor U1246 (N_1246,N_141,In_1571);
and U1247 (N_1247,In_1175,N_68);
nor U1248 (N_1248,N_690,In_750);
xnor U1249 (N_1249,In_1412,In_177);
nor U1250 (N_1250,In_1680,In_16);
and U1251 (N_1251,N_247,N_493);
and U1252 (N_1252,N_1071,In_1458);
nand U1253 (N_1253,In_102,N_1021);
nor U1254 (N_1254,N_741,In_267);
xnor U1255 (N_1255,N_594,N_553);
nor U1256 (N_1256,In_767,N_961);
nand U1257 (N_1257,N_189,N_986);
or U1258 (N_1258,In_1726,In_1524);
or U1259 (N_1259,N_566,N_84);
and U1260 (N_1260,N_1108,In_392);
nand U1261 (N_1261,N_1039,In_754);
or U1262 (N_1262,N_592,N_1078);
nor U1263 (N_1263,In_1156,N_436);
and U1264 (N_1264,N_865,N_910);
and U1265 (N_1265,N_804,N_1077);
or U1266 (N_1266,N_761,N_717);
nor U1267 (N_1267,N_320,N_718);
xnor U1268 (N_1268,In_1141,N_555);
or U1269 (N_1269,N_341,In_23);
nor U1270 (N_1270,N_1054,In_645);
or U1271 (N_1271,N_793,In_1732);
xor U1272 (N_1272,In_318,In_954);
or U1273 (N_1273,In_80,N_117);
nor U1274 (N_1274,In_1653,N_980);
nand U1275 (N_1275,N_1003,N_326);
xor U1276 (N_1276,N_792,In_667);
and U1277 (N_1277,N_1075,N_965);
xor U1278 (N_1278,N_596,N_907);
nor U1279 (N_1279,In_797,In_1331);
nor U1280 (N_1280,In_1139,In_451);
xnor U1281 (N_1281,In_545,In_1533);
xor U1282 (N_1282,N_1225,N_1155);
nor U1283 (N_1283,In_379,N_1175);
and U1284 (N_1284,N_193,In_216);
or U1285 (N_1285,N_83,N_181);
nor U1286 (N_1286,N_1207,N_1150);
xor U1287 (N_1287,N_1167,N_888);
or U1288 (N_1288,In_664,N_1177);
nor U1289 (N_1289,In_411,N_983);
xnor U1290 (N_1290,N_1230,N_1157);
or U1291 (N_1291,N_488,N_834);
or U1292 (N_1292,N_671,In_206);
nand U1293 (N_1293,N_1056,In_373);
or U1294 (N_1294,N_766,In_887);
xnor U1295 (N_1295,N_1038,N_496);
nor U1296 (N_1296,N_542,N_1123);
or U1297 (N_1297,N_1235,In_1896);
nor U1298 (N_1298,N_1000,N_509);
nand U1299 (N_1299,N_1153,N_1148);
xnor U1300 (N_1300,In_1020,N_1272);
xor U1301 (N_1301,N_1080,In_1363);
xnor U1302 (N_1302,N_872,In_67);
or U1303 (N_1303,N_982,N_1116);
and U1304 (N_1304,N_845,N_787);
nor U1305 (N_1305,N_684,N_623);
xnor U1306 (N_1306,In_15,N_1241);
nor U1307 (N_1307,N_813,N_989);
nand U1308 (N_1308,In_574,In_320);
nor U1309 (N_1309,In_1140,N_869);
and U1310 (N_1310,N_123,N_1223);
nor U1311 (N_1311,N_855,N_1105);
nor U1312 (N_1312,N_258,N_1042);
nor U1313 (N_1313,N_940,In_1705);
xor U1314 (N_1314,In_1699,N_1268);
or U1315 (N_1315,In_524,N_954);
or U1316 (N_1316,N_771,N_877);
xor U1317 (N_1317,N_435,N_973);
or U1318 (N_1318,In_778,N_549);
and U1319 (N_1319,N_367,In_458);
or U1320 (N_1320,N_1099,N_899);
and U1321 (N_1321,N_1205,N_944);
and U1322 (N_1322,In_1210,In_1364);
xor U1323 (N_1323,In_898,N_294);
nand U1324 (N_1324,N_1227,N_182);
nand U1325 (N_1325,N_796,In_125);
and U1326 (N_1326,N_960,N_1015);
xor U1327 (N_1327,In_1912,N_863);
and U1328 (N_1328,N_822,N_321);
or U1329 (N_1329,N_1209,N_539);
nor U1330 (N_1330,In_235,N_837);
or U1331 (N_1331,In_91,N_875);
nor U1332 (N_1332,N_1191,N_1222);
or U1333 (N_1333,In_1362,N_1023);
or U1334 (N_1334,In_1762,N_1245);
xnor U1335 (N_1335,N_587,N_46);
xor U1336 (N_1336,N_1137,N_1104);
nand U1337 (N_1337,In_47,N_1059);
and U1338 (N_1338,In_1914,In_116);
nand U1339 (N_1339,N_1164,N_1278);
nand U1340 (N_1340,N_682,N_58);
nor U1341 (N_1341,N_331,N_1127);
nor U1342 (N_1342,In_1686,N_658);
xnor U1343 (N_1343,In_1633,N_1037);
nand U1344 (N_1344,N_1183,N_782);
nand U1345 (N_1345,In_14,In_44);
xnor U1346 (N_1346,N_956,In_1221);
xnor U1347 (N_1347,In_624,N_634);
or U1348 (N_1348,N_678,N_773);
xnor U1349 (N_1349,N_1089,N_169);
nor U1350 (N_1350,In_1768,N_1204);
and U1351 (N_1351,In_188,N_1142);
nand U1352 (N_1352,N_1173,N_1258);
or U1353 (N_1353,N_1273,N_1066);
xor U1354 (N_1354,N_746,N_894);
or U1355 (N_1355,N_704,N_1264);
xor U1356 (N_1356,N_1244,N_1109);
xnor U1357 (N_1357,N_359,N_207);
and U1358 (N_1358,N_1259,N_722);
xor U1359 (N_1359,N_1254,In_1394);
or U1360 (N_1360,In_348,N_409);
nor U1361 (N_1361,N_1053,N_1208);
and U1362 (N_1362,N_210,N_1251);
or U1363 (N_1363,N_482,N_656);
or U1364 (N_1364,N_471,In_1819);
xnor U1365 (N_1365,In_870,N_974);
xnor U1366 (N_1366,N_1275,N_1174);
nor U1367 (N_1367,In_1767,N_911);
and U1368 (N_1368,N_998,In_1125);
and U1369 (N_1369,N_995,N_1199);
nor U1370 (N_1370,In_609,N_1001);
or U1371 (N_1371,N_1010,N_675);
and U1372 (N_1372,N_844,In_953);
nand U1373 (N_1373,N_1248,N_1118);
or U1374 (N_1374,N_759,N_1134);
xor U1375 (N_1375,N_25,N_1247);
and U1376 (N_1376,In_327,N_1172);
nand U1377 (N_1377,N_515,N_1036);
or U1378 (N_1378,N_1096,N_1187);
nand U1379 (N_1379,N_1091,In_126);
nand U1380 (N_1380,In_528,In_735);
and U1381 (N_1381,N_827,N_890);
xor U1382 (N_1382,N_1044,N_614);
and U1383 (N_1383,N_1147,In_1373);
nor U1384 (N_1384,N_1124,N_1166);
or U1385 (N_1385,N_399,N_856);
or U1386 (N_1386,In_1542,In_204);
or U1387 (N_1387,N_1031,N_1255);
nand U1388 (N_1388,N_951,In_998);
and U1389 (N_1389,N_360,N_1271);
nand U1390 (N_1390,N_0,N_595);
or U1391 (N_1391,N_937,In_1348);
nor U1392 (N_1392,N_1214,In_1631);
and U1393 (N_1393,N_1156,N_641);
or U1394 (N_1394,In_1982,N_196);
xor U1395 (N_1395,N_198,N_277);
nand U1396 (N_1396,N_823,N_705);
or U1397 (N_1397,N_1122,N_1072);
xor U1398 (N_1398,In_19,N_825);
and U1399 (N_1399,N_1160,N_1049);
and U1400 (N_1400,N_923,In_1609);
nor U1401 (N_1401,In_1276,In_1555);
nor U1402 (N_1402,N_130,N_1117);
and U1403 (N_1403,N_861,N_1262);
xor U1404 (N_1404,In_854,N_283);
nor U1405 (N_1405,In_1386,In_69);
nor U1406 (N_1406,N_1274,N_451);
nand U1407 (N_1407,N_880,N_1050);
and U1408 (N_1408,In_1117,N_702);
and U1409 (N_1409,N_175,In_525);
or U1410 (N_1410,N_1233,In_1298);
nor U1411 (N_1411,N_1246,In_1983);
nand U1412 (N_1412,In_1021,In_981);
or U1413 (N_1413,N_1263,N_1133);
xnor U1414 (N_1414,N_1185,N_1238);
nand U1415 (N_1415,N_962,N_1136);
and U1416 (N_1416,N_742,In_9);
nor U1417 (N_1417,N_1058,N_183);
and U1418 (N_1418,N_1193,N_1163);
xor U1419 (N_1419,N_138,N_177);
and U1420 (N_1420,N_627,N_560);
xor U1421 (N_1421,N_791,N_649);
nand U1422 (N_1422,N_1090,N_1110);
nor U1423 (N_1423,N_1236,N_267);
or U1424 (N_1424,N_632,In_1046);
xnor U1425 (N_1425,N_1211,N_1260);
and U1426 (N_1426,N_290,N_928);
and U1427 (N_1427,In_26,N_931);
xnor U1428 (N_1428,N_1220,N_1143);
or U1429 (N_1429,N_728,In_1852);
xor U1430 (N_1430,N_1261,N_991);
nor U1431 (N_1431,N_729,In_1805);
nor U1432 (N_1432,N_1242,In_1371);
nand U1433 (N_1433,N_1279,N_1154);
nor U1434 (N_1434,N_893,N_943);
xnor U1435 (N_1435,In_1274,N_906);
nor U1436 (N_1436,In_1677,N_129);
and U1437 (N_1437,N_1234,N_987);
nand U1438 (N_1438,In_484,N_1121);
and U1439 (N_1439,N_1192,N_234);
nand U1440 (N_1440,In_1965,N_730);
xor U1441 (N_1441,In_1814,In_1078);
or U1442 (N_1442,N_1434,N_1416);
nor U1443 (N_1443,N_1002,N_790);
nand U1444 (N_1444,In_1866,N_1318);
and U1445 (N_1445,N_819,In_1099);
and U1446 (N_1446,N_1311,In_819);
nor U1447 (N_1447,In_810,In_220);
and U1448 (N_1448,N_1081,N_16);
xnor U1449 (N_1449,N_1302,N_1297);
nand U1450 (N_1450,N_996,N_1184);
nor U1451 (N_1451,In_1287,In_312);
xnor U1452 (N_1452,N_1145,N_54);
or U1453 (N_1453,N_1344,In_952);
nand U1454 (N_1454,N_1141,N_1006);
nand U1455 (N_1455,N_276,N_719);
xnor U1456 (N_1456,N_1327,In_360);
or U1457 (N_1457,N_1337,In_468);
nor U1458 (N_1458,N_42,N_1404);
or U1459 (N_1459,N_1387,N_51);
xnor U1460 (N_1460,N_1436,N_1384);
xnor U1461 (N_1461,N_1128,N_1428);
or U1462 (N_1462,N_1432,N_1379);
xnor U1463 (N_1463,N_778,In_1589);
nor U1464 (N_1464,N_1399,N_384);
nand U1465 (N_1465,In_1882,N_767);
nor U1466 (N_1466,N_602,N_1400);
or U1467 (N_1467,N_1202,N_1309);
nor U1468 (N_1468,In_653,N_1418);
and U1469 (N_1469,In_1848,N_1282);
nand U1470 (N_1470,N_1398,N_624);
and U1471 (N_1471,N_841,N_1347);
nand U1472 (N_1472,N_798,N_1028);
and U1473 (N_1473,N_1394,In_1844);
nand U1474 (N_1474,N_1158,N_1402);
nand U1475 (N_1475,N_805,N_1349);
or U1476 (N_1476,N_1383,In_86);
or U1477 (N_1477,N_1338,N_1120);
xor U1478 (N_1478,N_456,N_1290);
or U1479 (N_1479,N_1417,In_1601);
nor U1480 (N_1480,N_166,In_1518);
and U1481 (N_1481,N_1267,N_1299);
xor U1482 (N_1482,N_668,N_1293);
and U1483 (N_1483,In_1224,N_1395);
nor U1484 (N_1484,N_621,In_309);
nor U1485 (N_1485,N_1397,N_920);
and U1486 (N_1486,N_1088,In_322);
nand U1487 (N_1487,N_1335,N_1283);
xor U1488 (N_1488,N_1291,N_655);
nand U1489 (N_1489,N_73,N_879);
nor U1490 (N_1490,N_449,In_428);
nand U1491 (N_1491,N_511,In_1817);
nor U1492 (N_1492,In_772,In_1488);
xor U1493 (N_1493,N_1102,N_1188);
or U1494 (N_1494,In_914,N_1422);
nand U1495 (N_1495,N_433,In_1829);
or U1496 (N_1496,N_107,N_1385);
and U1497 (N_1497,N_1367,In_485);
nor U1498 (N_1498,N_1312,N_1256);
nor U1499 (N_1499,N_1353,N_137);
nor U1500 (N_1500,N_1083,In_94);
xnor U1501 (N_1501,N_1178,N_368);
or U1502 (N_1502,N_1323,N_1414);
nor U1503 (N_1503,In_442,N_1011);
xor U1504 (N_1504,N_938,N_1082);
xnor U1505 (N_1505,N_1070,N_1303);
nand U1506 (N_1506,N_1041,N_1423);
and U1507 (N_1507,N_1285,N_968);
nor U1508 (N_1508,N_788,In_861);
or U1509 (N_1509,In_89,N_1030);
xor U1510 (N_1510,N_1328,N_852);
nand U1511 (N_1511,In_1043,N_1182);
and U1512 (N_1512,N_1427,N_898);
nand U1513 (N_1513,N_577,N_530);
xnor U1514 (N_1514,N_1144,N_1405);
or U1515 (N_1515,N_157,N_490);
or U1516 (N_1516,N_908,N_588);
nand U1517 (N_1517,N_955,N_1190);
nor U1518 (N_1518,N_651,N_1201);
nor U1519 (N_1519,N_786,N_1424);
and U1520 (N_1520,N_1249,N_988);
or U1521 (N_1521,N_273,N_1179);
and U1522 (N_1522,N_1094,N_1316);
or U1523 (N_1523,In_569,In_853);
nand U1524 (N_1524,N_1151,N_1198);
nor U1525 (N_1525,N_72,In_567);
nand U1526 (N_1526,N_1341,In_838);
xor U1527 (N_1527,N_1329,N_1065);
nor U1528 (N_1528,N_419,N_1289);
nand U1529 (N_1529,N_1357,N_835);
nor U1530 (N_1530,N_1130,In_1926);
or U1531 (N_1531,N_1033,N_1135);
and U1532 (N_1532,In_163,In_1454);
or U1533 (N_1533,N_692,N_1284);
and U1534 (N_1534,N_1350,In_736);
nor U1535 (N_1535,N_1364,N_165);
nor U1536 (N_1536,N_1281,N_1315);
and U1537 (N_1537,N_1186,N_739);
or U1538 (N_1538,N_716,N_316);
or U1539 (N_1539,N_1197,N_1401);
and U1540 (N_1540,N_697,N_1406);
and U1541 (N_1541,In_1059,N_1368);
or U1542 (N_1542,N_957,In_1050);
nand U1543 (N_1543,N_698,N_1296);
or U1544 (N_1544,N_1354,N_994);
and U1545 (N_1545,N_1221,N_1363);
or U1546 (N_1546,N_736,N_1439);
and U1547 (N_1547,N_1306,N_1294);
or U1548 (N_1548,N_1333,N_1420);
nor U1549 (N_1549,In_1219,N_1206);
xnor U1550 (N_1550,N_1232,N_1068);
nor U1551 (N_1551,N_512,N_281);
nor U1552 (N_1552,In_10,N_971);
xor U1553 (N_1553,N_1345,N_997);
nor U1554 (N_1554,N_1093,In_1133);
xnor U1555 (N_1555,N_864,N_912);
nor U1556 (N_1556,N_1213,N_1159);
or U1557 (N_1557,N_75,In_1949);
and U1558 (N_1558,N_1126,N_1196);
nand U1559 (N_1559,In_1294,N_1228);
nand U1560 (N_1560,N_1092,N_713);
or U1561 (N_1561,In_812,N_1376);
nor U1562 (N_1562,N_1381,N_748);
or U1563 (N_1563,N_862,N_1310);
nor U1564 (N_1564,In_148,N_1325);
xnor U1565 (N_1565,N_1307,N_1057);
nand U1566 (N_1566,N_306,N_1252);
or U1567 (N_1567,In_490,N_408);
or U1568 (N_1568,N_1438,N_1419);
nand U1569 (N_1569,N_801,N_900);
xnor U1570 (N_1570,N_745,In_1718);
and U1571 (N_1571,N_1426,N_1380);
nor U1572 (N_1572,N_457,N_209);
nor U1573 (N_1573,In_84,In_262);
xnor U1574 (N_1574,N_1301,N_1305);
nor U1575 (N_1575,N_468,In_555);
xor U1576 (N_1576,In_1944,N_1343);
nand U1577 (N_1577,N_1025,N_1351);
xnor U1578 (N_1578,N_1146,N_1111);
nand U1579 (N_1579,N_1162,N_715);
or U1580 (N_1580,In_209,N_478);
xor U1581 (N_1581,N_1339,N_1022);
nor U1582 (N_1582,N_1095,N_240);
nor U1583 (N_1583,N_700,N_492);
or U1584 (N_1584,N_672,In_1890);
nor U1585 (N_1585,N_1062,N_929);
nor U1586 (N_1586,N_1013,In_1055);
nor U1587 (N_1587,N_1269,N_1374);
or U1588 (N_1588,N_1431,In_1159);
xor U1589 (N_1589,N_933,N_1226);
nand U1590 (N_1590,In_1655,N_757);
nand U1591 (N_1591,N_1332,In_1313);
nor U1592 (N_1592,N_1168,N_1243);
or U1593 (N_1593,N_1369,N_1409);
nand U1594 (N_1594,N_1352,N_714);
nand U1595 (N_1595,N_1389,N_1217);
and U1596 (N_1596,N_1415,N_1300);
nand U1597 (N_1597,N_1288,N_1029);
xnor U1598 (N_1598,N_1020,N_749);
nand U1599 (N_1599,In_752,N_1009);
and U1600 (N_1600,N_1580,N_1590);
nand U1601 (N_1601,N_1407,N_1362);
xnor U1602 (N_1602,N_337,N_1342);
nor U1603 (N_1603,In_1761,N_1043);
nor U1604 (N_1604,N_1076,In_1100);
or U1605 (N_1605,N_1533,In_961);
xor U1606 (N_1606,In_1920,N_1579);
and U1607 (N_1607,N_328,N_1064);
and U1608 (N_1608,N_1466,N_1535);
or U1609 (N_1609,N_1578,N_760);
nor U1610 (N_1610,N_1319,N_1443);
and U1611 (N_1611,N_1355,N_1346);
xor U1612 (N_1612,N_1435,In_680);
nand U1613 (N_1613,N_1536,N_1139);
xor U1614 (N_1614,In_1280,N_1203);
nor U1615 (N_1615,N_1483,N_1014);
and U1616 (N_1616,N_1046,N_1456);
xor U1617 (N_1617,N_1497,N_1250);
nor U1618 (N_1618,N_1474,N_1480);
or U1619 (N_1619,N_160,N_1531);
xnor U1620 (N_1620,N_1371,In_457);
nor U1621 (N_1621,N_1373,N_1421);
or U1622 (N_1622,N_1138,In_1027);
and U1623 (N_1623,In_975,N_1561);
or U1624 (N_1624,N_1152,N_1140);
nor U1625 (N_1625,N_1500,N_1571);
and U1626 (N_1626,N_1595,In_610);
or U1627 (N_1627,In_1238,N_1448);
and U1628 (N_1628,N_1069,N_585);
and U1629 (N_1629,N_1461,N_1547);
xnor U1630 (N_1630,N_1149,N_1464);
or U1631 (N_1631,In_1970,N_1444);
nor U1632 (N_1632,N_1523,N_1529);
xnor U1633 (N_1633,N_1575,N_1455);
or U1634 (N_1634,N_1598,N_1537);
xor U1635 (N_1635,N_1482,N_1573);
xnor U1636 (N_1636,In_916,N_882);
nor U1637 (N_1637,N_818,N_809);
nand U1638 (N_1638,N_1170,N_1181);
xor U1639 (N_1639,N_1180,N_1132);
nand U1640 (N_1640,N_1487,N_1548);
and U1641 (N_1641,N_1592,N_1358);
xor U1642 (N_1642,N_1060,N_403);
and U1643 (N_1643,N_1189,In_448);
nand U1644 (N_1644,N_1452,N_1488);
or U1645 (N_1645,N_1229,In_872);
nand U1646 (N_1646,N_1563,N_1556);
nand U1647 (N_1647,N_1503,In_956);
xor U1648 (N_1648,In_1237,N_959);
and U1649 (N_1649,N_532,N_1441);
and U1650 (N_1650,N_1528,N_976);
nand U1651 (N_1651,N_1570,N_1507);
or U1652 (N_1652,N_1581,N_1599);
nand U1653 (N_1653,N_554,N_1509);
nor U1654 (N_1654,N_485,N_812);
nand U1655 (N_1655,In_627,N_483);
xnor U1656 (N_1656,N_1237,N_1200);
or U1657 (N_1657,N_1386,N_1462);
or U1658 (N_1658,N_1292,N_669);
nor U1659 (N_1659,N_1511,In_1350);
nand U1660 (N_1660,N_19,N_1378);
nor U1661 (N_1661,N_1433,N_1541);
xor U1662 (N_1662,N_886,N_1112);
or U1663 (N_1663,N_1304,In_1423);
and U1664 (N_1664,N_1587,N_1472);
nand U1665 (N_1665,N_1218,N_1565);
and U1666 (N_1666,N_1564,N_1554);
or U1667 (N_1667,N_1018,N_1265);
nor U1668 (N_1668,N_1594,N_1525);
xor U1669 (N_1669,N_1593,N_1557);
and U1670 (N_1670,N_1447,N_1451);
nand U1671 (N_1671,N_600,N_1390);
nand U1672 (N_1672,In_895,N_1489);
nand U1673 (N_1673,N_1521,N_1520);
and U1674 (N_1674,N_1257,N_1540);
nor U1675 (N_1675,N_1382,N_1485);
xor U1676 (N_1676,N_1210,N_1524);
nor U1677 (N_1677,N_703,N_1530);
or U1678 (N_1678,N_892,N_442);
nand U1679 (N_1679,N_1161,N_380);
nand U1680 (N_1680,In_849,N_1317);
xor U1681 (N_1681,N_946,N_1471);
nor U1682 (N_1682,N_1295,N_1024);
and U1683 (N_1683,N_1101,N_1457);
xor U1684 (N_1684,N_1320,In_883);
or U1685 (N_1685,N_1504,N_1321);
or U1686 (N_1686,N_663,N_494);
nand U1687 (N_1687,N_1277,N_1176);
nor U1688 (N_1688,N_1129,N_1216);
xor U1689 (N_1689,N_1550,N_1219);
nor U1690 (N_1690,N_1553,N_1516);
nor U1691 (N_1691,N_868,N_1560);
nand U1692 (N_1692,In_761,N_1494);
nand U1693 (N_1693,N_1195,N_1331);
nor U1694 (N_1694,N_1545,N_1576);
and U1695 (N_1695,N_1460,N_1440);
xor U1696 (N_1696,N_1079,In_166);
and U1697 (N_1697,N_891,N_795);
xnor U1698 (N_1698,N_1396,N_1391);
or U1699 (N_1699,N_1552,N_305);
xnor U1700 (N_1700,N_1393,N_540);
or U1701 (N_1701,N_1266,N_1502);
nor U1702 (N_1702,N_1106,N_1499);
xnor U1703 (N_1703,N_999,In_1290);
or U1704 (N_1704,N_905,N_233);
or U1705 (N_1705,N_876,N_1481);
nand U1706 (N_1706,N_1348,In_766);
nor U1707 (N_1707,N_1549,N_1286);
nand U1708 (N_1708,N_934,N_1392);
and U1709 (N_1709,In_827,N_1558);
xnor U1710 (N_1710,N_1470,N_1467);
nand U1711 (N_1711,In_985,N_1370);
nor U1712 (N_1712,N_1375,N_1298);
nor U1713 (N_1713,N_1577,N_1411);
or U1714 (N_1714,N_1459,N_1453);
nand U1715 (N_1715,N_1544,N_1388);
or U1716 (N_1716,In_1353,N_1479);
and U1717 (N_1717,N_1585,N_1253);
and U1718 (N_1718,N_1582,N_1539);
xnor U1719 (N_1719,N_1538,N_1486);
nor U1720 (N_1720,N_1495,N_1574);
nor U1721 (N_1721,N_1322,In_1679);
nand U1722 (N_1722,N_826,N_1568);
nand U1723 (N_1723,N_1169,N_1425);
nand U1724 (N_1724,N_1430,In_408);
and U1725 (N_1725,N_970,In_494);
or U1726 (N_1726,N_1463,N_1171);
nand U1727 (N_1727,N_1445,N_1506);
or U1728 (N_1728,N_1287,N_1410);
and U1729 (N_1729,N_1437,N_1098);
xnor U1730 (N_1730,N_272,N_932);
and U1731 (N_1731,In_1993,N_1403);
and U1732 (N_1732,N_1572,In_782);
xnor U1733 (N_1733,N_1498,N_1365);
nand U1734 (N_1734,N_1517,N_1519);
and U1735 (N_1735,N_1270,N_1336);
or U1736 (N_1736,N_1551,N_1583);
nand U1737 (N_1737,N_1449,N_1061);
and U1738 (N_1738,N_1477,N_1542);
or U1739 (N_1739,N_1591,N_1454);
nand U1740 (N_1740,N_1566,N_1491);
or U1741 (N_1741,In_439,N_1543);
nand U1742 (N_1742,N_1224,N_1165);
nand U1743 (N_1743,N_1326,N_584);
nor U1744 (N_1744,N_262,N_680);
xor U1745 (N_1745,N_606,N_1586);
and U1746 (N_1746,N_1324,In_1318);
or U1747 (N_1747,N_1114,N_1413);
or U1748 (N_1748,N_1505,N_1596);
and U1749 (N_1749,In_1776,In_871);
or U1750 (N_1750,N_1567,N_1584);
nand U1751 (N_1751,In_1820,N_1372);
nor U1752 (N_1752,N_1067,N_1588);
or U1753 (N_1753,N_1490,N_1513);
or U1754 (N_1754,N_979,In_727);
and U1755 (N_1755,N_1476,N_1515);
nand U1756 (N_1756,N_1493,In_1832);
and U1757 (N_1757,N_1330,N_1334);
and U1758 (N_1758,In_547,In_1730);
xnor U1759 (N_1759,N_1508,N_1308);
or U1760 (N_1760,N_1748,N_1686);
nor U1761 (N_1761,N_1412,N_1651);
nor U1762 (N_1762,N_1314,N_1719);
or U1763 (N_1763,N_1635,N_1740);
nand U1764 (N_1764,N_1693,N_1734);
nand U1765 (N_1765,N_1723,N_1600);
nand U1766 (N_1766,N_1612,N_1643);
or U1767 (N_1767,N_1610,N_1086);
nand U1768 (N_1768,N_1731,N_1692);
xnor U1769 (N_1769,N_1194,N_1510);
or U1770 (N_1770,N_1648,N_1361);
or U1771 (N_1771,N_1465,N_1625);
xor U1772 (N_1772,N_1700,N_1745);
and U1773 (N_1773,N_1702,N_1450);
and U1774 (N_1774,N_257,N_1722);
xor U1775 (N_1775,N_1360,N_1655);
or U1776 (N_1776,N_1688,N_1646);
and U1777 (N_1777,N_1678,N_1366);
and U1778 (N_1778,N_1514,N_1750);
xor U1779 (N_1779,N_1630,N_1017);
xor U1780 (N_1780,N_1657,N_1615);
or U1781 (N_1781,N_1532,N_1616);
nand U1782 (N_1782,N_1589,N_1641);
or U1783 (N_1783,N_1468,N_1710);
nand U1784 (N_1784,N_1496,N_1623);
nor U1785 (N_1785,N_1602,N_1619);
nor U1786 (N_1786,N_1280,N_1650);
or U1787 (N_1787,N_1753,N_1708);
or U1788 (N_1788,N_1704,N_1313);
xnor U1789 (N_1789,In_1490,N_1597);
or U1790 (N_1790,N_1694,N_1746);
nor U1791 (N_1791,N_1721,N_1622);
nor U1792 (N_1792,N_1669,N_1276);
or U1793 (N_1793,N_1626,N_1484);
or U1794 (N_1794,N_1658,N_811);
xor U1795 (N_1795,N_1640,N_1526);
xnor U1796 (N_1796,N_1614,In_1340);
or U1797 (N_1797,N_1726,N_1606);
or U1798 (N_1798,N_1697,N_1707);
or U1799 (N_1799,N_1733,N_1356);
nor U1800 (N_1800,In_55,N_1527);
xnor U1801 (N_1801,N_1555,N_1215);
nor U1802 (N_1802,N_1603,N_1667);
nor U1803 (N_1803,N_1751,N_1212);
xnor U1804 (N_1804,N_1627,N_1756);
nand U1805 (N_1805,N_1676,In_1044);
xor U1806 (N_1806,N_1716,N_1687);
nand U1807 (N_1807,N_1239,N_1749);
xnor U1808 (N_1808,N_1624,N_1605);
and U1809 (N_1809,N_1649,N_1681);
nand U1810 (N_1810,N_1609,In_758);
and U1811 (N_1811,N_1546,N_927);
and U1812 (N_1812,N_1644,N_1668);
and U1813 (N_1813,N_1473,N_1730);
or U1814 (N_1814,N_1738,N_949);
nand U1815 (N_1815,N_1632,N_1377);
and U1816 (N_1816,N_1559,N_1458);
or U1817 (N_1817,N_495,N_1663);
xnor U1818 (N_1818,N_1645,N_1629);
or U1819 (N_1819,N_1660,N_1755);
xnor U1820 (N_1820,N_1522,N_1712);
nor U1821 (N_1821,N_1628,N_1492);
nand U1822 (N_1822,N_1672,N_1621);
or U1823 (N_1823,N_1665,N_1429);
nor U1824 (N_1824,N_139,N_1469);
xor U1825 (N_1825,N_1703,N_1240);
nor U1826 (N_1826,N_1727,N_1656);
nor U1827 (N_1827,N_1636,N_1653);
nor U1828 (N_1828,N_1713,N_1720);
nor U1829 (N_1829,N_1618,N_1739);
xnor U1830 (N_1830,N_1518,N_1705);
nand U1831 (N_1831,N_1680,N_1670);
or U1832 (N_1832,N_1691,N_1478);
or U1833 (N_1833,N_1729,N_1743);
or U1834 (N_1834,N_1642,N_1696);
and U1835 (N_1835,N_1340,N_1074);
xor U1836 (N_1836,N_1718,N_1675);
xor U1837 (N_1837,N_1701,N_1359);
xor U1838 (N_1838,N_1638,N_1634);
nand U1839 (N_1839,In_804,In_995);
or U1840 (N_1840,N_1654,N_1717);
nor U1841 (N_1841,N_1752,N_505);
xnor U1842 (N_1842,N_1666,N_1671);
nor U1843 (N_1843,N_1534,N_1620);
nand U1844 (N_1844,N_1408,N_1742);
and U1845 (N_1845,N_1617,In_613);
and U1846 (N_1846,N_1744,N_1683);
xor U1847 (N_1847,N_1512,N_1689);
nor U1848 (N_1848,In_1654,N_1673);
xnor U1849 (N_1849,N_1735,N_1659);
xnor U1850 (N_1850,N_1711,N_1699);
xnor U1851 (N_1851,N_1737,N_1633);
and U1852 (N_1852,In_168,N_1637);
or U1853 (N_1853,N_1601,N_1732);
and U1854 (N_1854,N_1709,N_1714);
nor U1855 (N_1855,N_1715,In_106);
xor U1856 (N_1856,N_1662,N_1682);
nand U1857 (N_1857,N_1747,N_1759);
nand U1858 (N_1858,N_1639,N_1664);
nor U1859 (N_1859,In_1774,N_1631);
xor U1860 (N_1860,In_1427,N_1724);
or U1861 (N_1861,N_1695,N_935);
nor U1862 (N_1862,N_1706,N_1725);
and U1863 (N_1863,N_1684,N_1569);
xnor U1864 (N_1864,N_432,N_1736);
xor U1865 (N_1865,N_1125,N_1679);
nor U1866 (N_1866,N_836,N_1442);
nor U1867 (N_1867,N_1741,N_1652);
nor U1868 (N_1868,N_1131,N_1613);
or U1869 (N_1869,N_1611,N_1677);
or U1870 (N_1870,N_1475,N_1754);
or U1871 (N_1871,N_1501,In_740);
xor U1872 (N_1872,N_874,N_1685);
and U1873 (N_1873,N_1562,N_1661);
xnor U1874 (N_1874,N_1757,N_1446);
or U1875 (N_1875,N_1231,N_1647);
nor U1876 (N_1876,N_1607,N_1608);
nand U1877 (N_1877,N_1758,N_1698);
xor U1878 (N_1878,N_1728,N_1604);
and U1879 (N_1879,N_1674,N_1690);
and U1880 (N_1880,N_1473,N_1683);
and U1881 (N_1881,N_1684,N_1465);
nor U1882 (N_1882,N_1718,N_1644);
and U1883 (N_1883,N_1733,N_1632);
xor U1884 (N_1884,N_1617,N_1627);
or U1885 (N_1885,N_1602,N_1678);
or U1886 (N_1886,N_1745,N_1712);
nand U1887 (N_1887,N_1478,N_1231);
nand U1888 (N_1888,N_1662,N_1736);
and U1889 (N_1889,N_1510,N_1643);
nor U1890 (N_1890,N_1625,N_1703);
or U1891 (N_1891,N_1680,N_1737);
xor U1892 (N_1892,N_1473,N_1408);
or U1893 (N_1893,In_1774,N_1473);
nor U1894 (N_1894,In_1044,N_1478);
and U1895 (N_1895,N_1716,N_1736);
nand U1896 (N_1896,N_1534,N_874);
or U1897 (N_1897,N_1657,N_1646);
or U1898 (N_1898,N_1617,N_1670);
and U1899 (N_1899,N_1730,N_1615);
xor U1900 (N_1900,N_1484,N_1680);
and U1901 (N_1901,N_1635,N_1622);
nand U1902 (N_1902,N_1654,N_1314);
and U1903 (N_1903,N_1429,N_1759);
nor U1904 (N_1904,N_1740,N_1559);
and U1905 (N_1905,In_758,N_1648);
nor U1906 (N_1906,N_1704,In_55);
nor U1907 (N_1907,N_1715,N_1661);
nor U1908 (N_1908,N_1643,N_1650);
or U1909 (N_1909,N_1671,N_1732);
xnor U1910 (N_1910,N_1653,N_495);
nor U1911 (N_1911,N_1758,N_1613);
or U1912 (N_1912,N_1715,N_1601);
nor U1913 (N_1913,N_1657,N_1656);
xor U1914 (N_1914,N_1699,N_935);
and U1915 (N_1915,In_55,N_1276);
nor U1916 (N_1916,N_1608,N_1522);
and U1917 (N_1917,N_1620,N_1722);
nand U1918 (N_1918,N_1679,N_1707);
nor U1919 (N_1919,N_1724,N_1694);
xnor U1920 (N_1920,N_1874,N_1804);
nand U1921 (N_1921,N_1823,N_1770);
nor U1922 (N_1922,N_1894,N_1881);
and U1923 (N_1923,N_1807,N_1787);
and U1924 (N_1924,N_1789,N_1815);
nand U1925 (N_1925,N_1887,N_1898);
nor U1926 (N_1926,N_1909,N_1828);
nor U1927 (N_1927,N_1792,N_1783);
or U1928 (N_1928,N_1885,N_1912);
xnor U1929 (N_1929,N_1879,N_1833);
xnor U1930 (N_1930,N_1900,N_1777);
and U1931 (N_1931,N_1919,N_1808);
and U1932 (N_1932,N_1869,N_1877);
and U1933 (N_1933,N_1915,N_1764);
and U1934 (N_1934,N_1848,N_1886);
nor U1935 (N_1935,N_1847,N_1871);
nand U1936 (N_1936,N_1901,N_1802);
or U1937 (N_1937,N_1861,N_1809);
xor U1938 (N_1938,N_1910,N_1889);
nand U1939 (N_1939,N_1788,N_1902);
or U1940 (N_1940,N_1816,N_1820);
or U1941 (N_1941,N_1904,N_1813);
and U1942 (N_1942,N_1868,N_1858);
xor U1943 (N_1943,N_1841,N_1795);
and U1944 (N_1944,N_1782,N_1866);
xnor U1945 (N_1945,N_1878,N_1914);
nand U1946 (N_1946,N_1870,N_1846);
and U1947 (N_1947,N_1767,N_1806);
nand U1948 (N_1948,N_1850,N_1883);
xor U1949 (N_1949,N_1851,N_1880);
and U1950 (N_1950,N_1763,N_1906);
nand U1951 (N_1951,N_1760,N_1768);
and U1952 (N_1952,N_1891,N_1862);
nor U1953 (N_1953,N_1864,N_1786);
and U1954 (N_1954,N_1882,N_1840);
and U1955 (N_1955,N_1839,N_1772);
or U1956 (N_1956,N_1829,N_1849);
nand U1957 (N_1957,N_1825,N_1892);
xnor U1958 (N_1958,N_1824,N_1908);
nand U1959 (N_1959,N_1852,N_1875);
xnor U1960 (N_1960,N_1793,N_1794);
or U1961 (N_1961,N_1855,N_1844);
nor U1962 (N_1962,N_1798,N_1890);
xor U1963 (N_1963,N_1822,N_1790);
nor U1964 (N_1964,N_1873,N_1800);
and U1965 (N_1965,N_1854,N_1907);
xor U1966 (N_1966,N_1805,N_1888);
nor U1967 (N_1967,N_1860,N_1836);
nand U1968 (N_1968,N_1819,N_1784);
xnor U1969 (N_1969,N_1838,N_1776);
xnor U1970 (N_1970,N_1779,N_1876);
and U1971 (N_1971,N_1916,N_1801);
nor U1972 (N_1972,N_1778,N_1843);
and U1973 (N_1973,N_1766,N_1765);
or U1974 (N_1974,N_1799,N_1872);
nor U1975 (N_1975,N_1831,N_1837);
and U1976 (N_1976,N_1842,N_1785);
or U1977 (N_1977,N_1911,N_1811);
nand U1978 (N_1978,N_1780,N_1903);
nor U1979 (N_1979,N_1762,N_1796);
or U1980 (N_1980,N_1803,N_1863);
xnor U1981 (N_1981,N_1814,N_1865);
or U1982 (N_1982,N_1812,N_1884);
and U1983 (N_1983,N_1781,N_1818);
nor U1984 (N_1984,N_1774,N_1856);
or U1985 (N_1985,N_1769,N_1810);
nand U1986 (N_1986,N_1917,N_1857);
and U1987 (N_1987,N_1771,N_1834);
nor U1988 (N_1988,N_1821,N_1913);
xnor U1989 (N_1989,N_1895,N_1905);
or U1990 (N_1990,N_1845,N_1830);
and U1991 (N_1991,N_1918,N_1817);
nor U1992 (N_1992,N_1826,N_1797);
and U1993 (N_1993,N_1859,N_1827);
nand U1994 (N_1994,N_1773,N_1832);
or U1995 (N_1995,N_1897,N_1791);
and U1996 (N_1996,N_1896,N_1853);
xnor U1997 (N_1997,N_1761,N_1835);
or U1998 (N_1998,N_1899,N_1775);
xnor U1999 (N_1999,N_1893,N_1867);
and U2000 (N_2000,N_1914,N_1873);
and U2001 (N_2001,N_1778,N_1910);
or U2002 (N_2002,N_1888,N_1848);
xor U2003 (N_2003,N_1778,N_1819);
and U2004 (N_2004,N_1852,N_1794);
or U2005 (N_2005,N_1834,N_1817);
xnor U2006 (N_2006,N_1889,N_1821);
nand U2007 (N_2007,N_1850,N_1763);
xor U2008 (N_2008,N_1908,N_1776);
xnor U2009 (N_2009,N_1900,N_1878);
xor U2010 (N_2010,N_1787,N_1808);
xnor U2011 (N_2011,N_1863,N_1850);
nor U2012 (N_2012,N_1828,N_1760);
nor U2013 (N_2013,N_1796,N_1813);
or U2014 (N_2014,N_1800,N_1767);
nor U2015 (N_2015,N_1844,N_1875);
nand U2016 (N_2016,N_1772,N_1902);
or U2017 (N_2017,N_1869,N_1760);
nor U2018 (N_2018,N_1900,N_1826);
xor U2019 (N_2019,N_1812,N_1773);
xnor U2020 (N_2020,N_1822,N_1917);
xor U2021 (N_2021,N_1781,N_1841);
nand U2022 (N_2022,N_1767,N_1819);
xnor U2023 (N_2023,N_1908,N_1915);
or U2024 (N_2024,N_1795,N_1778);
xor U2025 (N_2025,N_1785,N_1820);
or U2026 (N_2026,N_1905,N_1775);
xnor U2027 (N_2027,N_1886,N_1794);
nand U2028 (N_2028,N_1869,N_1886);
xor U2029 (N_2029,N_1802,N_1800);
or U2030 (N_2030,N_1812,N_1804);
or U2031 (N_2031,N_1882,N_1857);
nor U2032 (N_2032,N_1894,N_1783);
and U2033 (N_2033,N_1859,N_1792);
and U2034 (N_2034,N_1834,N_1807);
and U2035 (N_2035,N_1910,N_1800);
nor U2036 (N_2036,N_1760,N_1885);
or U2037 (N_2037,N_1817,N_1895);
and U2038 (N_2038,N_1912,N_1873);
and U2039 (N_2039,N_1837,N_1792);
and U2040 (N_2040,N_1772,N_1862);
or U2041 (N_2041,N_1854,N_1911);
xnor U2042 (N_2042,N_1792,N_1829);
nand U2043 (N_2043,N_1823,N_1833);
xnor U2044 (N_2044,N_1791,N_1845);
and U2045 (N_2045,N_1800,N_1785);
nor U2046 (N_2046,N_1919,N_1910);
or U2047 (N_2047,N_1846,N_1813);
nand U2048 (N_2048,N_1843,N_1783);
and U2049 (N_2049,N_1891,N_1855);
and U2050 (N_2050,N_1911,N_1895);
nor U2051 (N_2051,N_1788,N_1914);
or U2052 (N_2052,N_1814,N_1886);
or U2053 (N_2053,N_1882,N_1893);
and U2054 (N_2054,N_1787,N_1847);
or U2055 (N_2055,N_1834,N_1769);
nand U2056 (N_2056,N_1914,N_1848);
or U2057 (N_2057,N_1907,N_1821);
and U2058 (N_2058,N_1806,N_1807);
xnor U2059 (N_2059,N_1832,N_1800);
xor U2060 (N_2060,N_1860,N_1767);
or U2061 (N_2061,N_1811,N_1804);
and U2062 (N_2062,N_1871,N_1807);
xor U2063 (N_2063,N_1799,N_1780);
and U2064 (N_2064,N_1826,N_1916);
nand U2065 (N_2065,N_1847,N_1777);
or U2066 (N_2066,N_1815,N_1778);
nor U2067 (N_2067,N_1906,N_1781);
and U2068 (N_2068,N_1792,N_1814);
or U2069 (N_2069,N_1806,N_1795);
and U2070 (N_2070,N_1792,N_1810);
xor U2071 (N_2071,N_1785,N_1770);
or U2072 (N_2072,N_1780,N_1918);
nor U2073 (N_2073,N_1846,N_1841);
xor U2074 (N_2074,N_1818,N_1801);
nor U2075 (N_2075,N_1848,N_1873);
nand U2076 (N_2076,N_1807,N_1912);
or U2077 (N_2077,N_1878,N_1917);
nand U2078 (N_2078,N_1899,N_1801);
xor U2079 (N_2079,N_1896,N_1881);
nand U2080 (N_2080,N_1945,N_1956);
xnor U2081 (N_2081,N_1968,N_1948);
xor U2082 (N_2082,N_1936,N_2044);
and U2083 (N_2083,N_1935,N_1987);
nand U2084 (N_2084,N_1960,N_2071);
nand U2085 (N_2085,N_1942,N_1924);
nand U2086 (N_2086,N_2028,N_1923);
xnor U2087 (N_2087,N_2007,N_1921);
nand U2088 (N_2088,N_2027,N_1978);
xor U2089 (N_2089,N_2038,N_2047);
or U2090 (N_2090,N_2043,N_1983);
nand U2091 (N_2091,N_2049,N_2032);
nand U2092 (N_2092,N_2021,N_2042);
nand U2093 (N_2093,N_1950,N_2054);
and U2094 (N_2094,N_1976,N_2008);
nor U2095 (N_2095,N_1937,N_2013);
nor U2096 (N_2096,N_1970,N_1999);
xnor U2097 (N_2097,N_2033,N_1995);
and U2098 (N_2098,N_2040,N_2072);
nand U2099 (N_2099,N_2031,N_2006);
nor U2100 (N_2100,N_1947,N_1979);
or U2101 (N_2101,N_1986,N_2046);
or U2102 (N_2102,N_1939,N_2037);
xnor U2103 (N_2103,N_1985,N_2005);
and U2104 (N_2104,N_2009,N_2024);
nand U2105 (N_2105,N_2056,N_2068);
nand U2106 (N_2106,N_1920,N_2012);
and U2107 (N_2107,N_1969,N_1959);
and U2108 (N_2108,N_1926,N_2077);
or U2109 (N_2109,N_2003,N_2051);
and U2110 (N_2110,N_1957,N_2075);
nand U2111 (N_2111,N_2030,N_1930);
and U2112 (N_2112,N_1952,N_1933);
or U2113 (N_2113,N_1994,N_2017);
and U2114 (N_2114,N_2069,N_1977);
xor U2115 (N_2115,N_2066,N_2070);
xnor U2116 (N_2116,N_1954,N_2023);
and U2117 (N_2117,N_2076,N_2015);
and U2118 (N_2118,N_1980,N_1934);
xnor U2119 (N_2119,N_1932,N_2018);
and U2120 (N_2120,N_1940,N_2052);
or U2121 (N_2121,N_2079,N_2064);
xor U2122 (N_2122,N_2026,N_1990);
or U2123 (N_2123,N_1955,N_2036);
xnor U2124 (N_2124,N_1925,N_2074);
or U2125 (N_2125,N_2061,N_2055);
nor U2126 (N_2126,N_1997,N_1966);
xnor U2127 (N_2127,N_2020,N_1949);
xor U2128 (N_2128,N_2019,N_1961);
nand U2129 (N_2129,N_1971,N_1962);
and U2130 (N_2130,N_2048,N_2004);
nand U2131 (N_2131,N_1993,N_1963);
and U2132 (N_2132,N_2029,N_1989);
or U2133 (N_2133,N_1975,N_2039);
nand U2134 (N_2134,N_1931,N_2010);
nand U2135 (N_2135,N_2022,N_2060);
xnor U2136 (N_2136,N_2065,N_2062);
and U2137 (N_2137,N_1973,N_2016);
or U2138 (N_2138,N_1964,N_1988);
nand U2139 (N_2139,N_2058,N_2057);
xor U2140 (N_2140,N_2041,N_2014);
nor U2141 (N_2141,N_1928,N_1922);
xnor U2142 (N_2142,N_1982,N_1998);
nor U2143 (N_2143,N_1929,N_2002);
nand U2144 (N_2144,N_2050,N_1941);
nand U2145 (N_2145,N_2001,N_2073);
or U2146 (N_2146,N_1992,N_1944);
xor U2147 (N_2147,N_1953,N_1951);
xnor U2148 (N_2148,N_2045,N_1974);
or U2149 (N_2149,N_2078,N_1991);
nand U2150 (N_2150,N_2034,N_1946);
or U2151 (N_2151,N_1965,N_1938);
nand U2152 (N_2152,N_2011,N_2063);
and U2153 (N_2153,N_1943,N_1967);
nor U2154 (N_2154,N_2025,N_1972);
xnor U2155 (N_2155,N_1958,N_2035);
or U2156 (N_2156,N_2059,N_1996);
xnor U2157 (N_2157,N_1981,N_2053);
or U2158 (N_2158,N_1927,N_2067);
nand U2159 (N_2159,N_1984,N_2000);
xor U2160 (N_2160,N_1980,N_2000);
nand U2161 (N_2161,N_2024,N_2067);
xnor U2162 (N_2162,N_2040,N_1980);
nand U2163 (N_2163,N_2014,N_1966);
nor U2164 (N_2164,N_1957,N_1926);
and U2165 (N_2165,N_1988,N_1927);
nand U2166 (N_2166,N_1968,N_2042);
nand U2167 (N_2167,N_1953,N_2031);
and U2168 (N_2168,N_2032,N_1935);
nor U2169 (N_2169,N_1970,N_2037);
xnor U2170 (N_2170,N_2047,N_1949);
and U2171 (N_2171,N_2039,N_2073);
and U2172 (N_2172,N_2040,N_1932);
or U2173 (N_2173,N_2077,N_2023);
or U2174 (N_2174,N_2041,N_1941);
xnor U2175 (N_2175,N_1978,N_1948);
xnor U2176 (N_2176,N_2025,N_2032);
nand U2177 (N_2177,N_2070,N_1980);
xnor U2178 (N_2178,N_2023,N_1997);
or U2179 (N_2179,N_2051,N_1934);
nor U2180 (N_2180,N_2051,N_1928);
and U2181 (N_2181,N_2007,N_1928);
nand U2182 (N_2182,N_1950,N_2006);
nand U2183 (N_2183,N_2062,N_2071);
xor U2184 (N_2184,N_2075,N_2049);
nand U2185 (N_2185,N_2063,N_2072);
or U2186 (N_2186,N_1963,N_1943);
nor U2187 (N_2187,N_2017,N_2012);
nor U2188 (N_2188,N_2045,N_1950);
and U2189 (N_2189,N_2009,N_1945);
xnor U2190 (N_2190,N_2064,N_2072);
and U2191 (N_2191,N_1995,N_1989);
nor U2192 (N_2192,N_2068,N_2026);
xnor U2193 (N_2193,N_2057,N_1950);
nor U2194 (N_2194,N_2068,N_2070);
xnor U2195 (N_2195,N_2065,N_2003);
nor U2196 (N_2196,N_2079,N_1952);
nor U2197 (N_2197,N_2016,N_2008);
xnor U2198 (N_2198,N_1948,N_1955);
nor U2199 (N_2199,N_2072,N_2050);
or U2200 (N_2200,N_2015,N_2004);
nand U2201 (N_2201,N_1958,N_1945);
nor U2202 (N_2202,N_2066,N_2009);
and U2203 (N_2203,N_1943,N_2074);
nand U2204 (N_2204,N_1973,N_2039);
or U2205 (N_2205,N_1938,N_1950);
and U2206 (N_2206,N_1945,N_2023);
xor U2207 (N_2207,N_1928,N_2064);
xnor U2208 (N_2208,N_1961,N_2003);
nand U2209 (N_2209,N_2033,N_2064);
and U2210 (N_2210,N_1936,N_2030);
nand U2211 (N_2211,N_1939,N_2005);
xnor U2212 (N_2212,N_1947,N_2027);
or U2213 (N_2213,N_2050,N_2052);
and U2214 (N_2214,N_1979,N_2072);
nor U2215 (N_2215,N_1973,N_2038);
nor U2216 (N_2216,N_2067,N_2049);
or U2217 (N_2217,N_1989,N_2067);
xnor U2218 (N_2218,N_1953,N_2063);
and U2219 (N_2219,N_2000,N_1990);
xor U2220 (N_2220,N_1986,N_1932);
or U2221 (N_2221,N_1968,N_1957);
nand U2222 (N_2222,N_2038,N_2042);
xor U2223 (N_2223,N_2002,N_1950);
nor U2224 (N_2224,N_1938,N_1975);
nor U2225 (N_2225,N_1987,N_1962);
and U2226 (N_2226,N_1960,N_2079);
nor U2227 (N_2227,N_2001,N_1995);
and U2228 (N_2228,N_2063,N_1940);
nor U2229 (N_2229,N_1949,N_1994);
xor U2230 (N_2230,N_2058,N_1967);
nor U2231 (N_2231,N_2015,N_1952);
xnor U2232 (N_2232,N_1982,N_2022);
nand U2233 (N_2233,N_1960,N_1942);
nor U2234 (N_2234,N_1929,N_2071);
or U2235 (N_2235,N_2076,N_1921);
and U2236 (N_2236,N_2011,N_1928);
and U2237 (N_2237,N_2071,N_1943);
nor U2238 (N_2238,N_2039,N_1993);
nor U2239 (N_2239,N_1925,N_2031);
or U2240 (N_2240,N_2165,N_2176);
nand U2241 (N_2241,N_2202,N_2148);
nor U2242 (N_2242,N_2187,N_2153);
nor U2243 (N_2243,N_2194,N_2114);
xnor U2244 (N_2244,N_2093,N_2096);
nand U2245 (N_2245,N_2110,N_2227);
nor U2246 (N_2246,N_2175,N_2112);
or U2247 (N_2247,N_2131,N_2235);
or U2248 (N_2248,N_2201,N_2119);
nand U2249 (N_2249,N_2220,N_2116);
nand U2250 (N_2250,N_2142,N_2206);
nor U2251 (N_2251,N_2212,N_2167);
nor U2252 (N_2252,N_2209,N_2132);
nor U2253 (N_2253,N_2180,N_2135);
or U2254 (N_2254,N_2103,N_2092);
or U2255 (N_2255,N_2216,N_2086);
or U2256 (N_2256,N_2098,N_2141);
or U2257 (N_2257,N_2203,N_2126);
nand U2258 (N_2258,N_2101,N_2123);
or U2259 (N_2259,N_2184,N_2236);
xnor U2260 (N_2260,N_2205,N_2106);
xor U2261 (N_2261,N_2087,N_2169);
xor U2262 (N_2262,N_2082,N_2197);
nor U2263 (N_2263,N_2160,N_2199);
and U2264 (N_2264,N_2178,N_2183);
and U2265 (N_2265,N_2228,N_2208);
nand U2266 (N_2266,N_2174,N_2102);
nand U2267 (N_2267,N_2164,N_2229);
nand U2268 (N_2268,N_2145,N_2193);
nand U2269 (N_2269,N_2127,N_2168);
xor U2270 (N_2270,N_2182,N_2237);
or U2271 (N_2271,N_2191,N_2083);
nor U2272 (N_2272,N_2214,N_2088);
and U2273 (N_2273,N_2188,N_2085);
and U2274 (N_2274,N_2166,N_2239);
xnor U2275 (N_2275,N_2151,N_2213);
or U2276 (N_2276,N_2080,N_2137);
xor U2277 (N_2277,N_2190,N_2172);
xor U2278 (N_2278,N_2221,N_2159);
nand U2279 (N_2279,N_2120,N_2136);
or U2280 (N_2280,N_2113,N_2143);
nor U2281 (N_2281,N_2100,N_2140);
or U2282 (N_2282,N_2224,N_2091);
xor U2283 (N_2283,N_2117,N_2161);
or U2284 (N_2284,N_2090,N_2222);
nand U2285 (N_2285,N_2121,N_2144);
or U2286 (N_2286,N_2130,N_2155);
nand U2287 (N_2287,N_2133,N_2134);
and U2288 (N_2288,N_2157,N_2238);
or U2289 (N_2289,N_2104,N_2118);
nor U2290 (N_2290,N_2192,N_2170);
nor U2291 (N_2291,N_2210,N_2207);
xor U2292 (N_2292,N_2163,N_2111);
nand U2293 (N_2293,N_2129,N_2125);
nand U2294 (N_2294,N_2179,N_2105);
and U2295 (N_2295,N_2099,N_2223);
xor U2296 (N_2296,N_2124,N_2226);
nand U2297 (N_2297,N_2158,N_2218);
nor U2298 (N_2298,N_2215,N_2162);
nor U2299 (N_2299,N_2107,N_2138);
and U2300 (N_2300,N_2156,N_2152);
nor U2301 (N_2301,N_2108,N_2186);
xnor U2302 (N_2302,N_2196,N_2233);
and U2303 (N_2303,N_2150,N_2225);
nand U2304 (N_2304,N_2139,N_2095);
nand U2305 (N_2305,N_2211,N_2122);
or U2306 (N_2306,N_2084,N_2232);
and U2307 (N_2307,N_2173,N_2147);
xnor U2308 (N_2308,N_2230,N_2198);
nor U2309 (N_2309,N_2185,N_2200);
and U2310 (N_2310,N_2231,N_2149);
or U2311 (N_2311,N_2234,N_2115);
xor U2312 (N_2312,N_2109,N_2081);
nand U2313 (N_2313,N_2128,N_2097);
or U2314 (N_2314,N_2089,N_2217);
and U2315 (N_2315,N_2195,N_2146);
nand U2316 (N_2316,N_2181,N_2177);
or U2317 (N_2317,N_2219,N_2171);
or U2318 (N_2318,N_2204,N_2154);
nor U2319 (N_2319,N_2189,N_2094);
nor U2320 (N_2320,N_2187,N_2185);
nor U2321 (N_2321,N_2190,N_2182);
and U2322 (N_2322,N_2234,N_2142);
nor U2323 (N_2323,N_2227,N_2081);
or U2324 (N_2324,N_2207,N_2150);
xnor U2325 (N_2325,N_2135,N_2161);
xnor U2326 (N_2326,N_2207,N_2105);
nand U2327 (N_2327,N_2222,N_2101);
nand U2328 (N_2328,N_2107,N_2206);
and U2329 (N_2329,N_2183,N_2184);
and U2330 (N_2330,N_2228,N_2157);
and U2331 (N_2331,N_2177,N_2140);
or U2332 (N_2332,N_2230,N_2165);
or U2333 (N_2333,N_2184,N_2134);
xnor U2334 (N_2334,N_2134,N_2119);
or U2335 (N_2335,N_2178,N_2215);
xor U2336 (N_2336,N_2125,N_2198);
and U2337 (N_2337,N_2182,N_2180);
xor U2338 (N_2338,N_2229,N_2190);
nor U2339 (N_2339,N_2189,N_2226);
nor U2340 (N_2340,N_2202,N_2166);
or U2341 (N_2341,N_2169,N_2180);
xnor U2342 (N_2342,N_2223,N_2194);
and U2343 (N_2343,N_2216,N_2147);
and U2344 (N_2344,N_2147,N_2187);
nand U2345 (N_2345,N_2151,N_2154);
xnor U2346 (N_2346,N_2187,N_2163);
xor U2347 (N_2347,N_2097,N_2124);
nand U2348 (N_2348,N_2205,N_2121);
nor U2349 (N_2349,N_2149,N_2189);
nor U2350 (N_2350,N_2219,N_2177);
xor U2351 (N_2351,N_2178,N_2232);
xnor U2352 (N_2352,N_2090,N_2113);
nor U2353 (N_2353,N_2130,N_2139);
nand U2354 (N_2354,N_2108,N_2190);
nand U2355 (N_2355,N_2139,N_2145);
xor U2356 (N_2356,N_2211,N_2170);
nand U2357 (N_2357,N_2082,N_2085);
nor U2358 (N_2358,N_2192,N_2199);
nor U2359 (N_2359,N_2098,N_2099);
or U2360 (N_2360,N_2130,N_2113);
and U2361 (N_2361,N_2116,N_2120);
and U2362 (N_2362,N_2239,N_2218);
or U2363 (N_2363,N_2114,N_2230);
nor U2364 (N_2364,N_2227,N_2091);
xor U2365 (N_2365,N_2174,N_2162);
xor U2366 (N_2366,N_2116,N_2087);
and U2367 (N_2367,N_2209,N_2117);
nor U2368 (N_2368,N_2179,N_2109);
nor U2369 (N_2369,N_2096,N_2108);
and U2370 (N_2370,N_2155,N_2176);
xor U2371 (N_2371,N_2121,N_2108);
nand U2372 (N_2372,N_2185,N_2196);
xor U2373 (N_2373,N_2193,N_2222);
xnor U2374 (N_2374,N_2185,N_2092);
and U2375 (N_2375,N_2224,N_2142);
or U2376 (N_2376,N_2205,N_2152);
or U2377 (N_2377,N_2104,N_2187);
and U2378 (N_2378,N_2080,N_2125);
or U2379 (N_2379,N_2092,N_2081);
or U2380 (N_2380,N_2201,N_2186);
xor U2381 (N_2381,N_2131,N_2090);
nor U2382 (N_2382,N_2147,N_2119);
and U2383 (N_2383,N_2218,N_2143);
and U2384 (N_2384,N_2111,N_2230);
and U2385 (N_2385,N_2161,N_2227);
nand U2386 (N_2386,N_2177,N_2129);
nand U2387 (N_2387,N_2143,N_2139);
xnor U2388 (N_2388,N_2143,N_2237);
nor U2389 (N_2389,N_2110,N_2216);
nand U2390 (N_2390,N_2089,N_2199);
xnor U2391 (N_2391,N_2127,N_2175);
and U2392 (N_2392,N_2183,N_2179);
and U2393 (N_2393,N_2130,N_2151);
nor U2394 (N_2394,N_2191,N_2096);
and U2395 (N_2395,N_2232,N_2116);
nand U2396 (N_2396,N_2108,N_2128);
and U2397 (N_2397,N_2145,N_2186);
xnor U2398 (N_2398,N_2156,N_2184);
xnor U2399 (N_2399,N_2218,N_2181);
nor U2400 (N_2400,N_2388,N_2391);
and U2401 (N_2401,N_2291,N_2346);
and U2402 (N_2402,N_2331,N_2271);
nor U2403 (N_2403,N_2371,N_2365);
and U2404 (N_2404,N_2304,N_2256);
nor U2405 (N_2405,N_2343,N_2330);
or U2406 (N_2406,N_2265,N_2281);
nand U2407 (N_2407,N_2298,N_2288);
and U2408 (N_2408,N_2351,N_2257);
xnor U2409 (N_2409,N_2325,N_2277);
or U2410 (N_2410,N_2251,N_2312);
xnor U2411 (N_2411,N_2374,N_2393);
and U2412 (N_2412,N_2320,N_2395);
and U2413 (N_2413,N_2369,N_2250);
xnor U2414 (N_2414,N_2302,N_2254);
or U2415 (N_2415,N_2295,N_2241);
nor U2416 (N_2416,N_2396,N_2287);
nand U2417 (N_2417,N_2384,N_2247);
and U2418 (N_2418,N_2379,N_2367);
nor U2419 (N_2419,N_2267,N_2318);
nand U2420 (N_2420,N_2337,N_2344);
nand U2421 (N_2421,N_2305,N_2336);
nor U2422 (N_2422,N_2268,N_2355);
or U2423 (N_2423,N_2249,N_2399);
nor U2424 (N_2424,N_2332,N_2273);
nor U2425 (N_2425,N_2259,N_2317);
nor U2426 (N_2426,N_2240,N_2263);
and U2427 (N_2427,N_2370,N_2276);
nand U2428 (N_2428,N_2313,N_2326);
or U2429 (N_2429,N_2359,N_2286);
xnor U2430 (N_2430,N_2368,N_2375);
nand U2431 (N_2431,N_2348,N_2269);
and U2432 (N_2432,N_2307,N_2342);
or U2433 (N_2433,N_2303,N_2309);
xnor U2434 (N_2434,N_2341,N_2306);
nand U2435 (N_2435,N_2258,N_2279);
nor U2436 (N_2436,N_2333,N_2293);
and U2437 (N_2437,N_2297,N_2386);
nor U2438 (N_2438,N_2296,N_2261);
xnor U2439 (N_2439,N_2382,N_2270);
and U2440 (N_2440,N_2262,N_2289);
and U2441 (N_2441,N_2278,N_2314);
nor U2442 (N_2442,N_2397,N_2358);
and U2443 (N_2443,N_2310,N_2315);
or U2444 (N_2444,N_2377,N_2274);
and U2445 (N_2445,N_2345,N_2383);
nand U2446 (N_2446,N_2373,N_2389);
nand U2447 (N_2447,N_2280,N_2316);
nand U2448 (N_2448,N_2311,N_2308);
nor U2449 (N_2449,N_2243,N_2329);
and U2450 (N_2450,N_2285,N_2275);
nor U2451 (N_2451,N_2248,N_2290);
and U2452 (N_2452,N_2380,N_2284);
nand U2453 (N_2453,N_2321,N_2398);
nand U2454 (N_2454,N_2323,N_2294);
and U2455 (N_2455,N_2299,N_2361);
xor U2456 (N_2456,N_2252,N_2354);
xor U2457 (N_2457,N_2327,N_2292);
or U2458 (N_2458,N_2264,N_2253);
nand U2459 (N_2459,N_2366,N_2272);
xor U2460 (N_2460,N_2363,N_2300);
xnor U2461 (N_2461,N_2376,N_2356);
xor U2462 (N_2462,N_2352,N_2378);
nor U2463 (N_2463,N_2357,N_2266);
and U2464 (N_2464,N_2334,N_2381);
nand U2465 (N_2465,N_2349,N_2372);
and U2466 (N_2466,N_2244,N_2260);
nor U2467 (N_2467,N_2283,N_2353);
or U2468 (N_2468,N_2347,N_2245);
nor U2469 (N_2469,N_2392,N_2385);
and U2470 (N_2470,N_2242,N_2324);
nand U2471 (N_2471,N_2301,N_2362);
nand U2472 (N_2472,N_2335,N_2394);
nor U2473 (N_2473,N_2282,N_2340);
and U2474 (N_2474,N_2319,N_2338);
nand U2475 (N_2475,N_2350,N_2328);
nor U2476 (N_2476,N_2390,N_2246);
and U2477 (N_2477,N_2255,N_2322);
and U2478 (N_2478,N_2387,N_2360);
xnor U2479 (N_2479,N_2339,N_2364);
xor U2480 (N_2480,N_2262,N_2285);
nand U2481 (N_2481,N_2304,N_2348);
nand U2482 (N_2482,N_2304,N_2331);
nand U2483 (N_2483,N_2295,N_2281);
or U2484 (N_2484,N_2360,N_2301);
nand U2485 (N_2485,N_2328,N_2390);
nand U2486 (N_2486,N_2304,N_2383);
xor U2487 (N_2487,N_2376,N_2398);
and U2488 (N_2488,N_2260,N_2347);
nor U2489 (N_2489,N_2356,N_2367);
nand U2490 (N_2490,N_2392,N_2253);
and U2491 (N_2491,N_2270,N_2255);
xnor U2492 (N_2492,N_2394,N_2308);
xnor U2493 (N_2493,N_2335,N_2247);
or U2494 (N_2494,N_2385,N_2368);
nand U2495 (N_2495,N_2263,N_2363);
nor U2496 (N_2496,N_2365,N_2370);
or U2497 (N_2497,N_2350,N_2335);
nor U2498 (N_2498,N_2383,N_2322);
xor U2499 (N_2499,N_2335,N_2311);
or U2500 (N_2500,N_2349,N_2241);
and U2501 (N_2501,N_2293,N_2260);
and U2502 (N_2502,N_2375,N_2328);
nand U2503 (N_2503,N_2354,N_2360);
nor U2504 (N_2504,N_2312,N_2302);
xnor U2505 (N_2505,N_2385,N_2343);
and U2506 (N_2506,N_2380,N_2353);
xor U2507 (N_2507,N_2399,N_2393);
and U2508 (N_2508,N_2260,N_2367);
nor U2509 (N_2509,N_2324,N_2337);
xnor U2510 (N_2510,N_2357,N_2271);
nor U2511 (N_2511,N_2259,N_2396);
nor U2512 (N_2512,N_2396,N_2348);
nor U2513 (N_2513,N_2276,N_2333);
nor U2514 (N_2514,N_2312,N_2396);
and U2515 (N_2515,N_2321,N_2362);
and U2516 (N_2516,N_2390,N_2388);
nand U2517 (N_2517,N_2272,N_2314);
nand U2518 (N_2518,N_2337,N_2302);
xor U2519 (N_2519,N_2321,N_2371);
nor U2520 (N_2520,N_2398,N_2307);
nor U2521 (N_2521,N_2328,N_2299);
nor U2522 (N_2522,N_2335,N_2244);
nand U2523 (N_2523,N_2250,N_2360);
xnor U2524 (N_2524,N_2249,N_2326);
xor U2525 (N_2525,N_2319,N_2330);
and U2526 (N_2526,N_2292,N_2281);
xor U2527 (N_2527,N_2286,N_2256);
or U2528 (N_2528,N_2352,N_2364);
nor U2529 (N_2529,N_2377,N_2297);
nand U2530 (N_2530,N_2371,N_2364);
xnor U2531 (N_2531,N_2245,N_2330);
nor U2532 (N_2532,N_2347,N_2310);
xor U2533 (N_2533,N_2245,N_2264);
nand U2534 (N_2534,N_2276,N_2350);
or U2535 (N_2535,N_2382,N_2272);
nand U2536 (N_2536,N_2322,N_2352);
nor U2537 (N_2537,N_2329,N_2386);
or U2538 (N_2538,N_2376,N_2304);
xor U2539 (N_2539,N_2359,N_2395);
and U2540 (N_2540,N_2303,N_2367);
or U2541 (N_2541,N_2301,N_2329);
nand U2542 (N_2542,N_2275,N_2386);
or U2543 (N_2543,N_2308,N_2359);
nor U2544 (N_2544,N_2356,N_2281);
xor U2545 (N_2545,N_2309,N_2310);
or U2546 (N_2546,N_2289,N_2285);
xnor U2547 (N_2547,N_2281,N_2276);
nand U2548 (N_2548,N_2247,N_2339);
or U2549 (N_2549,N_2373,N_2388);
and U2550 (N_2550,N_2342,N_2339);
nand U2551 (N_2551,N_2390,N_2301);
and U2552 (N_2552,N_2359,N_2370);
and U2553 (N_2553,N_2336,N_2357);
or U2554 (N_2554,N_2308,N_2327);
nor U2555 (N_2555,N_2321,N_2270);
and U2556 (N_2556,N_2298,N_2389);
and U2557 (N_2557,N_2393,N_2297);
and U2558 (N_2558,N_2388,N_2273);
xnor U2559 (N_2559,N_2242,N_2312);
xor U2560 (N_2560,N_2425,N_2505);
xor U2561 (N_2561,N_2531,N_2480);
xor U2562 (N_2562,N_2548,N_2522);
nor U2563 (N_2563,N_2420,N_2419);
or U2564 (N_2564,N_2513,N_2549);
xnor U2565 (N_2565,N_2557,N_2401);
nor U2566 (N_2566,N_2451,N_2430);
or U2567 (N_2567,N_2413,N_2539);
nand U2568 (N_2568,N_2551,N_2527);
or U2569 (N_2569,N_2544,N_2494);
and U2570 (N_2570,N_2418,N_2448);
or U2571 (N_2571,N_2538,N_2407);
and U2572 (N_2572,N_2443,N_2499);
nor U2573 (N_2573,N_2543,N_2450);
nand U2574 (N_2574,N_2445,N_2537);
nor U2575 (N_2575,N_2508,N_2486);
nor U2576 (N_2576,N_2502,N_2545);
or U2577 (N_2577,N_2492,N_2468);
or U2578 (N_2578,N_2403,N_2462);
or U2579 (N_2579,N_2410,N_2520);
and U2580 (N_2580,N_2481,N_2479);
xor U2581 (N_2581,N_2446,N_2510);
and U2582 (N_2582,N_2516,N_2536);
xnor U2583 (N_2583,N_2442,N_2409);
nand U2584 (N_2584,N_2421,N_2506);
or U2585 (N_2585,N_2554,N_2412);
nor U2586 (N_2586,N_2532,N_2438);
nor U2587 (N_2587,N_2555,N_2461);
and U2588 (N_2588,N_2435,N_2464);
nor U2589 (N_2589,N_2476,N_2535);
and U2590 (N_2590,N_2434,N_2427);
or U2591 (N_2591,N_2511,N_2541);
nor U2592 (N_2592,N_2433,N_2415);
and U2593 (N_2593,N_2416,N_2493);
nor U2594 (N_2594,N_2467,N_2422);
and U2595 (N_2595,N_2524,N_2424);
or U2596 (N_2596,N_2437,N_2517);
nor U2597 (N_2597,N_2463,N_2518);
xor U2598 (N_2598,N_2414,N_2485);
nor U2599 (N_2599,N_2455,N_2509);
nor U2600 (N_2600,N_2441,N_2503);
and U2601 (N_2601,N_2497,N_2496);
xor U2602 (N_2602,N_2552,N_2526);
nand U2603 (N_2603,N_2457,N_2498);
nand U2604 (N_2604,N_2491,N_2453);
or U2605 (N_2605,N_2533,N_2550);
or U2606 (N_2606,N_2515,N_2487);
nand U2607 (N_2607,N_2436,N_2473);
or U2608 (N_2608,N_2482,N_2556);
nor U2609 (N_2609,N_2547,N_2456);
or U2610 (N_2610,N_2472,N_2452);
xnor U2611 (N_2611,N_2404,N_2469);
or U2612 (N_2612,N_2426,N_2530);
xnor U2613 (N_2613,N_2558,N_2478);
or U2614 (N_2614,N_2460,N_2519);
nor U2615 (N_2615,N_2459,N_2559);
and U2616 (N_2616,N_2440,N_2408);
nand U2617 (N_2617,N_2484,N_2458);
and U2618 (N_2618,N_2449,N_2495);
or U2619 (N_2619,N_2504,N_2488);
or U2620 (N_2620,N_2411,N_2529);
or U2621 (N_2621,N_2444,N_2470);
nand U2622 (N_2622,N_2525,N_2507);
or U2623 (N_2623,N_2490,N_2534);
nand U2624 (N_2624,N_2501,N_2475);
nand U2625 (N_2625,N_2489,N_2432);
nor U2626 (N_2626,N_2454,N_2528);
and U2627 (N_2627,N_2429,N_2514);
or U2628 (N_2628,N_2540,N_2521);
nor U2629 (N_2629,N_2474,N_2406);
nand U2630 (N_2630,N_2546,N_2405);
xnor U2631 (N_2631,N_2542,N_2465);
and U2632 (N_2632,N_2431,N_2439);
xor U2633 (N_2633,N_2417,N_2428);
nand U2634 (N_2634,N_2400,N_2483);
and U2635 (N_2635,N_2553,N_2500);
nand U2636 (N_2636,N_2466,N_2477);
nor U2637 (N_2637,N_2423,N_2447);
nor U2638 (N_2638,N_2402,N_2471);
and U2639 (N_2639,N_2512,N_2523);
xnor U2640 (N_2640,N_2490,N_2438);
xor U2641 (N_2641,N_2502,N_2441);
xor U2642 (N_2642,N_2413,N_2430);
nor U2643 (N_2643,N_2526,N_2541);
or U2644 (N_2644,N_2460,N_2504);
nor U2645 (N_2645,N_2559,N_2529);
xnor U2646 (N_2646,N_2468,N_2464);
xor U2647 (N_2647,N_2477,N_2518);
and U2648 (N_2648,N_2454,N_2482);
or U2649 (N_2649,N_2447,N_2495);
and U2650 (N_2650,N_2453,N_2450);
nor U2651 (N_2651,N_2513,N_2476);
or U2652 (N_2652,N_2488,N_2419);
xor U2653 (N_2653,N_2431,N_2437);
nor U2654 (N_2654,N_2427,N_2499);
or U2655 (N_2655,N_2455,N_2553);
and U2656 (N_2656,N_2423,N_2555);
nor U2657 (N_2657,N_2480,N_2470);
or U2658 (N_2658,N_2541,N_2521);
nand U2659 (N_2659,N_2558,N_2462);
or U2660 (N_2660,N_2432,N_2426);
xnor U2661 (N_2661,N_2461,N_2403);
nor U2662 (N_2662,N_2467,N_2538);
nor U2663 (N_2663,N_2531,N_2509);
or U2664 (N_2664,N_2549,N_2412);
nor U2665 (N_2665,N_2443,N_2528);
and U2666 (N_2666,N_2520,N_2423);
and U2667 (N_2667,N_2502,N_2508);
nand U2668 (N_2668,N_2467,N_2493);
nor U2669 (N_2669,N_2436,N_2416);
and U2670 (N_2670,N_2479,N_2439);
nor U2671 (N_2671,N_2454,N_2538);
nand U2672 (N_2672,N_2401,N_2418);
nand U2673 (N_2673,N_2416,N_2490);
or U2674 (N_2674,N_2512,N_2440);
nand U2675 (N_2675,N_2499,N_2466);
xnor U2676 (N_2676,N_2426,N_2450);
xnor U2677 (N_2677,N_2551,N_2533);
nor U2678 (N_2678,N_2493,N_2473);
or U2679 (N_2679,N_2446,N_2474);
nor U2680 (N_2680,N_2478,N_2413);
nor U2681 (N_2681,N_2458,N_2548);
or U2682 (N_2682,N_2404,N_2455);
nor U2683 (N_2683,N_2482,N_2483);
nand U2684 (N_2684,N_2410,N_2508);
nor U2685 (N_2685,N_2412,N_2413);
or U2686 (N_2686,N_2546,N_2492);
nand U2687 (N_2687,N_2534,N_2443);
nor U2688 (N_2688,N_2552,N_2481);
or U2689 (N_2689,N_2512,N_2411);
nand U2690 (N_2690,N_2421,N_2482);
nand U2691 (N_2691,N_2451,N_2515);
nand U2692 (N_2692,N_2476,N_2480);
and U2693 (N_2693,N_2521,N_2538);
and U2694 (N_2694,N_2465,N_2458);
nor U2695 (N_2695,N_2488,N_2463);
nor U2696 (N_2696,N_2455,N_2447);
nand U2697 (N_2697,N_2443,N_2437);
nor U2698 (N_2698,N_2511,N_2465);
or U2699 (N_2699,N_2488,N_2431);
nand U2700 (N_2700,N_2530,N_2434);
nand U2701 (N_2701,N_2534,N_2435);
and U2702 (N_2702,N_2493,N_2486);
nor U2703 (N_2703,N_2422,N_2409);
xor U2704 (N_2704,N_2549,N_2419);
xor U2705 (N_2705,N_2522,N_2430);
xor U2706 (N_2706,N_2446,N_2454);
nor U2707 (N_2707,N_2424,N_2532);
and U2708 (N_2708,N_2476,N_2538);
xor U2709 (N_2709,N_2418,N_2438);
xnor U2710 (N_2710,N_2553,N_2423);
and U2711 (N_2711,N_2502,N_2485);
nor U2712 (N_2712,N_2454,N_2498);
nor U2713 (N_2713,N_2433,N_2452);
or U2714 (N_2714,N_2496,N_2426);
or U2715 (N_2715,N_2477,N_2559);
nand U2716 (N_2716,N_2452,N_2438);
nor U2717 (N_2717,N_2404,N_2422);
xor U2718 (N_2718,N_2482,N_2505);
and U2719 (N_2719,N_2556,N_2454);
xnor U2720 (N_2720,N_2695,N_2579);
nand U2721 (N_2721,N_2565,N_2657);
xnor U2722 (N_2722,N_2700,N_2696);
or U2723 (N_2723,N_2713,N_2701);
and U2724 (N_2724,N_2560,N_2603);
nand U2725 (N_2725,N_2660,N_2655);
or U2726 (N_2726,N_2654,N_2709);
xnor U2727 (N_2727,N_2704,N_2712);
nor U2728 (N_2728,N_2593,N_2635);
or U2729 (N_2729,N_2594,N_2698);
nand U2730 (N_2730,N_2685,N_2597);
xor U2731 (N_2731,N_2591,N_2581);
or U2732 (N_2732,N_2584,N_2681);
or U2733 (N_2733,N_2624,N_2562);
nor U2734 (N_2734,N_2566,N_2630);
or U2735 (N_2735,N_2610,N_2673);
xnor U2736 (N_2736,N_2592,N_2568);
nor U2737 (N_2737,N_2690,N_2598);
or U2738 (N_2738,N_2662,N_2634);
or U2739 (N_2739,N_2645,N_2602);
xnor U2740 (N_2740,N_2715,N_2661);
nor U2741 (N_2741,N_2621,N_2684);
and U2742 (N_2742,N_2649,N_2596);
xnor U2743 (N_2743,N_2650,N_2705);
xnor U2744 (N_2744,N_2719,N_2651);
xnor U2745 (N_2745,N_2615,N_2676);
and U2746 (N_2746,N_2692,N_2702);
and U2747 (N_2747,N_2699,N_2595);
nor U2748 (N_2748,N_2665,N_2711);
nand U2749 (N_2749,N_2672,N_2618);
and U2750 (N_2750,N_2613,N_2611);
nand U2751 (N_2751,N_2687,N_2664);
nor U2752 (N_2752,N_2653,N_2586);
xnor U2753 (N_2753,N_2628,N_2606);
or U2754 (N_2754,N_2648,N_2589);
or U2755 (N_2755,N_2638,N_2622);
or U2756 (N_2756,N_2605,N_2583);
nand U2757 (N_2757,N_2604,N_2639);
xnor U2758 (N_2758,N_2693,N_2626);
xnor U2759 (N_2759,N_2572,N_2563);
or U2760 (N_2760,N_2619,N_2679);
nor U2761 (N_2761,N_2683,N_2616);
or U2762 (N_2762,N_2682,N_2688);
or U2763 (N_2763,N_2674,N_2590);
xnor U2764 (N_2764,N_2620,N_2642);
nor U2765 (N_2765,N_2564,N_2625);
xor U2766 (N_2766,N_2675,N_2636);
and U2767 (N_2767,N_2580,N_2627);
nand U2768 (N_2768,N_2570,N_2710);
xnor U2769 (N_2769,N_2656,N_2680);
or U2770 (N_2770,N_2574,N_2718);
or U2771 (N_2771,N_2666,N_2678);
nand U2772 (N_2772,N_2641,N_2608);
or U2773 (N_2773,N_2575,N_2670);
nor U2774 (N_2774,N_2640,N_2631);
xor U2775 (N_2775,N_2647,N_2694);
nor U2776 (N_2776,N_2677,N_2609);
nor U2777 (N_2777,N_2629,N_2686);
nand U2778 (N_2778,N_2567,N_2714);
and U2779 (N_2779,N_2614,N_2703);
or U2780 (N_2780,N_2600,N_2617);
nand U2781 (N_2781,N_2599,N_2659);
nor U2782 (N_2782,N_2671,N_2646);
and U2783 (N_2783,N_2587,N_2668);
or U2784 (N_2784,N_2585,N_2578);
and U2785 (N_2785,N_2588,N_2667);
xor U2786 (N_2786,N_2577,N_2632);
and U2787 (N_2787,N_2644,N_2571);
nor U2788 (N_2788,N_2689,N_2569);
or U2789 (N_2789,N_2633,N_2717);
xor U2790 (N_2790,N_2582,N_2658);
and U2791 (N_2791,N_2637,N_2707);
or U2792 (N_2792,N_2669,N_2612);
xnor U2793 (N_2793,N_2697,N_2716);
and U2794 (N_2794,N_2652,N_2561);
and U2795 (N_2795,N_2623,N_2601);
xnor U2796 (N_2796,N_2576,N_2691);
and U2797 (N_2797,N_2643,N_2706);
nand U2798 (N_2798,N_2663,N_2607);
or U2799 (N_2799,N_2708,N_2573);
nand U2800 (N_2800,N_2670,N_2700);
nor U2801 (N_2801,N_2699,N_2676);
nand U2802 (N_2802,N_2611,N_2586);
nor U2803 (N_2803,N_2664,N_2646);
nor U2804 (N_2804,N_2682,N_2663);
and U2805 (N_2805,N_2598,N_2563);
and U2806 (N_2806,N_2705,N_2605);
nand U2807 (N_2807,N_2567,N_2687);
nand U2808 (N_2808,N_2715,N_2610);
and U2809 (N_2809,N_2700,N_2682);
nand U2810 (N_2810,N_2663,N_2679);
and U2811 (N_2811,N_2713,N_2646);
and U2812 (N_2812,N_2707,N_2656);
nor U2813 (N_2813,N_2630,N_2640);
xnor U2814 (N_2814,N_2710,N_2719);
or U2815 (N_2815,N_2616,N_2654);
and U2816 (N_2816,N_2683,N_2588);
nor U2817 (N_2817,N_2622,N_2603);
or U2818 (N_2818,N_2599,N_2696);
xor U2819 (N_2819,N_2627,N_2676);
and U2820 (N_2820,N_2681,N_2706);
xor U2821 (N_2821,N_2596,N_2678);
nor U2822 (N_2822,N_2663,N_2575);
nand U2823 (N_2823,N_2652,N_2666);
or U2824 (N_2824,N_2600,N_2692);
or U2825 (N_2825,N_2675,N_2587);
or U2826 (N_2826,N_2597,N_2622);
nand U2827 (N_2827,N_2665,N_2624);
xor U2828 (N_2828,N_2667,N_2626);
nand U2829 (N_2829,N_2658,N_2587);
xnor U2830 (N_2830,N_2693,N_2707);
xor U2831 (N_2831,N_2653,N_2584);
nor U2832 (N_2832,N_2680,N_2569);
nor U2833 (N_2833,N_2604,N_2584);
or U2834 (N_2834,N_2621,N_2579);
xnor U2835 (N_2835,N_2569,N_2660);
and U2836 (N_2836,N_2643,N_2702);
nand U2837 (N_2837,N_2571,N_2705);
xor U2838 (N_2838,N_2593,N_2671);
nor U2839 (N_2839,N_2635,N_2599);
nand U2840 (N_2840,N_2572,N_2643);
and U2841 (N_2841,N_2677,N_2628);
nor U2842 (N_2842,N_2705,N_2676);
and U2843 (N_2843,N_2622,N_2652);
nor U2844 (N_2844,N_2630,N_2598);
or U2845 (N_2845,N_2711,N_2717);
or U2846 (N_2846,N_2634,N_2686);
or U2847 (N_2847,N_2719,N_2677);
and U2848 (N_2848,N_2595,N_2684);
and U2849 (N_2849,N_2606,N_2686);
xnor U2850 (N_2850,N_2598,N_2620);
nor U2851 (N_2851,N_2563,N_2657);
nor U2852 (N_2852,N_2567,N_2683);
and U2853 (N_2853,N_2661,N_2704);
xnor U2854 (N_2854,N_2573,N_2603);
and U2855 (N_2855,N_2597,N_2626);
nor U2856 (N_2856,N_2648,N_2699);
or U2857 (N_2857,N_2610,N_2650);
xnor U2858 (N_2858,N_2711,N_2660);
or U2859 (N_2859,N_2616,N_2700);
nor U2860 (N_2860,N_2650,N_2678);
xnor U2861 (N_2861,N_2639,N_2704);
nor U2862 (N_2862,N_2632,N_2713);
nor U2863 (N_2863,N_2675,N_2669);
nand U2864 (N_2864,N_2644,N_2630);
xor U2865 (N_2865,N_2569,N_2717);
nor U2866 (N_2866,N_2676,N_2709);
nor U2867 (N_2867,N_2644,N_2703);
xnor U2868 (N_2868,N_2591,N_2622);
nand U2869 (N_2869,N_2659,N_2629);
nor U2870 (N_2870,N_2698,N_2560);
nor U2871 (N_2871,N_2687,N_2632);
or U2872 (N_2872,N_2601,N_2574);
or U2873 (N_2873,N_2620,N_2635);
or U2874 (N_2874,N_2614,N_2654);
and U2875 (N_2875,N_2700,N_2650);
nand U2876 (N_2876,N_2592,N_2586);
nand U2877 (N_2877,N_2606,N_2719);
xnor U2878 (N_2878,N_2696,N_2623);
or U2879 (N_2879,N_2560,N_2697);
and U2880 (N_2880,N_2878,N_2831);
xor U2881 (N_2881,N_2864,N_2736);
xor U2882 (N_2882,N_2861,N_2851);
xnor U2883 (N_2883,N_2769,N_2801);
and U2884 (N_2884,N_2839,N_2863);
xor U2885 (N_2885,N_2819,N_2722);
nand U2886 (N_2886,N_2744,N_2724);
xor U2887 (N_2887,N_2847,N_2782);
nor U2888 (N_2888,N_2866,N_2867);
nor U2889 (N_2889,N_2793,N_2879);
nand U2890 (N_2890,N_2747,N_2726);
or U2891 (N_2891,N_2737,N_2794);
xor U2892 (N_2892,N_2856,N_2799);
and U2893 (N_2893,N_2837,N_2750);
xnor U2894 (N_2894,N_2760,N_2781);
or U2895 (N_2895,N_2735,N_2874);
or U2896 (N_2896,N_2828,N_2830);
and U2897 (N_2897,N_2877,N_2823);
nor U2898 (N_2898,N_2870,N_2777);
or U2899 (N_2899,N_2836,N_2844);
nor U2900 (N_2900,N_2779,N_2809);
or U2901 (N_2901,N_2827,N_2751);
nor U2902 (N_2902,N_2846,N_2876);
xnor U2903 (N_2903,N_2774,N_2727);
or U2904 (N_2904,N_2868,N_2752);
and U2905 (N_2905,N_2756,N_2832);
nand U2906 (N_2906,N_2817,N_2725);
nand U2907 (N_2907,N_2768,N_2875);
or U2908 (N_2908,N_2742,N_2800);
nor U2909 (N_2909,N_2792,N_2869);
or U2910 (N_2910,N_2871,N_2865);
and U2911 (N_2911,N_2770,N_2841);
or U2912 (N_2912,N_2767,N_2842);
nand U2913 (N_2913,N_2743,N_2855);
or U2914 (N_2914,N_2732,N_2745);
nand U2915 (N_2915,N_2771,N_2807);
and U2916 (N_2916,N_2761,N_2860);
and U2917 (N_2917,N_2797,N_2787);
xnor U2918 (N_2918,N_2723,N_2813);
or U2919 (N_2919,N_2754,N_2795);
and U2920 (N_2920,N_2848,N_2729);
or U2921 (N_2921,N_2812,N_2757);
and U2922 (N_2922,N_2838,N_2721);
and U2923 (N_2923,N_2749,N_2766);
and U2924 (N_2924,N_2759,N_2720);
nand U2925 (N_2925,N_2746,N_2786);
and U2926 (N_2926,N_2840,N_2789);
xnor U2927 (N_2927,N_2784,N_2785);
or U2928 (N_2928,N_2825,N_2776);
or U2929 (N_2929,N_2820,N_2763);
or U2930 (N_2930,N_2740,N_2738);
and U2931 (N_2931,N_2730,N_2733);
nand U2932 (N_2932,N_2802,N_2858);
or U2933 (N_2933,N_2811,N_2857);
and U2934 (N_2934,N_2804,N_2778);
xor U2935 (N_2935,N_2748,N_2835);
or U2936 (N_2936,N_2833,N_2824);
nand U2937 (N_2937,N_2758,N_2826);
or U2938 (N_2938,N_2834,N_2859);
nand U2939 (N_2939,N_2814,N_2852);
nand U2940 (N_2940,N_2765,N_2796);
xor U2941 (N_2941,N_2822,N_2829);
xnor U2942 (N_2942,N_2783,N_2854);
nand U2943 (N_2943,N_2853,N_2788);
nand U2944 (N_2944,N_2808,N_2753);
xor U2945 (N_2945,N_2815,N_2798);
xnor U2946 (N_2946,N_2755,N_2762);
or U2947 (N_2947,N_2873,N_2790);
nand U2948 (N_2948,N_2741,N_2821);
xnor U2949 (N_2949,N_2803,N_2805);
xnor U2950 (N_2950,N_2772,N_2773);
and U2951 (N_2951,N_2791,N_2734);
and U2952 (N_2952,N_2780,N_2806);
or U2953 (N_2953,N_2849,N_2731);
or U2954 (N_2954,N_2728,N_2816);
and U2955 (N_2955,N_2818,N_2810);
or U2956 (N_2956,N_2843,N_2739);
or U2957 (N_2957,N_2862,N_2764);
nor U2958 (N_2958,N_2872,N_2850);
xnor U2959 (N_2959,N_2845,N_2775);
xor U2960 (N_2960,N_2845,N_2810);
xor U2961 (N_2961,N_2842,N_2867);
nand U2962 (N_2962,N_2870,N_2728);
nor U2963 (N_2963,N_2723,N_2748);
or U2964 (N_2964,N_2738,N_2846);
xor U2965 (N_2965,N_2809,N_2870);
xor U2966 (N_2966,N_2731,N_2855);
or U2967 (N_2967,N_2829,N_2857);
and U2968 (N_2968,N_2829,N_2819);
nor U2969 (N_2969,N_2779,N_2792);
and U2970 (N_2970,N_2752,N_2820);
or U2971 (N_2971,N_2872,N_2742);
nor U2972 (N_2972,N_2830,N_2862);
xor U2973 (N_2973,N_2862,N_2760);
nor U2974 (N_2974,N_2787,N_2875);
xor U2975 (N_2975,N_2766,N_2875);
or U2976 (N_2976,N_2863,N_2762);
or U2977 (N_2977,N_2771,N_2838);
xor U2978 (N_2978,N_2843,N_2798);
xnor U2979 (N_2979,N_2770,N_2775);
or U2980 (N_2980,N_2759,N_2844);
and U2981 (N_2981,N_2862,N_2775);
and U2982 (N_2982,N_2790,N_2821);
xor U2983 (N_2983,N_2834,N_2821);
xor U2984 (N_2984,N_2878,N_2730);
and U2985 (N_2985,N_2743,N_2868);
nand U2986 (N_2986,N_2815,N_2734);
or U2987 (N_2987,N_2867,N_2736);
xnor U2988 (N_2988,N_2784,N_2773);
or U2989 (N_2989,N_2816,N_2803);
nand U2990 (N_2990,N_2843,N_2815);
nor U2991 (N_2991,N_2722,N_2876);
nand U2992 (N_2992,N_2872,N_2739);
nor U2993 (N_2993,N_2804,N_2776);
nand U2994 (N_2994,N_2736,N_2808);
nand U2995 (N_2995,N_2878,N_2728);
xnor U2996 (N_2996,N_2767,N_2811);
and U2997 (N_2997,N_2744,N_2813);
xnor U2998 (N_2998,N_2805,N_2873);
nor U2999 (N_2999,N_2744,N_2741);
and U3000 (N_3000,N_2740,N_2793);
nor U3001 (N_3001,N_2848,N_2777);
nor U3002 (N_3002,N_2796,N_2741);
nor U3003 (N_3003,N_2769,N_2853);
xor U3004 (N_3004,N_2747,N_2869);
nor U3005 (N_3005,N_2783,N_2779);
nand U3006 (N_3006,N_2748,N_2760);
and U3007 (N_3007,N_2841,N_2781);
nand U3008 (N_3008,N_2759,N_2783);
xnor U3009 (N_3009,N_2835,N_2804);
nor U3010 (N_3010,N_2831,N_2835);
and U3011 (N_3011,N_2771,N_2784);
nor U3012 (N_3012,N_2865,N_2863);
nand U3013 (N_3013,N_2827,N_2723);
and U3014 (N_3014,N_2757,N_2794);
or U3015 (N_3015,N_2869,N_2814);
xor U3016 (N_3016,N_2752,N_2864);
or U3017 (N_3017,N_2872,N_2799);
or U3018 (N_3018,N_2756,N_2821);
nand U3019 (N_3019,N_2878,N_2750);
xnor U3020 (N_3020,N_2789,N_2820);
and U3021 (N_3021,N_2749,N_2794);
nand U3022 (N_3022,N_2773,N_2824);
nor U3023 (N_3023,N_2725,N_2864);
nor U3024 (N_3024,N_2842,N_2752);
nand U3025 (N_3025,N_2769,N_2878);
and U3026 (N_3026,N_2814,N_2782);
nand U3027 (N_3027,N_2851,N_2816);
or U3028 (N_3028,N_2743,N_2730);
and U3029 (N_3029,N_2873,N_2838);
nor U3030 (N_3030,N_2723,N_2793);
or U3031 (N_3031,N_2849,N_2864);
xor U3032 (N_3032,N_2877,N_2796);
and U3033 (N_3033,N_2875,N_2770);
or U3034 (N_3034,N_2832,N_2768);
nand U3035 (N_3035,N_2815,N_2745);
or U3036 (N_3036,N_2806,N_2805);
xor U3037 (N_3037,N_2840,N_2779);
nor U3038 (N_3038,N_2807,N_2732);
or U3039 (N_3039,N_2737,N_2777);
and U3040 (N_3040,N_2933,N_2883);
nand U3041 (N_3041,N_2992,N_2924);
nor U3042 (N_3042,N_3007,N_3023);
and U3043 (N_3043,N_3028,N_2891);
nand U3044 (N_3044,N_2984,N_2882);
nand U3045 (N_3045,N_2903,N_2918);
nor U3046 (N_3046,N_2970,N_3013);
nor U3047 (N_3047,N_2943,N_2885);
nand U3048 (N_3048,N_2990,N_2893);
xnor U3049 (N_3049,N_3027,N_2892);
xnor U3050 (N_3050,N_3006,N_3009);
nor U3051 (N_3051,N_2911,N_2922);
xor U3052 (N_3052,N_3024,N_2958);
and U3053 (N_3053,N_3016,N_2898);
or U3054 (N_3054,N_3026,N_2965);
and U3055 (N_3055,N_2960,N_2962);
xor U3056 (N_3056,N_3022,N_2988);
nand U3057 (N_3057,N_2953,N_3029);
and U3058 (N_3058,N_2944,N_3019);
nor U3059 (N_3059,N_3005,N_2904);
nor U3060 (N_3060,N_2895,N_2975);
and U3061 (N_3061,N_2951,N_2963);
nand U3062 (N_3062,N_2930,N_2952);
nor U3063 (N_3063,N_2914,N_2995);
nor U3064 (N_3064,N_3014,N_3017);
nand U3065 (N_3065,N_3039,N_2939);
nor U3066 (N_3066,N_2964,N_3034);
and U3067 (N_3067,N_3030,N_2957);
and U3068 (N_3068,N_3003,N_2881);
nor U3069 (N_3069,N_3025,N_2966);
or U3070 (N_3070,N_3011,N_2968);
nand U3071 (N_3071,N_2880,N_2982);
xnor U3072 (N_3072,N_3032,N_2997);
or U3073 (N_3073,N_3001,N_2907);
xor U3074 (N_3074,N_2999,N_2991);
nor U3075 (N_3075,N_2925,N_3031);
and U3076 (N_3076,N_2886,N_2902);
or U3077 (N_3077,N_2942,N_2905);
xnor U3078 (N_3078,N_2910,N_2938);
nor U3079 (N_3079,N_3033,N_3038);
or U3080 (N_3080,N_3035,N_2940);
xor U3081 (N_3081,N_2912,N_2976);
and U3082 (N_3082,N_2889,N_3021);
nand U3083 (N_3083,N_2916,N_3000);
nand U3084 (N_3084,N_2980,N_2989);
nor U3085 (N_3085,N_2927,N_2983);
or U3086 (N_3086,N_2979,N_2923);
nand U3087 (N_3087,N_2937,N_3002);
nand U3088 (N_3088,N_2974,N_2972);
or U3089 (N_3089,N_2906,N_2919);
xnor U3090 (N_3090,N_2948,N_2971);
and U3091 (N_3091,N_2977,N_2978);
nor U3092 (N_3092,N_2967,N_2993);
and U3093 (N_3093,N_2949,N_3004);
nand U3094 (N_3094,N_2956,N_2913);
xor U3095 (N_3095,N_2934,N_2920);
and U3096 (N_3096,N_2887,N_2955);
xnor U3097 (N_3097,N_2929,N_2896);
xor U3098 (N_3098,N_3020,N_3008);
or U3099 (N_3099,N_2909,N_2917);
xor U3100 (N_3100,N_2959,N_2946);
xor U3101 (N_3101,N_2994,N_3015);
nor U3102 (N_3102,N_2888,N_3010);
or U3103 (N_3103,N_2969,N_2973);
nor U3104 (N_3104,N_2915,N_2901);
nor U3105 (N_3105,N_2900,N_2897);
xnor U3106 (N_3106,N_2986,N_2981);
nand U3107 (N_3107,N_2954,N_2921);
xnor U3108 (N_3108,N_2926,N_3018);
xor U3109 (N_3109,N_2941,N_2935);
and U3110 (N_3110,N_2931,N_2884);
xor U3111 (N_3111,N_2932,N_2996);
nand U3112 (N_3112,N_2985,N_2945);
and U3113 (N_3113,N_2928,N_2890);
xor U3114 (N_3114,N_2998,N_2908);
nand U3115 (N_3115,N_2961,N_2987);
nor U3116 (N_3116,N_2899,N_2950);
nor U3117 (N_3117,N_2936,N_3036);
and U3118 (N_3118,N_3012,N_2894);
nor U3119 (N_3119,N_2947,N_3037);
xnor U3120 (N_3120,N_2922,N_2943);
and U3121 (N_3121,N_2977,N_2893);
nor U3122 (N_3122,N_2997,N_2991);
nor U3123 (N_3123,N_2914,N_3016);
or U3124 (N_3124,N_2883,N_2909);
nor U3125 (N_3125,N_2933,N_2959);
or U3126 (N_3126,N_2928,N_2964);
or U3127 (N_3127,N_2956,N_2899);
nor U3128 (N_3128,N_3022,N_2886);
or U3129 (N_3129,N_2910,N_2965);
or U3130 (N_3130,N_3026,N_3017);
and U3131 (N_3131,N_2894,N_3027);
nor U3132 (N_3132,N_3039,N_3009);
and U3133 (N_3133,N_2964,N_2923);
or U3134 (N_3134,N_3006,N_2925);
xnor U3135 (N_3135,N_2994,N_2888);
or U3136 (N_3136,N_2882,N_3022);
or U3137 (N_3137,N_3020,N_3031);
or U3138 (N_3138,N_2949,N_2902);
nor U3139 (N_3139,N_2894,N_2884);
and U3140 (N_3140,N_2882,N_2991);
or U3141 (N_3141,N_2936,N_2908);
xnor U3142 (N_3142,N_2886,N_2893);
nor U3143 (N_3143,N_2974,N_3009);
nand U3144 (N_3144,N_2898,N_2941);
nor U3145 (N_3145,N_2904,N_3029);
nor U3146 (N_3146,N_2908,N_3024);
nor U3147 (N_3147,N_3034,N_2999);
nand U3148 (N_3148,N_2971,N_2936);
nand U3149 (N_3149,N_2898,N_2964);
nor U3150 (N_3150,N_2986,N_2934);
nand U3151 (N_3151,N_2947,N_2972);
nor U3152 (N_3152,N_2984,N_2961);
and U3153 (N_3153,N_2992,N_2950);
nor U3154 (N_3154,N_2998,N_2894);
and U3155 (N_3155,N_3029,N_2935);
nor U3156 (N_3156,N_2930,N_2939);
and U3157 (N_3157,N_2989,N_3002);
nand U3158 (N_3158,N_2959,N_3020);
and U3159 (N_3159,N_3016,N_3037);
nand U3160 (N_3160,N_2936,N_2942);
or U3161 (N_3161,N_2997,N_2903);
or U3162 (N_3162,N_3023,N_3017);
nand U3163 (N_3163,N_3034,N_2904);
xor U3164 (N_3164,N_3000,N_2979);
nand U3165 (N_3165,N_2909,N_2980);
xnor U3166 (N_3166,N_2886,N_2995);
nor U3167 (N_3167,N_2969,N_3012);
nand U3168 (N_3168,N_2885,N_2976);
xnor U3169 (N_3169,N_2999,N_3014);
or U3170 (N_3170,N_2983,N_3030);
nor U3171 (N_3171,N_2908,N_2943);
nand U3172 (N_3172,N_2994,N_3004);
nor U3173 (N_3173,N_3008,N_2887);
xnor U3174 (N_3174,N_3015,N_2999);
nor U3175 (N_3175,N_2979,N_2888);
nor U3176 (N_3176,N_2993,N_3018);
nor U3177 (N_3177,N_2947,N_3029);
or U3178 (N_3178,N_2979,N_2913);
nand U3179 (N_3179,N_2942,N_2912);
nor U3180 (N_3180,N_2916,N_2948);
or U3181 (N_3181,N_2919,N_2926);
and U3182 (N_3182,N_3039,N_2970);
nand U3183 (N_3183,N_2901,N_2970);
xnor U3184 (N_3184,N_3026,N_2933);
nor U3185 (N_3185,N_3027,N_2947);
nor U3186 (N_3186,N_2974,N_2957);
nand U3187 (N_3187,N_2911,N_2956);
and U3188 (N_3188,N_2910,N_3022);
and U3189 (N_3189,N_2988,N_3011);
nor U3190 (N_3190,N_3015,N_2955);
xor U3191 (N_3191,N_3007,N_2919);
nor U3192 (N_3192,N_3032,N_2905);
xnor U3193 (N_3193,N_2943,N_2880);
xnor U3194 (N_3194,N_2954,N_3009);
nor U3195 (N_3195,N_2894,N_2917);
nor U3196 (N_3196,N_2902,N_2946);
or U3197 (N_3197,N_2951,N_2984);
nor U3198 (N_3198,N_2941,N_2922);
nand U3199 (N_3199,N_3016,N_2962);
nor U3200 (N_3200,N_3092,N_3090);
or U3201 (N_3201,N_3070,N_3048);
and U3202 (N_3202,N_3082,N_3069);
xnor U3203 (N_3203,N_3189,N_3076);
or U3204 (N_3204,N_3176,N_3079);
and U3205 (N_3205,N_3100,N_3058);
nand U3206 (N_3206,N_3049,N_3199);
xor U3207 (N_3207,N_3195,N_3112);
nor U3208 (N_3208,N_3173,N_3053);
or U3209 (N_3209,N_3085,N_3144);
and U3210 (N_3210,N_3096,N_3143);
and U3211 (N_3211,N_3141,N_3057);
or U3212 (N_3212,N_3073,N_3045);
xor U3213 (N_3213,N_3177,N_3043);
xor U3214 (N_3214,N_3044,N_3062);
nand U3215 (N_3215,N_3148,N_3155);
xor U3216 (N_3216,N_3198,N_3135);
or U3217 (N_3217,N_3133,N_3113);
nand U3218 (N_3218,N_3153,N_3160);
xor U3219 (N_3219,N_3136,N_3137);
xor U3220 (N_3220,N_3121,N_3061);
and U3221 (N_3221,N_3168,N_3186);
nand U3222 (N_3222,N_3099,N_3146);
nor U3223 (N_3223,N_3064,N_3193);
or U3224 (N_3224,N_3041,N_3169);
and U3225 (N_3225,N_3180,N_3042);
xor U3226 (N_3226,N_3179,N_3184);
or U3227 (N_3227,N_3107,N_3131);
or U3228 (N_3228,N_3157,N_3110);
or U3229 (N_3229,N_3103,N_3151);
and U3230 (N_3230,N_3194,N_3119);
or U3231 (N_3231,N_3139,N_3167);
or U3232 (N_3232,N_3094,N_3123);
and U3233 (N_3233,N_3166,N_3165);
nor U3234 (N_3234,N_3175,N_3040);
xnor U3235 (N_3235,N_3056,N_3197);
nor U3236 (N_3236,N_3074,N_3125);
nor U3237 (N_3237,N_3055,N_3185);
or U3238 (N_3238,N_3117,N_3170);
nor U3239 (N_3239,N_3083,N_3126);
xnor U3240 (N_3240,N_3124,N_3052);
nand U3241 (N_3241,N_3051,N_3102);
or U3242 (N_3242,N_3068,N_3071);
nor U3243 (N_3243,N_3191,N_3187);
nand U3244 (N_3244,N_3145,N_3089);
nand U3245 (N_3245,N_3084,N_3150);
nand U3246 (N_3246,N_3159,N_3080);
xor U3247 (N_3247,N_3075,N_3129);
xor U3248 (N_3248,N_3115,N_3059);
nand U3249 (N_3249,N_3087,N_3134);
and U3250 (N_3250,N_3060,N_3178);
or U3251 (N_3251,N_3183,N_3138);
or U3252 (N_3252,N_3158,N_3086);
nand U3253 (N_3253,N_3149,N_3046);
nor U3254 (N_3254,N_3127,N_3142);
xor U3255 (N_3255,N_3174,N_3120);
or U3256 (N_3256,N_3154,N_3098);
or U3257 (N_3257,N_3181,N_3072);
nand U3258 (N_3258,N_3161,N_3182);
nand U3259 (N_3259,N_3114,N_3140);
nand U3260 (N_3260,N_3130,N_3077);
and U3261 (N_3261,N_3152,N_3108);
or U3262 (N_3262,N_3081,N_3047);
nor U3263 (N_3263,N_3192,N_3162);
and U3264 (N_3264,N_3196,N_3097);
or U3265 (N_3265,N_3093,N_3109);
and U3266 (N_3266,N_3122,N_3132);
or U3267 (N_3267,N_3106,N_3147);
and U3268 (N_3268,N_3091,N_3156);
and U3269 (N_3269,N_3050,N_3172);
or U3270 (N_3270,N_3095,N_3088);
nor U3271 (N_3271,N_3171,N_3067);
and U3272 (N_3272,N_3190,N_3118);
nor U3273 (N_3273,N_3101,N_3065);
xnor U3274 (N_3274,N_3078,N_3063);
nand U3275 (N_3275,N_3105,N_3163);
or U3276 (N_3276,N_3066,N_3054);
and U3277 (N_3277,N_3128,N_3188);
nor U3278 (N_3278,N_3164,N_3116);
nor U3279 (N_3279,N_3111,N_3104);
and U3280 (N_3280,N_3111,N_3083);
nand U3281 (N_3281,N_3120,N_3086);
or U3282 (N_3282,N_3189,N_3185);
xor U3283 (N_3283,N_3111,N_3143);
xor U3284 (N_3284,N_3071,N_3163);
or U3285 (N_3285,N_3099,N_3138);
nand U3286 (N_3286,N_3118,N_3081);
nand U3287 (N_3287,N_3092,N_3111);
nor U3288 (N_3288,N_3128,N_3097);
or U3289 (N_3289,N_3076,N_3134);
nor U3290 (N_3290,N_3042,N_3076);
xnor U3291 (N_3291,N_3128,N_3167);
nand U3292 (N_3292,N_3074,N_3196);
xnor U3293 (N_3293,N_3075,N_3081);
nand U3294 (N_3294,N_3197,N_3129);
xor U3295 (N_3295,N_3085,N_3127);
nor U3296 (N_3296,N_3185,N_3176);
nor U3297 (N_3297,N_3190,N_3054);
and U3298 (N_3298,N_3065,N_3150);
xnor U3299 (N_3299,N_3185,N_3104);
or U3300 (N_3300,N_3071,N_3186);
nor U3301 (N_3301,N_3125,N_3164);
or U3302 (N_3302,N_3158,N_3143);
nor U3303 (N_3303,N_3134,N_3103);
or U3304 (N_3304,N_3189,N_3087);
nand U3305 (N_3305,N_3192,N_3116);
or U3306 (N_3306,N_3191,N_3062);
nand U3307 (N_3307,N_3176,N_3063);
nor U3308 (N_3308,N_3147,N_3067);
or U3309 (N_3309,N_3042,N_3169);
or U3310 (N_3310,N_3063,N_3040);
nand U3311 (N_3311,N_3124,N_3048);
nand U3312 (N_3312,N_3078,N_3164);
or U3313 (N_3313,N_3130,N_3125);
xnor U3314 (N_3314,N_3045,N_3065);
nand U3315 (N_3315,N_3172,N_3145);
and U3316 (N_3316,N_3115,N_3109);
xnor U3317 (N_3317,N_3156,N_3131);
xnor U3318 (N_3318,N_3081,N_3096);
or U3319 (N_3319,N_3153,N_3148);
xnor U3320 (N_3320,N_3054,N_3168);
and U3321 (N_3321,N_3086,N_3092);
and U3322 (N_3322,N_3168,N_3093);
nand U3323 (N_3323,N_3132,N_3068);
and U3324 (N_3324,N_3040,N_3110);
or U3325 (N_3325,N_3049,N_3068);
nor U3326 (N_3326,N_3146,N_3110);
and U3327 (N_3327,N_3080,N_3087);
or U3328 (N_3328,N_3074,N_3069);
xor U3329 (N_3329,N_3106,N_3064);
nand U3330 (N_3330,N_3061,N_3042);
and U3331 (N_3331,N_3116,N_3085);
or U3332 (N_3332,N_3048,N_3187);
or U3333 (N_3333,N_3148,N_3126);
and U3334 (N_3334,N_3133,N_3145);
xnor U3335 (N_3335,N_3160,N_3079);
xor U3336 (N_3336,N_3135,N_3137);
or U3337 (N_3337,N_3132,N_3115);
or U3338 (N_3338,N_3113,N_3088);
or U3339 (N_3339,N_3076,N_3184);
or U3340 (N_3340,N_3166,N_3133);
nand U3341 (N_3341,N_3186,N_3109);
xor U3342 (N_3342,N_3091,N_3067);
nor U3343 (N_3343,N_3101,N_3053);
xor U3344 (N_3344,N_3109,N_3108);
nand U3345 (N_3345,N_3185,N_3048);
and U3346 (N_3346,N_3114,N_3166);
nand U3347 (N_3347,N_3108,N_3073);
or U3348 (N_3348,N_3103,N_3198);
and U3349 (N_3349,N_3192,N_3143);
xor U3350 (N_3350,N_3095,N_3148);
xor U3351 (N_3351,N_3050,N_3101);
nand U3352 (N_3352,N_3154,N_3127);
and U3353 (N_3353,N_3101,N_3051);
nor U3354 (N_3354,N_3099,N_3066);
and U3355 (N_3355,N_3175,N_3195);
and U3356 (N_3356,N_3145,N_3162);
nand U3357 (N_3357,N_3052,N_3144);
xnor U3358 (N_3358,N_3161,N_3088);
xnor U3359 (N_3359,N_3096,N_3108);
or U3360 (N_3360,N_3274,N_3262);
and U3361 (N_3361,N_3242,N_3215);
xor U3362 (N_3362,N_3270,N_3205);
xnor U3363 (N_3363,N_3326,N_3206);
xor U3364 (N_3364,N_3298,N_3288);
nor U3365 (N_3365,N_3345,N_3208);
nand U3366 (N_3366,N_3325,N_3289);
nand U3367 (N_3367,N_3244,N_3328);
or U3368 (N_3368,N_3229,N_3341);
and U3369 (N_3369,N_3306,N_3304);
nor U3370 (N_3370,N_3269,N_3234);
xnor U3371 (N_3371,N_3231,N_3210);
xnor U3372 (N_3372,N_3209,N_3250);
nand U3373 (N_3373,N_3287,N_3236);
or U3374 (N_3374,N_3204,N_3358);
nor U3375 (N_3375,N_3214,N_3347);
nor U3376 (N_3376,N_3272,N_3299);
nand U3377 (N_3377,N_3310,N_3320);
nand U3378 (N_3378,N_3279,N_3213);
nand U3379 (N_3379,N_3337,N_3200);
or U3380 (N_3380,N_3255,N_3240);
nand U3381 (N_3381,N_3252,N_3261);
and U3382 (N_3382,N_3280,N_3251);
or U3383 (N_3383,N_3227,N_3247);
nand U3384 (N_3384,N_3327,N_3336);
and U3385 (N_3385,N_3237,N_3260);
or U3386 (N_3386,N_3254,N_3258);
nand U3387 (N_3387,N_3245,N_3217);
or U3388 (N_3388,N_3228,N_3201);
or U3389 (N_3389,N_3256,N_3330);
or U3390 (N_3390,N_3267,N_3243);
and U3391 (N_3391,N_3333,N_3313);
xnor U3392 (N_3392,N_3257,N_3216);
and U3393 (N_3393,N_3351,N_3221);
nor U3394 (N_3394,N_3321,N_3305);
and U3395 (N_3395,N_3334,N_3344);
xnor U3396 (N_3396,N_3284,N_3357);
or U3397 (N_3397,N_3352,N_3285);
and U3398 (N_3398,N_3293,N_3349);
nor U3399 (N_3399,N_3230,N_3212);
or U3400 (N_3400,N_3248,N_3238);
and U3401 (N_3401,N_3290,N_3219);
and U3402 (N_3402,N_3259,N_3355);
xor U3403 (N_3403,N_3241,N_3202);
xor U3404 (N_3404,N_3253,N_3331);
or U3405 (N_3405,N_3207,N_3233);
and U3406 (N_3406,N_3323,N_3307);
xnor U3407 (N_3407,N_3335,N_3222);
xnor U3408 (N_3408,N_3343,N_3291);
xnor U3409 (N_3409,N_3312,N_3356);
nand U3410 (N_3410,N_3308,N_3218);
or U3411 (N_3411,N_3354,N_3268);
or U3412 (N_3412,N_3235,N_3311);
nor U3413 (N_3413,N_3295,N_3294);
xor U3414 (N_3414,N_3232,N_3353);
xor U3415 (N_3415,N_3332,N_3338);
xnor U3416 (N_3416,N_3265,N_3342);
xor U3417 (N_3417,N_3226,N_3246);
nor U3418 (N_3418,N_3281,N_3224);
xnor U3419 (N_3419,N_3275,N_3220);
nor U3420 (N_3420,N_3264,N_3322);
xor U3421 (N_3421,N_3225,N_3346);
or U3422 (N_3422,N_3278,N_3314);
or U3423 (N_3423,N_3292,N_3211);
nor U3424 (N_3424,N_3283,N_3301);
and U3425 (N_3425,N_3329,N_3223);
nor U3426 (N_3426,N_3324,N_3339);
nand U3427 (N_3427,N_3303,N_3203);
nor U3428 (N_3428,N_3315,N_3249);
xnor U3429 (N_3429,N_3340,N_3239);
xor U3430 (N_3430,N_3359,N_3297);
and U3431 (N_3431,N_3302,N_3263);
and U3432 (N_3432,N_3296,N_3319);
or U3433 (N_3433,N_3266,N_3271);
nand U3434 (N_3434,N_3316,N_3277);
nand U3435 (N_3435,N_3348,N_3286);
xnor U3436 (N_3436,N_3317,N_3273);
xor U3437 (N_3437,N_3282,N_3300);
nor U3438 (N_3438,N_3350,N_3309);
xnor U3439 (N_3439,N_3318,N_3276);
and U3440 (N_3440,N_3253,N_3355);
or U3441 (N_3441,N_3241,N_3274);
and U3442 (N_3442,N_3330,N_3283);
and U3443 (N_3443,N_3300,N_3342);
and U3444 (N_3444,N_3352,N_3280);
and U3445 (N_3445,N_3289,N_3294);
and U3446 (N_3446,N_3243,N_3296);
and U3447 (N_3447,N_3317,N_3262);
nor U3448 (N_3448,N_3213,N_3352);
nand U3449 (N_3449,N_3331,N_3200);
or U3450 (N_3450,N_3346,N_3253);
xnor U3451 (N_3451,N_3245,N_3281);
and U3452 (N_3452,N_3311,N_3286);
xnor U3453 (N_3453,N_3278,N_3225);
nand U3454 (N_3454,N_3269,N_3311);
nor U3455 (N_3455,N_3328,N_3246);
nor U3456 (N_3456,N_3292,N_3228);
and U3457 (N_3457,N_3330,N_3246);
and U3458 (N_3458,N_3351,N_3339);
nor U3459 (N_3459,N_3281,N_3257);
nand U3460 (N_3460,N_3308,N_3347);
or U3461 (N_3461,N_3354,N_3264);
and U3462 (N_3462,N_3298,N_3348);
nor U3463 (N_3463,N_3218,N_3299);
xor U3464 (N_3464,N_3228,N_3338);
nor U3465 (N_3465,N_3309,N_3230);
or U3466 (N_3466,N_3212,N_3207);
and U3467 (N_3467,N_3208,N_3299);
nand U3468 (N_3468,N_3226,N_3266);
or U3469 (N_3469,N_3242,N_3323);
xor U3470 (N_3470,N_3274,N_3286);
xnor U3471 (N_3471,N_3282,N_3321);
xor U3472 (N_3472,N_3343,N_3334);
xor U3473 (N_3473,N_3317,N_3238);
xor U3474 (N_3474,N_3310,N_3256);
or U3475 (N_3475,N_3237,N_3292);
xnor U3476 (N_3476,N_3244,N_3268);
and U3477 (N_3477,N_3226,N_3249);
nand U3478 (N_3478,N_3308,N_3257);
nor U3479 (N_3479,N_3305,N_3276);
nor U3480 (N_3480,N_3318,N_3311);
or U3481 (N_3481,N_3332,N_3317);
or U3482 (N_3482,N_3204,N_3286);
xor U3483 (N_3483,N_3351,N_3220);
nand U3484 (N_3484,N_3334,N_3247);
xor U3485 (N_3485,N_3209,N_3276);
or U3486 (N_3486,N_3332,N_3203);
nand U3487 (N_3487,N_3218,N_3207);
nor U3488 (N_3488,N_3256,N_3295);
nand U3489 (N_3489,N_3303,N_3319);
nand U3490 (N_3490,N_3240,N_3266);
nor U3491 (N_3491,N_3302,N_3331);
or U3492 (N_3492,N_3201,N_3354);
nand U3493 (N_3493,N_3345,N_3254);
nor U3494 (N_3494,N_3317,N_3328);
xnor U3495 (N_3495,N_3258,N_3333);
xnor U3496 (N_3496,N_3252,N_3325);
and U3497 (N_3497,N_3215,N_3219);
xnor U3498 (N_3498,N_3326,N_3315);
xnor U3499 (N_3499,N_3333,N_3348);
nand U3500 (N_3500,N_3256,N_3216);
or U3501 (N_3501,N_3358,N_3276);
nand U3502 (N_3502,N_3201,N_3208);
nor U3503 (N_3503,N_3315,N_3244);
xor U3504 (N_3504,N_3296,N_3331);
or U3505 (N_3505,N_3245,N_3219);
nor U3506 (N_3506,N_3353,N_3266);
or U3507 (N_3507,N_3320,N_3237);
nand U3508 (N_3508,N_3216,N_3309);
nor U3509 (N_3509,N_3321,N_3232);
and U3510 (N_3510,N_3215,N_3246);
xnor U3511 (N_3511,N_3265,N_3300);
xnor U3512 (N_3512,N_3337,N_3272);
or U3513 (N_3513,N_3289,N_3261);
nor U3514 (N_3514,N_3250,N_3308);
or U3515 (N_3515,N_3293,N_3236);
nor U3516 (N_3516,N_3314,N_3227);
nand U3517 (N_3517,N_3235,N_3337);
nand U3518 (N_3518,N_3301,N_3203);
or U3519 (N_3519,N_3254,N_3311);
and U3520 (N_3520,N_3478,N_3507);
or U3521 (N_3521,N_3495,N_3406);
xor U3522 (N_3522,N_3421,N_3405);
nor U3523 (N_3523,N_3415,N_3445);
or U3524 (N_3524,N_3385,N_3463);
or U3525 (N_3525,N_3513,N_3437);
or U3526 (N_3526,N_3381,N_3432);
or U3527 (N_3527,N_3461,N_3470);
or U3528 (N_3528,N_3387,N_3492);
and U3529 (N_3529,N_3430,N_3364);
nand U3530 (N_3530,N_3429,N_3498);
or U3531 (N_3531,N_3469,N_3420);
and U3532 (N_3532,N_3365,N_3441);
or U3533 (N_3533,N_3378,N_3383);
nor U3534 (N_3534,N_3386,N_3447);
nor U3535 (N_3535,N_3403,N_3511);
nand U3536 (N_3536,N_3453,N_3512);
xnor U3537 (N_3537,N_3502,N_3506);
or U3538 (N_3538,N_3419,N_3484);
and U3539 (N_3539,N_3368,N_3393);
nand U3540 (N_3540,N_3398,N_3481);
and U3541 (N_3541,N_3457,N_3414);
and U3542 (N_3542,N_3450,N_3496);
nor U3543 (N_3543,N_3372,N_3407);
and U3544 (N_3544,N_3515,N_3411);
xnor U3545 (N_3545,N_3514,N_3443);
xor U3546 (N_3546,N_3412,N_3377);
xnor U3547 (N_3547,N_3487,N_3367);
and U3548 (N_3548,N_3362,N_3452);
nand U3549 (N_3549,N_3459,N_3360);
xor U3550 (N_3550,N_3425,N_3435);
or U3551 (N_3551,N_3401,N_3392);
nor U3552 (N_3552,N_3371,N_3423);
xnor U3553 (N_3553,N_3493,N_3490);
nor U3554 (N_3554,N_3460,N_3446);
nor U3555 (N_3555,N_3509,N_3501);
nor U3556 (N_3556,N_3465,N_3455);
nand U3557 (N_3557,N_3369,N_3456);
nand U3558 (N_3558,N_3382,N_3510);
nor U3559 (N_3559,N_3380,N_3436);
nor U3560 (N_3560,N_3384,N_3438);
nand U3561 (N_3561,N_3427,N_3444);
xnor U3562 (N_3562,N_3418,N_3395);
or U3563 (N_3563,N_3479,N_3413);
nor U3564 (N_3564,N_3467,N_3394);
nand U3565 (N_3565,N_3426,N_3476);
or U3566 (N_3566,N_3466,N_3416);
nand U3567 (N_3567,N_3431,N_3397);
nor U3568 (N_3568,N_3388,N_3374);
xor U3569 (N_3569,N_3500,N_3424);
nand U3570 (N_3570,N_3464,N_3508);
or U3571 (N_3571,N_3486,N_3376);
or U3572 (N_3572,N_3503,N_3442);
nand U3573 (N_3573,N_3370,N_3483);
and U3574 (N_3574,N_3391,N_3399);
and U3575 (N_3575,N_3390,N_3462);
nor U3576 (N_3576,N_3499,N_3458);
nor U3577 (N_3577,N_3410,N_3477);
or U3578 (N_3578,N_3428,N_3475);
and U3579 (N_3579,N_3408,N_3491);
nand U3580 (N_3580,N_3375,N_3404);
nor U3581 (N_3581,N_3505,N_3389);
xnor U3582 (N_3582,N_3449,N_3474);
nor U3583 (N_3583,N_3454,N_3472);
nor U3584 (N_3584,N_3366,N_3489);
nor U3585 (N_3585,N_3516,N_3400);
or U3586 (N_3586,N_3504,N_3480);
and U3587 (N_3587,N_3361,N_3451);
nand U3588 (N_3588,N_3471,N_3440);
nand U3589 (N_3589,N_3422,N_3519);
nor U3590 (N_3590,N_3482,N_3517);
and U3591 (N_3591,N_3494,N_3434);
and U3592 (N_3592,N_3396,N_3468);
xor U3593 (N_3593,N_3488,N_3439);
and U3594 (N_3594,N_3497,N_3485);
and U3595 (N_3595,N_3409,N_3373);
nor U3596 (N_3596,N_3402,N_3379);
xor U3597 (N_3597,N_3448,N_3518);
nor U3598 (N_3598,N_3417,N_3473);
or U3599 (N_3599,N_3363,N_3433);
nor U3600 (N_3600,N_3417,N_3364);
or U3601 (N_3601,N_3377,N_3493);
and U3602 (N_3602,N_3507,N_3411);
and U3603 (N_3603,N_3376,N_3439);
nand U3604 (N_3604,N_3371,N_3452);
xnor U3605 (N_3605,N_3514,N_3395);
or U3606 (N_3606,N_3442,N_3378);
and U3607 (N_3607,N_3466,N_3461);
or U3608 (N_3608,N_3465,N_3400);
and U3609 (N_3609,N_3426,N_3381);
nand U3610 (N_3610,N_3361,N_3479);
nand U3611 (N_3611,N_3486,N_3514);
nand U3612 (N_3612,N_3361,N_3385);
nand U3613 (N_3613,N_3466,N_3413);
and U3614 (N_3614,N_3506,N_3393);
nor U3615 (N_3615,N_3381,N_3445);
or U3616 (N_3616,N_3472,N_3413);
or U3617 (N_3617,N_3463,N_3464);
nand U3618 (N_3618,N_3498,N_3388);
and U3619 (N_3619,N_3473,N_3448);
nand U3620 (N_3620,N_3364,N_3420);
xor U3621 (N_3621,N_3472,N_3471);
or U3622 (N_3622,N_3362,N_3430);
and U3623 (N_3623,N_3445,N_3397);
nand U3624 (N_3624,N_3443,N_3481);
and U3625 (N_3625,N_3508,N_3496);
or U3626 (N_3626,N_3480,N_3508);
xnor U3627 (N_3627,N_3413,N_3451);
nor U3628 (N_3628,N_3498,N_3438);
and U3629 (N_3629,N_3408,N_3479);
and U3630 (N_3630,N_3459,N_3519);
nor U3631 (N_3631,N_3406,N_3391);
or U3632 (N_3632,N_3426,N_3398);
nand U3633 (N_3633,N_3439,N_3459);
nor U3634 (N_3634,N_3401,N_3403);
nor U3635 (N_3635,N_3463,N_3440);
nor U3636 (N_3636,N_3488,N_3400);
nand U3637 (N_3637,N_3418,N_3460);
or U3638 (N_3638,N_3465,N_3391);
or U3639 (N_3639,N_3428,N_3441);
xnor U3640 (N_3640,N_3410,N_3476);
or U3641 (N_3641,N_3368,N_3372);
and U3642 (N_3642,N_3363,N_3465);
nor U3643 (N_3643,N_3435,N_3513);
and U3644 (N_3644,N_3457,N_3490);
xor U3645 (N_3645,N_3449,N_3378);
nand U3646 (N_3646,N_3508,N_3366);
nor U3647 (N_3647,N_3471,N_3370);
and U3648 (N_3648,N_3450,N_3429);
nand U3649 (N_3649,N_3399,N_3361);
and U3650 (N_3650,N_3498,N_3389);
nor U3651 (N_3651,N_3460,N_3407);
xor U3652 (N_3652,N_3475,N_3445);
nor U3653 (N_3653,N_3494,N_3396);
nor U3654 (N_3654,N_3498,N_3448);
nor U3655 (N_3655,N_3405,N_3513);
nand U3656 (N_3656,N_3421,N_3461);
or U3657 (N_3657,N_3503,N_3516);
xnor U3658 (N_3658,N_3367,N_3420);
nor U3659 (N_3659,N_3460,N_3432);
and U3660 (N_3660,N_3400,N_3389);
nand U3661 (N_3661,N_3397,N_3394);
or U3662 (N_3662,N_3400,N_3421);
and U3663 (N_3663,N_3400,N_3483);
xor U3664 (N_3664,N_3465,N_3498);
or U3665 (N_3665,N_3508,N_3503);
nand U3666 (N_3666,N_3510,N_3363);
and U3667 (N_3667,N_3387,N_3460);
and U3668 (N_3668,N_3515,N_3381);
and U3669 (N_3669,N_3459,N_3431);
and U3670 (N_3670,N_3390,N_3362);
or U3671 (N_3671,N_3375,N_3372);
nand U3672 (N_3672,N_3515,N_3364);
nand U3673 (N_3673,N_3496,N_3444);
and U3674 (N_3674,N_3391,N_3364);
xor U3675 (N_3675,N_3439,N_3461);
nand U3676 (N_3676,N_3408,N_3374);
and U3677 (N_3677,N_3491,N_3392);
or U3678 (N_3678,N_3459,N_3449);
and U3679 (N_3679,N_3371,N_3394);
or U3680 (N_3680,N_3662,N_3623);
nor U3681 (N_3681,N_3608,N_3655);
nor U3682 (N_3682,N_3544,N_3600);
and U3683 (N_3683,N_3624,N_3556);
xor U3684 (N_3684,N_3589,N_3574);
or U3685 (N_3685,N_3529,N_3644);
nand U3686 (N_3686,N_3599,N_3635);
or U3687 (N_3687,N_3648,N_3679);
and U3688 (N_3688,N_3523,N_3546);
nor U3689 (N_3689,N_3560,N_3654);
or U3690 (N_3690,N_3548,N_3643);
xnor U3691 (N_3691,N_3580,N_3549);
or U3692 (N_3692,N_3611,N_3629);
nor U3693 (N_3693,N_3627,N_3524);
or U3694 (N_3694,N_3617,N_3551);
and U3695 (N_3695,N_3664,N_3613);
xnor U3696 (N_3696,N_3647,N_3552);
nor U3697 (N_3697,N_3542,N_3590);
or U3698 (N_3698,N_3669,N_3642);
or U3699 (N_3699,N_3625,N_3597);
nand U3700 (N_3700,N_3676,N_3576);
nand U3701 (N_3701,N_3603,N_3573);
or U3702 (N_3702,N_3615,N_3567);
or U3703 (N_3703,N_3530,N_3569);
nand U3704 (N_3704,N_3527,N_3536);
nand U3705 (N_3705,N_3656,N_3657);
nand U3706 (N_3706,N_3673,N_3564);
nor U3707 (N_3707,N_3637,N_3604);
or U3708 (N_3708,N_3652,N_3561);
nor U3709 (N_3709,N_3666,N_3612);
and U3710 (N_3710,N_3582,N_3521);
nand U3711 (N_3711,N_3593,N_3631);
or U3712 (N_3712,N_3663,N_3658);
or U3713 (N_3713,N_3607,N_3675);
and U3714 (N_3714,N_3609,N_3636);
nand U3715 (N_3715,N_3558,N_3539);
nand U3716 (N_3716,N_3661,N_3670);
nand U3717 (N_3717,N_3667,N_3565);
or U3718 (N_3718,N_3525,N_3598);
nor U3719 (N_3719,N_3614,N_3641);
or U3720 (N_3720,N_3602,N_3570);
or U3721 (N_3721,N_3659,N_3587);
xor U3722 (N_3722,N_3619,N_3550);
nand U3723 (N_3723,N_3522,N_3645);
and U3724 (N_3724,N_3665,N_3584);
nor U3725 (N_3725,N_3583,N_3630);
nor U3726 (N_3726,N_3566,N_3533);
nand U3727 (N_3727,N_3537,N_3581);
or U3728 (N_3728,N_3653,N_3639);
and U3729 (N_3729,N_3531,N_3534);
and U3730 (N_3730,N_3568,N_3575);
nor U3731 (N_3731,N_3591,N_3622);
and U3732 (N_3732,N_3660,N_3585);
nor U3733 (N_3733,N_3528,N_3606);
or U3734 (N_3734,N_3594,N_3555);
xor U3735 (N_3735,N_3601,N_3620);
xnor U3736 (N_3736,N_3541,N_3559);
xnor U3737 (N_3737,N_3571,N_3563);
nor U3738 (N_3738,N_3668,N_3632);
nor U3739 (N_3739,N_3532,N_3605);
and U3740 (N_3740,N_3595,N_3640);
and U3741 (N_3741,N_3554,N_3520);
nand U3742 (N_3742,N_3628,N_3678);
nand U3743 (N_3743,N_3535,N_3621);
and U3744 (N_3744,N_3578,N_3672);
xnor U3745 (N_3745,N_3650,N_3649);
nor U3746 (N_3746,N_3526,N_3572);
or U3747 (N_3747,N_3579,N_3547);
nand U3748 (N_3748,N_3586,N_3674);
nor U3749 (N_3749,N_3616,N_3618);
or U3750 (N_3750,N_3557,N_3626);
nand U3751 (N_3751,N_3634,N_3538);
nor U3752 (N_3752,N_3671,N_3638);
and U3753 (N_3753,N_3543,N_3540);
nand U3754 (N_3754,N_3553,N_3592);
and U3755 (N_3755,N_3677,N_3651);
nor U3756 (N_3756,N_3545,N_3588);
or U3757 (N_3757,N_3562,N_3633);
or U3758 (N_3758,N_3610,N_3577);
xor U3759 (N_3759,N_3646,N_3596);
nor U3760 (N_3760,N_3541,N_3616);
nand U3761 (N_3761,N_3568,N_3616);
xor U3762 (N_3762,N_3590,N_3527);
xnor U3763 (N_3763,N_3566,N_3652);
or U3764 (N_3764,N_3625,N_3679);
nor U3765 (N_3765,N_3574,N_3638);
xnor U3766 (N_3766,N_3672,N_3586);
nor U3767 (N_3767,N_3607,N_3610);
nand U3768 (N_3768,N_3594,N_3657);
and U3769 (N_3769,N_3557,N_3669);
and U3770 (N_3770,N_3594,N_3604);
and U3771 (N_3771,N_3610,N_3637);
xnor U3772 (N_3772,N_3588,N_3537);
nor U3773 (N_3773,N_3634,N_3621);
xor U3774 (N_3774,N_3639,N_3601);
xor U3775 (N_3775,N_3549,N_3566);
xor U3776 (N_3776,N_3599,N_3653);
nor U3777 (N_3777,N_3579,N_3616);
or U3778 (N_3778,N_3589,N_3569);
xor U3779 (N_3779,N_3626,N_3533);
and U3780 (N_3780,N_3625,N_3672);
nor U3781 (N_3781,N_3610,N_3542);
nand U3782 (N_3782,N_3641,N_3671);
nand U3783 (N_3783,N_3614,N_3552);
xor U3784 (N_3784,N_3616,N_3547);
or U3785 (N_3785,N_3527,N_3645);
nand U3786 (N_3786,N_3565,N_3587);
and U3787 (N_3787,N_3674,N_3676);
xor U3788 (N_3788,N_3582,N_3527);
or U3789 (N_3789,N_3528,N_3625);
nor U3790 (N_3790,N_3604,N_3646);
xnor U3791 (N_3791,N_3614,N_3658);
xor U3792 (N_3792,N_3655,N_3631);
or U3793 (N_3793,N_3573,N_3527);
and U3794 (N_3794,N_3588,N_3667);
xnor U3795 (N_3795,N_3546,N_3618);
and U3796 (N_3796,N_3536,N_3544);
or U3797 (N_3797,N_3617,N_3543);
xor U3798 (N_3798,N_3614,N_3629);
nand U3799 (N_3799,N_3575,N_3671);
xnor U3800 (N_3800,N_3548,N_3642);
nor U3801 (N_3801,N_3644,N_3531);
nor U3802 (N_3802,N_3644,N_3669);
nor U3803 (N_3803,N_3567,N_3595);
nand U3804 (N_3804,N_3678,N_3679);
nand U3805 (N_3805,N_3575,N_3576);
xnor U3806 (N_3806,N_3605,N_3615);
and U3807 (N_3807,N_3547,N_3679);
xnor U3808 (N_3808,N_3655,N_3622);
or U3809 (N_3809,N_3646,N_3599);
nor U3810 (N_3810,N_3547,N_3534);
nand U3811 (N_3811,N_3666,N_3543);
or U3812 (N_3812,N_3632,N_3622);
nor U3813 (N_3813,N_3545,N_3559);
nand U3814 (N_3814,N_3650,N_3571);
or U3815 (N_3815,N_3645,N_3631);
nor U3816 (N_3816,N_3553,N_3614);
nand U3817 (N_3817,N_3553,N_3618);
xnor U3818 (N_3818,N_3574,N_3648);
and U3819 (N_3819,N_3586,N_3567);
nor U3820 (N_3820,N_3656,N_3668);
and U3821 (N_3821,N_3636,N_3567);
and U3822 (N_3822,N_3619,N_3678);
nor U3823 (N_3823,N_3665,N_3667);
xnor U3824 (N_3824,N_3547,N_3602);
nor U3825 (N_3825,N_3617,N_3563);
nand U3826 (N_3826,N_3538,N_3547);
nor U3827 (N_3827,N_3543,N_3644);
xor U3828 (N_3828,N_3601,N_3525);
nand U3829 (N_3829,N_3551,N_3542);
or U3830 (N_3830,N_3674,N_3564);
or U3831 (N_3831,N_3575,N_3626);
xnor U3832 (N_3832,N_3541,N_3624);
nand U3833 (N_3833,N_3675,N_3550);
nor U3834 (N_3834,N_3605,N_3613);
nand U3835 (N_3835,N_3541,N_3531);
nand U3836 (N_3836,N_3622,N_3572);
and U3837 (N_3837,N_3665,N_3611);
nand U3838 (N_3838,N_3640,N_3543);
xnor U3839 (N_3839,N_3529,N_3597);
nand U3840 (N_3840,N_3718,N_3766);
nor U3841 (N_3841,N_3789,N_3818);
xnor U3842 (N_3842,N_3695,N_3782);
nand U3843 (N_3843,N_3781,N_3734);
xor U3844 (N_3844,N_3706,N_3836);
nand U3845 (N_3845,N_3827,N_3748);
nand U3846 (N_3846,N_3757,N_3685);
and U3847 (N_3847,N_3832,N_3773);
nor U3848 (N_3848,N_3787,N_3741);
nor U3849 (N_3849,N_3754,N_3777);
or U3850 (N_3850,N_3724,N_3687);
or U3851 (N_3851,N_3749,N_3705);
and U3852 (N_3852,N_3804,N_3716);
nor U3853 (N_3853,N_3736,N_3719);
or U3854 (N_3854,N_3830,N_3763);
xor U3855 (N_3855,N_3812,N_3732);
nand U3856 (N_3856,N_3725,N_3721);
nand U3857 (N_3857,N_3820,N_3809);
or U3858 (N_3858,N_3759,N_3765);
xor U3859 (N_3859,N_3834,N_3813);
nor U3860 (N_3860,N_3747,N_3802);
and U3861 (N_3861,N_3752,N_3703);
or U3862 (N_3862,N_3697,N_3738);
xor U3863 (N_3863,N_3701,N_3771);
xnor U3864 (N_3864,N_3710,N_3829);
or U3865 (N_3865,N_3760,N_3728);
xnor U3866 (N_3866,N_3723,N_3753);
nor U3867 (N_3867,N_3702,N_3808);
nor U3868 (N_3868,N_3735,N_3762);
nor U3869 (N_3869,N_3783,N_3810);
nand U3870 (N_3870,N_3814,N_3839);
or U3871 (N_3871,N_3713,N_3838);
xor U3872 (N_3872,N_3756,N_3796);
and U3873 (N_3873,N_3816,N_3835);
nand U3874 (N_3874,N_3704,N_3805);
and U3875 (N_3875,N_3815,N_3758);
or U3876 (N_3876,N_3731,N_3690);
nor U3877 (N_3877,N_3715,N_3730);
nor U3878 (N_3878,N_3791,N_3682);
nor U3879 (N_3879,N_3744,N_3775);
nor U3880 (N_3880,N_3683,N_3698);
nor U3881 (N_3881,N_3681,N_3691);
nor U3882 (N_3882,N_3807,N_3751);
xor U3883 (N_3883,N_3708,N_3729);
or U3884 (N_3884,N_3831,N_3764);
xnor U3885 (N_3885,N_3722,N_3699);
or U3886 (N_3886,N_3761,N_3746);
xor U3887 (N_3887,N_3711,N_3819);
or U3888 (N_3888,N_3779,N_3755);
nor U3889 (N_3889,N_3767,N_3792);
and U3890 (N_3890,N_3769,N_3720);
nor U3891 (N_3891,N_3709,N_3825);
and U3892 (N_3892,N_3811,N_3799);
xnor U3893 (N_3893,N_3837,N_3689);
nand U3894 (N_3894,N_3788,N_3717);
xor U3895 (N_3895,N_3733,N_3770);
or U3896 (N_3896,N_3774,N_3684);
nor U3897 (N_3897,N_3795,N_3712);
and U3898 (N_3898,N_3780,N_3828);
nor U3899 (N_3899,N_3822,N_3692);
xnor U3900 (N_3900,N_3785,N_3739);
nand U3901 (N_3901,N_3700,N_3806);
and U3902 (N_3902,N_3784,N_3740);
xnor U3903 (N_3903,N_3693,N_3824);
or U3904 (N_3904,N_3745,N_3694);
xor U3905 (N_3905,N_3778,N_3801);
xnor U3906 (N_3906,N_3750,N_3727);
or U3907 (N_3907,N_3817,N_3688);
and U3908 (N_3908,N_3707,N_3743);
xor U3909 (N_3909,N_3797,N_3786);
nand U3910 (N_3910,N_3686,N_3776);
xnor U3911 (N_3911,N_3772,N_3790);
nor U3912 (N_3912,N_3696,N_3826);
or U3913 (N_3913,N_3821,N_3737);
xnor U3914 (N_3914,N_3794,N_3714);
or U3915 (N_3915,N_3803,N_3823);
and U3916 (N_3916,N_3798,N_3742);
nand U3917 (N_3917,N_3800,N_3768);
nand U3918 (N_3918,N_3680,N_3726);
and U3919 (N_3919,N_3793,N_3833);
xor U3920 (N_3920,N_3728,N_3759);
nand U3921 (N_3921,N_3774,N_3693);
nor U3922 (N_3922,N_3725,N_3797);
or U3923 (N_3923,N_3806,N_3712);
nand U3924 (N_3924,N_3774,N_3826);
nand U3925 (N_3925,N_3784,N_3682);
nor U3926 (N_3926,N_3776,N_3772);
nand U3927 (N_3927,N_3837,N_3778);
or U3928 (N_3928,N_3743,N_3814);
xor U3929 (N_3929,N_3827,N_3813);
and U3930 (N_3930,N_3691,N_3718);
nand U3931 (N_3931,N_3784,N_3698);
nor U3932 (N_3932,N_3824,N_3717);
or U3933 (N_3933,N_3783,N_3780);
or U3934 (N_3934,N_3796,N_3776);
xnor U3935 (N_3935,N_3806,N_3749);
or U3936 (N_3936,N_3683,N_3739);
or U3937 (N_3937,N_3779,N_3737);
and U3938 (N_3938,N_3735,N_3746);
and U3939 (N_3939,N_3694,N_3777);
and U3940 (N_3940,N_3800,N_3739);
nor U3941 (N_3941,N_3792,N_3714);
xor U3942 (N_3942,N_3765,N_3728);
or U3943 (N_3943,N_3789,N_3741);
and U3944 (N_3944,N_3831,N_3824);
xor U3945 (N_3945,N_3759,N_3798);
nand U3946 (N_3946,N_3764,N_3779);
nor U3947 (N_3947,N_3810,N_3740);
and U3948 (N_3948,N_3725,N_3722);
nand U3949 (N_3949,N_3752,N_3727);
or U3950 (N_3950,N_3838,N_3818);
nor U3951 (N_3951,N_3716,N_3827);
nor U3952 (N_3952,N_3682,N_3831);
or U3953 (N_3953,N_3746,N_3804);
nor U3954 (N_3954,N_3754,N_3740);
xnor U3955 (N_3955,N_3792,N_3754);
nor U3956 (N_3956,N_3703,N_3809);
and U3957 (N_3957,N_3793,N_3691);
nand U3958 (N_3958,N_3729,N_3822);
or U3959 (N_3959,N_3776,N_3813);
nand U3960 (N_3960,N_3708,N_3759);
and U3961 (N_3961,N_3827,N_3719);
or U3962 (N_3962,N_3822,N_3782);
nand U3963 (N_3963,N_3804,N_3708);
and U3964 (N_3964,N_3697,N_3816);
and U3965 (N_3965,N_3811,N_3827);
nor U3966 (N_3966,N_3817,N_3729);
or U3967 (N_3967,N_3758,N_3724);
or U3968 (N_3968,N_3696,N_3774);
or U3969 (N_3969,N_3707,N_3773);
nor U3970 (N_3970,N_3748,N_3735);
nand U3971 (N_3971,N_3747,N_3832);
or U3972 (N_3972,N_3744,N_3788);
nor U3973 (N_3973,N_3774,N_3708);
and U3974 (N_3974,N_3829,N_3760);
xor U3975 (N_3975,N_3734,N_3763);
or U3976 (N_3976,N_3761,N_3684);
xor U3977 (N_3977,N_3733,N_3784);
and U3978 (N_3978,N_3694,N_3720);
xnor U3979 (N_3979,N_3811,N_3814);
nor U3980 (N_3980,N_3712,N_3731);
and U3981 (N_3981,N_3692,N_3726);
or U3982 (N_3982,N_3774,N_3789);
and U3983 (N_3983,N_3779,N_3723);
nor U3984 (N_3984,N_3754,N_3761);
nand U3985 (N_3985,N_3824,N_3838);
nor U3986 (N_3986,N_3835,N_3755);
nor U3987 (N_3987,N_3744,N_3684);
and U3988 (N_3988,N_3707,N_3765);
nand U3989 (N_3989,N_3777,N_3722);
or U3990 (N_3990,N_3692,N_3762);
nor U3991 (N_3991,N_3754,N_3772);
nand U3992 (N_3992,N_3710,N_3757);
nor U3993 (N_3993,N_3787,N_3811);
xnor U3994 (N_3994,N_3721,N_3802);
nand U3995 (N_3995,N_3697,N_3700);
nand U3996 (N_3996,N_3732,N_3757);
nor U3997 (N_3997,N_3724,N_3707);
or U3998 (N_3998,N_3732,N_3818);
and U3999 (N_3999,N_3817,N_3712);
and U4000 (N_4000,N_3916,N_3951);
or U4001 (N_4001,N_3998,N_3943);
and U4002 (N_4002,N_3979,N_3978);
nor U4003 (N_4003,N_3846,N_3920);
nor U4004 (N_4004,N_3992,N_3947);
or U4005 (N_4005,N_3880,N_3878);
xnor U4006 (N_4006,N_3892,N_3996);
or U4007 (N_4007,N_3926,N_3952);
or U4008 (N_4008,N_3965,N_3852);
and U4009 (N_4009,N_3844,N_3898);
nor U4010 (N_4010,N_3909,N_3985);
xnor U4011 (N_4011,N_3882,N_3956);
or U4012 (N_4012,N_3934,N_3859);
nor U4013 (N_4013,N_3912,N_3966);
or U4014 (N_4014,N_3913,N_3935);
or U4015 (N_4015,N_3967,N_3850);
nor U4016 (N_4016,N_3915,N_3964);
and U4017 (N_4017,N_3946,N_3847);
nand U4018 (N_4018,N_3928,N_3984);
and U4019 (N_4019,N_3879,N_3875);
and U4020 (N_4020,N_3988,N_3886);
nor U4021 (N_4021,N_3872,N_3867);
or U4022 (N_4022,N_3910,N_3974);
or U4023 (N_4023,N_3942,N_3927);
nor U4024 (N_4024,N_3884,N_3969);
xnor U4025 (N_4025,N_3895,N_3911);
and U4026 (N_4026,N_3863,N_3907);
nor U4027 (N_4027,N_3995,N_3976);
and U4028 (N_4028,N_3970,N_3871);
xor U4029 (N_4029,N_3873,N_3857);
nor U4030 (N_4030,N_3930,N_3991);
or U4031 (N_4031,N_3937,N_3861);
nand U4032 (N_4032,N_3963,N_3987);
xnor U4033 (N_4033,N_3868,N_3849);
nor U4034 (N_4034,N_3941,N_3982);
or U4035 (N_4035,N_3960,N_3989);
nor U4036 (N_4036,N_3874,N_3948);
or U4037 (N_4037,N_3864,N_3855);
and U4038 (N_4038,N_3841,N_3940);
nor U4039 (N_4039,N_3918,N_3980);
nand U4040 (N_4040,N_3923,N_3914);
xor U4041 (N_4041,N_3962,N_3896);
or U4042 (N_4042,N_3902,N_3845);
nor U4043 (N_4043,N_3993,N_3881);
and U4044 (N_4044,N_3939,N_3854);
or U4045 (N_4045,N_3889,N_3853);
and U4046 (N_4046,N_3919,N_3953);
and U4047 (N_4047,N_3973,N_3929);
or U4048 (N_4048,N_3840,N_3860);
or U4049 (N_4049,N_3869,N_3950);
and U4050 (N_4050,N_3894,N_3885);
nor U4051 (N_4051,N_3891,N_3958);
xnor U4052 (N_4052,N_3944,N_3971);
xor U4053 (N_4053,N_3917,N_3975);
or U4054 (N_4054,N_3904,N_3924);
and U4055 (N_4055,N_3877,N_3968);
xnor U4056 (N_4056,N_3870,N_3908);
nor U4057 (N_4057,N_3931,N_3899);
or U4058 (N_4058,N_3945,N_3938);
or U4059 (N_4059,N_3990,N_3851);
xnor U4060 (N_4060,N_3949,N_3997);
nand U4061 (N_4061,N_3876,N_3994);
nand U4062 (N_4062,N_3848,N_3866);
xnor U4063 (N_4063,N_3954,N_3883);
and U4064 (N_4064,N_3862,N_3900);
and U4065 (N_4065,N_3893,N_3981);
nor U4066 (N_4066,N_3977,N_3983);
and U4067 (N_4067,N_3887,N_3905);
nor U4068 (N_4068,N_3842,N_3906);
xor U4069 (N_4069,N_3890,N_3999);
or U4070 (N_4070,N_3961,N_3925);
and U4071 (N_4071,N_3856,N_3933);
xnor U4072 (N_4072,N_3955,N_3843);
nor U4073 (N_4073,N_3932,N_3957);
nor U4074 (N_4074,N_3922,N_3897);
nor U4075 (N_4075,N_3865,N_3986);
or U4076 (N_4076,N_3903,N_3888);
xor U4077 (N_4077,N_3936,N_3959);
xor U4078 (N_4078,N_3921,N_3858);
nor U4079 (N_4079,N_3972,N_3901);
nor U4080 (N_4080,N_3920,N_3945);
nor U4081 (N_4081,N_3988,N_3936);
or U4082 (N_4082,N_3988,N_3876);
nor U4083 (N_4083,N_3965,N_3997);
xor U4084 (N_4084,N_3844,N_3965);
or U4085 (N_4085,N_3984,N_3895);
and U4086 (N_4086,N_3910,N_3842);
xor U4087 (N_4087,N_3879,N_3885);
or U4088 (N_4088,N_3892,N_3866);
nor U4089 (N_4089,N_3842,N_3965);
xnor U4090 (N_4090,N_3951,N_3850);
or U4091 (N_4091,N_3935,N_3969);
nor U4092 (N_4092,N_3954,N_3841);
or U4093 (N_4093,N_3993,N_3842);
xnor U4094 (N_4094,N_3943,N_3950);
or U4095 (N_4095,N_3976,N_3953);
xnor U4096 (N_4096,N_3998,N_3872);
or U4097 (N_4097,N_3914,N_3948);
nand U4098 (N_4098,N_3898,N_3911);
nor U4099 (N_4099,N_3957,N_3940);
nand U4100 (N_4100,N_3923,N_3891);
nand U4101 (N_4101,N_3930,N_3922);
or U4102 (N_4102,N_3971,N_3995);
nand U4103 (N_4103,N_3843,N_3990);
or U4104 (N_4104,N_3957,N_3974);
xor U4105 (N_4105,N_3861,N_3878);
nand U4106 (N_4106,N_3971,N_3887);
nand U4107 (N_4107,N_3962,N_3909);
xnor U4108 (N_4108,N_3996,N_3956);
xor U4109 (N_4109,N_3996,N_3977);
nor U4110 (N_4110,N_3948,N_3871);
xnor U4111 (N_4111,N_3961,N_3908);
nor U4112 (N_4112,N_3918,N_3935);
and U4113 (N_4113,N_3910,N_3871);
nor U4114 (N_4114,N_3977,N_3938);
nor U4115 (N_4115,N_3862,N_3881);
nand U4116 (N_4116,N_3984,N_3870);
nand U4117 (N_4117,N_3952,N_3928);
nor U4118 (N_4118,N_3945,N_3929);
nand U4119 (N_4119,N_3843,N_3883);
xor U4120 (N_4120,N_3854,N_3929);
nand U4121 (N_4121,N_3944,N_3947);
and U4122 (N_4122,N_3975,N_3967);
or U4123 (N_4123,N_3862,N_3893);
xnor U4124 (N_4124,N_3928,N_3847);
and U4125 (N_4125,N_3965,N_3969);
or U4126 (N_4126,N_3953,N_3961);
nor U4127 (N_4127,N_3897,N_3946);
nand U4128 (N_4128,N_3990,N_3845);
nor U4129 (N_4129,N_3962,N_3945);
and U4130 (N_4130,N_3884,N_3876);
or U4131 (N_4131,N_3849,N_3990);
nand U4132 (N_4132,N_3861,N_3853);
and U4133 (N_4133,N_3946,N_3850);
and U4134 (N_4134,N_3929,N_3996);
xor U4135 (N_4135,N_3927,N_3873);
nand U4136 (N_4136,N_3953,N_3894);
nor U4137 (N_4137,N_3919,N_3882);
or U4138 (N_4138,N_3873,N_3879);
nand U4139 (N_4139,N_3879,N_3964);
xor U4140 (N_4140,N_3961,N_3921);
and U4141 (N_4141,N_3840,N_3914);
xor U4142 (N_4142,N_3843,N_3966);
and U4143 (N_4143,N_3945,N_3943);
xnor U4144 (N_4144,N_3846,N_3945);
nand U4145 (N_4145,N_3997,N_3984);
nand U4146 (N_4146,N_3840,N_3960);
xor U4147 (N_4147,N_3941,N_3894);
xor U4148 (N_4148,N_3922,N_3971);
or U4149 (N_4149,N_3898,N_3877);
xnor U4150 (N_4150,N_3854,N_3881);
nand U4151 (N_4151,N_3928,N_3868);
or U4152 (N_4152,N_3932,N_3993);
and U4153 (N_4153,N_3927,N_3862);
xor U4154 (N_4154,N_3855,N_3895);
nor U4155 (N_4155,N_3908,N_3994);
and U4156 (N_4156,N_3895,N_3886);
and U4157 (N_4157,N_3874,N_3954);
xor U4158 (N_4158,N_3856,N_3893);
xnor U4159 (N_4159,N_3973,N_3958);
and U4160 (N_4160,N_4003,N_4027);
xnor U4161 (N_4161,N_4081,N_4140);
and U4162 (N_4162,N_4141,N_4051);
nand U4163 (N_4163,N_4031,N_4015);
nor U4164 (N_4164,N_4073,N_4108);
or U4165 (N_4165,N_4138,N_4110);
or U4166 (N_4166,N_4012,N_4152);
and U4167 (N_4167,N_4028,N_4022);
nor U4168 (N_4168,N_4062,N_4066);
nor U4169 (N_4169,N_4047,N_4098);
and U4170 (N_4170,N_4041,N_4059);
nand U4171 (N_4171,N_4023,N_4053);
xnor U4172 (N_4172,N_4118,N_4016);
nand U4173 (N_4173,N_4033,N_4029);
and U4174 (N_4174,N_4013,N_4080);
xnor U4175 (N_4175,N_4144,N_4122);
and U4176 (N_4176,N_4109,N_4101);
and U4177 (N_4177,N_4125,N_4063);
nor U4178 (N_4178,N_4052,N_4032);
and U4179 (N_4179,N_4045,N_4020);
nand U4180 (N_4180,N_4034,N_4120);
and U4181 (N_4181,N_4078,N_4159);
and U4182 (N_4182,N_4007,N_4105);
nand U4183 (N_4183,N_4035,N_4021);
xnor U4184 (N_4184,N_4088,N_4093);
nor U4185 (N_4185,N_4157,N_4124);
or U4186 (N_4186,N_4100,N_4149);
and U4187 (N_4187,N_4116,N_4134);
xor U4188 (N_4188,N_4090,N_4004);
xnor U4189 (N_4189,N_4112,N_4074);
xnor U4190 (N_4190,N_4114,N_4057);
nor U4191 (N_4191,N_4133,N_4077);
xor U4192 (N_4192,N_4106,N_4038);
or U4193 (N_4193,N_4072,N_4000);
and U4194 (N_4194,N_4089,N_4084);
and U4195 (N_4195,N_4097,N_4131);
xor U4196 (N_4196,N_4130,N_4019);
xnor U4197 (N_4197,N_4070,N_4071);
or U4198 (N_4198,N_4076,N_4111);
nand U4199 (N_4199,N_4024,N_4129);
and U4200 (N_4200,N_4147,N_4086);
and U4201 (N_4201,N_4099,N_4127);
xnor U4202 (N_4202,N_4043,N_4067);
and U4203 (N_4203,N_4121,N_4126);
and U4204 (N_4204,N_4069,N_4154);
nor U4205 (N_4205,N_4049,N_4151);
and U4206 (N_4206,N_4018,N_4055);
and U4207 (N_4207,N_4039,N_4011);
nand U4208 (N_4208,N_4104,N_4006);
or U4209 (N_4209,N_4119,N_4046);
nand U4210 (N_4210,N_4058,N_4132);
or U4211 (N_4211,N_4095,N_4117);
and U4212 (N_4212,N_4153,N_4079);
nor U4213 (N_4213,N_4014,N_4158);
xnor U4214 (N_4214,N_4083,N_4136);
or U4215 (N_4215,N_4115,N_4128);
nor U4216 (N_4216,N_4001,N_4009);
nor U4217 (N_4217,N_4008,N_4146);
nand U4218 (N_4218,N_4087,N_4075);
and U4219 (N_4219,N_4085,N_4048);
and U4220 (N_4220,N_4143,N_4139);
or U4221 (N_4221,N_4137,N_4150);
and U4222 (N_4222,N_4037,N_4103);
and U4223 (N_4223,N_4017,N_4156);
or U4224 (N_4224,N_4056,N_4005);
and U4225 (N_4225,N_4054,N_4123);
or U4226 (N_4226,N_4060,N_4155);
or U4227 (N_4227,N_4107,N_4050);
and U4228 (N_4228,N_4010,N_4042);
xor U4229 (N_4229,N_4026,N_4044);
and U4230 (N_4230,N_4068,N_4040);
xor U4231 (N_4231,N_4102,N_4142);
and U4232 (N_4232,N_4091,N_4036);
nand U4233 (N_4233,N_4061,N_4064);
and U4234 (N_4234,N_4148,N_4096);
nor U4235 (N_4235,N_4113,N_4030);
xnor U4236 (N_4236,N_4082,N_4025);
xor U4237 (N_4237,N_4065,N_4002);
xnor U4238 (N_4238,N_4135,N_4145);
or U4239 (N_4239,N_4094,N_4092);
and U4240 (N_4240,N_4087,N_4109);
or U4241 (N_4241,N_4016,N_4043);
or U4242 (N_4242,N_4048,N_4157);
nor U4243 (N_4243,N_4155,N_4091);
or U4244 (N_4244,N_4021,N_4072);
and U4245 (N_4245,N_4013,N_4113);
and U4246 (N_4246,N_4016,N_4080);
nand U4247 (N_4247,N_4130,N_4049);
xnor U4248 (N_4248,N_4128,N_4042);
nor U4249 (N_4249,N_4027,N_4138);
or U4250 (N_4250,N_4079,N_4098);
xnor U4251 (N_4251,N_4006,N_4103);
nand U4252 (N_4252,N_4151,N_4026);
nor U4253 (N_4253,N_4156,N_4118);
xnor U4254 (N_4254,N_4070,N_4061);
or U4255 (N_4255,N_4103,N_4091);
xor U4256 (N_4256,N_4038,N_4020);
or U4257 (N_4257,N_4024,N_4037);
or U4258 (N_4258,N_4026,N_4063);
or U4259 (N_4259,N_4136,N_4089);
xor U4260 (N_4260,N_4062,N_4018);
and U4261 (N_4261,N_4072,N_4134);
xnor U4262 (N_4262,N_4016,N_4136);
nor U4263 (N_4263,N_4014,N_4093);
nand U4264 (N_4264,N_4020,N_4156);
nor U4265 (N_4265,N_4155,N_4050);
and U4266 (N_4266,N_4095,N_4061);
nor U4267 (N_4267,N_4156,N_4003);
or U4268 (N_4268,N_4130,N_4027);
nand U4269 (N_4269,N_4055,N_4006);
and U4270 (N_4270,N_4064,N_4099);
xor U4271 (N_4271,N_4159,N_4017);
nor U4272 (N_4272,N_4024,N_4139);
or U4273 (N_4273,N_4148,N_4008);
or U4274 (N_4274,N_4025,N_4112);
nor U4275 (N_4275,N_4044,N_4033);
xnor U4276 (N_4276,N_4037,N_4006);
or U4277 (N_4277,N_4078,N_4000);
and U4278 (N_4278,N_4044,N_4024);
nand U4279 (N_4279,N_4154,N_4051);
nor U4280 (N_4280,N_4071,N_4003);
and U4281 (N_4281,N_4007,N_4099);
nor U4282 (N_4282,N_4053,N_4037);
or U4283 (N_4283,N_4048,N_4034);
xnor U4284 (N_4284,N_4026,N_4098);
nor U4285 (N_4285,N_4119,N_4083);
nand U4286 (N_4286,N_4033,N_4040);
nand U4287 (N_4287,N_4025,N_4136);
nor U4288 (N_4288,N_4146,N_4088);
and U4289 (N_4289,N_4094,N_4006);
xnor U4290 (N_4290,N_4058,N_4066);
or U4291 (N_4291,N_4051,N_4123);
xor U4292 (N_4292,N_4092,N_4057);
and U4293 (N_4293,N_4079,N_4113);
nor U4294 (N_4294,N_4046,N_4152);
or U4295 (N_4295,N_4086,N_4010);
xor U4296 (N_4296,N_4089,N_4108);
xnor U4297 (N_4297,N_4127,N_4011);
nand U4298 (N_4298,N_4124,N_4148);
and U4299 (N_4299,N_4103,N_4102);
nand U4300 (N_4300,N_4031,N_4112);
or U4301 (N_4301,N_4070,N_4093);
nor U4302 (N_4302,N_4108,N_4064);
and U4303 (N_4303,N_4120,N_4124);
nor U4304 (N_4304,N_4072,N_4096);
nor U4305 (N_4305,N_4143,N_4057);
nor U4306 (N_4306,N_4025,N_4050);
and U4307 (N_4307,N_4068,N_4059);
xnor U4308 (N_4308,N_4075,N_4140);
and U4309 (N_4309,N_4129,N_4031);
and U4310 (N_4310,N_4061,N_4014);
or U4311 (N_4311,N_4094,N_4123);
and U4312 (N_4312,N_4005,N_4149);
nor U4313 (N_4313,N_4075,N_4091);
or U4314 (N_4314,N_4008,N_4100);
or U4315 (N_4315,N_4088,N_4110);
nor U4316 (N_4316,N_4054,N_4032);
xor U4317 (N_4317,N_4140,N_4157);
nor U4318 (N_4318,N_4135,N_4115);
xnor U4319 (N_4319,N_4133,N_4117);
nor U4320 (N_4320,N_4286,N_4273);
and U4321 (N_4321,N_4267,N_4216);
nand U4322 (N_4322,N_4227,N_4288);
nand U4323 (N_4323,N_4232,N_4229);
xnor U4324 (N_4324,N_4257,N_4287);
nor U4325 (N_4325,N_4181,N_4207);
nand U4326 (N_4326,N_4316,N_4255);
nand U4327 (N_4327,N_4217,N_4304);
and U4328 (N_4328,N_4311,N_4292);
and U4329 (N_4329,N_4302,N_4172);
or U4330 (N_4330,N_4289,N_4160);
nor U4331 (N_4331,N_4193,N_4163);
nand U4332 (N_4332,N_4263,N_4196);
nor U4333 (N_4333,N_4223,N_4260);
nand U4334 (N_4334,N_4310,N_4240);
xor U4335 (N_4335,N_4228,N_4164);
nand U4336 (N_4336,N_4202,N_4280);
and U4337 (N_4337,N_4269,N_4317);
or U4338 (N_4338,N_4275,N_4262);
and U4339 (N_4339,N_4241,N_4266);
nor U4340 (N_4340,N_4190,N_4186);
or U4341 (N_4341,N_4197,N_4220);
xor U4342 (N_4342,N_4191,N_4282);
nand U4343 (N_4343,N_4290,N_4301);
xor U4344 (N_4344,N_4252,N_4174);
and U4345 (N_4345,N_4278,N_4259);
nand U4346 (N_4346,N_4284,N_4265);
xnor U4347 (N_4347,N_4293,N_4246);
or U4348 (N_4348,N_4319,N_4224);
or U4349 (N_4349,N_4307,N_4291);
xnor U4350 (N_4350,N_4299,N_4218);
nor U4351 (N_4351,N_4165,N_4243);
xnor U4352 (N_4352,N_4188,N_4281);
xnor U4353 (N_4353,N_4214,N_4314);
or U4354 (N_4354,N_4251,N_4176);
nand U4355 (N_4355,N_4274,N_4247);
nand U4356 (N_4356,N_4200,N_4206);
nor U4357 (N_4357,N_4221,N_4180);
nand U4358 (N_4358,N_4279,N_4222);
nand U4359 (N_4359,N_4204,N_4199);
nor U4360 (N_4360,N_4212,N_4276);
and U4361 (N_4361,N_4238,N_4237);
nor U4362 (N_4362,N_4234,N_4272);
xnor U4363 (N_4363,N_4283,N_4225);
or U4364 (N_4364,N_4230,N_4318);
nor U4365 (N_4365,N_4203,N_4201);
and U4366 (N_4366,N_4185,N_4189);
or U4367 (N_4367,N_4305,N_4183);
or U4368 (N_4368,N_4177,N_4236);
nor U4369 (N_4369,N_4261,N_4270);
or U4370 (N_4370,N_4285,N_4297);
or U4371 (N_4371,N_4268,N_4303);
nor U4372 (N_4372,N_4208,N_4187);
or U4373 (N_4373,N_4226,N_4306);
nor U4374 (N_4374,N_4171,N_4248);
and U4375 (N_4375,N_4175,N_4161);
or U4376 (N_4376,N_4162,N_4231);
or U4377 (N_4377,N_4249,N_4277);
nor U4378 (N_4378,N_4245,N_4315);
nor U4379 (N_4379,N_4313,N_4179);
xor U4380 (N_4380,N_4312,N_4167);
xor U4381 (N_4381,N_4205,N_4296);
nor U4382 (N_4382,N_4173,N_4258);
and U4383 (N_4383,N_4300,N_4215);
xnor U4384 (N_4384,N_4253,N_4242);
xor U4385 (N_4385,N_4184,N_4254);
or U4386 (N_4386,N_4250,N_4182);
xnor U4387 (N_4387,N_4194,N_4192);
nor U4388 (N_4388,N_4235,N_4166);
nand U4389 (N_4389,N_4294,N_4198);
xor U4390 (N_4390,N_4219,N_4308);
xor U4391 (N_4391,N_4239,N_4264);
nand U4392 (N_4392,N_4210,N_4256);
or U4393 (N_4393,N_4178,N_4271);
and U4394 (N_4394,N_4211,N_4169);
or U4395 (N_4395,N_4209,N_4170);
xor U4396 (N_4396,N_4309,N_4295);
nor U4397 (N_4397,N_4195,N_4213);
xnor U4398 (N_4398,N_4168,N_4244);
nor U4399 (N_4399,N_4233,N_4298);
and U4400 (N_4400,N_4240,N_4266);
xor U4401 (N_4401,N_4165,N_4206);
or U4402 (N_4402,N_4294,N_4200);
or U4403 (N_4403,N_4268,N_4199);
nand U4404 (N_4404,N_4189,N_4290);
or U4405 (N_4405,N_4260,N_4174);
xnor U4406 (N_4406,N_4301,N_4183);
nor U4407 (N_4407,N_4271,N_4291);
xnor U4408 (N_4408,N_4303,N_4311);
and U4409 (N_4409,N_4192,N_4179);
xnor U4410 (N_4410,N_4265,N_4315);
and U4411 (N_4411,N_4251,N_4298);
and U4412 (N_4412,N_4198,N_4262);
or U4413 (N_4413,N_4277,N_4191);
xor U4414 (N_4414,N_4183,N_4179);
nor U4415 (N_4415,N_4239,N_4181);
nor U4416 (N_4416,N_4242,N_4195);
or U4417 (N_4417,N_4164,N_4248);
and U4418 (N_4418,N_4235,N_4180);
nor U4419 (N_4419,N_4303,N_4310);
nand U4420 (N_4420,N_4269,N_4252);
or U4421 (N_4421,N_4290,N_4227);
nor U4422 (N_4422,N_4306,N_4173);
xnor U4423 (N_4423,N_4280,N_4170);
xnor U4424 (N_4424,N_4317,N_4313);
nor U4425 (N_4425,N_4279,N_4192);
and U4426 (N_4426,N_4209,N_4272);
nor U4427 (N_4427,N_4304,N_4231);
nand U4428 (N_4428,N_4296,N_4249);
nor U4429 (N_4429,N_4205,N_4252);
nor U4430 (N_4430,N_4179,N_4284);
nand U4431 (N_4431,N_4277,N_4291);
nand U4432 (N_4432,N_4211,N_4215);
or U4433 (N_4433,N_4204,N_4316);
or U4434 (N_4434,N_4210,N_4259);
or U4435 (N_4435,N_4168,N_4308);
and U4436 (N_4436,N_4188,N_4275);
and U4437 (N_4437,N_4184,N_4163);
xnor U4438 (N_4438,N_4314,N_4259);
or U4439 (N_4439,N_4175,N_4302);
or U4440 (N_4440,N_4299,N_4233);
or U4441 (N_4441,N_4275,N_4175);
and U4442 (N_4442,N_4210,N_4309);
nand U4443 (N_4443,N_4288,N_4290);
nor U4444 (N_4444,N_4161,N_4277);
nand U4445 (N_4445,N_4253,N_4217);
nor U4446 (N_4446,N_4247,N_4253);
xor U4447 (N_4447,N_4266,N_4290);
nand U4448 (N_4448,N_4313,N_4221);
nor U4449 (N_4449,N_4201,N_4200);
nor U4450 (N_4450,N_4191,N_4224);
nand U4451 (N_4451,N_4289,N_4198);
xor U4452 (N_4452,N_4218,N_4165);
nand U4453 (N_4453,N_4190,N_4256);
nand U4454 (N_4454,N_4230,N_4246);
and U4455 (N_4455,N_4303,N_4196);
or U4456 (N_4456,N_4281,N_4280);
nand U4457 (N_4457,N_4274,N_4261);
and U4458 (N_4458,N_4162,N_4227);
xnor U4459 (N_4459,N_4314,N_4263);
nand U4460 (N_4460,N_4305,N_4260);
nand U4461 (N_4461,N_4213,N_4164);
nor U4462 (N_4462,N_4199,N_4283);
and U4463 (N_4463,N_4192,N_4246);
nand U4464 (N_4464,N_4220,N_4209);
nand U4465 (N_4465,N_4296,N_4223);
nor U4466 (N_4466,N_4312,N_4293);
xor U4467 (N_4467,N_4170,N_4213);
nand U4468 (N_4468,N_4302,N_4263);
nand U4469 (N_4469,N_4257,N_4286);
and U4470 (N_4470,N_4318,N_4201);
and U4471 (N_4471,N_4216,N_4208);
nor U4472 (N_4472,N_4272,N_4299);
xnor U4473 (N_4473,N_4171,N_4196);
nor U4474 (N_4474,N_4226,N_4179);
nand U4475 (N_4475,N_4311,N_4281);
nand U4476 (N_4476,N_4186,N_4251);
or U4477 (N_4477,N_4255,N_4300);
or U4478 (N_4478,N_4210,N_4241);
xor U4479 (N_4479,N_4308,N_4260);
or U4480 (N_4480,N_4385,N_4464);
or U4481 (N_4481,N_4346,N_4365);
or U4482 (N_4482,N_4403,N_4320);
xor U4483 (N_4483,N_4352,N_4387);
and U4484 (N_4484,N_4442,N_4359);
nand U4485 (N_4485,N_4366,N_4446);
nand U4486 (N_4486,N_4378,N_4321);
xnor U4487 (N_4487,N_4329,N_4324);
and U4488 (N_4488,N_4460,N_4423);
xor U4489 (N_4489,N_4374,N_4358);
and U4490 (N_4490,N_4475,N_4382);
nor U4491 (N_4491,N_4331,N_4344);
nor U4492 (N_4492,N_4419,N_4415);
xor U4493 (N_4493,N_4361,N_4407);
or U4494 (N_4494,N_4333,N_4369);
and U4495 (N_4495,N_4367,N_4342);
nor U4496 (N_4496,N_4398,N_4376);
nand U4497 (N_4497,N_4364,N_4345);
and U4498 (N_4498,N_4392,N_4455);
and U4499 (N_4499,N_4427,N_4356);
nor U4500 (N_4500,N_4472,N_4424);
nor U4501 (N_4501,N_4373,N_4405);
nand U4502 (N_4502,N_4441,N_4445);
xnor U4503 (N_4503,N_4452,N_4397);
and U4504 (N_4504,N_4395,N_4474);
nor U4505 (N_4505,N_4323,N_4335);
nor U4506 (N_4506,N_4443,N_4449);
or U4507 (N_4507,N_4383,N_4380);
nor U4508 (N_4508,N_4476,N_4447);
xnor U4509 (N_4509,N_4466,N_4340);
xnor U4510 (N_4510,N_4393,N_4370);
and U4511 (N_4511,N_4468,N_4347);
nor U4512 (N_4512,N_4325,N_4430);
and U4513 (N_4513,N_4371,N_4363);
nor U4514 (N_4514,N_4360,N_4357);
nand U4515 (N_4515,N_4432,N_4471);
or U4516 (N_4516,N_4428,N_4435);
or U4517 (N_4517,N_4326,N_4355);
and U4518 (N_4518,N_4413,N_4379);
xnor U4519 (N_4519,N_4422,N_4436);
nor U4520 (N_4520,N_4375,N_4394);
and U4521 (N_4521,N_4404,N_4479);
nand U4522 (N_4522,N_4334,N_4388);
nor U4523 (N_4523,N_4421,N_4339);
xnor U4524 (N_4524,N_4337,N_4399);
xnor U4525 (N_4525,N_4463,N_4332);
or U4526 (N_4526,N_4351,N_4450);
xor U4527 (N_4527,N_4377,N_4350);
xor U4528 (N_4528,N_4400,N_4448);
or U4529 (N_4529,N_4470,N_4429);
and U4530 (N_4530,N_4416,N_4389);
nand U4531 (N_4531,N_4402,N_4362);
xor U4532 (N_4532,N_4461,N_4336);
or U4533 (N_4533,N_4469,N_4438);
nand U4534 (N_4534,N_4354,N_4408);
or U4535 (N_4535,N_4386,N_4437);
nand U4536 (N_4536,N_4458,N_4425);
or U4537 (N_4537,N_4451,N_4417);
xor U4538 (N_4538,N_4462,N_4390);
and U4539 (N_4539,N_4330,N_4440);
nand U4540 (N_4540,N_4349,N_4456);
and U4541 (N_4541,N_4372,N_4411);
xnor U4542 (N_4542,N_4353,N_4391);
and U4543 (N_4543,N_4327,N_4348);
nand U4544 (N_4544,N_4396,N_4453);
and U4545 (N_4545,N_4434,N_4381);
nand U4546 (N_4546,N_4328,N_4341);
or U4547 (N_4547,N_4368,N_4420);
and U4548 (N_4548,N_4465,N_4467);
and U4549 (N_4549,N_4454,N_4439);
or U4550 (N_4550,N_4384,N_4473);
nand U4551 (N_4551,N_4418,N_4459);
nand U4552 (N_4552,N_4477,N_4412);
xnor U4553 (N_4553,N_4433,N_4343);
or U4554 (N_4554,N_4431,N_4426);
xnor U4555 (N_4555,N_4338,N_4322);
xor U4556 (N_4556,N_4401,N_4409);
nor U4557 (N_4557,N_4414,N_4457);
nor U4558 (N_4558,N_4444,N_4406);
and U4559 (N_4559,N_4478,N_4410);
and U4560 (N_4560,N_4385,N_4372);
nor U4561 (N_4561,N_4353,N_4337);
nor U4562 (N_4562,N_4374,N_4323);
nor U4563 (N_4563,N_4371,N_4327);
nand U4564 (N_4564,N_4384,N_4416);
or U4565 (N_4565,N_4413,N_4369);
and U4566 (N_4566,N_4327,N_4372);
xnor U4567 (N_4567,N_4382,N_4342);
nor U4568 (N_4568,N_4412,N_4387);
or U4569 (N_4569,N_4399,N_4346);
nor U4570 (N_4570,N_4367,N_4399);
or U4571 (N_4571,N_4352,N_4359);
nand U4572 (N_4572,N_4345,N_4435);
nand U4573 (N_4573,N_4477,N_4347);
nand U4574 (N_4574,N_4399,N_4405);
nor U4575 (N_4575,N_4352,N_4433);
nand U4576 (N_4576,N_4463,N_4471);
xor U4577 (N_4577,N_4331,N_4469);
or U4578 (N_4578,N_4324,N_4378);
xor U4579 (N_4579,N_4387,N_4473);
nor U4580 (N_4580,N_4470,N_4361);
xor U4581 (N_4581,N_4338,N_4377);
and U4582 (N_4582,N_4456,N_4474);
nor U4583 (N_4583,N_4384,N_4436);
and U4584 (N_4584,N_4410,N_4477);
or U4585 (N_4585,N_4401,N_4461);
nor U4586 (N_4586,N_4419,N_4384);
nand U4587 (N_4587,N_4360,N_4384);
or U4588 (N_4588,N_4326,N_4344);
xor U4589 (N_4589,N_4348,N_4376);
nand U4590 (N_4590,N_4339,N_4432);
nor U4591 (N_4591,N_4433,N_4321);
nor U4592 (N_4592,N_4451,N_4342);
and U4593 (N_4593,N_4321,N_4422);
nand U4594 (N_4594,N_4399,N_4468);
nand U4595 (N_4595,N_4424,N_4438);
nand U4596 (N_4596,N_4354,N_4346);
nor U4597 (N_4597,N_4330,N_4376);
or U4598 (N_4598,N_4461,N_4426);
and U4599 (N_4599,N_4331,N_4361);
or U4600 (N_4600,N_4392,N_4400);
or U4601 (N_4601,N_4385,N_4439);
nand U4602 (N_4602,N_4381,N_4326);
nand U4603 (N_4603,N_4426,N_4475);
nor U4604 (N_4604,N_4376,N_4458);
or U4605 (N_4605,N_4442,N_4327);
and U4606 (N_4606,N_4406,N_4443);
or U4607 (N_4607,N_4389,N_4395);
xor U4608 (N_4608,N_4438,N_4447);
xor U4609 (N_4609,N_4469,N_4413);
nand U4610 (N_4610,N_4445,N_4369);
nand U4611 (N_4611,N_4438,N_4419);
nand U4612 (N_4612,N_4347,N_4327);
or U4613 (N_4613,N_4409,N_4439);
and U4614 (N_4614,N_4353,N_4453);
nor U4615 (N_4615,N_4419,N_4374);
and U4616 (N_4616,N_4456,N_4415);
and U4617 (N_4617,N_4448,N_4413);
or U4618 (N_4618,N_4434,N_4356);
and U4619 (N_4619,N_4399,N_4371);
nand U4620 (N_4620,N_4421,N_4441);
nand U4621 (N_4621,N_4359,N_4393);
nand U4622 (N_4622,N_4364,N_4381);
nor U4623 (N_4623,N_4419,N_4435);
xor U4624 (N_4624,N_4402,N_4465);
nor U4625 (N_4625,N_4431,N_4410);
and U4626 (N_4626,N_4329,N_4443);
and U4627 (N_4627,N_4369,N_4443);
xor U4628 (N_4628,N_4448,N_4395);
nand U4629 (N_4629,N_4473,N_4477);
nand U4630 (N_4630,N_4413,N_4376);
and U4631 (N_4631,N_4413,N_4408);
or U4632 (N_4632,N_4381,N_4419);
nor U4633 (N_4633,N_4347,N_4395);
and U4634 (N_4634,N_4353,N_4379);
and U4635 (N_4635,N_4449,N_4415);
nor U4636 (N_4636,N_4395,N_4382);
xor U4637 (N_4637,N_4440,N_4428);
xnor U4638 (N_4638,N_4365,N_4420);
and U4639 (N_4639,N_4459,N_4370);
and U4640 (N_4640,N_4533,N_4541);
or U4641 (N_4641,N_4523,N_4580);
xor U4642 (N_4642,N_4601,N_4487);
and U4643 (N_4643,N_4520,N_4618);
xor U4644 (N_4644,N_4584,N_4581);
xnor U4645 (N_4645,N_4539,N_4612);
xnor U4646 (N_4646,N_4611,N_4518);
nor U4647 (N_4647,N_4583,N_4565);
or U4648 (N_4648,N_4592,N_4575);
or U4649 (N_4649,N_4628,N_4531);
and U4650 (N_4650,N_4627,N_4622);
or U4651 (N_4651,N_4486,N_4615);
xnor U4652 (N_4652,N_4516,N_4483);
nor U4653 (N_4653,N_4527,N_4495);
xnor U4654 (N_4654,N_4546,N_4543);
and U4655 (N_4655,N_4590,N_4536);
nor U4656 (N_4656,N_4578,N_4513);
and U4657 (N_4657,N_4600,N_4501);
or U4658 (N_4658,N_4639,N_4579);
nand U4659 (N_4659,N_4638,N_4571);
and U4660 (N_4660,N_4555,N_4561);
nand U4661 (N_4661,N_4493,N_4631);
and U4662 (N_4662,N_4537,N_4498);
xnor U4663 (N_4663,N_4564,N_4599);
nor U4664 (N_4664,N_4634,N_4551);
nor U4665 (N_4665,N_4485,N_4481);
or U4666 (N_4666,N_4549,N_4522);
and U4667 (N_4667,N_4614,N_4482);
nand U4668 (N_4668,N_4560,N_4530);
nand U4669 (N_4669,N_4598,N_4542);
xor U4670 (N_4670,N_4517,N_4604);
nor U4671 (N_4671,N_4635,N_4566);
xor U4672 (N_4672,N_4594,N_4607);
xor U4673 (N_4673,N_4507,N_4605);
or U4674 (N_4674,N_4608,N_4562);
and U4675 (N_4675,N_4509,N_4573);
nand U4676 (N_4676,N_4510,N_4621);
and U4677 (N_4677,N_4595,N_4609);
xnor U4678 (N_4678,N_4596,N_4557);
or U4679 (N_4679,N_4519,N_4526);
nor U4680 (N_4680,N_4589,N_4626);
xor U4681 (N_4681,N_4490,N_4494);
and U4682 (N_4682,N_4619,N_4524);
xor U4683 (N_4683,N_4624,N_4540);
xor U4684 (N_4684,N_4491,N_4528);
and U4685 (N_4685,N_4617,N_4512);
nor U4686 (N_4686,N_4552,N_4502);
nand U4687 (N_4687,N_4620,N_4633);
and U4688 (N_4688,N_4606,N_4497);
and U4689 (N_4689,N_4572,N_4484);
nand U4690 (N_4690,N_4496,N_4544);
nor U4691 (N_4691,N_4616,N_4480);
nand U4692 (N_4692,N_4503,N_4637);
and U4693 (N_4693,N_4489,N_4488);
or U4694 (N_4694,N_4567,N_4554);
xnor U4695 (N_4695,N_4587,N_4500);
nor U4696 (N_4696,N_4559,N_4603);
xnor U4697 (N_4697,N_4534,N_4563);
xor U4698 (N_4698,N_4574,N_4582);
xnor U4699 (N_4699,N_4553,N_4547);
nand U4700 (N_4700,N_4492,N_4556);
or U4701 (N_4701,N_4602,N_4506);
xor U4702 (N_4702,N_4632,N_4586);
nor U4703 (N_4703,N_4568,N_4535);
or U4704 (N_4704,N_4577,N_4504);
or U4705 (N_4705,N_4588,N_4514);
nor U4706 (N_4706,N_4591,N_4623);
xnor U4707 (N_4707,N_4521,N_4545);
and U4708 (N_4708,N_4570,N_4505);
or U4709 (N_4709,N_4630,N_4548);
nand U4710 (N_4710,N_4499,N_4593);
or U4711 (N_4711,N_4629,N_4585);
or U4712 (N_4712,N_4529,N_4597);
nor U4713 (N_4713,N_4508,N_4511);
nor U4714 (N_4714,N_4625,N_4576);
or U4715 (N_4715,N_4525,N_4532);
nand U4716 (N_4716,N_4515,N_4636);
or U4717 (N_4717,N_4538,N_4613);
nand U4718 (N_4718,N_4550,N_4610);
nor U4719 (N_4719,N_4569,N_4558);
nand U4720 (N_4720,N_4589,N_4621);
nand U4721 (N_4721,N_4549,N_4564);
nand U4722 (N_4722,N_4558,N_4524);
xor U4723 (N_4723,N_4618,N_4493);
or U4724 (N_4724,N_4618,N_4616);
xor U4725 (N_4725,N_4569,N_4481);
nand U4726 (N_4726,N_4573,N_4532);
nand U4727 (N_4727,N_4521,N_4582);
nor U4728 (N_4728,N_4536,N_4566);
or U4729 (N_4729,N_4630,N_4539);
and U4730 (N_4730,N_4607,N_4593);
or U4731 (N_4731,N_4536,N_4530);
or U4732 (N_4732,N_4558,N_4571);
nand U4733 (N_4733,N_4498,N_4628);
and U4734 (N_4734,N_4583,N_4524);
xnor U4735 (N_4735,N_4541,N_4576);
and U4736 (N_4736,N_4497,N_4610);
nor U4737 (N_4737,N_4614,N_4627);
and U4738 (N_4738,N_4502,N_4486);
nor U4739 (N_4739,N_4517,N_4639);
or U4740 (N_4740,N_4522,N_4552);
nor U4741 (N_4741,N_4582,N_4587);
nand U4742 (N_4742,N_4503,N_4570);
or U4743 (N_4743,N_4499,N_4480);
nand U4744 (N_4744,N_4602,N_4508);
nand U4745 (N_4745,N_4569,N_4546);
nand U4746 (N_4746,N_4559,N_4515);
and U4747 (N_4747,N_4608,N_4494);
xor U4748 (N_4748,N_4602,N_4491);
xnor U4749 (N_4749,N_4574,N_4575);
xnor U4750 (N_4750,N_4557,N_4492);
nor U4751 (N_4751,N_4499,N_4583);
xor U4752 (N_4752,N_4494,N_4638);
and U4753 (N_4753,N_4538,N_4545);
xor U4754 (N_4754,N_4535,N_4622);
or U4755 (N_4755,N_4605,N_4549);
and U4756 (N_4756,N_4551,N_4547);
or U4757 (N_4757,N_4570,N_4562);
and U4758 (N_4758,N_4573,N_4544);
xor U4759 (N_4759,N_4585,N_4566);
and U4760 (N_4760,N_4612,N_4602);
nor U4761 (N_4761,N_4519,N_4506);
or U4762 (N_4762,N_4576,N_4533);
and U4763 (N_4763,N_4631,N_4515);
nand U4764 (N_4764,N_4546,N_4512);
nor U4765 (N_4765,N_4614,N_4582);
xnor U4766 (N_4766,N_4556,N_4595);
nor U4767 (N_4767,N_4622,N_4618);
or U4768 (N_4768,N_4577,N_4535);
and U4769 (N_4769,N_4599,N_4562);
nor U4770 (N_4770,N_4508,N_4546);
nand U4771 (N_4771,N_4521,N_4511);
nor U4772 (N_4772,N_4603,N_4549);
or U4773 (N_4773,N_4571,N_4498);
or U4774 (N_4774,N_4634,N_4555);
nor U4775 (N_4775,N_4589,N_4495);
and U4776 (N_4776,N_4480,N_4510);
nor U4777 (N_4777,N_4572,N_4627);
or U4778 (N_4778,N_4530,N_4617);
xnor U4779 (N_4779,N_4608,N_4635);
nor U4780 (N_4780,N_4480,N_4537);
and U4781 (N_4781,N_4517,N_4598);
and U4782 (N_4782,N_4563,N_4579);
nand U4783 (N_4783,N_4558,N_4624);
nor U4784 (N_4784,N_4531,N_4615);
nand U4785 (N_4785,N_4481,N_4510);
or U4786 (N_4786,N_4610,N_4639);
xor U4787 (N_4787,N_4563,N_4639);
or U4788 (N_4788,N_4618,N_4599);
or U4789 (N_4789,N_4554,N_4516);
or U4790 (N_4790,N_4532,N_4536);
xnor U4791 (N_4791,N_4517,N_4509);
nor U4792 (N_4792,N_4555,N_4623);
nor U4793 (N_4793,N_4499,N_4615);
nor U4794 (N_4794,N_4565,N_4534);
nor U4795 (N_4795,N_4482,N_4525);
nand U4796 (N_4796,N_4551,N_4560);
xnor U4797 (N_4797,N_4529,N_4522);
nand U4798 (N_4798,N_4503,N_4518);
xor U4799 (N_4799,N_4554,N_4509);
nor U4800 (N_4800,N_4728,N_4650);
xnor U4801 (N_4801,N_4666,N_4794);
and U4802 (N_4802,N_4669,N_4747);
nand U4803 (N_4803,N_4661,N_4726);
or U4804 (N_4804,N_4693,N_4679);
and U4805 (N_4805,N_4695,N_4729);
and U4806 (N_4806,N_4767,N_4796);
and U4807 (N_4807,N_4741,N_4743);
and U4808 (N_4808,N_4668,N_4778);
xnor U4809 (N_4809,N_4694,N_4784);
xnor U4810 (N_4810,N_4783,N_4644);
and U4811 (N_4811,N_4643,N_4738);
or U4812 (N_4812,N_4671,N_4684);
or U4813 (N_4813,N_4721,N_4774);
and U4814 (N_4814,N_4762,N_4655);
or U4815 (N_4815,N_4710,N_4793);
and U4816 (N_4816,N_4775,N_4663);
nor U4817 (N_4817,N_4760,N_4786);
nor U4818 (N_4818,N_4697,N_4770);
and U4819 (N_4819,N_4727,N_4709);
nor U4820 (N_4820,N_4664,N_4753);
nand U4821 (N_4821,N_4702,N_4772);
xor U4822 (N_4822,N_4681,N_4674);
or U4823 (N_4823,N_4735,N_4676);
nor U4824 (N_4824,N_4717,N_4672);
and U4825 (N_4825,N_4649,N_4723);
and U4826 (N_4826,N_4665,N_4742);
nor U4827 (N_4827,N_4716,N_4788);
nand U4828 (N_4828,N_4799,N_4701);
nand U4829 (N_4829,N_4740,N_4759);
and U4830 (N_4830,N_4714,N_4641);
and U4831 (N_4831,N_4640,N_4752);
and U4832 (N_4832,N_4754,N_4703);
and U4833 (N_4833,N_4706,N_4699);
nor U4834 (N_4834,N_4686,N_4682);
xor U4835 (N_4835,N_4651,N_4696);
xor U4836 (N_4836,N_4779,N_4737);
or U4837 (N_4837,N_4751,N_4755);
and U4838 (N_4838,N_4654,N_4787);
nor U4839 (N_4839,N_4691,N_4781);
and U4840 (N_4840,N_4698,N_4647);
and U4841 (N_4841,N_4711,N_4648);
or U4842 (N_4842,N_4670,N_4790);
and U4843 (N_4843,N_4725,N_4705);
and U4844 (N_4844,N_4724,N_4746);
and U4845 (N_4845,N_4744,N_4687);
xor U4846 (N_4846,N_4761,N_4756);
or U4847 (N_4847,N_4777,N_4791);
and U4848 (N_4848,N_4704,N_4792);
nor U4849 (N_4849,N_4715,N_4734);
xor U4850 (N_4850,N_4678,N_4688);
nand U4851 (N_4851,N_4768,N_4731);
nand U4852 (N_4852,N_4749,N_4690);
xor U4853 (N_4853,N_4736,N_4773);
nor U4854 (N_4854,N_4733,N_4765);
nand U4855 (N_4855,N_4718,N_4713);
xnor U4856 (N_4856,N_4739,N_4667);
xnor U4857 (N_4857,N_4656,N_4782);
nor U4858 (N_4858,N_4795,N_4657);
or U4859 (N_4859,N_4662,N_4653);
and U4860 (N_4860,N_4645,N_4673);
nand U4861 (N_4861,N_4785,N_4677);
or U4862 (N_4862,N_4712,N_4764);
xnor U4863 (N_4863,N_4708,N_4750);
nand U4864 (N_4864,N_4642,N_4780);
and U4865 (N_4865,N_4789,N_4719);
and U4866 (N_4866,N_4748,N_4683);
or U4867 (N_4867,N_4675,N_4658);
xnor U4868 (N_4868,N_4692,N_4769);
or U4869 (N_4869,N_4758,N_4685);
nor U4870 (N_4870,N_4732,N_4766);
xnor U4871 (N_4871,N_4689,N_4722);
or U4872 (N_4872,N_4763,N_4652);
nand U4873 (N_4873,N_4720,N_4680);
and U4874 (N_4874,N_4646,N_4745);
nor U4875 (N_4875,N_4700,N_4730);
nand U4876 (N_4876,N_4776,N_4798);
nand U4877 (N_4877,N_4771,N_4757);
nand U4878 (N_4878,N_4659,N_4660);
nand U4879 (N_4879,N_4707,N_4797);
nand U4880 (N_4880,N_4681,N_4678);
or U4881 (N_4881,N_4785,N_4694);
and U4882 (N_4882,N_4690,N_4657);
nor U4883 (N_4883,N_4756,N_4743);
xor U4884 (N_4884,N_4703,N_4765);
and U4885 (N_4885,N_4666,N_4681);
or U4886 (N_4886,N_4738,N_4718);
and U4887 (N_4887,N_4790,N_4795);
xnor U4888 (N_4888,N_4764,N_4787);
xnor U4889 (N_4889,N_4768,N_4688);
nand U4890 (N_4890,N_4711,N_4680);
or U4891 (N_4891,N_4644,N_4770);
nor U4892 (N_4892,N_4769,N_4750);
xnor U4893 (N_4893,N_4734,N_4643);
and U4894 (N_4894,N_4707,N_4739);
and U4895 (N_4895,N_4671,N_4703);
or U4896 (N_4896,N_4777,N_4775);
nor U4897 (N_4897,N_4677,N_4767);
and U4898 (N_4898,N_4787,N_4774);
and U4899 (N_4899,N_4683,N_4778);
xor U4900 (N_4900,N_4698,N_4646);
xor U4901 (N_4901,N_4787,N_4712);
and U4902 (N_4902,N_4759,N_4787);
xor U4903 (N_4903,N_4798,N_4698);
and U4904 (N_4904,N_4767,N_4714);
or U4905 (N_4905,N_4771,N_4775);
and U4906 (N_4906,N_4669,N_4700);
xnor U4907 (N_4907,N_4797,N_4762);
nand U4908 (N_4908,N_4721,N_4664);
nand U4909 (N_4909,N_4696,N_4650);
nor U4910 (N_4910,N_4659,N_4698);
nand U4911 (N_4911,N_4726,N_4794);
and U4912 (N_4912,N_4777,N_4768);
and U4913 (N_4913,N_4721,N_4652);
xor U4914 (N_4914,N_4651,N_4662);
and U4915 (N_4915,N_4688,N_4796);
or U4916 (N_4916,N_4714,N_4640);
xnor U4917 (N_4917,N_4796,N_4722);
nor U4918 (N_4918,N_4731,N_4723);
and U4919 (N_4919,N_4684,N_4694);
or U4920 (N_4920,N_4704,N_4670);
nor U4921 (N_4921,N_4779,N_4754);
nor U4922 (N_4922,N_4757,N_4697);
nor U4923 (N_4923,N_4655,N_4737);
nor U4924 (N_4924,N_4655,N_4784);
and U4925 (N_4925,N_4654,N_4717);
nor U4926 (N_4926,N_4752,N_4797);
nor U4927 (N_4927,N_4665,N_4712);
and U4928 (N_4928,N_4652,N_4714);
xnor U4929 (N_4929,N_4792,N_4711);
nor U4930 (N_4930,N_4644,N_4790);
nand U4931 (N_4931,N_4799,N_4686);
or U4932 (N_4932,N_4663,N_4651);
and U4933 (N_4933,N_4766,N_4668);
nor U4934 (N_4934,N_4752,N_4683);
and U4935 (N_4935,N_4798,N_4689);
and U4936 (N_4936,N_4668,N_4701);
nor U4937 (N_4937,N_4766,N_4719);
nor U4938 (N_4938,N_4726,N_4645);
nand U4939 (N_4939,N_4703,N_4706);
nand U4940 (N_4940,N_4642,N_4772);
and U4941 (N_4941,N_4744,N_4773);
nor U4942 (N_4942,N_4669,N_4650);
nand U4943 (N_4943,N_4743,N_4663);
nor U4944 (N_4944,N_4659,N_4765);
nor U4945 (N_4945,N_4694,N_4739);
xnor U4946 (N_4946,N_4676,N_4780);
or U4947 (N_4947,N_4749,N_4662);
or U4948 (N_4948,N_4653,N_4794);
or U4949 (N_4949,N_4723,N_4651);
xnor U4950 (N_4950,N_4711,N_4732);
xor U4951 (N_4951,N_4775,N_4687);
or U4952 (N_4952,N_4739,N_4679);
and U4953 (N_4953,N_4680,N_4646);
xor U4954 (N_4954,N_4770,N_4663);
and U4955 (N_4955,N_4794,N_4738);
nand U4956 (N_4956,N_4708,N_4749);
or U4957 (N_4957,N_4774,N_4697);
xnor U4958 (N_4958,N_4691,N_4695);
xnor U4959 (N_4959,N_4687,N_4711);
nor U4960 (N_4960,N_4828,N_4808);
or U4961 (N_4961,N_4885,N_4934);
nand U4962 (N_4962,N_4865,N_4883);
nand U4963 (N_4963,N_4845,N_4857);
nand U4964 (N_4964,N_4878,N_4848);
or U4965 (N_4965,N_4953,N_4946);
nor U4966 (N_4966,N_4921,N_4899);
or U4967 (N_4967,N_4803,N_4952);
and U4968 (N_4968,N_4851,N_4884);
or U4969 (N_4969,N_4840,N_4954);
nor U4970 (N_4970,N_4866,N_4846);
nor U4971 (N_4971,N_4838,N_4829);
nor U4972 (N_4972,N_4825,N_4939);
nand U4973 (N_4973,N_4901,N_4912);
and U4974 (N_4974,N_4843,N_4852);
nand U4975 (N_4975,N_4872,N_4908);
xor U4976 (N_4976,N_4904,N_4919);
nand U4977 (N_4977,N_4940,N_4881);
xnor U4978 (N_4978,N_4859,N_4835);
nor U4979 (N_4979,N_4844,N_4943);
or U4980 (N_4980,N_4814,N_4900);
and U4981 (N_4981,N_4875,N_4930);
or U4982 (N_4982,N_4834,N_4874);
and U4983 (N_4983,N_4862,N_4896);
nand U4984 (N_4984,N_4891,N_4849);
xnor U4985 (N_4985,N_4842,N_4941);
nand U4986 (N_4986,N_4948,N_4922);
nand U4987 (N_4987,N_4817,N_4810);
and U4988 (N_4988,N_4898,N_4909);
nand U4989 (N_4989,N_4856,N_4932);
nor U4990 (N_4990,N_4928,N_4902);
or U4991 (N_4991,N_4906,N_4813);
and U4992 (N_4992,N_4812,N_4949);
nor U4993 (N_4993,N_4850,N_4889);
or U4994 (N_4994,N_4958,N_4839);
or U4995 (N_4995,N_4868,N_4876);
nand U4996 (N_4996,N_4860,N_4807);
nand U4997 (N_4997,N_4894,N_4947);
nor U4998 (N_4998,N_4867,N_4957);
and U4999 (N_4999,N_4925,N_4914);
and U5000 (N_5000,N_4927,N_4809);
xor U5001 (N_5001,N_4830,N_4800);
nor U5002 (N_5002,N_4879,N_4955);
nand U5003 (N_5003,N_4869,N_4805);
nand U5004 (N_5004,N_4826,N_4873);
nor U5005 (N_5005,N_4863,N_4815);
nor U5006 (N_5006,N_4847,N_4804);
nor U5007 (N_5007,N_4907,N_4951);
nor U5008 (N_5008,N_4819,N_4929);
or U5009 (N_5009,N_4905,N_4858);
and U5010 (N_5010,N_4924,N_4935);
nand U5011 (N_5011,N_4822,N_4841);
nand U5012 (N_5012,N_4910,N_4942);
and U5013 (N_5013,N_4811,N_4945);
nor U5014 (N_5014,N_4853,N_4824);
xor U5015 (N_5015,N_4897,N_4893);
xor U5016 (N_5016,N_4806,N_4821);
xnor U5017 (N_5017,N_4855,N_4833);
nor U5018 (N_5018,N_4836,N_4886);
nor U5019 (N_5019,N_4913,N_4818);
or U5020 (N_5020,N_4959,N_4917);
nand U5021 (N_5021,N_4820,N_4915);
or U5022 (N_5022,N_4880,N_4832);
xnor U5023 (N_5023,N_4837,N_4895);
xnor U5024 (N_5024,N_4861,N_4801);
and U5025 (N_5025,N_4916,N_4864);
xnor U5026 (N_5026,N_4918,N_4944);
nand U5027 (N_5027,N_4931,N_4933);
nor U5028 (N_5028,N_4854,N_4870);
xnor U5029 (N_5029,N_4938,N_4887);
xnor U5030 (N_5030,N_4802,N_4892);
nor U5031 (N_5031,N_4923,N_4827);
or U5032 (N_5032,N_4911,N_4890);
or U5033 (N_5033,N_4823,N_4956);
or U5034 (N_5034,N_4936,N_4926);
or U5035 (N_5035,N_4831,N_4950);
and U5036 (N_5036,N_4877,N_4882);
nor U5037 (N_5037,N_4871,N_4816);
and U5038 (N_5038,N_4888,N_4937);
xnor U5039 (N_5039,N_4920,N_4903);
xor U5040 (N_5040,N_4873,N_4924);
nor U5041 (N_5041,N_4922,N_4866);
or U5042 (N_5042,N_4813,N_4938);
nor U5043 (N_5043,N_4859,N_4921);
xnor U5044 (N_5044,N_4905,N_4856);
nor U5045 (N_5045,N_4924,N_4871);
nand U5046 (N_5046,N_4845,N_4849);
xnor U5047 (N_5047,N_4939,N_4919);
or U5048 (N_5048,N_4931,N_4926);
xnor U5049 (N_5049,N_4942,N_4892);
nor U5050 (N_5050,N_4862,N_4818);
xnor U5051 (N_5051,N_4843,N_4808);
nand U5052 (N_5052,N_4919,N_4874);
nand U5053 (N_5053,N_4902,N_4802);
or U5054 (N_5054,N_4812,N_4854);
or U5055 (N_5055,N_4946,N_4804);
xor U5056 (N_5056,N_4928,N_4952);
nand U5057 (N_5057,N_4884,N_4933);
nor U5058 (N_5058,N_4857,N_4851);
or U5059 (N_5059,N_4868,N_4801);
nand U5060 (N_5060,N_4939,N_4914);
or U5061 (N_5061,N_4885,N_4946);
and U5062 (N_5062,N_4811,N_4801);
xor U5063 (N_5063,N_4946,N_4819);
nand U5064 (N_5064,N_4879,N_4852);
xnor U5065 (N_5065,N_4920,N_4820);
and U5066 (N_5066,N_4951,N_4929);
nand U5067 (N_5067,N_4905,N_4880);
nand U5068 (N_5068,N_4805,N_4932);
nand U5069 (N_5069,N_4877,N_4863);
nand U5070 (N_5070,N_4904,N_4901);
xor U5071 (N_5071,N_4943,N_4922);
nor U5072 (N_5072,N_4870,N_4880);
nand U5073 (N_5073,N_4869,N_4826);
xor U5074 (N_5074,N_4921,N_4861);
and U5075 (N_5075,N_4917,N_4938);
nand U5076 (N_5076,N_4817,N_4904);
nand U5077 (N_5077,N_4871,N_4903);
or U5078 (N_5078,N_4911,N_4802);
xnor U5079 (N_5079,N_4820,N_4857);
and U5080 (N_5080,N_4899,N_4903);
nor U5081 (N_5081,N_4880,N_4946);
nor U5082 (N_5082,N_4824,N_4913);
nor U5083 (N_5083,N_4830,N_4924);
or U5084 (N_5084,N_4954,N_4816);
xnor U5085 (N_5085,N_4866,N_4939);
nor U5086 (N_5086,N_4888,N_4881);
or U5087 (N_5087,N_4894,N_4831);
xor U5088 (N_5088,N_4852,N_4800);
xor U5089 (N_5089,N_4922,N_4940);
nand U5090 (N_5090,N_4816,N_4951);
xor U5091 (N_5091,N_4858,N_4959);
or U5092 (N_5092,N_4890,N_4881);
xnor U5093 (N_5093,N_4856,N_4860);
nand U5094 (N_5094,N_4905,N_4921);
nor U5095 (N_5095,N_4856,N_4811);
and U5096 (N_5096,N_4831,N_4928);
and U5097 (N_5097,N_4886,N_4959);
nand U5098 (N_5098,N_4951,N_4874);
nor U5099 (N_5099,N_4949,N_4938);
and U5100 (N_5100,N_4942,N_4955);
nand U5101 (N_5101,N_4815,N_4939);
nor U5102 (N_5102,N_4847,N_4937);
nand U5103 (N_5103,N_4816,N_4844);
xnor U5104 (N_5104,N_4809,N_4896);
nand U5105 (N_5105,N_4802,N_4936);
and U5106 (N_5106,N_4885,N_4950);
or U5107 (N_5107,N_4860,N_4853);
or U5108 (N_5108,N_4862,N_4900);
nor U5109 (N_5109,N_4956,N_4953);
and U5110 (N_5110,N_4935,N_4931);
and U5111 (N_5111,N_4863,N_4816);
and U5112 (N_5112,N_4895,N_4852);
and U5113 (N_5113,N_4939,N_4910);
nor U5114 (N_5114,N_4928,N_4811);
nand U5115 (N_5115,N_4824,N_4919);
and U5116 (N_5116,N_4871,N_4918);
xnor U5117 (N_5117,N_4871,N_4875);
nor U5118 (N_5118,N_4881,N_4953);
nand U5119 (N_5119,N_4898,N_4838);
nand U5120 (N_5120,N_5048,N_5029);
xor U5121 (N_5121,N_4971,N_5014);
nor U5122 (N_5122,N_5106,N_5091);
xor U5123 (N_5123,N_5033,N_5026);
xor U5124 (N_5124,N_5018,N_5009);
and U5125 (N_5125,N_5101,N_4985);
or U5126 (N_5126,N_4975,N_5045);
xnor U5127 (N_5127,N_4982,N_5079);
nor U5128 (N_5128,N_5004,N_5052);
nor U5129 (N_5129,N_5050,N_5062);
and U5130 (N_5130,N_5070,N_5025);
and U5131 (N_5131,N_5035,N_4983);
and U5132 (N_5132,N_4963,N_4964);
xor U5133 (N_5133,N_5108,N_5042);
and U5134 (N_5134,N_5115,N_5080);
nand U5135 (N_5135,N_5051,N_5092);
and U5136 (N_5136,N_4968,N_5007);
and U5137 (N_5137,N_5107,N_4993);
or U5138 (N_5138,N_5093,N_5082);
nor U5139 (N_5139,N_5059,N_4994);
xor U5140 (N_5140,N_5038,N_4986);
nand U5141 (N_5141,N_5010,N_5077);
or U5142 (N_5142,N_4998,N_4979);
nor U5143 (N_5143,N_5008,N_5071);
nor U5144 (N_5144,N_5001,N_5020);
xnor U5145 (N_5145,N_5090,N_5023);
and U5146 (N_5146,N_5104,N_5072);
xnor U5147 (N_5147,N_5073,N_5114);
nand U5148 (N_5148,N_4996,N_5046);
xnor U5149 (N_5149,N_5064,N_4984);
nand U5150 (N_5150,N_5021,N_5099);
nor U5151 (N_5151,N_4980,N_5117);
or U5152 (N_5152,N_4967,N_4961);
nor U5153 (N_5153,N_5109,N_5089);
or U5154 (N_5154,N_5037,N_5016);
nand U5155 (N_5155,N_5030,N_5006);
and U5156 (N_5156,N_5031,N_5113);
nor U5157 (N_5157,N_4991,N_5118);
nand U5158 (N_5158,N_5061,N_5078);
nand U5159 (N_5159,N_5017,N_5103);
or U5160 (N_5160,N_5040,N_5024);
and U5161 (N_5161,N_4976,N_4977);
or U5162 (N_5162,N_5015,N_5000);
xor U5163 (N_5163,N_4969,N_5119);
nor U5164 (N_5164,N_5112,N_5067);
and U5165 (N_5165,N_5057,N_4988);
xor U5166 (N_5166,N_4973,N_4972);
and U5167 (N_5167,N_5027,N_5076);
or U5168 (N_5168,N_4970,N_5110);
nor U5169 (N_5169,N_5081,N_5098);
xor U5170 (N_5170,N_5083,N_5095);
nor U5171 (N_5171,N_4962,N_4966);
xor U5172 (N_5172,N_5039,N_4999);
xnor U5173 (N_5173,N_4978,N_5105);
or U5174 (N_5174,N_5075,N_5019);
nand U5175 (N_5175,N_5032,N_5111);
or U5176 (N_5176,N_5074,N_5013);
xnor U5177 (N_5177,N_4995,N_5066);
nor U5178 (N_5178,N_5058,N_5053);
xor U5179 (N_5179,N_4990,N_5049);
or U5180 (N_5180,N_5056,N_4987);
nor U5181 (N_5181,N_5116,N_5036);
and U5182 (N_5182,N_5096,N_5102);
nor U5183 (N_5183,N_4960,N_4997);
or U5184 (N_5184,N_5097,N_5086);
xor U5185 (N_5185,N_5044,N_4974);
nand U5186 (N_5186,N_5043,N_5047);
nor U5187 (N_5187,N_5055,N_5065);
xor U5188 (N_5188,N_5041,N_5012);
nand U5189 (N_5189,N_5094,N_5084);
or U5190 (N_5190,N_5063,N_5068);
nand U5191 (N_5191,N_4965,N_4989);
or U5192 (N_5192,N_5005,N_5011);
or U5193 (N_5193,N_5028,N_5022);
xor U5194 (N_5194,N_5034,N_5088);
xor U5195 (N_5195,N_5003,N_5002);
xor U5196 (N_5196,N_5060,N_5069);
xnor U5197 (N_5197,N_5087,N_5054);
nand U5198 (N_5198,N_4992,N_4981);
nor U5199 (N_5199,N_5085,N_5100);
and U5200 (N_5200,N_5077,N_4985);
xor U5201 (N_5201,N_5038,N_5021);
and U5202 (N_5202,N_5077,N_5030);
and U5203 (N_5203,N_4997,N_4975);
or U5204 (N_5204,N_5012,N_4999);
and U5205 (N_5205,N_5071,N_5029);
xor U5206 (N_5206,N_5095,N_5029);
xor U5207 (N_5207,N_5047,N_5073);
xnor U5208 (N_5208,N_5035,N_5075);
nand U5209 (N_5209,N_4994,N_5046);
nor U5210 (N_5210,N_5093,N_5100);
and U5211 (N_5211,N_5006,N_5013);
xor U5212 (N_5212,N_4969,N_5013);
nor U5213 (N_5213,N_4997,N_5082);
and U5214 (N_5214,N_5054,N_5069);
or U5215 (N_5215,N_5043,N_4976);
nor U5216 (N_5216,N_5065,N_5083);
and U5217 (N_5217,N_4984,N_4976);
or U5218 (N_5218,N_5093,N_5069);
xnor U5219 (N_5219,N_5098,N_5055);
nand U5220 (N_5220,N_5027,N_4966);
nand U5221 (N_5221,N_5017,N_5002);
and U5222 (N_5222,N_5065,N_5000);
xnor U5223 (N_5223,N_5062,N_5038);
nor U5224 (N_5224,N_4979,N_5053);
xor U5225 (N_5225,N_5034,N_5008);
or U5226 (N_5226,N_5040,N_5031);
xor U5227 (N_5227,N_4985,N_5010);
or U5228 (N_5228,N_5026,N_5071);
xor U5229 (N_5229,N_4981,N_4976);
and U5230 (N_5230,N_4989,N_5088);
or U5231 (N_5231,N_5069,N_5108);
nand U5232 (N_5232,N_5085,N_5018);
xnor U5233 (N_5233,N_4972,N_5072);
or U5234 (N_5234,N_5028,N_5077);
nor U5235 (N_5235,N_5012,N_5050);
or U5236 (N_5236,N_4966,N_4999);
or U5237 (N_5237,N_4991,N_5072);
nand U5238 (N_5238,N_5075,N_5027);
nor U5239 (N_5239,N_4988,N_5076);
nand U5240 (N_5240,N_4970,N_5031);
nand U5241 (N_5241,N_5033,N_5092);
xnor U5242 (N_5242,N_5038,N_5097);
nor U5243 (N_5243,N_4975,N_5009);
xor U5244 (N_5244,N_4995,N_5064);
nand U5245 (N_5245,N_5056,N_4975);
nand U5246 (N_5246,N_5082,N_5022);
and U5247 (N_5247,N_5092,N_4977);
nor U5248 (N_5248,N_4960,N_5078);
or U5249 (N_5249,N_5083,N_5036);
nor U5250 (N_5250,N_5059,N_5064);
or U5251 (N_5251,N_5080,N_4999);
or U5252 (N_5252,N_4996,N_5031);
and U5253 (N_5253,N_5115,N_4964);
xor U5254 (N_5254,N_5020,N_5024);
and U5255 (N_5255,N_5093,N_5114);
and U5256 (N_5256,N_5022,N_4979);
nor U5257 (N_5257,N_4961,N_5057);
xor U5258 (N_5258,N_5048,N_5052);
xnor U5259 (N_5259,N_5031,N_5010);
and U5260 (N_5260,N_5047,N_5057);
and U5261 (N_5261,N_5009,N_5081);
or U5262 (N_5262,N_5087,N_5075);
nor U5263 (N_5263,N_5073,N_5083);
and U5264 (N_5264,N_5007,N_4963);
and U5265 (N_5265,N_5052,N_5082);
nor U5266 (N_5266,N_4982,N_5063);
and U5267 (N_5267,N_5056,N_5061);
and U5268 (N_5268,N_5089,N_4990);
xnor U5269 (N_5269,N_5100,N_5094);
or U5270 (N_5270,N_5031,N_5117);
or U5271 (N_5271,N_4989,N_4984);
or U5272 (N_5272,N_5109,N_5008);
or U5273 (N_5273,N_5047,N_5011);
or U5274 (N_5274,N_5020,N_4999);
xnor U5275 (N_5275,N_5011,N_4974);
and U5276 (N_5276,N_4971,N_5040);
nor U5277 (N_5277,N_5007,N_5098);
nand U5278 (N_5278,N_5066,N_5067);
or U5279 (N_5279,N_5040,N_4997);
nor U5280 (N_5280,N_5145,N_5210);
and U5281 (N_5281,N_5257,N_5158);
and U5282 (N_5282,N_5196,N_5216);
and U5283 (N_5283,N_5156,N_5208);
xor U5284 (N_5284,N_5212,N_5134);
or U5285 (N_5285,N_5175,N_5231);
xor U5286 (N_5286,N_5150,N_5245);
xor U5287 (N_5287,N_5202,N_5143);
xor U5288 (N_5288,N_5181,N_5228);
and U5289 (N_5289,N_5203,N_5200);
xor U5290 (N_5290,N_5274,N_5130);
nand U5291 (N_5291,N_5224,N_5183);
xnor U5292 (N_5292,N_5180,N_5173);
and U5293 (N_5293,N_5213,N_5128);
or U5294 (N_5294,N_5138,N_5209);
xnor U5295 (N_5295,N_5243,N_5199);
or U5296 (N_5296,N_5148,N_5240);
or U5297 (N_5297,N_5265,N_5249);
nor U5298 (N_5298,N_5191,N_5162);
and U5299 (N_5299,N_5206,N_5258);
nand U5300 (N_5300,N_5169,N_5254);
nand U5301 (N_5301,N_5160,N_5253);
or U5302 (N_5302,N_5135,N_5272);
xor U5303 (N_5303,N_5126,N_5218);
nand U5304 (N_5304,N_5149,N_5230);
xor U5305 (N_5305,N_5262,N_5219);
and U5306 (N_5306,N_5174,N_5123);
and U5307 (N_5307,N_5211,N_5259);
nand U5308 (N_5308,N_5221,N_5263);
and U5309 (N_5309,N_5261,N_5185);
xnor U5310 (N_5310,N_5260,N_5251);
and U5311 (N_5311,N_5225,N_5141);
and U5312 (N_5312,N_5159,N_5131);
or U5313 (N_5313,N_5167,N_5176);
nand U5314 (N_5314,N_5255,N_5124);
xnor U5315 (N_5315,N_5279,N_5250);
or U5316 (N_5316,N_5151,N_5177);
nand U5317 (N_5317,N_5147,N_5195);
and U5318 (N_5318,N_5193,N_5188);
or U5319 (N_5319,N_5133,N_5222);
and U5320 (N_5320,N_5178,N_5121);
and U5321 (N_5321,N_5186,N_5152);
and U5322 (N_5322,N_5220,N_5217);
and U5323 (N_5323,N_5187,N_5248);
and U5324 (N_5324,N_5140,N_5223);
nor U5325 (N_5325,N_5125,N_5239);
nand U5326 (N_5326,N_5154,N_5215);
nand U5327 (N_5327,N_5242,N_5165);
xor U5328 (N_5328,N_5132,N_5236);
and U5329 (N_5329,N_5184,N_5157);
xor U5330 (N_5330,N_5146,N_5256);
or U5331 (N_5331,N_5198,N_5277);
xnor U5332 (N_5332,N_5172,N_5166);
xor U5333 (N_5333,N_5278,N_5275);
and U5334 (N_5334,N_5207,N_5170);
or U5335 (N_5335,N_5232,N_5182);
or U5336 (N_5336,N_5252,N_5204);
or U5337 (N_5337,N_5120,N_5247);
and U5338 (N_5338,N_5244,N_5136);
nand U5339 (N_5339,N_5234,N_5197);
or U5340 (N_5340,N_5189,N_5235);
and U5341 (N_5341,N_5139,N_5171);
xnor U5342 (N_5342,N_5142,N_5267);
or U5343 (N_5343,N_5194,N_5153);
or U5344 (N_5344,N_5168,N_5127);
nand U5345 (N_5345,N_5205,N_5155);
nand U5346 (N_5346,N_5129,N_5233);
or U5347 (N_5347,N_5273,N_5271);
xor U5348 (N_5348,N_5192,N_5179);
xor U5349 (N_5349,N_5214,N_5229);
nor U5350 (N_5350,N_5237,N_5276);
and U5351 (N_5351,N_5161,N_5268);
nand U5352 (N_5352,N_5190,N_5241);
xnor U5353 (N_5353,N_5246,N_5137);
xor U5354 (N_5354,N_5164,N_5201);
xnor U5355 (N_5355,N_5226,N_5144);
xnor U5356 (N_5356,N_5122,N_5270);
nand U5357 (N_5357,N_5264,N_5227);
xor U5358 (N_5358,N_5238,N_5269);
nand U5359 (N_5359,N_5266,N_5163);
xnor U5360 (N_5360,N_5253,N_5236);
or U5361 (N_5361,N_5123,N_5121);
and U5362 (N_5362,N_5129,N_5127);
nand U5363 (N_5363,N_5155,N_5240);
nand U5364 (N_5364,N_5190,N_5257);
nor U5365 (N_5365,N_5146,N_5169);
xnor U5366 (N_5366,N_5160,N_5125);
nor U5367 (N_5367,N_5235,N_5233);
xor U5368 (N_5368,N_5151,N_5132);
or U5369 (N_5369,N_5164,N_5235);
xor U5370 (N_5370,N_5271,N_5263);
and U5371 (N_5371,N_5223,N_5251);
and U5372 (N_5372,N_5265,N_5221);
nor U5373 (N_5373,N_5125,N_5143);
nand U5374 (N_5374,N_5215,N_5272);
or U5375 (N_5375,N_5232,N_5222);
or U5376 (N_5376,N_5223,N_5239);
xnor U5377 (N_5377,N_5263,N_5192);
nor U5378 (N_5378,N_5124,N_5168);
or U5379 (N_5379,N_5125,N_5142);
xnor U5380 (N_5380,N_5226,N_5231);
nand U5381 (N_5381,N_5181,N_5175);
and U5382 (N_5382,N_5224,N_5196);
and U5383 (N_5383,N_5128,N_5148);
nand U5384 (N_5384,N_5128,N_5176);
nor U5385 (N_5385,N_5195,N_5223);
and U5386 (N_5386,N_5180,N_5221);
and U5387 (N_5387,N_5214,N_5159);
xnor U5388 (N_5388,N_5253,N_5234);
and U5389 (N_5389,N_5268,N_5279);
nor U5390 (N_5390,N_5184,N_5126);
and U5391 (N_5391,N_5260,N_5120);
and U5392 (N_5392,N_5126,N_5140);
xnor U5393 (N_5393,N_5192,N_5150);
or U5394 (N_5394,N_5129,N_5199);
nor U5395 (N_5395,N_5244,N_5237);
and U5396 (N_5396,N_5174,N_5233);
xor U5397 (N_5397,N_5261,N_5196);
nand U5398 (N_5398,N_5158,N_5183);
nand U5399 (N_5399,N_5188,N_5222);
nor U5400 (N_5400,N_5126,N_5249);
xnor U5401 (N_5401,N_5197,N_5248);
xnor U5402 (N_5402,N_5189,N_5201);
and U5403 (N_5403,N_5216,N_5274);
nand U5404 (N_5404,N_5199,N_5258);
xor U5405 (N_5405,N_5120,N_5154);
or U5406 (N_5406,N_5258,N_5121);
xnor U5407 (N_5407,N_5269,N_5208);
nor U5408 (N_5408,N_5258,N_5142);
or U5409 (N_5409,N_5139,N_5277);
xnor U5410 (N_5410,N_5146,N_5183);
nand U5411 (N_5411,N_5163,N_5170);
nor U5412 (N_5412,N_5246,N_5164);
nor U5413 (N_5413,N_5133,N_5189);
and U5414 (N_5414,N_5131,N_5181);
xor U5415 (N_5415,N_5196,N_5187);
nor U5416 (N_5416,N_5255,N_5136);
xnor U5417 (N_5417,N_5277,N_5226);
nand U5418 (N_5418,N_5165,N_5273);
nor U5419 (N_5419,N_5159,N_5144);
nand U5420 (N_5420,N_5215,N_5222);
nand U5421 (N_5421,N_5180,N_5124);
nand U5422 (N_5422,N_5189,N_5126);
and U5423 (N_5423,N_5128,N_5129);
nand U5424 (N_5424,N_5162,N_5249);
and U5425 (N_5425,N_5154,N_5136);
or U5426 (N_5426,N_5278,N_5138);
nand U5427 (N_5427,N_5131,N_5129);
xnor U5428 (N_5428,N_5137,N_5179);
nand U5429 (N_5429,N_5125,N_5242);
and U5430 (N_5430,N_5123,N_5277);
xnor U5431 (N_5431,N_5218,N_5135);
nand U5432 (N_5432,N_5162,N_5189);
xor U5433 (N_5433,N_5161,N_5263);
nand U5434 (N_5434,N_5195,N_5275);
and U5435 (N_5435,N_5251,N_5124);
and U5436 (N_5436,N_5172,N_5156);
nand U5437 (N_5437,N_5140,N_5231);
nand U5438 (N_5438,N_5184,N_5233);
xnor U5439 (N_5439,N_5231,N_5203);
nand U5440 (N_5440,N_5398,N_5389);
or U5441 (N_5441,N_5325,N_5355);
nor U5442 (N_5442,N_5312,N_5302);
xor U5443 (N_5443,N_5284,N_5315);
nand U5444 (N_5444,N_5421,N_5333);
and U5445 (N_5445,N_5310,N_5380);
or U5446 (N_5446,N_5434,N_5290);
xor U5447 (N_5447,N_5388,N_5344);
or U5448 (N_5448,N_5385,N_5306);
nand U5449 (N_5449,N_5322,N_5350);
nand U5450 (N_5450,N_5349,N_5301);
nand U5451 (N_5451,N_5309,N_5362);
nor U5452 (N_5452,N_5416,N_5413);
xnor U5453 (N_5453,N_5293,N_5436);
nand U5454 (N_5454,N_5289,N_5294);
nor U5455 (N_5455,N_5299,N_5390);
or U5456 (N_5456,N_5336,N_5298);
xor U5457 (N_5457,N_5427,N_5366);
xnor U5458 (N_5458,N_5381,N_5324);
nand U5459 (N_5459,N_5411,N_5394);
nor U5460 (N_5460,N_5430,N_5297);
and U5461 (N_5461,N_5348,N_5371);
nand U5462 (N_5462,N_5410,N_5435);
or U5463 (N_5463,N_5401,N_5425);
or U5464 (N_5464,N_5281,N_5424);
and U5465 (N_5465,N_5379,N_5339);
xor U5466 (N_5466,N_5437,N_5288);
and U5467 (N_5467,N_5419,N_5395);
and U5468 (N_5468,N_5342,N_5300);
and U5469 (N_5469,N_5351,N_5354);
nand U5470 (N_5470,N_5326,N_5418);
and U5471 (N_5471,N_5353,N_5327);
or U5472 (N_5472,N_5358,N_5318);
or U5473 (N_5473,N_5340,N_5432);
nand U5474 (N_5474,N_5343,N_5397);
and U5475 (N_5475,N_5374,N_5357);
and U5476 (N_5476,N_5305,N_5408);
xnor U5477 (N_5477,N_5337,N_5363);
xor U5478 (N_5478,N_5328,N_5316);
xnor U5479 (N_5479,N_5378,N_5431);
nand U5480 (N_5480,N_5313,N_5311);
or U5481 (N_5481,N_5417,N_5283);
nor U5482 (N_5482,N_5341,N_5286);
nand U5483 (N_5483,N_5399,N_5314);
nor U5484 (N_5484,N_5422,N_5376);
nor U5485 (N_5485,N_5345,N_5308);
or U5486 (N_5486,N_5438,N_5368);
or U5487 (N_5487,N_5365,N_5404);
nand U5488 (N_5488,N_5393,N_5383);
xor U5489 (N_5489,N_5295,N_5321);
and U5490 (N_5490,N_5356,N_5361);
xor U5491 (N_5491,N_5375,N_5396);
nor U5492 (N_5492,N_5420,N_5287);
and U5493 (N_5493,N_5377,N_5303);
or U5494 (N_5494,N_5414,N_5439);
or U5495 (N_5495,N_5415,N_5307);
or U5496 (N_5496,N_5359,N_5406);
nand U5497 (N_5497,N_5373,N_5292);
nand U5498 (N_5498,N_5372,N_5347);
and U5499 (N_5499,N_5402,N_5291);
xnor U5500 (N_5500,N_5285,N_5391);
nor U5501 (N_5501,N_5405,N_5382);
xor U5502 (N_5502,N_5320,N_5407);
nor U5503 (N_5503,N_5329,N_5352);
xor U5504 (N_5504,N_5360,N_5334);
and U5505 (N_5505,N_5412,N_5282);
and U5506 (N_5506,N_5319,N_5384);
or U5507 (N_5507,N_5280,N_5296);
xor U5508 (N_5508,N_5433,N_5304);
nor U5509 (N_5509,N_5409,N_5338);
or U5510 (N_5510,N_5370,N_5426);
nor U5511 (N_5511,N_5387,N_5330);
or U5512 (N_5512,N_5332,N_5331);
or U5513 (N_5513,N_5367,N_5369);
or U5514 (N_5514,N_5428,N_5403);
or U5515 (N_5515,N_5386,N_5392);
nand U5516 (N_5516,N_5335,N_5400);
and U5517 (N_5517,N_5423,N_5364);
xor U5518 (N_5518,N_5429,N_5323);
nor U5519 (N_5519,N_5317,N_5346);
or U5520 (N_5520,N_5317,N_5323);
nor U5521 (N_5521,N_5349,N_5281);
and U5522 (N_5522,N_5327,N_5378);
nand U5523 (N_5523,N_5427,N_5344);
nand U5524 (N_5524,N_5432,N_5303);
xnor U5525 (N_5525,N_5430,N_5375);
or U5526 (N_5526,N_5357,N_5372);
or U5527 (N_5527,N_5384,N_5325);
nor U5528 (N_5528,N_5338,N_5397);
nor U5529 (N_5529,N_5325,N_5420);
or U5530 (N_5530,N_5329,N_5368);
nand U5531 (N_5531,N_5371,N_5294);
nand U5532 (N_5532,N_5337,N_5372);
or U5533 (N_5533,N_5320,N_5390);
xnor U5534 (N_5534,N_5436,N_5281);
nor U5535 (N_5535,N_5353,N_5384);
and U5536 (N_5536,N_5286,N_5365);
nand U5537 (N_5537,N_5392,N_5383);
nand U5538 (N_5538,N_5353,N_5368);
xnor U5539 (N_5539,N_5368,N_5330);
xor U5540 (N_5540,N_5327,N_5338);
or U5541 (N_5541,N_5308,N_5396);
or U5542 (N_5542,N_5302,N_5415);
nand U5543 (N_5543,N_5425,N_5341);
nand U5544 (N_5544,N_5417,N_5294);
and U5545 (N_5545,N_5425,N_5329);
nand U5546 (N_5546,N_5414,N_5400);
and U5547 (N_5547,N_5428,N_5384);
nor U5548 (N_5548,N_5432,N_5349);
and U5549 (N_5549,N_5371,N_5301);
xnor U5550 (N_5550,N_5383,N_5362);
and U5551 (N_5551,N_5439,N_5315);
nor U5552 (N_5552,N_5396,N_5382);
xor U5553 (N_5553,N_5309,N_5363);
nor U5554 (N_5554,N_5407,N_5311);
xor U5555 (N_5555,N_5299,N_5372);
and U5556 (N_5556,N_5407,N_5431);
nor U5557 (N_5557,N_5282,N_5289);
nor U5558 (N_5558,N_5355,N_5362);
xor U5559 (N_5559,N_5428,N_5390);
and U5560 (N_5560,N_5424,N_5407);
nor U5561 (N_5561,N_5367,N_5392);
nand U5562 (N_5562,N_5346,N_5367);
xor U5563 (N_5563,N_5417,N_5321);
nor U5564 (N_5564,N_5424,N_5318);
and U5565 (N_5565,N_5389,N_5294);
or U5566 (N_5566,N_5285,N_5407);
nor U5567 (N_5567,N_5394,N_5367);
and U5568 (N_5568,N_5401,N_5413);
xor U5569 (N_5569,N_5372,N_5331);
and U5570 (N_5570,N_5430,N_5332);
nor U5571 (N_5571,N_5342,N_5307);
xor U5572 (N_5572,N_5284,N_5379);
or U5573 (N_5573,N_5338,N_5301);
or U5574 (N_5574,N_5375,N_5344);
xor U5575 (N_5575,N_5405,N_5290);
or U5576 (N_5576,N_5381,N_5368);
and U5577 (N_5577,N_5369,N_5348);
and U5578 (N_5578,N_5347,N_5420);
xor U5579 (N_5579,N_5364,N_5306);
or U5580 (N_5580,N_5418,N_5317);
nand U5581 (N_5581,N_5351,N_5310);
or U5582 (N_5582,N_5359,N_5429);
nor U5583 (N_5583,N_5427,N_5429);
xor U5584 (N_5584,N_5359,N_5343);
and U5585 (N_5585,N_5398,N_5356);
xor U5586 (N_5586,N_5308,N_5408);
xor U5587 (N_5587,N_5437,N_5293);
and U5588 (N_5588,N_5354,N_5435);
nor U5589 (N_5589,N_5286,N_5428);
nand U5590 (N_5590,N_5374,N_5315);
xor U5591 (N_5591,N_5409,N_5421);
nor U5592 (N_5592,N_5413,N_5360);
nor U5593 (N_5593,N_5413,N_5370);
or U5594 (N_5594,N_5409,N_5343);
nand U5595 (N_5595,N_5359,N_5370);
or U5596 (N_5596,N_5395,N_5413);
or U5597 (N_5597,N_5301,N_5395);
and U5598 (N_5598,N_5411,N_5437);
xor U5599 (N_5599,N_5320,N_5381);
or U5600 (N_5600,N_5501,N_5557);
or U5601 (N_5601,N_5456,N_5593);
nand U5602 (N_5602,N_5475,N_5591);
or U5603 (N_5603,N_5527,N_5549);
or U5604 (N_5604,N_5493,N_5505);
and U5605 (N_5605,N_5490,N_5486);
xor U5606 (N_5606,N_5440,N_5455);
and U5607 (N_5607,N_5482,N_5503);
or U5608 (N_5608,N_5507,N_5592);
nand U5609 (N_5609,N_5524,N_5464);
or U5610 (N_5610,N_5515,N_5570);
nand U5611 (N_5611,N_5444,N_5536);
nor U5612 (N_5612,N_5573,N_5574);
and U5613 (N_5613,N_5467,N_5509);
or U5614 (N_5614,N_5492,N_5458);
or U5615 (N_5615,N_5508,N_5471);
or U5616 (N_5616,N_5531,N_5586);
xor U5617 (N_5617,N_5541,N_5452);
or U5618 (N_5618,N_5518,N_5495);
nor U5619 (N_5619,N_5576,N_5597);
xor U5620 (N_5620,N_5489,N_5584);
nor U5621 (N_5621,N_5529,N_5583);
xnor U5622 (N_5622,N_5460,N_5564);
and U5623 (N_5623,N_5555,N_5550);
nor U5624 (N_5624,N_5533,N_5551);
xor U5625 (N_5625,N_5449,N_5517);
nand U5626 (N_5626,N_5498,N_5461);
nand U5627 (N_5627,N_5512,N_5578);
xor U5628 (N_5628,N_5445,N_5559);
or U5629 (N_5629,N_5588,N_5441);
xnor U5630 (N_5630,N_5554,N_5526);
or U5631 (N_5631,N_5469,N_5568);
or U5632 (N_5632,N_5521,N_5539);
xor U5633 (N_5633,N_5480,N_5580);
nor U5634 (N_5634,N_5497,N_5514);
xnor U5635 (N_5635,N_5553,N_5516);
xnor U5636 (N_5636,N_5532,N_5589);
nand U5637 (N_5637,N_5544,N_5547);
nand U5638 (N_5638,N_5499,N_5511);
and U5639 (N_5639,N_5537,N_5459);
and U5640 (N_5640,N_5462,N_5535);
and U5641 (N_5641,N_5479,N_5569);
nand U5642 (N_5642,N_5481,N_5513);
or U5643 (N_5643,N_5447,N_5470);
nand U5644 (N_5644,N_5562,N_5540);
nand U5645 (N_5645,N_5478,N_5504);
and U5646 (N_5646,N_5494,N_5487);
nor U5647 (N_5647,N_5594,N_5457);
xnor U5648 (N_5648,N_5477,N_5561);
and U5649 (N_5649,N_5571,N_5476);
or U5650 (N_5650,N_5484,N_5448);
xor U5651 (N_5651,N_5523,N_5563);
nand U5652 (N_5652,N_5542,N_5528);
or U5653 (N_5653,N_5587,N_5510);
and U5654 (N_5654,N_5543,N_5585);
and U5655 (N_5655,N_5546,N_5519);
xor U5656 (N_5656,N_5582,N_5572);
nor U5657 (N_5657,N_5520,N_5558);
nor U5658 (N_5658,N_5453,N_5500);
or U5659 (N_5659,N_5560,N_5552);
or U5660 (N_5660,N_5483,N_5556);
xnor U5661 (N_5661,N_5506,N_5496);
xnor U5662 (N_5662,N_5522,N_5567);
nor U5663 (N_5663,N_5488,N_5565);
nand U5664 (N_5664,N_5525,N_5474);
nor U5665 (N_5665,N_5596,N_5485);
and U5666 (N_5666,N_5566,N_5442);
and U5667 (N_5667,N_5468,N_5598);
nor U5668 (N_5668,N_5545,N_5463);
or U5669 (N_5669,N_5530,N_5443);
nor U5670 (N_5670,N_5473,N_5575);
or U5671 (N_5671,N_5450,N_5590);
or U5672 (N_5672,N_5534,N_5451);
xnor U5673 (N_5673,N_5579,N_5472);
or U5674 (N_5674,N_5581,N_5502);
nand U5675 (N_5675,N_5446,N_5454);
nor U5676 (N_5676,N_5599,N_5466);
and U5677 (N_5677,N_5538,N_5548);
and U5678 (N_5678,N_5595,N_5465);
and U5679 (N_5679,N_5577,N_5491);
and U5680 (N_5680,N_5451,N_5502);
nand U5681 (N_5681,N_5545,N_5522);
nor U5682 (N_5682,N_5529,N_5491);
nand U5683 (N_5683,N_5461,N_5492);
xor U5684 (N_5684,N_5500,N_5542);
nor U5685 (N_5685,N_5563,N_5588);
nand U5686 (N_5686,N_5450,N_5442);
and U5687 (N_5687,N_5513,N_5467);
and U5688 (N_5688,N_5500,N_5494);
nand U5689 (N_5689,N_5457,N_5463);
nor U5690 (N_5690,N_5569,N_5544);
nand U5691 (N_5691,N_5592,N_5512);
nor U5692 (N_5692,N_5557,N_5583);
nor U5693 (N_5693,N_5441,N_5461);
nor U5694 (N_5694,N_5566,N_5552);
nor U5695 (N_5695,N_5483,N_5532);
nand U5696 (N_5696,N_5474,N_5578);
nor U5697 (N_5697,N_5497,N_5512);
nor U5698 (N_5698,N_5474,N_5469);
xor U5699 (N_5699,N_5461,N_5478);
nand U5700 (N_5700,N_5578,N_5486);
and U5701 (N_5701,N_5479,N_5481);
nand U5702 (N_5702,N_5504,N_5562);
xnor U5703 (N_5703,N_5537,N_5598);
or U5704 (N_5704,N_5502,N_5560);
nor U5705 (N_5705,N_5469,N_5484);
nor U5706 (N_5706,N_5501,N_5563);
nand U5707 (N_5707,N_5593,N_5567);
or U5708 (N_5708,N_5492,N_5519);
nor U5709 (N_5709,N_5463,N_5517);
nand U5710 (N_5710,N_5543,N_5444);
nand U5711 (N_5711,N_5453,N_5458);
xnor U5712 (N_5712,N_5528,N_5505);
nand U5713 (N_5713,N_5519,N_5594);
and U5714 (N_5714,N_5578,N_5484);
nor U5715 (N_5715,N_5513,N_5559);
xor U5716 (N_5716,N_5452,N_5489);
and U5717 (N_5717,N_5584,N_5552);
nand U5718 (N_5718,N_5539,N_5514);
nand U5719 (N_5719,N_5454,N_5511);
or U5720 (N_5720,N_5592,N_5447);
and U5721 (N_5721,N_5458,N_5510);
nand U5722 (N_5722,N_5489,N_5589);
nand U5723 (N_5723,N_5487,N_5477);
and U5724 (N_5724,N_5575,N_5468);
nor U5725 (N_5725,N_5488,N_5566);
xor U5726 (N_5726,N_5559,N_5599);
and U5727 (N_5727,N_5519,N_5467);
and U5728 (N_5728,N_5490,N_5592);
or U5729 (N_5729,N_5459,N_5553);
nand U5730 (N_5730,N_5535,N_5509);
or U5731 (N_5731,N_5579,N_5471);
nand U5732 (N_5732,N_5468,N_5559);
nand U5733 (N_5733,N_5578,N_5493);
and U5734 (N_5734,N_5594,N_5495);
xnor U5735 (N_5735,N_5563,N_5456);
xor U5736 (N_5736,N_5518,N_5461);
nor U5737 (N_5737,N_5451,N_5582);
nor U5738 (N_5738,N_5533,N_5497);
xnor U5739 (N_5739,N_5476,N_5470);
xor U5740 (N_5740,N_5563,N_5477);
nand U5741 (N_5741,N_5442,N_5588);
or U5742 (N_5742,N_5527,N_5475);
and U5743 (N_5743,N_5548,N_5480);
nor U5744 (N_5744,N_5451,N_5468);
or U5745 (N_5745,N_5510,N_5450);
nor U5746 (N_5746,N_5464,N_5562);
or U5747 (N_5747,N_5575,N_5480);
nand U5748 (N_5748,N_5491,N_5469);
nand U5749 (N_5749,N_5488,N_5480);
nand U5750 (N_5750,N_5526,N_5563);
xor U5751 (N_5751,N_5473,N_5502);
xor U5752 (N_5752,N_5516,N_5507);
nor U5753 (N_5753,N_5462,N_5518);
xor U5754 (N_5754,N_5443,N_5491);
nand U5755 (N_5755,N_5522,N_5596);
and U5756 (N_5756,N_5517,N_5578);
and U5757 (N_5757,N_5473,N_5464);
nor U5758 (N_5758,N_5564,N_5492);
nor U5759 (N_5759,N_5495,N_5569);
nor U5760 (N_5760,N_5690,N_5711);
nand U5761 (N_5761,N_5741,N_5727);
nor U5762 (N_5762,N_5616,N_5662);
and U5763 (N_5763,N_5730,N_5719);
and U5764 (N_5764,N_5679,N_5649);
nand U5765 (N_5765,N_5626,N_5706);
nand U5766 (N_5766,N_5735,N_5695);
nor U5767 (N_5767,N_5731,N_5618);
nand U5768 (N_5768,N_5652,N_5702);
xor U5769 (N_5769,N_5755,N_5605);
nor U5770 (N_5770,N_5659,N_5705);
and U5771 (N_5771,N_5632,N_5606);
or U5772 (N_5772,N_5749,N_5712);
and U5773 (N_5773,N_5740,N_5726);
and U5774 (N_5774,N_5674,N_5642);
or U5775 (N_5775,N_5658,N_5713);
nand U5776 (N_5776,N_5694,N_5654);
nand U5777 (N_5777,N_5700,N_5720);
xor U5778 (N_5778,N_5640,N_5644);
nand U5779 (N_5779,N_5672,N_5663);
nor U5780 (N_5780,N_5756,N_5624);
or U5781 (N_5781,N_5667,N_5688);
nand U5782 (N_5782,N_5691,N_5692);
nand U5783 (N_5783,N_5738,N_5607);
or U5784 (N_5784,N_5603,N_5609);
and U5785 (N_5785,N_5707,N_5634);
xnor U5786 (N_5786,N_5612,N_5724);
or U5787 (N_5787,N_5699,N_5664);
xor U5788 (N_5788,N_5710,N_5601);
nor U5789 (N_5789,N_5752,N_5701);
nor U5790 (N_5790,N_5647,N_5758);
xor U5791 (N_5791,N_5641,N_5717);
nor U5792 (N_5792,N_5681,N_5665);
and U5793 (N_5793,N_5604,N_5716);
and U5794 (N_5794,N_5636,N_5709);
xnor U5795 (N_5795,N_5668,N_5677);
xor U5796 (N_5796,N_5683,N_5620);
nor U5797 (N_5797,N_5734,N_5638);
and U5798 (N_5798,N_5622,N_5685);
or U5799 (N_5799,N_5715,N_5610);
nor U5800 (N_5800,N_5746,N_5613);
or U5801 (N_5801,N_5725,N_5687);
nor U5802 (N_5802,N_5703,N_5635);
xnor U5803 (N_5803,N_5625,N_5729);
or U5804 (N_5804,N_5660,N_5619);
nand U5805 (N_5805,N_5669,N_5682);
or U5806 (N_5806,N_5637,N_5708);
xor U5807 (N_5807,N_5739,N_5615);
xor U5808 (N_5808,N_5748,N_5743);
nand U5809 (N_5809,N_5721,N_5627);
nor U5810 (N_5810,N_5611,N_5600);
and U5811 (N_5811,N_5678,N_5675);
xnor U5812 (N_5812,N_5666,N_5754);
xor U5813 (N_5813,N_5623,N_5621);
or U5814 (N_5814,N_5653,N_5655);
nor U5815 (N_5815,N_5643,N_5757);
or U5816 (N_5816,N_5745,N_5733);
and U5817 (N_5817,N_5744,N_5670);
or U5818 (N_5818,N_5686,N_5608);
nor U5819 (N_5819,N_5656,N_5673);
nor U5820 (N_5820,N_5617,N_5718);
nand U5821 (N_5821,N_5639,N_5714);
xor U5822 (N_5822,N_5645,N_5657);
xnor U5823 (N_5823,N_5629,N_5747);
xor U5824 (N_5824,N_5696,N_5602);
or U5825 (N_5825,N_5751,N_5737);
xnor U5826 (N_5826,N_5698,N_5728);
nand U5827 (N_5827,N_5753,N_5680);
and U5828 (N_5828,N_5628,N_5722);
nand U5829 (N_5829,N_5661,N_5732);
nand U5830 (N_5830,N_5676,N_5614);
or U5831 (N_5831,N_5723,N_5689);
nand U5832 (N_5832,N_5704,N_5633);
and U5833 (N_5833,N_5736,N_5684);
and U5834 (N_5834,N_5671,N_5646);
nand U5835 (N_5835,N_5651,N_5631);
or U5836 (N_5836,N_5693,N_5742);
xnor U5837 (N_5837,N_5650,N_5759);
nor U5838 (N_5838,N_5648,N_5697);
nand U5839 (N_5839,N_5630,N_5750);
or U5840 (N_5840,N_5677,N_5750);
xnor U5841 (N_5841,N_5687,N_5604);
nand U5842 (N_5842,N_5689,N_5710);
and U5843 (N_5843,N_5685,N_5647);
and U5844 (N_5844,N_5674,N_5656);
nor U5845 (N_5845,N_5651,N_5757);
xor U5846 (N_5846,N_5708,N_5681);
or U5847 (N_5847,N_5671,N_5716);
nand U5848 (N_5848,N_5654,N_5627);
and U5849 (N_5849,N_5690,N_5688);
nand U5850 (N_5850,N_5647,N_5602);
xor U5851 (N_5851,N_5615,N_5606);
and U5852 (N_5852,N_5621,N_5699);
nor U5853 (N_5853,N_5686,N_5742);
nand U5854 (N_5854,N_5740,N_5678);
nor U5855 (N_5855,N_5638,N_5691);
nor U5856 (N_5856,N_5686,N_5616);
xor U5857 (N_5857,N_5684,N_5643);
nand U5858 (N_5858,N_5740,N_5701);
xnor U5859 (N_5859,N_5685,N_5752);
nand U5860 (N_5860,N_5695,N_5622);
nand U5861 (N_5861,N_5679,N_5701);
nor U5862 (N_5862,N_5725,N_5638);
nand U5863 (N_5863,N_5685,N_5601);
or U5864 (N_5864,N_5719,N_5654);
nand U5865 (N_5865,N_5710,N_5728);
nand U5866 (N_5866,N_5664,N_5645);
nand U5867 (N_5867,N_5605,N_5646);
xnor U5868 (N_5868,N_5727,N_5700);
nor U5869 (N_5869,N_5656,N_5758);
nor U5870 (N_5870,N_5712,N_5669);
and U5871 (N_5871,N_5677,N_5659);
and U5872 (N_5872,N_5733,N_5759);
and U5873 (N_5873,N_5752,N_5726);
and U5874 (N_5874,N_5726,N_5623);
nor U5875 (N_5875,N_5669,N_5664);
nand U5876 (N_5876,N_5738,N_5630);
and U5877 (N_5877,N_5672,N_5667);
xor U5878 (N_5878,N_5614,N_5610);
or U5879 (N_5879,N_5694,N_5665);
and U5880 (N_5880,N_5620,N_5676);
nand U5881 (N_5881,N_5687,N_5703);
xor U5882 (N_5882,N_5699,N_5644);
nor U5883 (N_5883,N_5621,N_5725);
xnor U5884 (N_5884,N_5684,N_5747);
xor U5885 (N_5885,N_5641,N_5670);
nor U5886 (N_5886,N_5659,N_5710);
or U5887 (N_5887,N_5640,N_5611);
xnor U5888 (N_5888,N_5618,N_5703);
or U5889 (N_5889,N_5709,N_5697);
or U5890 (N_5890,N_5642,N_5635);
xor U5891 (N_5891,N_5647,N_5754);
nand U5892 (N_5892,N_5704,N_5701);
nand U5893 (N_5893,N_5613,N_5605);
xnor U5894 (N_5894,N_5605,N_5602);
xor U5895 (N_5895,N_5647,N_5713);
xor U5896 (N_5896,N_5646,N_5743);
and U5897 (N_5897,N_5686,N_5610);
xnor U5898 (N_5898,N_5611,N_5693);
nand U5899 (N_5899,N_5662,N_5647);
nand U5900 (N_5900,N_5705,N_5681);
or U5901 (N_5901,N_5741,N_5756);
nor U5902 (N_5902,N_5697,N_5748);
nor U5903 (N_5903,N_5658,N_5719);
and U5904 (N_5904,N_5750,N_5703);
or U5905 (N_5905,N_5623,N_5740);
or U5906 (N_5906,N_5658,N_5644);
xnor U5907 (N_5907,N_5616,N_5613);
nor U5908 (N_5908,N_5682,N_5661);
or U5909 (N_5909,N_5653,N_5696);
or U5910 (N_5910,N_5624,N_5654);
xor U5911 (N_5911,N_5661,N_5692);
and U5912 (N_5912,N_5672,N_5644);
or U5913 (N_5913,N_5639,N_5666);
or U5914 (N_5914,N_5701,N_5705);
or U5915 (N_5915,N_5646,N_5659);
and U5916 (N_5916,N_5696,N_5735);
and U5917 (N_5917,N_5741,N_5604);
nor U5918 (N_5918,N_5699,N_5666);
nor U5919 (N_5919,N_5643,N_5724);
or U5920 (N_5920,N_5880,N_5826);
nor U5921 (N_5921,N_5893,N_5905);
and U5922 (N_5922,N_5868,N_5918);
nor U5923 (N_5923,N_5782,N_5803);
and U5924 (N_5924,N_5859,N_5879);
xnor U5925 (N_5925,N_5854,N_5769);
nor U5926 (N_5926,N_5786,N_5773);
and U5927 (N_5927,N_5915,N_5874);
nand U5928 (N_5928,N_5800,N_5873);
and U5929 (N_5929,N_5876,N_5855);
xor U5930 (N_5930,N_5818,N_5878);
and U5931 (N_5931,N_5914,N_5793);
nand U5932 (N_5932,N_5821,N_5767);
or U5933 (N_5933,N_5892,N_5819);
and U5934 (N_5934,N_5822,N_5775);
or U5935 (N_5935,N_5771,N_5815);
or U5936 (N_5936,N_5852,N_5788);
xor U5937 (N_5937,N_5898,N_5804);
xnor U5938 (N_5938,N_5789,N_5849);
nand U5939 (N_5939,N_5816,N_5882);
xor U5940 (N_5940,N_5838,N_5864);
and U5941 (N_5941,N_5802,N_5772);
or U5942 (N_5942,N_5825,N_5865);
or U5943 (N_5943,N_5843,N_5835);
nor U5944 (N_5944,N_5763,N_5853);
or U5945 (N_5945,N_5834,N_5888);
and U5946 (N_5946,N_5841,N_5850);
nand U5947 (N_5947,N_5883,N_5886);
and U5948 (N_5948,N_5832,N_5877);
or U5949 (N_5949,N_5761,N_5768);
and U5950 (N_5950,N_5848,N_5790);
or U5951 (N_5951,N_5817,N_5894);
nor U5952 (N_5952,N_5779,N_5907);
nand U5953 (N_5953,N_5828,N_5829);
nor U5954 (N_5954,N_5799,N_5766);
nor U5955 (N_5955,N_5846,N_5913);
xor U5956 (N_5956,N_5858,N_5807);
or U5957 (N_5957,N_5885,N_5871);
nor U5958 (N_5958,N_5806,N_5856);
or U5959 (N_5959,N_5770,N_5809);
or U5960 (N_5960,N_5774,N_5798);
and U5961 (N_5961,N_5824,N_5862);
nand U5962 (N_5962,N_5830,N_5794);
nand U5963 (N_5963,N_5884,N_5797);
nor U5964 (N_5964,N_5792,N_5881);
and U5965 (N_5965,N_5764,N_5777);
and U5966 (N_5966,N_5762,N_5908);
nor U5967 (N_5967,N_5904,N_5901);
nor U5968 (N_5968,N_5903,N_5900);
xor U5969 (N_5969,N_5776,N_5795);
nor U5970 (N_5970,N_5805,N_5781);
nand U5971 (N_5971,N_5840,N_5785);
or U5972 (N_5972,N_5813,N_5827);
and U5973 (N_5973,N_5895,N_5870);
and U5974 (N_5974,N_5796,N_5872);
and U5975 (N_5975,N_5814,N_5845);
nand U5976 (N_5976,N_5787,N_5866);
xor U5977 (N_5977,N_5844,N_5897);
or U5978 (N_5978,N_5860,N_5891);
xnor U5979 (N_5979,N_5812,N_5791);
and U5980 (N_5980,N_5875,N_5811);
or U5981 (N_5981,N_5760,N_5833);
nand U5982 (N_5982,N_5911,N_5863);
or U5983 (N_5983,N_5906,N_5837);
or U5984 (N_5984,N_5783,N_5851);
xor U5985 (N_5985,N_5836,N_5896);
xor U5986 (N_5986,N_5823,N_5857);
or U5987 (N_5987,N_5869,N_5765);
and U5988 (N_5988,N_5808,N_5917);
or U5989 (N_5989,N_5887,N_5839);
xnor U5990 (N_5990,N_5910,N_5890);
or U5991 (N_5991,N_5801,N_5778);
xor U5992 (N_5992,N_5867,N_5847);
xor U5993 (N_5993,N_5909,N_5919);
xnor U5994 (N_5994,N_5842,N_5820);
xnor U5995 (N_5995,N_5861,N_5831);
xor U5996 (N_5996,N_5780,N_5916);
xor U5997 (N_5997,N_5912,N_5889);
nor U5998 (N_5998,N_5902,N_5899);
xnor U5999 (N_5999,N_5784,N_5810);
nor U6000 (N_6000,N_5804,N_5816);
nor U6001 (N_6001,N_5768,N_5825);
or U6002 (N_6002,N_5812,N_5854);
nand U6003 (N_6003,N_5891,N_5842);
or U6004 (N_6004,N_5851,N_5850);
nand U6005 (N_6005,N_5894,N_5879);
nand U6006 (N_6006,N_5908,N_5782);
or U6007 (N_6007,N_5876,N_5808);
or U6008 (N_6008,N_5840,N_5802);
nand U6009 (N_6009,N_5843,N_5817);
xnor U6010 (N_6010,N_5881,N_5877);
nand U6011 (N_6011,N_5808,N_5859);
or U6012 (N_6012,N_5774,N_5764);
xor U6013 (N_6013,N_5783,N_5889);
nand U6014 (N_6014,N_5897,N_5783);
nand U6015 (N_6015,N_5890,N_5909);
xnor U6016 (N_6016,N_5846,N_5824);
nand U6017 (N_6017,N_5765,N_5818);
and U6018 (N_6018,N_5851,N_5849);
or U6019 (N_6019,N_5773,N_5851);
nor U6020 (N_6020,N_5876,N_5911);
nand U6021 (N_6021,N_5821,N_5855);
or U6022 (N_6022,N_5839,N_5838);
nand U6023 (N_6023,N_5870,N_5832);
xnor U6024 (N_6024,N_5889,N_5779);
xor U6025 (N_6025,N_5904,N_5891);
nand U6026 (N_6026,N_5775,N_5861);
or U6027 (N_6027,N_5913,N_5908);
and U6028 (N_6028,N_5914,N_5827);
and U6029 (N_6029,N_5868,N_5814);
nor U6030 (N_6030,N_5785,N_5875);
and U6031 (N_6031,N_5773,N_5848);
xnor U6032 (N_6032,N_5761,N_5882);
nor U6033 (N_6033,N_5778,N_5762);
and U6034 (N_6034,N_5835,N_5865);
xor U6035 (N_6035,N_5855,N_5858);
and U6036 (N_6036,N_5808,N_5866);
and U6037 (N_6037,N_5860,N_5801);
nand U6038 (N_6038,N_5892,N_5906);
nor U6039 (N_6039,N_5860,N_5841);
nand U6040 (N_6040,N_5813,N_5806);
nor U6041 (N_6041,N_5820,N_5864);
nand U6042 (N_6042,N_5897,N_5909);
nand U6043 (N_6043,N_5885,N_5893);
nor U6044 (N_6044,N_5799,N_5771);
and U6045 (N_6045,N_5860,N_5868);
or U6046 (N_6046,N_5911,N_5850);
and U6047 (N_6047,N_5888,N_5785);
nand U6048 (N_6048,N_5903,N_5832);
or U6049 (N_6049,N_5823,N_5843);
and U6050 (N_6050,N_5918,N_5810);
nor U6051 (N_6051,N_5861,N_5812);
nand U6052 (N_6052,N_5823,N_5850);
xnor U6053 (N_6053,N_5811,N_5864);
and U6054 (N_6054,N_5913,N_5886);
nand U6055 (N_6055,N_5917,N_5894);
and U6056 (N_6056,N_5914,N_5765);
or U6057 (N_6057,N_5763,N_5904);
nor U6058 (N_6058,N_5893,N_5896);
or U6059 (N_6059,N_5844,N_5794);
nand U6060 (N_6060,N_5789,N_5893);
and U6061 (N_6061,N_5907,N_5827);
nor U6062 (N_6062,N_5867,N_5874);
nor U6063 (N_6063,N_5882,N_5916);
nand U6064 (N_6064,N_5913,N_5797);
or U6065 (N_6065,N_5885,N_5781);
or U6066 (N_6066,N_5867,N_5792);
nand U6067 (N_6067,N_5886,N_5836);
xor U6068 (N_6068,N_5804,N_5760);
and U6069 (N_6069,N_5847,N_5870);
nor U6070 (N_6070,N_5787,N_5919);
xor U6071 (N_6071,N_5896,N_5910);
and U6072 (N_6072,N_5887,N_5769);
nor U6073 (N_6073,N_5832,N_5797);
nor U6074 (N_6074,N_5770,N_5811);
xor U6075 (N_6075,N_5918,N_5876);
or U6076 (N_6076,N_5829,N_5761);
or U6077 (N_6077,N_5772,N_5792);
nand U6078 (N_6078,N_5882,N_5803);
and U6079 (N_6079,N_5884,N_5800);
xor U6080 (N_6080,N_5958,N_5988);
nand U6081 (N_6081,N_5996,N_5936);
or U6082 (N_6082,N_6068,N_5948);
or U6083 (N_6083,N_5921,N_5923);
and U6084 (N_6084,N_6012,N_6051);
and U6085 (N_6085,N_6044,N_6047);
nor U6086 (N_6086,N_6000,N_5946);
nand U6087 (N_6087,N_5990,N_6073);
nor U6088 (N_6088,N_5922,N_6027);
nor U6089 (N_6089,N_5931,N_5972);
xor U6090 (N_6090,N_5989,N_5928);
nand U6091 (N_6091,N_5926,N_5984);
nor U6092 (N_6092,N_5940,N_5967);
nand U6093 (N_6093,N_5992,N_6011);
or U6094 (N_6094,N_6014,N_5935);
or U6095 (N_6095,N_5941,N_6053);
xnor U6096 (N_6096,N_6003,N_5987);
or U6097 (N_6097,N_6021,N_5999);
or U6098 (N_6098,N_6071,N_6060);
or U6099 (N_6099,N_5975,N_6077);
and U6100 (N_6100,N_5979,N_6006);
or U6101 (N_6101,N_6025,N_5964);
xnor U6102 (N_6102,N_6074,N_5938);
nand U6103 (N_6103,N_6046,N_5924);
xor U6104 (N_6104,N_6009,N_5963);
and U6105 (N_6105,N_6033,N_6045);
nand U6106 (N_6106,N_5944,N_6066);
or U6107 (N_6107,N_6023,N_6076);
and U6108 (N_6108,N_5920,N_6052);
xnor U6109 (N_6109,N_6048,N_6043);
nor U6110 (N_6110,N_6001,N_5991);
nand U6111 (N_6111,N_5970,N_6067);
xor U6112 (N_6112,N_6017,N_5985);
nor U6113 (N_6113,N_5949,N_6007);
nand U6114 (N_6114,N_5995,N_5962);
nand U6115 (N_6115,N_5952,N_6049);
xor U6116 (N_6116,N_6034,N_5956);
and U6117 (N_6117,N_5942,N_6072);
xor U6118 (N_6118,N_6026,N_5953);
xnor U6119 (N_6119,N_5934,N_5937);
and U6120 (N_6120,N_5957,N_5939);
nand U6121 (N_6121,N_6036,N_6016);
nand U6122 (N_6122,N_5966,N_5930);
and U6123 (N_6123,N_5961,N_6022);
nand U6124 (N_6124,N_6057,N_5959);
or U6125 (N_6125,N_6031,N_5965);
and U6126 (N_6126,N_5977,N_5976);
or U6127 (N_6127,N_6029,N_5960);
or U6128 (N_6128,N_5933,N_6038);
xnor U6129 (N_6129,N_5925,N_5983);
nand U6130 (N_6130,N_6075,N_5978);
and U6131 (N_6131,N_6063,N_6002);
and U6132 (N_6132,N_5981,N_6041);
xor U6133 (N_6133,N_5947,N_5993);
or U6134 (N_6134,N_6024,N_6079);
xor U6135 (N_6135,N_6028,N_6056);
or U6136 (N_6136,N_5955,N_5982);
nand U6137 (N_6137,N_5973,N_5927);
xor U6138 (N_6138,N_6032,N_6061);
nor U6139 (N_6139,N_6040,N_5951);
xor U6140 (N_6140,N_5971,N_6018);
xor U6141 (N_6141,N_5974,N_6050);
nand U6142 (N_6142,N_6019,N_6058);
or U6143 (N_6143,N_6069,N_6008);
or U6144 (N_6144,N_6042,N_6064);
and U6145 (N_6145,N_6078,N_5969);
nor U6146 (N_6146,N_6055,N_6010);
or U6147 (N_6147,N_5986,N_5968);
nor U6148 (N_6148,N_5929,N_5980);
nor U6149 (N_6149,N_5998,N_6062);
nand U6150 (N_6150,N_6013,N_5932);
nor U6151 (N_6151,N_6065,N_6004);
nor U6152 (N_6152,N_5945,N_6037);
and U6153 (N_6153,N_6070,N_5943);
and U6154 (N_6154,N_6054,N_6030);
xnor U6155 (N_6155,N_6005,N_6015);
xor U6156 (N_6156,N_6039,N_6059);
nor U6157 (N_6157,N_5950,N_5997);
nor U6158 (N_6158,N_6020,N_6035);
or U6159 (N_6159,N_5994,N_5954);
nand U6160 (N_6160,N_5954,N_5975);
nor U6161 (N_6161,N_6074,N_5964);
or U6162 (N_6162,N_5955,N_6033);
xnor U6163 (N_6163,N_6055,N_5971);
or U6164 (N_6164,N_5924,N_5962);
nand U6165 (N_6165,N_5956,N_6041);
nand U6166 (N_6166,N_6013,N_5954);
nor U6167 (N_6167,N_6002,N_6019);
and U6168 (N_6168,N_6019,N_6044);
nand U6169 (N_6169,N_5936,N_6002);
nand U6170 (N_6170,N_6012,N_5957);
and U6171 (N_6171,N_5925,N_6023);
xor U6172 (N_6172,N_6009,N_5958);
nand U6173 (N_6173,N_6035,N_5997);
nand U6174 (N_6174,N_5940,N_6060);
nor U6175 (N_6175,N_5923,N_6030);
and U6176 (N_6176,N_5972,N_5981);
nor U6177 (N_6177,N_5999,N_6031);
nand U6178 (N_6178,N_5946,N_5970);
nand U6179 (N_6179,N_5923,N_5959);
nor U6180 (N_6180,N_5950,N_5934);
xor U6181 (N_6181,N_6044,N_6067);
or U6182 (N_6182,N_5969,N_6057);
or U6183 (N_6183,N_5920,N_5966);
xnor U6184 (N_6184,N_5935,N_5967);
or U6185 (N_6185,N_5959,N_6047);
nand U6186 (N_6186,N_6015,N_6068);
nor U6187 (N_6187,N_5943,N_6038);
nor U6188 (N_6188,N_6044,N_5943);
nor U6189 (N_6189,N_6039,N_5970);
and U6190 (N_6190,N_5938,N_5946);
nor U6191 (N_6191,N_5988,N_5921);
nand U6192 (N_6192,N_5955,N_6014);
xnor U6193 (N_6193,N_5984,N_6041);
xor U6194 (N_6194,N_6031,N_5978);
nand U6195 (N_6195,N_5925,N_5985);
xor U6196 (N_6196,N_6049,N_6077);
xnor U6197 (N_6197,N_5992,N_5975);
xnor U6198 (N_6198,N_6066,N_6067);
and U6199 (N_6199,N_5925,N_5951);
or U6200 (N_6200,N_6035,N_6010);
nor U6201 (N_6201,N_6067,N_6064);
and U6202 (N_6202,N_6056,N_6026);
nor U6203 (N_6203,N_5964,N_6055);
or U6204 (N_6204,N_5973,N_6007);
or U6205 (N_6205,N_5958,N_6063);
or U6206 (N_6206,N_6050,N_5950);
and U6207 (N_6207,N_6001,N_5924);
nand U6208 (N_6208,N_5998,N_6053);
nor U6209 (N_6209,N_6007,N_6006);
nand U6210 (N_6210,N_6002,N_5923);
nand U6211 (N_6211,N_6070,N_5990);
nand U6212 (N_6212,N_5997,N_6032);
and U6213 (N_6213,N_5940,N_6053);
nand U6214 (N_6214,N_5978,N_5963);
xor U6215 (N_6215,N_5993,N_5974);
nor U6216 (N_6216,N_5963,N_6068);
nor U6217 (N_6217,N_5930,N_5933);
nor U6218 (N_6218,N_5954,N_6044);
or U6219 (N_6219,N_6058,N_6024);
nand U6220 (N_6220,N_5925,N_5929);
nand U6221 (N_6221,N_6040,N_5994);
and U6222 (N_6222,N_6012,N_6076);
nand U6223 (N_6223,N_6003,N_5926);
xnor U6224 (N_6224,N_6047,N_5996);
or U6225 (N_6225,N_5969,N_5958);
xor U6226 (N_6226,N_6040,N_6058);
nand U6227 (N_6227,N_6045,N_5938);
nand U6228 (N_6228,N_6065,N_5945);
or U6229 (N_6229,N_5929,N_5989);
nand U6230 (N_6230,N_6008,N_5995);
and U6231 (N_6231,N_5988,N_5920);
or U6232 (N_6232,N_5984,N_6078);
nand U6233 (N_6233,N_5953,N_5924);
nor U6234 (N_6234,N_5924,N_5947);
xor U6235 (N_6235,N_6054,N_6016);
or U6236 (N_6236,N_5975,N_6063);
or U6237 (N_6237,N_5999,N_6033);
nor U6238 (N_6238,N_6011,N_5941);
xnor U6239 (N_6239,N_6007,N_6050);
nor U6240 (N_6240,N_6228,N_6167);
nor U6241 (N_6241,N_6202,N_6207);
xnor U6242 (N_6242,N_6210,N_6162);
nor U6243 (N_6243,N_6187,N_6197);
and U6244 (N_6244,N_6203,N_6127);
or U6245 (N_6245,N_6174,N_6159);
or U6246 (N_6246,N_6110,N_6141);
or U6247 (N_6247,N_6222,N_6223);
or U6248 (N_6248,N_6115,N_6082);
xnor U6249 (N_6249,N_6112,N_6221);
nand U6250 (N_6250,N_6089,N_6151);
nand U6251 (N_6251,N_6209,N_6092);
xor U6252 (N_6252,N_6144,N_6198);
nand U6253 (N_6253,N_6143,N_6194);
nor U6254 (N_6254,N_6133,N_6208);
nor U6255 (N_6255,N_6091,N_6216);
nor U6256 (N_6256,N_6200,N_6190);
or U6257 (N_6257,N_6128,N_6196);
nand U6258 (N_6258,N_6142,N_6171);
or U6259 (N_6259,N_6175,N_6085);
nor U6260 (N_6260,N_6093,N_6149);
nand U6261 (N_6261,N_6163,N_6173);
and U6262 (N_6262,N_6113,N_6157);
nand U6263 (N_6263,N_6235,N_6121);
or U6264 (N_6264,N_6230,N_6238);
nor U6265 (N_6265,N_6080,N_6122);
xor U6266 (N_6266,N_6229,N_6137);
xnor U6267 (N_6267,N_6232,N_6226);
and U6268 (N_6268,N_6096,N_6183);
nor U6269 (N_6269,N_6125,N_6118);
xor U6270 (N_6270,N_6098,N_6087);
or U6271 (N_6271,N_6179,N_6180);
nand U6272 (N_6272,N_6129,N_6192);
xnor U6273 (N_6273,N_6131,N_6188);
nor U6274 (N_6274,N_6166,N_6145);
nor U6275 (N_6275,N_6099,N_6109);
nand U6276 (N_6276,N_6186,N_6160);
nor U6277 (N_6277,N_6195,N_6178);
or U6278 (N_6278,N_6153,N_6106);
nor U6279 (N_6279,N_6083,N_6204);
xnor U6280 (N_6280,N_6132,N_6193);
nand U6281 (N_6281,N_6100,N_6084);
xor U6282 (N_6282,N_6214,N_6182);
nand U6283 (N_6283,N_6172,N_6199);
and U6284 (N_6284,N_6205,N_6220);
xnor U6285 (N_6285,N_6212,N_6231);
or U6286 (N_6286,N_6102,N_6170);
xor U6287 (N_6287,N_6234,N_6225);
nor U6288 (N_6288,N_6123,N_6140);
or U6289 (N_6289,N_6134,N_6097);
nand U6290 (N_6290,N_6176,N_6177);
nand U6291 (N_6291,N_6138,N_6111);
and U6292 (N_6292,N_6114,N_6107);
nor U6293 (N_6293,N_6218,N_6239);
nand U6294 (N_6294,N_6136,N_6126);
nand U6295 (N_6295,N_6094,N_6227);
and U6296 (N_6296,N_6213,N_6103);
and U6297 (N_6297,N_6155,N_6189);
and U6298 (N_6298,N_6201,N_6211);
xor U6299 (N_6299,N_6165,N_6161);
nor U6300 (N_6300,N_6215,N_6148);
and U6301 (N_6301,N_6124,N_6147);
nand U6302 (N_6302,N_6168,N_6119);
xor U6303 (N_6303,N_6116,N_6081);
or U6304 (N_6304,N_6224,N_6206);
and U6305 (N_6305,N_6130,N_6169);
and U6306 (N_6306,N_6090,N_6135);
and U6307 (N_6307,N_6095,N_6154);
and U6308 (N_6308,N_6191,N_6181);
or U6309 (N_6309,N_6217,N_6120);
nor U6310 (N_6310,N_6185,N_6139);
xor U6311 (N_6311,N_6184,N_6236);
and U6312 (N_6312,N_6104,N_6088);
nor U6313 (N_6313,N_6150,N_6237);
or U6314 (N_6314,N_6117,N_6086);
and U6315 (N_6315,N_6105,N_6146);
xnor U6316 (N_6316,N_6164,N_6233);
nand U6317 (N_6317,N_6158,N_6219);
nand U6318 (N_6318,N_6108,N_6156);
or U6319 (N_6319,N_6101,N_6152);
xnor U6320 (N_6320,N_6181,N_6213);
or U6321 (N_6321,N_6155,N_6098);
nand U6322 (N_6322,N_6234,N_6082);
nand U6323 (N_6323,N_6157,N_6129);
and U6324 (N_6324,N_6084,N_6183);
nand U6325 (N_6325,N_6123,N_6109);
nand U6326 (N_6326,N_6189,N_6177);
or U6327 (N_6327,N_6154,N_6152);
or U6328 (N_6328,N_6161,N_6097);
nand U6329 (N_6329,N_6219,N_6152);
and U6330 (N_6330,N_6086,N_6150);
nand U6331 (N_6331,N_6136,N_6152);
xnor U6332 (N_6332,N_6106,N_6163);
xnor U6333 (N_6333,N_6086,N_6098);
xor U6334 (N_6334,N_6209,N_6150);
nor U6335 (N_6335,N_6192,N_6171);
nor U6336 (N_6336,N_6233,N_6223);
nor U6337 (N_6337,N_6148,N_6173);
and U6338 (N_6338,N_6102,N_6186);
or U6339 (N_6339,N_6120,N_6116);
nand U6340 (N_6340,N_6100,N_6229);
xor U6341 (N_6341,N_6086,N_6160);
nand U6342 (N_6342,N_6178,N_6136);
and U6343 (N_6343,N_6095,N_6177);
or U6344 (N_6344,N_6229,N_6192);
nand U6345 (N_6345,N_6217,N_6115);
or U6346 (N_6346,N_6082,N_6163);
and U6347 (N_6347,N_6101,N_6218);
nand U6348 (N_6348,N_6089,N_6201);
xnor U6349 (N_6349,N_6103,N_6126);
nand U6350 (N_6350,N_6106,N_6117);
or U6351 (N_6351,N_6151,N_6233);
or U6352 (N_6352,N_6196,N_6175);
nor U6353 (N_6353,N_6133,N_6095);
xor U6354 (N_6354,N_6153,N_6203);
nor U6355 (N_6355,N_6081,N_6083);
or U6356 (N_6356,N_6125,N_6237);
nor U6357 (N_6357,N_6192,N_6177);
or U6358 (N_6358,N_6140,N_6086);
or U6359 (N_6359,N_6199,N_6090);
nand U6360 (N_6360,N_6152,N_6127);
and U6361 (N_6361,N_6217,N_6091);
nor U6362 (N_6362,N_6099,N_6202);
nand U6363 (N_6363,N_6133,N_6179);
or U6364 (N_6364,N_6238,N_6128);
nand U6365 (N_6365,N_6105,N_6213);
xor U6366 (N_6366,N_6222,N_6211);
or U6367 (N_6367,N_6097,N_6137);
xnor U6368 (N_6368,N_6184,N_6207);
or U6369 (N_6369,N_6152,N_6099);
or U6370 (N_6370,N_6193,N_6155);
nor U6371 (N_6371,N_6164,N_6190);
and U6372 (N_6372,N_6082,N_6131);
xor U6373 (N_6373,N_6173,N_6159);
nand U6374 (N_6374,N_6157,N_6132);
nor U6375 (N_6375,N_6095,N_6138);
nand U6376 (N_6376,N_6187,N_6086);
and U6377 (N_6377,N_6108,N_6176);
xor U6378 (N_6378,N_6144,N_6211);
nor U6379 (N_6379,N_6096,N_6147);
or U6380 (N_6380,N_6182,N_6198);
nor U6381 (N_6381,N_6135,N_6137);
nand U6382 (N_6382,N_6158,N_6194);
nor U6383 (N_6383,N_6172,N_6145);
nor U6384 (N_6384,N_6181,N_6203);
or U6385 (N_6385,N_6118,N_6179);
xor U6386 (N_6386,N_6206,N_6232);
nor U6387 (N_6387,N_6218,N_6103);
nand U6388 (N_6388,N_6197,N_6168);
nor U6389 (N_6389,N_6119,N_6223);
xor U6390 (N_6390,N_6157,N_6164);
or U6391 (N_6391,N_6080,N_6196);
and U6392 (N_6392,N_6219,N_6237);
and U6393 (N_6393,N_6113,N_6170);
or U6394 (N_6394,N_6133,N_6224);
nand U6395 (N_6395,N_6228,N_6179);
nand U6396 (N_6396,N_6175,N_6169);
nand U6397 (N_6397,N_6224,N_6161);
or U6398 (N_6398,N_6218,N_6122);
nor U6399 (N_6399,N_6131,N_6102);
and U6400 (N_6400,N_6298,N_6357);
xnor U6401 (N_6401,N_6253,N_6274);
nor U6402 (N_6402,N_6359,N_6266);
or U6403 (N_6403,N_6251,N_6352);
nor U6404 (N_6404,N_6288,N_6310);
nor U6405 (N_6405,N_6291,N_6303);
and U6406 (N_6406,N_6327,N_6374);
and U6407 (N_6407,N_6351,N_6286);
nor U6408 (N_6408,N_6263,N_6382);
and U6409 (N_6409,N_6312,N_6325);
and U6410 (N_6410,N_6315,N_6330);
or U6411 (N_6411,N_6241,N_6247);
nor U6412 (N_6412,N_6262,N_6304);
nor U6413 (N_6413,N_6393,N_6248);
and U6414 (N_6414,N_6340,N_6392);
and U6415 (N_6415,N_6240,N_6378);
xnor U6416 (N_6416,N_6313,N_6388);
nor U6417 (N_6417,N_6326,N_6269);
nor U6418 (N_6418,N_6255,N_6394);
nor U6419 (N_6419,N_6387,N_6376);
nor U6420 (N_6420,N_6271,N_6391);
and U6421 (N_6421,N_6366,N_6329);
and U6422 (N_6422,N_6318,N_6301);
nand U6423 (N_6423,N_6333,N_6360);
nand U6424 (N_6424,N_6350,N_6314);
nor U6425 (N_6425,N_6324,N_6280);
xnor U6426 (N_6426,N_6368,N_6297);
nor U6427 (N_6427,N_6386,N_6305);
and U6428 (N_6428,N_6335,N_6367);
or U6429 (N_6429,N_6299,N_6284);
nor U6430 (N_6430,N_6295,N_6249);
nand U6431 (N_6431,N_6371,N_6296);
xnor U6432 (N_6432,N_6245,N_6328);
and U6433 (N_6433,N_6331,N_6375);
xor U6434 (N_6434,N_6283,N_6389);
or U6435 (N_6435,N_6373,N_6281);
or U6436 (N_6436,N_6289,N_6293);
nand U6437 (N_6437,N_6364,N_6347);
nor U6438 (N_6438,N_6307,N_6370);
and U6439 (N_6439,N_6267,N_6399);
or U6440 (N_6440,N_6337,N_6300);
nor U6441 (N_6441,N_6294,N_6259);
nand U6442 (N_6442,N_6287,N_6322);
nand U6443 (N_6443,N_6383,N_6302);
xor U6444 (N_6444,N_6344,N_6273);
nor U6445 (N_6445,N_6385,N_6356);
and U6446 (N_6446,N_6282,N_6365);
and U6447 (N_6447,N_6341,N_6290);
xor U6448 (N_6448,N_6363,N_6285);
and U6449 (N_6449,N_6342,N_6306);
and U6450 (N_6450,N_6264,N_6265);
xnor U6451 (N_6451,N_6254,N_6270);
and U6452 (N_6452,N_6321,N_6358);
nor U6453 (N_6453,N_6398,N_6292);
and U6454 (N_6454,N_6257,N_6345);
nor U6455 (N_6455,N_6354,N_6362);
nor U6456 (N_6456,N_6384,N_6319);
xnor U6457 (N_6457,N_6390,N_6381);
and U6458 (N_6458,N_6272,N_6380);
nand U6459 (N_6459,N_6334,N_6346);
and U6460 (N_6460,N_6343,N_6275);
nor U6461 (N_6461,N_6279,N_6317);
nor U6462 (N_6462,N_6396,N_6369);
xor U6463 (N_6463,N_6320,N_6377);
and U6464 (N_6464,N_6395,N_6277);
and U6465 (N_6465,N_6311,N_6268);
or U6466 (N_6466,N_6332,N_6397);
nand U6467 (N_6467,N_6349,N_6250);
and U6468 (N_6468,N_6379,N_6256);
nand U6469 (N_6469,N_6361,N_6242);
nand U6470 (N_6470,N_6353,N_6348);
nor U6471 (N_6471,N_6260,N_6278);
nor U6472 (N_6472,N_6246,N_6316);
nor U6473 (N_6473,N_6252,N_6339);
or U6474 (N_6474,N_6355,N_6309);
xnor U6475 (N_6475,N_6308,N_6338);
nand U6476 (N_6476,N_6258,N_6336);
nor U6477 (N_6477,N_6261,N_6372);
and U6478 (N_6478,N_6276,N_6323);
nand U6479 (N_6479,N_6243,N_6244);
or U6480 (N_6480,N_6310,N_6258);
nand U6481 (N_6481,N_6372,N_6259);
nor U6482 (N_6482,N_6386,N_6373);
nand U6483 (N_6483,N_6364,N_6323);
nor U6484 (N_6484,N_6268,N_6295);
xnor U6485 (N_6485,N_6246,N_6270);
nand U6486 (N_6486,N_6346,N_6356);
and U6487 (N_6487,N_6245,N_6351);
or U6488 (N_6488,N_6380,N_6355);
nand U6489 (N_6489,N_6329,N_6315);
nor U6490 (N_6490,N_6361,N_6257);
xnor U6491 (N_6491,N_6266,N_6369);
and U6492 (N_6492,N_6379,N_6392);
nor U6493 (N_6493,N_6385,N_6362);
xor U6494 (N_6494,N_6250,N_6309);
nand U6495 (N_6495,N_6311,N_6334);
xnor U6496 (N_6496,N_6325,N_6349);
and U6497 (N_6497,N_6285,N_6395);
or U6498 (N_6498,N_6254,N_6392);
or U6499 (N_6499,N_6287,N_6332);
nand U6500 (N_6500,N_6246,N_6273);
nor U6501 (N_6501,N_6367,N_6374);
xnor U6502 (N_6502,N_6297,N_6315);
nor U6503 (N_6503,N_6304,N_6339);
nor U6504 (N_6504,N_6353,N_6266);
nor U6505 (N_6505,N_6258,N_6303);
and U6506 (N_6506,N_6351,N_6319);
xnor U6507 (N_6507,N_6395,N_6300);
and U6508 (N_6508,N_6298,N_6346);
nor U6509 (N_6509,N_6299,N_6349);
and U6510 (N_6510,N_6277,N_6308);
xor U6511 (N_6511,N_6341,N_6244);
nor U6512 (N_6512,N_6282,N_6307);
nand U6513 (N_6513,N_6287,N_6260);
xnor U6514 (N_6514,N_6258,N_6362);
xnor U6515 (N_6515,N_6253,N_6301);
nor U6516 (N_6516,N_6301,N_6369);
nand U6517 (N_6517,N_6380,N_6266);
xnor U6518 (N_6518,N_6327,N_6395);
nand U6519 (N_6519,N_6270,N_6348);
nand U6520 (N_6520,N_6312,N_6324);
or U6521 (N_6521,N_6335,N_6393);
nor U6522 (N_6522,N_6299,N_6274);
and U6523 (N_6523,N_6269,N_6337);
nand U6524 (N_6524,N_6240,N_6314);
nor U6525 (N_6525,N_6261,N_6282);
xnor U6526 (N_6526,N_6261,N_6290);
and U6527 (N_6527,N_6350,N_6395);
xnor U6528 (N_6528,N_6360,N_6367);
and U6529 (N_6529,N_6330,N_6256);
xnor U6530 (N_6530,N_6310,N_6342);
and U6531 (N_6531,N_6292,N_6301);
or U6532 (N_6532,N_6282,N_6384);
xnor U6533 (N_6533,N_6260,N_6366);
or U6534 (N_6534,N_6396,N_6242);
xor U6535 (N_6535,N_6277,N_6300);
xnor U6536 (N_6536,N_6318,N_6287);
or U6537 (N_6537,N_6273,N_6274);
nor U6538 (N_6538,N_6397,N_6337);
nor U6539 (N_6539,N_6285,N_6259);
nor U6540 (N_6540,N_6363,N_6384);
and U6541 (N_6541,N_6348,N_6298);
or U6542 (N_6542,N_6257,N_6254);
or U6543 (N_6543,N_6300,N_6264);
nor U6544 (N_6544,N_6341,N_6292);
xnor U6545 (N_6545,N_6303,N_6242);
and U6546 (N_6546,N_6329,N_6374);
xor U6547 (N_6547,N_6300,N_6379);
nor U6548 (N_6548,N_6372,N_6279);
xor U6549 (N_6549,N_6396,N_6298);
nand U6550 (N_6550,N_6340,N_6318);
and U6551 (N_6551,N_6317,N_6345);
or U6552 (N_6552,N_6364,N_6371);
and U6553 (N_6553,N_6323,N_6395);
nand U6554 (N_6554,N_6244,N_6314);
and U6555 (N_6555,N_6342,N_6346);
nand U6556 (N_6556,N_6389,N_6286);
nand U6557 (N_6557,N_6245,N_6370);
or U6558 (N_6558,N_6350,N_6321);
nand U6559 (N_6559,N_6263,N_6357);
xnor U6560 (N_6560,N_6522,N_6557);
nor U6561 (N_6561,N_6466,N_6472);
nand U6562 (N_6562,N_6482,N_6511);
or U6563 (N_6563,N_6480,N_6493);
xor U6564 (N_6564,N_6449,N_6497);
and U6565 (N_6565,N_6525,N_6537);
xor U6566 (N_6566,N_6413,N_6555);
nand U6567 (N_6567,N_6477,N_6468);
nor U6568 (N_6568,N_6403,N_6441);
xnor U6569 (N_6569,N_6431,N_6454);
xor U6570 (N_6570,N_6505,N_6438);
xor U6571 (N_6571,N_6410,N_6479);
nor U6572 (N_6572,N_6459,N_6427);
or U6573 (N_6573,N_6415,N_6519);
nand U6574 (N_6574,N_6420,N_6538);
nand U6575 (N_6575,N_6458,N_6423);
nand U6576 (N_6576,N_6416,N_6409);
nor U6577 (N_6577,N_6526,N_6447);
or U6578 (N_6578,N_6434,N_6451);
and U6579 (N_6579,N_6556,N_6474);
xor U6580 (N_6580,N_6510,N_6456);
nor U6581 (N_6581,N_6504,N_6455);
nand U6582 (N_6582,N_6498,N_6514);
xnor U6583 (N_6583,N_6520,N_6412);
nand U6584 (N_6584,N_6443,N_6503);
xnor U6585 (N_6585,N_6542,N_6533);
nand U6586 (N_6586,N_6461,N_6559);
or U6587 (N_6587,N_6436,N_6445);
or U6588 (N_6588,N_6418,N_6453);
nand U6589 (N_6589,N_6545,N_6463);
nor U6590 (N_6590,N_6536,N_6489);
xor U6591 (N_6591,N_6554,N_6541);
or U6592 (N_6592,N_6491,N_6444);
and U6593 (N_6593,N_6457,N_6547);
nand U6594 (N_6594,N_6496,N_6475);
xor U6595 (N_6595,N_6551,N_6476);
and U6596 (N_6596,N_6524,N_6539);
nor U6597 (N_6597,N_6512,N_6473);
xor U6598 (N_6598,N_6478,N_6535);
and U6599 (N_6599,N_6486,N_6552);
or U6600 (N_6600,N_6408,N_6513);
or U6601 (N_6601,N_6499,N_6470);
and U6602 (N_6602,N_6528,N_6465);
or U6603 (N_6603,N_6417,N_6501);
nor U6604 (N_6604,N_6448,N_6532);
nor U6605 (N_6605,N_6471,N_6419);
and U6606 (N_6606,N_6428,N_6500);
or U6607 (N_6607,N_6549,N_6421);
nand U6608 (N_6608,N_6523,N_6432);
and U6609 (N_6609,N_6492,N_6546);
nor U6610 (N_6610,N_6517,N_6508);
nor U6611 (N_6611,N_6540,N_6507);
nand U6612 (N_6612,N_6485,N_6506);
or U6613 (N_6613,N_6548,N_6429);
nand U6614 (N_6614,N_6442,N_6467);
and U6615 (N_6615,N_6516,N_6422);
nor U6616 (N_6616,N_6515,N_6462);
nor U6617 (N_6617,N_6404,N_6435);
or U6618 (N_6618,N_6464,N_6484);
and U6619 (N_6619,N_6450,N_6490);
nand U6620 (N_6620,N_6406,N_6527);
nor U6621 (N_6621,N_6530,N_6469);
nand U6622 (N_6622,N_6487,N_6534);
and U6623 (N_6623,N_6544,N_6531);
and U6624 (N_6624,N_6405,N_6502);
nand U6625 (N_6625,N_6402,N_6411);
or U6626 (N_6626,N_6529,N_6452);
or U6627 (N_6627,N_6481,N_6424);
nor U6628 (N_6628,N_6446,N_6400);
nor U6629 (N_6629,N_6437,N_6553);
xnor U6630 (N_6630,N_6426,N_6401);
and U6631 (N_6631,N_6494,N_6509);
xor U6632 (N_6632,N_6460,N_6495);
and U6633 (N_6633,N_6518,N_6440);
nand U6634 (N_6634,N_6543,N_6488);
or U6635 (N_6635,N_6433,N_6558);
nor U6636 (N_6636,N_6483,N_6425);
nor U6637 (N_6637,N_6414,N_6430);
nand U6638 (N_6638,N_6439,N_6521);
nand U6639 (N_6639,N_6407,N_6550);
nor U6640 (N_6640,N_6463,N_6551);
nand U6641 (N_6641,N_6558,N_6531);
and U6642 (N_6642,N_6493,N_6450);
xnor U6643 (N_6643,N_6487,N_6462);
nor U6644 (N_6644,N_6403,N_6452);
xnor U6645 (N_6645,N_6497,N_6434);
nand U6646 (N_6646,N_6518,N_6411);
nor U6647 (N_6647,N_6482,N_6522);
nand U6648 (N_6648,N_6513,N_6425);
and U6649 (N_6649,N_6453,N_6450);
or U6650 (N_6650,N_6522,N_6502);
and U6651 (N_6651,N_6404,N_6432);
xor U6652 (N_6652,N_6466,N_6477);
nor U6653 (N_6653,N_6550,N_6465);
nor U6654 (N_6654,N_6530,N_6527);
or U6655 (N_6655,N_6537,N_6408);
and U6656 (N_6656,N_6444,N_6552);
nand U6657 (N_6657,N_6479,N_6552);
nor U6658 (N_6658,N_6408,N_6533);
nor U6659 (N_6659,N_6499,N_6424);
nand U6660 (N_6660,N_6462,N_6416);
xor U6661 (N_6661,N_6465,N_6437);
nor U6662 (N_6662,N_6523,N_6494);
nand U6663 (N_6663,N_6412,N_6516);
or U6664 (N_6664,N_6503,N_6454);
or U6665 (N_6665,N_6439,N_6468);
xnor U6666 (N_6666,N_6534,N_6441);
xnor U6667 (N_6667,N_6405,N_6538);
and U6668 (N_6668,N_6542,N_6448);
nor U6669 (N_6669,N_6411,N_6432);
xor U6670 (N_6670,N_6477,N_6441);
xor U6671 (N_6671,N_6534,N_6440);
nor U6672 (N_6672,N_6537,N_6495);
nand U6673 (N_6673,N_6510,N_6532);
xnor U6674 (N_6674,N_6431,N_6524);
xnor U6675 (N_6675,N_6462,N_6465);
xnor U6676 (N_6676,N_6505,N_6418);
xor U6677 (N_6677,N_6504,N_6409);
nor U6678 (N_6678,N_6425,N_6447);
and U6679 (N_6679,N_6458,N_6438);
xor U6680 (N_6680,N_6471,N_6477);
or U6681 (N_6681,N_6491,N_6484);
and U6682 (N_6682,N_6444,N_6529);
nand U6683 (N_6683,N_6535,N_6485);
or U6684 (N_6684,N_6401,N_6520);
or U6685 (N_6685,N_6524,N_6409);
nand U6686 (N_6686,N_6411,N_6410);
nand U6687 (N_6687,N_6450,N_6521);
xor U6688 (N_6688,N_6458,N_6462);
nor U6689 (N_6689,N_6457,N_6473);
nor U6690 (N_6690,N_6456,N_6501);
nor U6691 (N_6691,N_6400,N_6466);
nand U6692 (N_6692,N_6408,N_6479);
or U6693 (N_6693,N_6413,N_6424);
or U6694 (N_6694,N_6404,N_6506);
and U6695 (N_6695,N_6444,N_6520);
or U6696 (N_6696,N_6507,N_6470);
nor U6697 (N_6697,N_6538,N_6485);
and U6698 (N_6698,N_6543,N_6409);
nor U6699 (N_6699,N_6414,N_6506);
xnor U6700 (N_6700,N_6473,N_6462);
or U6701 (N_6701,N_6419,N_6421);
and U6702 (N_6702,N_6406,N_6547);
nand U6703 (N_6703,N_6477,N_6465);
xor U6704 (N_6704,N_6541,N_6418);
nor U6705 (N_6705,N_6546,N_6503);
and U6706 (N_6706,N_6497,N_6405);
and U6707 (N_6707,N_6425,N_6536);
nor U6708 (N_6708,N_6474,N_6510);
and U6709 (N_6709,N_6453,N_6511);
or U6710 (N_6710,N_6499,N_6437);
or U6711 (N_6711,N_6529,N_6407);
nand U6712 (N_6712,N_6485,N_6500);
nand U6713 (N_6713,N_6462,N_6559);
nand U6714 (N_6714,N_6478,N_6540);
or U6715 (N_6715,N_6420,N_6498);
nand U6716 (N_6716,N_6513,N_6459);
and U6717 (N_6717,N_6556,N_6555);
or U6718 (N_6718,N_6535,N_6415);
or U6719 (N_6719,N_6532,N_6401);
or U6720 (N_6720,N_6594,N_6701);
nand U6721 (N_6721,N_6641,N_6651);
nor U6722 (N_6722,N_6607,N_6636);
and U6723 (N_6723,N_6596,N_6566);
and U6724 (N_6724,N_6684,N_6635);
or U6725 (N_6725,N_6603,N_6655);
xor U6726 (N_6726,N_6698,N_6662);
xnor U6727 (N_6727,N_6626,N_6611);
nor U6728 (N_6728,N_6644,N_6614);
xor U6729 (N_6729,N_6714,N_6599);
and U6730 (N_6730,N_6664,N_6674);
or U6731 (N_6731,N_6693,N_6653);
nor U6732 (N_6732,N_6672,N_6629);
or U6733 (N_6733,N_6627,N_6657);
and U6734 (N_6734,N_6583,N_6719);
nand U6735 (N_6735,N_6678,N_6703);
xor U6736 (N_6736,N_6562,N_6597);
xnor U6737 (N_6737,N_6691,N_6625);
and U6738 (N_6738,N_6681,N_6579);
nand U6739 (N_6739,N_6669,N_6668);
xor U6740 (N_6740,N_6659,N_6652);
nor U6741 (N_6741,N_6648,N_6577);
nor U6742 (N_6742,N_6717,N_6595);
and U6743 (N_6743,N_6619,N_6604);
nand U6744 (N_6744,N_6598,N_6689);
and U6745 (N_6745,N_6613,N_6621);
nor U6746 (N_6746,N_6565,N_6576);
nor U6747 (N_6747,N_6661,N_6665);
nor U6748 (N_6748,N_6682,N_6571);
and U6749 (N_6749,N_6649,N_6718);
xnor U6750 (N_6750,N_6575,N_6704);
or U6751 (N_6751,N_6707,N_6697);
or U6752 (N_6752,N_6676,N_6679);
and U6753 (N_6753,N_6694,N_6609);
or U6754 (N_6754,N_6706,N_6573);
nand U6755 (N_6755,N_6570,N_6567);
xor U6756 (N_6756,N_6622,N_6645);
xor U6757 (N_6757,N_6630,N_6708);
and U6758 (N_6758,N_6580,N_6685);
or U6759 (N_6759,N_6581,N_6601);
nand U6760 (N_6760,N_6624,N_6585);
xnor U6761 (N_6761,N_6637,N_6688);
xor U6762 (N_6762,N_6673,N_6713);
nand U6763 (N_6763,N_6660,N_6591);
xor U6764 (N_6764,N_6574,N_6643);
or U6765 (N_6765,N_6561,N_6610);
and U6766 (N_6766,N_6560,N_6587);
or U6767 (N_6767,N_6666,N_6690);
or U6768 (N_6768,N_6692,N_6638);
xnor U6769 (N_6769,N_6620,N_6588);
xor U6770 (N_6770,N_6646,N_6650);
nor U6771 (N_6771,N_6564,N_6677);
nand U6772 (N_6772,N_6670,N_6584);
nor U6773 (N_6773,N_6616,N_6586);
or U6774 (N_6774,N_6634,N_6615);
and U6775 (N_6775,N_6578,N_6605);
nand U6776 (N_6776,N_6592,N_6715);
and U6777 (N_6777,N_6686,N_6608);
xor U6778 (N_6778,N_6632,N_6656);
xnor U6779 (N_6779,N_6675,N_6658);
nand U6780 (N_6780,N_6590,N_6623);
xor U6781 (N_6781,N_6618,N_6600);
and U6782 (N_6782,N_6642,N_6640);
xnor U6783 (N_6783,N_6639,N_6617);
nand U6784 (N_6784,N_6569,N_6582);
or U6785 (N_6785,N_6716,N_6711);
nor U6786 (N_6786,N_6606,N_6712);
nand U6787 (N_6787,N_6654,N_6696);
nor U6788 (N_6788,N_6702,N_6568);
xnor U6789 (N_6789,N_6647,N_6671);
nor U6790 (N_6790,N_6687,N_6563);
and U6791 (N_6791,N_6705,N_6695);
or U6792 (N_6792,N_6700,N_6709);
and U6793 (N_6793,N_6612,N_6683);
xnor U6794 (N_6794,N_6699,N_6667);
nand U6795 (N_6795,N_6710,N_6631);
and U6796 (N_6796,N_6602,N_6680);
nor U6797 (N_6797,N_6633,N_6593);
xor U6798 (N_6798,N_6663,N_6572);
and U6799 (N_6799,N_6628,N_6589);
xnor U6800 (N_6800,N_6573,N_6660);
or U6801 (N_6801,N_6579,N_6614);
and U6802 (N_6802,N_6587,N_6692);
and U6803 (N_6803,N_6640,N_6579);
and U6804 (N_6804,N_6568,N_6654);
nor U6805 (N_6805,N_6594,N_6602);
or U6806 (N_6806,N_6620,N_6678);
nor U6807 (N_6807,N_6706,N_6606);
xnor U6808 (N_6808,N_6594,N_6638);
or U6809 (N_6809,N_6709,N_6708);
xor U6810 (N_6810,N_6635,N_6592);
or U6811 (N_6811,N_6616,N_6668);
xor U6812 (N_6812,N_6639,N_6703);
xnor U6813 (N_6813,N_6573,N_6670);
nand U6814 (N_6814,N_6567,N_6599);
nand U6815 (N_6815,N_6600,N_6629);
nand U6816 (N_6816,N_6695,N_6696);
nand U6817 (N_6817,N_6685,N_6601);
nand U6818 (N_6818,N_6623,N_6576);
nand U6819 (N_6819,N_6642,N_6657);
xnor U6820 (N_6820,N_6572,N_6662);
xnor U6821 (N_6821,N_6577,N_6639);
nand U6822 (N_6822,N_6675,N_6690);
or U6823 (N_6823,N_6652,N_6580);
nand U6824 (N_6824,N_6575,N_6677);
and U6825 (N_6825,N_6694,N_6662);
or U6826 (N_6826,N_6673,N_6636);
or U6827 (N_6827,N_6692,N_6660);
xor U6828 (N_6828,N_6650,N_6591);
nor U6829 (N_6829,N_6653,N_6618);
xor U6830 (N_6830,N_6635,N_6659);
and U6831 (N_6831,N_6575,N_6641);
and U6832 (N_6832,N_6702,N_6655);
or U6833 (N_6833,N_6691,N_6699);
nor U6834 (N_6834,N_6703,N_6615);
and U6835 (N_6835,N_6632,N_6592);
nor U6836 (N_6836,N_6677,N_6708);
xnor U6837 (N_6837,N_6568,N_6622);
nand U6838 (N_6838,N_6640,N_6702);
nand U6839 (N_6839,N_6609,N_6701);
and U6840 (N_6840,N_6622,N_6705);
xnor U6841 (N_6841,N_6585,N_6680);
and U6842 (N_6842,N_6667,N_6681);
or U6843 (N_6843,N_6712,N_6590);
nor U6844 (N_6844,N_6656,N_6657);
or U6845 (N_6845,N_6572,N_6615);
nand U6846 (N_6846,N_6691,N_6636);
and U6847 (N_6847,N_6677,N_6714);
or U6848 (N_6848,N_6701,N_6703);
nand U6849 (N_6849,N_6630,N_6598);
nor U6850 (N_6850,N_6644,N_6656);
nor U6851 (N_6851,N_6674,N_6675);
nand U6852 (N_6852,N_6594,N_6687);
nand U6853 (N_6853,N_6560,N_6712);
or U6854 (N_6854,N_6677,N_6685);
or U6855 (N_6855,N_6612,N_6657);
or U6856 (N_6856,N_6628,N_6682);
or U6857 (N_6857,N_6615,N_6623);
xor U6858 (N_6858,N_6610,N_6697);
nor U6859 (N_6859,N_6671,N_6667);
nor U6860 (N_6860,N_6659,N_6571);
nand U6861 (N_6861,N_6685,N_6701);
or U6862 (N_6862,N_6617,N_6578);
nand U6863 (N_6863,N_6688,N_6591);
or U6864 (N_6864,N_6609,N_6624);
xnor U6865 (N_6865,N_6715,N_6573);
xnor U6866 (N_6866,N_6599,N_6642);
nand U6867 (N_6867,N_6567,N_6713);
nor U6868 (N_6868,N_6602,N_6585);
or U6869 (N_6869,N_6608,N_6719);
xnor U6870 (N_6870,N_6614,N_6707);
nand U6871 (N_6871,N_6698,N_6595);
nand U6872 (N_6872,N_6616,N_6697);
nand U6873 (N_6873,N_6681,N_6672);
nand U6874 (N_6874,N_6560,N_6642);
nand U6875 (N_6875,N_6632,N_6569);
or U6876 (N_6876,N_6661,N_6710);
and U6877 (N_6877,N_6584,N_6595);
xnor U6878 (N_6878,N_6584,N_6627);
nand U6879 (N_6879,N_6692,N_6693);
xor U6880 (N_6880,N_6852,N_6722);
or U6881 (N_6881,N_6875,N_6736);
nor U6882 (N_6882,N_6832,N_6851);
nor U6883 (N_6883,N_6828,N_6754);
nand U6884 (N_6884,N_6799,N_6780);
nand U6885 (N_6885,N_6784,N_6858);
nand U6886 (N_6886,N_6820,N_6819);
nand U6887 (N_6887,N_6783,N_6788);
and U6888 (N_6888,N_6815,N_6738);
xor U6889 (N_6889,N_6791,N_6794);
nand U6890 (N_6890,N_6721,N_6813);
or U6891 (N_6891,N_6795,N_6823);
nor U6892 (N_6892,N_6779,N_6760);
nor U6893 (N_6893,N_6732,N_6860);
nand U6894 (N_6894,N_6727,N_6796);
or U6895 (N_6895,N_6809,N_6731);
nand U6896 (N_6896,N_6763,N_6730);
nand U6897 (N_6897,N_6720,N_6774);
or U6898 (N_6898,N_6868,N_6803);
xnor U6899 (N_6899,N_6829,N_6733);
nand U6900 (N_6900,N_6808,N_6846);
nor U6901 (N_6901,N_6740,N_6790);
and U6902 (N_6902,N_6853,N_6729);
nand U6903 (N_6903,N_6806,N_6804);
nor U6904 (N_6904,N_6800,N_6747);
xor U6905 (N_6905,N_6855,N_6792);
nor U6906 (N_6906,N_6811,N_6807);
and U6907 (N_6907,N_6746,N_6769);
nor U6908 (N_6908,N_6762,N_6742);
xor U6909 (N_6909,N_6781,N_6728);
or U6910 (N_6910,N_6756,N_6830);
nand U6911 (N_6911,N_6825,N_6859);
xor U6912 (N_6912,N_6751,N_6785);
xnor U6913 (N_6913,N_6757,N_6782);
nand U6914 (N_6914,N_6865,N_6827);
or U6915 (N_6915,N_6798,N_6818);
and U6916 (N_6916,N_6725,N_6843);
nor U6917 (N_6917,N_6761,N_6869);
and U6918 (N_6918,N_6770,N_6759);
nor U6919 (N_6919,N_6836,N_6876);
and U6920 (N_6920,N_6743,N_6831);
or U6921 (N_6921,N_6873,N_6816);
xnor U6922 (N_6922,N_6771,N_6864);
nor U6923 (N_6923,N_6739,N_6750);
xnor U6924 (N_6924,N_6723,N_6817);
nand U6925 (N_6925,N_6870,N_6837);
nor U6926 (N_6926,N_6879,N_6741);
xnor U6927 (N_6927,N_6856,N_6764);
nand U6928 (N_6928,N_6850,N_6824);
nor U6929 (N_6929,N_6862,N_6765);
and U6930 (N_6930,N_6734,N_6812);
nor U6931 (N_6931,N_6776,N_6787);
nand U6932 (N_6932,N_6821,N_6768);
xnor U6933 (N_6933,N_6745,N_6871);
or U6934 (N_6934,N_6872,N_6801);
and U6935 (N_6935,N_6874,N_6838);
or U6936 (N_6936,N_6749,N_6878);
and U6937 (N_6937,N_6834,N_6767);
nor U6938 (N_6938,N_6744,N_6842);
nor U6939 (N_6939,N_6845,N_6752);
or U6940 (N_6940,N_6835,N_6866);
nor U6941 (N_6941,N_6863,N_6810);
and U6942 (N_6942,N_6786,N_6849);
nor U6943 (N_6943,N_6726,N_6814);
xor U6944 (N_6944,N_6753,N_6867);
nor U6945 (N_6945,N_6775,N_6797);
xor U6946 (N_6946,N_6840,N_6826);
and U6947 (N_6947,N_6772,N_6778);
or U6948 (N_6948,N_6822,N_6766);
or U6949 (N_6949,N_6857,N_6724);
or U6950 (N_6950,N_6777,N_6841);
or U6951 (N_6951,N_6748,N_6854);
and U6952 (N_6952,N_6848,N_6844);
and U6953 (N_6953,N_6839,N_6861);
nand U6954 (N_6954,N_6833,N_6758);
xor U6955 (N_6955,N_6735,N_6789);
or U6956 (N_6956,N_6847,N_6877);
xor U6957 (N_6957,N_6793,N_6805);
or U6958 (N_6958,N_6802,N_6773);
nor U6959 (N_6959,N_6737,N_6755);
and U6960 (N_6960,N_6756,N_6753);
nor U6961 (N_6961,N_6797,N_6828);
and U6962 (N_6962,N_6793,N_6759);
or U6963 (N_6963,N_6852,N_6750);
nor U6964 (N_6964,N_6744,N_6815);
nor U6965 (N_6965,N_6778,N_6834);
and U6966 (N_6966,N_6809,N_6862);
or U6967 (N_6967,N_6757,N_6725);
nor U6968 (N_6968,N_6742,N_6775);
or U6969 (N_6969,N_6875,N_6721);
nor U6970 (N_6970,N_6747,N_6737);
nand U6971 (N_6971,N_6750,N_6783);
or U6972 (N_6972,N_6798,N_6831);
xnor U6973 (N_6973,N_6794,N_6798);
or U6974 (N_6974,N_6806,N_6749);
and U6975 (N_6975,N_6829,N_6800);
or U6976 (N_6976,N_6876,N_6873);
and U6977 (N_6977,N_6868,N_6851);
and U6978 (N_6978,N_6778,N_6856);
nand U6979 (N_6979,N_6745,N_6775);
and U6980 (N_6980,N_6761,N_6805);
nand U6981 (N_6981,N_6842,N_6792);
nand U6982 (N_6982,N_6859,N_6752);
xor U6983 (N_6983,N_6818,N_6775);
nand U6984 (N_6984,N_6814,N_6787);
nor U6985 (N_6985,N_6791,N_6869);
and U6986 (N_6986,N_6817,N_6854);
nor U6987 (N_6987,N_6787,N_6878);
nor U6988 (N_6988,N_6794,N_6821);
xor U6989 (N_6989,N_6874,N_6830);
or U6990 (N_6990,N_6826,N_6853);
or U6991 (N_6991,N_6832,N_6876);
or U6992 (N_6992,N_6875,N_6806);
nor U6993 (N_6993,N_6779,N_6724);
xor U6994 (N_6994,N_6751,N_6828);
or U6995 (N_6995,N_6870,N_6726);
nor U6996 (N_6996,N_6752,N_6766);
or U6997 (N_6997,N_6730,N_6777);
nand U6998 (N_6998,N_6856,N_6799);
xnor U6999 (N_6999,N_6757,N_6811);
or U7000 (N_7000,N_6874,N_6776);
xor U7001 (N_7001,N_6781,N_6848);
nor U7002 (N_7002,N_6785,N_6798);
and U7003 (N_7003,N_6796,N_6739);
or U7004 (N_7004,N_6783,N_6769);
nand U7005 (N_7005,N_6822,N_6806);
xor U7006 (N_7006,N_6864,N_6795);
or U7007 (N_7007,N_6832,N_6763);
nand U7008 (N_7008,N_6741,N_6845);
xor U7009 (N_7009,N_6754,N_6764);
and U7010 (N_7010,N_6722,N_6846);
nand U7011 (N_7011,N_6778,N_6861);
or U7012 (N_7012,N_6759,N_6796);
xor U7013 (N_7013,N_6842,N_6730);
or U7014 (N_7014,N_6803,N_6857);
or U7015 (N_7015,N_6761,N_6851);
or U7016 (N_7016,N_6794,N_6812);
or U7017 (N_7017,N_6762,N_6796);
nor U7018 (N_7018,N_6867,N_6803);
nand U7019 (N_7019,N_6741,N_6818);
nor U7020 (N_7020,N_6856,N_6751);
xor U7021 (N_7021,N_6756,N_6734);
and U7022 (N_7022,N_6749,N_6809);
or U7023 (N_7023,N_6779,N_6877);
xnor U7024 (N_7024,N_6751,N_6734);
or U7025 (N_7025,N_6825,N_6748);
and U7026 (N_7026,N_6877,N_6750);
and U7027 (N_7027,N_6864,N_6745);
nand U7028 (N_7028,N_6813,N_6749);
nand U7029 (N_7029,N_6759,N_6867);
or U7030 (N_7030,N_6854,N_6855);
and U7031 (N_7031,N_6833,N_6845);
and U7032 (N_7032,N_6753,N_6848);
or U7033 (N_7033,N_6729,N_6837);
nor U7034 (N_7034,N_6810,N_6756);
nand U7035 (N_7035,N_6845,N_6757);
xor U7036 (N_7036,N_6860,N_6740);
xor U7037 (N_7037,N_6767,N_6758);
and U7038 (N_7038,N_6745,N_6721);
xnor U7039 (N_7039,N_6812,N_6750);
xnor U7040 (N_7040,N_7025,N_6937);
and U7041 (N_7041,N_7027,N_6958);
or U7042 (N_7042,N_6895,N_6894);
and U7043 (N_7043,N_6927,N_6943);
nand U7044 (N_7044,N_7020,N_6970);
xor U7045 (N_7045,N_6880,N_6977);
nor U7046 (N_7046,N_6948,N_6892);
or U7047 (N_7047,N_7005,N_6889);
and U7048 (N_7048,N_6964,N_7006);
or U7049 (N_7049,N_6941,N_7004);
and U7050 (N_7050,N_7026,N_7031);
nor U7051 (N_7051,N_6994,N_7023);
nor U7052 (N_7052,N_6966,N_6909);
xor U7053 (N_7053,N_7000,N_7034);
nor U7054 (N_7054,N_6979,N_7003);
or U7055 (N_7055,N_7028,N_6896);
and U7056 (N_7056,N_6899,N_6959);
nand U7057 (N_7057,N_7011,N_6933);
nand U7058 (N_7058,N_7001,N_7009);
nand U7059 (N_7059,N_6919,N_6939);
xor U7060 (N_7060,N_6913,N_7008);
xor U7061 (N_7061,N_7039,N_7015);
and U7062 (N_7062,N_6972,N_6984);
or U7063 (N_7063,N_6934,N_7035);
nor U7064 (N_7064,N_6921,N_6952);
or U7065 (N_7065,N_6942,N_6932);
and U7066 (N_7066,N_6949,N_7024);
and U7067 (N_7067,N_6882,N_6957);
nor U7068 (N_7068,N_6967,N_6950);
nor U7069 (N_7069,N_6980,N_6983);
and U7070 (N_7070,N_7016,N_7019);
xor U7071 (N_7071,N_6961,N_6993);
nor U7072 (N_7072,N_7029,N_6914);
xor U7073 (N_7073,N_6908,N_6885);
and U7074 (N_7074,N_6883,N_6881);
and U7075 (N_7075,N_6995,N_6965);
nand U7076 (N_7076,N_7022,N_6900);
xor U7077 (N_7077,N_7014,N_6886);
nand U7078 (N_7078,N_6951,N_6998);
and U7079 (N_7079,N_6955,N_6987);
nor U7080 (N_7080,N_6935,N_6944);
xor U7081 (N_7081,N_6911,N_7032);
nand U7082 (N_7082,N_6903,N_6923);
nor U7083 (N_7083,N_6905,N_6907);
nor U7084 (N_7084,N_7002,N_6985);
nor U7085 (N_7085,N_6891,N_7038);
nor U7086 (N_7086,N_6890,N_6929);
or U7087 (N_7087,N_7037,N_6904);
xnor U7088 (N_7088,N_7030,N_6947);
nand U7089 (N_7089,N_6924,N_6960);
and U7090 (N_7090,N_7036,N_6938);
nand U7091 (N_7091,N_6946,N_6975);
and U7092 (N_7092,N_6884,N_6969);
xor U7093 (N_7093,N_6974,N_6918);
xnor U7094 (N_7094,N_6930,N_7012);
xnor U7095 (N_7095,N_7017,N_6992);
nor U7096 (N_7096,N_6953,N_6954);
nand U7097 (N_7097,N_6997,N_6981);
or U7098 (N_7098,N_6915,N_6888);
nor U7099 (N_7099,N_6931,N_7021);
nor U7100 (N_7100,N_7018,N_6956);
nor U7101 (N_7101,N_7007,N_6916);
nor U7102 (N_7102,N_6945,N_6968);
xnor U7103 (N_7103,N_6973,N_6996);
xor U7104 (N_7104,N_6906,N_6990);
and U7105 (N_7105,N_6920,N_6912);
and U7106 (N_7106,N_6925,N_6898);
and U7107 (N_7107,N_6897,N_6902);
or U7108 (N_7108,N_6936,N_7033);
xor U7109 (N_7109,N_6926,N_6917);
and U7110 (N_7110,N_6986,N_6978);
nor U7111 (N_7111,N_6940,N_6963);
nand U7112 (N_7112,N_6988,N_6928);
and U7113 (N_7113,N_6887,N_6976);
or U7114 (N_7114,N_6893,N_7013);
or U7115 (N_7115,N_6971,N_6982);
nand U7116 (N_7116,N_6991,N_6901);
nor U7117 (N_7117,N_6999,N_6989);
nor U7118 (N_7118,N_7010,N_6962);
and U7119 (N_7119,N_6922,N_6910);
and U7120 (N_7120,N_6937,N_7030);
nor U7121 (N_7121,N_6934,N_6984);
or U7122 (N_7122,N_7006,N_6930);
and U7123 (N_7123,N_6949,N_6982);
and U7124 (N_7124,N_6988,N_7017);
and U7125 (N_7125,N_6999,N_6956);
nor U7126 (N_7126,N_6977,N_6920);
xor U7127 (N_7127,N_7018,N_7017);
nand U7128 (N_7128,N_6881,N_6922);
nor U7129 (N_7129,N_6887,N_6955);
xnor U7130 (N_7130,N_6921,N_7018);
and U7131 (N_7131,N_7038,N_6969);
and U7132 (N_7132,N_7032,N_6918);
and U7133 (N_7133,N_6962,N_7033);
and U7134 (N_7134,N_7034,N_7020);
xnor U7135 (N_7135,N_6945,N_6985);
xnor U7136 (N_7136,N_6936,N_6886);
nor U7137 (N_7137,N_6966,N_6948);
and U7138 (N_7138,N_6981,N_6915);
xnor U7139 (N_7139,N_6965,N_7035);
xor U7140 (N_7140,N_6975,N_6988);
and U7141 (N_7141,N_6902,N_6999);
nand U7142 (N_7142,N_7030,N_7031);
nor U7143 (N_7143,N_6880,N_6892);
and U7144 (N_7144,N_7022,N_7029);
xnor U7145 (N_7145,N_7016,N_6964);
nor U7146 (N_7146,N_6981,N_7037);
and U7147 (N_7147,N_7008,N_6970);
or U7148 (N_7148,N_7037,N_7000);
and U7149 (N_7149,N_6914,N_6892);
or U7150 (N_7150,N_6911,N_6941);
nor U7151 (N_7151,N_6979,N_6936);
nand U7152 (N_7152,N_6923,N_6953);
nand U7153 (N_7153,N_6983,N_6905);
nand U7154 (N_7154,N_6919,N_7007);
nor U7155 (N_7155,N_6940,N_6934);
xor U7156 (N_7156,N_6885,N_6994);
nor U7157 (N_7157,N_6887,N_6999);
xor U7158 (N_7158,N_6919,N_6929);
or U7159 (N_7159,N_6937,N_6968);
xor U7160 (N_7160,N_6885,N_7000);
and U7161 (N_7161,N_7007,N_6922);
or U7162 (N_7162,N_6966,N_6905);
and U7163 (N_7163,N_6928,N_7031);
nand U7164 (N_7164,N_7002,N_6998);
and U7165 (N_7165,N_6955,N_6978);
and U7166 (N_7166,N_7038,N_6894);
and U7167 (N_7167,N_6894,N_6982);
and U7168 (N_7168,N_6986,N_6962);
xnor U7169 (N_7169,N_6968,N_6959);
nor U7170 (N_7170,N_6987,N_6937);
nor U7171 (N_7171,N_6973,N_6901);
nor U7172 (N_7172,N_6954,N_6983);
nand U7173 (N_7173,N_6964,N_7021);
nand U7174 (N_7174,N_6901,N_6922);
nand U7175 (N_7175,N_7011,N_6881);
nand U7176 (N_7176,N_6971,N_7030);
nand U7177 (N_7177,N_6931,N_6897);
and U7178 (N_7178,N_6981,N_6911);
nand U7179 (N_7179,N_6988,N_6885);
and U7180 (N_7180,N_6996,N_7038);
nand U7181 (N_7181,N_6956,N_6932);
or U7182 (N_7182,N_6925,N_7035);
nor U7183 (N_7183,N_6890,N_6906);
nand U7184 (N_7184,N_7008,N_6907);
or U7185 (N_7185,N_6887,N_7011);
xnor U7186 (N_7186,N_6958,N_6903);
or U7187 (N_7187,N_6971,N_7001);
or U7188 (N_7188,N_6890,N_6983);
nor U7189 (N_7189,N_7003,N_6948);
xnor U7190 (N_7190,N_7010,N_6884);
xor U7191 (N_7191,N_6904,N_7016);
or U7192 (N_7192,N_7019,N_6999);
nand U7193 (N_7193,N_6899,N_6976);
or U7194 (N_7194,N_7021,N_7037);
nor U7195 (N_7195,N_7012,N_6927);
nor U7196 (N_7196,N_6932,N_7007);
xor U7197 (N_7197,N_6991,N_7018);
nand U7198 (N_7198,N_6923,N_6918);
and U7199 (N_7199,N_6962,N_6889);
and U7200 (N_7200,N_7055,N_7156);
nor U7201 (N_7201,N_7071,N_7087);
xnor U7202 (N_7202,N_7153,N_7118);
xnor U7203 (N_7203,N_7061,N_7143);
xnor U7204 (N_7204,N_7115,N_7050);
nor U7205 (N_7205,N_7127,N_7101);
nand U7206 (N_7206,N_7178,N_7180);
nor U7207 (N_7207,N_7167,N_7102);
nand U7208 (N_7208,N_7095,N_7058);
and U7209 (N_7209,N_7040,N_7150);
or U7210 (N_7210,N_7138,N_7179);
and U7211 (N_7211,N_7124,N_7199);
or U7212 (N_7212,N_7099,N_7163);
or U7213 (N_7213,N_7084,N_7152);
nand U7214 (N_7214,N_7186,N_7164);
nor U7215 (N_7215,N_7046,N_7129);
and U7216 (N_7216,N_7045,N_7073);
nand U7217 (N_7217,N_7159,N_7052);
xnor U7218 (N_7218,N_7145,N_7091);
xor U7219 (N_7219,N_7075,N_7113);
and U7220 (N_7220,N_7069,N_7169);
or U7221 (N_7221,N_7173,N_7122);
xor U7222 (N_7222,N_7047,N_7187);
nor U7223 (N_7223,N_7108,N_7165);
and U7224 (N_7224,N_7192,N_7133);
nand U7225 (N_7225,N_7147,N_7132);
or U7226 (N_7226,N_7111,N_7126);
and U7227 (N_7227,N_7080,N_7121);
or U7228 (N_7228,N_7086,N_7157);
nand U7229 (N_7229,N_7175,N_7104);
or U7230 (N_7230,N_7172,N_7181);
nor U7231 (N_7231,N_7131,N_7062);
or U7232 (N_7232,N_7161,N_7171);
and U7233 (N_7233,N_7096,N_7148);
and U7234 (N_7234,N_7144,N_7074);
or U7235 (N_7235,N_7160,N_7125);
or U7236 (N_7236,N_7154,N_7106);
xnor U7237 (N_7237,N_7198,N_7140);
or U7238 (N_7238,N_7098,N_7182);
and U7239 (N_7239,N_7112,N_7059);
nor U7240 (N_7240,N_7097,N_7066);
nand U7241 (N_7241,N_7130,N_7117);
nor U7242 (N_7242,N_7195,N_7142);
and U7243 (N_7243,N_7166,N_7170);
or U7244 (N_7244,N_7146,N_7056);
or U7245 (N_7245,N_7191,N_7094);
nand U7246 (N_7246,N_7105,N_7070);
or U7247 (N_7247,N_7107,N_7067);
nand U7248 (N_7248,N_7088,N_7188);
xor U7249 (N_7249,N_7193,N_7076);
or U7250 (N_7250,N_7064,N_7123);
or U7251 (N_7251,N_7119,N_7089);
xor U7252 (N_7252,N_7054,N_7065);
xor U7253 (N_7253,N_7158,N_7110);
nand U7254 (N_7254,N_7141,N_7139);
xnor U7255 (N_7255,N_7184,N_7063);
xor U7256 (N_7256,N_7149,N_7077);
xnor U7257 (N_7257,N_7083,N_7043);
xor U7258 (N_7258,N_7041,N_7197);
xnor U7259 (N_7259,N_7168,N_7044);
nor U7260 (N_7260,N_7151,N_7053);
xor U7261 (N_7261,N_7079,N_7177);
or U7262 (N_7262,N_7136,N_7090);
nor U7263 (N_7263,N_7174,N_7093);
and U7264 (N_7264,N_7116,N_7060);
nor U7265 (N_7265,N_7068,N_7103);
nand U7266 (N_7266,N_7185,N_7081);
nor U7267 (N_7267,N_7109,N_7194);
nand U7268 (N_7268,N_7162,N_7114);
or U7269 (N_7269,N_7092,N_7120);
nand U7270 (N_7270,N_7134,N_7072);
nor U7271 (N_7271,N_7082,N_7176);
or U7272 (N_7272,N_7057,N_7135);
or U7273 (N_7273,N_7137,N_7100);
nand U7274 (N_7274,N_7128,N_7078);
nand U7275 (N_7275,N_7190,N_7048);
xor U7276 (N_7276,N_7042,N_7155);
nand U7277 (N_7277,N_7183,N_7051);
and U7278 (N_7278,N_7189,N_7085);
or U7279 (N_7279,N_7049,N_7196);
nand U7280 (N_7280,N_7073,N_7144);
or U7281 (N_7281,N_7135,N_7177);
nand U7282 (N_7282,N_7159,N_7080);
nor U7283 (N_7283,N_7115,N_7116);
nand U7284 (N_7284,N_7050,N_7059);
nor U7285 (N_7285,N_7148,N_7185);
nor U7286 (N_7286,N_7177,N_7088);
xor U7287 (N_7287,N_7165,N_7129);
or U7288 (N_7288,N_7174,N_7146);
and U7289 (N_7289,N_7190,N_7042);
and U7290 (N_7290,N_7197,N_7134);
and U7291 (N_7291,N_7153,N_7158);
nand U7292 (N_7292,N_7071,N_7133);
nor U7293 (N_7293,N_7054,N_7051);
nor U7294 (N_7294,N_7116,N_7048);
or U7295 (N_7295,N_7063,N_7130);
nor U7296 (N_7296,N_7055,N_7069);
or U7297 (N_7297,N_7070,N_7180);
xor U7298 (N_7298,N_7116,N_7107);
and U7299 (N_7299,N_7089,N_7172);
xnor U7300 (N_7300,N_7067,N_7104);
xnor U7301 (N_7301,N_7191,N_7068);
nor U7302 (N_7302,N_7167,N_7148);
xor U7303 (N_7303,N_7051,N_7107);
and U7304 (N_7304,N_7050,N_7092);
xnor U7305 (N_7305,N_7199,N_7080);
or U7306 (N_7306,N_7101,N_7123);
nand U7307 (N_7307,N_7193,N_7059);
nand U7308 (N_7308,N_7164,N_7182);
xor U7309 (N_7309,N_7140,N_7065);
or U7310 (N_7310,N_7105,N_7051);
xor U7311 (N_7311,N_7181,N_7096);
xnor U7312 (N_7312,N_7193,N_7060);
nor U7313 (N_7313,N_7160,N_7115);
and U7314 (N_7314,N_7077,N_7096);
or U7315 (N_7315,N_7150,N_7115);
nor U7316 (N_7316,N_7081,N_7058);
nand U7317 (N_7317,N_7049,N_7127);
nor U7318 (N_7318,N_7076,N_7077);
nor U7319 (N_7319,N_7106,N_7178);
xor U7320 (N_7320,N_7178,N_7143);
or U7321 (N_7321,N_7085,N_7041);
nor U7322 (N_7322,N_7116,N_7139);
xnor U7323 (N_7323,N_7170,N_7129);
or U7324 (N_7324,N_7055,N_7173);
xnor U7325 (N_7325,N_7115,N_7088);
nor U7326 (N_7326,N_7150,N_7174);
xor U7327 (N_7327,N_7192,N_7072);
xor U7328 (N_7328,N_7178,N_7105);
and U7329 (N_7329,N_7180,N_7159);
and U7330 (N_7330,N_7100,N_7170);
xor U7331 (N_7331,N_7043,N_7185);
xnor U7332 (N_7332,N_7049,N_7138);
nand U7333 (N_7333,N_7128,N_7139);
xor U7334 (N_7334,N_7073,N_7100);
nor U7335 (N_7335,N_7096,N_7130);
or U7336 (N_7336,N_7106,N_7144);
nand U7337 (N_7337,N_7064,N_7156);
nor U7338 (N_7338,N_7048,N_7191);
nor U7339 (N_7339,N_7042,N_7196);
nand U7340 (N_7340,N_7041,N_7161);
or U7341 (N_7341,N_7042,N_7137);
nand U7342 (N_7342,N_7073,N_7093);
and U7343 (N_7343,N_7041,N_7128);
and U7344 (N_7344,N_7053,N_7092);
and U7345 (N_7345,N_7183,N_7122);
nand U7346 (N_7346,N_7142,N_7152);
nor U7347 (N_7347,N_7173,N_7069);
or U7348 (N_7348,N_7137,N_7077);
nor U7349 (N_7349,N_7189,N_7186);
xor U7350 (N_7350,N_7040,N_7049);
nor U7351 (N_7351,N_7083,N_7181);
and U7352 (N_7352,N_7182,N_7192);
or U7353 (N_7353,N_7066,N_7112);
and U7354 (N_7354,N_7138,N_7162);
xnor U7355 (N_7355,N_7104,N_7195);
or U7356 (N_7356,N_7188,N_7098);
xor U7357 (N_7357,N_7075,N_7060);
xor U7358 (N_7358,N_7113,N_7144);
xnor U7359 (N_7359,N_7154,N_7185);
nand U7360 (N_7360,N_7218,N_7313);
nand U7361 (N_7361,N_7331,N_7232);
or U7362 (N_7362,N_7231,N_7282);
and U7363 (N_7363,N_7341,N_7271);
xor U7364 (N_7364,N_7298,N_7201);
nor U7365 (N_7365,N_7322,N_7328);
and U7366 (N_7366,N_7250,N_7208);
or U7367 (N_7367,N_7343,N_7333);
or U7368 (N_7368,N_7294,N_7321);
and U7369 (N_7369,N_7327,N_7253);
nor U7370 (N_7370,N_7312,N_7292);
or U7371 (N_7371,N_7290,N_7257);
xor U7372 (N_7372,N_7222,N_7200);
and U7373 (N_7373,N_7269,N_7285);
and U7374 (N_7374,N_7265,N_7230);
or U7375 (N_7375,N_7238,N_7348);
and U7376 (N_7376,N_7239,N_7235);
and U7377 (N_7377,N_7284,N_7317);
and U7378 (N_7378,N_7288,N_7246);
and U7379 (N_7379,N_7309,N_7251);
or U7380 (N_7380,N_7261,N_7260);
nor U7381 (N_7381,N_7241,N_7338);
nand U7382 (N_7382,N_7283,N_7264);
and U7383 (N_7383,N_7248,N_7214);
and U7384 (N_7384,N_7259,N_7274);
or U7385 (N_7385,N_7217,N_7223);
or U7386 (N_7386,N_7273,N_7345);
or U7387 (N_7387,N_7306,N_7307);
or U7388 (N_7388,N_7209,N_7267);
nor U7389 (N_7389,N_7236,N_7354);
nor U7390 (N_7390,N_7330,N_7320);
nand U7391 (N_7391,N_7213,N_7359);
nor U7392 (N_7392,N_7226,N_7340);
xnor U7393 (N_7393,N_7229,N_7356);
and U7394 (N_7394,N_7324,N_7314);
and U7395 (N_7395,N_7352,N_7203);
nand U7396 (N_7396,N_7240,N_7323);
or U7397 (N_7397,N_7270,N_7207);
nor U7398 (N_7398,N_7210,N_7202);
and U7399 (N_7399,N_7268,N_7242);
nand U7400 (N_7400,N_7302,N_7278);
nor U7401 (N_7401,N_7256,N_7287);
and U7402 (N_7402,N_7311,N_7303);
xnor U7403 (N_7403,N_7219,N_7295);
or U7404 (N_7404,N_7332,N_7315);
xor U7405 (N_7405,N_7335,N_7216);
and U7406 (N_7406,N_7205,N_7351);
nor U7407 (N_7407,N_7289,N_7221);
or U7408 (N_7408,N_7224,N_7255);
xnor U7409 (N_7409,N_7225,N_7349);
nand U7410 (N_7410,N_7279,N_7275);
nand U7411 (N_7411,N_7308,N_7228);
nand U7412 (N_7412,N_7300,N_7249);
and U7413 (N_7413,N_7212,N_7245);
or U7414 (N_7414,N_7339,N_7318);
xnor U7415 (N_7415,N_7244,N_7297);
or U7416 (N_7416,N_7305,N_7234);
nand U7417 (N_7417,N_7350,N_7299);
or U7418 (N_7418,N_7304,N_7263);
nor U7419 (N_7419,N_7342,N_7206);
nand U7420 (N_7420,N_7204,N_7310);
and U7421 (N_7421,N_7291,N_7277);
or U7422 (N_7422,N_7334,N_7296);
and U7423 (N_7423,N_7227,N_7262);
xor U7424 (N_7424,N_7272,N_7286);
nand U7425 (N_7425,N_7266,N_7215);
or U7426 (N_7426,N_7252,N_7258);
nor U7427 (N_7427,N_7316,N_7254);
or U7428 (N_7428,N_7357,N_7329);
and U7429 (N_7429,N_7358,N_7220);
nor U7430 (N_7430,N_7276,N_7280);
nor U7431 (N_7431,N_7237,N_7233);
nor U7432 (N_7432,N_7326,N_7325);
nand U7433 (N_7433,N_7243,N_7301);
xnor U7434 (N_7434,N_7353,N_7344);
nor U7435 (N_7435,N_7336,N_7355);
or U7436 (N_7436,N_7211,N_7247);
nor U7437 (N_7437,N_7293,N_7346);
nor U7438 (N_7438,N_7337,N_7281);
nor U7439 (N_7439,N_7347,N_7319);
nor U7440 (N_7440,N_7350,N_7228);
xor U7441 (N_7441,N_7341,N_7333);
nand U7442 (N_7442,N_7266,N_7315);
nand U7443 (N_7443,N_7353,N_7331);
xnor U7444 (N_7444,N_7312,N_7227);
nor U7445 (N_7445,N_7321,N_7208);
nor U7446 (N_7446,N_7347,N_7236);
xnor U7447 (N_7447,N_7239,N_7340);
or U7448 (N_7448,N_7234,N_7275);
xor U7449 (N_7449,N_7332,N_7228);
nand U7450 (N_7450,N_7202,N_7330);
or U7451 (N_7451,N_7282,N_7358);
or U7452 (N_7452,N_7311,N_7253);
nor U7453 (N_7453,N_7220,N_7292);
nand U7454 (N_7454,N_7258,N_7279);
and U7455 (N_7455,N_7224,N_7234);
xor U7456 (N_7456,N_7301,N_7351);
or U7457 (N_7457,N_7348,N_7346);
nor U7458 (N_7458,N_7305,N_7215);
and U7459 (N_7459,N_7260,N_7304);
or U7460 (N_7460,N_7278,N_7267);
nor U7461 (N_7461,N_7320,N_7341);
xnor U7462 (N_7462,N_7252,N_7358);
and U7463 (N_7463,N_7280,N_7358);
and U7464 (N_7464,N_7207,N_7214);
xor U7465 (N_7465,N_7272,N_7266);
and U7466 (N_7466,N_7266,N_7345);
or U7467 (N_7467,N_7289,N_7234);
xor U7468 (N_7468,N_7255,N_7222);
xor U7469 (N_7469,N_7211,N_7205);
xnor U7470 (N_7470,N_7204,N_7234);
xor U7471 (N_7471,N_7230,N_7231);
and U7472 (N_7472,N_7336,N_7339);
xor U7473 (N_7473,N_7207,N_7290);
xor U7474 (N_7474,N_7250,N_7248);
nand U7475 (N_7475,N_7293,N_7269);
nor U7476 (N_7476,N_7342,N_7223);
and U7477 (N_7477,N_7212,N_7206);
and U7478 (N_7478,N_7206,N_7277);
nor U7479 (N_7479,N_7301,N_7252);
nand U7480 (N_7480,N_7311,N_7305);
nand U7481 (N_7481,N_7204,N_7239);
xnor U7482 (N_7482,N_7292,N_7224);
or U7483 (N_7483,N_7207,N_7321);
or U7484 (N_7484,N_7260,N_7312);
xnor U7485 (N_7485,N_7256,N_7251);
nand U7486 (N_7486,N_7236,N_7206);
and U7487 (N_7487,N_7275,N_7259);
nor U7488 (N_7488,N_7262,N_7230);
xnor U7489 (N_7489,N_7214,N_7255);
nor U7490 (N_7490,N_7227,N_7336);
and U7491 (N_7491,N_7250,N_7202);
or U7492 (N_7492,N_7354,N_7266);
and U7493 (N_7493,N_7258,N_7338);
nand U7494 (N_7494,N_7306,N_7345);
and U7495 (N_7495,N_7266,N_7281);
and U7496 (N_7496,N_7258,N_7326);
xnor U7497 (N_7497,N_7253,N_7283);
or U7498 (N_7498,N_7214,N_7312);
nor U7499 (N_7499,N_7290,N_7273);
or U7500 (N_7500,N_7207,N_7263);
nand U7501 (N_7501,N_7245,N_7261);
xor U7502 (N_7502,N_7336,N_7262);
nand U7503 (N_7503,N_7288,N_7282);
nor U7504 (N_7504,N_7264,N_7311);
xor U7505 (N_7505,N_7202,N_7281);
or U7506 (N_7506,N_7336,N_7247);
or U7507 (N_7507,N_7242,N_7273);
xnor U7508 (N_7508,N_7204,N_7274);
xor U7509 (N_7509,N_7260,N_7262);
or U7510 (N_7510,N_7350,N_7224);
xnor U7511 (N_7511,N_7350,N_7342);
and U7512 (N_7512,N_7262,N_7274);
and U7513 (N_7513,N_7245,N_7228);
nor U7514 (N_7514,N_7346,N_7272);
xnor U7515 (N_7515,N_7321,N_7231);
xnor U7516 (N_7516,N_7342,N_7332);
nand U7517 (N_7517,N_7249,N_7352);
nand U7518 (N_7518,N_7319,N_7327);
xor U7519 (N_7519,N_7324,N_7290);
nor U7520 (N_7520,N_7363,N_7481);
nand U7521 (N_7521,N_7453,N_7479);
or U7522 (N_7522,N_7503,N_7424);
nor U7523 (N_7523,N_7448,N_7394);
nor U7524 (N_7524,N_7421,N_7459);
or U7525 (N_7525,N_7402,N_7434);
or U7526 (N_7526,N_7413,N_7464);
nand U7527 (N_7527,N_7405,N_7447);
nand U7528 (N_7528,N_7371,N_7417);
nand U7529 (N_7529,N_7437,N_7468);
nand U7530 (N_7530,N_7399,N_7460);
or U7531 (N_7531,N_7418,N_7389);
nor U7532 (N_7532,N_7400,N_7515);
nor U7533 (N_7533,N_7375,N_7487);
or U7534 (N_7534,N_7452,N_7480);
and U7535 (N_7535,N_7461,N_7378);
nor U7536 (N_7536,N_7443,N_7469);
or U7537 (N_7537,N_7428,N_7438);
or U7538 (N_7538,N_7495,N_7426);
nor U7539 (N_7539,N_7384,N_7407);
or U7540 (N_7540,N_7387,N_7516);
or U7541 (N_7541,N_7411,N_7390);
nor U7542 (N_7542,N_7497,N_7466);
and U7543 (N_7543,N_7485,N_7456);
xor U7544 (N_7544,N_7444,N_7510);
xor U7545 (N_7545,N_7397,N_7431);
or U7546 (N_7546,N_7361,N_7360);
nand U7547 (N_7547,N_7395,N_7376);
or U7548 (N_7548,N_7398,N_7475);
nor U7549 (N_7549,N_7379,N_7490);
nand U7550 (N_7550,N_7500,N_7473);
xor U7551 (N_7551,N_7429,N_7436);
nor U7552 (N_7552,N_7442,N_7514);
and U7553 (N_7553,N_7446,N_7409);
xnor U7554 (N_7554,N_7440,N_7502);
and U7555 (N_7555,N_7435,N_7474);
and U7556 (N_7556,N_7372,N_7408);
and U7557 (N_7557,N_7385,N_7496);
nand U7558 (N_7558,N_7476,N_7513);
nor U7559 (N_7559,N_7369,N_7506);
xnor U7560 (N_7560,N_7454,N_7465);
xor U7561 (N_7561,N_7362,N_7494);
and U7562 (N_7562,N_7427,N_7511);
nand U7563 (N_7563,N_7470,N_7471);
nand U7564 (N_7564,N_7457,N_7463);
nand U7565 (N_7565,N_7396,N_7406);
nand U7566 (N_7566,N_7388,N_7462);
and U7567 (N_7567,N_7493,N_7374);
nor U7568 (N_7568,N_7404,N_7439);
or U7569 (N_7569,N_7489,N_7472);
nor U7570 (N_7570,N_7412,N_7482);
xor U7571 (N_7571,N_7365,N_7508);
xnor U7572 (N_7572,N_7370,N_7512);
nor U7573 (N_7573,N_7403,N_7451);
xnor U7574 (N_7574,N_7519,N_7380);
or U7575 (N_7575,N_7391,N_7455);
nand U7576 (N_7576,N_7393,N_7507);
and U7577 (N_7577,N_7501,N_7505);
nand U7578 (N_7578,N_7416,N_7483);
or U7579 (N_7579,N_7410,N_7386);
or U7580 (N_7580,N_7382,N_7419);
nor U7581 (N_7581,N_7367,N_7458);
nor U7582 (N_7582,N_7478,N_7420);
or U7583 (N_7583,N_7517,N_7377);
and U7584 (N_7584,N_7477,N_7491);
nand U7585 (N_7585,N_7432,N_7498);
xnor U7586 (N_7586,N_7518,N_7488);
or U7587 (N_7587,N_7509,N_7450);
nor U7588 (N_7588,N_7504,N_7441);
or U7589 (N_7589,N_7415,N_7368);
or U7590 (N_7590,N_7392,N_7364);
nand U7591 (N_7591,N_7433,N_7467);
or U7592 (N_7592,N_7449,N_7486);
or U7593 (N_7593,N_7422,N_7425);
and U7594 (N_7594,N_7423,N_7445);
and U7595 (N_7595,N_7366,N_7373);
and U7596 (N_7596,N_7414,N_7499);
or U7597 (N_7597,N_7381,N_7492);
or U7598 (N_7598,N_7430,N_7484);
or U7599 (N_7599,N_7383,N_7401);
and U7600 (N_7600,N_7387,N_7476);
nand U7601 (N_7601,N_7471,N_7518);
xnor U7602 (N_7602,N_7414,N_7481);
nor U7603 (N_7603,N_7470,N_7515);
xnor U7604 (N_7604,N_7371,N_7518);
or U7605 (N_7605,N_7459,N_7485);
or U7606 (N_7606,N_7415,N_7452);
xnor U7607 (N_7607,N_7428,N_7365);
xor U7608 (N_7608,N_7437,N_7389);
nor U7609 (N_7609,N_7455,N_7404);
and U7610 (N_7610,N_7444,N_7515);
nand U7611 (N_7611,N_7493,N_7366);
nor U7612 (N_7612,N_7445,N_7484);
xor U7613 (N_7613,N_7418,N_7425);
nor U7614 (N_7614,N_7516,N_7485);
nand U7615 (N_7615,N_7452,N_7417);
xnor U7616 (N_7616,N_7404,N_7480);
nand U7617 (N_7617,N_7472,N_7504);
xnor U7618 (N_7618,N_7384,N_7495);
or U7619 (N_7619,N_7518,N_7498);
or U7620 (N_7620,N_7424,N_7389);
or U7621 (N_7621,N_7487,N_7416);
xor U7622 (N_7622,N_7440,N_7474);
or U7623 (N_7623,N_7395,N_7385);
nand U7624 (N_7624,N_7498,N_7468);
or U7625 (N_7625,N_7429,N_7379);
and U7626 (N_7626,N_7453,N_7419);
nand U7627 (N_7627,N_7432,N_7455);
and U7628 (N_7628,N_7497,N_7474);
and U7629 (N_7629,N_7387,N_7375);
or U7630 (N_7630,N_7511,N_7461);
or U7631 (N_7631,N_7448,N_7396);
or U7632 (N_7632,N_7404,N_7486);
or U7633 (N_7633,N_7452,N_7493);
or U7634 (N_7634,N_7372,N_7435);
nand U7635 (N_7635,N_7457,N_7371);
xnor U7636 (N_7636,N_7399,N_7441);
or U7637 (N_7637,N_7443,N_7393);
xor U7638 (N_7638,N_7395,N_7432);
nand U7639 (N_7639,N_7405,N_7434);
and U7640 (N_7640,N_7386,N_7485);
and U7641 (N_7641,N_7404,N_7378);
xor U7642 (N_7642,N_7408,N_7425);
and U7643 (N_7643,N_7407,N_7433);
xor U7644 (N_7644,N_7401,N_7404);
nor U7645 (N_7645,N_7417,N_7512);
nand U7646 (N_7646,N_7387,N_7457);
or U7647 (N_7647,N_7472,N_7382);
nand U7648 (N_7648,N_7423,N_7363);
nor U7649 (N_7649,N_7437,N_7466);
nand U7650 (N_7650,N_7409,N_7440);
nor U7651 (N_7651,N_7453,N_7493);
or U7652 (N_7652,N_7380,N_7454);
xnor U7653 (N_7653,N_7513,N_7362);
nor U7654 (N_7654,N_7362,N_7499);
nand U7655 (N_7655,N_7399,N_7513);
or U7656 (N_7656,N_7408,N_7443);
nor U7657 (N_7657,N_7398,N_7463);
nor U7658 (N_7658,N_7442,N_7470);
and U7659 (N_7659,N_7492,N_7505);
and U7660 (N_7660,N_7376,N_7425);
nor U7661 (N_7661,N_7411,N_7441);
nor U7662 (N_7662,N_7469,N_7459);
and U7663 (N_7663,N_7445,N_7427);
and U7664 (N_7664,N_7381,N_7402);
nor U7665 (N_7665,N_7404,N_7379);
or U7666 (N_7666,N_7457,N_7411);
or U7667 (N_7667,N_7480,N_7492);
or U7668 (N_7668,N_7451,N_7408);
nor U7669 (N_7669,N_7361,N_7363);
xor U7670 (N_7670,N_7388,N_7474);
xor U7671 (N_7671,N_7368,N_7505);
nand U7672 (N_7672,N_7437,N_7425);
nand U7673 (N_7673,N_7370,N_7466);
nor U7674 (N_7674,N_7432,N_7465);
xor U7675 (N_7675,N_7362,N_7485);
or U7676 (N_7676,N_7453,N_7410);
xor U7677 (N_7677,N_7377,N_7450);
nor U7678 (N_7678,N_7420,N_7448);
nor U7679 (N_7679,N_7441,N_7494);
nand U7680 (N_7680,N_7611,N_7573);
and U7681 (N_7681,N_7564,N_7527);
or U7682 (N_7682,N_7531,N_7536);
xor U7683 (N_7683,N_7667,N_7670);
nand U7684 (N_7684,N_7594,N_7553);
or U7685 (N_7685,N_7577,N_7605);
or U7686 (N_7686,N_7547,N_7622);
xor U7687 (N_7687,N_7574,N_7650);
or U7688 (N_7688,N_7677,N_7628);
or U7689 (N_7689,N_7606,N_7627);
or U7690 (N_7690,N_7621,N_7642);
xor U7691 (N_7691,N_7539,N_7661);
xor U7692 (N_7692,N_7637,N_7619);
and U7693 (N_7693,N_7588,N_7595);
xor U7694 (N_7694,N_7676,N_7644);
nand U7695 (N_7695,N_7610,N_7585);
and U7696 (N_7696,N_7530,N_7623);
nand U7697 (N_7697,N_7598,N_7602);
or U7698 (N_7698,N_7571,N_7581);
xor U7699 (N_7699,N_7678,N_7630);
and U7700 (N_7700,N_7641,N_7674);
and U7701 (N_7701,N_7651,N_7659);
or U7702 (N_7702,N_7638,N_7616);
or U7703 (N_7703,N_7652,N_7620);
nand U7704 (N_7704,N_7523,N_7569);
nand U7705 (N_7705,N_7604,N_7657);
and U7706 (N_7706,N_7563,N_7525);
xor U7707 (N_7707,N_7656,N_7584);
nand U7708 (N_7708,N_7607,N_7566);
or U7709 (N_7709,N_7540,N_7590);
and U7710 (N_7710,N_7646,N_7636);
nand U7711 (N_7711,N_7561,N_7609);
nor U7712 (N_7712,N_7532,N_7624);
xor U7713 (N_7713,N_7649,N_7583);
nand U7714 (N_7714,N_7666,N_7662);
or U7715 (N_7715,N_7675,N_7664);
xnor U7716 (N_7716,N_7552,N_7555);
nand U7717 (N_7717,N_7669,N_7556);
or U7718 (N_7718,N_7615,N_7568);
nand U7719 (N_7719,N_7679,N_7520);
or U7720 (N_7720,N_7625,N_7632);
nor U7721 (N_7721,N_7586,N_7560);
or U7722 (N_7722,N_7597,N_7647);
or U7723 (N_7723,N_7591,N_7589);
nand U7724 (N_7724,N_7576,N_7645);
and U7725 (N_7725,N_7582,N_7565);
or U7726 (N_7726,N_7543,N_7640);
or U7727 (N_7727,N_7613,N_7596);
xnor U7728 (N_7728,N_7562,N_7551);
or U7729 (N_7729,N_7614,N_7528);
nand U7730 (N_7730,N_7592,N_7559);
or U7731 (N_7731,N_7660,N_7668);
xor U7732 (N_7732,N_7545,N_7626);
and U7733 (N_7733,N_7542,N_7618);
and U7734 (N_7734,N_7524,N_7541);
and U7735 (N_7735,N_7600,N_7575);
or U7736 (N_7736,N_7534,N_7634);
nor U7737 (N_7737,N_7554,N_7535);
nand U7738 (N_7738,N_7633,N_7673);
nor U7739 (N_7739,N_7631,N_7663);
xnor U7740 (N_7740,N_7558,N_7671);
or U7741 (N_7741,N_7579,N_7617);
and U7742 (N_7742,N_7544,N_7538);
nor U7743 (N_7743,N_7572,N_7612);
xnor U7744 (N_7744,N_7522,N_7557);
nor U7745 (N_7745,N_7548,N_7549);
nor U7746 (N_7746,N_7599,N_7635);
and U7747 (N_7747,N_7648,N_7665);
xnor U7748 (N_7748,N_7537,N_7643);
xor U7749 (N_7749,N_7601,N_7653);
and U7750 (N_7750,N_7550,N_7578);
nor U7751 (N_7751,N_7639,N_7546);
nor U7752 (N_7752,N_7580,N_7658);
or U7753 (N_7753,N_7521,N_7526);
nor U7754 (N_7754,N_7587,N_7593);
nor U7755 (N_7755,N_7567,N_7533);
or U7756 (N_7756,N_7629,N_7655);
or U7757 (N_7757,N_7654,N_7672);
or U7758 (N_7758,N_7608,N_7529);
nor U7759 (N_7759,N_7570,N_7603);
xnor U7760 (N_7760,N_7558,N_7568);
and U7761 (N_7761,N_7646,N_7658);
and U7762 (N_7762,N_7674,N_7604);
nand U7763 (N_7763,N_7659,N_7662);
nand U7764 (N_7764,N_7533,N_7566);
and U7765 (N_7765,N_7679,N_7534);
nand U7766 (N_7766,N_7652,N_7648);
xor U7767 (N_7767,N_7587,N_7619);
and U7768 (N_7768,N_7605,N_7521);
xnor U7769 (N_7769,N_7617,N_7639);
nand U7770 (N_7770,N_7525,N_7594);
nor U7771 (N_7771,N_7530,N_7643);
or U7772 (N_7772,N_7538,N_7575);
and U7773 (N_7773,N_7535,N_7533);
or U7774 (N_7774,N_7599,N_7612);
nor U7775 (N_7775,N_7551,N_7653);
xnor U7776 (N_7776,N_7549,N_7522);
nand U7777 (N_7777,N_7564,N_7590);
or U7778 (N_7778,N_7631,N_7671);
or U7779 (N_7779,N_7573,N_7638);
nand U7780 (N_7780,N_7616,N_7624);
nand U7781 (N_7781,N_7545,N_7675);
nor U7782 (N_7782,N_7538,N_7625);
nand U7783 (N_7783,N_7575,N_7626);
or U7784 (N_7784,N_7531,N_7666);
xnor U7785 (N_7785,N_7668,N_7546);
nand U7786 (N_7786,N_7663,N_7666);
or U7787 (N_7787,N_7621,N_7587);
and U7788 (N_7788,N_7647,N_7646);
or U7789 (N_7789,N_7538,N_7534);
xor U7790 (N_7790,N_7608,N_7599);
nor U7791 (N_7791,N_7564,N_7603);
xor U7792 (N_7792,N_7586,N_7650);
and U7793 (N_7793,N_7602,N_7660);
or U7794 (N_7794,N_7607,N_7637);
nor U7795 (N_7795,N_7542,N_7560);
xor U7796 (N_7796,N_7589,N_7631);
and U7797 (N_7797,N_7576,N_7539);
nor U7798 (N_7798,N_7622,N_7530);
or U7799 (N_7799,N_7587,N_7578);
and U7800 (N_7800,N_7663,N_7676);
nor U7801 (N_7801,N_7605,N_7574);
or U7802 (N_7802,N_7521,N_7659);
nand U7803 (N_7803,N_7550,N_7634);
xnor U7804 (N_7804,N_7574,N_7655);
nand U7805 (N_7805,N_7626,N_7544);
nor U7806 (N_7806,N_7554,N_7652);
or U7807 (N_7807,N_7597,N_7640);
xor U7808 (N_7808,N_7580,N_7570);
nor U7809 (N_7809,N_7677,N_7626);
or U7810 (N_7810,N_7649,N_7576);
xnor U7811 (N_7811,N_7627,N_7596);
nand U7812 (N_7812,N_7543,N_7592);
or U7813 (N_7813,N_7647,N_7531);
or U7814 (N_7814,N_7577,N_7568);
and U7815 (N_7815,N_7532,N_7576);
nor U7816 (N_7816,N_7563,N_7585);
xor U7817 (N_7817,N_7526,N_7614);
nor U7818 (N_7818,N_7666,N_7536);
or U7819 (N_7819,N_7623,N_7587);
xor U7820 (N_7820,N_7643,N_7653);
and U7821 (N_7821,N_7663,N_7645);
nand U7822 (N_7822,N_7579,N_7625);
and U7823 (N_7823,N_7597,N_7669);
xnor U7824 (N_7824,N_7650,N_7646);
and U7825 (N_7825,N_7679,N_7666);
nand U7826 (N_7826,N_7610,N_7606);
or U7827 (N_7827,N_7563,N_7659);
and U7828 (N_7828,N_7526,N_7673);
nand U7829 (N_7829,N_7599,N_7534);
or U7830 (N_7830,N_7611,N_7521);
xnor U7831 (N_7831,N_7520,N_7555);
nand U7832 (N_7832,N_7544,N_7520);
nor U7833 (N_7833,N_7675,N_7661);
nor U7834 (N_7834,N_7596,N_7663);
and U7835 (N_7835,N_7620,N_7550);
and U7836 (N_7836,N_7532,N_7643);
or U7837 (N_7837,N_7649,N_7548);
xnor U7838 (N_7838,N_7551,N_7622);
xnor U7839 (N_7839,N_7675,N_7672);
and U7840 (N_7840,N_7752,N_7832);
nor U7841 (N_7841,N_7827,N_7763);
or U7842 (N_7842,N_7804,N_7688);
or U7843 (N_7843,N_7825,N_7834);
xnor U7844 (N_7844,N_7720,N_7819);
or U7845 (N_7845,N_7811,N_7812);
and U7846 (N_7846,N_7707,N_7683);
nor U7847 (N_7847,N_7725,N_7754);
nand U7848 (N_7848,N_7830,N_7705);
nor U7849 (N_7849,N_7839,N_7799);
or U7850 (N_7850,N_7735,N_7787);
nor U7851 (N_7851,N_7822,N_7816);
xnor U7852 (N_7852,N_7691,N_7712);
nor U7853 (N_7853,N_7807,N_7794);
nand U7854 (N_7854,N_7802,N_7739);
or U7855 (N_7855,N_7779,N_7771);
xor U7856 (N_7856,N_7814,N_7744);
xor U7857 (N_7857,N_7758,N_7750);
nor U7858 (N_7858,N_7826,N_7701);
nor U7859 (N_7859,N_7784,N_7741);
xor U7860 (N_7860,N_7745,N_7737);
or U7861 (N_7861,N_7797,N_7680);
or U7862 (N_7862,N_7682,N_7789);
nand U7863 (N_7863,N_7767,N_7738);
xnor U7864 (N_7864,N_7690,N_7836);
nor U7865 (N_7865,N_7791,N_7709);
xnor U7866 (N_7866,N_7728,N_7694);
and U7867 (N_7867,N_7731,N_7716);
nand U7868 (N_7868,N_7717,N_7788);
or U7869 (N_7869,N_7740,N_7734);
nand U7870 (N_7870,N_7753,N_7743);
and U7871 (N_7871,N_7700,N_7782);
xnor U7872 (N_7872,N_7837,N_7747);
xnor U7873 (N_7873,N_7706,N_7761);
nand U7874 (N_7874,N_7838,N_7818);
or U7875 (N_7875,N_7724,N_7685);
nor U7876 (N_7876,N_7833,N_7684);
nand U7877 (N_7877,N_7775,N_7770);
and U7878 (N_7878,N_7813,N_7736);
and U7879 (N_7879,N_7764,N_7790);
or U7880 (N_7880,N_7697,N_7769);
xor U7881 (N_7881,N_7722,N_7803);
and U7882 (N_7882,N_7695,N_7783);
and U7883 (N_7883,N_7801,N_7773);
or U7884 (N_7884,N_7726,N_7687);
nand U7885 (N_7885,N_7828,N_7692);
and U7886 (N_7886,N_7792,N_7729);
nor U7887 (N_7887,N_7766,N_7686);
and U7888 (N_7888,N_7795,N_7681);
nor U7889 (N_7889,N_7806,N_7719);
and U7890 (N_7890,N_7808,N_7824);
nor U7891 (N_7891,N_7796,N_7702);
or U7892 (N_7892,N_7781,N_7708);
xnor U7893 (N_7893,N_7732,N_7730);
and U7894 (N_7894,N_7821,N_7746);
and U7895 (N_7895,N_7756,N_7698);
nand U7896 (N_7896,N_7786,N_7823);
and U7897 (N_7897,N_7815,N_7757);
and U7898 (N_7898,N_7809,N_7798);
and U7899 (N_7899,N_7772,N_7765);
and U7900 (N_7900,N_7714,N_7693);
xnor U7901 (N_7901,N_7748,N_7689);
or U7902 (N_7902,N_7800,N_7776);
xor U7903 (N_7903,N_7723,N_7835);
and U7904 (N_7904,N_7760,N_7696);
and U7905 (N_7905,N_7703,N_7749);
xnor U7906 (N_7906,N_7755,N_7727);
or U7907 (N_7907,N_7768,N_7810);
and U7908 (N_7908,N_7817,N_7733);
or U7909 (N_7909,N_7831,N_7805);
nor U7910 (N_7910,N_7713,N_7715);
xnor U7911 (N_7911,N_7704,N_7762);
xor U7912 (N_7912,N_7742,N_7751);
and U7913 (N_7913,N_7711,N_7721);
nand U7914 (N_7914,N_7777,N_7759);
or U7915 (N_7915,N_7774,N_7785);
or U7916 (N_7916,N_7829,N_7699);
nor U7917 (N_7917,N_7793,N_7820);
nand U7918 (N_7918,N_7718,N_7710);
nor U7919 (N_7919,N_7778,N_7780);
nand U7920 (N_7920,N_7789,N_7686);
nand U7921 (N_7921,N_7724,N_7787);
nand U7922 (N_7922,N_7711,N_7823);
xor U7923 (N_7923,N_7790,N_7716);
nand U7924 (N_7924,N_7813,N_7729);
nor U7925 (N_7925,N_7791,N_7796);
nand U7926 (N_7926,N_7729,N_7745);
nand U7927 (N_7927,N_7765,N_7809);
or U7928 (N_7928,N_7784,N_7775);
and U7929 (N_7929,N_7796,N_7706);
nand U7930 (N_7930,N_7690,N_7799);
or U7931 (N_7931,N_7755,N_7831);
and U7932 (N_7932,N_7707,N_7735);
xnor U7933 (N_7933,N_7826,N_7794);
and U7934 (N_7934,N_7763,N_7692);
nand U7935 (N_7935,N_7772,N_7777);
nand U7936 (N_7936,N_7771,N_7727);
nor U7937 (N_7937,N_7703,N_7766);
xnor U7938 (N_7938,N_7763,N_7716);
xnor U7939 (N_7939,N_7680,N_7817);
and U7940 (N_7940,N_7758,N_7732);
nor U7941 (N_7941,N_7740,N_7782);
nor U7942 (N_7942,N_7698,N_7703);
nor U7943 (N_7943,N_7816,N_7749);
and U7944 (N_7944,N_7783,N_7759);
and U7945 (N_7945,N_7767,N_7822);
and U7946 (N_7946,N_7805,N_7816);
and U7947 (N_7947,N_7720,N_7755);
nand U7948 (N_7948,N_7811,N_7713);
or U7949 (N_7949,N_7694,N_7746);
xnor U7950 (N_7950,N_7691,N_7725);
nand U7951 (N_7951,N_7787,N_7775);
or U7952 (N_7952,N_7723,N_7793);
and U7953 (N_7953,N_7684,N_7819);
nor U7954 (N_7954,N_7719,N_7810);
nor U7955 (N_7955,N_7812,N_7704);
xor U7956 (N_7956,N_7779,N_7688);
or U7957 (N_7957,N_7808,N_7684);
and U7958 (N_7958,N_7809,N_7801);
xnor U7959 (N_7959,N_7773,N_7804);
nor U7960 (N_7960,N_7751,N_7836);
nand U7961 (N_7961,N_7823,N_7798);
and U7962 (N_7962,N_7770,N_7757);
xor U7963 (N_7963,N_7760,N_7758);
xor U7964 (N_7964,N_7807,N_7698);
or U7965 (N_7965,N_7723,N_7688);
xnor U7966 (N_7966,N_7741,N_7731);
and U7967 (N_7967,N_7790,N_7721);
nor U7968 (N_7968,N_7767,N_7776);
or U7969 (N_7969,N_7808,N_7756);
xnor U7970 (N_7970,N_7831,N_7832);
xnor U7971 (N_7971,N_7784,N_7808);
xor U7972 (N_7972,N_7764,N_7716);
xor U7973 (N_7973,N_7710,N_7725);
nor U7974 (N_7974,N_7834,N_7804);
or U7975 (N_7975,N_7683,N_7777);
nand U7976 (N_7976,N_7743,N_7795);
xor U7977 (N_7977,N_7831,N_7766);
nor U7978 (N_7978,N_7785,N_7768);
or U7979 (N_7979,N_7814,N_7780);
nand U7980 (N_7980,N_7788,N_7752);
xor U7981 (N_7981,N_7838,N_7731);
and U7982 (N_7982,N_7701,N_7712);
nor U7983 (N_7983,N_7825,N_7751);
nor U7984 (N_7984,N_7736,N_7775);
and U7985 (N_7985,N_7830,N_7834);
xnor U7986 (N_7986,N_7754,N_7684);
and U7987 (N_7987,N_7784,N_7812);
nand U7988 (N_7988,N_7734,N_7825);
or U7989 (N_7989,N_7737,N_7790);
and U7990 (N_7990,N_7746,N_7711);
or U7991 (N_7991,N_7806,N_7788);
and U7992 (N_7992,N_7687,N_7689);
xor U7993 (N_7993,N_7722,N_7734);
and U7994 (N_7994,N_7773,N_7833);
nor U7995 (N_7995,N_7697,N_7725);
and U7996 (N_7996,N_7716,N_7753);
nor U7997 (N_7997,N_7763,N_7762);
nor U7998 (N_7998,N_7768,N_7737);
or U7999 (N_7999,N_7703,N_7779);
or U8000 (N_8000,N_7930,N_7894);
nor U8001 (N_8001,N_7969,N_7867);
nor U8002 (N_8002,N_7879,N_7875);
and U8003 (N_8003,N_7948,N_7863);
and U8004 (N_8004,N_7874,N_7895);
and U8005 (N_8005,N_7960,N_7962);
or U8006 (N_8006,N_7887,N_7847);
and U8007 (N_8007,N_7936,N_7876);
nor U8008 (N_8008,N_7989,N_7952);
or U8009 (N_8009,N_7956,N_7888);
nand U8010 (N_8010,N_7853,N_7920);
nand U8011 (N_8011,N_7859,N_7893);
or U8012 (N_8012,N_7951,N_7983);
nand U8013 (N_8013,N_7923,N_7844);
nand U8014 (N_8014,N_7947,N_7987);
nor U8015 (N_8015,N_7881,N_7885);
xor U8016 (N_8016,N_7850,N_7896);
or U8017 (N_8017,N_7916,N_7858);
nor U8018 (N_8018,N_7998,N_7890);
or U8019 (N_8019,N_7946,N_7980);
and U8020 (N_8020,N_7979,N_7883);
nand U8021 (N_8021,N_7984,N_7981);
or U8022 (N_8022,N_7900,N_7935);
nor U8023 (N_8023,N_7907,N_7878);
xor U8024 (N_8024,N_7910,N_7843);
nand U8025 (N_8025,N_7848,N_7868);
or U8026 (N_8026,N_7892,N_7889);
xor U8027 (N_8027,N_7912,N_7938);
nor U8028 (N_8028,N_7995,N_7841);
xnor U8029 (N_8029,N_7957,N_7925);
nand U8030 (N_8030,N_7922,N_7954);
nor U8031 (N_8031,N_7880,N_7861);
xnor U8032 (N_8032,N_7917,N_7905);
nor U8033 (N_8033,N_7985,N_7919);
xor U8034 (N_8034,N_7908,N_7852);
xor U8035 (N_8035,N_7891,N_7904);
nor U8036 (N_8036,N_7988,N_7871);
nand U8037 (N_8037,N_7967,N_7903);
nor U8038 (N_8038,N_7856,N_7991);
nand U8039 (N_8039,N_7924,N_7864);
or U8040 (N_8040,N_7884,N_7928);
and U8041 (N_8041,N_7877,N_7972);
nand U8042 (N_8042,N_7975,N_7950);
or U8043 (N_8043,N_7986,N_7932);
nor U8044 (N_8044,N_7913,N_7971);
or U8045 (N_8045,N_7933,N_7978);
xnor U8046 (N_8046,N_7921,N_7939);
xor U8047 (N_8047,N_7965,N_7997);
or U8048 (N_8048,N_7973,N_7845);
or U8049 (N_8049,N_7992,N_7964);
xnor U8050 (N_8050,N_7993,N_7943);
or U8051 (N_8051,N_7840,N_7902);
or U8052 (N_8052,N_7918,N_7970);
xnor U8053 (N_8053,N_7842,N_7857);
nand U8054 (N_8054,N_7909,N_7977);
nor U8055 (N_8055,N_7851,N_7994);
nand U8056 (N_8056,N_7914,N_7849);
or U8057 (N_8057,N_7897,N_7942);
or U8058 (N_8058,N_7869,N_7882);
xor U8059 (N_8059,N_7931,N_7860);
xor U8060 (N_8060,N_7898,N_7899);
nand U8061 (N_8061,N_7865,N_7944);
nor U8062 (N_8062,N_7955,N_7866);
and U8063 (N_8063,N_7982,N_7934);
or U8064 (N_8064,N_7945,N_7937);
or U8065 (N_8065,N_7873,N_7974);
xor U8066 (N_8066,N_7926,N_7901);
xor U8067 (N_8067,N_7959,N_7958);
xnor U8068 (N_8068,N_7940,N_7929);
or U8069 (N_8069,N_7996,N_7872);
and U8070 (N_8070,N_7963,N_7886);
and U8071 (N_8071,N_7855,N_7961);
xnor U8072 (N_8072,N_7953,N_7915);
nor U8073 (N_8073,N_7968,N_7854);
and U8074 (N_8074,N_7976,N_7906);
nor U8075 (N_8075,N_7862,N_7990);
and U8076 (N_8076,N_7966,N_7941);
xnor U8077 (N_8077,N_7911,N_7846);
or U8078 (N_8078,N_7870,N_7927);
nand U8079 (N_8079,N_7949,N_7999);
and U8080 (N_8080,N_7963,N_7999);
or U8081 (N_8081,N_7844,N_7955);
nand U8082 (N_8082,N_7950,N_7909);
xnor U8083 (N_8083,N_7993,N_7900);
nand U8084 (N_8084,N_7945,N_7949);
nand U8085 (N_8085,N_7927,N_7910);
nand U8086 (N_8086,N_7964,N_7925);
xnor U8087 (N_8087,N_7892,N_7878);
or U8088 (N_8088,N_7920,N_7871);
nor U8089 (N_8089,N_7871,N_7980);
or U8090 (N_8090,N_7886,N_7987);
nor U8091 (N_8091,N_7980,N_7956);
or U8092 (N_8092,N_7947,N_7990);
and U8093 (N_8093,N_7872,N_7910);
nor U8094 (N_8094,N_7877,N_7949);
nand U8095 (N_8095,N_7992,N_7989);
xnor U8096 (N_8096,N_7933,N_7971);
and U8097 (N_8097,N_7990,N_7930);
xor U8098 (N_8098,N_7967,N_7976);
xnor U8099 (N_8099,N_7860,N_7993);
or U8100 (N_8100,N_7998,N_7970);
xnor U8101 (N_8101,N_7941,N_7908);
nor U8102 (N_8102,N_7895,N_7889);
nor U8103 (N_8103,N_7848,N_7882);
nand U8104 (N_8104,N_7908,N_7841);
or U8105 (N_8105,N_7965,N_7891);
nor U8106 (N_8106,N_7851,N_7972);
or U8107 (N_8107,N_7866,N_7929);
or U8108 (N_8108,N_7899,N_7936);
nand U8109 (N_8109,N_7980,N_7922);
and U8110 (N_8110,N_7941,N_7857);
nor U8111 (N_8111,N_7878,N_7977);
nand U8112 (N_8112,N_7871,N_7955);
or U8113 (N_8113,N_7855,N_7896);
and U8114 (N_8114,N_7918,N_7892);
or U8115 (N_8115,N_7956,N_7951);
and U8116 (N_8116,N_7972,N_7938);
or U8117 (N_8117,N_7851,N_7871);
or U8118 (N_8118,N_7862,N_7917);
or U8119 (N_8119,N_7906,N_7873);
and U8120 (N_8120,N_7901,N_7956);
nor U8121 (N_8121,N_7860,N_7949);
and U8122 (N_8122,N_7947,N_7950);
and U8123 (N_8123,N_7926,N_7871);
or U8124 (N_8124,N_7913,N_7895);
and U8125 (N_8125,N_7865,N_7882);
or U8126 (N_8126,N_7902,N_7845);
xor U8127 (N_8127,N_7893,N_7941);
nor U8128 (N_8128,N_7947,N_7943);
and U8129 (N_8129,N_7993,N_7921);
or U8130 (N_8130,N_7959,N_7995);
or U8131 (N_8131,N_7882,N_7871);
or U8132 (N_8132,N_7970,N_7957);
nand U8133 (N_8133,N_7953,N_7938);
nor U8134 (N_8134,N_7863,N_7883);
and U8135 (N_8135,N_7882,N_7917);
or U8136 (N_8136,N_7947,N_7883);
or U8137 (N_8137,N_7951,N_7844);
nand U8138 (N_8138,N_7963,N_7869);
nand U8139 (N_8139,N_7930,N_7864);
or U8140 (N_8140,N_7845,N_7877);
or U8141 (N_8141,N_7931,N_7977);
nand U8142 (N_8142,N_7959,N_7996);
or U8143 (N_8143,N_7982,N_7841);
nor U8144 (N_8144,N_7872,N_7988);
nand U8145 (N_8145,N_7980,N_7895);
nor U8146 (N_8146,N_7937,N_7982);
and U8147 (N_8147,N_7993,N_7970);
nor U8148 (N_8148,N_7999,N_7905);
xnor U8149 (N_8149,N_7951,N_7930);
and U8150 (N_8150,N_7928,N_7859);
nand U8151 (N_8151,N_7927,N_7889);
xnor U8152 (N_8152,N_7892,N_7920);
or U8153 (N_8153,N_7957,N_7918);
and U8154 (N_8154,N_7841,N_7899);
nand U8155 (N_8155,N_7858,N_7932);
and U8156 (N_8156,N_7953,N_7894);
and U8157 (N_8157,N_7929,N_7946);
nand U8158 (N_8158,N_7992,N_7927);
nand U8159 (N_8159,N_7950,N_7994);
xnor U8160 (N_8160,N_8056,N_8071);
xnor U8161 (N_8161,N_8020,N_8095);
or U8162 (N_8162,N_8128,N_8016);
and U8163 (N_8163,N_8048,N_8066);
and U8164 (N_8164,N_8011,N_8129);
or U8165 (N_8165,N_8030,N_8050);
nor U8166 (N_8166,N_8058,N_8151);
or U8167 (N_8167,N_8049,N_8127);
nand U8168 (N_8168,N_8099,N_8035);
and U8169 (N_8169,N_8087,N_8106);
xor U8170 (N_8170,N_8122,N_8069);
nor U8171 (N_8171,N_8021,N_8028);
nand U8172 (N_8172,N_8076,N_8144);
and U8173 (N_8173,N_8132,N_8065);
and U8174 (N_8174,N_8155,N_8159);
nand U8175 (N_8175,N_8022,N_8033);
nand U8176 (N_8176,N_8001,N_8133);
xor U8177 (N_8177,N_8123,N_8039);
xor U8178 (N_8178,N_8027,N_8024);
xnor U8179 (N_8179,N_8103,N_8079);
or U8180 (N_8180,N_8114,N_8112);
nand U8181 (N_8181,N_8002,N_8148);
xnor U8182 (N_8182,N_8052,N_8067);
nand U8183 (N_8183,N_8149,N_8141);
and U8184 (N_8184,N_8029,N_8038);
or U8185 (N_8185,N_8060,N_8040);
nand U8186 (N_8186,N_8037,N_8094);
and U8187 (N_8187,N_8131,N_8117);
and U8188 (N_8188,N_8135,N_8009);
or U8189 (N_8189,N_8104,N_8089);
xor U8190 (N_8190,N_8000,N_8010);
and U8191 (N_8191,N_8093,N_8057);
xnor U8192 (N_8192,N_8088,N_8047);
and U8193 (N_8193,N_8018,N_8108);
or U8194 (N_8194,N_8072,N_8098);
nand U8195 (N_8195,N_8143,N_8032);
nor U8196 (N_8196,N_8077,N_8019);
and U8197 (N_8197,N_8115,N_8031);
nor U8198 (N_8198,N_8078,N_8005);
and U8199 (N_8199,N_8041,N_8012);
nor U8200 (N_8200,N_8017,N_8102);
or U8201 (N_8201,N_8053,N_8097);
or U8202 (N_8202,N_8084,N_8013);
xnor U8203 (N_8203,N_8147,N_8157);
nor U8204 (N_8204,N_8063,N_8119);
and U8205 (N_8205,N_8139,N_8026);
nor U8206 (N_8206,N_8105,N_8023);
or U8207 (N_8207,N_8015,N_8156);
or U8208 (N_8208,N_8107,N_8025);
xnor U8209 (N_8209,N_8046,N_8140);
nor U8210 (N_8210,N_8064,N_8154);
nand U8211 (N_8211,N_8134,N_8138);
xnor U8212 (N_8212,N_8090,N_8153);
nor U8213 (N_8213,N_8113,N_8003);
or U8214 (N_8214,N_8130,N_8006);
and U8215 (N_8215,N_8074,N_8062);
and U8216 (N_8216,N_8096,N_8075);
or U8217 (N_8217,N_8083,N_8121);
xor U8218 (N_8218,N_8124,N_8142);
nor U8219 (N_8219,N_8100,N_8126);
xor U8220 (N_8220,N_8061,N_8158);
xor U8221 (N_8221,N_8152,N_8118);
nor U8222 (N_8222,N_8101,N_8073);
nand U8223 (N_8223,N_8081,N_8110);
or U8224 (N_8224,N_8004,N_8109);
nand U8225 (N_8225,N_8085,N_8014);
xor U8226 (N_8226,N_8042,N_8120);
and U8227 (N_8227,N_8086,N_8059);
xnor U8228 (N_8228,N_8007,N_8137);
xor U8229 (N_8229,N_8125,N_8043);
or U8230 (N_8230,N_8045,N_8068);
nor U8231 (N_8231,N_8008,N_8082);
or U8232 (N_8232,N_8111,N_8054);
nor U8233 (N_8233,N_8150,N_8055);
xor U8234 (N_8234,N_8070,N_8080);
nand U8235 (N_8235,N_8145,N_8036);
or U8236 (N_8236,N_8034,N_8136);
nor U8237 (N_8237,N_8051,N_8091);
and U8238 (N_8238,N_8092,N_8044);
and U8239 (N_8239,N_8146,N_8116);
xnor U8240 (N_8240,N_8102,N_8044);
nand U8241 (N_8241,N_8080,N_8123);
nand U8242 (N_8242,N_8078,N_8054);
and U8243 (N_8243,N_8029,N_8094);
xnor U8244 (N_8244,N_8042,N_8141);
or U8245 (N_8245,N_8021,N_8118);
nand U8246 (N_8246,N_8045,N_8041);
and U8247 (N_8247,N_8033,N_8039);
nor U8248 (N_8248,N_8083,N_8155);
and U8249 (N_8249,N_8011,N_8139);
or U8250 (N_8250,N_8077,N_8065);
and U8251 (N_8251,N_8111,N_8098);
nand U8252 (N_8252,N_8128,N_8079);
nor U8253 (N_8253,N_8107,N_8143);
nor U8254 (N_8254,N_8151,N_8044);
or U8255 (N_8255,N_8020,N_8050);
and U8256 (N_8256,N_8032,N_8084);
xor U8257 (N_8257,N_8110,N_8036);
xor U8258 (N_8258,N_8037,N_8009);
nor U8259 (N_8259,N_8054,N_8029);
xor U8260 (N_8260,N_8024,N_8084);
or U8261 (N_8261,N_8019,N_8057);
or U8262 (N_8262,N_8008,N_8052);
nand U8263 (N_8263,N_8032,N_8099);
and U8264 (N_8264,N_8146,N_8097);
and U8265 (N_8265,N_8035,N_8119);
nand U8266 (N_8266,N_8022,N_8138);
and U8267 (N_8267,N_8061,N_8040);
xnor U8268 (N_8268,N_8115,N_8076);
xor U8269 (N_8269,N_8043,N_8106);
or U8270 (N_8270,N_8057,N_8107);
xnor U8271 (N_8271,N_8075,N_8095);
nand U8272 (N_8272,N_8004,N_8133);
nor U8273 (N_8273,N_8100,N_8127);
or U8274 (N_8274,N_8003,N_8013);
nor U8275 (N_8275,N_8100,N_8059);
and U8276 (N_8276,N_8068,N_8115);
xor U8277 (N_8277,N_8119,N_8073);
or U8278 (N_8278,N_8149,N_8115);
xor U8279 (N_8279,N_8118,N_8033);
or U8280 (N_8280,N_8028,N_8141);
nand U8281 (N_8281,N_8022,N_8038);
nand U8282 (N_8282,N_8074,N_8150);
xor U8283 (N_8283,N_8054,N_8075);
xor U8284 (N_8284,N_8132,N_8070);
and U8285 (N_8285,N_8031,N_8079);
xnor U8286 (N_8286,N_8145,N_8102);
and U8287 (N_8287,N_8003,N_8102);
nor U8288 (N_8288,N_8041,N_8032);
and U8289 (N_8289,N_8123,N_8007);
or U8290 (N_8290,N_8031,N_8157);
nor U8291 (N_8291,N_8090,N_8140);
nand U8292 (N_8292,N_8153,N_8059);
or U8293 (N_8293,N_8150,N_8090);
nand U8294 (N_8294,N_8024,N_8149);
and U8295 (N_8295,N_8062,N_8004);
xor U8296 (N_8296,N_8117,N_8020);
or U8297 (N_8297,N_8006,N_8092);
nor U8298 (N_8298,N_8095,N_8130);
and U8299 (N_8299,N_8100,N_8129);
xnor U8300 (N_8300,N_8112,N_8125);
xor U8301 (N_8301,N_8007,N_8091);
or U8302 (N_8302,N_8128,N_8049);
xnor U8303 (N_8303,N_8085,N_8059);
or U8304 (N_8304,N_8129,N_8060);
xor U8305 (N_8305,N_8054,N_8040);
nor U8306 (N_8306,N_8009,N_8128);
nor U8307 (N_8307,N_8067,N_8151);
or U8308 (N_8308,N_8108,N_8134);
nand U8309 (N_8309,N_8153,N_8088);
nor U8310 (N_8310,N_8109,N_8046);
and U8311 (N_8311,N_8017,N_8111);
nor U8312 (N_8312,N_8022,N_8083);
nand U8313 (N_8313,N_8058,N_8054);
or U8314 (N_8314,N_8150,N_8130);
or U8315 (N_8315,N_8026,N_8002);
nor U8316 (N_8316,N_8037,N_8127);
and U8317 (N_8317,N_8009,N_8114);
and U8318 (N_8318,N_8027,N_8125);
nand U8319 (N_8319,N_8073,N_8106);
and U8320 (N_8320,N_8227,N_8311);
nor U8321 (N_8321,N_8235,N_8212);
nor U8322 (N_8322,N_8228,N_8248);
nor U8323 (N_8323,N_8195,N_8202);
nor U8324 (N_8324,N_8167,N_8260);
xor U8325 (N_8325,N_8190,N_8205);
and U8326 (N_8326,N_8261,N_8225);
or U8327 (N_8327,N_8312,N_8299);
xor U8328 (N_8328,N_8296,N_8279);
nor U8329 (N_8329,N_8174,N_8181);
or U8330 (N_8330,N_8295,N_8274);
and U8331 (N_8331,N_8307,N_8276);
nor U8332 (N_8332,N_8189,N_8303);
or U8333 (N_8333,N_8229,N_8291);
nand U8334 (N_8334,N_8187,N_8314);
nor U8335 (N_8335,N_8270,N_8188);
xnor U8336 (N_8336,N_8161,N_8170);
nand U8337 (N_8337,N_8317,N_8297);
and U8338 (N_8338,N_8253,N_8176);
nor U8339 (N_8339,N_8204,N_8237);
nand U8340 (N_8340,N_8263,N_8254);
xnor U8341 (N_8341,N_8268,N_8293);
or U8342 (N_8342,N_8177,N_8209);
nand U8343 (N_8343,N_8304,N_8316);
or U8344 (N_8344,N_8232,N_8319);
xor U8345 (N_8345,N_8172,N_8219);
xor U8346 (N_8346,N_8288,N_8192);
and U8347 (N_8347,N_8179,N_8160);
or U8348 (N_8348,N_8271,N_8309);
xor U8349 (N_8349,N_8182,N_8216);
and U8350 (N_8350,N_8285,N_8221);
nor U8351 (N_8351,N_8186,N_8223);
nand U8352 (N_8352,N_8166,N_8163);
nand U8353 (N_8353,N_8290,N_8215);
nor U8354 (N_8354,N_8220,N_8218);
xnor U8355 (N_8355,N_8208,N_8214);
xnor U8356 (N_8356,N_8287,N_8178);
nand U8357 (N_8357,N_8318,N_8191);
nand U8358 (N_8358,N_8213,N_8245);
or U8359 (N_8359,N_8247,N_8238);
or U8360 (N_8360,N_8206,N_8203);
nand U8361 (N_8361,N_8284,N_8301);
nand U8362 (N_8362,N_8257,N_8164);
nor U8363 (N_8363,N_8241,N_8175);
xnor U8364 (N_8364,N_8226,N_8173);
nor U8365 (N_8365,N_8242,N_8306);
and U8366 (N_8366,N_8267,N_8162);
xnor U8367 (N_8367,N_8244,N_8243);
and U8368 (N_8368,N_8250,N_8278);
xor U8369 (N_8369,N_8255,N_8280);
or U8370 (N_8370,N_8310,N_8193);
nand U8371 (N_8371,N_8222,N_8198);
or U8372 (N_8372,N_8275,N_8252);
nand U8373 (N_8373,N_8169,N_8281);
and U8374 (N_8374,N_8183,N_8256);
nor U8375 (N_8375,N_8294,N_8300);
nor U8376 (N_8376,N_8308,N_8185);
xnor U8377 (N_8377,N_8233,N_8194);
nand U8378 (N_8378,N_8302,N_8230);
and U8379 (N_8379,N_8234,N_8211);
or U8380 (N_8380,N_8283,N_8289);
and U8381 (N_8381,N_8246,N_8266);
xnor U8382 (N_8382,N_8207,N_8292);
or U8383 (N_8383,N_8249,N_8262);
or U8384 (N_8384,N_8200,N_8282);
nor U8385 (N_8385,N_8277,N_8240);
or U8386 (N_8386,N_8286,N_8196);
and U8387 (N_8387,N_8305,N_8180);
nand U8388 (N_8388,N_8197,N_8315);
xor U8389 (N_8389,N_8168,N_8210);
or U8390 (N_8390,N_8224,N_8272);
or U8391 (N_8391,N_8171,N_8201);
and U8392 (N_8392,N_8298,N_8269);
or U8393 (N_8393,N_8313,N_8273);
nor U8394 (N_8394,N_8265,N_8236);
and U8395 (N_8395,N_8264,N_8184);
or U8396 (N_8396,N_8239,N_8199);
and U8397 (N_8397,N_8259,N_8231);
and U8398 (N_8398,N_8165,N_8258);
or U8399 (N_8399,N_8217,N_8251);
nor U8400 (N_8400,N_8317,N_8160);
xnor U8401 (N_8401,N_8213,N_8190);
and U8402 (N_8402,N_8307,N_8251);
nand U8403 (N_8403,N_8223,N_8295);
nor U8404 (N_8404,N_8251,N_8233);
and U8405 (N_8405,N_8298,N_8230);
xnor U8406 (N_8406,N_8203,N_8178);
nor U8407 (N_8407,N_8179,N_8241);
nor U8408 (N_8408,N_8198,N_8303);
xor U8409 (N_8409,N_8194,N_8187);
nand U8410 (N_8410,N_8206,N_8257);
nand U8411 (N_8411,N_8318,N_8250);
or U8412 (N_8412,N_8242,N_8316);
and U8413 (N_8413,N_8236,N_8287);
nor U8414 (N_8414,N_8174,N_8317);
and U8415 (N_8415,N_8208,N_8180);
and U8416 (N_8416,N_8243,N_8214);
or U8417 (N_8417,N_8295,N_8177);
or U8418 (N_8418,N_8180,N_8190);
or U8419 (N_8419,N_8218,N_8232);
and U8420 (N_8420,N_8257,N_8292);
nand U8421 (N_8421,N_8190,N_8259);
or U8422 (N_8422,N_8238,N_8271);
nor U8423 (N_8423,N_8312,N_8257);
nor U8424 (N_8424,N_8294,N_8277);
xor U8425 (N_8425,N_8291,N_8222);
and U8426 (N_8426,N_8274,N_8269);
and U8427 (N_8427,N_8315,N_8246);
and U8428 (N_8428,N_8231,N_8207);
nor U8429 (N_8429,N_8291,N_8225);
nor U8430 (N_8430,N_8229,N_8215);
nand U8431 (N_8431,N_8172,N_8189);
nor U8432 (N_8432,N_8165,N_8238);
nor U8433 (N_8433,N_8282,N_8246);
xnor U8434 (N_8434,N_8307,N_8206);
nor U8435 (N_8435,N_8307,N_8243);
or U8436 (N_8436,N_8188,N_8293);
nor U8437 (N_8437,N_8169,N_8181);
nor U8438 (N_8438,N_8289,N_8217);
or U8439 (N_8439,N_8174,N_8306);
and U8440 (N_8440,N_8192,N_8185);
nor U8441 (N_8441,N_8191,N_8238);
nand U8442 (N_8442,N_8191,N_8269);
and U8443 (N_8443,N_8178,N_8165);
xnor U8444 (N_8444,N_8242,N_8304);
or U8445 (N_8445,N_8307,N_8218);
nand U8446 (N_8446,N_8244,N_8225);
and U8447 (N_8447,N_8214,N_8234);
xnor U8448 (N_8448,N_8179,N_8246);
xor U8449 (N_8449,N_8181,N_8213);
or U8450 (N_8450,N_8232,N_8197);
nor U8451 (N_8451,N_8279,N_8294);
xnor U8452 (N_8452,N_8244,N_8245);
and U8453 (N_8453,N_8189,N_8250);
nor U8454 (N_8454,N_8188,N_8294);
nor U8455 (N_8455,N_8247,N_8276);
and U8456 (N_8456,N_8287,N_8235);
and U8457 (N_8457,N_8164,N_8245);
nand U8458 (N_8458,N_8289,N_8264);
nor U8459 (N_8459,N_8198,N_8319);
nor U8460 (N_8460,N_8251,N_8319);
or U8461 (N_8461,N_8211,N_8180);
nor U8462 (N_8462,N_8177,N_8293);
nand U8463 (N_8463,N_8245,N_8196);
xor U8464 (N_8464,N_8228,N_8305);
xor U8465 (N_8465,N_8167,N_8267);
xnor U8466 (N_8466,N_8169,N_8191);
or U8467 (N_8467,N_8229,N_8210);
xor U8468 (N_8468,N_8238,N_8234);
or U8469 (N_8469,N_8242,N_8204);
nor U8470 (N_8470,N_8245,N_8227);
or U8471 (N_8471,N_8191,N_8163);
and U8472 (N_8472,N_8189,N_8226);
xor U8473 (N_8473,N_8245,N_8310);
nor U8474 (N_8474,N_8313,N_8304);
nor U8475 (N_8475,N_8284,N_8219);
or U8476 (N_8476,N_8294,N_8170);
nand U8477 (N_8477,N_8198,N_8313);
and U8478 (N_8478,N_8170,N_8237);
or U8479 (N_8479,N_8219,N_8278);
nor U8480 (N_8480,N_8360,N_8358);
nand U8481 (N_8481,N_8343,N_8408);
nand U8482 (N_8482,N_8401,N_8476);
and U8483 (N_8483,N_8432,N_8330);
or U8484 (N_8484,N_8448,N_8454);
or U8485 (N_8485,N_8465,N_8374);
xnor U8486 (N_8486,N_8472,N_8362);
and U8487 (N_8487,N_8403,N_8364);
and U8488 (N_8488,N_8439,N_8413);
or U8489 (N_8489,N_8477,N_8386);
nor U8490 (N_8490,N_8450,N_8421);
or U8491 (N_8491,N_8412,N_8451);
and U8492 (N_8492,N_8449,N_8428);
and U8493 (N_8493,N_8361,N_8387);
nand U8494 (N_8494,N_8388,N_8347);
and U8495 (N_8495,N_8329,N_8372);
xor U8496 (N_8496,N_8411,N_8395);
nand U8497 (N_8497,N_8431,N_8427);
and U8498 (N_8498,N_8334,N_8475);
nand U8499 (N_8499,N_8442,N_8468);
nand U8500 (N_8500,N_8393,N_8389);
nand U8501 (N_8501,N_8379,N_8337);
nor U8502 (N_8502,N_8333,N_8325);
xnor U8503 (N_8503,N_8456,N_8383);
and U8504 (N_8504,N_8338,N_8416);
xnor U8505 (N_8505,N_8406,N_8396);
nor U8506 (N_8506,N_8459,N_8400);
and U8507 (N_8507,N_8366,N_8385);
nand U8508 (N_8508,N_8422,N_8430);
xnor U8509 (N_8509,N_8446,N_8352);
or U8510 (N_8510,N_8391,N_8326);
nor U8511 (N_8511,N_8417,N_8384);
xnor U8512 (N_8512,N_8353,N_8405);
xor U8513 (N_8513,N_8322,N_8356);
nor U8514 (N_8514,N_8328,N_8320);
and U8515 (N_8515,N_8373,N_8369);
or U8516 (N_8516,N_8368,N_8398);
and U8517 (N_8517,N_8340,N_8467);
or U8518 (N_8518,N_8321,N_8453);
nand U8519 (N_8519,N_8470,N_8447);
nor U8520 (N_8520,N_8350,N_8429);
and U8521 (N_8521,N_8363,N_8457);
nand U8522 (N_8522,N_8335,N_8354);
or U8523 (N_8523,N_8378,N_8415);
xnor U8524 (N_8524,N_8365,N_8377);
nor U8525 (N_8525,N_8332,N_8436);
nor U8526 (N_8526,N_8443,N_8473);
nor U8527 (N_8527,N_8357,N_8445);
nand U8528 (N_8528,N_8458,N_8380);
nor U8529 (N_8529,N_8419,N_8435);
nand U8530 (N_8530,N_8424,N_8370);
or U8531 (N_8531,N_8463,N_8423);
xnor U8532 (N_8532,N_8402,N_8323);
or U8533 (N_8533,N_8351,N_8336);
nor U8534 (N_8534,N_8414,N_8381);
nand U8535 (N_8535,N_8474,N_8461);
and U8536 (N_8536,N_8460,N_8425);
nor U8537 (N_8537,N_8437,N_8466);
nand U8538 (N_8538,N_8394,N_8342);
xor U8539 (N_8539,N_8444,N_8348);
nor U8540 (N_8540,N_8410,N_8355);
xnor U8541 (N_8541,N_8382,N_8464);
and U8542 (N_8542,N_8359,N_8438);
nor U8543 (N_8543,N_8349,N_8397);
xnor U8544 (N_8544,N_8478,N_8469);
or U8545 (N_8545,N_8471,N_8455);
nor U8546 (N_8546,N_8341,N_8399);
xor U8547 (N_8547,N_8392,N_8404);
and U8548 (N_8548,N_8371,N_8440);
nand U8549 (N_8549,N_8434,N_8367);
nand U8550 (N_8550,N_8433,N_8479);
nand U8551 (N_8551,N_8418,N_8462);
or U8552 (N_8552,N_8376,N_8409);
nor U8553 (N_8553,N_8345,N_8331);
and U8554 (N_8554,N_8346,N_8407);
nand U8555 (N_8555,N_8390,N_8324);
and U8556 (N_8556,N_8344,N_8420);
xnor U8557 (N_8557,N_8339,N_8327);
nand U8558 (N_8558,N_8441,N_8375);
nand U8559 (N_8559,N_8426,N_8452);
xnor U8560 (N_8560,N_8347,N_8396);
and U8561 (N_8561,N_8433,N_8336);
nor U8562 (N_8562,N_8447,N_8393);
nand U8563 (N_8563,N_8432,N_8420);
nand U8564 (N_8564,N_8459,N_8466);
nor U8565 (N_8565,N_8350,N_8451);
xor U8566 (N_8566,N_8399,N_8385);
xor U8567 (N_8567,N_8404,N_8446);
or U8568 (N_8568,N_8471,N_8472);
or U8569 (N_8569,N_8454,N_8376);
xnor U8570 (N_8570,N_8381,N_8379);
or U8571 (N_8571,N_8471,N_8426);
or U8572 (N_8572,N_8324,N_8456);
nor U8573 (N_8573,N_8378,N_8402);
and U8574 (N_8574,N_8431,N_8398);
nand U8575 (N_8575,N_8418,N_8345);
nand U8576 (N_8576,N_8361,N_8416);
and U8577 (N_8577,N_8344,N_8403);
xnor U8578 (N_8578,N_8427,N_8434);
or U8579 (N_8579,N_8371,N_8429);
or U8580 (N_8580,N_8464,N_8328);
and U8581 (N_8581,N_8420,N_8466);
nor U8582 (N_8582,N_8380,N_8468);
nor U8583 (N_8583,N_8387,N_8451);
and U8584 (N_8584,N_8321,N_8430);
nor U8585 (N_8585,N_8359,N_8477);
xor U8586 (N_8586,N_8321,N_8342);
nand U8587 (N_8587,N_8425,N_8331);
or U8588 (N_8588,N_8440,N_8460);
xnor U8589 (N_8589,N_8327,N_8362);
or U8590 (N_8590,N_8360,N_8474);
xnor U8591 (N_8591,N_8449,N_8377);
xnor U8592 (N_8592,N_8409,N_8415);
xor U8593 (N_8593,N_8363,N_8376);
nand U8594 (N_8594,N_8347,N_8389);
and U8595 (N_8595,N_8427,N_8403);
nor U8596 (N_8596,N_8329,N_8413);
and U8597 (N_8597,N_8385,N_8429);
or U8598 (N_8598,N_8348,N_8451);
or U8599 (N_8599,N_8390,N_8351);
and U8600 (N_8600,N_8376,N_8404);
or U8601 (N_8601,N_8445,N_8415);
xnor U8602 (N_8602,N_8419,N_8339);
xnor U8603 (N_8603,N_8351,N_8380);
xor U8604 (N_8604,N_8432,N_8320);
xnor U8605 (N_8605,N_8332,N_8406);
nor U8606 (N_8606,N_8451,N_8340);
nand U8607 (N_8607,N_8387,N_8450);
nand U8608 (N_8608,N_8419,N_8380);
xnor U8609 (N_8609,N_8390,N_8405);
or U8610 (N_8610,N_8407,N_8386);
or U8611 (N_8611,N_8369,N_8399);
nand U8612 (N_8612,N_8412,N_8380);
or U8613 (N_8613,N_8340,N_8394);
xnor U8614 (N_8614,N_8349,N_8378);
nand U8615 (N_8615,N_8441,N_8382);
nor U8616 (N_8616,N_8373,N_8477);
nand U8617 (N_8617,N_8447,N_8367);
and U8618 (N_8618,N_8414,N_8409);
and U8619 (N_8619,N_8404,N_8469);
xnor U8620 (N_8620,N_8457,N_8386);
nand U8621 (N_8621,N_8360,N_8424);
nor U8622 (N_8622,N_8384,N_8477);
and U8623 (N_8623,N_8415,N_8389);
nor U8624 (N_8624,N_8349,N_8433);
nand U8625 (N_8625,N_8411,N_8424);
or U8626 (N_8626,N_8367,N_8413);
or U8627 (N_8627,N_8472,N_8431);
and U8628 (N_8628,N_8389,N_8441);
nand U8629 (N_8629,N_8371,N_8478);
nand U8630 (N_8630,N_8468,N_8401);
nor U8631 (N_8631,N_8377,N_8350);
xnor U8632 (N_8632,N_8409,N_8386);
xor U8633 (N_8633,N_8410,N_8450);
nand U8634 (N_8634,N_8413,N_8405);
xnor U8635 (N_8635,N_8346,N_8357);
xnor U8636 (N_8636,N_8469,N_8343);
or U8637 (N_8637,N_8432,N_8449);
nor U8638 (N_8638,N_8454,N_8473);
or U8639 (N_8639,N_8429,N_8363);
nor U8640 (N_8640,N_8562,N_8543);
xor U8641 (N_8641,N_8531,N_8589);
nor U8642 (N_8642,N_8503,N_8547);
nor U8643 (N_8643,N_8594,N_8614);
nand U8644 (N_8644,N_8621,N_8525);
xor U8645 (N_8645,N_8528,N_8590);
nor U8646 (N_8646,N_8526,N_8540);
xnor U8647 (N_8647,N_8625,N_8495);
xnor U8648 (N_8648,N_8502,N_8609);
and U8649 (N_8649,N_8511,N_8581);
and U8650 (N_8650,N_8558,N_8494);
xnor U8651 (N_8651,N_8480,N_8600);
and U8652 (N_8652,N_8573,N_8607);
nand U8653 (N_8653,N_8497,N_8588);
nor U8654 (N_8654,N_8582,N_8535);
or U8655 (N_8655,N_8563,N_8623);
and U8656 (N_8656,N_8510,N_8541);
nand U8657 (N_8657,N_8513,N_8626);
nor U8658 (N_8658,N_8529,N_8604);
or U8659 (N_8659,N_8586,N_8548);
nor U8660 (N_8660,N_8555,N_8617);
or U8661 (N_8661,N_8556,N_8633);
nand U8662 (N_8662,N_8568,N_8501);
nand U8663 (N_8663,N_8591,N_8552);
nor U8664 (N_8664,N_8485,N_8632);
and U8665 (N_8665,N_8606,N_8585);
or U8666 (N_8666,N_8598,N_8489);
nor U8667 (N_8667,N_8553,N_8611);
nand U8668 (N_8668,N_8618,N_8629);
and U8669 (N_8669,N_8544,N_8539);
nand U8670 (N_8670,N_8508,N_8549);
nand U8671 (N_8671,N_8559,N_8596);
nor U8672 (N_8672,N_8515,N_8496);
nand U8673 (N_8673,N_8532,N_8577);
nor U8674 (N_8674,N_8487,N_8619);
nor U8675 (N_8675,N_8634,N_8512);
nand U8676 (N_8676,N_8639,N_8624);
nand U8677 (N_8677,N_8516,N_8514);
or U8678 (N_8678,N_8498,N_8627);
nand U8679 (N_8679,N_8550,N_8538);
xnor U8680 (N_8680,N_8576,N_8530);
or U8681 (N_8681,N_8564,N_8527);
nand U8682 (N_8682,N_8599,N_8488);
nand U8683 (N_8683,N_8481,N_8620);
nand U8684 (N_8684,N_8579,N_8580);
xor U8685 (N_8685,N_8493,N_8524);
nand U8686 (N_8686,N_8520,N_8631);
nand U8687 (N_8687,N_8638,N_8584);
nor U8688 (N_8688,N_8482,N_8536);
nor U8689 (N_8689,N_8551,N_8570);
and U8690 (N_8690,N_8509,N_8593);
nor U8691 (N_8691,N_8571,N_8505);
or U8692 (N_8692,N_8612,N_8546);
nand U8693 (N_8693,N_8613,N_8597);
nor U8694 (N_8694,N_8635,N_8557);
and U8695 (N_8695,N_8605,N_8572);
xor U8696 (N_8696,N_8484,N_8545);
xor U8697 (N_8697,N_8565,N_8575);
nand U8698 (N_8698,N_8587,N_8592);
or U8699 (N_8699,N_8630,N_8534);
nor U8700 (N_8700,N_8506,N_8523);
xor U8701 (N_8701,N_8637,N_8491);
and U8702 (N_8702,N_8628,N_8595);
nand U8703 (N_8703,N_8533,N_8492);
and U8704 (N_8704,N_8500,N_8507);
and U8705 (N_8705,N_8517,N_8560);
nand U8706 (N_8706,N_8522,N_8622);
nor U8707 (N_8707,N_8574,N_8537);
nand U8708 (N_8708,N_8567,N_8499);
xnor U8709 (N_8709,N_8601,N_8542);
nor U8710 (N_8710,N_8636,N_8608);
xnor U8711 (N_8711,N_8490,N_8519);
nor U8712 (N_8712,N_8483,N_8566);
and U8713 (N_8713,N_8504,N_8554);
nor U8714 (N_8714,N_8583,N_8578);
nand U8715 (N_8715,N_8486,N_8518);
nor U8716 (N_8716,N_8561,N_8610);
xnor U8717 (N_8717,N_8603,N_8521);
nor U8718 (N_8718,N_8615,N_8602);
and U8719 (N_8719,N_8569,N_8616);
nand U8720 (N_8720,N_8495,N_8534);
and U8721 (N_8721,N_8557,N_8582);
nor U8722 (N_8722,N_8561,N_8629);
nor U8723 (N_8723,N_8497,N_8609);
nor U8724 (N_8724,N_8529,N_8556);
or U8725 (N_8725,N_8570,N_8559);
nor U8726 (N_8726,N_8588,N_8548);
or U8727 (N_8727,N_8533,N_8521);
xnor U8728 (N_8728,N_8609,N_8577);
nor U8729 (N_8729,N_8624,N_8619);
xnor U8730 (N_8730,N_8532,N_8637);
xnor U8731 (N_8731,N_8614,N_8587);
and U8732 (N_8732,N_8519,N_8616);
or U8733 (N_8733,N_8534,N_8518);
and U8734 (N_8734,N_8636,N_8594);
nand U8735 (N_8735,N_8617,N_8488);
or U8736 (N_8736,N_8598,N_8515);
nor U8737 (N_8737,N_8609,N_8574);
nor U8738 (N_8738,N_8566,N_8556);
nand U8739 (N_8739,N_8529,N_8577);
nand U8740 (N_8740,N_8627,N_8572);
and U8741 (N_8741,N_8585,N_8580);
nor U8742 (N_8742,N_8501,N_8485);
or U8743 (N_8743,N_8598,N_8529);
nor U8744 (N_8744,N_8621,N_8519);
nor U8745 (N_8745,N_8623,N_8604);
xnor U8746 (N_8746,N_8494,N_8540);
and U8747 (N_8747,N_8482,N_8606);
nor U8748 (N_8748,N_8597,N_8587);
xnor U8749 (N_8749,N_8546,N_8541);
xor U8750 (N_8750,N_8482,N_8596);
nor U8751 (N_8751,N_8502,N_8509);
and U8752 (N_8752,N_8494,N_8603);
nor U8753 (N_8753,N_8549,N_8553);
xor U8754 (N_8754,N_8489,N_8604);
or U8755 (N_8755,N_8607,N_8588);
xor U8756 (N_8756,N_8523,N_8616);
nor U8757 (N_8757,N_8495,N_8493);
nor U8758 (N_8758,N_8595,N_8493);
nand U8759 (N_8759,N_8592,N_8483);
nand U8760 (N_8760,N_8610,N_8614);
nor U8761 (N_8761,N_8562,N_8502);
or U8762 (N_8762,N_8575,N_8619);
xor U8763 (N_8763,N_8624,N_8553);
xor U8764 (N_8764,N_8626,N_8531);
or U8765 (N_8765,N_8605,N_8528);
xnor U8766 (N_8766,N_8543,N_8547);
xnor U8767 (N_8767,N_8519,N_8558);
and U8768 (N_8768,N_8519,N_8557);
xor U8769 (N_8769,N_8583,N_8500);
or U8770 (N_8770,N_8615,N_8596);
nor U8771 (N_8771,N_8635,N_8547);
or U8772 (N_8772,N_8555,N_8610);
or U8773 (N_8773,N_8608,N_8512);
nand U8774 (N_8774,N_8513,N_8541);
or U8775 (N_8775,N_8608,N_8563);
xnor U8776 (N_8776,N_8515,N_8577);
xor U8777 (N_8777,N_8565,N_8604);
nor U8778 (N_8778,N_8551,N_8532);
or U8779 (N_8779,N_8518,N_8606);
nand U8780 (N_8780,N_8589,N_8506);
and U8781 (N_8781,N_8602,N_8512);
xnor U8782 (N_8782,N_8639,N_8591);
or U8783 (N_8783,N_8561,N_8537);
and U8784 (N_8784,N_8613,N_8496);
xor U8785 (N_8785,N_8615,N_8528);
nand U8786 (N_8786,N_8492,N_8616);
and U8787 (N_8787,N_8604,N_8504);
and U8788 (N_8788,N_8602,N_8481);
and U8789 (N_8789,N_8576,N_8515);
nand U8790 (N_8790,N_8598,N_8483);
and U8791 (N_8791,N_8591,N_8551);
nand U8792 (N_8792,N_8543,N_8496);
and U8793 (N_8793,N_8515,N_8520);
or U8794 (N_8794,N_8519,N_8586);
xnor U8795 (N_8795,N_8494,N_8505);
xnor U8796 (N_8796,N_8553,N_8595);
nor U8797 (N_8797,N_8525,N_8595);
nor U8798 (N_8798,N_8493,N_8548);
xor U8799 (N_8799,N_8531,N_8632);
and U8800 (N_8800,N_8783,N_8717);
nor U8801 (N_8801,N_8721,N_8715);
and U8802 (N_8802,N_8693,N_8722);
nand U8803 (N_8803,N_8656,N_8736);
nor U8804 (N_8804,N_8664,N_8667);
and U8805 (N_8805,N_8741,N_8742);
nor U8806 (N_8806,N_8697,N_8740);
or U8807 (N_8807,N_8671,N_8676);
or U8808 (N_8808,N_8642,N_8658);
nand U8809 (N_8809,N_8669,N_8773);
and U8810 (N_8810,N_8746,N_8756);
xnor U8811 (N_8811,N_8744,N_8644);
nor U8812 (N_8812,N_8657,N_8668);
xor U8813 (N_8813,N_8731,N_8729);
or U8814 (N_8814,N_8753,N_8739);
and U8815 (N_8815,N_8789,N_8705);
nand U8816 (N_8816,N_8788,N_8701);
nor U8817 (N_8817,N_8771,N_8776);
xnor U8818 (N_8818,N_8647,N_8772);
and U8819 (N_8819,N_8646,N_8686);
nand U8820 (N_8820,N_8790,N_8640);
nor U8821 (N_8821,N_8681,N_8648);
or U8822 (N_8822,N_8711,N_8723);
or U8823 (N_8823,N_8700,N_8682);
nand U8824 (N_8824,N_8651,N_8779);
nor U8825 (N_8825,N_8679,N_8743);
xor U8826 (N_8826,N_8734,N_8794);
nand U8827 (N_8827,N_8785,N_8685);
or U8828 (N_8828,N_8735,N_8643);
nor U8829 (N_8829,N_8799,N_8662);
xnor U8830 (N_8830,N_8732,N_8653);
or U8831 (N_8831,N_8696,N_8798);
or U8832 (N_8832,N_8687,N_8708);
and U8833 (N_8833,N_8752,N_8792);
or U8834 (N_8834,N_8703,N_8720);
or U8835 (N_8835,N_8689,N_8751);
nor U8836 (N_8836,N_8672,N_8778);
xor U8837 (N_8837,N_8787,N_8795);
or U8838 (N_8838,N_8650,N_8791);
nand U8839 (N_8839,N_8652,N_8737);
and U8840 (N_8840,N_8678,N_8713);
xor U8841 (N_8841,N_8663,N_8692);
nand U8842 (N_8842,N_8674,N_8754);
nor U8843 (N_8843,N_8762,N_8680);
xnor U8844 (N_8844,N_8774,N_8641);
nand U8845 (N_8845,N_8649,N_8768);
or U8846 (N_8846,N_8780,N_8777);
or U8847 (N_8847,N_8695,N_8767);
and U8848 (N_8848,N_8698,N_8738);
nor U8849 (N_8849,N_8770,N_8645);
nor U8850 (N_8850,N_8726,N_8784);
nor U8851 (N_8851,N_8745,N_8718);
nand U8852 (N_8852,N_8786,N_8728);
or U8853 (N_8853,N_8706,N_8699);
and U8854 (N_8854,N_8782,N_8796);
nor U8855 (N_8855,N_8691,N_8714);
nand U8856 (N_8856,N_8704,N_8763);
and U8857 (N_8857,N_8750,N_8707);
xnor U8858 (N_8858,N_8716,N_8766);
nor U8859 (N_8859,N_8690,N_8765);
or U8860 (N_8860,N_8659,N_8725);
and U8861 (N_8861,N_8665,N_8775);
xor U8862 (N_8862,N_8655,N_8709);
or U8863 (N_8863,N_8673,N_8702);
xor U8864 (N_8864,N_8666,N_8760);
nor U8865 (N_8865,N_8755,N_8683);
and U8866 (N_8866,N_8797,N_8661);
nand U8867 (N_8867,N_8660,N_8694);
nor U8868 (N_8868,N_8684,N_8710);
xnor U8869 (N_8869,N_8793,N_8688);
nor U8870 (N_8870,N_8677,N_8758);
and U8871 (N_8871,N_8724,N_8654);
xor U8872 (N_8872,N_8670,N_8761);
and U8873 (N_8873,N_8764,N_8712);
xor U8874 (N_8874,N_8730,N_8759);
nor U8875 (N_8875,N_8781,N_8675);
nor U8876 (N_8876,N_8769,N_8757);
nand U8877 (N_8877,N_8733,N_8749);
or U8878 (N_8878,N_8719,N_8747);
nand U8879 (N_8879,N_8727,N_8748);
xor U8880 (N_8880,N_8792,N_8789);
or U8881 (N_8881,N_8783,N_8735);
and U8882 (N_8882,N_8794,N_8705);
xnor U8883 (N_8883,N_8686,N_8707);
xor U8884 (N_8884,N_8792,N_8684);
nor U8885 (N_8885,N_8720,N_8661);
and U8886 (N_8886,N_8676,N_8759);
nand U8887 (N_8887,N_8663,N_8795);
xor U8888 (N_8888,N_8682,N_8784);
and U8889 (N_8889,N_8730,N_8762);
and U8890 (N_8890,N_8752,N_8723);
nand U8891 (N_8891,N_8771,N_8792);
or U8892 (N_8892,N_8765,N_8748);
or U8893 (N_8893,N_8659,N_8748);
or U8894 (N_8894,N_8677,N_8774);
and U8895 (N_8895,N_8654,N_8764);
xnor U8896 (N_8896,N_8731,N_8684);
and U8897 (N_8897,N_8661,N_8771);
xor U8898 (N_8898,N_8763,N_8692);
or U8899 (N_8899,N_8787,N_8793);
xor U8900 (N_8900,N_8663,N_8797);
xor U8901 (N_8901,N_8668,N_8661);
or U8902 (N_8902,N_8779,N_8727);
and U8903 (N_8903,N_8713,N_8662);
or U8904 (N_8904,N_8705,N_8755);
and U8905 (N_8905,N_8794,N_8733);
nand U8906 (N_8906,N_8692,N_8671);
or U8907 (N_8907,N_8665,N_8699);
and U8908 (N_8908,N_8711,N_8646);
and U8909 (N_8909,N_8782,N_8703);
nor U8910 (N_8910,N_8795,N_8652);
or U8911 (N_8911,N_8754,N_8717);
nand U8912 (N_8912,N_8786,N_8652);
xor U8913 (N_8913,N_8710,N_8667);
xor U8914 (N_8914,N_8755,N_8773);
xor U8915 (N_8915,N_8773,N_8718);
and U8916 (N_8916,N_8647,N_8715);
xnor U8917 (N_8917,N_8797,N_8788);
xor U8918 (N_8918,N_8798,N_8685);
xor U8919 (N_8919,N_8682,N_8725);
nand U8920 (N_8920,N_8713,N_8744);
or U8921 (N_8921,N_8767,N_8764);
and U8922 (N_8922,N_8761,N_8724);
xnor U8923 (N_8923,N_8678,N_8792);
or U8924 (N_8924,N_8754,N_8731);
nand U8925 (N_8925,N_8793,N_8712);
or U8926 (N_8926,N_8714,N_8668);
or U8927 (N_8927,N_8669,N_8651);
nor U8928 (N_8928,N_8677,N_8760);
xnor U8929 (N_8929,N_8732,N_8670);
nor U8930 (N_8930,N_8718,N_8721);
xor U8931 (N_8931,N_8708,N_8744);
or U8932 (N_8932,N_8695,N_8762);
nand U8933 (N_8933,N_8651,N_8799);
or U8934 (N_8934,N_8651,N_8745);
nand U8935 (N_8935,N_8751,N_8726);
nand U8936 (N_8936,N_8685,N_8711);
or U8937 (N_8937,N_8772,N_8753);
or U8938 (N_8938,N_8795,N_8699);
nand U8939 (N_8939,N_8725,N_8775);
or U8940 (N_8940,N_8703,N_8739);
nor U8941 (N_8941,N_8788,N_8727);
and U8942 (N_8942,N_8740,N_8686);
and U8943 (N_8943,N_8796,N_8645);
or U8944 (N_8944,N_8777,N_8691);
xnor U8945 (N_8945,N_8707,N_8780);
xor U8946 (N_8946,N_8701,N_8642);
and U8947 (N_8947,N_8778,N_8723);
and U8948 (N_8948,N_8674,N_8667);
or U8949 (N_8949,N_8656,N_8700);
and U8950 (N_8950,N_8707,N_8736);
xor U8951 (N_8951,N_8728,N_8675);
and U8952 (N_8952,N_8770,N_8663);
xor U8953 (N_8953,N_8701,N_8781);
nor U8954 (N_8954,N_8753,N_8664);
nand U8955 (N_8955,N_8702,N_8681);
xor U8956 (N_8956,N_8675,N_8697);
and U8957 (N_8957,N_8789,N_8759);
or U8958 (N_8958,N_8792,N_8769);
xnor U8959 (N_8959,N_8648,N_8767);
and U8960 (N_8960,N_8817,N_8922);
nor U8961 (N_8961,N_8928,N_8881);
or U8962 (N_8962,N_8816,N_8924);
nand U8963 (N_8963,N_8810,N_8906);
nand U8964 (N_8964,N_8857,N_8902);
nor U8965 (N_8965,N_8806,N_8892);
xnor U8966 (N_8966,N_8899,N_8813);
xnor U8967 (N_8967,N_8869,N_8855);
nand U8968 (N_8968,N_8845,N_8933);
or U8969 (N_8969,N_8829,N_8936);
or U8970 (N_8970,N_8894,N_8858);
xnor U8971 (N_8971,N_8887,N_8925);
nor U8972 (N_8972,N_8865,N_8826);
or U8973 (N_8973,N_8853,N_8907);
xor U8974 (N_8974,N_8909,N_8864);
nand U8975 (N_8975,N_8957,N_8875);
and U8976 (N_8976,N_8841,N_8884);
xnor U8977 (N_8977,N_8918,N_8898);
xor U8978 (N_8978,N_8901,N_8812);
and U8979 (N_8979,N_8867,N_8821);
or U8980 (N_8980,N_8904,N_8929);
or U8981 (N_8981,N_8866,N_8913);
nor U8982 (N_8982,N_8872,N_8800);
and U8983 (N_8983,N_8815,N_8863);
nand U8984 (N_8984,N_8886,N_8868);
and U8985 (N_8985,N_8830,N_8944);
nor U8986 (N_8986,N_8959,N_8940);
nor U8987 (N_8987,N_8951,N_8814);
or U8988 (N_8988,N_8860,N_8942);
nor U8989 (N_8989,N_8828,N_8953);
or U8990 (N_8990,N_8905,N_8958);
or U8991 (N_8991,N_8923,N_8948);
or U8992 (N_8992,N_8839,N_8874);
nand U8993 (N_8993,N_8859,N_8804);
nor U8994 (N_8994,N_8947,N_8949);
xnor U8995 (N_8995,N_8952,N_8896);
xor U8996 (N_8996,N_8917,N_8808);
xor U8997 (N_8997,N_8823,N_8803);
or U8998 (N_8998,N_8921,N_8811);
nor U8999 (N_8999,N_8908,N_8911);
nor U9000 (N_9000,N_8879,N_8843);
or U9001 (N_9001,N_8819,N_8895);
nand U9002 (N_9002,N_8851,N_8870);
nand U9003 (N_9003,N_8897,N_8846);
and U9004 (N_9004,N_8941,N_8801);
nand U9005 (N_9005,N_8877,N_8932);
nor U9006 (N_9006,N_8805,N_8945);
nand U9007 (N_9007,N_8890,N_8840);
nand U9008 (N_9008,N_8827,N_8834);
nand U9009 (N_9009,N_8883,N_8835);
nor U9010 (N_9010,N_8935,N_8893);
and U9011 (N_9011,N_8850,N_8842);
nand U9012 (N_9012,N_8856,N_8919);
and U9013 (N_9013,N_8861,N_8956);
and U9014 (N_9014,N_8854,N_8836);
xor U9015 (N_9015,N_8912,N_8888);
or U9016 (N_9016,N_8891,N_8809);
or U9017 (N_9017,N_8833,N_8954);
or U9018 (N_9018,N_8926,N_8910);
or U9019 (N_9019,N_8903,N_8914);
nand U9020 (N_9020,N_8915,N_8943);
xnor U9021 (N_9021,N_8950,N_8882);
nand U9022 (N_9022,N_8802,N_8832);
and U9023 (N_9023,N_8889,N_8820);
and U9024 (N_9024,N_8852,N_8927);
nand U9025 (N_9025,N_8876,N_8844);
xor U9026 (N_9026,N_8825,N_8838);
and U9027 (N_9027,N_8930,N_8939);
nand U9028 (N_9028,N_8831,N_8822);
and U9029 (N_9029,N_8862,N_8847);
nor U9030 (N_9030,N_8818,N_8878);
or U9031 (N_9031,N_8938,N_8934);
xor U9032 (N_9032,N_8873,N_8937);
and U9033 (N_9033,N_8946,N_8880);
or U9034 (N_9034,N_8849,N_8871);
or U9035 (N_9035,N_8916,N_8824);
nor U9036 (N_9036,N_8931,N_8848);
nand U9037 (N_9037,N_8955,N_8900);
nand U9038 (N_9038,N_8885,N_8837);
and U9039 (N_9039,N_8920,N_8807);
nor U9040 (N_9040,N_8872,N_8945);
xor U9041 (N_9041,N_8940,N_8840);
xnor U9042 (N_9042,N_8917,N_8854);
nand U9043 (N_9043,N_8870,N_8944);
or U9044 (N_9044,N_8891,N_8834);
or U9045 (N_9045,N_8843,N_8934);
and U9046 (N_9046,N_8831,N_8874);
nand U9047 (N_9047,N_8931,N_8882);
nand U9048 (N_9048,N_8887,N_8890);
nand U9049 (N_9049,N_8833,N_8819);
and U9050 (N_9050,N_8877,N_8948);
and U9051 (N_9051,N_8812,N_8949);
xnor U9052 (N_9052,N_8869,N_8840);
xnor U9053 (N_9053,N_8943,N_8929);
nand U9054 (N_9054,N_8958,N_8953);
and U9055 (N_9055,N_8915,N_8870);
xor U9056 (N_9056,N_8858,N_8907);
xnor U9057 (N_9057,N_8876,N_8943);
and U9058 (N_9058,N_8957,N_8918);
nor U9059 (N_9059,N_8936,N_8947);
or U9060 (N_9060,N_8947,N_8896);
and U9061 (N_9061,N_8821,N_8931);
nor U9062 (N_9062,N_8869,N_8892);
nor U9063 (N_9063,N_8900,N_8847);
nand U9064 (N_9064,N_8911,N_8830);
xnor U9065 (N_9065,N_8810,N_8823);
xor U9066 (N_9066,N_8905,N_8934);
or U9067 (N_9067,N_8959,N_8908);
nor U9068 (N_9068,N_8830,N_8879);
nor U9069 (N_9069,N_8837,N_8858);
nor U9070 (N_9070,N_8804,N_8866);
xor U9071 (N_9071,N_8950,N_8895);
or U9072 (N_9072,N_8878,N_8877);
or U9073 (N_9073,N_8950,N_8899);
or U9074 (N_9074,N_8876,N_8869);
nor U9075 (N_9075,N_8861,N_8901);
xnor U9076 (N_9076,N_8829,N_8848);
nand U9077 (N_9077,N_8821,N_8811);
or U9078 (N_9078,N_8845,N_8802);
or U9079 (N_9079,N_8852,N_8859);
nand U9080 (N_9080,N_8850,N_8948);
and U9081 (N_9081,N_8904,N_8933);
or U9082 (N_9082,N_8867,N_8909);
and U9083 (N_9083,N_8816,N_8913);
and U9084 (N_9084,N_8956,N_8824);
xnor U9085 (N_9085,N_8912,N_8812);
or U9086 (N_9086,N_8897,N_8841);
nor U9087 (N_9087,N_8914,N_8801);
and U9088 (N_9088,N_8898,N_8810);
or U9089 (N_9089,N_8908,N_8953);
nor U9090 (N_9090,N_8931,N_8914);
xor U9091 (N_9091,N_8845,N_8825);
nor U9092 (N_9092,N_8900,N_8925);
and U9093 (N_9093,N_8869,N_8810);
and U9094 (N_9094,N_8858,N_8926);
nand U9095 (N_9095,N_8870,N_8945);
or U9096 (N_9096,N_8821,N_8823);
nand U9097 (N_9097,N_8929,N_8867);
nand U9098 (N_9098,N_8897,N_8895);
nor U9099 (N_9099,N_8897,N_8809);
and U9100 (N_9100,N_8862,N_8819);
or U9101 (N_9101,N_8819,N_8942);
nand U9102 (N_9102,N_8951,N_8931);
xor U9103 (N_9103,N_8927,N_8933);
nor U9104 (N_9104,N_8848,N_8864);
and U9105 (N_9105,N_8905,N_8837);
nor U9106 (N_9106,N_8815,N_8836);
and U9107 (N_9107,N_8819,N_8866);
nor U9108 (N_9108,N_8894,N_8939);
nand U9109 (N_9109,N_8872,N_8885);
xor U9110 (N_9110,N_8833,N_8896);
nand U9111 (N_9111,N_8866,N_8850);
and U9112 (N_9112,N_8848,N_8807);
xnor U9113 (N_9113,N_8848,N_8946);
xnor U9114 (N_9114,N_8924,N_8903);
or U9115 (N_9115,N_8894,N_8838);
nor U9116 (N_9116,N_8857,N_8843);
nand U9117 (N_9117,N_8948,N_8900);
nand U9118 (N_9118,N_8948,N_8868);
nand U9119 (N_9119,N_8857,N_8809);
or U9120 (N_9120,N_9042,N_9004);
nor U9121 (N_9121,N_9009,N_9047);
or U9122 (N_9122,N_9039,N_9083);
and U9123 (N_9123,N_8975,N_9102);
or U9124 (N_9124,N_9029,N_9017);
nand U9125 (N_9125,N_9057,N_9091);
or U9126 (N_9126,N_9041,N_8977);
nor U9127 (N_9127,N_8991,N_9117);
and U9128 (N_9128,N_8980,N_8982);
xor U9129 (N_9129,N_9020,N_8993);
nor U9130 (N_9130,N_9115,N_8970);
nor U9131 (N_9131,N_9006,N_9081);
nand U9132 (N_9132,N_9074,N_9079);
nor U9133 (N_9133,N_9080,N_9109);
xnor U9134 (N_9134,N_9075,N_9108);
nor U9135 (N_9135,N_9067,N_9056);
and U9136 (N_9136,N_8983,N_9024);
or U9137 (N_9137,N_9048,N_9101);
nand U9138 (N_9138,N_9051,N_9107);
and U9139 (N_9139,N_9016,N_8986);
or U9140 (N_9140,N_8969,N_9070);
or U9141 (N_9141,N_9007,N_9104);
or U9142 (N_9142,N_9049,N_9045);
or U9143 (N_9143,N_9010,N_9071);
nor U9144 (N_9144,N_9046,N_8998);
nor U9145 (N_9145,N_9001,N_9060);
xor U9146 (N_9146,N_9072,N_9069);
nor U9147 (N_9147,N_9052,N_8979);
nand U9148 (N_9148,N_9105,N_8989);
nand U9149 (N_9149,N_8971,N_9002);
and U9150 (N_9150,N_9058,N_8963);
xor U9151 (N_9151,N_9003,N_9030);
or U9152 (N_9152,N_9095,N_9078);
nor U9153 (N_9153,N_9094,N_9027);
xnor U9154 (N_9154,N_8995,N_9014);
nor U9155 (N_9155,N_9037,N_9062);
nor U9156 (N_9156,N_8987,N_9077);
or U9157 (N_9157,N_9053,N_9100);
nor U9158 (N_9158,N_9096,N_9011);
and U9159 (N_9159,N_9054,N_9015);
xnor U9160 (N_9160,N_9012,N_9000);
xor U9161 (N_9161,N_9119,N_8985);
and U9162 (N_9162,N_9092,N_9086);
nor U9163 (N_9163,N_8968,N_9018);
and U9164 (N_9164,N_9084,N_9065);
nor U9165 (N_9165,N_9050,N_8999);
nand U9166 (N_9166,N_9043,N_9111);
nor U9167 (N_9167,N_9040,N_9044);
or U9168 (N_9168,N_9021,N_8996);
xnor U9169 (N_9169,N_9035,N_9066);
nor U9170 (N_9170,N_8966,N_9097);
xor U9171 (N_9171,N_9068,N_8992);
xor U9172 (N_9172,N_9114,N_8978);
nor U9173 (N_9173,N_9118,N_9090);
nand U9174 (N_9174,N_9088,N_8984);
or U9175 (N_9175,N_9098,N_9089);
or U9176 (N_9176,N_8964,N_9061);
nand U9177 (N_9177,N_8973,N_8997);
and U9178 (N_9178,N_8965,N_9038);
nor U9179 (N_9179,N_8988,N_9032);
xor U9180 (N_9180,N_9019,N_9023);
and U9181 (N_9181,N_9036,N_8962);
nor U9182 (N_9182,N_9063,N_9112);
nand U9183 (N_9183,N_9028,N_8976);
or U9184 (N_9184,N_9008,N_9005);
nand U9185 (N_9185,N_9110,N_9022);
xnor U9186 (N_9186,N_9106,N_8990);
or U9187 (N_9187,N_9034,N_9025);
and U9188 (N_9188,N_8981,N_8974);
or U9189 (N_9189,N_9055,N_8967);
xor U9190 (N_9190,N_9073,N_8994);
or U9191 (N_9191,N_8960,N_9033);
xor U9192 (N_9192,N_8972,N_9076);
nand U9193 (N_9193,N_8961,N_9093);
and U9194 (N_9194,N_9064,N_9082);
nand U9195 (N_9195,N_9059,N_9031);
nand U9196 (N_9196,N_9103,N_9013);
or U9197 (N_9197,N_9087,N_9085);
xnor U9198 (N_9198,N_9026,N_9113);
nor U9199 (N_9199,N_9099,N_9116);
xor U9200 (N_9200,N_9033,N_9027);
xor U9201 (N_9201,N_9030,N_9065);
or U9202 (N_9202,N_9042,N_9048);
xnor U9203 (N_9203,N_9087,N_9084);
xor U9204 (N_9204,N_9029,N_9044);
xor U9205 (N_9205,N_9033,N_9099);
nor U9206 (N_9206,N_8998,N_8984);
nor U9207 (N_9207,N_9111,N_8999);
nand U9208 (N_9208,N_9023,N_9064);
nand U9209 (N_9209,N_9104,N_9027);
nor U9210 (N_9210,N_8966,N_8975);
xor U9211 (N_9211,N_8980,N_9057);
nand U9212 (N_9212,N_9056,N_9049);
nor U9213 (N_9213,N_9036,N_8986);
nand U9214 (N_9214,N_9055,N_9029);
nand U9215 (N_9215,N_9108,N_9083);
xor U9216 (N_9216,N_9113,N_9023);
nor U9217 (N_9217,N_9071,N_8968);
nand U9218 (N_9218,N_9111,N_8987);
nor U9219 (N_9219,N_8988,N_9023);
nand U9220 (N_9220,N_8960,N_9091);
nand U9221 (N_9221,N_9114,N_9094);
or U9222 (N_9222,N_9050,N_9027);
nand U9223 (N_9223,N_9031,N_9002);
or U9224 (N_9224,N_9029,N_9028);
xor U9225 (N_9225,N_9076,N_9097);
and U9226 (N_9226,N_8993,N_9047);
nor U9227 (N_9227,N_8993,N_9015);
and U9228 (N_9228,N_9047,N_9118);
xnor U9229 (N_9229,N_8976,N_9107);
or U9230 (N_9230,N_9092,N_9006);
xor U9231 (N_9231,N_9050,N_9052);
or U9232 (N_9232,N_9075,N_9058);
xor U9233 (N_9233,N_9072,N_8989);
nand U9234 (N_9234,N_9113,N_8981);
or U9235 (N_9235,N_9065,N_9075);
xor U9236 (N_9236,N_9036,N_8983);
and U9237 (N_9237,N_9039,N_8983);
nand U9238 (N_9238,N_9020,N_8988);
nor U9239 (N_9239,N_8966,N_9070);
and U9240 (N_9240,N_8984,N_8977);
nand U9241 (N_9241,N_9083,N_9026);
and U9242 (N_9242,N_9098,N_9006);
xor U9243 (N_9243,N_9048,N_9110);
xnor U9244 (N_9244,N_9003,N_9004);
nand U9245 (N_9245,N_9095,N_8989);
and U9246 (N_9246,N_9062,N_9060);
nand U9247 (N_9247,N_8965,N_9095);
and U9248 (N_9248,N_9000,N_9074);
nand U9249 (N_9249,N_9066,N_9081);
nand U9250 (N_9250,N_9011,N_8971);
nand U9251 (N_9251,N_8979,N_8986);
nor U9252 (N_9252,N_9020,N_9096);
nand U9253 (N_9253,N_8974,N_9027);
and U9254 (N_9254,N_9009,N_9112);
nand U9255 (N_9255,N_9024,N_9071);
or U9256 (N_9256,N_9001,N_9112);
and U9257 (N_9257,N_9076,N_9082);
and U9258 (N_9258,N_9119,N_9085);
and U9259 (N_9259,N_9041,N_9047);
and U9260 (N_9260,N_8976,N_9003);
and U9261 (N_9261,N_8998,N_9007);
nor U9262 (N_9262,N_8977,N_8975);
and U9263 (N_9263,N_9059,N_8965);
and U9264 (N_9264,N_9075,N_9002);
or U9265 (N_9265,N_8985,N_9012);
xor U9266 (N_9266,N_8980,N_9062);
nand U9267 (N_9267,N_8966,N_8998);
xnor U9268 (N_9268,N_9074,N_9033);
or U9269 (N_9269,N_8990,N_8979);
or U9270 (N_9270,N_9109,N_9092);
nand U9271 (N_9271,N_8969,N_9083);
nor U9272 (N_9272,N_9085,N_8993);
or U9273 (N_9273,N_9096,N_8985);
xor U9274 (N_9274,N_9089,N_9035);
and U9275 (N_9275,N_8983,N_8973);
xor U9276 (N_9276,N_9041,N_8994);
nand U9277 (N_9277,N_9111,N_9030);
nand U9278 (N_9278,N_9032,N_9112);
nor U9279 (N_9279,N_8965,N_9047);
and U9280 (N_9280,N_9125,N_9200);
nand U9281 (N_9281,N_9203,N_9217);
xnor U9282 (N_9282,N_9173,N_9177);
xor U9283 (N_9283,N_9127,N_9252);
xnor U9284 (N_9284,N_9141,N_9261);
or U9285 (N_9285,N_9209,N_9153);
nor U9286 (N_9286,N_9249,N_9128);
xnor U9287 (N_9287,N_9198,N_9157);
nand U9288 (N_9288,N_9210,N_9253);
nor U9289 (N_9289,N_9175,N_9189);
nor U9290 (N_9290,N_9133,N_9241);
nand U9291 (N_9291,N_9220,N_9256);
or U9292 (N_9292,N_9235,N_9138);
xor U9293 (N_9293,N_9183,N_9123);
and U9294 (N_9294,N_9264,N_9242);
nand U9295 (N_9295,N_9196,N_9258);
nand U9296 (N_9296,N_9171,N_9159);
nand U9297 (N_9297,N_9169,N_9135);
nor U9298 (N_9298,N_9162,N_9254);
nand U9299 (N_9299,N_9181,N_9160);
and U9300 (N_9300,N_9168,N_9120);
nand U9301 (N_9301,N_9201,N_9166);
and U9302 (N_9302,N_9211,N_9260);
or U9303 (N_9303,N_9224,N_9272);
or U9304 (N_9304,N_9208,N_9202);
nor U9305 (N_9305,N_9223,N_9197);
or U9306 (N_9306,N_9247,N_9179);
nand U9307 (N_9307,N_9155,N_9279);
nor U9308 (N_9308,N_9273,N_9124);
and U9309 (N_9309,N_9184,N_9228);
and U9310 (N_9310,N_9246,N_9262);
and U9311 (N_9311,N_9182,N_9165);
nor U9312 (N_9312,N_9158,N_9143);
nand U9313 (N_9313,N_9271,N_9192);
or U9314 (N_9314,N_9234,N_9219);
xnor U9315 (N_9315,N_9164,N_9151);
nand U9316 (N_9316,N_9240,N_9222);
xnor U9317 (N_9317,N_9188,N_9195);
nand U9318 (N_9318,N_9191,N_9259);
nand U9319 (N_9319,N_9176,N_9238);
or U9320 (N_9320,N_9214,N_9140);
or U9321 (N_9321,N_9226,N_9145);
and U9322 (N_9322,N_9244,N_9190);
xnor U9323 (N_9323,N_9215,N_9237);
and U9324 (N_9324,N_9274,N_9265);
nand U9325 (N_9325,N_9199,N_9152);
or U9326 (N_9326,N_9144,N_9122);
xor U9327 (N_9327,N_9231,N_9239);
and U9328 (N_9328,N_9178,N_9174);
or U9329 (N_9329,N_9269,N_9263);
or U9330 (N_9330,N_9193,N_9180);
or U9331 (N_9331,N_9278,N_9221);
nand U9332 (N_9332,N_9205,N_9277);
xnor U9333 (N_9333,N_9185,N_9245);
nor U9334 (N_9334,N_9121,N_9150);
nor U9335 (N_9335,N_9147,N_9204);
nand U9336 (N_9336,N_9167,N_9227);
and U9337 (N_9337,N_9267,N_9156);
and U9338 (N_9338,N_9154,N_9139);
nand U9339 (N_9339,N_9213,N_9186);
nand U9340 (N_9340,N_9268,N_9229);
nand U9341 (N_9341,N_9194,N_9233);
or U9342 (N_9342,N_9212,N_9270);
xor U9343 (N_9343,N_9126,N_9170);
xor U9344 (N_9344,N_9149,N_9216);
or U9345 (N_9345,N_9148,N_9187);
or U9346 (N_9346,N_9257,N_9172);
xnor U9347 (N_9347,N_9206,N_9131);
nor U9348 (N_9348,N_9146,N_9243);
xor U9349 (N_9349,N_9132,N_9163);
and U9350 (N_9350,N_9230,N_9255);
xnor U9351 (N_9351,N_9275,N_9137);
xnor U9352 (N_9352,N_9276,N_9218);
nor U9353 (N_9353,N_9248,N_9250);
xor U9354 (N_9354,N_9136,N_9266);
nand U9355 (N_9355,N_9225,N_9232);
nand U9356 (N_9356,N_9207,N_9142);
nor U9357 (N_9357,N_9130,N_9161);
or U9358 (N_9358,N_9251,N_9134);
nand U9359 (N_9359,N_9129,N_9236);
xnor U9360 (N_9360,N_9259,N_9202);
nor U9361 (N_9361,N_9218,N_9211);
or U9362 (N_9362,N_9230,N_9172);
xnor U9363 (N_9363,N_9129,N_9155);
nor U9364 (N_9364,N_9142,N_9176);
nor U9365 (N_9365,N_9162,N_9175);
nand U9366 (N_9366,N_9131,N_9260);
nor U9367 (N_9367,N_9130,N_9205);
or U9368 (N_9368,N_9230,N_9180);
nor U9369 (N_9369,N_9194,N_9142);
or U9370 (N_9370,N_9191,N_9238);
or U9371 (N_9371,N_9249,N_9221);
or U9372 (N_9372,N_9267,N_9205);
nor U9373 (N_9373,N_9163,N_9170);
or U9374 (N_9374,N_9272,N_9255);
or U9375 (N_9375,N_9198,N_9258);
nor U9376 (N_9376,N_9184,N_9232);
xnor U9377 (N_9377,N_9231,N_9259);
nand U9378 (N_9378,N_9279,N_9243);
nor U9379 (N_9379,N_9188,N_9261);
nand U9380 (N_9380,N_9250,N_9277);
nor U9381 (N_9381,N_9137,N_9167);
nand U9382 (N_9382,N_9178,N_9158);
nand U9383 (N_9383,N_9134,N_9164);
or U9384 (N_9384,N_9248,N_9133);
nor U9385 (N_9385,N_9232,N_9141);
and U9386 (N_9386,N_9126,N_9187);
or U9387 (N_9387,N_9159,N_9194);
nand U9388 (N_9388,N_9175,N_9208);
and U9389 (N_9389,N_9167,N_9228);
xor U9390 (N_9390,N_9266,N_9172);
or U9391 (N_9391,N_9260,N_9152);
nor U9392 (N_9392,N_9245,N_9222);
xor U9393 (N_9393,N_9161,N_9177);
and U9394 (N_9394,N_9141,N_9263);
or U9395 (N_9395,N_9236,N_9189);
xor U9396 (N_9396,N_9187,N_9168);
nor U9397 (N_9397,N_9201,N_9134);
nand U9398 (N_9398,N_9200,N_9164);
or U9399 (N_9399,N_9175,N_9165);
nor U9400 (N_9400,N_9159,N_9213);
xor U9401 (N_9401,N_9213,N_9255);
and U9402 (N_9402,N_9147,N_9198);
xor U9403 (N_9403,N_9164,N_9191);
and U9404 (N_9404,N_9159,N_9158);
or U9405 (N_9405,N_9183,N_9273);
or U9406 (N_9406,N_9272,N_9200);
and U9407 (N_9407,N_9140,N_9272);
nor U9408 (N_9408,N_9220,N_9254);
or U9409 (N_9409,N_9160,N_9253);
nor U9410 (N_9410,N_9141,N_9237);
or U9411 (N_9411,N_9242,N_9150);
nand U9412 (N_9412,N_9232,N_9132);
and U9413 (N_9413,N_9153,N_9155);
or U9414 (N_9414,N_9122,N_9230);
nor U9415 (N_9415,N_9159,N_9140);
nand U9416 (N_9416,N_9223,N_9241);
nor U9417 (N_9417,N_9210,N_9172);
and U9418 (N_9418,N_9135,N_9261);
nand U9419 (N_9419,N_9191,N_9180);
or U9420 (N_9420,N_9253,N_9192);
nand U9421 (N_9421,N_9233,N_9235);
nand U9422 (N_9422,N_9254,N_9228);
nor U9423 (N_9423,N_9192,N_9153);
or U9424 (N_9424,N_9229,N_9187);
xnor U9425 (N_9425,N_9133,N_9161);
or U9426 (N_9426,N_9278,N_9167);
nor U9427 (N_9427,N_9222,N_9214);
and U9428 (N_9428,N_9254,N_9273);
xor U9429 (N_9429,N_9185,N_9217);
and U9430 (N_9430,N_9123,N_9269);
or U9431 (N_9431,N_9196,N_9187);
xnor U9432 (N_9432,N_9185,N_9122);
and U9433 (N_9433,N_9258,N_9125);
or U9434 (N_9434,N_9234,N_9209);
or U9435 (N_9435,N_9245,N_9272);
xnor U9436 (N_9436,N_9187,N_9207);
nand U9437 (N_9437,N_9267,N_9171);
nand U9438 (N_9438,N_9182,N_9192);
nand U9439 (N_9439,N_9183,N_9276);
nor U9440 (N_9440,N_9322,N_9405);
and U9441 (N_9441,N_9289,N_9365);
nor U9442 (N_9442,N_9417,N_9284);
nor U9443 (N_9443,N_9375,N_9280);
nor U9444 (N_9444,N_9385,N_9304);
nand U9445 (N_9445,N_9401,N_9368);
xnor U9446 (N_9446,N_9302,N_9306);
xor U9447 (N_9447,N_9395,N_9373);
xnor U9448 (N_9448,N_9419,N_9340);
nor U9449 (N_9449,N_9420,N_9319);
xnor U9450 (N_9450,N_9379,N_9351);
and U9451 (N_9451,N_9317,N_9394);
xnor U9452 (N_9452,N_9371,N_9335);
xor U9453 (N_9453,N_9424,N_9349);
or U9454 (N_9454,N_9303,N_9356);
or U9455 (N_9455,N_9337,N_9418);
or U9456 (N_9456,N_9377,N_9430);
xor U9457 (N_9457,N_9288,N_9406);
nand U9458 (N_9458,N_9363,N_9286);
and U9459 (N_9459,N_9438,N_9372);
nand U9460 (N_9460,N_9411,N_9345);
and U9461 (N_9461,N_9376,N_9325);
xor U9462 (N_9462,N_9310,N_9431);
and U9463 (N_9463,N_9374,N_9344);
nand U9464 (N_9464,N_9314,N_9383);
and U9465 (N_9465,N_9364,N_9397);
and U9466 (N_9466,N_9293,N_9329);
or U9467 (N_9467,N_9300,N_9318);
or U9468 (N_9468,N_9358,N_9414);
xnor U9469 (N_9469,N_9307,N_9410);
and U9470 (N_9470,N_9426,N_9336);
and U9471 (N_9471,N_9416,N_9433);
nor U9472 (N_9472,N_9295,N_9332);
and U9473 (N_9473,N_9381,N_9367);
and U9474 (N_9474,N_9309,N_9323);
xor U9475 (N_9475,N_9361,N_9382);
xnor U9476 (N_9476,N_9287,N_9330);
or U9477 (N_9477,N_9437,N_9353);
or U9478 (N_9478,N_9392,N_9281);
nand U9479 (N_9479,N_9359,N_9360);
xnor U9480 (N_9480,N_9386,N_9327);
nor U9481 (N_9481,N_9400,N_9393);
and U9482 (N_9482,N_9347,N_9290);
or U9483 (N_9483,N_9357,N_9296);
or U9484 (N_9484,N_9404,N_9331);
or U9485 (N_9485,N_9320,N_9352);
and U9486 (N_9486,N_9355,N_9333);
or U9487 (N_9487,N_9422,N_9312);
nor U9488 (N_9488,N_9412,N_9338);
or U9489 (N_9489,N_9316,N_9328);
xor U9490 (N_9490,N_9427,N_9348);
and U9491 (N_9491,N_9423,N_9370);
or U9492 (N_9492,N_9380,N_9409);
nand U9493 (N_9493,N_9402,N_9434);
nand U9494 (N_9494,N_9403,N_9384);
or U9495 (N_9495,N_9362,N_9390);
nor U9496 (N_9496,N_9439,N_9342);
nor U9497 (N_9497,N_9294,N_9339);
and U9498 (N_9498,N_9291,N_9387);
nor U9499 (N_9499,N_9301,N_9399);
xnor U9500 (N_9500,N_9396,N_9298);
or U9501 (N_9501,N_9292,N_9369);
or U9502 (N_9502,N_9428,N_9324);
xnor U9503 (N_9503,N_9408,N_9389);
nor U9504 (N_9504,N_9343,N_9297);
nor U9505 (N_9505,N_9315,N_9313);
and U9506 (N_9506,N_9366,N_9388);
nor U9507 (N_9507,N_9413,N_9326);
xor U9508 (N_9508,N_9398,N_9429);
and U9509 (N_9509,N_9283,N_9432);
nand U9510 (N_9510,N_9311,N_9282);
nand U9511 (N_9511,N_9334,N_9305);
nor U9512 (N_9512,N_9407,N_9299);
nor U9513 (N_9513,N_9346,N_9354);
nand U9514 (N_9514,N_9350,N_9378);
xor U9515 (N_9515,N_9421,N_9435);
xnor U9516 (N_9516,N_9436,N_9415);
and U9517 (N_9517,N_9425,N_9391);
or U9518 (N_9518,N_9341,N_9285);
and U9519 (N_9519,N_9321,N_9308);
or U9520 (N_9520,N_9405,N_9404);
or U9521 (N_9521,N_9392,N_9438);
or U9522 (N_9522,N_9330,N_9420);
nand U9523 (N_9523,N_9429,N_9318);
nand U9524 (N_9524,N_9341,N_9383);
xnor U9525 (N_9525,N_9328,N_9415);
nor U9526 (N_9526,N_9358,N_9361);
nand U9527 (N_9527,N_9429,N_9305);
or U9528 (N_9528,N_9346,N_9294);
nor U9529 (N_9529,N_9301,N_9319);
or U9530 (N_9530,N_9395,N_9286);
xnor U9531 (N_9531,N_9349,N_9405);
xor U9532 (N_9532,N_9318,N_9395);
nand U9533 (N_9533,N_9423,N_9296);
or U9534 (N_9534,N_9292,N_9433);
and U9535 (N_9535,N_9327,N_9387);
and U9536 (N_9536,N_9373,N_9418);
or U9537 (N_9537,N_9375,N_9417);
or U9538 (N_9538,N_9413,N_9349);
nand U9539 (N_9539,N_9393,N_9362);
nor U9540 (N_9540,N_9370,N_9425);
nand U9541 (N_9541,N_9428,N_9348);
and U9542 (N_9542,N_9330,N_9352);
and U9543 (N_9543,N_9384,N_9378);
xor U9544 (N_9544,N_9412,N_9411);
or U9545 (N_9545,N_9320,N_9365);
nand U9546 (N_9546,N_9308,N_9346);
or U9547 (N_9547,N_9430,N_9355);
or U9548 (N_9548,N_9381,N_9300);
xnor U9549 (N_9549,N_9378,N_9295);
and U9550 (N_9550,N_9412,N_9422);
xor U9551 (N_9551,N_9367,N_9351);
xnor U9552 (N_9552,N_9357,N_9406);
xor U9553 (N_9553,N_9350,N_9370);
nand U9554 (N_9554,N_9368,N_9318);
and U9555 (N_9555,N_9396,N_9343);
nand U9556 (N_9556,N_9345,N_9386);
xnor U9557 (N_9557,N_9286,N_9411);
and U9558 (N_9558,N_9309,N_9406);
xnor U9559 (N_9559,N_9390,N_9407);
and U9560 (N_9560,N_9297,N_9336);
nor U9561 (N_9561,N_9406,N_9334);
and U9562 (N_9562,N_9409,N_9431);
xnor U9563 (N_9563,N_9302,N_9403);
or U9564 (N_9564,N_9369,N_9332);
and U9565 (N_9565,N_9423,N_9368);
and U9566 (N_9566,N_9306,N_9364);
nand U9567 (N_9567,N_9306,N_9359);
and U9568 (N_9568,N_9358,N_9421);
and U9569 (N_9569,N_9358,N_9398);
nand U9570 (N_9570,N_9344,N_9323);
xor U9571 (N_9571,N_9400,N_9390);
nor U9572 (N_9572,N_9315,N_9337);
and U9573 (N_9573,N_9347,N_9395);
nor U9574 (N_9574,N_9390,N_9409);
xnor U9575 (N_9575,N_9373,N_9357);
xnor U9576 (N_9576,N_9374,N_9404);
xnor U9577 (N_9577,N_9367,N_9431);
and U9578 (N_9578,N_9295,N_9326);
xor U9579 (N_9579,N_9331,N_9430);
or U9580 (N_9580,N_9369,N_9398);
nor U9581 (N_9581,N_9389,N_9360);
nand U9582 (N_9582,N_9430,N_9406);
nand U9583 (N_9583,N_9410,N_9387);
xor U9584 (N_9584,N_9432,N_9287);
nor U9585 (N_9585,N_9334,N_9327);
nand U9586 (N_9586,N_9282,N_9393);
nand U9587 (N_9587,N_9367,N_9369);
and U9588 (N_9588,N_9330,N_9281);
and U9589 (N_9589,N_9327,N_9281);
nand U9590 (N_9590,N_9367,N_9340);
and U9591 (N_9591,N_9370,N_9320);
nand U9592 (N_9592,N_9342,N_9358);
nor U9593 (N_9593,N_9371,N_9379);
or U9594 (N_9594,N_9423,N_9373);
and U9595 (N_9595,N_9431,N_9293);
nand U9596 (N_9596,N_9438,N_9418);
nor U9597 (N_9597,N_9366,N_9303);
or U9598 (N_9598,N_9397,N_9305);
nand U9599 (N_9599,N_9361,N_9416);
nand U9600 (N_9600,N_9456,N_9583);
and U9601 (N_9601,N_9596,N_9577);
nor U9602 (N_9602,N_9522,N_9575);
xor U9603 (N_9603,N_9441,N_9538);
nor U9604 (N_9604,N_9526,N_9510);
or U9605 (N_9605,N_9449,N_9590);
nand U9606 (N_9606,N_9545,N_9592);
nor U9607 (N_9607,N_9565,N_9528);
or U9608 (N_9608,N_9547,N_9527);
nor U9609 (N_9609,N_9591,N_9554);
or U9610 (N_9610,N_9470,N_9549);
or U9611 (N_9611,N_9494,N_9579);
nand U9612 (N_9612,N_9541,N_9486);
nand U9613 (N_9613,N_9587,N_9542);
xnor U9614 (N_9614,N_9440,N_9462);
and U9615 (N_9615,N_9457,N_9524);
nand U9616 (N_9616,N_9557,N_9552);
nor U9617 (N_9617,N_9562,N_9567);
nor U9618 (N_9618,N_9515,N_9513);
nand U9619 (N_9619,N_9588,N_9523);
xor U9620 (N_9620,N_9502,N_9455);
nand U9621 (N_9621,N_9525,N_9478);
nand U9622 (N_9622,N_9546,N_9569);
nor U9623 (N_9623,N_9458,N_9492);
or U9624 (N_9624,N_9593,N_9580);
or U9625 (N_9625,N_9509,N_9466);
and U9626 (N_9626,N_9508,N_9564);
nand U9627 (N_9627,N_9558,N_9551);
xnor U9628 (N_9628,N_9481,N_9531);
and U9629 (N_9629,N_9533,N_9543);
or U9630 (N_9630,N_9582,N_9514);
xnor U9631 (N_9631,N_9489,N_9536);
and U9632 (N_9632,N_9594,N_9453);
and U9633 (N_9633,N_9573,N_9501);
xor U9634 (N_9634,N_9471,N_9459);
and U9635 (N_9635,N_9468,N_9472);
or U9636 (N_9636,N_9589,N_9556);
and U9637 (N_9637,N_9559,N_9535);
nand U9638 (N_9638,N_9530,N_9480);
and U9639 (N_9639,N_9448,N_9497);
or U9640 (N_9640,N_9443,N_9447);
nand U9641 (N_9641,N_9483,N_9519);
or U9642 (N_9642,N_9571,N_9445);
xnor U9643 (N_9643,N_9506,N_9585);
nand U9644 (N_9644,N_9487,N_9477);
or U9645 (N_9645,N_9532,N_9469);
nor U9646 (N_9646,N_9442,N_9544);
or U9647 (N_9647,N_9581,N_9467);
and U9648 (N_9648,N_9452,N_9463);
and U9649 (N_9649,N_9599,N_9490);
xor U9650 (N_9650,N_9495,N_9507);
nor U9651 (N_9651,N_9465,N_9518);
nand U9652 (N_9652,N_9566,N_9598);
xor U9653 (N_9653,N_9488,N_9568);
and U9654 (N_9654,N_9553,N_9493);
and U9655 (N_9655,N_9464,N_9548);
nand U9656 (N_9656,N_9516,N_9555);
nand U9657 (N_9657,N_9444,N_9496);
and U9658 (N_9658,N_9505,N_9451);
and U9659 (N_9659,N_9460,N_9504);
nor U9660 (N_9660,N_9540,N_9473);
xnor U9661 (N_9661,N_9500,N_9474);
xor U9662 (N_9662,N_9521,N_9482);
or U9663 (N_9663,N_9529,N_9550);
or U9664 (N_9664,N_9485,N_9476);
and U9665 (N_9665,N_9560,N_9484);
or U9666 (N_9666,N_9446,N_9517);
nand U9667 (N_9667,N_9586,N_9570);
xor U9668 (N_9668,N_9534,N_9454);
or U9669 (N_9669,N_9595,N_9574);
or U9670 (N_9670,N_9561,N_9537);
and U9671 (N_9671,N_9578,N_9563);
nor U9672 (N_9672,N_9475,N_9520);
nor U9673 (N_9673,N_9584,N_9498);
nor U9674 (N_9674,N_9479,N_9597);
nand U9675 (N_9675,N_9450,N_9461);
nand U9676 (N_9676,N_9499,N_9539);
nor U9677 (N_9677,N_9512,N_9511);
and U9678 (N_9678,N_9491,N_9576);
xor U9679 (N_9679,N_9503,N_9572);
nor U9680 (N_9680,N_9585,N_9469);
nand U9681 (N_9681,N_9452,N_9592);
xnor U9682 (N_9682,N_9530,N_9577);
nor U9683 (N_9683,N_9483,N_9531);
nand U9684 (N_9684,N_9460,N_9454);
or U9685 (N_9685,N_9574,N_9448);
or U9686 (N_9686,N_9441,N_9581);
nand U9687 (N_9687,N_9518,N_9578);
and U9688 (N_9688,N_9592,N_9558);
and U9689 (N_9689,N_9515,N_9552);
nor U9690 (N_9690,N_9459,N_9500);
and U9691 (N_9691,N_9571,N_9575);
nand U9692 (N_9692,N_9447,N_9595);
nor U9693 (N_9693,N_9532,N_9561);
xor U9694 (N_9694,N_9491,N_9503);
nand U9695 (N_9695,N_9492,N_9550);
nor U9696 (N_9696,N_9510,N_9540);
or U9697 (N_9697,N_9518,N_9511);
nor U9698 (N_9698,N_9547,N_9574);
xor U9699 (N_9699,N_9501,N_9448);
xnor U9700 (N_9700,N_9470,N_9505);
or U9701 (N_9701,N_9453,N_9529);
and U9702 (N_9702,N_9532,N_9484);
or U9703 (N_9703,N_9468,N_9574);
xnor U9704 (N_9704,N_9451,N_9469);
and U9705 (N_9705,N_9531,N_9576);
nand U9706 (N_9706,N_9548,N_9488);
and U9707 (N_9707,N_9553,N_9557);
nand U9708 (N_9708,N_9564,N_9579);
nor U9709 (N_9709,N_9457,N_9586);
nor U9710 (N_9710,N_9590,N_9551);
and U9711 (N_9711,N_9506,N_9517);
xnor U9712 (N_9712,N_9586,N_9541);
xor U9713 (N_9713,N_9455,N_9485);
xor U9714 (N_9714,N_9475,N_9594);
nand U9715 (N_9715,N_9564,N_9594);
nor U9716 (N_9716,N_9502,N_9477);
and U9717 (N_9717,N_9508,N_9544);
nor U9718 (N_9718,N_9529,N_9580);
nand U9719 (N_9719,N_9538,N_9468);
or U9720 (N_9720,N_9576,N_9537);
nand U9721 (N_9721,N_9457,N_9485);
and U9722 (N_9722,N_9519,N_9582);
and U9723 (N_9723,N_9531,N_9529);
and U9724 (N_9724,N_9497,N_9452);
nor U9725 (N_9725,N_9527,N_9541);
xor U9726 (N_9726,N_9443,N_9579);
nor U9727 (N_9727,N_9551,N_9515);
nand U9728 (N_9728,N_9533,N_9573);
and U9729 (N_9729,N_9446,N_9568);
nor U9730 (N_9730,N_9490,N_9555);
nand U9731 (N_9731,N_9583,N_9445);
and U9732 (N_9732,N_9550,N_9468);
or U9733 (N_9733,N_9590,N_9492);
or U9734 (N_9734,N_9537,N_9513);
and U9735 (N_9735,N_9488,N_9494);
nor U9736 (N_9736,N_9515,N_9534);
or U9737 (N_9737,N_9491,N_9465);
nor U9738 (N_9738,N_9578,N_9547);
or U9739 (N_9739,N_9569,N_9563);
nor U9740 (N_9740,N_9477,N_9534);
or U9741 (N_9741,N_9530,N_9551);
nand U9742 (N_9742,N_9569,N_9480);
or U9743 (N_9743,N_9578,N_9529);
nand U9744 (N_9744,N_9538,N_9461);
nand U9745 (N_9745,N_9474,N_9584);
or U9746 (N_9746,N_9575,N_9530);
xor U9747 (N_9747,N_9476,N_9539);
nor U9748 (N_9748,N_9447,N_9501);
nor U9749 (N_9749,N_9599,N_9509);
or U9750 (N_9750,N_9536,N_9573);
nor U9751 (N_9751,N_9583,N_9554);
nor U9752 (N_9752,N_9469,N_9453);
xnor U9753 (N_9753,N_9480,N_9490);
xor U9754 (N_9754,N_9544,N_9566);
or U9755 (N_9755,N_9572,N_9504);
or U9756 (N_9756,N_9468,N_9585);
or U9757 (N_9757,N_9444,N_9493);
and U9758 (N_9758,N_9477,N_9574);
or U9759 (N_9759,N_9522,N_9444);
or U9760 (N_9760,N_9616,N_9630);
and U9761 (N_9761,N_9612,N_9638);
and U9762 (N_9762,N_9665,N_9708);
or U9763 (N_9763,N_9656,N_9692);
nor U9764 (N_9764,N_9704,N_9695);
xnor U9765 (N_9765,N_9603,N_9647);
or U9766 (N_9766,N_9736,N_9660);
and U9767 (N_9767,N_9699,N_9719);
xnor U9768 (N_9768,N_9654,N_9730);
nand U9769 (N_9769,N_9661,N_9717);
xor U9770 (N_9770,N_9614,N_9711);
xor U9771 (N_9771,N_9663,N_9637);
nand U9772 (N_9772,N_9607,N_9731);
xnor U9773 (N_9773,N_9713,N_9696);
xor U9774 (N_9774,N_9685,N_9720);
nor U9775 (N_9775,N_9608,N_9678);
and U9776 (N_9776,N_9681,N_9675);
xnor U9777 (N_9777,N_9738,N_9600);
or U9778 (N_9778,N_9709,N_9657);
or U9779 (N_9779,N_9721,N_9702);
xnor U9780 (N_9780,N_9714,N_9621);
and U9781 (N_9781,N_9715,N_9739);
or U9782 (N_9782,N_9635,N_9673);
xor U9783 (N_9783,N_9634,N_9758);
nor U9784 (N_9784,N_9750,N_9606);
and U9785 (N_9785,N_9655,N_9674);
nor U9786 (N_9786,N_9601,N_9740);
xnor U9787 (N_9787,N_9633,N_9615);
nand U9788 (N_9788,N_9744,N_9602);
xnor U9789 (N_9789,N_9712,N_9753);
or U9790 (N_9790,N_9684,N_9722);
or U9791 (N_9791,N_9664,N_9718);
and U9792 (N_9792,N_9625,N_9624);
xor U9793 (N_9793,N_9705,N_9698);
or U9794 (N_9794,N_9703,N_9680);
nand U9795 (N_9795,N_9687,N_9748);
and U9796 (N_9796,N_9693,N_9682);
or U9797 (N_9797,N_9757,N_9737);
nand U9798 (N_9798,N_9746,N_9641);
nand U9799 (N_9799,N_9728,N_9623);
or U9800 (N_9800,N_9632,N_9651);
or U9801 (N_9801,N_9672,N_9686);
nor U9802 (N_9802,N_9611,N_9754);
or U9803 (N_9803,N_9690,N_9667);
xor U9804 (N_9804,N_9646,N_9751);
nand U9805 (N_9805,N_9752,N_9742);
nand U9806 (N_9806,N_9676,N_9658);
nand U9807 (N_9807,N_9735,N_9723);
xnor U9808 (N_9808,N_9645,N_9662);
xor U9809 (N_9809,N_9613,N_9636);
nand U9810 (N_9810,N_9609,N_9727);
or U9811 (N_9811,N_9644,N_9670);
nor U9812 (N_9812,N_9610,N_9683);
or U9813 (N_9813,N_9749,N_9741);
nand U9814 (N_9814,N_9648,N_9733);
xor U9815 (N_9815,N_9659,N_9724);
or U9816 (N_9816,N_9726,N_9707);
and U9817 (N_9817,N_9706,N_9631);
xnor U9818 (N_9818,N_9649,N_9747);
nand U9819 (N_9819,N_9669,N_9622);
nand U9820 (N_9820,N_9679,N_9643);
or U9821 (N_9821,N_9710,N_9701);
nor U9822 (N_9822,N_9650,N_9697);
nor U9823 (N_9823,N_9639,N_9640);
nor U9824 (N_9824,N_9604,N_9700);
or U9825 (N_9825,N_9732,N_9691);
and U9826 (N_9826,N_9677,N_9617);
and U9827 (N_9827,N_9618,N_9620);
nor U9828 (N_9828,N_9745,N_9629);
xnor U9829 (N_9829,N_9619,N_9668);
xnor U9830 (N_9830,N_9626,N_9605);
or U9831 (N_9831,N_9716,N_9689);
nand U9832 (N_9832,N_9666,N_9729);
nor U9833 (N_9833,N_9628,N_9756);
and U9834 (N_9834,N_9694,N_9688);
and U9835 (N_9835,N_9652,N_9642);
nor U9836 (N_9836,N_9743,N_9759);
or U9837 (N_9837,N_9755,N_9627);
xor U9838 (N_9838,N_9734,N_9725);
xnor U9839 (N_9839,N_9671,N_9653);
and U9840 (N_9840,N_9714,N_9600);
nand U9841 (N_9841,N_9654,N_9617);
nor U9842 (N_9842,N_9692,N_9629);
nand U9843 (N_9843,N_9696,N_9738);
or U9844 (N_9844,N_9747,N_9625);
and U9845 (N_9845,N_9709,N_9632);
nor U9846 (N_9846,N_9674,N_9611);
or U9847 (N_9847,N_9614,N_9608);
nand U9848 (N_9848,N_9704,N_9635);
xnor U9849 (N_9849,N_9657,N_9663);
xor U9850 (N_9850,N_9614,N_9759);
nor U9851 (N_9851,N_9713,N_9685);
nand U9852 (N_9852,N_9749,N_9639);
xor U9853 (N_9853,N_9658,N_9667);
and U9854 (N_9854,N_9610,N_9655);
xor U9855 (N_9855,N_9638,N_9699);
and U9856 (N_9856,N_9644,N_9685);
xor U9857 (N_9857,N_9696,N_9681);
nor U9858 (N_9858,N_9695,N_9630);
and U9859 (N_9859,N_9631,N_9708);
nor U9860 (N_9860,N_9695,N_9736);
nand U9861 (N_9861,N_9668,N_9697);
or U9862 (N_9862,N_9628,N_9739);
nand U9863 (N_9863,N_9755,N_9668);
nand U9864 (N_9864,N_9618,N_9657);
nor U9865 (N_9865,N_9672,N_9736);
nor U9866 (N_9866,N_9662,N_9727);
and U9867 (N_9867,N_9640,N_9631);
nand U9868 (N_9868,N_9745,N_9632);
nand U9869 (N_9869,N_9713,N_9622);
nand U9870 (N_9870,N_9642,N_9635);
or U9871 (N_9871,N_9680,N_9613);
nand U9872 (N_9872,N_9637,N_9610);
nand U9873 (N_9873,N_9698,N_9708);
xnor U9874 (N_9874,N_9719,N_9707);
xor U9875 (N_9875,N_9657,N_9632);
nor U9876 (N_9876,N_9624,N_9759);
xor U9877 (N_9877,N_9696,N_9638);
or U9878 (N_9878,N_9658,N_9612);
and U9879 (N_9879,N_9742,N_9719);
or U9880 (N_9880,N_9704,N_9698);
nand U9881 (N_9881,N_9659,N_9727);
xor U9882 (N_9882,N_9644,N_9743);
nor U9883 (N_9883,N_9689,N_9623);
xnor U9884 (N_9884,N_9682,N_9747);
nor U9885 (N_9885,N_9633,N_9668);
xnor U9886 (N_9886,N_9699,N_9600);
or U9887 (N_9887,N_9635,N_9613);
nor U9888 (N_9888,N_9710,N_9655);
or U9889 (N_9889,N_9636,N_9667);
nor U9890 (N_9890,N_9628,N_9718);
xor U9891 (N_9891,N_9743,N_9748);
or U9892 (N_9892,N_9741,N_9756);
nor U9893 (N_9893,N_9735,N_9676);
xor U9894 (N_9894,N_9657,N_9698);
or U9895 (N_9895,N_9610,N_9729);
xor U9896 (N_9896,N_9732,N_9730);
and U9897 (N_9897,N_9725,N_9747);
xor U9898 (N_9898,N_9615,N_9619);
or U9899 (N_9899,N_9736,N_9641);
and U9900 (N_9900,N_9621,N_9707);
nand U9901 (N_9901,N_9656,N_9733);
nand U9902 (N_9902,N_9726,N_9688);
and U9903 (N_9903,N_9615,N_9673);
nand U9904 (N_9904,N_9600,N_9657);
nor U9905 (N_9905,N_9657,N_9641);
xnor U9906 (N_9906,N_9720,N_9709);
or U9907 (N_9907,N_9624,N_9721);
and U9908 (N_9908,N_9711,N_9647);
or U9909 (N_9909,N_9631,N_9720);
or U9910 (N_9910,N_9698,N_9636);
nor U9911 (N_9911,N_9750,N_9658);
nand U9912 (N_9912,N_9620,N_9738);
or U9913 (N_9913,N_9607,N_9684);
nor U9914 (N_9914,N_9722,N_9609);
xnor U9915 (N_9915,N_9687,N_9647);
and U9916 (N_9916,N_9748,N_9659);
xnor U9917 (N_9917,N_9615,N_9654);
xor U9918 (N_9918,N_9635,N_9747);
nor U9919 (N_9919,N_9717,N_9677);
nor U9920 (N_9920,N_9806,N_9858);
or U9921 (N_9921,N_9821,N_9835);
or U9922 (N_9922,N_9765,N_9784);
nor U9923 (N_9923,N_9823,N_9890);
nand U9924 (N_9924,N_9868,N_9767);
and U9925 (N_9925,N_9844,N_9810);
and U9926 (N_9926,N_9853,N_9902);
nor U9927 (N_9927,N_9769,N_9917);
nand U9928 (N_9928,N_9781,N_9838);
and U9929 (N_9929,N_9881,N_9870);
xor U9930 (N_9930,N_9908,N_9856);
xnor U9931 (N_9931,N_9895,N_9860);
nor U9932 (N_9932,N_9776,N_9825);
and U9933 (N_9933,N_9845,N_9905);
or U9934 (N_9934,N_9787,N_9885);
or U9935 (N_9935,N_9774,N_9777);
nand U9936 (N_9936,N_9872,N_9826);
nor U9937 (N_9937,N_9848,N_9880);
xor U9938 (N_9938,N_9873,N_9813);
nand U9939 (N_9939,N_9915,N_9893);
and U9940 (N_9940,N_9795,N_9918);
xnor U9941 (N_9941,N_9883,N_9879);
nand U9942 (N_9942,N_9789,N_9830);
nand U9943 (N_9943,N_9862,N_9906);
or U9944 (N_9944,N_9778,N_9863);
nand U9945 (N_9945,N_9807,N_9779);
nor U9946 (N_9946,N_9907,N_9783);
and U9947 (N_9947,N_9865,N_9819);
nand U9948 (N_9948,N_9891,N_9843);
nand U9949 (N_9949,N_9909,N_9803);
nor U9950 (N_9950,N_9800,N_9761);
xor U9951 (N_9951,N_9898,N_9816);
or U9952 (N_9952,N_9916,N_9822);
nand U9953 (N_9953,N_9910,N_9874);
nor U9954 (N_9954,N_9846,N_9839);
nor U9955 (N_9955,N_9794,N_9801);
and U9956 (N_9956,N_9831,N_9798);
nor U9957 (N_9957,N_9892,N_9901);
nand U9958 (N_9958,N_9896,N_9833);
nand U9959 (N_9959,N_9887,N_9850);
and U9960 (N_9960,N_9799,N_9882);
xnor U9961 (N_9961,N_9809,N_9876);
and U9962 (N_9962,N_9857,N_9912);
and U9963 (N_9963,N_9802,N_9849);
and U9964 (N_9964,N_9842,N_9832);
nor U9965 (N_9965,N_9820,N_9837);
nand U9966 (N_9966,N_9897,N_9866);
nor U9967 (N_9967,N_9869,N_9836);
nand U9968 (N_9968,N_9796,N_9886);
and U9969 (N_9969,N_9797,N_9770);
or U9970 (N_9970,N_9847,N_9851);
xnor U9971 (N_9971,N_9815,N_9911);
nor U9972 (N_9972,N_9829,N_9864);
nand U9973 (N_9973,N_9824,N_9877);
nand U9974 (N_9974,N_9904,N_9760);
xor U9975 (N_9975,N_9808,N_9780);
xnor U9976 (N_9976,N_9817,N_9900);
or U9977 (N_9977,N_9859,N_9899);
or U9978 (N_9978,N_9827,N_9790);
and U9979 (N_9979,N_9884,N_9878);
xnor U9980 (N_9980,N_9788,N_9818);
nor U9981 (N_9981,N_9792,N_9762);
nand U9982 (N_9982,N_9773,N_9894);
or U9983 (N_9983,N_9841,N_9854);
or U9984 (N_9984,N_9867,N_9814);
and U9985 (N_9985,N_9775,N_9840);
and U9986 (N_9986,N_9914,N_9804);
and U9987 (N_9987,N_9768,N_9834);
xnor U9988 (N_9988,N_9903,N_9771);
or U9989 (N_9989,N_9828,N_9782);
nor U9990 (N_9990,N_9919,N_9811);
xnor U9991 (N_9991,N_9888,N_9889);
nor U9992 (N_9992,N_9855,N_9861);
xor U9993 (N_9993,N_9791,N_9913);
and U9994 (N_9994,N_9852,N_9805);
and U9995 (N_9995,N_9871,N_9766);
nor U9996 (N_9996,N_9772,N_9785);
and U9997 (N_9997,N_9812,N_9786);
xnor U9998 (N_9998,N_9764,N_9763);
xor U9999 (N_9999,N_9793,N_9875);
xor U10000 (N_10000,N_9885,N_9874);
nor U10001 (N_10001,N_9795,N_9821);
or U10002 (N_10002,N_9766,N_9913);
xor U10003 (N_10003,N_9868,N_9807);
and U10004 (N_10004,N_9838,N_9848);
nor U10005 (N_10005,N_9799,N_9762);
nand U10006 (N_10006,N_9801,N_9821);
and U10007 (N_10007,N_9877,N_9829);
or U10008 (N_10008,N_9828,N_9791);
nand U10009 (N_10009,N_9827,N_9825);
or U10010 (N_10010,N_9848,N_9915);
nand U10011 (N_10011,N_9851,N_9907);
nand U10012 (N_10012,N_9811,N_9851);
and U10013 (N_10013,N_9826,N_9828);
nand U10014 (N_10014,N_9837,N_9859);
and U10015 (N_10015,N_9902,N_9780);
xor U10016 (N_10016,N_9782,N_9842);
and U10017 (N_10017,N_9880,N_9876);
xor U10018 (N_10018,N_9797,N_9809);
nor U10019 (N_10019,N_9796,N_9871);
xnor U10020 (N_10020,N_9843,N_9815);
or U10021 (N_10021,N_9906,N_9857);
or U10022 (N_10022,N_9829,N_9868);
or U10023 (N_10023,N_9832,N_9806);
or U10024 (N_10024,N_9851,N_9862);
or U10025 (N_10025,N_9861,N_9856);
or U10026 (N_10026,N_9787,N_9763);
xor U10027 (N_10027,N_9832,N_9912);
and U10028 (N_10028,N_9777,N_9765);
nor U10029 (N_10029,N_9857,N_9877);
nor U10030 (N_10030,N_9911,N_9899);
nand U10031 (N_10031,N_9865,N_9908);
and U10032 (N_10032,N_9903,N_9906);
xnor U10033 (N_10033,N_9877,N_9900);
and U10034 (N_10034,N_9824,N_9768);
xnor U10035 (N_10035,N_9777,N_9776);
nand U10036 (N_10036,N_9863,N_9764);
xnor U10037 (N_10037,N_9796,N_9825);
nand U10038 (N_10038,N_9870,N_9772);
nor U10039 (N_10039,N_9839,N_9898);
and U10040 (N_10040,N_9768,N_9818);
xor U10041 (N_10041,N_9867,N_9908);
xor U10042 (N_10042,N_9845,N_9827);
nand U10043 (N_10043,N_9823,N_9812);
nand U10044 (N_10044,N_9876,N_9918);
nand U10045 (N_10045,N_9806,N_9822);
or U10046 (N_10046,N_9785,N_9856);
xor U10047 (N_10047,N_9781,N_9773);
nand U10048 (N_10048,N_9818,N_9766);
nand U10049 (N_10049,N_9896,N_9821);
nand U10050 (N_10050,N_9799,N_9893);
nand U10051 (N_10051,N_9919,N_9918);
or U10052 (N_10052,N_9878,N_9792);
and U10053 (N_10053,N_9875,N_9848);
nand U10054 (N_10054,N_9887,N_9818);
nor U10055 (N_10055,N_9863,N_9855);
nand U10056 (N_10056,N_9814,N_9839);
and U10057 (N_10057,N_9764,N_9868);
or U10058 (N_10058,N_9828,N_9769);
nor U10059 (N_10059,N_9919,N_9836);
nand U10060 (N_10060,N_9904,N_9889);
xor U10061 (N_10061,N_9815,N_9906);
nand U10062 (N_10062,N_9855,N_9828);
nand U10063 (N_10063,N_9784,N_9892);
nor U10064 (N_10064,N_9848,N_9784);
and U10065 (N_10065,N_9875,N_9796);
and U10066 (N_10066,N_9868,N_9904);
nor U10067 (N_10067,N_9853,N_9779);
nor U10068 (N_10068,N_9905,N_9805);
nor U10069 (N_10069,N_9828,N_9851);
and U10070 (N_10070,N_9818,N_9882);
xor U10071 (N_10071,N_9797,N_9804);
and U10072 (N_10072,N_9788,N_9857);
nor U10073 (N_10073,N_9889,N_9878);
and U10074 (N_10074,N_9786,N_9798);
xnor U10075 (N_10075,N_9789,N_9841);
xor U10076 (N_10076,N_9763,N_9872);
nand U10077 (N_10077,N_9876,N_9883);
or U10078 (N_10078,N_9854,N_9805);
or U10079 (N_10079,N_9907,N_9884);
or U10080 (N_10080,N_9957,N_10045);
nand U10081 (N_10081,N_9940,N_9967);
and U10082 (N_10082,N_10017,N_9982);
nand U10083 (N_10083,N_10000,N_9937);
nor U10084 (N_10084,N_10043,N_9976);
xnor U10085 (N_10085,N_10077,N_9991);
xor U10086 (N_10086,N_10065,N_9938);
nand U10087 (N_10087,N_9941,N_10008);
nor U10088 (N_10088,N_10032,N_9958);
nor U10089 (N_10089,N_9949,N_9960);
or U10090 (N_10090,N_9920,N_9954);
nand U10091 (N_10091,N_9948,N_10010);
nand U10092 (N_10092,N_9943,N_10067);
xnor U10093 (N_10093,N_9966,N_10029);
nand U10094 (N_10094,N_9961,N_10057);
nor U10095 (N_10095,N_10042,N_10049);
xnor U10096 (N_10096,N_10073,N_9980);
or U10097 (N_10097,N_10076,N_9995);
nor U10098 (N_10098,N_10040,N_9968);
or U10099 (N_10099,N_9933,N_9931);
nor U10100 (N_10100,N_10002,N_10005);
or U10101 (N_10101,N_10062,N_10051);
nor U10102 (N_10102,N_10035,N_10059);
xnor U10103 (N_10103,N_9977,N_10011);
nor U10104 (N_10104,N_9956,N_9946);
or U10105 (N_10105,N_10023,N_9984);
nand U10106 (N_10106,N_9923,N_9924);
and U10107 (N_10107,N_10009,N_9925);
and U10108 (N_10108,N_10014,N_10075);
xnor U10109 (N_10109,N_9998,N_10007);
nor U10110 (N_10110,N_10066,N_10046);
xnor U10111 (N_10111,N_10064,N_9971);
nor U10112 (N_10112,N_9993,N_10034);
xor U10113 (N_10113,N_9988,N_9947);
or U10114 (N_10114,N_9939,N_9985);
and U10115 (N_10115,N_10061,N_9996);
nand U10116 (N_10116,N_9962,N_10025);
nor U10117 (N_10117,N_9978,N_9932);
nand U10118 (N_10118,N_9944,N_10074);
nand U10119 (N_10119,N_10052,N_9928);
nor U10120 (N_10120,N_10050,N_9952);
nor U10121 (N_10121,N_10047,N_10036);
xor U10122 (N_10122,N_9992,N_9974);
nand U10123 (N_10123,N_9945,N_9972);
nand U10124 (N_10124,N_10015,N_10022);
xor U10125 (N_10125,N_10006,N_10033);
and U10126 (N_10126,N_10013,N_9986);
xnor U10127 (N_10127,N_10060,N_9951);
or U10128 (N_10128,N_10078,N_9989);
or U10129 (N_10129,N_9994,N_10021);
xnor U10130 (N_10130,N_9953,N_9929);
nor U10131 (N_10131,N_9927,N_9983);
and U10132 (N_10132,N_10038,N_10055);
or U10133 (N_10133,N_9921,N_10018);
xor U10134 (N_10134,N_9981,N_9970);
xor U10135 (N_10135,N_10027,N_10016);
xnor U10136 (N_10136,N_10012,N_9935);
nand U10137 (N_10137,N_10037,N_9964);
and U10138 (N_10138,N_10028,N_10069);
or U10139 (N_10139,N_9999,N_9963);
or U10140 (N_10140,N_10058,N_9973);
xor U10141 (N_10141,N_9934,N_10044);
or U10142 (N_10142,N_9936,N_10004);
nor U10143 (N_10143,N_10031,N_10079);
or U10144 (N_10144,N_9950,N_9955);
nor U10145 (N_10145,N_10048,N_10030);
xor U10146 (N_10146,N_9979,N_10003);
nand U10147 (N_10147,N_10054,N_10068);
nor U10148 (N_10148,N_10063,N_9997);
or U10149 (N_10149,N_10024,N_9965);
nor U10150 (N_10150,N_9987,N_9969);
and U10151 (N_10151,N_9990,N_10070);
nand U10152 (N_10152,N_9942,N_10041);
nand U10153 (N_10153,N_10026,N_9922);
and U10154 (N_10154,N_10056,N_10001);
xor U10155 (N_10155,N_10019,N_10053);
or U10156 (N_10156,N_10020,N_9930);
and U10157 (N_10157,N_9959,N_9926);
or U10158 (N_10158,N_10071,N_10072);
nor U10159 (N_10159,N_9975,N_10039);
nor U10160 (N_10160,N_10067,N_9983);
nor U10161 (N_10161,N_10071,N_10009);
nand U10162 (N_10162,N_10038,N_9968);
and U10163 (N_10163,N_10079,N_9994);
and U10164 (N_10164,N_10075,N_9995);
or U10165 (N_10165,N_9973,N_10015);
nor U10166 (N_10166,N_9930,N_9964);
nor U10167 (N_10167,N_9940,N_10049);
nor U10168 (N_10168,N_10029,N_10028);
nor U10169 (N_10169,N_10071,N_9953);
or U10170 (N_10170,N_10043,N_9967);
nor U10171 (N_10171,N_10052,N_9992);
nand U10172 (N_10172,N_10060,N_9969);
nand U10173 (N_10173,N_10022,N_9928);
nand U10174 (N_10174,N_10051,N_9950);
nor U10175 (N_10175,N_10038,N_10020);
or U10176 (N_10176,N_10015,N_10073);
and U10177 (N_10177,N_9966,N_9954);
nor U10178 (N_10178,N_9996,N_10008);
xor U10179 (N_10179,N_9998,N_10056);
xor U10180 (N_10180,N_9954,N_10007);
and U10181 (N_10181,N_9990,N_9936);
or U10182 (N_10182,N_10068,N_10043);
and U10183 (N_10183,N_10052,N_9968);
and U10184 (N_10184,N_10001,N_9966);
nand U10185 (N_10185,N_9996,N_10020);
xnor U10186 (N_10186,N_9948,N_9975);
xor U10187 (N_10187,N_10002,N_10038);
or U10188 (N_10188,N_9990,N_9964);
nand U10189 (N_10189,N_10004,N_10014);
nor U10190 (N_10190,N_10044,N_9946);
or U10191 (N_10191,N_10046,N_9973);
xnor U10192 (N_10192,N_9927,N_10020);
nor U10193 (N_10193,N_10067,N_9961);
and U10194 (N_10194,N_10058,N_9985);
xnor U10195 (N_10195,N_9983,N_9931);
and U10196 (N_10196,N_10003,N_10026);
nand U10197 (N_10197,N_9985,N_10013);
nor U10198 (N_10198,N_10044,N_9985);
or U10199 (N_10199,N_9939,N_10007);
nor U10200 (N_10200,N_10025,N_10002);
and U10201 (N_10201,N_9986,N_10027);
xnor U10202 (N_10202,N_10051,N_9941);
and U10203 (N_10203,N_10012,N_10010);
nand U10204 (N_10204,N_10020,N_10057);
xor U10205 (N_10205,N_9938,N_10004);
or U10206 (N_10206,N_9957,N_10030);
nand U10207 (N_10207,N_9958,N_9998);
and U10208 (N_10208,N_10052,N_9954);
xnor U10209 (N_10209,N_10027,N_9975);
and U10210 (N_10210,N_9999,N_9982);
nand U10211 (N_10211,N_10039,N_9980);
nor U10212 (N_10212,N_9925,N_9960);
nor U10213 (N_10213,N_9990,N_9920);
xor U10214 (N_10214,N_9933,N_9999);
and U10215 (N_10215,N_9936,N_9920);
xor U10216 (N_10216,N_10003,N_10029);
and U10217 (N_10217,N_10059,N_9997);
or U10218 (N_10218,N_9973,N_9993);
xor U10219 (N_10219,N_10000,N_10066);
and U10220 (N_10220,N_10008,N_9923);
nand U10221 (N_10221,N_9985,N_9965);
and U10222 (N_10222,N_10067,N_10015);
nor U10223 (N_10223,N_10039,N_9944);
nand U10224 (N_10224,N_10021,N_10016);
or U10225 (N_10225,N_10025,N_9999);
or U10226 (N_10226,N_9930,N_9947);
or U10227 (N_10227,N_10059,N_9936);
or U10228 (N_10228,N_9925,N_10024);
and U10229 (N_10229,N_9962,N_10043);
nand U10230 (N_10230,N_10027,N_9959);
nand U10231 (N_10231,N_9954,N_9975);
or U10232 (N_10232,N_10023,N_9978);
xnor U10233 (N_10233,N_10043,N_9995);
nor U10234 (N_10234,N_9951,N_9921);
nor U10235 (N_10235,N_10002,N_9942);
and U10236 (N_10236,N_10047,N_9943);
and U10237 (N_10237,N_9923,N_9954);
nor U10238 (N_10238,N_9980,N_10065);
xor U10239 (N_10239,N_9990,N_9925);
or U10240 (N_10240,N_10161,N_10203);
nand U10241 (N_10241,N_10129,N_10138);
and U10242 (N_10242,N_10159,N_10177);
or U10243 (N_10243,N_10124,N_10175);
xnor U10244 (N_10244,N_10090,N_10216);
xnor U10245 (N_10245,N_10081,N_10088);
nor U10246 (N_10246,N_10233,N_10231);
nand U10247 (N_10247,N_10179,N_10082);
xnor U10248 (N_10248,N_10100,N_10181);
nor U10249 (N_10249,N_10136,N_10080);
nand U10250 (N_10250,N_10191,N_10118);
xor U10251 (N_10251,N_10120,N_10164);
nand U10252 (N_10252,N_10105,N_10224);
nor U10253 (N_10253,N_10193,N_10152);
xnor U10254 (N_10254,N_10104,N_10102);
xor U10255 (N_10255,N_10218,N_10110);
xnor U10256 (N_10256,N_10239,N_10083);
and U10257 (N_10257,N_10204,N_10156);
and U10258 (N_10258,N_10207,N_10173);
xor U10259 (N_10259,N_10126,N_10232);
xnor U10260 (N_10260,N_10148,N_10225);
or U10261 (N_10261,N_10157,N_10205);
and U10262 (N_10262,N_10167,N_10116);
or U10263 (N_10263,N_10214,N_10108);
and U10264 (N_10264,N_10133,N_10095);
nand U10265 (N_10265,N_10230,N_10189);
xor U10266 (N_10266,N_10112,N_10234);
nand U10267 (N_10267,N_10132,N_10135);
xor U10268 (N_10268,N_10220,N_10211);
xor U10269 (N_10269,N_10227,N_10187);
and U10270 (N_10270,N_10163,N_10221);
nor U10271 (N_10271,N_10125,N_10178);
or U10272 (N_10272,N_10172,N_10155);
or U10273 (N_10273,N_10229,N_10144);
xor U10274 (N_10274,N_10085,N_10113);
xnor U10275 (N_10275,N_10131,N_10091);
and U10276 (N_10276,N_10117,N_10228);
nor U10277 (N_10277,N_10139,N_10168);
and U10278 (N_10278,N_10196,N_10141);
nor U10279 (N_10279,N_10162,N_10096);
and U10280 (N_10280,N_10174,N_10166);
nor U10281 (N_10281,N_10182,N_10160);
or U10282 (N_10282,N_10198,N_10123);
nor U10283 (N_10283,N_10119,N_10109);
or U10284 (N_10284,N_10171,N_10194);
nand U10285 (N_10285,N_10098,N_10183);
nand U10286 (N_10286,N_10208,N_10143);
or U10287 (N_10287,N_10145,N_10215);
xor U10288 (N_10288,N_10237,N_10190);
xor U10289 (N_10289,N_10169,N_10130);
and U10290 (N_10290,N_10217,N_10092);
or U10291 (N_10291,N_10128,N_10222);
nand U10292 (N_10292,N_10201,N_10127);
xnor U10293 (N_10293,N_10086,N_10101);
or U10294 (N_10294,N_10165,N_10195);
xnor U10295 (N_10295,N_10140,N_10223);
nor U10296 (N_10296,N_10235,N_10106);
and U10297 (N_10297,N_10122,N_10226);
or U10298 (N_10298,N_10137,N_10202);
xnor U10299 (N_10299,N_10115,N_10154);
nand U10300 (N_10300,N_10093,N_10121);
and U10301 (N_10301,N_10134,N_10153);
nor U10302 (N_10302,N_10111,N_10180);
or U10303 (N_10303,N_10114,N_10236);
and U10304 (N_10304,N_10199,N_10099);
nand U10305 (N_10305,N_10089,N_10185);
nor U10306 (N_10306,N_10097,N_10147);
or U10307 (N_10307,N_10192,N_10213);
xnor U10308 (N_10308,N_10158,N_10146);
xnor U10309 (N_10309,N_10087,N_10206);
xor U10310 (N_10310,N_10197,N_10219);
or U10311 (N_10311,N_10107,N_10150);
nor U10312 (N_10312,N_10200,N_10149);
xnor U10313 (N_10313,N_10238,N_10094);
nand U10314 (N_10314,N_10212,N_10176);
nor U10315 (N_10315,N_10151,N_10142);
or U10316 (N_10316,N_10188,N_10186);
and U10317 (N_10317,N_10103,N_10209);
nand U10318 (N_10318,N_10184,N_10170);
nor U10319 (N_10319,N_10210,N_10084);
and U10320 (N_10320,N_10212,N_10180);
nor U10321 (N_10321,N_10209,N_10085);
nand U10322 (N_10322,N_10226,N_10173);
nor U10323 (N_10323,N_10160,N_10188);
or U10324 (N_10324,N_10169,N_10111);
nand U10325 (N_10325,N_10168,N_10223);
nor U10326 (N_10326,N_10231,N_10202);
and U10327 (N_10327,N_10215,N_10182);
and U10328 (N_10328,N_10201,N_10119);
or U10329 (N_10329,N_10088,N_10156);
or U10330 (N_10330,N_10142,N_10099);
xnor U10331 (N_10331,N_10221,N_10205);
and U10332 (N_10332,N_10223,N_10164);
nor U10333 (N_10333,N_10140,N_10155);
nand U10334 (N_10334,N_10139,N_10101);
or U10335 (N_10335,N_10118,N_10096);
nor U10336 (N_10336,N_10192,N_10155);
and U10337 (N_10337,N_10234,N_10085);
nand U10338 (N_10338,N_10094,N_10188);
xor U10339 (N_10339,N_10104,N_10148);
and U10340 (N_10340,N_10134,N_10105);
and U10341 (N_10341,N_10149,N_10094);
or U10342 (N_10342,N_10221,N_10239);
nand U10343 (N_10343,N_10218,N_10176);
nand U10344 (N_10344,N_10191,N_10164);
nand U10345 (N_10345,N_10143,N_10183);
xnor U10346 (N_10346,N_10229,N_10131);
and U10347 (N_10347,N_10148,N_10187);
and U10348 (N_10348,N_10149,N_10099);
or U10349 (N_10349,N_10155,N_10179);
nand U10350 (N_10350,N_10221,N_10155);
nor U10351 (N_10351,N_10082,N_10141);
nor U10352 (N_10352,N_10222,N_10116);
nor U10353 (N_10353,N_10095,N_10149);
nand U10354 (N_10354,N_10204,N_10228);
nand U10355 (N_10355,N_10161,N_10134);
or U10356 (N_10356,N_10121,N_10116);
nor U10357 (N_10357,N_10135,N_10189);
nor U10358 (N_10358,N_10121,N_10106);
and U10359 (N_10359,N_10237,N_10125);
and U10360 (N_10360,N_10151,N_10088);
nand U10361 (N_10361,N_10203,N_10121);
nand U10362 (N_10362,N_10204,N_10210);
nand U10363 (N_10363,N_10147,N_10208);
xor U10364 (N_10364,N_10091,N_10121);
nand U10365 (N_10365,N_10120,N_10177);
nand U10366 (N_10366,N_10127,N_10216);
nand U10367 (N_10367,N_10188,N_10126);
and U10368 (N_10368,N_10161,N_10167);
and U10369 (N_10369,N_10120,N_10111);
or U10370 (N_10370,N_10184,N_10157);
and U10371 (N_10371,N_10224,N_10229);
and U10372 (N_10372,N_10203,N_10141);
and U10373 (N_10373,N_10173,N_10121);
nand U10374 (N_10374,N_10188,N_10147);
xor U10375 (N_10375,N_10115,N_10193);
and U10376 (N_10376,N_10177,N_10140);
and U10377 (N_10377,N_10185,N_10194);
and U10378 (N_10378,N_10156,N_10219);
nand U10379 (N_10379,N_10232,N_10237);
and U10380 (N_10380,N_10103,N_10084);
and U10381 (N_10381,N_10199,N_10168);
nor U10382 (N_10382,N_10206,N_10113);
xnor U10383 (N_10383,N_10117,N_10124);
and U10384 (N_10384,N_10237,N_10208);
or U10385 (N_10385,N_10119,N_10118);
xor U10386 (N_10386,N_10183,N_10089);
or U10387 (N_10387,N_10188,N_10088);
nand U10388 (N_10388,N_10081,N_10106);
nand U10389 (N_10389,N_10220,N_10199);
nand U10390 (N_10390,N_10093,N_10131);
xnor U10391 (N_10391,N_10088,N_10083);
nor U10392 (N_10392,N_10206,N_10144);
xor U10393 (N_10393,N_10108,N_10221);
and U10394 (N_10394,N_10147,N_10235);
nand U10395 (N_10395,N_10228,N_10088);
nor U10396 (N_10396,N_10219,N_10182);
xnor U10397 (N_10397,N_10126,N_10124);
xnor U10398 (N_10398,N_10154,N_10219);
and U10399 (N_10399,N_10204,N_10229);
nand U10400 (N_10400,N_10387,N_10318);
nor U10401 (N_10401,N_10345,N_10365);
nor U10402 (N_10402,N_10248,N_10357);
xnor U10403 (N_10403,N_10351,N_10290);
xor U10404 (N_10404,N_10257,N_10291);
nor U10405 (N_10405,N_10322,N_10298);
and U10406 (N_10406,N_10399,N_10320);
nor U10407 (N_10407,N_10358,N_10346);
and U10408 (N_10408,N_10374,N_10330);
nand U10409 (N_10409,N_10258,N_10262);
nand U10410 (N_10410,N_10370,N_10356);
nor U10411 (N_10411,N_10388,N_10244);
xnor U10412 (N_10412,N_10284,N_10323);
or U10413 (N_10413,N_10361,N_10375);
nand U10414 (N_10414,N_10255,N_10354);
xor U10415 (N_10415,N_10285,N_10302);
and U10416 (N_10416,N_10315,N_10347);
nor U10417 (N_10417,N_10334,N_10281);
and U10418 (N_10418,N_10329,N_10383);
xnor U10419 (N_10419,N_10277,N_10276);
and U10420 (N_10420,N_10381,N_10293);
or U10421 (N_10421,N_10327,N_10335);
nor U10422 (N_10422,N_10376,N_10336);
nand U10423 (N_10423,N_10397,N_10314);
and U10424 (N_10424,N_10270,N_10317);
nor U10425 (N_10425,N_10379,N_10288);
nand U10426 (N_10426,N_10274,N_10352);
nand U10427 (N_10427,N_10325,N_10266);
and U10428 (N_10428,N_10259,N_10303);
or U10429 (N_10429,N_10313,N_10287);
nor U10430 (N_10430,N_10342,N_10280);
or U10431 (N_10431,N_10344,N_10312);
and U10432 (N_10432,N_10349,N_10389);
nand U10433 (N_10433,N_10242,N_10273);
nand U10434 (N_10434,N_10307,N_10385);
or U10435 (N_10435,N_10260,N_10319);
or U10436 (N_10436,N_10264,N_10382);
and U10437 (N_10437,N_10377,N_10331);
and U10438 (N_10438,N_10240,N_10275);
and U10439 (N_10439,N_10250,N_10321);
or U10440 (N_10440,N_10295,N_10360);
and U10441 (N_10441,N_10338,N_10324);
nor U10442 (N_10442,N_10359,N_10343);
or U10443 (N_10443,N_10341,N_10305);
nor U10444 (N_10444,N_10328,N_10371);
or U10445 (N_10445,N_10333,N_10332);
or U10446 (N_10446,N_10363,N_10390);
xor U10447 (N_10447,N_10378,N_10380);
and U10448 (N_10448,N_10392,N_10367);
nand U10449 (N_10449,N_10391,N_10311);
or U10450 (N_10450,N_10394,N_10362);
nand U10451 (N_10451,N_10246,N_10369);
nand U10452 (N_10452,N_10304,N_10272);
and U10453 (N_10453,N_10241,N_10355);
nand U10454 (N_10454,N_10339,N_10310);
nand U10455 (N_10455,N_10300,N_10297);
nor U10456 (N_10456,N_10271,N_10373);
xnor U10457 (N_10457,N_10309,N_10251);
and U10458 (N_10458,N_10366,N_10350);
nand U10459 (N_10459,N_10348,N_10254);
xor U10460 (N_10460,N_10286,N_10252);
and U10461 (N_10461,N_10268,N_10279);
xor U10462 (N_10462,N_10294,N_10353);
xor U10463 (N_10463,N_10316,N_10278);
nand U10464 (N_10464,N_10249,N_10398);
xnor U10465 (N_10465,N_10253,N_10292);
and U10466 (N_10466,N_10364,N_10368);
and U10467 (N_10467,N_10372,N_10395);
or U10468 (N_10468,N_10261,N_10393);
or U10469 (N_10469,N_10243,N_10263);
and U10470 (N_10470,N_10308,N_10384);
nor U10471 (N_10471,N_10296,N_10265);
nand U10472 (N_10472,N_10282,N_10245);
nand U10473 (N_10473,N_10267,N_10337);
and U10474 (N_10474,N_10306,N_10326);
nor U10475 (N_10475,N_10396,N_10301);
nor U10476 (N_10476,N_10289,N_10340);
or U10477 (N_10477,N_10256,N_10269);
nor U10478 (N_10478,N_10283,N_10299);
xor U10479 (N_10479,N_10386,N_10247);
nor U10480 (N_10480,N_10301,N_10351);
or U10481 (N_10481,N_10271,N_10364);
and U10482 (N_10482,N_10250,N_10265);
xor U10483 (N_10483,N_10290,N_10268);
nor U10484 (N_10484,N_10363,N_10351);
nand U10485 (N_10485,N_10323,N_10381);
xor U10486 (N_10486,N_10312,N_10331);
xor U10487 (N_10487,N_10340,N_10305);
or U10488 (N_10488,N_10271,N_10298);
xnor U10489 (N_10489,N_10307,N_10347);
or U10490 (N_10490,N_10329,N_10259);
or U10491 (N_10491,N_10376,N_10360);
and U10492 (N_10492,N_10379,N_10364);
or U10493 (N_10493,N_10300,N_10358);
nor U10494 (N_10494,N_10368,N_10390);
and U10495 (N_10495,N_10297,N_10375);
and U10496 (N_10496,N_10293,N_10394);
nand U10497 (N_10497,N_10382,N_10245);
nand U10498 (N_10498,N_10276,N_10270);
nand U10499 (N_10499,N_10243,N_10318);
xnor U10500 (N_10500,N_10348,N_10310);
nand U10501 (N_10501,N_10272,N_10328);
or U10502 (N_10502,N_10319,N_10344);
xor U10503 (N_10503,N_10254,N_10363);
xor U10504 (N_10504,N_10292,N_10247);
xnor U10505 (N_10505,N_10244,N_10243);
and U10506 (N_10506,N_10342,N_10381);
or U10507 (N_10507,N_10377,N_10370);
xnor U10508 (N_10508,N_10353,N_10276);
nand U10509 (N_10509,N_10246,N_10372);
xnor U10510 (N_10510,N_10250,N_10394);
nand U10511 (N_10511,N_10388,N_10262);
nand U10512 (N_10512,N_10250,N_10393);
nor U10513 (N_10513,N_10362,N_10311);
nand U10514 (N_10514,N_10359,N_10399);
nor U10515 (N_10515,N_10389,N_10324);
xnor U10516 (N_10516,N_10243,N_10292);
or U10517 (N_10517,N_10275,N_10269);
and U10518 (N_10518,N_10263,N_10369);
and U10519 (N_10519,N_10399,N_10266);
xnor U10520 (N_10520,N_10324,N_10298);
and U10521 (N_10521,N_10358,N_10288);
nor U10522 (N_10522,N_10284,N_10382);
and U10523 (N_10523,N_10282,N_10260);
and U10524 (N_10524,N_10278,N_10277);
nor U10525 (N_10525,N_10294,N_10392);
nand U10526 (N_10526,N_10325,N_10350);
and U10527 (N_10527,N_10331,N_10346);
xnor U10528 (N_10528,N_10292,N_10312);
or U10529 (N_10529,N_10284,N_10290);
or U10530 (N_10530,N_10293,N_10335);
xor U10531 (N_10531,N_10279,N_10243);
and U10532 (N_10532,N_10264,N_10384);
xor U10533 (N_10533,N_10339,N_10306);
and U10534 (N_10534,N_10345,N_10342);
or U10535 (N_10535,N_10241,N_10286);
and U10536 (N_10536,N_10364,N_10352);
nand U10537 (N_10537,N_10365,N_10363);
nand U10538 (N_10538,N_10303,N_10328);
and U10539 (N_10539,N_10359,N_10249);
or U10540 (N_10540,N_10252,N_10270);
and U10541 (N_10541,N_10366,N_10275);
nand U10542 (N_10542,N_10359,N_10335);
xor U10543 (N_10543,N_10357,N_10306);
nand U10544 (N_10544,N_10339,N_10254);
and U10545 (N_10545,N_10367,N_10373);
xor U10546 (N_10546,N_10345,N_10302);
nor U10547 (N_10547,N_10261,N_10389);
nand U10548 (N_10548,N_10320,N_10263);
nor U10549 (N_10549,N_10263,N_10240);
nor U10550 (N_10550,N_10372,N_10282);
xor U10551 (N_10551,N_10278,N_10269);
nand U10552 (N_10552,N_10385,N_10315);
nand U10553 (N_10553,N_10360,N_10277);
or U10554 (N_10554,N_10308,N_10275);
and U10555 (N_10555,N_10302,N_10280);
nor U10556 (N_10556,N_10267,N_10327);
nand U10557 (N_10557,N_10261,N_10290);
and U10558 (N_10558,N_10317,N_10256);
xor U10559 (N_10559,N_10247,N_10333);
xnor U10560 (N_10560,N_10407,N_10473);
and U10561 (N_10561,N_10444,N_10455);
xor U10562 (N_10562,N_10467,N_10459);
nand U10563 (N_10563,N_10556,N_10442);
or U10564 (N_10564,N_10410,N_10424);
nand U10565 (N_10565,N_10477,N_10534);
nand U10566 (N_10566,N_10532,N_10509);
xnor U10567 (N_10567,N_10480,N_10557);
and U10568 (N_10568,N_10506,N_10525);
xnor U10569 (N_10569,N_10460,N_10402);
nor U10570 (N_10570,N_10436,N_10443);
nor U10571 (N_10571,N_10471,N_10415);
nand U10572 (N_10572,N_10423,N_10470);
or U10573 (N_10573,N_10517,N_10430);
nor U10574 (N_10574,N_10513,N_10466);
xnor U10575 (N_10575,N_10511,N_10457);
and U10576 (N_10576,N_10544,N_10403);
nand U10577 (N_10577,N_10540,N_10552);
nand U10578 (N_10578,N_10492,N_10405);
and U10579 (N_10579,N_10510,N_10411);
nor U10580 (N_10580,N_10418,N_10422);
and U10581 (N_10581,N_10536,N_10496);
xnor U10582 (N_10582,N_10531,N_10554);
nand U10583 (N_10583,N_10523,N_10401);
nor U10584 (N_10584,N_10538,N_10522);
nand U10585 (N_10585,N_10499,N_10553);
nor U10586 (N_10586,N_10468,N_10518);
nand U10587 (N_10587,N_10482,N_10551);
xnor U10588 (N_10588,N_10452,N_10539);
xnor U10589 (N_10589,N_10537,N_10484);
nand U10590 (N_10590,N_10400,N_10507);
nor U10591 (N_10591,N_10555,N_10475);
nand U10592 (N_10592,N_10488,N_10498);
nand U10593 (N_10593,N_10541,N_10426);
and U10594 (N_10594,N_10524,N_10514);
or U10595 (N_10595,N_10417,N_10446);
nand U10596 (N_10596,N_10515,N_10527);
nor U10597 (N_10597,N_10439,N_10487);
nand U10598 (N_10598,N_10420,N_10469);
nor U10599 (N_10599,N_10433,N_10429);
nor U10600 (N_10600,N_10500,N_10472);
nor U10601 (N_10601,N_10535,N_10558);
and U10602 (N_10602,N_10456,N_10427);
or U10603 (N_10603,N_10462,N_10516);
nor U10604 (N_10604,N_10497,N_10485);
nand U10605 (N_10605,N_10489,N_10440);
nand U10606 (N_10606,N_10445,N_10476);
xnor U10607 (N_10607,N_10463,N_10448);
nor U10608 (N_10608,N_10512,N_10451);
and U10609 (N_10609,N_10409,N_10533);
nand U10610 (N_10610,N_10449,N_10412);
nand U10611 (N_10611,N_10406,N_10493);
xnor U10612 (N_10612,N_10559,N_10437);
nor U10613 (N_10613,N_10431,N_10414);
nand U10614 (N_10614,N_10547,N_10545);
xnor U10615 (N_10615,N_10421,N_10491);
nand U10616 (N_10616,N_10546,N_10419);
and U10617 (N_10617,N_10425,N_10479);
or U10618 (N_10618,N_10501,N_10408);
and U10619 (N_10619,N_10526,N_10504);
xnor U10620 (N_10620,N_10495,N_10543);
and U10621 (N_10621,N_10478,N_10486);
nand U10622 (N_10622,N_10505,N_10416);
xnor U10623 (N_10623,N_10483,N_10454);
and U10624 (N_10624,N_10503,N_10494);
xor U10625 (N_10625,N_10465,N_10549);
and U10626 (N_10626,N_10413,N_10490);
and U10627 (N_10627,N_10404,N_10548);
or U10628 (N_10628,N_10508,N_10550);
nor U10629 (N_10629,N_10428,N_10502);
or U10630 (N_10630,N_10474,N_10529);
or U10631 (N_10631,N_10453,N_10521);
and U10632 (N_10632,N_10481,N_10542);
nand U10633 (N_10633,N_10438,N_10530);
nand U10634 (N_10634,N_10432,N_10435);
xor U10635 (N_10635,N_10519,N_10528);
or U10636 (N_10636,N_10520,N_10461);
nand U10637 (N_10637,N_10434,N_10441);
and U10638 (N_10638,N_10458,N_10450);
nor U10639 (N_10639,N_10447,N_10464);
nor U10640 (N_10640,N_10527,N_10476);
nand U10641 (N_10641,N_10536,N_10451);
or U10642 (N_10642,N_10431,N_10516);
nand U10643 (N_10643,N_10501,N_10499);
nand U10644 (N_10644,N_10468,N_10506);
and U10645 (N_10645,N_10408,N_10513);
and U10646 (N_10646,N_10549,N_10457);
nor U10647 (N_10647,N_10435,N_10444);
nor U10648 (N_10648,N_10411,N_10506);
or U10649 (N_10649,N_10515,N_10453);
and U10650 (N_10650,N_10478,N_10523);
xnor U10651 (N_10651,N_10462,N_10429);
xor U10652 (N_10652,N_10493,N_10485);
or U10653 (N_10653,N_10551,N_10400);
or U10654 (N_10654,N_10408,N_10412);
nand U10655 (N_10655,N_10528,N_10433);
nor U10656 (N_10656,N_10433,N_10450);
nor U10657 (N_10657,N_10405,N_10488);
xnor U10658 (N_10658,N_10523,N_10558);
or U10659 (N_10659,N_10405,N_10464);
xnor U10660 (N_10660,N_10403,N_10441);
and U10661 (N_10661,N_10460,N_10547);
nand U10662 (N_10662,N_10483,N_10476);
and U10663 (N_10663,N_10449,N_10411);
or U10664 (N_10664,N_10489,N_10421);
nand U10665 (N_10665,N_10526,N_10441);
nand U10666 (N_10666,N_10496,N_10524);
xnor U10667 (N_10667,N_10487,N_10520);
or U10668 (N_10668,N_10416,N_10457);
or U10669 (N_10669,N_10423,N_10434);
nand U10670 (N_10670,N_10530,N_10490);
and U10671 (N_10671,N_10542,N_10507);
nand U10672 (N_10672,N_10445,N_10441);
or U10673 (N_10673,N_10456,N_10511);
or U10674 (N_10674,N_10422,N_10521);
or U10675 (N_10675,N_10528,N_10466);
nand U10676 (N_10676,N_10554,N_10539);
nand U10677 (N_10677,N_10491,N_10552);
or U10678 (N_10678,N_10493,N_10461);
nor U10679 (N_10679,N_10522,N_10408);
nor U10680 (N_10680,N_10532,N_10521);
and U10681 (N_10681,N_10526,N_10501);
xor U10682 (N_10682,N_10405,N_10486);
or U10683 (N_10683,N_10419,N_10558);
nand U10684 (N_10684,N_10508,N_10528);
or U10685 (N_10685,N_10537,N_10505);
or U10686 (N_10686,N_10494,N_10541);
nor U10687 (N_10687,N_10487,N_10450);
and U10688 (N_10688,N_10432,N_10545);
xor U10689 (N_10689,N_10513,N_10551);
or U10690 (N_10690,N_10518,N_10411);
nand U10691 (N_10691,N_10534,N_10498);
nor U10692 (N_10692,N_10416,N_10490);
xor U10693 (N_10693,N_10546,N_10455);
and U10694 (N_10694,N_10468,N_10417);
or U10695 (N_10695,N_10519,N_10414);
xor U10696 (N_10696,N_10454,N_10492);
and U10697 (N_10697,N_10413,N_10500);
or U10698 (N_10698,N_10510,N_10527);
nor U10699 (N_10699,N_10482,N_10553);
or U10700 (N_10700,N_10408,N_10403);
or U10701 (N_10701,N_10514,N_10456);
xnor U10702 (N_10702,N_10502,N_10407);
and U10703 (N_10703,N_10508,N_10492);
nor U10704 (N_10704,N_10415,N_10552);
and U10705 (N_10705,N_10468,N_10512);
and U10706 (N_10706,N_10449,N_10432);
nand U10707 (N_10707,N_10466,N_10404);
or U10708 (N_10708,N_10437,N_10502);
nor U10709 (N_10709,N_10465,N_10539);
or U10710 (N_10710,N_10537,N_10503);
nand U10711 (N_10711,N_10417,N_10454);
xor U10712 (N_10712,N_10420,N_10412);
xnor U10713 (N_10713,N_10527,N_10442);
nor U10714 (N_10714,N_10473,N_10408);
nor U10715 (N_10715,N_10527,N_10447);
nor U10716 (N_10716,N_10492,N_10412);
nand U10717 (N_10717,N_10490,N_10447);
xor U10718 (N_10718,N_10444,N_10456);
xnor U10719 (N_10719,N_10544,N_10434);
nand U10720 (N_10720,N_10626,N_10645);
nand U10721 (N_10721,N_10687,N_10657);
xnor U10722 (N_10722,N_10624,N_10633);
nand U10723 (N_10723,N_10673,N_10702);
or U10724 (N_10724,N_10595,N_10677);
xnor U10725 (N_10725,N_10605,N_10713);
nand U10726 (N_10726,N_10719,N_10565);
or U10727 (N_10727,N_10576,N_10639);
nand U10728 (N_10728,N_10616,N_10563);
nor U10729 (N_10729,N_10609,N_10591);
nor U10730 (N_10730,N_10636,N_10588);
xor U10731 (N_10731,N_10665,N_10675);
and U10732 (N_10732,N_10668,N_10647);
and U10733 (N_10733,N_10715,N_10669);
xnor U10734 (N_10734,N_10688,N_10602);
nand U10735 (N_10735,N_10663,N_10598);
or U10736 (N_10736,N_10597,N_10603);
nor U10737 (N_10737,N_10651,N_10580);
nor U10738 (N_10738,N_10694,N_10573);
xor U10739 (N_10739,N_10672,N_10579);
or U10740 (N_10740,N_10604,N_10705);
nor U10741 (N_10741,N_10666,N_10637);
nor U10742 (N_10742,N_10708,N_10640);
nand U10743 (N_10743,N_10569,N_10601);
and U10744 (N_10744,N_10634,N_10593);
xor U10745 (N_10745,N_10681,N_10600);
nand U10746 (N_10746,N_10589,N_10700);
or U10747 (N_10747,N_10627,N_10667);
or U10748 (N_10748,N_10630,N_10623);
and U10749 (N_10749,N_10676,N_10693);
or U10750 (N_10750,N_10707,N_10586);
and U10751 (N_10751,N_10578,N_10615);
and U10752 (N_10752,N_10562,N_10661);
xor U10753 (N_10753,N_10712,N_10680);
xor U10754 (N_10754,N_10607,N_10568);
nand U10755 (N_10755,N_10585,N_10711);
or U10756 (N_10756,N_10574,N_10660);
and U10757 (N_10757,N_10691,N_10653);
nand U10758 (N_10758,N_10686,N_10618);
nand U10759 (N_10759,N_10575,N_10621);
or U10760 (N_10760,N_10583,N_10709);
nand U10761 (N_10761,N_10596,N_10678);
xnor U10762 (N_10762,N_10664,N_10570);
or U10763 (N_10763,N_10572,N_10577);
nand U10764 (N_10764,N_10679,N_10650);
nand U10765 (N_10765,N_10692,N_10701);
nand U10766 (N_10766,N_10685,N_10625);
nand U10767 (N_10767,N_10683,N_10646);
nand U10768 (N_10768,N_10614,N_10635);
and U10769 (N_10769,N_10581,N_10674);
nand U10770 (N_10770,N_10699,N_10710);
nor U10771 (N_10771,N_10622,N_10584);
or U10772 (N_10772,N_10695,N_10567);
and U10773 (N_10773,N_10696,N_10662);
nand U10774 (N_10774,N_10590,N_10611);
nand U10775 (N_10775,N_10631,N_10690);
nand U10776 (N_10776,N_10698,N_10587);
nand U10777 (N_10777,N_10717,N_10564);
nor U10778 (N_10778,N_10638,N_10689);
or U10779 (N_10779,N_10671,N_10617);
and U10780 (N_10780,N_10697,N_10682);
xnor U10781 (N_10781,N_10655,N_10610);
xnor U10782 (N_10782,N_10658,N_10608);
or U10783 (N_10783,N_10632,N_10670);
or U10784 (N_10784,N_10659,N_10654);
xor U10785 (N_10785,N_10703,N_10706);
nor U10786 (N_10786,N_10612,N_10652);
or U10787 (N_10787,N_10648,N_10716);
nor U10788 (N_10788,N_10620,N_10649);
or U10789 (N_10789,N_10641,N_10560);
xor U10790 (N_10790,N_10592,N_10594);
nand U10791 (N_10791,N_10644,N_10582);
nor U10792 (N_10792,N_10619,N_10561);
nor U10793 (N_10793,N_10718,N_10642);
nand U10794 (N_10794,N_10704,N_10566);
or U10795 (N_10795,N_10684,N_10656);
or U10796 (N_10796,N_10714,N_10629);
xor U10797 (N_10797,N_10606,N_10628);
nand U10798 (N_10798,N_10613,N_10571);
nand U10799 (N_10799,N_10643,N_10599);
and U10800 (N_10800,N_10586,N_10593);
and U10801 (N_10801,N_10580,N_10577);
nand U10802 (N_10802,N_10668,N_10695);
nand U10803 (N_10803,N_10620,N_10646);
xnor U10804 (N_10804,N_10621,N_10605);
nand U10805 (N_10805,N_10686,N_10571);
nand U10806 (N_10806,N_10714,N_10589);
xnor U10807 (N_10807,N_10605,N_10708);
nand U10808 (N_10808,N_10639,N_10682);
and U10809 (N_10809,N_10708,N_10658);
or U10810 (N_10810,N_10591,N_10632);
nand U10811 (N_10811,N_10564,N_10601);
and U10812 (N_10812,N_10687,N_10594);
nor U10813 (N_10813,N_10566,N_10620);
or U10814 (N_10814,N_10615,N_10691);
xnor U10815 (N_10815,N_10686,N_10636);
or U10816 (N_10816,N_10693,N_10625);
xor U10817 (N_10817,N_10589,N_10681);
nor U10818 (N_10818,N_10671,N_10619);
nor U10819 (N_10819,N_10719,N_10677);
xor U10820 (N_10820,N_10715,N_10652);
or U10821 (N_10821,N_10687,N_10605);
xor U10822 (N_10822,N_10625,N_10565);
nand U10823 (N_10823,N_10561,N_10704);
and U10824 (N_10824,N_10714,N_10562);
nor U10825 (N_10825,N_10668,N_10672);
and U10826 (N_10826,N_10715,N_10695);
and U10827 (N_10827,N_10688,N_10561);
nand U10828 (N_10828,N_10582,N_10705);
nor U10829 (N_10829,N_10664,N_10581);
or U10830 (N_10830,N_10718,N_10594);
or U10831 (N_10831,N_10707,N_10565);
xor U10832 (N_10832,N_10580,N_10643);
and U10833 (N_10833,N_10601,N_10719);
or U10834 (N_10834,N_10625,N_10649);
or U10835 (N_10835,N_10617,N_10677);
nand U10836 (N_10836,N_10710,N_10596);
and U10837 (N_10837,N_10691,N_10656);
nor U10838 (N_10838,N_10642,N_10681);
xnor U10839 (N_10839,N_10685,N_10697);
xnor U10840 (N_10840,N_10635,N_10600);
and U10841 (N_10841,N_10657,N_10640);
xnor U10842 (N_10842,N_10618,N_10715);
and U10843 (N_10843,N_10696,N_10712);
or U10844 (N_10844,N_10660,N_10652);
nand U10845 (N_10845,N_10669,N_10635);
and U10846 (N_10846,N_10684,N_10685);
or U10847 (N_10847,N_10572,N_10609);
nand U10848 (N_10848,N_10585,N_10651);
xor U10849 (N_10849,N_10609,N_10669);
nand U10850 (N_10850,N_10697,N_10574);
xnor U10851 (N_10851,N_10655,N_10628);
and U10852 (N_10852,N_10580,N_10574);
nor U10853 (N_10853,N_10633,N_10643);
and U10854 (N_10854,N_10596,N_10692);
nor U10855 (N_10855,N_10695,N_10656);
nand U10856 (N_10856,N_10659,N_10590);
or U10857 (N_10857,N_10703,N_10682);
xor U10858 (N_10858,N_10665,N_10623);
and U10859 (N_10859,N_10662,N_10625);
xor U10860 (N_10860,N_10670,N_10602);
nand U10861 (N_10861,N_10650,N_10609);
nand U10862 (N_10862,N_10665,N_10691);
nand U10863 (N_10863,N_10697,N_10670);
or U10864 (N_10864,N_10633,N_10578);
nor U10865 (N_10865,N_10716,N_10616);
nor U10866 (N_10866,N_10671,N_10664);
nor U10867 (N_10867,N_10578,N_10590);
xor U10868 (N_10868,N_10645,N_10617);
and U10869 (N_10869,N_10701,N_10574);
nor U10870 (N_10870,N_10607,N_10691);
nand U10871 (N_10871,N_10663,N_10679);
nand U10872 (N_10872,N_10608,N_10613);
nand U10873 (N_10873,N_10609,N_10585);
or U10874 (N_10874,N_10679,N_10651);
and U10875 (N_10875,N_10644,N_10664);
or U10876 (N_10876,N_10685,N_10629);
and U10877 (N_10877,N_10694,N_10675);
and U10878 (N_10878,N_10670,N_10668);
xnor U10879 (N_10879,N_10562,N_10627);
or U10880 (N_10880,N_10746,N_10765);
xor U10881 (N_10881,N_10806,N_10851);
xnor U10882 (N_10882,N_10727,N_10723);
or U10883 (N_10883,N_10733,N_10748);
or U10884 (N_10884,N_10737,N_10828);
nand U10885 (N_10885,N_10834,N_10730);
xor U10886 (N_10886,N_10790,N_10845);
nor U10887 (N_10887,N_10831,N_10796);
xor U10888 (N_10888,N_10773,N_10844);
nand U10889 (N_10889,N_10752,N_10755);
nand U10890 (N_10890,N_10780,N_10736);
or U10891 (N_10891,N_10801,N_10740);
and U10892 (N_10892,N_10819,N_10876);
nor U10893 (N_10893,N_10820,N_10782);
or U10894 (N_10894,N_10875,N_10829);
or U10895 (N_10895,N_10784,N_10843);
or U10896 (N_10896,N_10741,N_10821);
nand U10897 (N_10897,N_10735,N_10751);
and U10898 (N_10898,N_10877,N_10745);
or U10899 (N_10899,N_10814,N_10721);
and U10900 (N_10900,N_10857,N_10731);
and U10901 (N_10901,N_10793,N_10785);
nor U10902 (N_10902,N_10832,N_10766);
or U10903 (N_10903,N_10842,N_10783);
nor U10904 (N_10904,N_10817,N_10836);
and U10905 (N_10905,N_10826,N_10879);
nand U10906 (N_10906,N_10874,N_10769);
nand U10907 (N_10907,N_10799,N_10760);
nand U10908 (N_10908,N_10815,N_10781);
nand U10909 (N_10909,N_10865,N_10747);
xor U10910 (N_10910,N_10768,N_10792);
xor U10911 (N_10911,N_10763,N_10838);
xor U10912 (N_10912,N_10761,N_10724);
xnor U10913 (N_10913,N_10872,N_10795);
or U10914 (N_10914,N_10870,N_10802);
and U10915 (N_10915,N_10830,N_10762);
nand U10916 (N_10916,N_10774,N_10776);
or U10917 (N_10917,N_10812,N_10859);
nor U10918 (N_10918,N_10871,N_10854);
nor U10919 (N_10919,N_10850,N_10798);
xnor U10920 (N_10920,N_10811,N_10800);
or U10921 (N_10921,N_10777,N_10729);
xnor U10922 (N_10922,N_10726,N_10846);
or U10923 (N_10923,N_10804,N_10813);
nand U10924 (N_10924,N_10852,N_10770);
xnor U10925 (N_10925,N_10840,N_10861);
or U10926 (N_10926,N_10791,N_10873);
nand U10927 (N_10927,N_10771,N_10772);
and U10928 (N_10928,N_10858,N_10722);
nor U10929 (N_10929,N_10756,N_10786);
nand U10930 (N_10930,N_10767,N_10849);
xnor U10931 (N_10931,N_10827,N_10837);
nor U10932 (N_10932,N_10856,N_10808);
xor U10933 (N_10933,N_10810,N_10788);
nor U10934 (N_10934,N_10725,N_10853);
xnor U10935 (N_10935,N_10822,N_10742);
and U10936 (N_10936,N_10863,N_10744);
nand U10937 (N_10937,N_10758,N_10789);
nand U10938 (N_10938,N_10855,N_10732);
nor U10939 (N_10939,N_10720,N_10866);
xor U10940 (N_10940,N_10862,N_10809);
nor U10941 (N_10941,N_10841,N_10759);
and U10942 (N_10942,N_10816,N_10825);
or U10943 (N_10943,N_10867,N_10835);
nand U10944 (N_10944,N_10757,N_10860);
xor U10945 (N_10945,N_10794,N_10805);
and U10946 (N_10946,N_10864,N_10728);
or U10947 (N_10947,N_10847,N_10818);
nand U10948 (N_10948,N_10869,N_10807);
nor U10949 (N_10949,N_10787,N_10833);
nor U10950 (N_10950,N_10739,N_10848);
nand U10951 (N_10951,N_10749,N_10778);
and U10952 (N_10952,N_10868,N_10754);
xnor U10953 (N_10953,N_10839,N_10738);
nor U10954 (N_10954,N_10803,N_10775);
nand U10955 (N_10955,N_10823,N_10753);
xor U10956 (N_10956,N_10750,N_10764);
xor U10957 (N_10957,N_10824,N_10734);
and U10958 (N_10958,N_10797,N_10743);
and U10959 (N_10959,N_10878,N_10779);
and U10960 (N_10960,N_10758,N_10802);
nor U10961 (N_10961,N_10820,N_10836);
or U10962 (N_10962,N_10850,N_10826);
and U10963 (N_10963,N_10854,N_10804);
nor U10964 (N_10964,N_10838,N_10798);
nor U10965 (N_10965,N_10796,N_10737);
xnor U10966 (N_10966,N_10755,N_10753);
or U10967 (N_10967,N_10875,N_10848);
nand U10968 (N_10968,N_10747,N_10748);
xor U10969 (N_10969,N_10768,N_10830);
nor U10970 (N_10970,N_10778,N_10825);
or U10971 (N_10971,N_10788,N_10871);
nand U10972 (N_10972,N_10764,N_10836);
xnor U10973 (N_10973,N_10744,N_10729);
nand U10974 (N_10974,N_10724,N_10753);
xor U10975 (N_10975,N_10816,N_10851);
nor U10976 (N_10976,N_10735,N_10758);
nand U10977 (N_10977,N_10723,N_10776);
and U10978 (N_10978,N_10742,N_10834);
or U10979 (N_10979,N_10822,N_10776);
xnor U10980 (N_10980,N_10721,N_10769);
and U10981 (N_10981,N_10830,N_10834);
or U10982 (N_10982,N_10758,N_10820);
nand U10983 (N_10983,N_10830,N_10839);
nand U10984 (N_10984,N_10828,N_10731);
xor U10985 (N_10985,N_10758,N_10833);
or U10986 (N_10986,N_10858,N_10818);
xnor U10987 (N_10987,N_10801,N_10765);
xnor U10988 (N_10988,N_10765,N_10737);
and U10989 (N_10989,N_10790,N_10773);
nand U10990 (N_10990,N_10763,N_10795);
xor U10991 (N_10991,N_10812,N_10782);
nand U10992 (N_10992,N_10836,N_10731);
nand U10993 (N_10993,N_10753,N_10780);
and U10994 (N_10994,N_10775,N_10812);
xor U10995 (N_10995,N_10792,N_10824);
and U10996 (N_10996,N_10877,N_10842);
and U10997 (N_10997,N_10764,N_10841);
nor U10998 (N_10998,N_10785,N_10756);
nand U10999 (N_10999,N_10755,N_10858);
and U11000 (N_11000,N_10737,N_10797);
nor U11001 (N_11001,N_10753,N_10775);
nor U11002 (N_11002,N_10756,N_10738);
and U11003 (N_11003,N_10740,N_10815);
nand U11004 (N_11004,N_10875,N_10812);
nand U11005 (N_11005,N_10819,N_10738);
and U11006 (N_11006,N_10855,N_10783);
or U11007 (N_11007,N_10727,N_10869);
xor U11008 (N_11008,N_10725,N_10865);
and U11009 (N_11009,N_10792,N_10813);
xnor U11010 (N_11010,N_10871,N_10730);
nor U11011 (N_11011,N_10760,N_10740);
or U11012 (N_11012,N_10826,N_10818);
nor U11013 (N_11013,N_10721,N_10834);
xnor U11014 (N_11014,N_10770,N_10738);
and U11015 (N_11015,N_10722,N_10761);
nand U11016 (N_11016,N_10840,N_10747);
or U11017 (N_11017,N_10755,N_10870);
or U11018 (N_11018,N_10756,N_10859);
nand U11019 (N_11019,N_10752,N_10828);
or U11020 (N_11020,N_10871,N_10777);
and U11021 (N_11021,N_10841,N_10833);
nor U11022 (N_11022,N_10795,N_10779);
nand U11023 (N_11023,N_10866,N_10822);
and U11024 (N_11024,N_10731,N_10739);
or U11025 (N_11025,N_10852,N_10872);
or U11026 (N_11026,N_10773,N_10783);
and U11027 (N_11027,N_10795,N_10825);
xnor U11028 (N_11028,N_10739,N_10815);
xor U11029 (N_11029,N_10779,N_10818);
and U11030 (N_11030,N_10759,N_10737);
nand U11031 (N_11031,N_10856,N_10824);
or U11032 (N_11032,N_10876,N_10851);
nand U11033 (N_11033,N_10738,N_10816);
and U11034 (N_11034,N_10729,N_10796);
and U11035 (N_11035,N_10835,N_10770);
or U11036 (N_11036,N_10723,N_10810);
nand U11037 (N_11037,N_10735,N_10837);
nand U11038 (N_11038,N_10753,N_10838);
or U11039 (N_11039,N_10789,N_10740);
nand U11040 (N_11040,N_11039,N_10986);
nor U11041 (N_11041,N_10976,N_10983);
and U11042 (N_11042,N_10919,N_11006);
and U11043 (N_11043,N_10920,N_10972);
xor U11044 (N_11044,N_10934,N_10961);
nand U11045 (N_11045,N_10997,N_11012);
nor U11046 (N_11046,N_10977,N_10951);
xnor U11047 (N_11047,N_10954,N_10946);
or U11048 (N_11048,N_10894,N_11013);
nand U11049 (N_11049,N_10947,N_10962);
or U11050 (N_11050,N_10912,N_10999);
xor U11051 (N_11051,N_10922,N_11023);
nand U11052 (N_11052,N_10949,N_10939);
xor U11053 (N_11053,N_10896,N_10904);
and U11054 (N_11054,N_11036,N_10953);
nor U11055 (N_11055,N_10943,N_10930);
or U11056 (N_11056,N_10993,N_11015);
xor U11057 (N_11057,N_10979,N_10970);
or U11058 (N_11058,N_11030,N_11004);
nor U11059 (N_11059,N_10955,N_10906);
nand U11060 (N_11060,N_10917,N_11005);
xnor U11061 (N_11061,N_10909,N_10967);
nor U11062 (N_11062,N_10992,N_11033);
nand U11063 (N_11063,N_10888,N_10956);
nand U11064 (N_11064,N_11032,N_10968);
nand U11065 (N_11065,N_11018,N_10892);
xnor U11066 (N_11066,N_11034,N_10937);
nor U11067 (N_11067,N_11008,N_10925);
and U11068 (N_11068,N_11011,N_10938);
nand U11069 (N_11069,N_11035,N_10915);
and U11070 (N_11070,N_10959,N_10895);
nor U11071 (N_11071,N_11017,N_10964);
nor U11072 (N_11072,N_11037,N_10998);
xor U11073 (N_11073,N_11038,N_11024);
nor U11074 (N_11074,N_10990,N_10890);
nor U11075 (N_11075,N_10981,N_10884);
or U11076 (N_11076,N_10882,N_10980);
nor U11077 (N_11077,N_10881,N_11014);
nor U11078 (N_11078,N_11025,N_10901);
or U11079 (N_11079,N_10965,N_11022);
and U11080 (N_11080,N_10950,N_10978);
and U11081 (N_11081,N_10898,N_11019);
nor U11082 (N_11082,N_11016,N_11009);
nand U11083 (N_11083,N_11003,N_10933);
xor U11084 (N_11084,N_10916,N_10893);
nor U11085 (N_11085,N_10926,N_10987);
or U11086 (N_11086,N_10995,N_10982);
nand U11087 (N_11087,N_10929,N_11007);
or U11088 (N_11088,N_10908,N_10994);
nor U11089 (N_11089,N_10942,N_10897);
nand U11090 (N_11090,N_10910,N_10974);
and U11091 (N_11091,N_10928,N_10966);
xor U11092 (N_11092,N_10932,N_11021);
and U11093 (N_11093,N_11026,N_10945);
and U11094 (N_11094,N_11000,N_10958);
or U11095 (N_11095,N_11001,N_10944);
nand U11096 (N_11096,N_10921,N_10989);
and U11097 (N_11097,N_10940,N_11002);
xor U11098 (N_11098,N_10913,N_10960);
or U11099 (N_11099,N_10996,N_10885);
xor U11100 (N_11100,N_11031,N_10927);
or U11101 (N_11101,N_10911,N_10948);
nand U11102 (N_11102,N_10963,N_10936);
nand U11103 (N_11103,N_10952,N_10889);
or U11104 (N_11104,N_10887,N_10905);
and U11105 (N_11105,N_11029,N_10899);
nor U11106 (N_11106,N_10918,N_10886);
nor U11107 (N_11107,N_10984,N_11010);
and U11108 (N_11108,N_10891,N_10902);
nor U11109 (N_11109,N_10900,N_10969);
nor U11110 (N_11110,N_10880,N_10903);
nand U11111 (N_11111,N_10914,N_11027);
xor U11112 (N_11112,N_10991,N_10924);
xnor U11113 (N_11113,N_10957,N_10907);
and U11114 (N_11114,N_10931,N_10988);
nand U11115 (N_11115,N_10883,N_10923);
nand U11116 (N_11116,N_10985,N_10935);
or U11117 (N_11117,N_10941,N_10971);
xor U11118 (N_11118,N_11028,N_10973);
or U11119 (N_11119,N_11020,N_10975);
nand U11120 (N_11120,N_11036,N_10964);
xnor U11121 (N_11121,N_11026,N_10922);
or U11122 (N_11122,N_10881,N_11024);
nor U11123 (N_11123,N_10891,N_10885);
nand U11124 (N_11124,N_10921,N_10924);
nor U11125 (N_11125,N_10938,N_10906);
xnor U11126 (N_11126,N_11024,N_10963);
nor U11127 (N_11127,N_10941,N_10897);
or U11128 (N_11128,N_10957,N_10906);
or U11129 (N_11129,N_10901,N_10887);
xnor U11130 (N_11130,N_10975,N_11019);
xnor U11131 (N_11131,N_10959,N_11039);
nor U11132 (N_11132,N_10957,N_11017);
and U11133 (N_11133,N_10922,N_10891);
and U11134 (N_11134,N_11005,N_10892);
xnor U11135 (N_11135,N_10889,N_11010);
xnor U11136 (N_11136,N_11008,N_10887);
nand U11137 (N_11137,N_11036,N_11030);
nand U11138 (N_11138,N_10929,N_10972);
xnor U11139 (N_11139,N_11028,N_10895);
xnor U11140 (N_11140,N_10952,N_10986);
nor U11141 (N_11141,N_11015,N_11032);
nand U11142 (N_11142,N_10974,N_10905);
or U11143 (N_11143,N_10977,N_10962);
nor U11144 (N_11144,N_10881,N_10886);
nor U11145 (N_11145,N_11022,N_10915);
nor U11146 (N_11146,N_11033,N_10883);
and U11147 (N_11147,N_11030,N_11003);
xnor U11148 (N_11148,N_10931,N_10936);
or U11149 (N_11149,N_10964,N_10908);
nand U11150 (N_11150,N_10955,N_11020);
nor U11151 (N_11151,N_10971,N_10901);
and U11152 (N_11152,N_11039,N_10924);
and U11153 (N_11153,N_10911,N_11030);
nand U11154 (N_11154,N_10982,N_10975);
xnor U11155 (N_11155,N_10983,N_10909);
or U11156 (N_11156,N_11017,N_10951);
xnor U11157 (N_11157,N_10961,N_10937);
nand U11158 (N_11158,N_11022,N_10986);
nand U11159 (N_11159,N_10926,N_10920);
xor U11160 (N_11160,N_10886,N_10973);
and U11161 (N_11161,N_10981,N_10999);
or U11162 (N_11162,N_11020,N_11012);
xnor U11163 (N_11163,N_10915,N_10887);
xnor U11164 (N_11164,N_10895,N_10948);
nor U11165 (N_11165,N_10881,N_11002);
and U11166 (N_11166,N_10910,N_10941);
nand U11167 (N_11167,N_10932,N_10969);
or U11168 (N_11168,N_11019,N_10893);
xnor U11169 (N_11169,N_10932,N_10924);
xor U11170 (N_11170,N_10950,N_10895);
or U11171 (N_11171,N_11034,N_10997);
or U11172 (N_11172,N_10954,N_11036);
or U11173 (N_11173,N_10915,N_11028);
xnor U11174 (N_11174,N_11003,N_10906);
nand U11175 (N_11175,N_11007,N_10935);
nand U11176 (N_11176,N_10957,N_10890);
and U11177 (N_11177,N_10922,N_10974);
or U11178 (N_11178,N_10981,N_10917);
nand U11179 (N_11179,N_11038,N_10888);
nor U11180 (N_11180,N_10904,N_10969);
and U11181 (N_11181,N_10994,N_11002);
xor U11182 (N_11182,N_11008,N_10978);
nor U11183 (N_11183,N_11018,N_10981);
and U11184 (N_11184,N_10902,N_10911);
or U11185 (N_11185,N_10935,N_10979);
nor U11186 (N_11186,N_10949,N_10942);
and U11187 (N_11187,N_10904,N_10981);
nor U11188 (N_11188,N_10982,N_10933);
nor U11189 (N_11189,N_10979,N_10917);
or U11190 (N_11190,N_10950,N_11006);
or U11191 (N_11191,N_10892,N_10951);
nor U11192 (N_11192,N_11021,N_10916);
xor U11193 (N_11193,N_10904,N_10975);
xor U11194 (N_11194,N_11028,N_10997);
and U11195 (N_11195,N_10970,N_11008);
nor U11196 (N_11196,N_10993,N_11031);
nor U11197 (N_11197,N_10992,N_10964);
xor U11198 (N_11198,N_10994,N_11023);
and U11199 (N_11199,N_10907,N_10901);
and U11200 (N_11200,N_11048,N_11184);
xnor U11201 (N_11201,N_11138,N_11142);
nand U11202 (N_11202,N_11161,N_11108);
xnor U11203 (N_11203,N_11044,N_11090);
and U11204 (N_11204,N_11117,N_11118);
nand U11205 (N_11205,N_11174,N_11162);
nor U11206 (N_11206,N_11116,N_11065);
nand U11207 (N_11207,N_11169,N_11072);
and U11208 (N_11208,N_11140,N_11113);
nor U11209 (N_11209,N_11058,N_11144);
and U11210 (N_11210,N_11066,N_11198);
nor U11211 (N_11211,N_11163,N_11087);
and U11212 (N_11212,N_11127,N_11145);
or U11213 (N_11213,N_11130,N_11069);
and U11214 (N_11214,N_11085,N_11181);
and U11215 (N_11215,N_11155,N_11139);
and U11216 (N_11216,N_11153,N_11175);
or U11217 (N_11217,N_11125,N_11171);
xor U11218 (N_11218,N_11047,N_11056);
or U11219 (N_11219,N_11049,N_11149);
nor U11220 (N_11220,N_11061,N_11043);
nand U11221 (N_11221,N_11052,N_11192);
xor U11222 (N_11222,N_11167,N_11185);
xor U11223 (N_11223,N_11180,N_11176);
and U11224 (N_11224,N_11148,N_11107);
xor U11225 (N_11225,N_11099,N_11147);
and U11226 (N_11226,N_11096,N_11080);
xor U11227 (N_11227,N_11071,N_11088);
nand U11228 (N_11228,N_11098,N_11199);
xnor U11229 (N_11229,N_11103,N_11115);
and U11230 (N_11230,N_11154,N_11068);
nand U11231 (N_11231,N_11160,N_11150);
nand U11232 (N_11232,N_11134,N_11188);
and U11233 (N_11233,N_11093,N_11119);
nand U11234 (N_11234,N_11110,N_11050);
and U11235 (N_11235,N_11158,N_11053);
and U11236 (N_11236,N_11156,N_11121);
xnor U11237 (N_11237,N_11132,N_11194);
or U11238 (N_11238,N_11041,N_11124);
xor U11239 (N_11239,N_11126,N_11054);
xnor U11240 (N_11240,N_11191,N_11059);
xor U11241 (N_11241,N_11089,N_11091);
nand U11242 (N_11242,N_11081,N_11057);
and U11243 (N_11243,N_11045,N_11083);
and U11244 (N_11244,N_11106,N_11143);
nand U11245 (N_11245,N_11135,N_11094);
nand U11246 (N_11246,N_11128,N_11131);
or U11247 (N_11247,N_11101,N_11196);
xnor U11248 (N_11248,N_11120,N_11152);
or U11249 (N_11249,N_11170,N_11178);
xor U11250 (N_11250,N_11164,N_11082);
xor U11251 (N_11251,N_11197,N_11055);
and U11252 (N_11252,N_11064,N_11042);
xor U11253 (N_11253,N_11165,N_11187);
nor U11254 (N_11254,N_11129,N_11070);
and U11255 (N_11255,N_11146,N_11092);
nand U11256 (N_11256,N_11095,N_11190);
xnor U11257 (N_11257,N_11104,N_11151);
nand U11258 (N_11258,N_11136,N_11172);
nand U11259 (N_11259,N_11040,N_11189);
and U11260 (N_11260,N_11075,N_11166);
and U11261 (N_11261,N_11168,N_11097);
nand U11262 (N_11262,N_11074,N_11062);
nand U11263 (N_11263,N_11111,N_11079);
xor U11264 (N_11264,N_11137,N_11073);
nand U11265 (N_11265,N_11077,N_11122);
or U11266 (N_11266,N_11123,N_11102);
xor U11267 (N_11267,N_11195,N_11105);
and U11268 (N_11268,N_11063,N_11078);
nand U11269 (N_11269,N_11159,N_11133);
and U11270 (N_11270,N_11086,N_11112);
nor U11271 (N_11271,N_11177,N_11060);
nand U11272 (N_11272,N_11183,N_11186);
xor U11273 (N_11273,N_11109,N_11114);
xnor U11274 (N_11274,N_11067,N_11051);
nand U11275 (N_11275,N_11076,N_11141);
or U11276 (N_11276,N_11179,N_11046);
nand U11277 (N_11277,N_11157,N_11193);
nand U11278 (N_11278,N_11182,N_11100);
nor U11279 (N_11279,N_11173,N_11084);
nand U11280 (N_11280,N_11085,N_11136);
or U11281 (N_11281,N_11135,N_11153);
nand U11282 (N_11282,N_11168,N_11181);
nor U11283 (N_11283,N_11080,N_11150);
xor U11284 (N_11284,N_11067,N_11144);
and U11285 (N_11285,N_11068,N_11115);
or U11286 (N_11286,N_11162,N_11089);
nand U11287 (N_11287,N_11189,N_11128);
or U11288 (N_11288,N_11043,N_11077);
and U11289 (N_11289,N_11148,N_11059);
or U11290 (N_11290,N_11113,N_11107);
or U11291 (N_11291,N_11053,N_11049);
and U11292 (N_11292,N_11076,N_11078);
nand U11293 (N_11293,N_11184,N_11096);
xnor U11294 (N_11294,N_11132,N_11190);
or U11295 (N_11295,N_11075,N_11188);
nand U11296 (N_11296,N_11144,N_11147);
xnor U11297 (N_11297,N_11111,N_11069);
or U11298 (N_11298,N_11074,N_11152);
and U11299 (N_11299,N_11118,N_11052);
xnor U11300 (N_11300,N_11163,N_11166);
nand U11301 (N_11301,N_11164,N_11188);
nor U11302 (N_11302,N_11091,N_11181);
nor U11303 (N_11303,N_11077,N_11167);
xor U11304 (N_11304,N_11095,N_11169);
and U11305 (N_11305,N_11063,N_11097);
or U11306 (N_11306,N_11117,N_11167);
xnor U11307 (N_11307,N_11129,N_11056);
or U11308 (N_11308,N_11168,N_11164);
and U11309 (N_11309,N_11059,N_11135);
nand U11310 (N_11310,N_11139,N_11052);
nand U11311 (N_11311,N_11149,N_11157);
nor U11312 (N_11312,N_11189,N_11102);
and U11313 (N_11313,N_11059,N_11094);
nand U11314 (N_11314,N_11155,N_11097);
xnor U11315 (N_11315,N_11081,N_11109);
or U11316 (N_11316,N_11105,N_11077);
and U11317 (N_11317,N_11112,N_11188);
and U11318 (N_11318,N_11166,N_11140);
nand U11319 (N_11319,N_11128,N_11140);
xor U11320 (N_11320,N_11163,N_11097);
or U11321 (N_11321,N_11140,N_11079);
xor U11322 (N_11322,N_11107,N_11165);
or U11323 (N_11323,N_11196,N_11041);
or U11324 (N_11324,N_11085,N_11067);
or U11325 (N_11325,N_11081,N_11046);
and U11326 (N_11326,N_11151,N_11171);
nor U11327 (N_11327,N_11149,N_11064);
or U11328 (N_11328,N_11087,N_11118);
and U11329 (N_11329,N_11156,N_11046);
nor U11330 (N_11330,N_11132,N_11158);
xor U11331 (N_11331,N_11103,N_11053);
nor U11332 (N_11332,N_11199,N_11129);
nand U11333 (N_11333,N_11058,N_11151);
nand U11334 (N_11334,N_11128,N_11062);
nor U11335 (N_11335,N_11089,N_11111);
xnor U11336 (N_11336,N_11117,N_11155);
or U11337 (N_11337,N_11040,N_11129);
or U11338 (N_11338,N_11136,N_11061);
nor U11339 (N_11339,N_11067,N_11100);
or U11340 (N_11340,N_11134,N_11168);
nand U11341 (N_11341,N_11061,N_11047);
and U11342 (N_11342,N_11194,N_11118);
and U11343 (N_11343,N_11043,N_11086);
and U11344 (N_11344,N_11134,N_11095);
or U11345 (N_11345,N_11087,N_11055);
or U11346 (N_11346,N_11169,N_11150);
nor U11347 (N_11347,N_11048,N_11043);
or U11348 (N_11348,N_11086,N_11056);
and U11349 (N_11349,N_11156,N_11194);
nor U11350 (N_11350,N_11166,N_11098);
and U11351 (N_11351,N_11123,N_11044);
nand U11352 (N_11352,N_11113,N_11068);
or U11353 (N_11353,N_11127,N_11104);
and U11354 (N_11354,N_11166,N_11053);
xnor U11355 (N_11355,N_11146,N_11172);
and U11356 (N_11356,N_11112,N_11145);
nor U11357 (N_11357,N_11049,N_11181);
nand U11358 (N_11358,N_11190,N_11079);
xor U11359 (N_11359,N_11118,N_11113);
xnor U11360 (N_11360,N_11281,N_11344);
xor U11361 (N_11361,N_11222,N_11276);
nor U11362 (N_11362,N_11262,N_11261);
or U11363 (N_11363,N_11334,N_11238);
nand U11364 (N_11364,N_11308,N_11207);
or U11365 (N_11365,N_11215,N_11335);
xnor U11366 (N_11366,N_11309,N_11275);
or U11367 (N_11367,N_11211,N_11303);
and U11368 (N_11368,N_11305,N_11359);
nor U11369 (N_11369,N_11214,N_11205);
nand U11370 (N_11370,N_11299,N_11298);
nand U11371 (N_11371,N_11340,N_11267);
nand U11372 (N_11372,N_11322,N_11280);
and U11373 (N_11373,N_11239,N_11278);
nand U11374 (N_11374,N_11286,N_11225);
xor U11375 (N_11375,N_11354,N_11296);
and U11376 (N_11376,N_11217,N_11328);
nand U11377 (N_11377,N_11216,N_11333);
or U11378 (N_11378,N_11218,N_11332);
or U11379 (N_11379,N_11293,N_11264);
nor U11380 (N_11380,N_11345,N_11233);
or U11381 (N_11381,N_11337,N_11229);
and U11382 (N_11382,N_11226,N_11282);
nand U11383 (N_11383,N_11343,N_11350);
nor U11384 (N_11384,N_11237,N_11249);
nor U11385 (N_11385,N_11292,N_11266);
nor U11386 (N_11386,N_11324,N_11268);
nand U11387 (N_11387,N_11240,N_11279);
xor U11388 (N_11388,N_11304,N_11244);
nand U11389 (N_11389,N_11273,N_11269);
xnor U11390 (N_11390,N_11341,N_11212);
nand U11391 (N_11391,N_11355,N_11259);
nor U11392 (N_11392,N_11245,N_11295);
or U11393 (N_11393,N_11353,N_11256);
nor U11394 (N_11394,N_11310,N_11289);
nand U11395 (N_11395,N_11277,N_11321);
and U11396 (N_11396,N_11357,N_11231);
and U11397 (N_11397,N_11202,N_11342);
nand U11398 (N_11398,N_11203,N_11291);
nor U11399 (N_11399,N_11314,N_11301);
and U11400 (N_11400,N_11272,N_11250);
and U11401 (N_11401,N_11252,N_11336);
nand U11402 (N_11402,N_11297,N_11283);
and U11403 (N_11403,N_11230,N_11356);
nor U11404 (N_11404,N_11228,N_11204);
xor U11405 (N_11405,N_11316,N_11241);
and U11406 (N_11406,N_11320,N_11329);
and U11407 (N_11407,N_11294,N_11235);
nor U11408 (N_11408,N_11234,N_11288);
and U11409 (N_11409,N_11247,N_11220);
xnor U11410 (N_11410,N_11248,N_11223);
nor U11411 (N_11411,N_11284,N_11209);
nor U11412 (N_11412,N_11348,N_11274);
nor U11413 (N_11413,N_11253,N_11300);
or U11414 (N_11414,N_11349,N_11287);
xnor U11415 (N_11415,N_11257,N_11285);
or U11416 (N_11416,N_11346,N_11201);
nor U11417 (N_11417,N_11210,N_11260);
and U11418 (N_11418,N_11221,N_11254);
nand U11419 (N_11419,N_11246,N_11302);
nand U11420 (N_11420,N_11263,N_11312);
and U11421 (N_11421,N_11255,N_11347);
nand U11422 (N_11422,N_11315,N_11206);
nor U11423 (N_11423,N_11331,N_11325);
xnor U11424 (N_11424,N_11339,N_11352);
xnor U11425 (N_11425,N_11330,N_11271);
nand U11426 (N_11426,N_11213,N_11227);
or U11427 (N_11427,N_11326,N_11208);
or U11428 (N_11428,N_11338,N_11323);
nor U11429 (N_11429,N_11224,N_11306);
and U11430 (N_11430,N_11258,N_11200);
nor U11431 (N_11431,N_11251,N_11313);
or U11432 (N_11432,N_11219,N_11265);
xnor U11433 (N_11433,N_11307,N_11358);
xor U11434 (N_11434,N_11327,N_11351);
nand U11435 (N_11435,N_11318,N_11270);
nand U11436 (N_11436,N_11243,N_11311);
nor U11437 (N_11437,N_11236,N_11232);
xor U11438 (N_11438,N_11290,N_11242);
and U11439 (N_11439,N_11319,N_11317);
xnor U11440 (N_11440,N_11341,N_11210);
or U11441 (N_11441,N_11248,N_11340);
or U11442 (N_11442,N_11250,N_11212);
xnor U11443 (N_11443,N_11302,N_11201);
and U11444 (N_11444,N_11276,N_11251);
and U11445 (N_11445,N_11352,N_11305);
xnor U11446 (N_11446,N_11338,N_11354);
nor U11447 (N_11447,N_11332,N_11238);
and U11448 (N_11448,N_11334,N_11212);
or U11449 (N_11449,N_11271,N_11311);
nor U11450 (N_11450,N_11238,N_11221);
nor U11451 (N_11451,N_11310,N_11312);
nand U11452 (N_11452,N_11287,N_11247);
and U11453 (N_11453,N_11325,N_11279);
xnor U11454 (N_11454,N_11275,N_11333);
nand U11455 (N_11455,N_11291,N_11256);
nor U11456 (N_11456,N_11218,N_11310);
xor U11457 (N_11457,N_11315,N_11231);
and U11458 (N_11458,N_11331,N_11280);
nor U11459 (N_11459,N_11316,N_11202);
and U11460 (N_11460,N_11327,N_11239);
or U11461 (N_11461,N_11344,N_11234);
and U11462 (N_11462,N_11276,N_11249);
xnor U11463 (N_11463,N_11280,N_11219);
or U11464 (N_11464,N_11323,N_11210);
nand U11465 (N_11465,N_11336,N_11283);
or U11466 (N_11466,N_11218,N_11355);
nand U11467 (N_11467,N_11290,N_11289);
nor U11468 (N_11468,N_11300,N_11306);
and U11469 (N_11469,N_11350,N_11296);
nand U11470 (N_11470,N_11304,N_11291);
nor U11471 (N_11471,N_11321,N_11355);
or U11472 (N_11472,N_11309,N_11204);
and U11473 (N_11473,N_11337,N_11318);
and U11474 (N_11474,N_11228,N_11356);
nor U11475 (N_11475,N_11335,N_11297);
xnor U11476 (N_11476,N_11308,N_11313);
or U11477 (N_11477,N_11215,N_11260);
and U11478 (N_11478,N_11245,N_11228);
nand U11479 (N_11479,N_11333,N_11292);
or U11480 (N_11480,N_11317,N_11267);
or U11481 (N_11481,N_11204,N_11306);
xnor U11482 (N_11482,N_11216,N_11264);
nand U11483 (N_11483,N_11282,N_11219);
or U11484 (N_11484,N_11308,N_11258);
nor U11485 (N_11485,N_11234,N_11321);
and U11486 (N_11486,N_11288,N_11284);
xor U11487 (N_11487,N_11339,N_11321);
nand U11488 (N_11488,N_11336,N_11313);
nand U11489 (N_11489,N_11359,N_11264);
and U11490 (N_11490,N_11236,N_11280);
or U11491 (N_11491,N_11237,N_11357);
xnor U11492 (N_11492,N_11286,N_11253);
nor U11493 (N_11493,N_11213,N_11351);
and U11494 (N_11494,N_11268,N_11332);
and U11495 (N_11495,N_11202,N_11324);
nor U11496 (N_11496,N_11230,N_11304);
and U11497 (N_11497,N_11216,N_11254);
or U11498 (N_11498,N_11252,N_11311);
nand U11499 (N_11499,N_11249,N_11229);
nor U11500 (N_11500,N_11263,N_11310);
and U11501 (N_11501,N_11228,N_11343);
and U11502 (N_11502,N_11306,N_11280);
and U11503 (N_11503,N_11221,N_11320);
or U11504 (N_11504,N_11347,N_11318);
xnor U11505 (N_11505,N_11239,N_11221);
xnor U11506 (N_11506,N_11215,N_11281);
xnor U11507 (N_11507,N_11215,N_11213);
or U11508 (N_11508,N_11241,N_11332);
and U11509 (N_11509,N_11234,N_11302);
nand U11510 (N_11510,N_11308,N_11336);
or U11511 (N_11511,N_11280,N_11259);
xor U11512 (N_11512,N_11218,N_11209);
nor U11513 (N_11513,N_11249,N_11251);
or U11514 (N_11514,N_11233,N_11258);
nand U11515 (N_11515,N_11303,N_11276);
or U11516 (N_11516,N_11259,N_11267);
nand U11517 (N_11517,N_11259,N_11337);
nor U11518 (N_11518,N_11293,N_11302);
nor U11519 (N_11519,N_11350,N_11251);
xnor U11520 (N_11520,N_11497,N_11381);
and U11521 (N_11521,N_11452,N_11385);
and U11522 (N_11522,N_11370,N_11390);
or U11523 (N_11523,N_11489,N_11415);
or U11524 (N_11524,N_11514,N_11487);
xor U11525 (N_11525,N_11361,N_11365);
nor U11526 (N_11526,N_11461,N_11417);
or U11527 (N_11527,N_11379,N_11471);
xor U11528 (N_11528,N_11469,N_11380);
nand U11529 (N_11529,N_11445,N_11388);
nor U11530 (N_11530,N_11393,N_11446);
nand U11531 (N_11531,N_11439,N_11456);
nor U11532 (N_11532,N_11401,N_11421);
nand U11533 (N_11533,N_11396,N_11402);
xnor U11534 (N_11534,N_11389,N_11427);
xor U11535 (N_11535,N_11504,N_11400);
nor U11536 (N_11536,N_11418,N_11428);
or U11537 (N_11537,N_11425,N_11476);
xnor U11538 (N_11538,N_11500,N_11440);
nand U11539 (N_11539,N_11369,N_11399);
nor U11540 (N_11540,N_11431,N_11458);
nor U11541 (N_11541,N_11491,N_11515);
nor U11542 (N_11542,N_11477,N_11416);
nor U11543 (N_11543,N_11387,N_11368);
and U11544 (N_11544,N_11442,N_11486);
xor U11545 (N_11545,N_11375,N_11395);
and U11546 (N_11546,N_11510,N_11473);
or U11547 (N_11547,N_11429,N_11502);
nand U11548 (N_11548,N_11419,N_11362);
nor U11549 (N_11549,N_11466,N_11403);
xor U11550 (N_11550,N_11482,N_11410);
xor U11551 (N_11551,N_11516,N_11413);
and U11552 (N_11552,N_11468,N_11488);
nor U11553 (N_11553,N_11414,N_11411);
nand U11554 (N_11554,N_11437,N_11503);
or U11555 (N_11555,N_11378,N_11371);
or U11556 (N_11556,N_11518,N_11360);
nand U11557 (N_11557,N_11433,N_11470);
nand U11558 (N_11558,N_11441,N_11465);
nor U11559 (N_11559,N_11459,N_11506);
nand U11560 (N_11560,N_11480,N_11447);
nor U11561 (N_11561,N_11397,N_11454);
xor U11562 (N_11562,N_11460,N_11478);
nor U11563 (N_11563,N_11484,N_11376);
nor U11564 (N_11564,N_11505,N_11511);
nand U11565 (N_11565,N_11386,N_11485);
xor U11566 (N_11566,N_11422,N_11435);
and U11567 (N_11567,N_11404,N_11426);
xor U11568 (N_11568,N_11382,N_11507);
and U11569 (N_11569,N_11374,N_11408);
and U11570 (N_11570,N_11453,N_11443);
and U11571 (N_11571,N_11392,N_11501);
nand U11572 (N_11572,N_11517,N_11519);
and U11573 (N_11573,N_11444,N_11366);
nand U11574 (N_11574,N_11512,N_11508);
or U11575 (N_11575,N_11479,N_11457);
xor U11576 (N_11576,N_11436,N_11490);
nor U11577 (N_11577,N_11430,N_11463);
and U11578 (N_11578,N_11492,N_11407);
and U11579 (N_11579,N_11405,N_11409);
xnor U11580 (N_11580,N_11451,N_11391);
nand U11581 (N_11581,N_11495,N_11412);
xnor U11582 (N_11582,N_11432,N_11394);
or U11583 (N_11583,N_11467,N_11464);
xor U11584 (N_11584,N_11398,N_11367);
or U11585 (N_11585,N_11373,N_11496);
xnor U11586 (N_11586,N_11450,N_11494);
and U11587 (N_11587,N_11474,N_11434);
nand U11588 (N_11588,N_11462,N_11483);
nor U11589 (N_11589,N_11481,N_11383);
xor U11590 (N_11590,N_11509,N_11475);
nand U11591 (N_11591,N_11363,N_11438);
and U11592 (N_11592,N_11377,N_11406);
xor U11593 (N_11593,N_11455,N_11513);
xor U11594 (N_11594,N_11448,N_11372);
nand U11595 (N_11595,N_11424,N_11423);
nand U11596 (N_11596,N_11472,N_11384);
and U11597 (N_11597,N_11498,N_11364);
nor U11598 (N_11598,N_11499,N_11493);
and U11599 (N_11599,N_11449,N_11420);
and U11600 (N_11600,N_11382,N_11426);
or U11601 (N_11601,N_11404,N_11364);
xor U11602 (N_11602,N_11393,N_11365);
and U11603 (N_11603,N_11478,N_11386);
nor U11604 (N_11604,N_11426,N_11386);
xnor U11605 (N_11605,N_11380,N_11503);
or U11606 (N_11606,N_11421,N_11452);
or U11607 (N_11607,N_11383,N_11423);
or U11608 (N_11608,N_11478,N_11459);
nand U11609 (N_11609,N_11382,N_11433);
or U11610 (N_11610,N_11379,N_11416);
nand U11611 (N_11611,N_11380,N_11398);
or U11612 (N_11612,N_11436,N_11392);
xnor U11613 (N_11613,N_11487,N_11504);
and U11614 (N_11614,N_11388,N_11489);
and U11615 (N_11615,N_11369,N_11403);
nor U11616 (N_11616,N_11470,N_11390);
xor U11617 (N_11617,N_11474,N_11478);
xor U11618 (N_11618,N_11486,N_11434);
and U11619 (N_11619,N_11385,N_11382);
and U11620 (N_11620,N_11373,N_11423);
nand U11621 (N_11621,N_11370,N_11426);
nor U11622 (N_11622,N_11504,N_11464);
xor U11623 (N_11623,N_11405,N_11386);
and U11624 (N_11624,N_11391,N_11470);
and U11625 (N_11625,N_11501,N_11382);
nor U11626 (N_11626,N_11373,N_11405);
nor U11627 (N_11627,N_11459,N_11495);
and U11628 (N_11628,N_11385,N_11376);
xnor U11629 (N_11629,N_11447,N_11381);
nand U11630 (N_11630,N_11439,N_11494);
or U11631 (N_11631,N_11385,N_11506);
nand U11632 (N_11632,N_11394,N_11452);
nand U11633 (N_11633,N_11494,N_11513);
nand U11634 (N_11634,N_11491,N_11468);
xnor U11635 (N_11635,N_11366,N_11424);
or U11636 (N_11636,N_11398,N_11435);
nand U11637 (N_11637,N_11477,N_11430);
nand U11638 (N_11638,N_11429,N_11475);
xnor U11639 (N_11639,N_11512,N_11455);
nor U11640 (N_11640,N_11400,N_11456);
xnor U11641 (N_11641,N_11422,N_11415);
xnor U11642 (N_11642,N_11364,N_11371);
xor U11643 (N_11643,N_11410,N_11369);
or U11644 (N_11644,N_11427,N_11377);
nor U11645 (N_11645,N_11461,N_11386);
or U11646 (N_11646,N_11504,N_11441);
nor U11647 (N_11647,N_11436,N_11443);
nand U11648 (N_11648,N_11444,N_11368);
and U11649 (N_11649,N_11456,N_11393);
xnor U11650 (N_11650,N_11495,N_11364);
xor U11651 (N_11651,N_11500,N_11381);
xor U11652 (N_11652,N_11449,N_11424);
nand U11653 (N_11653,N_11485,N_11399);
and U11654 (N_11654,N_11491,N_11405);
nor U11655 (N_11655,N_11421,N_11367);
or U11656 (N_11656,N_11421,N_11455);
nand U11657 (N_11657,N_11402,N_11427);
xor U11658 (N_11658,N_11486,N_11378);
xnor U11659 (N_11659,N_11507,N_11504);
nand U11660 (N_11660,N_11512,N_11424);
nor U11661 (N_11661,N_11455,N_11503);
nand U11662 (N_11662,N_11396,N_11496);
xor U11663 (N_11663,N_11509,N_11393);
nor U11664 (N_11664,N_11361,N_11394);
nand U11665 (N_11665,N_11388,N_11435);
nor U11666 (N_11666,N_11468,N_11510);
or U11667 (N_11667,N_11438,N_11472);
or U11668 (N_11668,N_11483,N_11461);
nand U11669 (N_11669,N_11505,N_11492);
nor U11670 (N_11670,N_11448,N_11397);
xnor U11671 (N_11671,N_11511,N_11437);
or U11672 (N_11672,N_11406,N_11448);
or U11673 (N_11673,N_11435,N_11417);
or U11674 (N_11674,N_11484,N_11486);
or U11675 (N_11675,N_11472,N_11425);
nand U11676 (N_11676,N_11504,N_11467);
nand U11677 (N_11677,N_11401,N_11431);
and U11678 (N_11678,N_11442,N_11409);
nand U11679 (N_11679,N_11438,N_11406);
nor U11680 (N_11680,N_11537,N_11555);
nand U11681 (N_11681,N_11656,N_11668);
and U11682 (N_11682,N_11593,N_11523);
or U11683 (N_11683,N_11526,N_11679);
nand U11684 (N_11684,N_11569,N_11650);
nand U11685 (N_11685,N_11578,N_11662);
nand U11686 (N_11686,N_11648,N_11675);
xnor U11687 (N_11687,N_11587,N_11597);
nand U11688 (N_11688,N_11592,N_11619);
nor U11689 (N_11689,N_11577,N_11630);
nand U11690 (N_11690,N_11584,N_11653);
nor U11691 (N_11691,N_11628,N_11599);
xor U11692 (N_11692,N_11548,N_11525);
or U11693 (N_11693,N_11557,N_11612);
or U11694 (N_11694,N_11573,N_11571);
and U11695 (N_11695,N_11524,N_11589);
and U11696 (N_11696,N_11546,N_11608);
or U11697 (N_11697,N_11620,N_11545);
nor U11698 (N_11698,N_11536,N_11605);
nor U11699 (N_11699,N_11576,N_11530);
nor U11700 (N_11700,N_11561,N_11601);
nor U11701 (N_11701,N_11666,N_11638);
nor U11702 (N_11702,N_11583,N_11582);
nand U11703 (N_11703,N_11618,N_11538);
and U11704 (N_11704,N_11520,N_11640);
nor U11705 (N_11705,N_11636,N_11560);
nor U11706 (N_11706,N_11678,N_11667);
or U11707 (N_11707,N_11602,N_11609);
and U11708 (N_11708,N_11529,N_11623);
nor U11709 (N_11709,N_11615,N_11659);
and U11710 (N_11710,N_11598,N_11677);
and U11711 (N_11711,N_11532,N_11559);
xnor U11712 (N_11712,N_11616,N_11629);
xor U11713 (N_11713,N_11527,N_11558);
or U11714 (N_11714,N_11676,N_11534);
nand U11715 (N_11715,N_11551,N_11544);
or U11716 (N_11716,N_11586,N_11617);
or U11717 (N_11717,N_11625,N_11565);
nand U11718 (N_11718,N_11541,N_11531);
and U11719 (N_11719,N_11591,N_11624);
nor U11720 (N_11720,N_11632,N_11654);
or U11721 (N_11721,N_11631,N_11674);
or U11722 (N_11722,N_11610,N_11580);
and U11723 (N_11723,N_11658,N_11622);
nor U11724 (N_11724,N_11600,N_11581);
xnor U11725 (N_11725,N_11673,N_11595);
nor U11726 (N_11726,N_11594,N_11626);
or U11727 (N_11727,N_11566,N_11661);
xnor U11728 (N_11728,N_11547,N_11554);
nand U11729 (N_11729,N_11647,N_11635);
nand U11730 (N_11730,N_11613,N_11564);
nor U11731 (N_11731,N_11549,N_11649);
and U11732 (N_11732,N_11611,N_11671);
and U11733 (N_11733,N_11634,N_11552);
or U11734 (N_11734,N_11535,N_11563);
nor U11735 (N_11735,N_11579,N_11642);
nor U11736 (N_11736,N_11663,N_11540);
and U11737 (N_11737,N_11596,N_11539);
xnor U11738 (N_11738,N_11521,N_11657);
nor U11739 (N_11739,N_11572,N_11655);
xnor U11740 (N_11740,N_11543,N_11669);
nor U11741 (N_11741,N_11585,N_11588);
or U11742 (N_11742,N_11652,N_11570);
nor U11743 (N_11743,N_11550,N_11533);
or U11744 (N_11744,N_11574,N_11651);
nor U11745 (N_11745,N_11633,N_11621);
nand U11746 (N_11746,N_11604,N_11562);
xor U11747 (N_11747,N_11603,N_11670);
and U11748 (N_11748,N_11641,N_11644);
xor U11749 (N_11749,N_11664,N_11522);
xnor U11750 (N_11750,N_11643,N_11553);
xnor U11751 (N_11751,N_11660,N_11567);
nand U11752 (N_11752,N_11639,N_11590);
xor U11753 (N_11753,N_11528,N_11672);
xnor U11754 (N_11754,N_11665,N_11556);
nor U11755 (N_11755,N_11627,N_11606);
or U11756 (N_11756,N_11645,N_11614);
nand U11757 (N_11757,N_11637,N_11568);
and U11758 (N_11758,N_11646,N_11542);
and U11759 (N_11759,N_11575,N_11607);
or U11760 (N_11760,N_11574,N_11584);
nor U11761 (N_11761,N_11606,N_11641);
and U11762 (N_11762,N_11662,N_11631);
and U11763 (N_11763,N_11676,N_11599);
xor U11764 (N_11764,N_11658,N_11621);
nor U11765 (N_11765,N_11586,N_11618);
nor U11766 (N_11766,N_11602,N_11560);
or U11767 (N_11767,N_11539,N_11664);
and U11768 (N_11768,N_11554,N_11558);
nand U11769 (N_11769,N_11620,N_11574);
or U11770 (N_11770,N_11595,N_11535);
and U11771 (N_11771,N_11621,N_11654);
nand U11772 (N_11772,N_11652,N_11581);
xor U11773 (N_11773,N_11613,N_11621);
nand U11774 (N_11774,N_11546,N_11559);
nand U11775 (N_11775,N_11522,N_11676);
or U11776 (N_11776,N_11575,N_11622);
nand U11777 (N_11777,N_11565,N_11578);
or U11778 (N_11778,N_11602,N_11611);
or U11779 (N_11779,N_11580,N_11543);
and U11780 (N_11780,N_11649,N_11551);
nor U11781 (N_11781,N_11678,N_11553);
nor U11782 (N_11782,N_11565,N_11566);
nand U11783 (N_11783,N_11526,N_11676);
and U11784 (N_11784,N_11633,N_11608);
and U11785 (N_11785,N_11568,N_11589);
or U11786 (N_11786,N_11558,N_11648);
xnor U11787 (N_11787,N_11607,N_11678);
and U11788 (N_11788,N_11561,N_11566);
xor U11789 (N_11789,N_11606,N_11664);
and U11790 (N_11790,N_11618,N_11559);
nand U11791 (N_11791,N_11634,N_11535);
nand U11792 (N_11792,N_11590,N_11598);
nor U11793 (N_11793,N_11613,N_11522);
or U11794 (N_11794,N_11585,N_11650);
nor U11795 (N_11795,N_11523,N_11618);
nand U11796 (N_11796,N_11670,N_11605);
xor U11797 (N_11797,N_11567,N_11613);
and U11798 (N_11798,N_11573,N_11643);
nand U11799 (N_11799,N_11633,N_11593);
nand U11800 (N_11800,N_11659,N_11568);
xor U11801 (N_11801,N_11619,N_11611);
or U11802 (N_11802,N_11659,N_11580);
or U11803 (N_11803,N_11654,N_11552);
nor U11804 (N_11804,N_11659,N_11602);
or U11805 (N_11805,N_11664,N_11626);
and U11806 (N_11806,N_11638,N_11675);
xor U11807 (N_11807,N_11616,N_11591);
xor U11808 (N_11808,N_11523,N_11647);
nand U11809 (N_11809,N_11612,N_11657);
or U11810 (N_11810,N_11611,N_11525);
or U11811 (N_11811,N_11641,N_11653);
nor U11812 (N_11812,N_11614,N_11572);
nand U11813 (N_11813,N_11536,N_11656);
nor U11814 (N_11814,N_11524,N_11650);
nor U11815 (N_11815,N_11623,N_11556);
and U11816 (N_11816,N_11644,N_11527);
nand U11817 (N_11817,N_11629,N_11580);
or U11818 (N_11818,N_11544,N_11669);
nor U11819 (N_11819,N_11548,N_11625);
xnor U11820 (N_11820,N_11569,N_11591);
and U11821 (N_11821,N_11534,N_11603);
xnor U11822 (N_11822,N_11638,N_11546);
and U11823 (N_11823,N_11596,N_11607);
nor U11824 (N_11824,N_11591,N_11582);
and U11825 (N_11825,N_11676,N_11669);
nand U11826 (N_11826,N_11601,N_11541);
and U11827 (N_11827,N_11634,N_11551);
and U11828 (N_11828,N_11664,N_11631);
xnor U11829 (N_11829,N_11592,N_11659);
nand U11830 (N_11830,N_11643,N_11530);
nand U11831 (N_11831,N_11642,N_11526);
nand U11832 (N_11832,N_11561,N_11557);
nand U11833 (N_11833,N_11595,N_11598);
nand U11834 (N_11834,N_11596,N_11594);
and U11835 (N_11835,N_11579,N_11626);
nor U11836 (N_11836,N_11535,N_11667);
xor U11837 (N_11837,N_11645,N_11578);
nand U11838 (N_11838,N_11622,N_11675);
nor U11839 (N_11839,N_11600,N_11617);
or U11840 (N_11840,N_11767,N_11768);
and U11841 (N_11841,N_11839,N_11809);
nand U11842 (N_11842,N_11755,N_11723);
nor U11843 (N_11843,N_11731,N_11813);
and U11844 (N_11844,N_11729,N_11690);
xor U11845 (N_11845,N_11707,N_11700);
xnor U11846 (N_11846,N_11834,N_11792);
nand U11847 (N_11847,N_11769,N_11753);
or U11848 (N_11848,N_11796,N_11742);
xor U11849 (N_11849,N_11681,N_11757);
xnor U11850 (N_11850,N_11746,N_11697);
xnor U11851 (N_11851,N_11737,N_11775);
or U11852 (N_11852,N_11763,N_11682);
or U11853 (N_11853,N_11725,N_11803);
and U11854 (N_11854,N_11806,N_11710);
and U11855 (N_11855,N_11774,N_11754);
or U11856 (N_11856,N_11777,N_11801);
nand U11857 (N_11857,N_11705,N_11693);
or U11858 (N_11858,N_11751,N_11822);
nor U11859 (N_11859,N_11815,N_11764);
xor U11860 (N_11860,N_11817,N_11699);
or U11861 (N_11861,N_11683,N_11685);
and U11862 (N_11862,N_11738,N_11826);
nor U11863 (N_11863,N_11706,N_11837);
xnor U11864 (N_11864,N_11836,N_11788);
nor U11865 (N_11865,N_11692,N_11807);
and U11866 (N_11866,N_11712,N_11698);
nand U11867 (N_11867,N_11745,N_11714);
nor U11868 (N_11868,N_11695,N_11829);
nor U11869 (N_11869,N_11747,N_11821);
xnor U11870 (N_11870,N_11684,N_11736);
nand U11871 (N_11871,N_11761,N_11766);
xor U11872 (N_11872,N_11790,N_11818);
nand U11873 (N_11873,N_11743,N_11770);
or U11874 (N_11874,N_11716,N_11730);
nor U11875 (N_11875,N_11687,N_11835);
xor U11876 (N_11876,N_11734,N_11794);
xor U11877 (N_11877,N_11711,N_11787);
nor U11878 (N_11878,N_11779,N_11782);
and U11879 (N_11879,N_11820,N_11810);
nor U11880 (N_11880,N_11830,N_11696);
nor U11881 (N_11881,N_11781,N_11776);
nor U11882 (N_11882,N_11748,N_11709);
or U11883 (N_11883,N_11694,N_11728);
nand U11884 (N_11884,N_11828,N_11702);
or U11885 (N_11885,N_11780,N_11739);
or U11886 (N_11886,N_11726,N_11772);
nand U11887 (N_11887,N_11758,N_11733);
or U11888 (N_11888,N_11811,N_11759);
and U11889 (N_11889,N_11816,N_11715);
nand U11890 (N_11890,N_11804,N_11778);
nor U11891 (N_11891,N_11823,N_11785);
xnor U11892 (N_11892,N_11740,N_11691);
nand U11893 (N_11893,N_11784,N_11686);
nor U11894 (N_11894,N_11773,N_11741);
nor U11895 (N_11895,N_11720,N_11832);
or U11896 (N_11896,N_11833,N_11744);
nor U11897 (N_11897,N_11762,N_11789);
or U11898 (N_11898,N_11689,N_11795);
nand U11899 (N_11899,N_11808,N_11708);
nand U11900 (N_11900,N_11812,N_11749);
xnor U11901 (N_11901,N_11799,N_11713);
or U11902 (N_11902,N_11831,N_11838);
and U11903 (N_11903,N_11722,N_11819);
nand U11904 (N_11904,N_11703,N_11824);
nor U11905 (N_11905,N_11814,N_11756);
or U11906 (N_11906,N_11805,N_11750);
or U11907 (N_11907,N_11793,N_11727);
nor U11908 (N_11908,N_11771,N_11798);
or U11909 (N_11909,N_11802,N_11800);
or U11910 (N_11910,N_11797,N_11791);
nand U11911 (N_11911,N_11721,N_11825);
and U11912 (N_11912,N_11732,N_11704);
nor U11913 (N_11913,N_11786,N_11719);
nand U11914 (N_11914,N_11717,N_11765);
xnor U11915 (N_11915,N_11752,N_11688);
and U11916 (N_11916,N_11724,N_11760);
nor U11917 (N_11917,N_11783,N_11701);
nor U11918 (N_11918,N_11718,N_11827);
nand U11919 (N_11919,N_11735,N_11680);
and U11920 (N_11920,N_11791,N_11710);
xnor U11921 (N_11921,N_11790,N_11687);
xor U11922 (N_11922,N_11838,N_11726);
and U11923 (N_11923,N_11800,N_11723);
and U11924 (N_11924,N_11815,N_11684);
nand U11925 (N_11925,N_11748,N_11715);
and U11926 (N_11926,N_11785,N_11734);
xor U11927 (N_11927,N_11747,N_11759);
nand U11928 (N_11928,N_11777,N_11715);
xnor U11929 (N_11929,N_11716,N_11739);
nand U11930 (N_11930,N_11826,N_11765);
or U11931 (N_11931,N_11824,N_11806);
nor U11932 (N_11932,N_11722,N_11831);
or U11933 (N_11933,N_11736,N_11700);
nand U11934 (N_11934,N_11689,N_11783);
or U11935 (N_11935,N_11706,N_11780);
and U11936 (N_11936,N_11801,N_11832);
xor U11937 (N_11937,N_11783,N_11780);
or U11938 (N_11938,N_11791,N_11796);
and U11939 (N_11939,N_11794,N_11720);
nor U11940 (N_11940,N_11705,N_11730);
or U11941 (N_11941,N_11685,N_11827);
nor U11942 (N_11942,N_11740,N_11753);
nand U11943 (N_11943,N_11784,N_11772);
xor U11944 (N_11944,N_11823,N_11753);
nand U11945 (N_11945,N_11806,N_11766);
nor U11946 (N_11946,N_11828,N_11680);
nand U11947 (N_11947,N_11750,N_11753);
xor U11948 (N_11948,N_11800,N_11773);
nor U11949 (N_11949,N_11823,N_11811);
and U11950 (N_11950,N_11757,N_11735);
and U11951 (N_11951,N_11698,N_11743);
and U11952 (N_11952,N_11771,N_11745);
and U11953 (N_11953,N_11738,N_11686);
and U11954 (N_11954,N_11685,N_11736);
and U11955 (N_11955,N_11821,N_11824);
or U11956 (N_11956,N_11771,N_11692);
and U11957 (N_11957,N_11773,N_11751);
or U11958 (N_11958,N_11788,N_11729);
nand U11959 (N_11959,N_11738,N_11740);
xnor U11960 (N_11960,N_11794,N_11698);
nand U11961 (N_11961,N_11715,N_11732);
or U11962 (N_11962,N_11687,N_11822);
nor U11963 (N_11963,N_11817,N_11690);
or U11964 (N_11964,N_11813,N_11693);
nor U11965 (N_11965,N_11798,N_11723);
or U11966 (N_11966,N_11798,N_11833);
nand U11967 (N_11967,N_11740,N_11704);
or U11968 (N_11968,N_11790,N_11745);
or U11969 (N_11969,N_11723,N_11754);
nor U11970 (N_11970,N_11778,N_11766);
and U11971 (N_11971,N_11722,N_11715);
and U11972 (N_11972,N_11805,N_11722);
or U11973 (N_11973,N_11695,N_11783);
or U11974 (N_11974,N_11787,N_11775);
nor U11975 (N_11975,N_11680,N_11781);
and U11976 (N_11976,N_11715,N_11779);
and U11977 (N_11977,N_11718,N_11817);
or U11978 (N_11978,N_11784,N_11781);
nand U11979 (N_11979,N_11734,N_11827);
xnor U11980 (N_11980,N_11814,N_11807);
nand U11981 (N_11981,N_11790,N_11726);
and U11982 (N_11982,N_11826,N_11832);
and U11983 (N_11983,N_11828,N_11731);
and U11984 (N_11984,N_11742,N_11838);
nor U11985 (N_11985,N_11682,N_11710);
xor U11986 (N_11986,N_11771,N_11814);
xor U11987 (N_11987,N_11696,N_11804);
nor U11988 (N_11988,N_11819,N_11689);
nor U11989 (N_11989,N_11805,N_11767);
xnor U11990 (N_11990,N_11720,N_11788);
nand U11991 (N_11991,N_11722,N_11701);
nand U11992 (N_11992,N_11700,N_11837);
and U11993 (N_11993,N_11824,N_11747);
xor U11994 (N_11994,N_11702,N_11746);
nand U11995 (N_11995,N_11833,N_11803);
or U11996 (N_11996,N_11751,N_11810);
or U11997 (N_11997,N_11709,N_11762);
and U11998 (N_11998,N_11722,N_11783);
and U11999 (N_11999,N_11696,N_11712);
and U12000 (N_12000,N_11916,N_11942);
nor U12001 (N_12001,N_11968,N_11992);
nand U12002 (N_12002,N_11840,N_11884);
nor U12003 (N_12003,N_11872,N_11876);
xnor U12004 (N_12004,N_11981,N_11874);
and U12005 (N_12005,N_11856,N_11920);
and U12006 (N_12006,N_11950,N_11843);
and U12007 (N_12007,N_11993,N_11890);
and U12008 (N_12008,N_11980,N_11955);
nand U12009 (N_12009,N_11889,N_11854);
and U12010 (N_12010,N_11989,N_11937);
nand U12011 (N_12011,N_11912,N_11978);
nor U12012 (N_12012,N_11859,N_11971);
and U12013 (N_12013,N_11998,N_11897);
and U12014 (N_12014,N_11936,N_11844);
or U12015 (N_12015,N_11893,N_11963);
nor U12016 (N_12016,N_11932,N_11858);
and U12017 (N_12017,N_11903,N_11848);
and U12018 (N_12018,N_11841,N_11952);
nor U12019 (N_12019,N_11961,N_11883);
nor U12020 (N_12020,N_11923,N_11985);
nor U12021 (N_12021,N_11852,N_11954);
or U12022 (N_12022,N_11972,N_11970);
and U12023 (N_12023,N_11875,N_11924);
or U12024 (N_12024,N_11886,N_11973);
nor U12025 (N_12025,N_11965,N_11927);
nand U12026 (N_12026,N_11966,N_11990);
nor U12027 (N_12027,N_11846,N_11995);
and U12028 (N_12028,N_11987,N_11899);
xor U12029 (N_12029,N_11896,N_11901);
nor U12030 (N_12030,N_11929,N_11917);
xor U12031 (N_12031,N_11911,N_11957);
and U12032 (N_12032,N_11845,N_11918);
nor U12033 (N_12033,N_11898,N_11958);
or U12034 (N_12034,N_11847,N_11914);
or U12035 (N_12035,N_11870,N_11947);
nand U12036 (N_12036,N_11956,N_11988);
nor U12037 (N_12037,N_11888,N_11865);
and U12038 (N_12038,N_11913,N_11930);
or U12039 (N_12039,N_11976,N_11895);
or U12040 (N_12040,N_11967,N_11868);
nand U12041 (N_12041,N_11850,N_11964);
and U12042 (N_12042,N_11991,N_11938);
nor U12043 (N_12043,N_11842,N_11994);
and U12044 (N_12044,N_11922,N_11941);
xnor U12045 (N_12045,N_11984,N_11935);
nand U12046 (N_12046,N_11919,N_11879);
nor U12047 (N_12047,N_11860,N_11887);
xnor U12048 (N_12048,N_11880,N_11939);
nand U12049 (N_12049,N_11864,N_11974);
or U12050 (N_12050,N_11905,N_11885);
nor U12051 (N_12051,N_11851,N_11892);
or U12052 (N_12052,N_11933,N_11982);
or U12053 (N_12053,N_11910,N_11960);
nor U12054 (N_12054,N_11902,N_11873);
and U12055 (N_12055,N_11959,N_11948);
nand U12056 (N_12056,N_11849,N_11869);
or U12057 (N_12057,N_11857,N_11943);
nor U12058 (N_12058,N_11878,N_11909);
xor U12059 (N_12059,N_11866,N_11940);
xor U12060 (N_12060,N_11953,N_11894);
nor U12061 (N_12061,N_11977,N_11906);
nand U12062 (N_12062,N_11983,N_11945);
or U12063 (N_12063,N_11962,N_11997);
and U12064 (N_12064,N_11877,N_11881);
nor U12065 (N_12065,N_11855,N_11979);
xnor U12066 (N_12066,N_11951,N_11928);
or U12067 (N_12067,N_11867,N_11931);
nand U12068 (N_12068,N_11871,N_11969);
and U12069 (N_12069,N_11853,N_11949);
nand U12070 (N_12070,N_11861,N_11934);
or U12071 (N_12071,N_11891,N_11926);
or U12072 (N_12072,N_11863,N_11915);
nor U12073 (N_12073,N_11986,N_11862);
and U12074 (N_12074,N_11904,N_11975);
nor U12075 (N_12075,N_11946,N_11907);
nand U12076 (N_12076,N_11999,N_11921);
xor U12077 (N_12077,N_11900,N_11944);
nand U12078 (N_12078,N_11908,N_11882);
nor U12079 (N_12079,N_11925,N_11996);
and U12080 (N_12080,N_11980,N_11922);
nand U12081 (N_12081,N_11995,N_11930);
nor U12082 (N_12082,N_11889,N_11960);
and U12083 (N_12083,N_11847,N_11876);
nor U12084 (N_12084,N_11916,N_11917);
xnor U12085 (N_12085,N_11990,N_11980);
nor U12086 (N_12086,N_11875,N_11904);
nand U12087 (N_12087,N_11851,N_11923);
and U12088 (N_12088,N_11979,N_11985);
or U12089 (N_12089,N_11880,N_11960);
nand U12090 (N_12090,N_11915,N_11996);
and U12091 (N_12091,N_11952,N_11960);
or U12092 (N_12092,N_11851,N_11960);
xnor U12093 (N_12093,N_11880,N_11847);
or U12094 (N_12094,N_11920,N_11937);
or U12095 (N_12095,N_11988,N_11963);
or U12096 (N_12096,N_11949,N_11935);
or U12097 (N_12097,N_11976,N_11907);
xor U12098 (N_12098,N_11863,N_11860);
nor U12099 (N_12099,N_11973,N_11862);
nor U12100 (N_12100,N_11953,N_11974);
or U12101 (N_12101,N_11905,N_11926);
nor U12102 (N_12102,N_11999,N_11988);
nor U12103 (N_12103,N_11844,N_11842);
or U12104 (N_12104,N_11888,N_11993);
or U12105 (N_12105,N_11890,N_11989);
xnor U12106 (N_12106,N_11996,N_11942);
nor U12107 (N_12107,N_11929,N_11992);
or U12108 (N_12108,N_11953,N_11986);
or U12109 (N_12109,N_11979,N_11916);
xor U12110 (N_12110,N_11876,N_11954);
or U12111 (N_12111,N_11927,N_11895);
or U12112 (N_12112,N_11981,N_11949);
and U12113 (N_12113,N_11880,N_11954);
nand U12114 (N_12114,N_11974,N_11944);
xnor U12115 (N_12115,N_11881,N_11974);
xnor U12116 (N_12116,N_11920,N_11843);
or U12117 (N_12117,N_11992,N_11919);
or U12118 (N_12118,N_11951,N_11850);
nand U12119 (N_12119,N_11853,N_11851);
or U12120 (N_12120,N_11878,N_11898);
and U12121 (N_12121,N_11890,N_11933);
or U12122 (N_12122,N_11951,N_11996);
and U12123 (N_12123,N_11875,N_11994);
xor U12124 (N_12124,N_11958,N_11963);
nand U12125 (N_12125,N_11840,N_11926);
xnor U12126 (N_12126,N_11859,N_11988);
and U12127 (N_12127,N_11872,N_11986);
and U12128 (N_12128,N_11849,N_11999);
nand U12129 (N_12129,N_11856,N_11894);
nand U12130 (N_12130,N_11851,N_11898);
or U12131 (N_12131,N_11987,N_11843);
nor U12132 (N_12132,N_11967,N_11910);
nor U12133 (N_12133,N_11860,N_11877);
or U12134 (N_12134,N_11912,N_11869);
or U12135 (N_12135,N_11870,N_11845);
xor U12136 (N_12136,N_11868,N_11891);
nor U12137 (N_12137,N_11974,N_11885);
nor U12138 (N_12138,N_11945,N_11840);
xnor U12139 (N_12139,N_11878,N_11928);
and U12140 (N_12140,N_11906,N_11973);
nand U12141 (N_12141,N_11916,N_11897);
or U12142 (N_12142,N_11985,N_11867);
xor U12143 (N_12143,N_11909,N_11970);
and U12144 (N_12144,N_11973,N_11888);
nand U12145 (N_12145,N_11906,N_11985);
nor U12146 (N_12146,N_11846,N_11844);
and U12147 (N_12147,N_11976,N_11861);
nand U12148 (N_12148,N_11899,N_11890);
xnor U12149 (N_12149,N_11964,N_11961);
or U12150 (N_12150,N_11993,N_11978);
nand U12151 (N_12151,N_11925,N_11844);
nor U12152 (N_12152,N_11975,N_11890);
nand U12153 (N_12153,N_11921,N_11973);
xor U12154 (N_12154,N_11936,N_11974);
nor U12155 (N_12155,N_11849,N_11858);
and U12156 (N_12156,N_11872,N_11979);
and U12157 (N_12157,N_11972,N_11883);
xnor U12158 (N_12158,N_11900,N_11850);
xor U12159 (N_12159,N_11865,N_11937);
or U12160 (N_12160,N_12143,N_12157);
nor U12161 (N_12161,N_12005,N_12061);
nor U12162 (N_12162,N_12091,N_12104);
xnor U12163 (N_12163,N_12011,N_12036);
or U12164 (N_12164,N_12093,N_12046);
or U12165 (N_12165,N_12045,N_12142);
or U12166 (N_12166,N_12136,N_12101);
nand U12167 (N_12167,N_12065,N_12001);
or U12168 (N_12168,N_12112,N_12014);
nand U12169 (N_12169,N_12057,N_12135);
xor U12170 (N_12170,N_12123,N_12009);
xnor U12171 (N_12171,N_12152,N_12090);
xnor U12172 (N_12172,N_12086,N_12035);
nor U12173 (N_12173,N_12103,N_12037);
or U12174 (N_12174,N_12017,N_12121);
nor U12175 (N_12175,N_12146,N_12062);
or U12176 (N_12176,N_12088,N_12099);
and U12177 (N_12177,N_12117,N_12085);
nand U12178 (N_12178,N_12108,N_12008);
and U12179 (N_12179,N_12052,N_12056);
xor U12180 (N_12180,N_12082,N_12126);
and U12181 (N_12181,N_12129,N_12138);
xnor U12182 (N_12182,N_12071,N_12111);
nor U12183 (N_12183,N_12154,N_12026);
nor U12184 (N_12184,N_12076,N_12107);
xnor U12185 (N_12185,N_12075,N_12092);
or U12186 (N_12186,N_12084,N_12125);
xnor U12187 (N_12187,N_12079,N_12033);
nor U12188 (N_12188,N_12119,N_12128);
or U12189 (N_12189,N_12127,N_12055);
nand U12190 (N_12190,N_12069,N_12042);
xor U12191 (N_12191,N_12087,N_12053);
xor U12192 (N_12192,N_12124,N_12106);
nor U12193 (N_12193,N_12156,N_12151);
or U12194 (N_12194,N_12081,N_12133);
and U12195 (N_12195,N_12067,N_12066);
nand U12196 (N_12196,N_12020,N_12004);
or U12197 (N_12197,N_12145,N_12027);
nand U12198 (N_12198,N_12019,N_12010);
xnor U12199 (N_12199,N_12043,N_12131);
xnor U12200 (N_12200,N_12050,N_12058);
nand U12201 (N_12201,N_12149,N_12102);
nand U12202 (N_12202,N_12049,N_12158);
or U12203 (N_12203,N_12115,N_12024);
nand U12204 (N_12204,N_12021,N_12083);
nor U12205 (N_12205,N_12132,N_12063);
nand U12206 (N_12206,N_12038,N_12059);
and U12207 (N_12207,N_12113,N_12002);
xor U12208 (N_12208,N_12064,N_12012);
and U12209 (N_12209,N_12007,N_12013);
nor U12210 (N_12210,N_12122,N_12095);
nor U12211 (N_12211,N_12097,N_12006);
and U12212 (N_12212,N_12144,N_12039);
and U12213 (N_12213,N_12034,N_12100);
nand U12214 (N_12214,N_12077,N_12048);
or U12215 (N_12215,N_12047,N_12070);
xnor U12216 (N_12216,N_12110,N_12016);
and U12217 (N_12217,N_12148,N_12023);
or U12218 (N_12218,N_12096,N_12015);
xor U12219 (N_12219,N_12018,N_12028);
xor U12220 (N_12220,N_12098,N_12022);
and U12221 (N_12221,N_12051,N_12155);
nor U12222 (N_12222,N_12060,N_12032);
nor U12223 (N_12223,N_12147,N_12078);
and U12224 (N_12224,N_12109,N_12031);
nand U12225 (N_12225,N_12040,N_12130);
or U12226 (N_12226,N_12068,N_12072);
or U12227 (N_12227,N_12141,N_12118);
xnor U12228 (N_12228,N_12139,N_12041);
or U12229 (N_12229,N_12120,N_12105);
nor U12230 (N_12230,N_12044,N_12080);
nor U12231 (N_12231,N_12116,N_12000);
or U12232 (N_12232,N_12140,N_12159);
nand U12233 (N_12233,N_12089,N_12134);
xor U12234 (N_12234,N_12054,N_12025);
or U12235 (N_12235,N_12074,N_12003);
nand U12236 (N_12236,N_12094,N_12030);
and U12237 (N_12237,N_12029,N_12150);
nand U12238 (N_12238,N_12153,N_12073);
nand U12239 (N_12239,N_12137,N_12114);
or U12240 (N_12240,N_12028,N_12138);
nor U12241 (N_12241,N_12099,N_12127);
or U12242 (N_12242,N_12052,N_12007);
or U12243 (N_12243,N_12061,N_12102);
nand U12244 (N_12244,N_12112,N_12141);
nand U12245 (N_12245,N_12020,N_12027);
or U12246 (N_12246,N_12007,N_12106);
and U12247 (N_12247,N_12047,N_12029);
and U12248 (N_12248,N_12100,N_12124);
xor U12249 (N_12249,N_12053,N_12041);
nor U12250 (N_12250,N_12055,N_12051);
nor U12251 (N_12251,N_12075,N_12019);
and U12252 (N_12252,N_12080,N_12154);
xor U12253 (N_12253,N_12048,N_12020);
xor U12254 (N_12254,N_12115,N_12102);
nand U12255 (N_12255,N_12036,N_12054);
nor U12256 (N_12256,N_12056,N_12066);
nand U12257 (N_12257,N_12120,N_12137);
nor U12258 (N_12258,N_12111,N_12038);
or U12259 (N_12259,N_12054,N_12092);
nor U12260 (N_12260,N_12042,N_12002);
xnor U12261 (N_12261,N_12118,N_12102);
xnor U12262 (N_12262,N_12018,N_12001);
nor U12263 (N_12263,N_12154,N_12043);
xor U12264 (N_12264,N_12002,N_12117);
nor U12265 (N_12265,N_12053,N_12068);
nor U12266 (N_12266,N_12152,N_12080);
xor U12267 (N_12267,N_12062,N_12139);
and U12268 (N_12268,N_12135,N_12098);
xor U12269 (N_12269,N_12004,N_12071);
nand U12270 (N_12270,N_12141,N_12032);
nor U12271 (N_12271,N_12025,N_12115);
nand U12272 (N_12272,N_12158,N_12084);
nor U12273 (N_12273,N_12123,N_12043);
or U12274 (N_12274,N_12139,N_12049);
nor U12275 (N_12275,N_12044,N_12053);
nor U12276 (N_12276,N_12059,N_12105);
nor U12277 (N_12277,N_12017,N_12032);
nor U12278 (N_12278,N_12146,N_12148);
or U12279 (N_12279,N_12072,N_12150);
xnor U12280 (N_12280,N_12057,N_12147);
or U12281 (N_12281,N_12062,N_12044);
nand U12282 (N_12282,N_12130,N_12030);
nor U12283 (N_12283,N_12039,N_12031);
and U12284 (N_12284,N_12057,N_12034);
nand U12285 (N_12285,N_12122,N_12033);
nor U12286 (N_12286,N_12145,N_12016);
or U12287 (N_12287,N_12082,N_12072);
and U12288 (N_12288,N_12056,N_12046);
xor U12289 (N_12289,N_12101,N_12047);
and U12290 (N_12290,N_12053,N_12064);
nor U12291 (N_12291,N_12062,N_12070);
or U12292 (N_12292,N_12154,N_12010);
and U12293 (N_12293,N_12104,N_12029);
and U12294 (N_12294,N_12071,N_12105);
nor U12295 (N_12295,N_12090,N_12030);
nor U12296 (N_12296,N_12123,N_12070);
and U12297 (N_12297,N_12002,N_12043);
nor U12298 (N_12298,N_12071,N_12045);
nand U12299 (N_12299,N_12155,N_12073);
nor U12300 (N_12300,N_12049,N_12083);
nor U12301 (N_12301,N_12129,N_12062);
or U12302 (N_12302,N_12126,N_12014);
or U12303 (N_12303,N_12004,N_12001);
xor U12304 (N_12304,N_12156,N_12090);
or U12305 (N_12305,N_12056,N_12023);
nor U12306 (N_12306,N_12064,N_12010);
or U12307 (N_12307,N_12005,N_12157);
nand U12308 (N_12308,N_12060,N_12113);
or U12309 (N_12309,N_12028,N_12134);
nand U12310 (N_12310,N_12141,N_12106);
nand U12311 (N_12311,N_12117,N_12154);
xor U12312 (N_12312,N_12149,N_12017);
or U12313 (N_12313,N_12025,N_12122);
xor U12314 (N_12314,N_12102,N_12146);
or U12315 (N_12315,N_12144,N_12102);
nand U12316 (N_12316,N_12055,N_12047);
and U12317 (N_12317,N_12093,N_12070);
nand U12318 (N_12318,N_12067,N_12151);
xnor U12319 (N_12319,N_12051,N_12007);
or U12320 (N_12320,N_12182,N_12298);
nor U12321 (N_12321,N_12227,N_12264);
nor U12322 (N_12322,N_12190,N_12274);
nor U12323 (N_12323,N_12308,N_12186);
and U12324 (N_12324,N_12316,N_12241);
or U12325 (N_12325,N_12305,N_12251);
or U12326 (N_12326,N_12166,N_12300);
nand U12327 (N_12327,N_12319,N_12236);
xor U12328 (N_12328,N_12267,N_12215);
xnor U12329 (N_12329,N_12259,N_12185);
nor U12330 (N_12330,N_12205,N_12208);
nor U12331 (N_12331,N_12278,N_12169);
and U12332 (N_12332,N_12188,N_12244);
and U12333 (N_12333,N_12191,N_12230);
or U12334 (N_12334,N_12297,N_12223);
or U12335 (N_12335,N_12204,N_12282);
nor U12336 (N_12336,N_12195,N_12292);
nor U12337 (N_12337,N_12187,N_12285);
or U12338 (N_12338,N_12288,N_12279);
xor U12339 (N_12339,N_12162,N_12280);
and U12340 (N_12340,N_12229,N_12211);
or U12341 (N_12341,N_12167,N_12286);
xor U12342 (N_12342,N_12184,N_12299);
nand U12343 (N_12343,N_12224,N_12283);
nand U12344 (N_12344,N_12234,N_12265);
nor U12345 (N_12345,N_12249,N_12312);
xnor U12346 (N_12346,N_12216,N_12261);
or U12347 (N_12347,N_12172,N_12276);
or U12348 (N_12348,N_12318,N_12281);
nand U12349 (N_12349,N_12189,N_12257);
and U12350 (N_12350,N_12235,N_12161);
xor U12351 (N_12351,N_12201,N_12198);
or U12352 (N_12352,N_12262,N_12221);
nor U12353 (N_12353,N_12213,N_12217);
and U12354 (N_12354,N_12165,N_12302);
nor U12355 (N_12355,N_12199,N_12294);
and U12356 (N_12356,N_12232,N_12180);
and U12357 (N_12357,N_12266,N_12317);
nor U12358 (N_12358,N_12310,N_12219);
xor U12359 (N_12359,N_12228,N_12237);
nor U12360 (N_12360,N_12290,N_12209);
and U12361 (N_12361,N_12175,N_12193);
and U12362 (N_12362,N_12270,N_12203);
and U12363 (N_12363,N_12295,N_12311);
xnor U12364 (N_12364,N_12173,N_12178);
xnor U12365 (N_12365,N_12287,N_12194);
nand U12366 (N_12366,N_12246,N_12253);
or U12367 (N_12367,N_12170,N_12239);
nand U12368 (N_12368,N_12268,N_12163);
and U12369 (N_12369,N_12252,N_12260);
nand U12370 (N_12370,N_12207,N_12258);
xor U12371 (N_12371,N_12181,N_12256);
nor U12372 (N_12372,N_12171,N_12160);
nor U12373 (N_12373,N_12306,N_12197);
xor U12374 (N_12374,N_12164,N_12218);
nor U12375 (N_12375,N_12225,N_12248);
nor U12376 (N_12376,N_12233,N_12231);
nor U12377 (N_12377,N_12240,N_12247);
nand U12378 (N_12378,N_12168,N_12238);
or U12379 (N_12379,N_12314,N_12275);
and U12380 (N_12380,N_12200,N_12220);
or U12381 (N_12381,N_12250,N_12254);
or U12382 (N_12382,N_12289,N_12183);
nand U12383 (N_12383,N_12309,N_12303);
nor U12384 (N_12384,N_12304,N_12263);
or U12385 (N_12385,N_12315,N_12202);
xor U12386 (N_12386,N_12301,N_12313);
and U12387 (N_12387,N_12307,N_12214);
nand U12388 (N_12388,N_12222,N_12291);
or U12389 (N_12389,N_12192,N_12255);
xor U12390 (N_12390,N_12179,N_12277);
or U12391 (N_12391,N_12212,N_12210);
xnor U12392 (N_12392,N_12174,N_12273);
nand U12393 (N_12393,N_12242,N_12296);
or U12394 (N_12394,N_12243,N_12226);
nand U12395 (N_12395,N_12271,N_12272);
nor U12396 (N_12396,N_12196,N_12206);
and U12397 (N_12397,N_12284,N_12177);
nand U12398 (N_12398,N_12176,N_12245);
nor U12399 (N_12399,N_12293,N_12269);
nand U12400 (N_12400,N_12270,N_12214);
xor U12401 (N_12401,N_12197,N_12309);
nand U12402 (N_12402,N_12267,N_12271);
nor U12403 (N_12403,N_12225,N_12221);
nor U12404 (N_12404,N_12312,N_12307);
and U12405 (N_12405,N_12173,N_12282);
xor U12406 (N_12406,N_12293,N_12249);
and U12407 (N_12407,N_12260,N_12305);
nor U12408 (N_12408,N_12276,N_12261);
nor U12409 (N_12409,N_12310,N_12190);
nor U12410 (N_12410,N_12267,N_12227);
or U12411 (N_12411,N_12247,N_12292);
xnor U12412 (N_12412,N_12224,N_12252);
xor U12413 (N_12413,N_12191,N_12277);
nor U12414 (N_12414,N_12296,N_12258);
or U12415 (N_12415,N_12297,N_12225);
or U12416 (N_12416,N_12233,N_12299);
and U12417 (N_12417,N_12234,N_12232);
xnor U12418 (N_12418,N_12301,N_12276);
and U12419 (N_12419,N_12269,N_12242);
or U12420 (N_12420,N_12265,N_12171);
or U12421 (N_12421,N_12238,N_12316);
nand U12422 (N_12422,N_12243,N_12257);
or U12423 (N_12423,N_12247,N_12170);
nand U12424 (N_12424,N_12310,N_12168);
nor U12425 (N_12425,N_12221,N_12192);
xnor U12426 (N_12426,N_12197,N_12239);
nor U12427 (N_12427,N_12289,N_12207);
or U12428 (N_12428,N_12221,N_12239);
nor U12429 (N_12429,N_12208,N_12299);
and U12430 (N_12430,N_12230,N_12161);
nor U12431 (N_12431,N_12219,N_12193);
nor U12432 (N_12432,N_12177,N_12206);
xnor U12433 (N_12433,N_12258,N_12284);
or U12434 (N_12434,N_12271,N_12233);
and U12435 (N_12435,N_12171,N_12261);
nand U12436 (N_12436,N_12215,N_12318);
xnor U12437 (N_12437,N_12187,N_12170);
and U12438 (N_12438,N_12245,N_12297);
or U12439 (N_12439,N_12221,N_12189);
or U12440 (N_12440,N_12263,N_12253);
nor U12441 (N_12441,N_12228,N_12298);
and U12442 (N_12442,N_12270,N_12179);
xnor U12443 (N_12443,N_12280,N_12220);
and U12444 (N_12444,N_12313,N_12208);
and U12445 (N_12445,N_12275,N_12300);
xnor U12446 (N_12446,N_12172,N_12264);
xor U12447 (N_12447,N_12174,N_12276);
nand U12448 (N_12448,N_12265,N_12309);
or U12449 (N_12449,N_12249,N_12314);
or U12450 (N_12450,N_12306,N_12274);
nand U12451 (N_12451,N_12210,N_12205);
xnor U12452 (N_12452,N_12197,N_12245);
xor U12453 (N_12453,N_12169,N_12253);
or U12454 (N_12454,N_12208,N_12301);
and U12455 (N_12455,N_12192,N_12197);
nand U12456 (N_12456,N_12230,N_12222);
nor U12457 (N_12457,N_12318,N_12164);
nor U12458 (N_12458,N_12302,N_12266);
and U12459 (N_12459,N_12228,N_12299);
nand U12460 (N_12460,N_12189,N_12263);
or U12461 (N_12461,N_12270,N_12315);
and U12462 (N_12462,N_12254,N_12165);
xnor U12463 (N_12463,N_12168,N_12220);
xor U12464 (N_12464,N_12206,N_12197);
nand U12465 (N_12465,N_12235,N_12228);
nor U12466 (N_12466,N_12218,N_12227);
xor U12467 (N_12467,N_12282,N_12258);
or U12468 (N_12468,N_12219,N_12251);
and U12469 (N_12469,N_12315,N_12279);
xnor U12470 (N_12470,N_12168,N_12274);
nand U12471 (N_12471,N_12262,N_12242);
xor U12472 (N_12472,N_12180,N_12240);
nor U12473 (N_12473,N_12303,N_12194);
xnor U12474 (N_12474,N_12230,N_12177);
nor U12475 (N_12475,N_12281,N_12173);
or U12476 (N_12476,N_12185,N_12220);
or U12477 (N_12477,N_12260,N_12166);
xor U12478 (N_12478,N_12217,N_12283);
nor U12479 (N_12479,N_12259,N_12279);
and U12480 (N_12480,N_12460,N_12479);
and U12481 (N_12481,N_12360,N_12399);
nand U12482 (N_12482,N_12470,N_12427);
or U12483 (N_12483,N_12331,N_12372);
xnor U12484 (N_12484,N_12467,N_12448);
and U12485 (N_12485,N_12373,N_12377);
and U12486 (N_12486,N_12408,N_12346);
xnor U12487 (N_12487,N_12387,N_12330);
and U12488 (N_12488,N_12350,N_12418);
and U12489 (N_12489,N_12381,N_12347);
and U12490 (N_12490,N_12471,N_12345);
xnor U12491 (N_12491,N_12461,N_12378);
nor U12492 (N_12492,N_12341,N_12391);
and U12493 (N_12493,N_12478,N_12351);
xnor U12494 (N_12494,N_12375,N_12396);
and U12495 (N_12495,N_12338,N_12324);
nand U12496 (N_12496,N_12366,N_12328);
xor U12497 (N_12497,N_12322,N_12343);
nand U12498 (N_12498,N_12385,N_12365);
nor U12499 (N_12499,N_12443,N_12432);
xor U12500 (N_12500,N_12383,N_12397);
and U12501 (N_12501,N_12428,N_12363);
xor U12502 (N_12502,N_12336,N_12473);
and U12503 (N_12503,N_12401,N_12425);
nand U12504 (N_12504,N_12409,N_12386);
nor U12505 (N_12505,N_12453,N_12332);
nand U12506 (N_12506,N_12392,N_12416);
xnor U12507 (N_12507,N_12367,N_12413);
nand U12508 (N_12508,N_12433,N_12451);
xor U12509 (N_12509,N_12325,N_12415);
or U12510 (N_12510,N_12388,N_12394);
nor U12511 (N_12511,N_12362,N_12430);
nor U12512 (N_12512,N_12356,N_12339);
and U12513 (N_12513,N_12445,N_12431);
xnor U12514 (N_12514,N_12329,N_12402);
nand U12515 (N_12515,N_12442,N_12333);
or U12516 (N_12516,N_12390,N_12452);
nand U12517 (N_12517,N_12466,N_12454);
or U12518 (N_12518,N_12437,N_12417);
nand U12519 (N_12519,N_12406,N_12426);
and U12520 (N_12520,N_12374,N_12465);
nand U12521 (N_12521,N_12436,N_12334);
nand U12522 (N_12522,N_12327,N_12455);
or U12523 (N_12523,N_12477,N_12410);
or U12524 (N_12524,N_12352,N_12440);
xor U12525 (N_12525,N_12380,N_12355);
nor U12526 (N_12526,N_12419,N_12458);
nand U12527 (N_12527,N_12423,N_12361);
and U12528 (N_12528,N_12342,N_12472);
and U12529 (N_12529,N_12337,N_12435);
or U12530 (N_12530,N_12405,N_12393);
or U12531 (N_12531,N_12326,N_12463);
nand U12532 (N_12532,N_12434,N_12369);
xnor U12533 (N_12533,N_12450,N_12439);
xor U12534 (N_12534,N_12469,N_12447);
nor U12535 (N_12535,N_12359,N_12400);
nor U12536 (N_12536,N_12382,N_12323);
xor U12537 (N_12537,N_12404,N_12371);
xor U12538 (N_12538,N_12321,N_12420);
nand U12539 (N_12539,N_12348,N_12358);
or U12540 (N_12540,N_12357,N_12344);
nor U12541 (N_12541,N_12475,N_12414);
or U12542 (N_12542,N_12474,N_12468);
and U12543 (N_12543,N_12376,N_12389);
nand U12544 (N_12544,N_12449,N_12412);
nor U12545 (N_12545,N_12398,N_12441);
nor U12546 (N_12546,N_12403,N_12446);
or U12547 (N_12547,N_12411,N_12340);
nor U12548 (N_12548,N_12320,N_12459);
nand U12549 (N_12549,N_12407,N_12457);
xnor U12550 (N_12550,N_12422,N_12353);
and U12551 (N_12551,N_12438,N_12349);
and U12552 (N_12552,N_12395,N_12444);
nand U12553 (N_12553,N_12370,N_12424);
nor U12554 (N_12554,N_12379,N_12476);
nand U12555 (N_12555,N_12464,N_12456);
xnor U12556 (N_12556,N_12335,N_12368);
or U12557 (N_12557,N_12421,N_12462);
or U12558 (N_12558,N_12429,N_12384);
nand U12559 (N_12559,N_12364,N_12354);
and U12560 (N_12560,N_12425,N_12380);
and U12561 (N_12561,N_12416,N_12468);
nor U12562 (N_12562,N_12342,N_12423);
nand U12563 (N_12563,N_12414,N_12399);
xor U12564 (N_12564,N_12411,N_12321);
or U12565 (N_12565,N_12330,N_12333);
or U12566 (N_12566,N_12447,N_12434);
xor U12567 (N_12567,N_12423,N_12400);
nor U12568 (N_12568,N_12429,N_12364);
xnor U12569 (N_12569,N_12427,N_12478);
nand U12570 (N_12570,N_12413,N_12427);
and U12571 (N_12571,N_12326,N_12478);
nand U12572 (N_12572,N_12383,N_12421);
xnor U12573 (N_12573,N_12387,N_12350);
xor U12574 (N_12574,N_12422,N_12364);
and U12575 (N_12575,N_12341,N_12327);
xor U12576 (N_12576,N_12438,N_12442);
nor U12577 (N_12577,N_12380,N_12337);
and U12578 (N_12578,N_12411,N_12391);
nor U12579 (N_12579,N_12397,N_12417);
nor U12580 (N_12580,N_12422,N_12395);
nor U12581 (N_12581,N_12401,N_12426);
nand U12582 (N_12582,N_12396,N_12437);
nand U12583 (N_12583,N_12359,N_12416);
and U12584 (N_12584,N_12386,N_12451);
nor U12585 (N_12585,N_12401,N_12453);
nand U12586 (N_12586,N_12326,N_12444);
and U12587 (N_12587,N_12417,N_12459);
nor U12588 (N_12588,N_12412,N_12399);
xor U12589 (N_12589,N_12444,N_12386);
xnor U12590 (N_12590,N_12434,N_12420);
xnor U12591 (N_12591,N_12324,N_12415);
or U12592 (N_12592,N_12355,N_12341);
nor U12593 (N_12593,N_12442,N_12458);
or U12594 (N_12594,N_12347,N_12447);
and U12595 (N_12595,N_12473,N_12413);
xor U12596 (N_12596,N_12421,N_12362);
and U12597 (N_12597,N_12465,N_12421);
and U12598 (N_12598,N_12340,N_12354);
nor U12599 (N_12599,N_12381,N_12478);
and U12600 (N_12600,N_12390,N_12440);
and U12601 (N_12601,N_12343,N_12441);
or U12602 (N_12602,N_12462,N_12445);
nor U12603 (N_12603,N_12342,N_12332);
nand U12604 (N_12604,N_12358,N_12350);
nor U12605 (N_12605,N_12344,N_12326);
nand U12606 (N_12606,N_12404,N_12337);
or U12607 (N_12607,N_12386,N_12392);
xor U12608 (N_12608,N_12479,N_12340);
xor U12609 (N_12609,N_12471,N_12320);
nor U12610 (N_12610,N_12337,N_12345);
xor U12611 (N_12611,N_12402,N_12396);
xnor U12612 (N_12612,N_12406,N_12366);
nand U12613 (N_12613,N_12344,N_12466);
or U12614 (N_12614,N_12334,N_12465);
and U12615 (N_12615,N_12396,N_12466);
and U12616 (N_12616,N_12397,N_12443);
nor U12617 (N_12617,N_12395,N_12417);
xor U12618 (N_12618,N_12335,N_12457);
xor U12619 (N_12619,N_12347,N_12378);
or U12620 (N_12620,N_12321,N_12478);
and U12621 (N_12621,N_12459,N_12440);
nor U12622 (N_12622,N_12358,N_12412);
and U12623 (N_12623,N_12459,N_12341);
and U12624 (N_12624,N_12355,N_12333);
or U12625 (N_12625,N_12336,N_12334);
and U12626 (N_12626,N_12348,N_12440);
or U12627 (N_12627,N_12363,N_12375);
or U12628 (N_12628,N_12440,N_12410);
nand U12629 (N_12629,N_12453,N_12477);
nand U12630 (N_12630,N_12357,N_12371);
nand U12631 (N_12631,N_12456,N_12390);
xor U12632 (N_12632,N_12327,N_12389);
nand U12633 (N_12633,N_12335,N_12343);
nand U12634 (N_12634,N_12467,N_12469);
and U12635 (N_12635,N_12349,N_12442);
nor U12636 (N_12636,N_12380,N_12404);
nand U12637 (N_12637,N_12323,N_12335);
xnor U12638 (N_12638,N_12340,N_12390);
and U12639 (N_12639,N_12425,N_12446);
and U12640 (N_12640,N_12541,N_12487);
nand U12641 (N_12641,N_12573,N_12593);
nand U12642 (N_12642,N_12635,N_12583);
or U12643 (N_12643,N_12568,N_12588);
nand U12644 (N_12644,N_12491,N_12632);
and U12645 (N_12645,N_12601,N_12544);
nand U12646 (N_12646,N_12562,N_12598);
nor U12647 (N_12647,N_12516,N_12580);
or U12648 (N_12648,N_12550,N_12513);
and U12649 (N_12649,N_12579,N_12483);
and U12650 (N_12650,N_12484,N_12631);
or U12651 (N_12651,N_12636,N_12595);
or U12652 (N_12652,N_12522,N_12524);
nor U12653 (N_12653,N_12608,N_12553);
nand U12654 (N_12654,N_12480,N_12528);
or U12655 (N_12655,N_12489,N_12607);
nor U12656 (N_12656,N_12603,N_12597);
or U12657 (N_12657,N_12546,N_12574);
nor U12658 (N_12658,N_12566,N_12545);
nor U12659 (N_12659,N_12616,N_12493);
and U12660 (N_12660,N_12497,N_12509);
nor U12661 (N_12661,N_12514,N_12496);
or U12662 (N_12662,N_12581,N_12515);
or U12663 (N_12663,N_12628,N_12532);
or U12664 (N_12664,N_12611,N_12561);
xor U12665 (N_12665,N_12547,N_12525);
nand U12666 (N_12666,N_12582,N_12506);
nand U12667 (N_12667,N_12576,N_12610);
or U12668 (N_12668,N_12594,N_12508);
and U12669 (N_12669,N_12572,N_12626);
xnor U12670 (N_12670,N_12485,N_12565);
nor U12671 (N_12671,N_12502,N_12575);
or U12672 (N_12672,N_12555,N_12585);
nor U12673 (N_12673,N_12490,N_12578);
or U12674 (N_12674,N_12557,N_12512);
xnor U12675 (N_12675,N_12517,N_12596);
xnor U12676 (N_12676,N_12634,N_12589);
nand U12677 (N_12677,N_12494,N_12498);
or U12678 (N_12678,N_12543,N_12570);
xnor U12679 (N_12679,N_12519,N_12518);
or U12680 (N_12680,N_12501,N_12542);
or U12681 (N_12681,N_12529,N_12560);
nor U12682 (N_12682,N_12551,N_12619);
nor U12683 (N_12683,N_12540,N_12600);
nand U12684 (N_12684,N_12624,N_12630);
and U12685 (N_12685,N_12638,N_12536);
xor U12686 (N_12686,N_12621,N_12613);
nand U12687 (N_12687,N_12505,N_12590);
xnor U12688 (N_12688,N_12526,N_12627);
xor U12689 (N_12689,N_12606,N_12510);
or U12690 (N_12690,N_12495,N_12612);
nor U12691 (N_12691,N_12617,N_12567);
and U12692 (N_12692,N_12556,N_12486);
nand U12693 (N_12693,N_12520,N_12569);
and U12694 (N_12694,N_12587,N_12559);
nor U12695 (N_12695,N_12623,N_12535);
nor U12696 (N_12696,N_12622,N_12488);
or U12697 (N_12697,N_12615,N_12527);
or U12698 (N_12698,N_12523,N_12625);
or U12699 (N_12699,N_12577,N_12591);
or U12700 (N_12700,N_12500,N_12637);
or U12701 (N_12701,N_12618,N_12602);
nor U12702 (N_12702,N_12620,N_12492);
nor U12703 (N_12703,N_12592,N_12629);
nor U12704 (N_12704,N_12503,N_12564);
nand U12705 (N_12705,N_12534,N_12614);
xnor U12706 (N_12706,N_12548,N_12531);
nor U12707 (N_12707,N_12539,N_12558);
nand U12708 (N_12708,N_12571,N_12538);
nor U12709 (N_12709,N_12586,N_12507);
xnor U12710 (N_12710,N_12563,N_12499);
nor U12711 (N_12711,N_12584,N_12504);
or U12712 (N_12712,N_12549,N_12554);
or U12713 (N_12713,N_12605,N_12537);
nand U12714 (N_12714,N_12604,N_12639);
nand U12715 (N_12715,N_12511,N_12533);
or U12716 (N_12716,N_12530,N_12599);
nand U12717 (N_12717,N_12633,N_12521);
xor U12718 (N_12718,N_12481,N_12609);
and U12719 (N_12719,N_12552,N_12482);
xnor U12720 (N_12720,N_12636,N_12614);
nand U12721 (N_12721,N_12580,N_12592);
or U12722 (N_12722,N_12584,N_12578);
xor U12723 (N_12723,N_12484,N_12500);
nand U12724 (N_12724,N_12558,N_12497);
xor U12725 (N_12725,N_12583,N_12577);
nand U12726 (N_12726,N_12528,N_12576);
xor U12727 (N_12727,N_12625,N_12638);
or U12728 (N_12728,N_12518,N_12532);
nand U12729 (N_12729,N_12590,N_12604);
or U12730 (N_12730,N_12591,N_12639);
nor U12731 (N_12731,N_12524,N_12482);
xor U12732 (N_12732,N_12603,N_12627);
nor U12733 (N_12733,N_12636,N_12533);
xnor U12734 (N_12734,N_12610,N_12557);
nor U12735 (N_12735,N_12617,N_12615);
nor U12736 (N_12736,N_12634,N_12596);
nand U12737 (N_12737,N_12489,N_12619);
and U12738 (N_12738,N_12492,N_12609);
nor U12739 (N_12739,N_12611,N_12593);
or U12740 (N_12740,N_12560,N_12566);
xnor U12741 (N_12741,N_12618,N_12539);
nor U12742 (N_12742,N_12606,N_12632);
xnor U12743 (N_12743,N_12634,N_12496);
nand U12744 (N_12744,N_12624,N_12594);
and U12745 (N_12745,N_12490,N_12548);
or U12746 (N_12746,N_12531,N_12490);
nor U12747 (N_12747,N_12618,N_12568);
nand U12748 (N_12748,N_12519,N_12605);
and U12749 (N_12749,N_12523,N_12593);
nand U12750 (N_12750,N_12625,N_12627);
nor U12751 (N_12751,N_12606,N_12590);
and U12752 (N_12752,N_12630,N_12563);
nand U12753 (N_12753,N_12558,N_12639);
xnor U12754 (N_12754,N_12498,N_12540);
nor U12755 (N_12755,N_12503,N_12481);
and U12756 (N_12756,N_12482,N_12506);
and U12757 (N_12757,N_12633,N_12491);
xnor U12758 (N_12758,N_12617,N_12630);
xnor U12759 (N_12759,N_12593,N_12615);
and U12760 (N_12760,N_12633,N_12539);
nor U12761 (N_12761,N_12488,N_12506);
and U12762 (N_12762,N_12587,N_12588);
nor U12763 (N_12763,N_12605,N_12544);
and U12764 (N_12764,N_12622,N_12543);
nand U12765 (N_12765,N_12563,N_12600);
or U12766 (N_12766,N_12572,N_12588);
or U12767 (N_12767,N_12584,N_12609);
and U12768 (N_12768,N_12480,N_12529);
or U12769 (N_12769,N_12550,N_12607);
nor U12770 (N_12770,N_12488,N_12632);
and U12771 (N_12771,N_12500,N_12591);
or U12772 (N_12772,N_12514,N_12598);
nand U12773 (N_12773,N_12517,N_12621);
nand U12774 (N_12774,N_12601,N_12499);
nand U12775 (N_12775,N_12636,N_12546);
nand U12776 (N_12776,N_12530,N_12512);
or U12777 (N_12777,N_12607,N_12570);
and U12778 (N_12778,N_12619,N_12485);
nand U12779 (N_12779,N_12582,N_12550);
nor U12780 (N_12780,N_12624,N_12623);
or U12781 (N_12781,N_12496,N_12511);
nor U12782 (N_12782,N_12570,N_12550);
or U12783 (N_12783,N_12571,N_12555);
nor U12784 (N_12784,N_12486,N_12544);
and U12785 (N_12785,N_12625,N_12521);
nand U12786 (N_12786,N_12531,N_12610);
or U12787 (N_12787,N_12504,N_12606);
or U12788 (N_12788,N_12520,N_12553);
nor U12789 (N_12789,N_12612,N_12555);
xnor U12790 (N_12790,N_12561,N_12515);
and U12791 (N_12791,N_12637,N_12598);
nand U12792 (N_12792,N_12511,N_12552);
and U12793 (N_12793,N_12556,N_12580);
or U12794 (N_12794,N_12615,N_12565);
xnor U12795 (N_12795,N_12613,N_12570);
xnor U12796 (N_12796,N_12521,N_12612);
nor U12797 (N_12797,N_12498,N_12566);
nand U12798 (N_12798,N_12527,N_12505);
nand U12799 (N_12799,N_12585,N_12605);
or U12800 (N_12800,N_12713,N_12657);
nand U12801 (N_12801,N_12654,N_12741);
and U12802 (N_12802,N_12663,N_12708);
xnor U12803 (N_12803,N_12715,N_12707);
xor U12804 (N_12804,N_12673,N_12648);
nand U12805 (N_12805,N_12796,N_12752);
nand U12806 (N_12806,N_12795,N_12729);
and U12807 (N_12807,N_12798,N_12678);
nand U12808 (N_12808,N_12655,N_12700);
nand U12809 (N_12809,N_12656,N_12722);
nand U12810 (N_12810,N_12701,N_12792);
xnor U12811 (N_12811,N_12664,N_12688);
xor U12812 (N_12812,N_12661,N_12647);
or U12813 (N_12813,N_12706,N_12751);
nand U12814 (N_12814,N_12774,N_12649);
xor U12815 (N_12815,N_12763,N_12651);
and U12816 (N_12816,N_12784,N_12702);
and U12817 (N_12817,N_12735,N_12775);
xor U12818 (N_12818,N_12726,N_12720);
and U12819 (N_12819,N_12643,N_12666);
nand U12820 (N_12820,N_12744,N_12732);
nand U12821 (N_12821,N_12731,N_12717);
and U12822 (N_12822,N_12768,N_12780);
nand U12823 (N_12823,N_12671,N_12723);
or U12824 (N_12824,N_12642,N_12681);
and U12825 (N_12825,N_12736,N_12719);
nand U12826 (N_12826,N_12690,N_12640);
or U12827 (N_12827,N_12788,N_12765);
xor U12828 (N_12828,N_12756,N_12769);
nand U12829 (N_12829,N_12710,N_12703);
nand U12830 (N_12830,N_12746,N_12753);
xnor U12831 (N_12831,N_12645,N_12691);
and U12832 (N_12832,N_12770,N_12740);
nor U12833 (N_12833,N_12658,N_12725);
nand U12834 (N_12834,N_12669,N_12737);
nand U12835 (N_12835,N_12714,N_12758);
nand U12836 (N_12836,N_12660,N_12653);
nor U12837 (N_12837,N_12705,N_12683);
or U12838 (N_12838,N_12682,N_12668);
or U12839 (N_12839,N_12783,N_12692);
and U12840 (N_12840,N_12716,N_12687);
nand U12841 (N_12841,N_12799,N_12665);
or U12842 (N_12842,N_12761,N_12779);
nor U12843 (N_12843,N_12733,N_12730);
or U12844 (N_12844,N_12662,N_12644);
or U12845 (N_12845,N_12759,N_12787);
and U12846 (N_12846,N_12650,N_12772);
nor U12847 (N_12847,N_12641,N_12771);
nand U12848 (N_12848,N_12694,N_12652);
or U12849 (N_12849,N_12724,N_12785);
xor U12850 (N_12850,N_12699,N_12711);
xor U12851 (N_12851,N_12762,N_12738);
or U12852 (N_12852,N_12667,N_12760);
nand U12853 (N_12853,N_12739,N_12755);
nor U12854 (N_12854,N_12646,N_12698);
and U12855 (N_12855,N_12743,N_12749);
xnor U12856 (N_12856,N_12742,N_12686);
and U12857 (N_12857,N_12689,N_12748);
xor U12858 (N_12858,N_12672,N_12728);
nor U12859 (N_12859,N_12790,N_12777);
or U12860 (N_12860,N_12764,N_12794);
xor U12861 (N_12861,N_12696,N_12679);
and U12862 (N_12862,N_12766,N_12754);
or U12863 (N_12863,N_12695,N_12791);
nor U12864 (N_12864,N_12676,N_12734);
xor U12865 (N_12865,N_12685,N_12789);
nand U12866 (N_12866,N_12778,N_12727);
nor U12867 (N_12867,N_12793,N_12712);
nor U12868 (N_12868,N_12781,N_12674);
or U12869 (N_12869,N_12786,N_12709);
nand U12870 (N_12870,N_12670,N_12721);
nand U12871 (N_12871,N_12776,N_12747);
nor U12872 (N_12872,N_12767,N_12782);
nand U12873 (N_12873,N_12659,N_12680);
nand U12874 (N_12874,N_12684,N_12697);
xor U12875 (N_12875,N_12675,N_12773);
and U12876 (N_12876,N_12797,N_12693);
nor U12877 (N_12877,N_12745,N_12718);
nor U12878 (N_12878,N_12757,N_12704);
or U12879 (N_12879,N_12677,N_12750);
nor U12880 (N_12880,N_12733,N_12736);
or U12881 (N_12881,N_12710,N_12657);
nand U12882 (N_12882,N_12779,N_12697);
nand U12883 (N_12883,N_12669,N_12709);
xnor U12884 (N_12884,N_12671,N_12779);
xnor U12885 (N_12885,N_12714,N_12654);
nand U12886 (N_12886,N_12776,N_12733);
and U12887 (N_12887,N_12781,N_12773);
nand U12888 (N_12888,N_12723,N_12688);
nor U12889 (N_12889,N_12653,N_12686);
nand U12890 (N_12890,N_12741,N_12678);
or U12891 (N_12891,N_12778,N_12662);
xor U12892 (N_12892,N_12720,N_12715);
xor U12893 (N_12893,N_12726,N_12754);
nor U12894 (N_12894,N_12726,N_12735);
or U12895 (N_12895,N_12665,N_12789);
nand U12896 (N_12896,N_12715,N_12760);
and U12897 (N_12897,N_12649,N_12692);
nand U12898 (N_12898,N_12714,N_12736);
and U12899 (N_12899,N_12764,N_12781);
or U12900 (N_12900,N_12756,N_12761);
or U12901 (N_12901,N_12796,N_12656);
nor U12902 (N_12902,N_12648,N_12678);
or U12903 (N_12903,N_12784,N_12751);
nand U12904 (N_12904,N_12727,N_12730);
xor U12905 (N_12905,N_12657,N_12733);
xnor U12906 (N_12906,N_12796,N_12758);
and U12907 (N_12907,N_12697,N_12790);
nor U12908 (N_12908,N_12740,N_12687);
or U12909 (N_12909,N_12705,N_12782);
nand U12910 (N_12910,N_12756,N_12678);
and U12911 (N_12911,N_12756,N_12725);
nand U12912 (N_12912,N_12732,N_12749);
nor U12913 (N_12913,N_12781,N_12669);
or U12914 (N_12914,N_12681,N_12781);
or U12915 (N_12915,N_12665,N_12705);
and U12916 (N_12916,N_12640,N_12701);
nor U12917 (N_12917,N_12755,N_12673);
or U12918 (N_12918,N_12724,N_12735);
nor U12919 (N_12919,N_12670,N_12667);
nand U12920 (N_12920,N_12778,N_12725);
or U12921 (N_12921,N_12739,N_12703);
or U12922 (N_12922,N_12709,N_12702);
nand U12923 (N_12923,N_12774,N_12685);
or U12924 (N_12924,N_12741,N_12656);
xnor U12925 (N_12925,N_12745,N_12751);
nor U12926 (N_12926,N_12770,N_12675);
nor U12927 (N_12927,N_12673,N_12740);
nor U12928 (N_12928,N_12771,N_12736);
nor U12929 (N_12929,N_12762,N_12687);
or U12930 (N_12930,N_12755,N_12652);
nor U12931 (N_12931,N_12788,N_12661);
nor U12932 (N_12932,N_12716,N_12780);
xor U12933 (N_12933,N_12748,N_12691);
xor U12934 (N_12934,N_12780,N_12692);
xnor U12935 (N_12935,N_12730,N_12729);
xnor U12936 (N_12936,N_12798,N_12694);
nand U12937 (N_12937,N_12742,N_12729);
nand U12938 (N_12938,N_12798,N_12781);
nor U12939 (N_12939,N_12664,N_12713);
nand U12940 (N_12940,N_12763,N_12758);
and U12941 (N_12941,N_12764,N_12663);
or U12942 (N_12942,N_12648,N_12706);
and U12943 (N_12943,N_12736,N_12789);
or U12944 (N_12944,N_12667,N_12714);
nor U12945 (N_12945,N_12651,N_12640);
xor U12946 (N_12946,N_12692,N_12768);
nor U12947 (N_12947,N_12703,N_12760);
or U12948 (N_12948,N_12692,N_12708);
nand U12949 (N_12949,N_12725,N_12797);
nand U12950 (N_12950,N_12763,N_12769);
nand U12951 (N_12951,N_12774,N_12741);
or U12952 (N_12952,N_12771,N_12755);
nand U12953 (N_12953,N_12691,N_12673);
xnor U12954 (N_12954,N_12797,N_12679);
and U12955 (N_12955,N_12668,N_12694);
and U12956 (N_12956,N_12661,N_12663);
xor U12957 (N_12957,N_12755,N_12778);
xnor U12958 (N_12958,N_12798,N_12746);
nor U12959 (N_12959,N_12758,N_12785);
or U12960 (N_12960,N_12883,N_12842);
and U12961 (N_12961,N_12932,N_12894);
nand U12962 (N_12962,N_12875,N_12936);
xor U12963 (N_12963,N_12893,N_12857);
and U12964 (N_12964,N_12854,N_12814);
xor U12965 (N_12965,N_12810,N_12909);
nor U12966 (N_12966,N_12855,N_12874);
and U12967 (N_12967,N_12844,N_12885);
xor U12968 (N_12968,N_12907,N_12811);
and U12969 (N_12969,N_12869,N_12902);
xnor U12970 (N_12970,N_12850,N_12879);
nand U12971 (N_12971,N_12940,N_12953);
and U12972 (N_12972,N_12878,N_12821);
and U12973 (N_12973,N_12897,N_12950);
nor U12974 (N_12974,N_12937,N_12840);
xor U12975 (N_12975,N_12828,N_12852);
xor U12976 (N_12976,N_12918,N_12867);
xor U12977 (N_12977,N_12815,N_12862);
xnor U12978 (N_12978,N_12957,N_12880);
nand U12979 (N_12979,N_12818,N_12866);
and U12980 (N_12980,N_12845,N_12823);
and U12981 (N_12981,N_12830,N_12933);
or U12982 (N_12982,N_12832,N_12872);
and U12983 (N_12983,N_12876,N_12889);
nand U12984 (N_12984,N_12915,N_12824);
and U12985 (N_12985,N_12834,N_12816);
xnor U12986 (N_12986,N_12849,N_12943);
and U12987 (N_12987,N_12836,N_12853);
and U12988 (N_12988,N_12809,N_12805);
nand U12989 (N_12989,N_12813,N_12922);
nand U12990 (N_12990,N_12861,N_12921);
or U12991 (N_12991,N_12947,N_12860);
nand U12992 (N_12992,N_12892,N_12865);
nand U12993 (N_12993,N_12864,N_12939);
nand U12994 (N_12994,N_12919,N_12858);
nand U12995 (N_12995,N_12917,N_12835);
and U12996 (N_12996,N_12884,N_12911);
or U12997 (N_12997,N_12946,N_12873);
or U12998 (N_12998,N_12800,N_12806);
nor U12999 (N_12999,N_12941,N_12890);
xnor U13000 (N_13000,N_12820,N_12929);
nor U13001 (N_13001,N_12931,N_12901);
nor U13002 (N_13002,N_12863,N_12877);
xnor U13003 (N_13003,N_12831,N_12944);
or U13004 (N_13004,N_12881,N_12851);
nand U13005 (N_13005,N_12895,N_12908);
or U13006 (N_13006,N_12801,N_12930);
nor U13007 (N_13007,N_12942,N_12868);
or U13008 (N_13008,N_12959,N_12938);
nand U13009 (N_13009,N_12920,N_12804);
nor U13010 (N_13010,N_12887,N_12948);
xnor U13011 (N_13011,N_12954,N_12934);
nand U13012 (N_13012,N_12871,N_12927);
nor U13013 (N_13013,N_12945,N_12952);
nor U13014 (N_13014,N_12825,N_12949);
nand U13015 (N_13015,N_12841,N_12838);
xnor U13016 (N_13016,N_12827,N_12808);
or U13017 (N_13017,N_12856,N_12839);
and U13018 (N_13018,N_12846,N_12903);
nand U13019 (N_13019,N_12912,N_12822);
xor U13020 (N_13020,N_12848,N_12928);
or U13021 (N_13021,N_12896,N_12870);
xnor U13022 (N_13022,N_12925,N_12833);
or U13023 (N_13023,N_12905,N_12900);
xnor U13024 (N_13024,N_12847,N_12956);
xnor U13025 (N_13025,N_12888,N_12882);
or U13026 (N_13026,N_12904,N_12899);
or U13027 (N_13027,N_12914,N_12886);
nand U13028 (N_13028,N_12913,N_12819);
nand U13029 (N_13029,N_12916,N_12803);
xor U13030 (N_13030,N_12935,N_12829);
nand U13031 (N_13031,N_12923,N_12802);
xor U13032 (N_13032,N_12926,N_12898);
nand U13033 (N_13033,N_12812,N_12891);
or U13034 (N_13034,N_12859,N_12843);
xnor U13035 (N_13035,N_12807,N_12951);
nand U13036 (N_13036,N_12817,N_12906);
nand U13037 (N_13037,N_12924,N_12958);
nor U13038 (N_13038,N_12910,N_12826);
nor U13039 (N_13039,N_12955,N_12837);
or U13040 (N_13040,N_12919,N_12879);
xor U13041 (N_13041,N_12863,N_12917);
xor U13042 (N_13042,N_12876,N_12881);
xor U13043 (N_13043,N_12896,N_12958);
nand U13044 (N_13044,N_12901,N_12941);
or U13045 (N_13045,N_12859,N_12876);
xor U13046 (N_13046,N_12802,N_12800);
nand U13047 (N_13047,N_12901,N_12801);
and U13048 (N_13048,N_12865,N_12931);
nor U13049 (N_13049,N_12928,N_12882);
nand U13050 (N_13050,N_12881,N_12869);
and U13051 (N_13051,N_12891,N_12840);
xnor U13052 (N_13052,N_12819,N_12936);
nor U13053 (N_13053,N_12901,N_12836);
or U13054 (N_13054,N_12894,N_12852);
xnor U13055 (N_13055,N_12920,N_12936);
and U13056 (N_13056,N_12949,N_12912);
or U13057 (N_13057,N_12875,N_12823);
or U13058 (N_13058,N_12922,N_12866);
or U13059 (N_13059,N_12823,N_12830);
and U13060 (N_13060,N_12865,N_12810);
and U13061 (N_13061,N_12859,N_12902);
or U13062 (N_13062,N_12958,N_12861);
and U13063 (N_13063,N_12835,N_12890);
nand U13064 (N_13064,N_12862,N_12846);
and U13065 (N_13065,N_12945,N_12810);
or U13066 (N_13066,N_12841,N_12800);
nand U13067 (N_13067,N_12859,N_12885);
or U13068 (N_13068,N_12894,N_12886);
or U13069 (N_13069,N_12841,N_12833);
and U13070 (N_13070,N_12932,N_12947);
and U13071 (N_13071,N_12834,N_12926);
and U13072 (N_13072,N_12825,N_12809);
nand U13073 (N_13073,N_12885,N_12910);
xor U13074 (N_13074,N_12814,N_12954);
and U13075 (N_13075,N_12936,N_12854);
or U13076 (N_13076,N_12876,N_12807);
and U13077 (N_13077,N_12831,N_12826);
and U13078 (N_13078,N_12923,N_12871);
xor U13079 (N_13079,N_12814,N_12827);
xnor U13080 (N_13080,N_12957,N_12913);
and U13081 (N_13081,N_12889,N_12865);
nor U13082 (N_13082,N_12949,N_12837);
nor U13083 (N_13083,N_12830,N_12833);
and U13084 (N_13084,N_12895,N_12927);
or U13085 (N_13085,N_12909,N_12922);
or U13086 (N_13086,N_12853,N_12948);
xnor U13087 (N_13087,N_12885,N_12935);
and U13088 (N_13088,N_12875,N_12932);
and U13089 (N_13089,N_12849,N_12856);
and U13090 (N_13090,N_12956,N_12813);
nand U13091 (N_13091,N_12883,N_12942);
or U13092 (N_13092,N_12909,N_12842);
nor U13093 (N_13093,N_12806,N_12945);
and U13094 (N_13094,N_12886,N_12809);
and U13095 (N_13095,N_12851,N_12876);
and U13096 (N_13096,N_12910,N_12814);
nor U13097 (N_13097,N_12902,N_12809);
nor U13098 (N_13098,N_12956,N_12822);
and U13099 (N_13099,N_12931,N_12839);
xnor U13100 (N_13100,N_12948,N_12890);
nand U13101 (N_13101,N_12910,N_12876);
nor U13102 (N_13102,N_12831,N_12837);
nor U13103 (N_13103,N_12895,N_12910);
nor U13104 (N_13104,N_12828,N_12873);
or U13105 (N_13105,N_12920,N_12932);
or U13106 (N_13106,N_12872,N_12824);
nor U13107 (N_13107,N_12811,N_12824);
or U13108 (N_13108,N_12837,N_12817);
xor U13109 (N_13109,N_12947,N_12885);
xnor U13110 (N_13110,N_12850,N_12868);
and U13111 (N_13111,N_12890,N_12806);
and U13112 (N_13112,N_12882,N_12895);
xor U13113 (N_13113,N_12902,N_12931);
nand U13114 (N_13114,N_12949,N_12817);
xor U13115 (N_13115,N_12920,N_12843);
xor U13116 (N_13116,N_12897,N_12941);
and U13117 (N_13117,N_12851,N_12803);
and U13118 (N_13118,N_12859,N_12852);
nor U13119 (N_13119,N_12860,N_12917);
nand U13120 (N_13120,N_13050,N_13105);
xnor U13121 (N_13121,N_13043,N_13052);
xnor U13122 (N_13122,N_13030,N_13077);
nor U13123 (N_13123,N_13051,N_13085);
nor U13124 (N_13124,N_13060,N_13112);
nand U13125 (N_13125,N_13019,N_13041);
and U13126 (N_13126,N_13028,N_12972);
and U13127 (N_13127,N_12970,N_13038);
xor U13128 (N_13128,N_13114,N_13118);
or U13129 (N_13129,N_13040,N_13097);
and U13130 (N_13130,N_13109,N_13018);
and U13131 (N_13131,N_12986,N_13042);
or U13132 (N_13132,N_12989,N_13011);
xnor U13133 (N_13133,N_13070,N_13088);
nor U13134 (N_13134,N_13069,N_13061);
nand U13135 (N_13135,N_13101,N_13017);
or U13136 (N_13136,N_12964,N_13044);
and U13137 (N_13137,N_12990,N_13004);
nor U13138 (N_13138,N_13053,N_12965);
or U13139 (N_13139,N_13020,N_13115);
nor U13140 (N_13140,N_13031,N_13036);
nand U13141 (N_13141,N_12981,N_13087);
nor U13142 (N_13142,N_12963,N_12967);
or U13143 (N_13143,N_12962,N_13015);
xnor U13144 (N_13144,N_13078,N_13048);
nand U13145 (N_13145,N_13116,N_12975);
or U13146 (N_13146,N_13055,N_13063);
xor U13147 (N_13147,N_13056,N_13094);
xor U13148 (N_13148,N_12994,N_13079);
nand U13149 (N_13149,N_13065,N_13033);
and U13150 (N_13150,N_13026,N_13027);
xor U13151 (N_13151,N_13023,N_12966);
xor U13152 (N_13152,N_12968,N_13025);
or U13153 (N_13153,N_12977,N_13107);
or U13154 (N_13154,N_13119,N_13099);
nor U13155 (N_13155,N_12991,N_13104);
xor U13156 (N_13156,N_13001,N_12998);
and U13157 (N_13157,N_13012,N_13083);
and U13158 (N_13158,N_13059,N_13074);
and U13159 (N_13159,N_13013,N_13005);
xor U13160 (N_13160,N_12996,N_13096);
nand U13161 (N_13161,N_13000,N_13103);
nor U13162 (N_13162,N_12974,N_12983);
nand U13163 (N_13163,N_13071,N_13003);
and U13164 (N_13164,N_12984,N_13067);
xnor U13165 (N_13165,N_13076,N_13022);
nor U13166 (N_13166,N_13080,N_12969);
and U13167 (N_13167,N_13024,N_13032);
nand U13168 (N_13168,N_13081,N_13106);
xor U13169 (N_13169,N_12978,N_13095);
nor U13170 (N_13170,N_12995,N_13089);
nand U13171 (N_13171,N_13113,N_12961);
and U13172 (N_13172,N_12960,N_12979);
or U13173 (N_13173,N_13062,N_13035);
nor U13174 (N_13174,N_13084,N_12993);
nand U13175 (N_13175,N_13047,N_12971);
xnor U13176 (N_13176,N_13093,N_12980);
or U13177 (N_13177,N_13086,N_13098);
nand U13178 (N_13178,N_13064,N_12997);
xor U13179 (N_13179,N_13037,N_13068);
xor U13180 (N_13180,N_13039,N_13045);
nor U13181 (N_13181,N_13082,N_13029);
nor U13182 (N_13182,N_13057,N_13016);
nor U13183 (N_13183,N_13006,N_13049);
or U13184 (N_13184,N_13090,N_12987);
xnor U13185 (N_13185,N_12973,N_13108);
nand U13186 (N_13186,N_13073,N_13100);
and U13187 (N_13187,N_13102,N_13021);
and U13188 (N_13188,N_13117,N_13007);
nand U13189 (N_13189,N_13046,N_13054);
and U13190 (N_13190,N_12976,N_13008);
xnor U13191 (N_13191,N_12982,N_13091);
xor U13192 (N_13192,N_13058,N_12985);
nand U13193 (N_13193,N_13010,N_13014);
nand U13194 (N_13194,N_13034,N_12988);
xor U13195 (N_13195,N_13002,N_13092);
nor U13196 (N_13196,N_12992,N_13075);
nand U13197 (N_13197,N_13009,N_13072);
and U13198 (N_13198,N_13110,N_12999);
nor U13199 (N_13199,N_13111,N_13066);
xnor U13200 (N_13200,N_13015,N_13065);
or U13201 (N_13201,N_13106,N_12986);
and U13202 (N_13202,N_12975,N_13022);
or U13203 (N_13203,N_12962,N_13002);
and U13204 (N_13204,N_13027,N_12970);
or U13205 (N_13205,N_13093,N_13057);
nand U13206 (N_13206,N_13070,N_13055);
xor U13207 (N_13207,N_12983,N_13094);
and U13208 (N_13208,N_13073,N_13103);
nand U13209 (N_13209,N_12967,N_13076);
and U13210 (N_13210,N_12998,N_12989);
nor U13211 (N_13211,N_13041,N_13000);
nor U13212 (N_13212,N_12995,N_12963);
xnor U13213 (N_13213,N_13109,N_13062);
xnor U13214 (N_13214,N_13022,N_13003);
and U13215 (N_13215,N_13109,N_13045);
xnor U13216 (N_13216,N_13113,N_12993);
nor U13217 (N_13217,N_13102,N_13022);
and U13218 (N_13218,N_13010,N_13051);
and U13219 (N_13219,N_12969,N_13094);
nor U13220 (N_13220,N_13107,N_13064);
nand U13221 (N_13221,N_13040,N_12981);
nor U13222 (N_13222,N_13054,N_13103);
and U13223 (N_13223,N_12986,N_13054);
xor U13224 (N_13224,N_13019,N_13023);
nand U13225 (N_13225,N_13030,N_13078);
nor U13226 (N_13226,N_12987,N_13067);
nor U13227 (N_13227,N_13111,N_13070);
or U13228 (N_13228,N_12989,N_13091);
and U13229 (N_13229,N_13031,N_12966);
xor U13230 (N_13230,N_13004,N_13043);
and U13231 (N_13231,N_13089,N_13064);
nand U13232 (N_13232,N_13024,N_13086);
nand U13233 (N_13233,N_13056,N_13095);
xor U13234 (N_13234,N_12971,N_12985);
nand U13235 (N_13235,N_13102,N_13013);
nor U13236 (N_13236,N_12970,N_12964);
xnor U13237 (N_13237,N_13102,N_13008);
and U13238 (N_13238,N_13051,N_13097);
nand U13239 (N_13239,N_13001,N_13011);
or U13240 (N_13240,N_13085,N_12982);
nand U13241 (N_13241,N_13056,N_13087);
and U13242 (N_13242,N_12987,N_13075);
and U13243 (N_13243,N_13041,N_13103);
and U13244 (N_13244,N_12976,N_13016);
nor U13245 (N_13245,N_12968,N_13056);
xor U13246 (N_13246,N_13028,N_12963);
nand U13247 (N_13247,N_13091,N_12980);
or U13248 (N_13248,N_13111,N_13080);
nor U13249 (N_13249,N_13079,N_13073);
xnor U13250 (N_13250,N_13024,N_13101);
or U13251 (N_13251,N_13078,N_13070);
or U13252 (N_13252,N_13044,N_13056);
nor U13253 (N_13253,N_13029,N_13024);
nor U13254 (N_13254,N_12965,N_12980);
nor U13255 (N_13255,N_12972,N_12973);
or U13256 (N_13256,N_12978,N_13059);
nor U13257 (N_13257,N_13060,N_13096);
or U13258 (N_13258,N_13007,N_13026);
nand U13259 (N_13259,N_13084,N_13014);
xor U13260 (N_13260,N_13080,N_12978);
or U13261 (N_13261,N_13022,N_13042);
xnor U13262 (N_13262,N_12974,N_12972);
nand U13263 (N_13263,N_13047,N_13079);
or U13264 (N_13264,N_12967,N_12975);
nor U13265 (N_13265,N_12989,N_13019);
nor U13266 (N_13266,N_13088,N_12967);
or U13267 (N_13267,N_13001,N_13074);
or U13268 (N_13268,N_12980,N_13089);
nor U13269 (N_13269,N_13081,N_13043);
nand U13270 (N_13270,N_13094,N_13011);
and U13271 (N_13271,N_13025,N_12972);
nand U13272 (N_13272,N_13085,N_13094);
or U13273 (N_13273,N_12997,N_13020);
xor U13274 (N_13274,N_13040,N_13100);
or U13275 (N_13275,N_13068,N_13039);
nand U13276 (N_13276,N_13087,N_13084);
nor U13277 (N_13277,N_13012,N_13078);
nand U13278 (N_13278,N_12977,N_13053);
nand U13279 (N_13279,N_12961,N_12981);
or U13280 (N_13280,N_13123,N_13222);
and U13281 (N_13281,N_13148,N_13133);
nand U13282 (N_13282,N_13151,N_13269);
or U13283 (N_13283,N_13214,N_13232);
xor U13284 (N_13284,N_13272,N_13152);
and U13285 (N_13285,N_13244,N_13169);
xnor U13286 (N_13286,N_13263,N_13258);
nand U13287 (N_13287,N_13185,N_13177);
or U13288 (N_13288,N_13196,N_13271);
nor U13289 (N_13289,N_13203,N_13229);
nand U13290 (N_13290,N_13187,N_13250);
and U13291 (N_13291,N_13202,N_13210);
and U13292 (N_13292,N_13184,N_13255);
or U13293 (N_13293,N_13267,N_13209);
or U13294 (N_13294,N_13197,N_13163);
xnor U13295 (N_13295,N_13162,N_13147);
nor U13296 (N_13296,N_13275,N_13273);
xor U13297 (N_13297,N_13191,N_13259);
or U13298 (N_13298,N_13215,N_13135);
nand U13299 (N_13299,N_13270,N_13276);
nor U13300 (N_13300,N_13132,N_13134);
nand U13301 (N_13301,N_13125,N_13246);
and U13302 (N_13302,N_13160,N_13142);
or U13303 (N_13303,N_13128,N_13236);
nor U13304 (N_13304,N_13240,N_13188);
and U13305 (N_13305,N_13129,N_13216);
nor U13306 (N_13306,N_13159,N_13206);
xnor U13307 (N_13307,N_13278,N_13130);
xnor U13308 (N_13308,N_13178,N_13235);
nor U13309 (N_13309,N_13181,N_13158);
nor U13310 (N_13310,N_13239,N_13265);
or U13311 (N_13311,N_13228,N_13277);
xnor U13312 (N_13312,N_13190,N_13204);
nand U13313 (N_13313,N_13260,N_13268);
and U13314 (N_13314,N_13153,N_13121);
or U13315 (N_13315,N_13221,N_13224);
nand U13316 (N_13316,N_13157,N_13251);
xnor U13317 (N_13317,N_13183,N_13233);
xor U13318 (N_13318,N_13266,N_13168);
and U13319 (N_13319,N_13124,N_13242);
xnor U13320 (N_13320,N_13264,N_13200);
or U13321 (N_13321,N_13249,N_13149);
nand U13322 (N_13322,N_13226,N_13207);
xor U13323 (N_13323,N_13274,N_13213);
nand U13324 (N_13324,N_13253,N_13223);
xnor U13325 (N_13325,N_13165,N_13208);
xor U13326 (N_13326,N_13231,N_13212);
xnor U13327 (N_13327,N_13120,N_13179);
nand U13328 (N_13328,N_13241,N_13131);
nor U13329 (N_13329,N_13127,N_13138);
xor U13330 (N_13330,N_13256,N_13180);
nor U13331 (N_13331,N_13144,N_13211);
and U13332 (N_13332,N_13122,N_13195);
and U13333 (N_13333,N_13175,N_13192);
or U13334 (N_13334,N_13243,N_13166);
or U13335 (N_13335,N_13227,N_13150);
xnor U13336 (N_13336,N_13146,N_13254);
and U13337 (N_13337,N_13182,N_13193);
nand U13338 (N_13338,N_13247,N_13126);
or U13339 (N_13339,N_13248,N_13262);
or U13340 (N_13340,N_13167,N_13219);
and U13341 (N_13341,N_13145,N_13174);
and U13342 (N_13342,N_13156,N_13279);
or U13343 (N_13343,N_13234,N_13170);
nor U13344 (N_13344,N_13161,N_13137);
and U13345 (N_13345,N_13245,N_13257);
xnor U13346 (N_13346,N_13172,N_13217);
or U13347 (N_13347,N_13164,N_13198);
nand U13348 (N_13348,N_13136,N_13237);
xor U13349 (N_13349,N_13176,N_13194);
xnor U13350 (N_13350,N_13141,N_13189);
and U13351 (N_13351,N_13238,N_13155);
and U13352 (N_13352,N_13139,N_13201);
nand U13353 (N_13353,N_13140,N_13225);
nor U13354 (N_13354,N_13186,N_13218);
or U13355 (N_13355,N_13143,N_13261);
xnor U13356 (N_13356,N_13205,N_13199);
xnor U13357 (N_13357,N_13171,N_13173);
or U13358 (N_13358,N_13154,N_13252);
nor U13359 (N_13359,N_13230,N_13220);
or U13360 (N_13360,N_13126,N_13165);
or U13361 (N_13361,N_13208,N_13161);
and U13362 (N_13362,N_13129,N_13209);
nor U13363 (N_13363,N_13197,N_13261);
or U13364 (N_13364,N_13161,N_13194);
and U13365 (N_13365,N_13181,N_13160);
and U13366 (N_13366,N_13207,N_13275);
or U13367 (N_13367,N_13177,N_13257);
and U13368 (N_13368,N_13252,N_13266);
and U13369 (N_13369,N_13145,N_13275);
nor U13370 (N_13370,N_13189,N_13210);
xor U13371 (N_13371,N_13262,N_13205);
xnor U13372 (N_13372,N_13186,N_13230);
nor U13373 (N_13373,N_13174,N_13250);
xor U13374 (N_13374,N_13257,N_13125);
nand U13375 (N_13375,N_13256,N_13222);
xor U13376 (N_13376,N_13218,N_13205);
nand U13377 (N_13377,N_13132,N_13220);
or U13378 (N_13378,N_13167,N_13239);
or U13379 (N_13379,N_13245,N_13162);
or U13380 (N_13380,N_13203,N_13141);
xor U13381 (N_13381,N_13203,N_13146);
xor U13382 (N_13382,N_13256,N_13146);
or U13383 (N_13383,N_13153,N_13203);
xor U13384 (N_13384,N_13264,N_13181);
nor U13385 (N_13385,N_13268,N_13169);
or U13386 (N_13386,N_13167,N_13136);
nand U13387 (N_13387,N_13253,N_13249);
or U13388 (N_13388,N_13129,N_13225);
xnor U13389 (N_13389,N_13263,N_13234);
xor U13390 (N_13390,N_13123,N_13160);
and U13391 (N_13391,N_13218,N_13207);
and U13392 (N_13392,N_13242,N_13178);
nor U13393 (N_13393,N_13126,N_13264);
and U13394 (N_13394,N_13222,N_13257);
nand U13395 (N_13395,N_13125,N_13148);
or U13396 (N_13396,N_13268,N_13256);
and U13397 (N_13397,N_13261,N_13180);
and U13398 (N_13398,N_13234,N_13179);
xor U13399 (N_13399,N_13208,N_13274);
or U13400 (N_13400,N_13246,N_13216);
or U13401 (N_13401,N_13175,N_13122);
or U13402 (N_13402,N_13190,N_13260);
or U13403 (N_13403,N_13239,N_13146);
and U13404 (N_13404,N_13135,N_13175);
or U13405 (N_13405,N_13273,N_13274);
and U13406 (N_13406,N_13124,N_13248);
or U13407 (N_13407,N_13177,N_13183);
nand U13408 (N_13408,N_13181,N_13204);
or U13409 (N_13409,N_13184,N_13149);
nand U13410 (N_13410,N_13244,N_13161);
and U13411 (N_13411,N_13134,N_13240);
nand U13412 (N_13412,N_13164,N_13245);
or U13413 (N_13413,N_13235,N_13204);
or U13414 (N_13414,N_13130,N_13186);
nor U13415 (N_13415,N_13130,N_13159);
nand U13416 (N_13416,N_13188,N_13207);
or U13417 (N_13417,N_13238,N_13204);
nand U13418 (N_13418,N_13257,N_13200);
nor U13419 (N_13419,N_13173,N_13142);
xor U13420 (N_13420,N_13177,N_13152);
nor U13421 (N_13421,N_13278,N_13190);
xnor U13422 (N_13422,N_13158,N_13120);
and U13423 (N_13423,N_13249,N_13259);
xnor U13424 (N_13424,N_13231,N_13144);
xor U13425 (N_13425,N_13196,N_13243);
and U13426 (N_13426,N_13249,N_13189);
and U13427 (N_13427,N_13183,N_13277);
and U13428 (N_13428,N_13141,N_13149);
and U13429 (N_13429,N_13133,N_13197);
nor U13430 (N_13430,N_13230,N_13123);
and U13431 (N_13431,N_13163,N_13210);
xnor U13432 (N_13432,N_13159,N_13235);
xnor U13433 (N_13433,N_13225,N_13275);
nor U13434 (N_13434,N_13263,N_13242);
xnor U13435 (N_13435,N_13237,N_13142);
xnor U13436 (N_13436,N_13210,N_13141);
nor U13437 (N_13437,N_13248,N_13205);
nand U13438 (N_13438,N_13215,N_13267);
and U13439 (N_13439,N_13145,N_13254);
and U13440 (N_13440,N_13372,N_13301);
xnor U13441 (N_13441,N_13416,N_13360);
nand U13442 (N_13442,N_13341,N_13370);
or U13443 (N_13443,N_13354,N_13292);
and U13444 (N_13444,N_13328,N_13388);
and U13445 (N_13445,N_13433,N_13411);
and U13446 (N_13446,N_13408,N_13400);
xor U13447 (N_13447,N_13280,N_13306);
nor U13448 (N_13448,N_13300,N_13347);
nand U13449 (N_13449,N_13415,N_13373);
xor U13450 (N_13450,N_13351,N_13285);
nor U13451 (N_13451,N_13417,N_13382);
nand U13452 (N_13452,N_13439,N_13409);
or U13453 (N_13453,N_13323,N_13368);
nand U13454 (N_13454,N_13325,N_13294);
and U13455 (N_13455,N_13378,N_13299);
nand U13456 (N_13456,N_13402,N_13377);
nor U13457 (N_13457,N_13349,N_13421);
xor U13458 (N_13458,N_13304,N_13381);
or U13459 (N_13459,N_13380,N_13362);
and U13460 (N_13460,N_13406,N_13432);
nand U13461 (N_13461,N_13399,N_13437);
nand U13462 (N_13462,N_13392,N_13394);
xor U13463 (N_13463,N_13289,N_13283);
xnor U13464 (N_13464,N_13308,N_13383);
xor U13465 (N_13465,N_13295,N_13396);
nand U13466 (N_13466,N_13314,N_13288);
xor U13467 (N_13467,N_13311,N_13307);
nand U13468 (N_13468,N_13329,N_13375);
xnor U13469 (N_13469,N_13350,N_13356);
nand U13470 (N_13470,N_13365,N_13296);
xor U13471 (N_13471,N_13355,N_13357);
nand U13472 (N_13472,N_13391,N_13371);
nand U13473 (N_13473,N_13390,N_13290);
and U13474 (N_13474,N_13425,N_13309);
nand U13475 (N_13475,N_13403,N_13389);
nand U13476 (N_13476,N_13320,N_13340);
and U13477 (N_13477,N_13324,N_13282);
nand U13478 (N_13478,N_13423,N_13404);
xor U13479 (N_13479,N_13366,N_13374);
and U13480 (N_13480,N_13286,N_13318);
or U13481 (N_13481,N_13331,N_13332);
and U13482 (N_13482,N_13313,N_13322);
nor U13483 (N_13483,N_13435,N_13401);
or U13484 (N_13484,N_13407,N_13405);
xnor U13485 (N_13485,N_13312,N_13337);
nand U13486 (N_13486,N_13291,N_13413);
nand U13487 (N_13487,N_13353,N_13348);
nand U13488 (N_13488,N_13339,N_13398);
nand U13489 (N_13489,N_13412,N_13336);
nor U13490 (N_13490,N_13395,N_13376);
nor U13491 (N_13491,N_13321,N_13305);
and U13492 (N_13492,N_13369,N_13386);
or U13493 (N_13493,N_13345,N_13310);
xnor U13494 (N_13494,N_13420,N_13419);
or U13495 (N_13495,N_13287,N_13387);
and U13496 (N_13496,N_13297,N_13342);
and U13497 (N_13497,N_13393,N_13335);
xnor U13498 (N_13498,N_13361,N_13281);
and U13499 (N_13499,N_13293,N_13426);
and U13500 (N_13500,N_13316,N_13428);
and U13501 (N_13501,N_13397,N_13326);
nor U13502 (N_13502,N_13422,N_13330);
nand U13503 (N_13503,N_13363,N_13385);
xnor U13504 (N_13504,N_13364,N_13359);
or U13505 (N_13505,N_13315,N_13334);
xnor U13506 (N_13506,N_13358,N_13430);
and U13507 (N_13507,N_13317,N_13429);
nor U13508 (N_13508,N_13431,N_13338);
nor U13509 (N_13509,N_13410,N_13436);
or U13510 (N_13510,N_13384,N_13418);
or U13511 (N_13511,N_13327,N_13438);
nor U13512 (N_13512,N_13344,N_13427);
or U13513 (N_13513,N_13434,N_13303);
and U13514 (N_13514,N_13333,N_13414);
and U13515 (N_13515,N_13284,N_13352);
or U13516 (N_13516,N_13367,N_13346);
xor U13517 (N_13517,N_13302,N_13319);
nor U13518 (N_13518,N_13298,N_13379);
xor U13519 (N_13519,N_13343,N_13424);
or U13520 (N_13520,N_13406,N_13437);
and U13521 (N_13521,N_13368,N_13435);
nor U13522 (N_13522,N_13298,N_13339);
and U13523 (N_13523,N_13343,N_13388);
xnor U13524 (N_13524,N_13337,N_13369);
or U13525 (N_13525,N_13404,N_13375);
and U13526 (N_13526,N_13300,N_13428);
xnor U13527 (N_13527,N_13365,N_13330);
nand U13528 (N_13528,N_13429,N_13435);
nand U13529 (N_13529,N_13355,N_13336);
or U13530 (N_13530,N_13384,N_13363);
and U13531 (N_13531,N_13415,N_13289);
or U13532 (N_13532,N_13415,N_13355);
or U13533 (N_13533,N_13435,N_13325);
xnor U13534 (N_13534,N_13369,N_13330);
xor U13535 (N_13535,N_13296,N_13352);
xnor U13536 (N_13536,N_13313,N_13332);
nor U13537 (N_13537,N_13409,N_13306);
xnor U13538 (N_13538,N_13301,N_13304);
nand U13539 (N_13539,N_13338,N_13352);
nor U13540 (N_13540,N_13338,N_13419);
nand U13541 (N_13541,N_13349,N_13339);
xor U13542 (N_13542,N_13378,N_13425);
and U13543 (N_13543,N_13435,N_13326);
nor U13544 (N_13544,N_13437,N_13387);
nor U13545 (N_13545,N_13303,N_13362);
or U13546 (N_13546,N_13292,N_13421);
nand U13547 (N_13547,N_13340,N_13415);
xnor U13548 (N_13548,N_13418,N_13383);
and U13549 (N_13549,N_13325,N_13317);
and U13550 (N_13550,N_13302,N_13407);
and U13551 (N_13551,N_13352,N_13379);
nor U13552 (N_13552,N_13415,N_13332);
and U13553 (N_13553,N_13331,N_13439);
and U13554 (N_13554,N_13287,N_13401);
nand U13555 (N_13555,N_13322,N_13348);
and U13556 (N_13556,N_13396,N_13374);
nor U13557 (N_13557,N_13289,N_13410);
nor U13558 (N_13558,N_13430,N_13360);
xnor U13559 (N_13559,N_13387,N_13400);
or U13560 (N_13560,N_13353,N_13370);
or U13561 (N_13561,N_13323,N_13396);
nand U13562 (N_13562,N_13353,N_13435);
nor U13563 (N_13563,N_13289,N_13371);
and U13564 (N_13564,N_13398,N_13403);
xnor U13565 (N_13565,N_13435,N_13301);
nand U13566 (N_13566,N_13296,N_13380);
nor U13567 (N_13567,N_13372,N_13381);
and U13568 (N_13568,N_13324,N_13375);
nor U13569 (N_13569,N_13425,N_13346);
or U13570 (N_13570,N_13329,N_13320);
or U13571 (N_13571,N_13390,N_13351);
nor U13572 (N_13572,N_13302,N_13344);
nand U13573 (N_13573,N_13428,N_13410);
or U13574 (N_13574,N_13388,N_13284);
nor U13575 (N_13575,N_13344,N_13434);
or U13576 (N_13576,N_13422,N_13381);
xor U13577 (N_13577,N_13354,N_13356);
or U13578 (N_13578,N_13307,N_13347);
or U13579 (N_13579,N_13370,N_13384);
nand U13580 (N_13580,N_13416,N_13383);
nand U13581 (N_13581,N_13436,N_13425);
nor U13582 (N_13582,N_13288,N_13370);
and U13583 (N_13583,N_13372,N_13346);
or U13584 (N_13584,N_13438,N_13435);
or U13585 (N_13585,N_13308,N_13385);
nor U13586 (N_13586,N_13425,N_13403);
and U13587 (N_13587,N_13355,N_13366);
nand U13588 (N_13588,N_13294,N_13380);
nand U13589 (N_13589,N_13323,N_13326);
and U13590 (N_13590,N_13381,N_13290);
or U13591 (N_13591,N_13435,N_13319);
nor U13592 (N_13592,N_13294,N_13303);
and U13593 (N_13593,N_13410,N_13312);
nor U13594 (N_13594,N_13292,N_13317);
nor U13595 (N_13595,N_13362,N_13425);
xnor U13596 (N_13596,N_13416,N_13401);
nand U13597 (N_13597,N_13439,N_13297);
xor U13598 (N_13598,N_13368,N_13288);
and U13599 (N_13599,N_13380,N_13428);
nor U13600 (N_13600,N_13472,N_13444);
nand U13601 (N_13601,N_13538,N_13542);
xnor U13602 (N_13602,N_13479,N_13595);
xnor U13603 (N_13603,N_13578,N_13586);
or U13604 (N_13604,N_13574,N_13478);
nand U13605 (N_13605,N_13598,N_13445);
xnor U13606 (N_13606,N_13446,N_13463);
nand U13607 (N_13607,N_13487,N_13523);
and U13608 (N_13608,N_13459,N_13453);
or U13609 (N_13609,N_13525,N_13469);
and U13610 (N_13610,N_13468,N_13488);
nand U13611 (N_13611,N_13599,N_13510);
nand U13612 (N_13612,N_13502,N_13499);
nor U13613 (N_13613,N_13485,N_13577);
nor U13614 (N_13614,N_13455,N_13591);
or U13615 (N_13615,N_13547,N_13451);
nand U13616 (N_13616,N_13458,N_13569);
nand U13617 (N_13617,N_13592,N_13442);
nand U13618 (N_13618,N_13526,N_13562);
xor U13619 (N_13619,N_13518,N_13536);
or U13620 (N_13620,N_13593,N_13597);
nor U13621 (N_13621,N_13564,N_13483);
or U13622 (N_13622,N_13447,N_13549);
and U13623 (N_13623,N_13529,N_13568);
nand U13624 (N_13624,N_13482,N_13579);
xor U13625 (N_13625,N_13519,N_13589);
or U13626 (N_13626,N_13594,N_13557);
or U13627 (N_13627,N_13491,N_13516);
nor U13628 (N_13628,N_13546,N_13558);
nor U13629 (N_13629,N_13489,N_13484);
or U13630 (N_13630,N_13587,N_13545);
xnor U13631 (N_13631,N_13573,N_13456);
and U13632 (N_13632,N_13582,N_13501);
nor U13633 (N_13633,N_13532,N_13596);
or U13634 (N_13634,N_13555,N_13521);
and U13635 (N_13635,N_13454,N_13535);
and U13636 (N_13636,N_13551,N_13560);
and U13637 (N_13637,N_13513,N_13503);
nor U13638 (N_13638,N_13567,N_13512);
and U13639 (N_13639,N_13580,N_13490);
nand U13640 (N_13640,N_13584,N_13576);
xor U13641 (N_13641,N_13511,N_13466);
or U13642 (N_13642,N_13553,N_13481);
nor U13643 (N_13643,N_13505,N_13540);
nand U13644 (N_13644,N_13480,N_13470);
and U13645 (N_13645,N_13515,N_13533);
xnor U13646 (N_13646,N_13443,N_13572);
nand U13647 (N_13647,N_13448,N_13552);
nand U13648 (N_13648,N_13575,N_13530);
nor U13649 (N_13649,N_13506,N_13517);
or U13650 (N_13650,N_13590,N_13556);
nand U13651 (N_13651,N_13477,N_13441);
or U13652 (N_13652,N_13462,N_13585);
or U13653 (N_13653,N_13570,N_13500);
or U13654 (N_13654,N_13522,N_13581);
nand U13655 (N_13655,N_13507,N_13457);
nor U13656 (N_13656,N_13550,N_13498);
xnor U13657 (N_13657,N_13514,N_13492);
nor U13658 (N_13658,N_13583,N_13493);
nor U13659 (N_13659,N_13565,N_13508);
nand U13660 (N_13660,N_13537,N_13476);
or U13661 (N_13661,N_13528,N_13527);
or U13662 (N_13662,N_13534,N_13495);
and U13663 (N_13663,N_13475,N_13524);
and U13664 (N_13664,N_13520,N_13509);
xnor U13665 (N_13665,N_13465,N_13473);
or U13666 (N_13666,N_13486,N_13543);
or U13667 (N_13667,N_13467,N_13449);
nand U13668 (N_13668,N_13559,N_13539);
nor U13669 (N_13669,N_13494,N_13541);
and U13670 (N_13670,N_13554,N_13531);
or U13671 (N_13671,N_13461,N_13548);
nand U13672 (N_13672,N_13440,N_13504);
nor U13673 (N_13673,N_13497,N_13561);
and U13674 (N_13674,N_13464,N_13544);
nand U13675 (N_13675,N_13471,N_13460);
or U13676 (N_13676,N_13588,N_13496);
and U13677 (N_13677,N_13450,N_13563);
or U13678 (N_13678,N_13452,N_13571);
and U13679 (N_13679,N_13566,N_13474);
or U13680 (N_13680,N_13594,N_13467);
nor U13681 (N_13681,N_13533,N_13442);
nand U13682 (N_13682,N_13455,N_13474);
nand U13683 (N_13683,N_13532,N_13563);
and U13684 (N_13684,N_13543,N_13448);
and U13685 (N_13685,N_13453,N_13528);
or U13686 (N_13686,N_13474,N_13531);
nand U13687 (N_13687,N_13560,N_13507);
nand U13688 (N_13688,N_13463,N_13518);
nand U13689 (N_13689,N_13525,N_13464);
xnor U13690 (N_13690,N_13552,N_13597);
nand U13691 (N_13691,N_13448,N_13528);
nand U13692 (N_13692,N_13469,N_13455);
and U13693 (N_13693,N_13481,N_13544);
nor U13694 (N_13694,N_13566,N_13481);
and U13695 (N_13695,N_13490,N_13494);
xnor U13696 (N_13696,N_13536,N_13578);
nor U13697 (N_13697,N_13543,N_13496);
nand U13698 (N_13698,N_13553,N_13557);
nand U13699 (N_13699,N_13573,N_13558);
and U13700 (N_13700,N_13472,N_13499);
nand U13701 (N_13701,N_13498,N_13496);
nor U13702 (N_13702,N_13489,N_13535);
xor U13703 (N_13703,N_13549,N_13525);
nor U13704 (N_13704,N_13587,N_13597);
and U13705 (N_13705,N_13520,N_13483);
nand U13706 (N_13706,N_13444,N_13565);
and U13707 (N_13707,N_13484,N_13504);
and U13708 (N_13708,N_13459,N_13468);
nand U13709 (N_13709,N_13559,N_13533);
or U13710 (N_13710,N_13457,N_13513);
and U13711 (N_13711,N_13467,N_13497);
nor U13712 (N_13712,N_13442,N_13446);
xnor U13713 (N_13713,N_13492,N_13494);
xor U13714 (N_13714,N_13581,N_13484);
and U13715 (N_13715,N_13477,N_13540);
nand U13716 (N_13716,N_13575,N_13482);
nand U13717 (N_13717,N_13499,N_13455);
nor U13718 (N_13718,N_13559,N_13535);
and U13719 (N_13719,N_13519,N_13461);
xnor U13720 (N_13720,N_13486,N_13445);
nor U13721 (N_13721,N_13586,N_13501);
nor U13722 (N_13722,N_13588,N_13597);
or U13723 (N_13723,N_13447,N_13451);
or U13724 (N_13724,N_13568,N_13547);
nor U13725 (N_13725,N_13576,N_13440);
or U13726 (N_13726,N_13532,N_13455);
or U13727 (N_13727,N_13461,N_13596);
xor U13728 (N_13728,N_13519,N_13495);
or U13729 (N_13729,N_13526,N_13575);
nand U13730 (N_13730,N_13458,N_13502);
xnor U13731 (N_13731,N_13540,N_13499);
xnor U13732 (N_13732,N_13511,N_13565);
xor U13733 (N_13733,N_13451,N_13499);
and U13734 (N_13734,N_13478,N_13586);
nand U13735 (N_13735,N_13471,N_13504);
or U13736 (N_13736,N_13541,N_13565);
nor U13737 (N_13737,N_13572,N_13555);
nor U13738 (N_13738,N_13496,N_13515);
xor U13739 (N_13739,N_13573,N_13591);
xor U13740 (N_13740,N_13516,N_13543);
xnor U13741 (N_13741,N_13561,N_13534);
or U13742 (N_13742,N_13441,N_13522);
nor U13743 (N_13743,N_13470,N_13518);
nor U13744 (N_13744,N_13506,N_13521);
or U13745 (N_13745,N_13503,N_13453);
nand U13746 (N_13746,N_13482,N_13571);
and U13747 (N_13747,N_13494,N_13590);
or U13748 (N_13748,N_13550,N_13478);
nor U13749 (N_13749,N_13546,N_13509);
nand U13750 (N_13750,N_13530,N_13452);
or U13751 (N_13751,N_13498,N_13553);
nor U13752 (N_13752,N_13526,N_13598);
nand U13753 (N_13753,N_13592,N_13578);
and U13754 (N_13754,N_13596,N_13471);
and U13755 (N_13755,N_13500,N_13487);
nor U13756 (N_13756,N_13533,N_13482);
or U13757 (N_13757,N_13542,N_13449);
xor U13758 (N_13758,N_13561,N_13592);
nand U13759 (N_13759,N_13512,N_13482);
or U13760 (N_13760,N_13658,N_13629);
nor U13761 (N_13761,N_13738,N_13612);
nand U13762 (N_13762,N_13633,N_13666);
and U13763 (N_13763,N_13683,N_13635);
xor U13764 (N_13764,N_13747,N_13695);
nand U13765 (N_13765,N_13631,N_13718);
nand U13766 (N_13766,N_13724,N_13620);
and U13767 (N_13767,N_13609,N_13674);
or U13768 (N_13768,N_13676,N_13726);
xnor U13769 (N_13769,N_13709,N_13693);
and U13770 (N_13770,N_13702,N_13696);
and U13771 (N_13771,N_13686,N_13737);
nor U13772 (N_13772,N_13735,N_13721);
or U13773 (N_13773,N_13741,N_13627);
nor U13774 (N_13774,N_13700,N_13719);
xnor U13775 (N_13775,N_13630,N_13757);
nor U13776 (N_13776,N_13649,N_13754);
and U13777 (N_13777,N_13714,N_13756);
nor U13778 (N_13778,N_13697,N_13680);
nor U13779 (N_13779,N_13672,N_13600);
nor U13780 (N_13780,N_13653,N_13643);
nor U13781 (N_13781,N_13698,N_13660);
xnor U13782 (N_13782,N_13728,N_13692);
or U13783 (N_13783,N_13716,N_13617);
nand U13784 (N_13784,N_13694,N_13717);
nand U13785 (N_13785,N_13740,N_13688);
nor U13786 (N_13786,N_13748,N_13750);
xor U13787 (N_13787,N_13759,N_13712);
nand U13788 (N_13788,N_13638,N_13689);
or U13789 (N_13789,N_13647,N_13713);
or U13790 (N_13790,N_13632,N_13704);
and U13791 (N_13791,N_13613,N_13668);
xor U13792 (N_13792,N_13691,N_13652);
or U13793 (N_13793,N_13755,N_13670);
nor U13794 (N_13794,N_13651,N_13644);
or U13795 (N_13795,N_13752,N_13710);
or U13796 (N_13796,N_13646,N_13677);
and U13797 (N_13797,N_13628,N_13634);
nor U13798 (N_13798,N_13687,N_13707);
nor U13799 (N_13799,N_13655,N_13679);
and U13800 (N_13800,N_13682,N_13673);
and U13801 (N_13801,N_13641,N_13640);
nand U13802 (N_13802,N_13690,N_13648);
or U13803 (N_13803,N_13711,N_13624);
or U13804 (N_13804,N_13732,N_13684);
nor U13805 (N_13805,N_13720,N_13608);
nand U13806 (N_13806,N_13731,N_13730);
and U13807 (N_13807,N_13619,N_13739);
nand U13808 (N_13808,N_13725,N_13722);
or U13809 (N_13809,N_13699,N_13605);
xor U13810 (N_13810,N_13749,N_13606);
nand U13811 (N_13811,N_13656,N_13667);
nor U13812 (N_13812,N_13715,N_13746);
nor U13813 (N_13813,N_13642,N_13745);
or U13814 (N_13814,N_13602,N_13681);
xor U13815 (N_13815,N_13729,N_13678);
and U13816 (N_13816,N_13614,N_13671);
and U13817 (N_13817,N_13703,N_13744);
and U13818 (N_13818,N_13625,N_13661);
nor U13819 (N_13819,N_13705,N_13663);
and U13820 (N_13820,N_13637,N_13751);
nor U13821 (N_13821,N_13618,N_13616);
or U13822 (N_13822,N_13607,N_13639);
nand U13823 (N_13823,N_13601,N_13742);
xor U13824 (N_13824,N_13622,N_13733);
xnor U13825 (N_13825,N_13664,N_13753);
nor U13826 (N_13826,N_13662,N_13723);
nand U13827 (N_13827,N_13685,N_13758);
and U13828 (N_13828,N_13659,N_13604);
nand U13829 (N_13829,N_13708,N_13675);
xnor U13830 (N_13830,N_13654,N_13603);
or U13831 (N_13831,N_13706,N_13743);
xnor U13832 (N_13832,N_13626,N_13701);
xnor U13833 (N_13833,N_13615,N_13636);
nor U13834 (N_13834,N_13665,N_13611);
xor U13835 (N_13835,N_13734,N_13610);
nand U13836 (N_13836,N_13669,N_13727);
or U13837 (N_13837,N_13645,N_13657);
xor U13838 (N_13838,N_13650,N_13736);
nand U13839 (N_13839,N_13623,N_13621);
or U13840 (N_13840,N_13726,N_13655);
or U13841 (N_13841,N_13675,N_13697);
xnor U13842 (N_13842,N_13700,N_13666);
and U13843 (N_13843,N_13653,N_13677);
nand U13844 (N_13844,N_13691,N_13727);
nor U13845 (N_13845,N_13633,N_13649);
or U13846 (N_13846,N_13672,N_13702);
or U13847 (N_13847,N_13647,N_13659);
nand U13848 (N_13848,N_13631,N_13609);
xor U13849 (N_13849,N_13620,N_13659);
xor U13850 (N_13850,N_13714,N_13669);
and U13851 (N_13851,N_13756,N_13695);
and U13852 (N_13852,N_13684,N_13644);
nor U13853 (N_13853,N_13616,N_13717);
nor U13854 (N_13854,N_13677,N_13674);
nand U13855 (N_13855,N_13677,N_13721);
nand U13856 (N_13856,N_13757,N_13702);
or U13857 (N_13857,N_13706,N_13652);
xor U13858 (N_13858,N_13612,N_13710);
nand U13859 (N_13859,N_13683,N_13612);
or U13860 (N_13860,N_13624,N_13646);
nand U13861 (N_13861,N_13694,N_13684);
xor U13862 (N_13862,N_13685,N_13695);
nand U13863 (N_13863,N_13695,N_13642);
xor U13864 (N_13864,N_13663,N_13716);
nand U13865 (N_13865,N_13692,N_13673);
nand U13866 (N_13866,N_13639,N_13673);
nand U13867 (N_13867,N_13687,N_13619);
and U13868 (N_13868,N_13677,N_13683);
nand U13869 (N_13869,N_13603,N_13635);
nor U13870 (N_13870,N_13701,N_13683);
and U13871 (N_13871,N_13741,N_13683);
nor U13872 (N_13872,N_13633,N_13702);
or U13873 (N_13873,N_13635,N_13653);
xnor U13874 (N_13874,N_13736,N_13719);
and U13875 (N_13875,N_13736,N_13682);
or U13876 (N_13876,N_13673,N_13626);
or U13877 (N_13877,N_13723,N_13740);
nand U13878 (N_13878,N_13657,N_13642);
and U13879 (N_13879,N_13742,N_13715);
and U13880 (N_13880,N_13673,N_13661);
and U13881 (N_13881,N_13667,N_13679);
or U13882 (N_13882,N_13658,N_13759);
nand U13883 (N_13883,N_13754,N_13759);
nor U13884 (N_13884,N_13744,N_13708);
nand U13885 (N_13885,N_13690,N_13718);
xnor U13886 (N_13886,N_13681,N_13621);
nor U13887 (N_13887,N_13737,N_13654);
nor U13888 (N_13888,N_13700,N_13702);
nand U13889 (N_13889,N_13686,N_13699);
or U13890 (N_13890,N_13641,N_13651);
xor U13891 (N_13891,N_13658,N_13630);
and U13892 (N_13892,N_13621,N_13633);
xnor U13893 (N_13893,N_13666,N_13747);
nand U13894 (N_13894,N_13686,N_13605);
or U13895 (N_13895,N_13714,N_13703);
and U13896 (N_13896,N_13742,N_13753);
or U13897 (N_13897,N_13694,N_13622);
nor U13898 (N_13898,N_13703,N_13650);
xor U13899 (N_13899,N_13627,N_13604);
nand U13900 (N_13900,N_13753,N_13696);
and U13901 (N_13901,N_13750,N_13630);
xnor U13902 (N_13902,N_13619,N_13682);
nor U13903 (N_13903,N_13739,N_13755);
nand U13904 (N_13904,N_13669,N_13746);
or U13905 (N_13905,N_13670,N_13611);
nor U13906 (N_13906,N_13701,N_13700);
nand U13907 (N_13907,N_13660,N_13648);
nor U13908 (N_13908,N_13704,N_13721);
xor U13909 (N_13909,N_13627,N_13722);
nor U13910 (N_13910,N_13659,N_13657);
nand U13911 (N_13911,N_13724,N_13756);
nor U13912 (N_13912,N_13732,N_13635);
xnor U13913 (N_13913,N_13689,N_13724);
nand U13914 (N_13914,N_13659,N_13686);
and U13915 (N_13915,N_13611,N_13733);
or U13916 (N_13916,N_13640,N_13667);
and U13917 (N_13917,N_13608,N_13642);
or U13918 (N_13918,N_13703,N_13600);
and U13919 (N_13919,N_13721,N_13659);
xor U13920 (N_13920,N_13827,N_13849);
nand U13921 (N_13921,N_13803,N_13864);
nand U13922 (N_13922,N_13823,N_13835);
nor U13923 (N_13923,N_13866,N_13824);
and U13924 (N_13924,N_13764,N_13858);
or U13925 (N_13925,N_13867,N_13839);
nor U13926 (N_13926,N_13848,N_13777);
nor U13927 (N_13927,N_13880,N_13818);
xnor U13928 (N_13928,N_13798,N_13837);
nand U13929 (N_13929,N_13822,N_13903);
or U13930 (N_13930,N_13860,N_13846);
and U13931 (N_13931,N_13801,N_13871);
nand U13932 (N_13932,N_13789,N_13865);
nand U13933 (N_13933,N_13895,N_13815);
xnor U13934 (N_13934,N_13853,N_13766);
nand U13935 (N_13935,N_13886,N_13857);
nor U13936 (N_13936,N_13917,N_13773);
nand U13937 (N_13937,N_13795,N_13770);
xor U13938 (N_13938,N_13778,N_13782);
and U13939 (N_13939,N_13807,N_13787);
xnor U13940 (N_13940,N_13873,N_13877);
nor U13941 (N_13941,N_13768,N_13916);
or U13942 (N_13942,N_13902,N_13898);
and U13943 (N_13943,N_13878,N_13881);
or U13944 (N_13944,N_13804,N_13841);
or U13945 (N_13945,N_13914,N_13887);
and U13946 (N_13946,N_13771,N_13809);
and U13947 (N_13947,N_13834,N_13876);
xor U13948 (N_13948,N_13911,N_13859);
or U13949 (N_13949,N_13765,N_13825);
xor U13950 (N_13950,N_13769,N_13780);
xor U13951 (N_13951,N_13790,N_13872);
or U13952 (N_13952,N_13893,N_13806);
and U13953 (N_13953,N_13775,N_13863);
and U13954 (N_13954,N_13861,N_13868);
and U13955 (N_13955,N_13796,N_13802);
and U13956 (N_13956,N_13833,N_13910);
nor U13957 (N_13957,N_13840,N_13897);
or U13958 (N_13958,N_13847,N_13811);
nand U13959 (N_13959,N_13781,N_13786);
and U13960 (N_13960,N_13767,N_13772);
or U13961 (N_13961,N_13843,N_13820);
and U13962 (N_13962,N_13819,N_13913);
xnor U13963 (N_13963,N_13792,N_13828);
or U13964 (N_13964,N_13912,N_13892);
or U13965 (N_13965,N_13875,N_13826);
or U13966 (N_13966,N_13762,N_13785);
or U13967 (N_13967,N_13810,N_13883);
and U13968 (N_13968,N_13908,N_13882);
xor U13969 (N_13969,N_13900,N_13905);
xnor U13970 (N_13970,N_13919,N_13797);
and U13971 (N_13971,N_13832,N_13836);
and U13972 (N_13972,N_13906,N_13844);
nand U13973 (N_13973,N_13808,N_13854);
and U13974 (N_13974,N_13788,N_13830);
nor U13975 (N_13975,N_13852,N_13793);
or U13976 (N_13976,N_13890,N_13885);
nand U13977 (N_13977,N_13821,N_13884);
nor U13978 (N_13978,N_13894,N_13845);
xor U13979 (N_13979,N_13869,N_13891);
xnor U13980 (N_13980,N_13889,N_13888);
xnor U13981 (N_13981,N_13784,N_13805);
nor U13982 (N_13982,N_13850,N_13831);
and U13983 (N_13983,N_13774,N_13915);
xnor U13984 (N_13984,N_13870,N_13776);
nor U13985 (N_13985,N_13761,N_13838);
and U13986 (N_13986,N_13896,N_13817);
or U13987 (N_13987,N_13874,N_13856);
nor U13988 (N_13988,N_13899,N_13842);
xnor U13989 (N_13989,N_13794,N_13816);
xor U13990 (N_13990,N_13800,N_13791);
or U13991 (N_13991,N_13879,N_13909);
nand U13992 (N_13992,N_13862,N_13829);
xnor U13993 (N_13993,N_13918,N_13799);
nand U13994 (N_13994,N_13763,N_13814);
nor U13995 (N_13995,N_13779,N_13760);
or U13996 (N_13996,N_13813,N_13855);
or U13997 (N_13997,N_13783,N_13851);
xnor U13998 (N_13998,N_13907,N_13901);
and U13999 (N_13999,N_13812,N_13904);
xnor U14000 (N_14000,N_13816,N_13842);
nor U14001 (N_14001,N_13815,N_13817);
xor U14002 (N_14002,N_13833,N_13774);
nor U14003 (N_14003,N_13901,N_13850);
nor U14004 (N_14004,N_13864,N_13880);
or U14005 (N_14005,N_13853,N_13810);
and U14006 (N_14006,N_13833,N_13907);
nor U14007 (N_14007,N_13916,N_13777);
nor U14008 (N_14008,N_13771,N_13904);
or U14009 (N_14009,N_13818,N_13809);
or U14010 (N_14010,N_13874,N_13824);
xor U14011 (N_14011,N_13808,N_13862);
and U14012 (N_14012,N_13847,N_13884);
nand U14013 (N_14013,N_13828,N_13801);
nor U14014 (N_14014,N_13917,N_13860);
nand U14015 (N_14015,N_13785,N_13796);
or U14016 (N_14016,N_13919,N_13871);
and U14017 (N_14017,N_13868,N_13869);
nand U14018 (N_14018,N_13912,N_13784);
nand U14019 (N_14019,N_13845,N_13841);
nor U14020 (N_14020,N_13831,N_13800);
nor U14021 (N_14021,N_13854,N_13836);
and U14022 (N_14022,N_13861,N_13903);
xnor U14023 (N_14023,N_13771,N_13876);
nor U14024 (N_14024,N_13769,N_13862);
nor U14025 (N_14025,N_13875,N_13902);
nand U14026 (N_14026,N_13800,N_13799);
nand U14027 (N_14027,N_13848,N_13828);
or U14028 (N_14028,N_13901,N_13875);
and U14029 (N_14029,N_13894,N_13806);
nand U14030 (N_14030,N_13908,N_13839);
xnor U14031 (N_14031,N_13826,N_13767);
nand U14032 (N_14032,N_13826,N_13888);
nand U14033 (N_14033,N_13788,N_13885);
nand U14034 (N_14034,N_13774,N_13837);
nand U14035 (N_14035,N_13794,N_13764);
and U14036 (N_14036,N_13804,N_13877);
and U14037 (N_14037,N_13866,N_13836);
nor U14038 (N_14038,N_13820,N_13835);
and U14039 (N_14039,N_13824,N_13800);
and U14040 (N_14040,N_13820,N_13813);
and U14041 (N_14041,N_13775,N_13850);
or U14042 (N_14042,N_13913,N_13784);
xor U14043 (N_14043,N_13826,N_13892);
or U14044 (N_14044,N_13764,N_13772);
and U14045 (N_14045,N_13898,N_13815);
or U14046 (N_14046,N_13781,N_13854);
nand U14047 (N_14047,N_13863,N_13793);
and U14048 (N_14048,N_13868,N_13807);
or U14049 (N_14049,N_13851,N_13876);
nor U14050 (N_14050,N_13791,N_13891);
nand U14051 (N_14051,N_13819,N_13875);
xor U14052 (N_14052,N_13786,N_13762);
xor U14053 (N_14053,N_13895,N_13760);
nand U14054 (N_14054,N_13902,N_13828);
xor U14055 (N_14055,N_13834,N_13853);
xor U14056 (N_14056,N_13779,N_13909);
xor U14057 (N_14057,N_13788,N_13890);
nor U14058 (N_14058,N_13912,N_13897);
and U14059 (N_14059,N_13794,N_13914);
nor U14060 (N_14060,N_13912,N_13836);
nand U14061 (N_14061,N_13894,N_13849);
xor U14062 (N_14062,N_13819,N_13843);
or U14063 (N_14063,N_13904,N_13914);
or U14064 (N_14064,N_13791,N_13784);
and U14065 (N_14065,N_13883,N_13880);
xnor U14066 (N_14066,N_13845,N_13777);
or U14067 (N_14067,N_13902,N_13824);
and U14068 (N_14068,N_13829,N_13913);
and U14069 (N_14069,N_13849,N_13787);
nand U14070 (N_14070,N_13911,N_13802);
or U14071 (N_14071,N_13837,N_13836);
or U14072 (N_14072,N_13845,N_13826);
xor U14073 (N_14073,N_13897,N_13820);
nand U14074 (N_14074,N_13915,N_13864);
nand U14075 (N_14075,N_13861,N_13810);
or U14076 (N_14076,N_13795,N_13820);
xnor U14077 (N_14077,N_13761,N_13778);
nand U14078 (N_14078,N_13858,N_13830);
xnor U14079 (N_14079,N_13842,N_13908);
nand U14080 (N_14080,N_14067,N_13927);
xnor U14081 (N_14081,N_14006,N_14075);
nand U14082 (N_14082,N_13924,N_14073);
xor U14083 (N_14083,N_14061,N_13967);
and U14084 (N_14084,N_14029,N_13979);
xor U14085 (N_14085,N_13998,N_14017);
nand U14086 (N_14086,N_13984,N_14036);
nor U14087 (N_14087,N_14062,N_14039);
nor U14088 (N_14088,N_14070,N_13943);
nor U14089 (N_14089,N_14027,N_13997);
xor U14090 (N_14090,N_14026,N_14009);
xor U14091 (N_14091,N_13937,N_13964);
nor U14092 (N_14092,N_14045,N_14037);
and U14093 (N_14093,N_13951,N_13952);
or U14094 (N_14094,N_14044,N_14066);
xnor U14095 (N_14095,N_14005,N_13935);
xnor U14096 (N_14096,N_13978,N_14031);
or U14097 (N_14097,N_13988,N_13939);
xor U14098 (N_14098,N_13940,N_14003);
nand U14099 (N_14099,N_14065,N_14025);
or U14100 (N_14100,N_13932,N_14016);
xor U14101 (N_14101,N_14004,N_14000);
or U14102 (N_14102,N_14057,N_13921);
or U14103 (N_14103,N_14068,N_13972);
nand U14104 (N_14104,N_14058,N_13945);
and U14105 (N_14105,N_13980,N_14072);
nand U14106 (N_14106,N_14040,N_14022);
or U14107 (N_14107,N_13962,N_14043);
xor U14108 (N_14108,N_14020,N_13969);
nor U14109 (N_14109,N_13987,N_14069);
or U14110 (N_14110,N_13983,N_14013);
or U14111 (N_14111,N_13966,N_13993);
nand U14112 (N_14112,N_13973,N_14010);
and U14113 (N_14113,N_13938,N_14055);
xor U14114 (N_14114,N_14063,N_13958);
nor U14115 (N_14115,N_14001,N_13928);
xor U14116 (N_14116,N_13934,N_14028);
xor U14117 (N_14117,N_14012,N_13959);
and U14118 (N_14118,N_13981,N_13991);
nor U14119 (N_14119,N_13968,N_13941);
xor U14120 (N_14120,N_13996,N_13965);
or U14121 (N_14121,N_13986,N_14011);
nor U14122 (N_14122,N_13930,N_13953);
nor U14123 (N_14123,N_13944,N_13925);
nand U14124 (N_14124,N_13922,N_13961);
nor U14125 (N_14125,N_13975,N_13946);
nand U14126 (N_14126,N_13957,N_14007);
and U14127 (N_14127,N_14079,N_13926);
and U14128 (N_14128,N_13950,N_13999);
xor U14129 (N_14129,N_14023,N_13936);
nand U14130 (N_14130,N_14035,N_13923);
nor U14131 (N_14131,N_14019,N_13955);
xor U14132 (N_14132,N_14078,N_13929);
nand U14133 (N_14133,N_14018,N_14048);
and U14134 (N_14134,N_13994,N_14033);
nor U14135 (N_14135,N_14064,N_13977);
nor U14136 (N_14136,N_13942,N_14002);
nor U14137 (N_14137,N_14024,N_14074);
nor U14138 (N_14138,N_13982,N_14034);
xnor U14139 (N_14139,N_13947,N_14076);
nand U14140 (N_14140,N_14047,N_13971);
or U14141 (N_14141,N_14021,N_13956);
nor U14142 (N_14142,N_14059,N_13974);
and U14143 (N_14143,N_14051,N_14014);
or U14144 (N_14144,N_13931,N_14052);
xnor U14145 (N_14145,N_13963,N_14050);
and U14146 (N_14146,N_14032,N_14030);
and U14147 (N_14147,N_13949,N_14041);
and U14148 (N_14148,N_13954,N_14008);
xor U14149 (N_14149,N_14049,N_14053);
and U14150 (N_14150,N_14054,N_14015);
nand U14151 (N_14151,N_13992,N_13960);
nor U14152 (N_14152,N_13920,N_14071);
nand U14153 (N_14153,N_14077,N_13970);
xnor U14154 (N_14154,N_14056,N_13948);
xnor U14155 (N_14155,N_13990,N_13995);
nand U14156 (N_14156,N_14042,N_13989);
nor U14157 (N_14157,N_14038,N_14046);
and U14158 (N_14158,N_13985,N_14060);
xor U14159 (N_14159,N_13933,N_13976);
and U14160 (N_14160,N_14053,N_13923);
nor U14161 (N_14161,N_14028,N_14061);
nor U14162 (N_14162,N_13932,N_14073);
nor U14163 (N_14163,N_14014,N_13951);
nand U14164 (N_14164,N_14072,N_13949);
and U14165 (N_14165,N_14006,N_14008);
nand U14166 (N_14166,N_14073,N_14064);
nand U14167 (N_14167,N_13968,N_14062);
or U14168 (N_14168,N_14020,N_13991);
and U14169 (N_14169,N_13994,N_13956);
and U14170 (N_14170,N_13932,N_14046);
nor U14171 (N_14171,N_13944,N_13974);
nor U14172 (N_14172,N_13959,N_14018);
xnor U14173 (N_14173,N_13941,N_14010);
nand U14174 (N_14174,N_14004,N_14056);
or U14175 (N_14175,N_13989,N_13956);
xor U14176 (N_14176,N_14025,N_13995);
xnor U14177 (N_14177,N_14029,N_13976);
xnor U14178 (N_14178,N_13981,N_14007);
nor U14179 (N_14179,N_14079,N_14050);
nor U14180 (N_14180,N_13991,N_14076);
and U14181 (N_14181,N_13929,N_13988);
or U14182 (N_14182,N_14035,N_13962);
and U14183 (N_14183,N_14074,N_14056);
xnor U14184 (N_14184,N_13972,N_13924);
and U14185 (N_14185,N_13992,N_14013);
xor U14186 (N_14186,N_13969,N_14046);
nand U14187 (N_14187,N_13966,N_14010);
or U14188 (N_14188,N_13953,N_14060);
nand U14189 (N_14189,N_14050,N_13941);
nor U14190 (N_14190,N_13937,N_13921);
xor U14191 (N_14191,N_13986,N_14037);
xnor U14192 (N_14192,N_14030,N_14057);
or U14193 (N_14193,N_14047,N_14020);
and U14194 (N_14194,N_13933,N_13927);
nand U14195 (N_14195,N_13963,N_14067);
nand U14196 (N_14196,N_14067,N_13955);
nor U14197 (N_14197,N_14005,N_13934);
nand U14198 (N_14198,N_14025,N_13994);
nor U14199 (N_14199,N_14043,N_13988);
nor U14200 (N_14200,N_13985,N_13968);
nor U14201 (N_14201,N_13997,N_13971);
and U14202 (N_14202,N_13974,N_14006);
and U14203 (N_14203,N_13930,N_13992);
nand U14204 (N_14204,N_13924,N_13988);
nand U14205 (N_14205,N_13979,N_13968);
xor U14206 (N_14206,N_13949,N_14034);
and U14207 (N_14207,N_13987,N_13945);
nor U14208 (N_14208,N_14035,N_14072);
or U14209 (N_14209,N_14009,N_14039);
nor U14210 (N_14210,N_14009,N_13925);
and U14211 (N_14211,N_13963,N_14073);
or U14212 (N_14212,N_13930,N_14072);
nand U14213 (N_14213,N_14024,N_13942);
or U14214 (N_14214,N_13963,N_14012);
nand U14215 (N_14215,N_14053,N_13991);
nor U14216 (N_14216,N_13964,N_13945);
nor U14217 (N_14217,N_14021,N_13988);
nand U14218 (N_14218,N_14010,N_13949);
and U14219 (N_14219,N_14019,N_14012);
and U14220 (N_14220,N_14024,N_13995);
nand U14221 (N_14221,N_14043,N_14006);
nor U14222 (N_14222,N_14070,N_14010);
and U14223 (N_14223,N_14003,N_13961);
nor U14224 (N_14224,N_14047,N_13970);
nor U14225 (N_14225,N_13970,N_13961);
or U14226 (N_14226,N_13993,N_14062);
and U14227 (N_14227,N_14036,N_13960);
xor U14228 (N_14228,N_13998,N_13984);
nor U14229 (N_14229,N_14031,N_14003);
xor U14230 (N_14230,N_14060,N_14062);
xnor U14231 (N_14231,N_14053,N_14037);
xor U14232 (N_14232,N_13956,N_14050);
nand U14233 (N_14233,N_13971,N_14035);
nand U14234 (N_14234,N_13994,N_13984);
or U14235 (N_14235,N_13976,N_14046);
nand U14236 (N_14236,N_14010,N_13980);
nand U14237 (N_14237,N_14052,N_14000);
xnor U14238 (N_14238,N_14041,N_14010);
or U14239 (N_14239,N_13985,N_13925);
or U14240 (N_14240,N_14172,N_14198);
or U14241 (N_14241,N_14201,N_14167);
and U14242 (N_14242,N_14139,N_14118);
and U14243 (N_14243,N_14238,N_14227);
or U14244 (N_14244,N_14206,N_14181);
xnor U14245 (N_14245,N_14123,N_14218);
or U14246 (N_14246,N_14237,N_14086);
and U14247 (N_14247,N_14203,N_14222);
nand U14248 (N_14248,N_14131,N_14183);
xnor U14249 (N_14249,N_14213,N_14124);
xnor U14250 (N_14250,N_14192,N_14148);
or U14251 (N_14251,N_14169,N_14219);
nor U14252 (N_14252,N_14158,N_14157);
xor U14253 (N_14253,N_14239,N_14221);
nor U14254 (N_14254,N_14188,N_14128);
and U14255 (N_14255,N_14120,N_14101);
nand U14256 (N_14256,N_14085,N_14164);
nand U14257 (N_14257,N_14134,N_14080);
xor U14258 (N_14258,N_14092,N_14230);
nand U14259 (N_14259,N_14149,N_14145);
nor U14260 (N_14260,N_14187,N_14116);
nor U14261 (N_14261,N_14212,N_14153);
nor U14262 (N_14262,N_14178,N_14174);
xor U14263 (N_14263,N_14171,N_14126);
xnor U14264 (N_14264,N_14205,N_14229);
or U14265 (N_14265,N_14224,N_14106);
nand U14266 (N_14266,N_14179,N_14210);
nand U14267 (N_14267,N_14163,N_14108);
xnor U14268 (N_14268,N_14127,N_14235);
nor U14269 (N_14269,N_14095,N_14132);
xor U14270 (N_14270,N_14115,N_14119);
nor U14271 (N_14271,N_14236,N_14091);
and U14272 (N_14272,N_14193,N_14105);
xnor U14273 (N_14273,N_14215,N_14090);
nand U14274 (N_14274,N_14110,N_14113);
nor U14275 (N_14275,N_14151,N_14098);
nand U14276 (N_14276,N_14159,N_14234);
xnor U14277 (N_14277,N_14112,N_14209);
xor U14278 (N_14278,N_14087,N_14117);
or U14279 (N_14279,N_14084,N_14141);
nand U14280 (N_14280,N_14114,N_14088);
nor U14281 (N_14281,N_14082,N_14096);
nand U14282 (N_14282,N_14161,N_14223);
and U14283 (N_14283,N_14100,N_14190);
nor U14284 (N_14284,N_14177,N_14160);
and U14285 (N_14285,N_14099,N_14097);
nor U14286 (N_14286,N_14226,N_14137);
nor U14287 (N_14287,N_14156,N_14103);
and U14288 (N_14288,N_14152,N_14173);
or U14289 (N_14289,N_14143,N_14217);
or U14290 (N_14290,N_14136,N_14155);
xnor U14291 (N_14291,N_14165,N_14083);
or U14292 (N_14292,N_14199,N_14191);
or U14293 (N_14293,N_14202,N_14166);
nand U14294 (N_14294,N_14228,N_14204);
or U14295 (N_14295,N_14189,N_14184);
or U14296 (N_14296,N_14233,N_14130);
xor U14297 (N_14297,N_14081,N_14207);
and U14298 (N_14298,N_14109,N_14231);
and U14299 (N_14299,N_14122,N_14211);
nand U14300 (N_14300,N_14225,N_14176);
xnor U14301 (N_14301,N_14093,N_14144);
and U14302 (N_14302,N_14194,N_14182);
nand U14303 (N_14303,N_14142,N_14138);
nor U14304 (N_14304,N_14107,N_14168);
or U14305 (N_14305,N_14135,N_14162);
nand U14306 (N_14306,N_14214,N_14175);
and U14307 (N_14307,N_14133,N_14129);
or U14308 (N_14308,N_14185,N_14125);
or U14309 (N_14309,N_14180,N_14216);
nor U14310 (N_14310,N_14146,N_14197);
and U14311 (N_14311,N_14140,N_14104);
and U14312 (N_14312,N_14195,N_14121);
nor U14313 (N_14313,N_14232,N_14154);
or U14314 (N_14314,N_14196,N_14089);
nor U14315 (N_14315,N_14150,N_14170);
nor U14316 (N_14316,N_14094,N_14186);
nor U14317 (N_14317,N_14208,N_14111);
nor U14318 (N_14318,N_14102,N_14200);
xor U14319 (N_14319,N_14147,N_14220);
nor U14320 (N_14320,N_14216,N_14140);
or U14321 (N_14321,N_14125,N_14082);
nand U14322 (N_14322,N_14101,N_14164);
or U14323 (N_14323,N_14203,N_14130);
nor U14324 (N_14324,N_14158,N_14235);
xor U14325 (N_14325,N_14137,N_14230);
nand U14326 (N_14326,N_14193,N_14205);
xnor U14327 (N_14327,N_14092,N_14145);
nand U14328 (N_14328,N_14223,N_14231);
and U14329 (N_14329,N_14148,N_14190);
or U14330 (N_14330,N_14084,N_14114);
or U14331 (N_14331,N_14099,N_14095);
nand U14332 (N_14332,N_14235,N_14199);
xor U14333 (N_14333,N_14225,N_14093);
or U14334 (N_14334,N_14114,N_14097);
and U14335 (N_14335,N_14164,N_14215);
xnor U14336 (N_14336,N_14167,N_14207);
or U14337 (N_14337,N_14150,N_14100);
xor U14338 (N_14338,N_14229,N_14132);
and U14339 (N_14339,N_14093,N_14084);
xnor U14340 (N_14340,N_14101,N_14146);
nand U14341 (N_14341,N_14080,N_14205);
or U14342 (N_14342,N_14165,N_14186);
and U14343 (N_14343,N_14214,N_14138);
and U14344 (N_14344,N_14127,N_14222);
nor U14345 (N_14345,N_14165,N_14171);
or U14346 (N_14346,N_14098,N_14083);
nor U14347 (N_14347,N_14155,N_14149);
and U14348 (N_14348,N_14132,N_14143);
nor U14349 (N_14349,N_14087,N_14123);
and U14350 (N_14350,N_14178,N_14107);
nor U14351 (N_14351,N_14174,N_14168);
and U14352 (N_14352,N_14120,N_14150);
nand U14353 (N_14353,N_14167,N_14220);
or U14354 (N_14354,N_14193,N_14204);
nor U14355 (N_14355,N_14229,N_14210);
and U14356 (N_14356,N_14144,N_14083);
nor U14357 (N_14357,N_14196,N_14096);
xor U14358 (N_14358,N_14237,N_14214);
xnor U14359 (N_14359,N_14169,N_14199);
or U14360 (N_14360,N_14187,N_14167);
nand U14361 (N_14361,N_14222,N_14206);
and U14362 (N_14362,N_14162,N_14238);
or U14363 (N_14363,N_14110,N_14202);
xnor U14364 (N_14364,N_14104,N_14222);
or U14365 (N_14365,N_14208,N_14195);
or U14366 (N_14366,N_14226,N_14104);
xor U14367 (N_14367,N_14197,N_14081);
or U14368 (N_14368,N_14161,N_14194);
xor U14369 (N_14369,N_14175,N_14202);
nor U14370 (N_14370,N_14090,N_14112);
and U14371 (N_14371,N_14186,N_14223);
nand U14372 (N_14372,N_14152,N_14181);
or U14373 (N_14373,N_14084,N_14230);
nand U14374 (N_14374,N_14220,N_14106);
xor U14375 (N_14375,N_14129,N_14213);
nor U14376 (N_14376,N_14096,N_14090);
nor U14377 (N_14377,N_14169,N_14151);
and U14378 (N_14378,N_14170,N_14227);
or U14379 (N_14379,N_14239,N_14117);
xnor U14380 (N_14380,N_14142,N_14213);
nand U14381 (N_14381,N_14099,N_14209);
or U14382 (N_14382,N_14199,N_14187);
nand U14383 (N_14383,N_14221,N_14217);
nand U14384 (N_14384,N_14085,N_14215);
or U14385 (N_14385,N_14221,N_14137);
or U14386 (N_14386,N_14130,N_14168);
nor U14387 (N_14387,N_14143,N_14145);
and U14388 (N_14388,N_14226,N_14191);
xnor U14389 (N_14389,N_14100,N_14234);
xor U14390 (N_14390,N_14212,N_14221);
nand U14391 (N_14391,N_14234,N_14102);
and U14392 (N_14392,N_14228,N_14132);
nand U14393 (N_14393,N_14223,N_14119);
xnor U14394 (N_14394,N_14174,N_14213);
or U14395 (N_14395,N_14088,N_14185);
xnor U14396 (N_14396,N_14133,N_14104);
xor U14397 (N_14397,N_14232,N_14201);
or U14398 (N_14398,N_14205,N_14110);
xor U14399 (N_14399,N_14170,N_14165);
nor U14400 (N_14400,N_14311,N_14302);
xnor U14401 (N_14401,N_14268,N_14252);
or U14402 (N_14402,N_14299,N_14366);
nor U14403 (N_14403,N_14258,N_14261);
and U14404 (N_14404,N_14384,N_14244);
nand U14405 (N_14405,N_14246,N_14391);
or U14406 (N_14406,N_14398,N_14367);
nor U14407 (N_14407,N_14313,N_14322);
or U14408 (N_14408,N_14285,N_14346);
nand U14409 (N_14409,N_14308,N_14396);
xnor U14410 (N_14410,N_14303,N_14377);
and U14411 (N_14411,N_14245,N_14343);
and U14412 (N_14412,N_14386,N_14354);
nor U14413 (N_14413,N_14341,N_14318);
or U14414 (N_14414,N_14369,N_14390);
nor U14415 (N_14415,N_14315,N_14266);
nor U14416 (N_14416,N_14375,N_14382);
nor U14417 (N_14417,N_14286,N_14321);
or U14418 (N_14418,N_14264,N_14290);
and U14419 (N_14419,N_14278,N_14277);
and U14420 (N_14420,N_14339,N_14304);
and U14421 (N_14421,N_14371,N_14338);
or U14422 (N_14422,N_14323,N_14262);
and U14423 (N_14423,N_14353,N_14392);
and U14424 (N_14424,N_14331,N_14325);
or U14425 (N_14425,N_14309,N_14280);
xor U14426 (N_14426,N_14281,N_14360);
xnor U14427 (N_14427,N_14256,N_14255);
and U14428 (N_14428,N_14342,N_14276);
and U14429 (N_14429,N_14329,N_14296);
nand U14430 (N_14430,N_14379,N_14373);
xor U14431 (N_14431,N_14389,N_14388);
xor U14432 (N_14432,N_14399,N_14279);
nor U14433 (N_14433,N_14283,N_14327);
xnor U14434 (N_14434,N_14293,N_14269);
nor U14435 (N_14435,N_14365,N_14272);
or U14436 (N_14436,N_14328,N_14270);
nor U14437 (N_14437,N_14330,N_14305);
and U14438 (N_14438,N_14297,N_14291);
nor U14439 (N_14439,N_14372,N_14242);
nand U14440 (N_14440,N_14292,N_14385);
nand U14441 (N_14441,N_14394,N_14294);
or U14442 (N_14442,N_14250,N_14254);
nand U14443 (N_14443,N_14301,N_14345);
and U14444 (N_14444,N_14306,N_14348);
nand U14445 (N_14445,N_14320,N_14350);
or U14446 (N_14446,N_14312,N_14307);
and U14447 (N_14447,N_14374,N_14380);
nor U14448 (N_14448,N_14317,N_14257);
xor U14449 (N_14449,N_14295,N_14326);
nor U14450 (N_14450,N_14359,N_14259);
nor U14451 (N_14451,N_14247,N_14361);
and U14452 (N_14452,N_14378,N_14273);
xor U14453 (N_14453,N_14243,N_14282);
xor U14454 (N_14454,N_14351,N_14289);
nand U14455 (N_14455,N_14368,N_14275);
xor U14456 (N_14456,N_14319,N_14383);
nor U14457 (N_14457,N_14333,N_14334);
and U14458 (N_14458,N_14253,N_14387);
and U14459 (N_14459,N_14355,N_14340);
xnor U14460 (N_14460,N_14241,N_14265);
nand U14461 (N_14461,N_14381,N_14248);
or U14462 (N_14462,N_14362,N_14344);
and U14463 (N_14463,N_14284,N_14310);
and U14464 (N_14464,N_14352,N_14274);
or U14465 (N_14465,N_14240,N_14370);
xor U14466 (N_14466,N_14267,N_14314);
and U14467 (N_14467,N_14287,N_14251);
nor U14468 (N_14468,N_14336,N_14337);
nor U14469 (N_14469,N_14335,N_14260);
and U14470 (N_14470,N_14356,N_14316);
or U14471 (N_14471,N_14332,N_14271);
or U14472 (N_14472,N_14358,N_14249);
nand U14473 (N_14473,N_14300,N_14357);
nor U14474 (N_14474,N_14288,N_14364);
xor U14475 (N_14475,N_14263,N_14363);
xor U14476 (N_14476,N_14376,N_14397);
and U14477 (N_14477,N_14393,N_14298);
xor U14478 (N_14478,N_14349,N_14347);
xor U14479 (N_14479,N_14324,N_14395);
or U14480 (N_14480,N_14394,N_14380);
nor U14481 (N_14481,N_14394,N_14248);
nor U14482 (N_14482,N_14379,N_14287);
nor U14483 (N_14483,N_14380,N_14301);
and U14484 (N_14484,N_14344,N_14375);
nand U14485 (N_14485,N_14355,N_14373);
xor U14486 (N_14486,N_14244,N_14383);
and U14487 (N_14487,N_14295,N_14399);
nor U14488 (N_14488,N_14266,N_14380);
or U14489 (N_14489,N_14289,N_14260);
or U14490 (N_14490,N_14259,N_14269);
xor U14491 (N_14491,N_14274,N_14315);
xnor U14492 (N_14492,N_14293,N_14246);
or U14493 (N_14493,N_14241,N_14358);
nand U14494 (N_14494,N_14392,N_14341);
nor U14495 (N_14495,N_14293,N_14329);
xor U14496 (N_14496,N_14356,N_14306);
and U14497 (N_14497,N_14263,N_14354);
nor U14498 (N_14498,N_14326,N_14277);
xnor U14499 (N_14499,N_14302,N_14305);
xnor U14500 (N_14500,N_14245,N_14377);
and U14501 (N_14501,N_14270,N_14298);
or U14502 (N_14502,N_14266,N_14366);
nor U14503 (N_14503,N_14339,N_14343);
nand U14504 (N_14504,N_14327,N_14282);
nor U14505 (N_14505,N_14399,N_14315);
nand U14506 (N_14506,N_14317,N_14286);
xnor U14507 (N_14507,N_14389,N_14262);
nor U14508 (N_14508,N_14259,N_14368);
xor U14509 (N_14509,N_14255,N_14248);
nand U14510 (N_14510,N_14325,N_14281);
xor U14511 (N_14511,N_14343,N_14259);
xnor U14512 (N_14512,N_14257,N_14353);
nor U14513 (N_14513,N_14353,N_14326);
and U14514 (N_14514,N_14243,N_14381);
nand U14515 (N_14515,N_14333,N_14252);
and U14516 (N_14516,N_14292,N_14243);
nor U14517 (N_14517,N_14286,N_14373);
xnor U14518 (N_14518,N_14281,N_14277);
nor U14519 (N_14519,N_14359,N_14348);
and U14520 (N_14520,N_14383,N_14357);
and U14521 (N_14521,N_14396,N_14345);
xnor U14522 (N_14522,N_14291,N_14364);
or U14523 (N_14523,N_14392,N_14390);
nor U14524 (N_14524,N_14256,N_14384);
xor U14525 (N_14525,N_14375,N_14308);
and U14526 (N_14526,N_14350,N_14282);
xnor U14527 (N_14527,N_14298,N_14374);
nor U14528 (N_14528,N_14344,N_14259);
nor U14529 (N_14529,N_14309,N_14386);
nor U14530 (N_14530,N_14269,N_14279);
nand U14531 (N_14531,N_14340,N_14319);
nor U14532 (N_14532,N_14295,N_14388);
xnor U14533 (N_14533,N_14369,N_14240);
and U14534 (N_14534,N_14292,N_14257);
nand U14535 (N_14535,N_14270,N_14260);
nor U14536 (N_14536,N_14264,N_14349);
and U14537 (N_14537,N_14282,N_14345);
or U14538 (N_14538,N_14298,N_14247);
and U14539 (N_14539,N_14395,N_14275);
xor U14540 (N_14540,N_14246,N_14299);
nand U14541 (N_14541,N_14268,N_14389);
nand U14542 (N_14542,N_14259,N_14374);
nor U14543 (N_14543,N_14317,N_14301);
and U14544 (N_14544,N_14307,N_14263);
nand U14545 (N_14545,N_14356,N_14377);
xor U14546 (N_14546,N_14263,N_14294);
xor U14547 (N_14547,N_14280,N_14327);
xor U14548 (N_14548,N_14255,N_14378);
nor U14549 (N_14549,N_14319,N_14356);
nand U14550 (N_14550,N_14265,N_14347);
and U14551 (N_14551,N_14392,N_14362);
or U14552 (N_14552,N_14361,N_14245);
nand U14553 (N_14553,N_14340,N_14333);
or U14554 (N_14554,N_14313,N_14347);
nor U14555 (N_14555,N_14361,N_14249);
or U14556 (N_14556,N_14383,N_14358);
nand U14557 (N_14557,N_14312,N_14324);
and U14558 (N_14558,N_14369,N_14336);
or U14559 (N_14559,N_14281,N_14327);
xor U14560 (N_14560,N_14511,N_14535);
or U14561 (N_14561,N_14405,N_14400);
nor U14562 (N_14562,N_14502,N_14411);
and U14563 (N_14563,N_14525,N_14495);
nor U14564 (N_14564,N_14509,N_14449);
or U14565 (N_14565,N_14413,N_14516);
and U14566 (N_14566,N_14455,N_14542);
and U14567 (N_14567,N_14540,N_14483);
xnor U14568 (N_14568,N_14425,N_14503);
nand U14569 (N_14569,N_14420,N_14491);
or U14570 (N_14570,N_14510,N_14485);
nand U14571 (N_14571,N_14518,N_14472);
nand U14572 (N_14572,N_14436,N_14528);
and U14573 (N_14573,N_14498,N_14532);
nor U14574 (N_14574,N_14442,N_14433);
and U14575 (N_14575,N_14484,N_14448);
nand U14576 (N_14576,N_14427,N_14429);
and U14577 (N_14577,N_14408,N_14454);
nand U14578 (N_14578,N_14521,N_14551);
nand U14579 (N_14579,N_14554,N_14437);
and U14580 (N_14580,N_14496,N_14479);
nor U14581 (N_14581,N_14407,N_14468);
and U14582 (N_14582,N_14499,N_14545);
nand U14583 (N_14583,N_14506,N_14515);
xnor U14584 (N_14584,N_14497,N_14475);
and U14585 (N_14585,N_14536,N_14558);
nand U14586 (N_14586,N_14533,N_14527);
and U14587 (N_14587,N_14410,N_14401);
xnor U14588 (N_14588,N_14412,N_14451);
nand U14589 (N_14589,N_14466,N_14463);
and U14590 (N_14590,N_14476,N_14546);
or U14591 (N_14591,N_14488,N_14526);
or U14592 (N_14592,N_14460,N_14461);
nand U14593 (N_14593,N_14409,N_14553);
or U14594 (N_14594,N_14416,N_14406);
or U14595 (N_14595,N_14555,N_14426);
xor U14596 (N_14596,N_14493,N_14492);
nand U14597 (N_14597,N_14477,N_14529);
nand U14598 (N_14598,N_14441,N_14444);
or U14599 (N_14599,N_14539,N_14524);
nor U14600 (N_14600,N_14487,N_14470);
nor U14601 (N_14601,N_14469,N_14538);
or U14602 (N_14602,N_14514,N_14435);
or U14603 (N_14603,N_14467,N_14462);
nand U14604 (N_14604,N_14486,N_14523);
nor U14605 (N_14605,N_14458,N_14445);
nand U14606 (N_14606,N_14517,N_14443);
and U14607 (N_14607,N_14531,N_14402);
nand U14608 (N_14608,N_14559,N_14422);
nand U14609 (N_14609,N_14430,N_14431);
nor U14610 (N_14610,N_14440,N_14534);
and U14611 (N_14611,N_14415,N_14417);
nand U14612 (N_14612,N_14480,N_14403);
nor U14613 (N_14613,N_14482,N_14423);
or U14614 (N_14614,N_14456,N_14543);
nor U14615 (N_14615,N_14452,N_14522);
and U14616 (N_14616,N_14519,N_14494);
or U14617 (N_14617,N_14453,N_14548);
nand U14618 (N_14618,N_14520,N_14537);
nand U14619 (N_14619,N_14457,N_14428);
and U14620 (N_14620,N_14464,N_14552);
nand U14621 (N_14621,N_14504,N_14471);
nand U14622 (N_14622,N_14500,N_14547);
or U14623 (N_14623,N_14513,N_14512);
xnor U14624 (N_14624,N_14418,N_14505);
or U14625 (N_14625,N_14414,N_14481);
and U14626 (N_14626,N_14501,N_14438);
nor U14627 (N_14627,N_14465,N_14556);
nand U14628 (N_14628,N_14549,N_14473);
xnor U14629 (N_14629,N_14550,N_14419);
xor U14630 (N_14630,N_14421,N_14459);
nand U14631 (N_14631,N_14508,N_14490);
xor U14632 (N_14632,N_14404,N_14530);
xor U14633 (N_14633,N_14507,N_14447);
and U14634 (N_14634,N_14489,N_14446);
xnor U14635 (N_14635,N_14432,N_14541);
and U14636 (N_14636,N_14434,N_14474);
nand U14637 (N_14637,N_14544,N_14424);
nand U14638 (N_14638,N_14450,N_14557);
and U14639 (N_14639,N_14478,N_14439);
nand U14640 (N_14640,N_14513,N_14457);
and U14641 (N_14641,N_14502,N_14508);
nand U14642 (N_14642,N_14508,N_14476);
nand U14643 (N_14643,N_14528,N_14549);
and U14644 (N_14644,N_14497,N_14408);
or U14645 (N_14645,N_14531,N_14539);
nor U14646 (N_14646,N_14424,N_14413);
nor U14647 (N_14647,N_14480,N_14466);
xnor U14648 (N_14648,N_14477,N_14548);
nor U14649 (N_14649,N_14526,N_14429);
nor U14650 (N_14650,N_14430,N_14488);
or U14651 (N_14651,N_14486,N_14402);
nand U14652 (N_14652,N_14402,N_14494);
nor U14653 (N_14653,N_14505,N_14541);
xnor U14654 (N_14654,N_14478,N_14485);
and U14655 (N_14655,N_14524,N_14426);
and U14656 (N_14656,N_14554,N_14461);
nor U14657 (N_14657,N_14443,N_14504);
or U14658 (N_14658,N_14432,N_14408);
nand U14659 (N_14659,N_14405,N_14453);
nor U14660 (N_14660,N_14486,N_14488);
xnor U14661 (N_14661,N_14514,N_14429);
nand U14662 (N_14662,N_14414,N_14437);
nor U14663 (N_14663,N_14467,N_14552);
or U14664 (N_14664,N_14541,N_14509);
and U14665 (N_14665,N_14509,N_14463);
and U14666 (N_14666,N_14404,N_14408);
nor U14667 (N_14667,N_14401,N_14478);
and U14668 (N_14668,N_14551,N_14419);
nor U14669 (N_14669,N_14496,N_14525);
and U14670 (N_14670,N_14481,N_14434);
or U14671 (N_14671,N_14412,N_14464);
xor U14672 (N_14672,N_14541,N_14473);
or U14673 (N_14673,N_14439,N_14547);
and U14674 (N_14674,N_14529,N_14432);
and U14675 (N_14675,N_14471,N_14411);
or U14676 (N_14676,N_14431,N_14434);
xor U14677 (N_14677,N_14437,N_14534);
nand U14678 (N_14678,N_14530,N_14420);
nor U14679 (N_14679,N_14422,N_14426);
nand U14680 (N_14680,N_14522,N_14441);
or U14681 (N_14681,N_14497,N_14545);
nand U14682 (N_14682,N_14515,N_14521);
or U14683 (N_14683,N_14475,N_14501);
xor U14684 (N_14684,N_14525,N_14549);
nand U14685 (N_14685,N_14526,N_14535);
xor U14686 (N_14686,N_14548,N_14551);
and U14687 (N_14687,N_14513,N_14501);
or U14688 (N_14688,N_14442,N_14539);
nand U14689 (N_14689,N_14415,N_14508);
and U14690 (N_14690,N_14490,N_14515);
and U14691 (N_14691,N_14522,N_14440);
nor U14692 (N_14692,N_14536,N_14462);
or U14693 (N_14693,N_14526,N_14546);
nand U14694 (N_14694,N_14536,N_14479);
or U14695 (N_14695,N_14520,N_14548);
or U14696 (N_14696,N_14474,N_14554);
or U14697 (N_14697,N_14415,N_14544);
nand U14698 (N_14698,N_14404,N_14518);
nand U14699 (N_14699,N_14466,N_14460);
or U14700 (N_14700,N_14403,N_14542);
nor U14701 (N_14701,N_14538,N_14418);
or U14702 (N_14702,N_14423,N_14526);
and U14703 (N_14703,N_14425,N_14525);
or U14704 (N_14704,N_14454,N_14503);
and U14705 (N_14705,N_14409,N_14426);
or U14706 (N_14706,N_14448,N_14426);
xor U14707 (N_14707,N_14419,N_14521);
nor U14708 (N_14708,N_14469,N_14449);
xnor U14709 (N_14709,N_14502,N_14504);
nand U14710 (N_14710,N_14409,N_14420);
xnor U14711 (N_14711,N_14559,N_14461);
nand U14712 (N_14712,N_14408,N_14449);
nand U14713 (N_14713,N_14430,N_14458);
nor U14714 (N_14714,N_14485,N_14539);
nor U14715 (N_14715,N_14549,N_14469);
or U14716 (N_14716,N_14513,N_14463);
xnor U14717 (N_14717,N_14489,N_14467);
xnor U14718 (N_14718,N_14545,N_14445);
nor U14719 (N_14719,N_14495,N_14454);
nand U14720 (N_14720,N_14624,N_14715);
or U14721 (N_14721,N_14587,N_14712);
nor U14722 (N_14722,N_14679,N_14704);
xnor U14723 (N_14723,N_14643,N_14631);
nor U14724 (N_14724,N_14687,N_14669);
or U14725 (N_14725,N_14586,N_14597);
or U14726 (N_14726,N_14700,N_14705);
xnor U14727 (N_14727,N_14697,N_14717);
or U14728 (N_14728,N_14634,N_14571);
or U14729 (N_14729,N_14567,N_14668);
xor U14730 (N_14730,N_14646,N_14616);
and U14731 (N_14731,N_14692,N_14657);
nor U14732 (N_14732,N_14607,N_14645);
nor U14733 (N_14733,N_14699,N_14610);
and U14734 (N_14734,N_14676,N_14653);
nand U14735 (N_14735,N_14606,N_14652);
and U14736 (N_14736,N_14590,N_14633);
xnor U14737 (N_14737,N_14570,N_14600);
xnor U14738 (N_14738,N_14703,N_14661);
xor U14739 (N_14739,N_14589,N_14591);
or U14740 (N_14740,N_14560,N_14648);
xnor U14741 (N_14741,N_14581,N_14663);
xnor U14742 (N_14742,N_14611,N_14626);
or U14743 (N_14743,N_14632,N_14706);
nor U14744 (N_14744,N_14622,N_14592);
xor U14745 (N_14745,N_14662,N_14671);
nor U14746 (N_14746,N_14566,N_14714);
xnor U14747 (N_14747,N_14674,N_14677);
xnor U14748 (N_14748,N_14609,N_14627);
and U14749 (N_14749,N_14672,N_14628);
xor U14750 (N_14750,N_14576,N_14686);
nor U14751 (N_14751,N_14564,N_14650);
nand U14752 (N_14752,N_14618,N_14693);
nor U14753 (N_14753,N_14639,N_14695);
or U14754 (N_14754,N_14635,N_14637);
xnor U14755 (N_14755,N_14574,N_14630);
and U14756 (N_14756,N_14608,N_14573);
xnor U14757 (N_14757,N_14649,N_14593);
or U14758 (N_14758,N_14580,N_14654);
nor U14759 (N_14759,N_14602,N_14615);
and U14760 (N_14760,N_14613,N_14579);
or U14761 (N_14761,N_14667,N_14660);
or U14762 (N_14762,N_14572,N_14582);
or U14763 (N_14763,N_14623,N_14701);
or U14764 (N_14764,N_14619,N_14664);
or U14765 (N_14765,N_14563,N_14708);
xnor U14766 (N_14766,N_14599,N_14681);
or U14767 (N_14767,N_14604,N_14698);
or U14768 (N_14768,N_14584,N_14641);
nand U14769 (N_14769,N_14675,N_14665);
or U14770 (N_14770,N_14575,N_14655);
nor U14771 (N_14771,N_14696,N_14702);
or U14772 (N_14772,N_14561,N_14588);
or U14773 (N_14773,N_14689,N_14659);
xnor U14774 (N_14774,N_14638,N_14598);
nand U14775 (N_14775,N_14569,N_14568);
nand U14776 (N_14776,N_14658,N_14680);
xor U14777 (N_14777,N_14640,N_14711);
nor U14778 (N_14778,N_14644,N_14718);
nand U14779 (N_14779,N_14625,N_14614);
or U14780 (N_14780,N_14578,N_14678);
nor U14781 (N_14781,N_14673,N_14683);
nor U14782 (N_14782,N_14684,N_14691);
nand U14783 (N_14783,N_14596,N_14594);
nor U14784 (N_14784,N_14565,N_14583);
or U14785 (N_14785,N_14694,N_14601);
and U14786 (N_14786,N_14651,N_14636);
or U14787 (N_14787,N_14585,N_14647);
nand U14788 (N_14788,N_14719,N_14685);
nand U14789 (N_14789,N_14620,N_14688);
xor U14790 (N_14790,N_14621,N_14642);
or U14791 (N_14791,N_14682,N_14605);
and U14792 (N_14792,N_14577,N_14690);
or U14793 (N_14793,N_14603,N_14710);
xor U14794 (N_14794,N_14716,N_14670);
nor U14795 (N_14795,N_14562,N_14595);
nand U14796 (N_14796,N_14656,N_14629);
nand U14797 (N_14797,N_14666,N_14707);
xor U14798 (N_14798,N_14709,N_14612);
xor U14799 (N_14799,N_14713,N_14617);
and U14800 (N_14800,N_14595,N_14607);
and U14801 (N_14801,N_14589,N_14703);
nand U14802 (N_14802,N_14651,N_14649);
and U14803 (N_14803,N_14705,N_14703);
and U14804 (N_14804,N_14617,N_14676);
or U14805 (N_14805,N_14607,N_14651);
and U14806 (N_14806,N_14634,N_14569);
and U14807 (N_14807,N_14697,N_14703);
nor U14808 (N_14808,N_14575,N_14614);
or U14809 (N_14809,N_14601,N_14660);
nand U14810 (N_14810,N_14646,N_14619);
nand U14811 (N_14811,N_14572,N_14658);
or U14812 (N_14812,N_14668,N_14697);
and U14813 (N_14813,N_14588,N_14610);
or U14814 (N_14814,N_14606,N_14635);
nand U14815 (N_14815,N_14717,N_14674);
nand U14816 (N_14816,N_14604,N_14708);
and U14817 (N_14817,N_14651,N_14719);
and U14818 (N_14818,N_14654,N_14704);
nand U14819 (N_14819,N_14654,N_14665);
and U14820 (N_14820,N_14692,N_14668);
xnor U14821 (N_14821,N_14707,N_14621);
or U14822 (N_14822,N_14620,N_14561);
xor U14823 (N_14823,N_14676,N_14622);
nor U14824 (N_14824,N_14670,N_14700);
and U14825 (N_14825,N_14621,N_14560);
and U14826 (N_14826,N_14632,N_14688);
and U14827 (N_14827,N_14629,N_14676);
nor U14828 (N_14828,N_14562,N_14704);
xnor U14829 (N_14829,N_14610,N_14576);
nand U14830 (N_14830,N_14603,N_14580);
nand U14831 (N_14831,N_14706,N_14637);
xor U14832 (N_14832,N_14689,N_14653);
or U14833 (N_14833,N_14576,N_14650);
xnor U14834 (N_14834,N_14622,N_14660);
and U14835 (N_14835,N_14636,N_14667);
xor U14836 (N_14836,N_14656,N_14673);
nor U14837 (N_14837,N_14662,N_14571);
xnor U14838 (N_14838,N_14606,N_14702);
or U14839 (N_14839,N_14680,N_14690);
nand U14840 (N_14840,N_14712,N_14715);
or U14841 (N_14841,N_14595,N_14661);
nand U14842 (N_14842,N_14689,N_14703);
and U14843 (N_14843,N_14640,N_14713);
and U14844 (N_14844,N_14719,N_14636);
or U14845 (N_14845,N_14672,N_14651);
nand U14846 (N_14846,N_14635,N_14672);
or U14847 (N_14847,N_14634,N_14639);
and U14848 (N_14848,N_14648,N_14603);
nand U14849 (N_14849,N_14660,N_14689);
nand U14850 (N_14850,N_14662,N_14618);
nand U14851 (N_14851,N_14707,N_14697);
and U14852 (N_14852,N_14597,N_14574);
nor U14853 (N_14853,N_14643,N_14637);
nand U14854 (N_14854,N_14717,N_14590);
or U14855 (N_14855,N_14563,N_14582);
and U14856 (N_14856,N_14620,N_14649);
nor U14857 (N_14857,N_14595,N_14574);
nor U14858 (N_14858,N_14692,N_14681);
nor U14859 (N_14859,N_14660,N_14712);
nor U14860 (N_14860,N_14629,N_14607);
xor U14861 (N_14861,N_14686,N_14568);
nand U14862 (N_14862,N_14572,N_14574);
nand U14863 (N_14863,N_14640,N_14670);
or U14864 (N_14864,N_14689,N_14625);
or U14865 (N_14865,N_14581,N_14676);
nor U14866 (N_14866,N_14680,N_14572);
and U14867 (N_14867,N_14586,N_14665);
nor U14868 (N_14868,N_14662,N_14595);
and U14869 (N_14869,N_14631,N_14674);
xor U14870 (N_14870,N_14661,N_14685);
or U14871 (N_14871,N_14583,N_14702);
nor U14872 (N_14872,N_14663,N_14708);
and U14873 (N_14873,N_14588,N_14699);
or U14874 (N_14874,N_14591,N_14636);
or U14875 (N_14875,N_14591,N_14641);
nor U14876 (N_14876,N_14619,N_14616);
nand U14877 (N_14877,N_14596,N_14569);
nand U14878 (N_14878,N_14694,N_14620);
and U14879 (N_14879,N_14650,N_14599);
or U14880 (N_14880,N_14807,N_14782);
xnor U14881 (N_14881,N_14811,N_14861);
xor U14882 (N_14882,N_14790,N_14796);
xor U14883 (N_14883,N_14860,N_14750);
and U14884 (N_14884,N_14776,N_14873);
nand U14885 (N_14885,N_14842,N_14856);
nor U14886 (N_14886,N_14818,N_14826);
and U14887 (N_14887,N_14788,N_14876);
or U14888 (N_14888,N_14748,N_14760);
nor U14889 (N_14889,N_14813,N_14768);
and U14890 (N_14890,N_14743,N_14835);
xor U14891 (N_14891,N_14799,N_14852);
nor U14892 (N_14892,N_14735,N_14867);
xnor U14893 (N_14893,N_14774,N_14849);
and U14894 (N_14894,N_14803,N_14822);
or U14895 (N_14895,N_14756,N_14823);
nand U14896 (N_14896,N_14850,N_14720);
nor U14897 (N_14897,N_14833,N_14859);
nand U14898 (N_14898,N_14779,N_14812);
or U14899 (N_14899,N_14846,N_14877);
nand U14900 (N_14900,N_14764,N_14769);
and U14901 (N_14901,N_14864,N_14798);
or U14902 (N_14902,N_14809,N_14829);
nand U14903 (N_14903,N_14847,N_14840);
and U14904 (N_14904,N_14858,N_14737);
nand U14905 (N_14905,N_14772,N_14815);
xor U14906 (N_14906,N_14729,N_14739);
and U14907 (N_14907,N_14757,N_14728);
or U14908 (N_14908,N_14787,N_14797);
and U14909 (N_14909,N_14879,N_14872);
or U14910 (N_14910,N_14843,N_14830);
or U14911 (N_14911,N_14730,N_14834);
xnor U14912 (N_14912,N_14758,N_14724);
nor U14913 (N_14913,N_14791,N_14853);
or U14914 (N_14914,N_14854,N_14839);
or U14915 (N_14915,N_14736,N_14817);
xor U14916 (N_14916,N_14751,N_14862);
or U14917 (N_14917,N_14740,N_14857);
nor U14918 (N_14918,N_14848,N_14802);
and U14919 (N_14919,N_14754,N_14868);
and U14920 (N_14920,N_14816,N_14837);
nor U14921 (N_14921,N_14875,N_14783);
xor U14922 (N_14922,N_14746,N_14821);
nand U14923 (N_14923,N_14795,N_14742);
or U14924 (N_14924,N_14814,N_14755);
or U14925 (N_14925,N_14874,N_14771);
nor U14926 (N_14926,N_14784,N_14808);
or U14927 (N_14927,N_14789,N_14785);
xor U14928 (N_14928,N_14801,N_14869);
nor U14929 (N_14929,N_14726,N_14722);
nor U14930 (N_14930,N_14844,N_14819);
or U14931 (N_14931,N_14734,N_14747);
nor U14932 (N_14932,N_14800,N_14805);
and U14933 (N_14933,N_14832,N_14744);
nor U14934 (N_14934,N_14723,N_14767);
and U14935 (N_14935,N_14761,N_14721);
xor U14936 (N_14936,N_14851,N_14773);
xnor U14937 (N_14937,N_14727,N_14745);
nand U14938 (N_14938,N_14824,N_14731);
nor U14939 (N_14939,N_14752,N_14863);
nand U14940 (N_14940,N_14841,N_14738);
nand U14941 (N_14941,N_14878,N_14810);
and U14942 (N_14942,N_14793,N_14780);
and U14943 (N_14943,N_14804,N_14820);
nand U14944 (N_14944,N_14845,N_14870);
or U14945 (N_14945,N_14749,N_14759);
and U14946 (N_14946,N_14792,N_14732);
nor U14947 (N_14947,N_14733,N_14765);
xor U14948 (N_14948,N_14786,N_14775);
nor U14949 (N_14949,N_14763,N_14855);
nor U14950 (N_14950,N_14766,N_14770);
nand U14951 (N_14951,N_14827,N_14866);
and U14952 (N_14952,N_14794,N_14753);
nor U14953 (N_14953,N_14741,N_14828);
nor U14954 (N_14954,N_14725,N_14838);
xor U14955 (N_14955,N_14806,N_14781);
or U14956 (N_14956,N_14825,N_14778);
and U14957 (N_14957,N_14865,N_14831);
xor U14958 (N_14958,N_14836,N_14777);
nor U14959 (N_14959,N_14871,N_14762);
or U14960 (N_14960,N_14818,N_14730);
and U14961 (N_14961,N_14829,N_14754);
nor U14962 (N_14962,N_14734,N_14825);
nand U14963 (N_14963,N_14843,N_14747);
or U14964 (N_14964,N_14829,N_14875);
or U14965 (N_14965,N_14733,N_14843);
or U14966 (N_14966,N_14798,N_14854);
nor U14967 (N_14967,N_14847,N_14796);
nand U14968 (N_14968,N_14856,N_14754);
or U14969 (N_14969,N_14855,N_14769);
nand U14970 (N_14970,N_14773,N_14753);
nor U14971 (N_14971,N_14754,N_14801);
xor U14972 (N_14972,N_14836,N_14790);
and U14973 (N_14973,N_14794,N_14856);
xnor U14974 (N_14974,N_14807,N_14803);
xor U14975 (N_14975,N_14776,N_14842);
and U14976 (N_14976,N_14822,N_14791);
nor U14977 (N_14977,N_14842,N_14845);
nor U14978 (N_14978,N_14726,N_14867);
or U14979 (N_14979,N_14853,N_14797);
or U14980 (N_14980,N_14773,N_14776);
or U14981 (N_14981,N_14735,N_14865);
xnor U14982 (N_14982,N_14749,N_14863);
and U14983 (N_14983,N_14727,N_14823);
nor U14984 (N_14984,N_14796,N_14791);
and U14985 (N_14985,N_14860,N_14879);
xor U14986 (N_14986,N_14774,N_14828);
nand U14987 (N_14987,N_14828,N_14813);
and U14988 (N_14988,N_14866,N_14758);
xnor U14989 (N_14989,N_14720,N_14804);
xnor U14990 (N_14990,N_14743,N_14734);
nor U14991 (N_14991,N_14878,N_14725);
xnor U14992 (N_14992,N_14758,N_14873);
or U14993 (N_14993,N_14837,N_14760);
or U14994 (N_14994,N_14784,N_14805);
or U14995 (N_14995,N_14787,N_14872);
and U14996 (N_14996,N_14751,N_14764);
xor U14997 (N_14997,N_14847,N_14751);
nor U14998 (N_14998,N_14843,N_14812);
or U14999 (N_14999,N_14786,N_14751);
xnor U15000 (N_15000,N_14785,N_14803);
nor U15001 (N_15001,N_14833,N_14824);
nand U15002 (N_15002,N_14818,N_14878);
nand U15003 (N_15003,N_14736,N_14827);
or U15004 (N_15004,N_14759,N_14848);
and U15005 (N_15005,N_14749,N_14792);
xnor U15006 (N_15006,N_14779,N_14815);
and U15007 (N_15007,N_14868,N_14829);
or U15008 (N_15008,N_14823,N_14789);
and U15009 (N_15009,N_14787,N_14824);
xor U15010 (N_15010,N_14728,N_14789);
nand U15011 (N_15011,N_14779,N_14870);
xnor U15012 (N_15012,N_14754,N_14724);
and U15013 (N_15013,N_14748,N_14863);
xnor U15014 (N_15014,N_14817,N_14801);
and U15015 (N_15015,N_14876,N_14813);
nor U15016 (N_15016,N_14817,N_14803);
nand U15017 (N_15017,N_14836,N_14815);
and U15018 (N_15018,N_14792,N_14877);
nand U15019 (N_15019,N_14852,N_14798);
nand U15020 (N_15020,N_14756,N_14726);
nor U15021 (N_15021,N_14747,N_14848);
xor U15022 (N_15022,N_14721,N_14792);
nand U15023 (N_15023,N_14861,N_14738);
xnor U15024 (N_15024,N_14875,N_14748);
and U15025 (N_15025,N_14832,N_14877);
xor U15026 (N_15026,N_14854,N_14849);
nor U15027 (N_15027,N_14827,N_14792);
xnor U15028 (N_15028,N_14776,N_14791);
nand U15029 (N_15029,N_14878,N_14797);
or U15030 (N_15030,N_14852,N_14807);
nand U15031 (N_15031,N_14750,N_14807);
nand U15032 (N_15032,N_14851,N_14815);
and U15033 (N_15033,N_14822,N_14828);
nand U15034 (N_15034,N_14777,N_14748);
nand U15035 (N_15035,N_14771,N_14802);
or U15036 (N_15036,N_14790,N_14831);
xor U15037 (N_15037,N_14758,N_14786);
nor U15038 (N_15038,N_14844,N_14799);
and U15039 (N_15039,N_14789,N_14878);
or U15040 (N_15040,N_14990,N_14971);
nor U15041 (N_15041,N_14967,N_14982);
or U15042 (N_15042,N_14927,N_14898);
or U15043 (N_15043,N_14998,N_14880);
nand U15044 (N_15044,N_14956,N_14906);
xnor U15045 (N_15045,N_14981,N_14993);
nand U15046 (N_15046,N_14976,N_14946);
or U15047 (N_15047,N_14974,N_14948);
and U15048 (N_15048,N_14962,N_14922);
nand U15049 (N_15049,N_14970,N_14923);
and U15050 (N_15050,N_14949,N_14975);
and U15051 (N_15051,N_15023,N_14938);
nand U15052 (N_15052,N_14904,N_14964);
and U15053 (N_15053,N_15029,N_14947);
or U15054 (N_15054,N_15027,N_14983);
and U15055 (N_15055,N_15036,N_14914);
nor U15056 (N_15056,N_14959,N_15030);
nand U15057 (N_15057,N_14917,N_14991);
nand U15058 (N_15058,N_14908,N_15038);
xnor U15059 (N_15059,N_14932,N_14887);
xor U15060 (N_15060,N_15019,N_15008);
and U15061 (N_15061,N_14900,N_14913);
nor U15062 (N_15062,N_14940,N_14954);
or U15063 (N_15063,N_14955,N_15032);
xor U15064 (N_15064,N_14907,N_14915);
nand U15065 (N_15065,N_15031,N_14989);
nor U15066 (N_15066,N_14951,N_15022);
xor U15067 (N_15067,N_15018,N_14937);
nor U15068 (N_15068,N_15005,N_15021);
nand U15069 (N_15069,N_14918,N_14901);
xor U15070 (N_15070,N_14952,N_14945);
nand U15071 (N_15071,N_14886,N_14939);
nand U15072 (N_15072,N_15035,N_14889);
xor U15073 (N_15073,N_14979,N_15001);
xor U15074 (N_15074,N_14925,N_14920);
nor U15075 (N_15075,N_14926,N_15000);
nor U15076 (N_15076,N_14896,N_15034);
nand U15077 (N_15077,N_15013,N_15015);
and U15078 (N_15078,N_15039,N_14958);
and U15079 (N_15079,N_14953,N_14966);
and U15080 (N_15080,N_14881,N_14895);
nand U15081 (N_15081,N_14894,N_14933);
and U15082 (N_15082,N_14930,N_14995);
nor U15083 (N_15083,N_14890,N_14882);
nand U15084 (N_15084,N_14935,N_14987);
or U15085 (N_15085,N_14921,N_14919);
and U15086 (N_15086,N_14944,N_14903);
or U15087 (N_15087,N_14988,N_14984);
nand U15088 (N_15088,N_14884,N_14897);
and U15089 (N_15089,N_14941,N_14973);
or U15090 (N_15090,N_14961,N_15020);
nand U15091 (N_15091,N_14978,N_14986);
nand U15092 (N_15092,N_15002,N_14950);
xor U15093 (N_15093,N_14916,N_14996);
and U15094 (N_15094,N_15006,N_15025);
xor U15095 (N_15095,N_14994,N_14997);
or U15096 (N_15096,N_15014,N_14892);
nor U15097 (N_15097,N_15007,N_14969);
xor U15098 (N_15098,N_15028,N_14972);
nor U15099 (N_15099,N_14893,N_15026);
and U15100 (N_15100,N_15012,N_14929);
nor U15101 (N_15101,N_14911,N_14965);
nand U15102 (N_15102,N_14899,N_15011);
nor U15103 (N_15103,N_14977,N_14888);
nand U15104 (N_15104,N_15017,N_14980);
nor U15105 (N_15105,N_14963,N_15016);
or U15106 (N_15106,N_14909,N_14883);
or U15107 (N_15107,N_14936,N_14910);
and U15108 (N_15108,N_14912,N_14931);
and U15109 (N_15109,N_14924,N_14992);
nand U15110 (N_15110,N_14968,N_14960);
or U15111 (N_15111,N_14928,N_14957);
and U15112 (N_15112,N_15004,N_14985);
and U15113 (N_15113,N_14905,N_15010);
nor U15114 (N_15114,N_14943,N_14885);
and U15115 (N_15115,N_15033,N_14891);
nor U15116 (N_15116,N_15037,N_15003);
nor U15117 (N_15117,N_14934,N_14902);
nand U15118 (N_15118,N_14942,N_15024);
nand U15119 (N_15119,N_14999,N_15009);
xnor U15120 (N_15120,N_14913,N_14932);
and U15121 (N_15121,N_14979,N_15039);
nor U15122 (N_15122,N_15033,N_14941);
xor U15123 (N_15123,N_14934,N_14898);
nand U15124 (N_15124,N_14939,N_14936);
or U15125 (N_15125,N_14919,N_14997);
nor U15126 (N_15126,N_14929,N_14992);
and U15127 (N_15127,N_14914,N_15030);
nor U15128 (N_15128,N_14960,N_14974);
nor U15129 (N_15129,N_15036,N_14985);
xor U15130 (N_15130,N_15037,N_14882);
xnor U15131 (N_15131,N_14968,N_15000);
and U15132 (N_15132,N_14888,N_14971);
and U15133 (N_15133,N_15011,N_14995);
nand U15134 (N_15134,N_14927,N_14982);
xnor U15135 (N_15135,N_14996,N_14999);
and U15136 (N_15136,N_14994,N_14926);
and U15137 (N_15137,N_14882,N_14964);
nand U15138 (N_15138,N_14996,N_14908);
and U15139 (N_15139,N_14895,N_14901);
xnor U15140 (N_15140,N_14973,N_14943);
xnor U15141 (N_15141,N_14951,N_14929);
and U15142 (N_15142,N_15025,N_14981);
nand U15143 (N_15143,N_14924,N_14942);
and U15144 (N_15144,N_15029,N_14920);
nor U15145 (N_15145,N_14907,N_14888);
or U15146 (N_15146,N_14910,N_14933);
nor U15147 (N_15147,N_14948,N_15002);
nor U15148 (N_15148,N_14964,N_15022);
nand U15149 (N_15149,N_15035,N_15006);
xnor U15150 (N_15150,N_14956,N_14964);
xor U15151 (N_15151,N_14901,N_14961);
and U15152 (N_15152,N_14915,N_15039);
or U15153 (N_15153,N_15021,N_14932);
nand U15154 (N_15154,N_14986,N_15035);
xnor U15155 (N_15155,N_14945,N_14880);
nor U15156 (N_15156,N_14996,N_14983);
or U15157 (N_15157,N_14886,N_15011);
or U15158 (N_15158,N_15013,N_14989);
or U15159 (N_15159,N_14999,N_15007);
nor U15160 (N_15160,N_14947,N_14942);
nor U15161 (N_15161,N_14955,N_14999);
xor U15162 (N_15162,N_14965,N_14880);
nand U15163 (N_15163,N_15038,N_14985);
and U15164 (N_15164,N_14919,N_14947);
xnor U15165 (N_15165,N_14931,N_14925);
nand U15166 (N_15166,N_14882,N_14983);
nand U15167 (N_15167,N_14992,N_14979);
xor U15168 (N_15168,N_14949,N_14966);
xnor U15169 (N_15169,N_14911,N_15008);
or U15170 (N_15170,N_14926,N_14973);
nand U15171 (N_15171,N_15003,N_14981);
xor U15172 (N_15172,N_14969,N_14998);
xnor U15173 (N_15173,N_14933,N_14966);
or U15174 (N_15174,N_14883,N_14946);
nand U15175 (N_15175,N_14984,N_14990);
nand U15176 (N_15176,N_14885,N_14896);
or U15177 (N_15177,N_15024,N_14983);
and U15178 (N_15178,N_14920,N_14984);
or U15179 (N_15179,N_14930,N_14994);
and U15180 (N_15180,N_15004,N_14944);
nand U15181 (N_15181,N_15021,N_14896);
nand U15182 (N_15182,N_15013,N_14945);
nor U15183 (N_15183,N_14940,N_14944);
and U15184 (N_15184,N_15012,N_14969);
nor U15185 (N_15185,N_14899,N_15020);
xor U15186 (N_15186,N_14992,N_15026);
or U15187 (N_15187,N_14952,N_14943);
xor U15188 (N_15188,N_14914,N_15005);
xnor U15189 (N_15189,N_15033,N_14895);
nand U15190 (N_15190,N_14953,N_14898);
and U15191 (N_15191,N_14978,N_14939);
xnor U15192 (N_15192,N_14884,N_14970);
nand U15193 (N_15193,N_14895,N_14915);
nor U15194 (N_15194,N_14925,N_14894);
nor U15195 (N_15195,N_14999,N_14970);
xor U15196 (N_15196,N_15036,N_14973);
or U15197 (N_15197,N_14986,N_14991);
or U15198 (N_15198,N_14940,N_14992);
nor U15199 (N_15199,N_15028,N_15010);
and U15200 (N_15200,N_15059,N_15156);
xor U15201 (N_15201,N_15187,N_15066);
xnor U15202 (N_15202,N_15115,N_15199);
nor U15203 (N_15203,N_15182,N_15108);
and U15204 (N_15204,N_15192,N_15152);
xor U15205 (N_15205,N_15137,N_15077);
and U15206 (N_15206,N_15147,N_15061);
nand U15207 (N_15207,N_15073,N_15136);
nor U15208 (N_15208,N_15106,N_15103);
nor U15209 (N_15209,N_15111,N_15185);
or U15210 (N_15210,N_15054,N_15101);
and U15211 (N_15211,N_15072,N_15180);
nand U15212 (N_15212,N_15160,N_15090);
or U15213 (N_15213,N_15172,N_15138);
nor U15214 (N_15214,N_15048,N_15041);
or U15215 (N_15215,N_15087,N_15083);
nand U15216 (N_15216,N_15196,N_15092);
xnor U15217 (N_15217,N_15150,N_15052);
or U15218 (N_15218,N_15181,N_15190);
and U15219 (N_15219,N_15088,N_15155);
nand U15220 (N_15220,N_15120,N_15085);
and U15221 (N_15221,N_15091,N_15056);
nor U15222 (N_15222,N_15107,N_15164);
nand U15223 (N_15223,N_15166,N_15131);
nand U15224 (N_15224,N_15157,N_15114);
xnor U15225 (N_15225,N_15173,N_15098);
nor U15226 (N_15226,N_15141,N_15125);
nand U15227 (N_15227,N_15133,N_15153);
xnor U15228 (N_15228,N_15070,N_15096);
xnor U15229 (N_15229,N_15169,N_15165);
xnor U15230 (N_15230,N_15129,N_15176);
xor U15231 (N_15231,N_15068,N_15163);
nor U15232 (N_15232,N_15174,N_15195);
xor U15233 (N_15233,N_15134,N_15105);
xnor U15234 (N_15234,N_15127,N_15122);
and U15235 (N_15235,N_15112,N_15058);
and U15236 (N_15236,N_15167,N_15093);
xor U15237 (N_15237,N_15045,N_15135);
and U15238 (N_15238,N_15154,N_15080);
nor U15239 (N_15239,N_15062,N_15064);
xnor U15240 (N_15240,N_15158,N_15099);
nor U15241 (N_15241,N_15116,N_15118);
nor U15242 (N_15242,N_15132,N_15145);
xnor U15243 (N_15243,N_15184,N_15097);
nand U15244 (N_15244,N_15124,N_15113);
or U15245 (N_15245,N_15143,N_15142);
nand U15246 (N_15246,N_15086,N_15089);
and U15247 (N_15247,N_15100,N_15119);
xnor U15248 (N_15248,N_15071,N_15102);
nor U15249 (N_15249,N_15130,N_15046);
or U15250 (N_15250,N_15050,N_15067);
nor U15251 (N_15251,N_15191,N_15128);
nand U15252 (N_15252,N_15123,N_15186);
nand U15253 (N_15253,N_15140,N_15162);
and U15254 (N_15254,N_15040,N_15110);
nor U15255 (N_15255,N_15055,N_15074);
xor U15256 (N_15256,N_15104,N_15159);
or U15257 (N_15257,N_15177,N_15063);
or U15258 (N_15258,N_15069,N_15047);
xnor U15259 (N_15259,N_15149,N_15075);
and U15260 (N_15260,N_15117,N_15084);
xor U15261 (N_15261,N_15065,N_15178);
or U15262 (N_15262,N_15161,N_15194);
xor U15263 (N_15263,N_15189,N_15126);
or U15264 (N_15264,N_15170,N_15193);
and U15265 (N_15265,N_15148,N_15144);
xnor U15266 (N_15266,N_15049,N_15151);
and U15267 (N_15267,N_15042,N_15044);
or U15268 (N_15268,N_15043,N_15121);
or U15269 (N_15269,N_15095,N_15082);
xor U15270 (N_15270,N_15168,N_15076);
and U15271 (N_15271,N_15109,N_15183);
or U15272 (N_15272,N_15198,N_15057);
nor U15273 (N_15273,N_15079,N_15179);
and U15274 (N_15274,N_15139,N_15094);
xor U15275 (N_15275,N_15081,N_15171);
or U15276 (N_15276,N_15051,N_15197);
nand U15277 (N_15277,N_15060,N_15175);
xnor U15278 (N_15278,N_15188,N_15078);
nand U15279 (N_15279,N_15053,N_15146);
nand U15280 (N_15280,N_15147,N_15118);
or U15281 (N_15281,N_15117,N_15093);
xnor U15282 (N_15282,N_15074,N_15136);
xnor U15283 (N_15283,N_15044,N_15113);
nor U15284 (N_15284,N_15094,N_15194);
and U15285 (N_15285,N_15095,N_15050);
xnor U15286 (N_15286,N_15163,N_15041);
xnor U15287 (N_15287,N_15165,N_15152);
and U15288 (N_15288,N_15192,N_15172);
and U15289 (N_15289,N_15086,N_15151);
nor U15290 (N_15290,N_15088,N_15178);
nor U15291 (N_15291,N_15147,N_15172);
or U15292 (N_15292,N_15094,N_15151);
and U15293 (N_15293,N_15114,N_15145);
nand U15294 (N_15294,N_15198,N_15134);
nor U15295 (N_15295,N_15143,N_15050);
nand U15296 (N_15296,N_15175,N_15093);
xor U15297 (N_15297,N_15119,N_15112);
xnor U15298 (N_15298,N_15134,N_15179);
and U15299 (N_15299,N_15115,N_15130);
or U15300 (N_15300,N_15173,N_15077);
nor U15301 (N_15301,N_15148,N_15154);
or U15302 (N_15302,N_15118,N_15098);
nand U15303 (N_15303,N_15052,N_15175);
nand U15304 (N_15304,N_15055,N_15138);
and U15305 (N_15305,N_15059,N_15088);
or U15306 (N_15306,N_15040,N_15091);
xor U15307 (N_15307,N_15197,N_15041);
nor U15308 (N_15308,N_15107,N_15140);
or U15309 (N_15309,N_15147,N_15075);
and U15310 (N_15310,N_15138,N_15071);
nor U15311 (N_15311,N_15119,N_15188);
xor U15312 (N_15312,N_15140,N_15156);
nand U15313 (N_15313,N_15132,N_15198);
nand U15314 (N_15314,N_15118,N_15048);
or U15315 (N_15315,N_15079,N_15130);
xor U15316 (N_15316,N_15125,N_15177);
xnor U15317 (N_15317,N_15049,N_15162);
nand U15318 (N_15318,N_15073,N_15174);
or U15319 (N_15319,N_15166,N_15139);
and U15320 (N_15320,N_15137,N_15082);
or U15321 (N_15321,N_15073,N_15194);
xnor U15322 (N_15322,N_15121,N_15042);
nor U15323 (N_15323,N_15175,N_15071);
nor U15324 (N_15324,N_15170,N_15054);
or U15325 (N_15325,N_15076,N_15146);
nor U15326 (N_15326,N_15188,N_15176);
xor U15327 (N_15327,N_15156,N_15183);
xor U15328 (N_15328,N_15116,N_15105);
and U15329 (N_15329,N_15140,N_15153);
and U15330 (N_15330,N_15111,N_15170);
nor U15331 (N_15331,N_15103,N_15145);
nand U15332 (N_15332,N_15082,N_15141);
xnor U15333 (N_15333,N_15097,N_15108);
or U15334 (N_15334,N_15189,N_15188);
nand U15335 (N_15335,N_15191,N_15141);
or U15336 (N_15336,N_15198,N_15188);
nor U15337 (N_15337,N_15127,N_15145);
xnor U15338 (N_15338,N_15192,N_15050);
nand U15339 (N_15339,N_15139,N_15045);
xnor U15340 (N_15340,N_15085,N_15108);
or U15341 (N_15341,N_15158,N_15179);
nand U15342 (N_15342,N_15190,N_15176);
and U15343 (N_15343,N_15068,N_15169);
xnor U15344 (N_15344,N_15051,N_15131);
nand U15345 (N_15345,N_15063,N_15199);
xor U15346 (N_15346,N_15091,N_15184);
or U15347 (N_15347,N_15136,N_15157);
nand U15348 (N_15348,N_15111,N_15053);
nand U15349 (N_15349,N_15133,N_15120);
nand U15350 (N_15350,N_15144,N_15117);
xnor U15351 (N_15351,N_15065,N_15072);
nor U15352 (N_15352,N_15185,N_15183);
nand U15353 (N_15353,N_15130,N_15091);
or U15354 (N_15354,N_15136,N_15199);
xor U15355 (N_15355,N_15120,N_15043);
and U15356 (N_15356,N_15074,N_15064);
nor U15357 (N_15357,N_15068,N_15054);
nand U15358 (N_15358,N_15175,N_15187);
nand U15359 (N_15359,N_15074,N_15043);
nor U15360 (N_15360,N_15219,N_15256);
nor U15361 (N_15361,N_15354,N_15206);
and U15362 (N_15362,N_15216,N_15287);
nand U15363 (N_15363,N_15238,N_15343);
and U15364 (N_15364,N_15244,N_15297);
nand U15365 (N_15365,N_15284,N_15241);
nand U15366 (N_15366,N_15351,N_15347);
xor U15367 (N_15367,N_15357,N_15242);
nand U15368 (N_15368,N_15295,N_15235);
and U15369 (N_15369,N_15263,N_15274);
nor U15370 (N_15370,N_15303,N_15337);
and U15371 (N_15371,N_15340,N_15232);
nor U15372 (N_15372,N_15278,N_15272);
nand U15373 (N_15373,N_15260,N_15285);
xor U15374 (N_15374,N_15356,N_15246);
nor U15375 (N_15375,N_15248,N_15240);
or U15376 (N_15376,N_15214,N_15298);
and U15377 (N_15377,N_15210,N_15275);
or U15378 (N_15378,N_15330,N_15209);
or U15379 (N_15379,N_15223,N_15341);
or U15380 (N_15380,N_15325,N_15282);
and U15381 (N_15381,N_15332,N_15290);
xnor U15382 (N_15382,N_15220,N_15301);
nand U15383 (N_15383,N_15315,N_15213);
and U15384 (N_15384,N_15236,N_15279);
nor U15385 (N_15385,N_15268,N_15212);
nand U15386 (N_15386,N_15336,N_15321);
nor U15387 (N_15387,N_15229,N_15237);
and U15388 (N_15388,N_15286,N_15227);
xnor U15389 (N_15389,N_15313,N_15322);
or U15390 (N_15390,N_15342,N_15353);
nor U15391 (N_15391,N_15231,N_15273);
nor U15392 (N_15392,N_15333,N_15252);
xor U15393 (N_15393,N_15239,N_15344);
or U15394 (N_15394,N_15225,N_15348);
nor U15395 (N_15395,N_15207,N_15312);
xor U15396 (N_15396,N_15277,N_15211);
nand U15397 (N_15397,N_15304,N_15265);
or U15398 (N_15398,N_15226,N_15250);
and U15399 (N_15399,N_15318,N_15291);
or U15400 (N_15400,N_15326,N_15281);
and U15401 (N_15401,N_15300,N_15305);
or U15402 (N_15402,N_15289,N_15251);
and U15403 (N_15403,N_15302,N_15316);
and U15404 (N_15404,N_15259,N_15205);
and U15405 (N_15405,N_15253,N_15270);
nor U15406 (N_15406,N_15247,N_15215);
and U15407 (N_15407,N_15255,N_15320);
nor U15408 (N_15408,N_15234,N_15352);
nor U15409 (N_15409,N_15307,N_15355);
nor U15410 (N_15410,N_15293,N_15319);
xnor U15411 (N_15411,N_15292,N_15224);
xor U15412 (N_15412,N_15262,N_15311);
and U15413 (N_15413,N_15296,N_15217);
or U15414 (N_15414,N_15254,N_15308);
and U15415 (N_15415,N_15331,N_15328);
xnor U15416 (N_15416,N_15338,N_15314);
and U15417 (N_15417,N_15266,N_15280);
xnor U15418 (N_15418,N_15245,N_15257);
nor U15419 (N_15419,N_15334,N_15269);
nand U15420 (N_15420,N_15267,N_15339);
xor U15421 (N_15421,N_15218,N_15323);
or U15422 (N_15422,N_15276,N_15261);
nor U15423 (N_15423,N_15324,N_15335);
or U15424 (N_15424,N_15200,N_15222);
or U15425 (N_15425,N_15299,N_15201);
and U15426 (N_15426,N_15358,N_15249);
nor U15427 (N_15427,N_15258,N_15310);
or U15428 (N_15428,N_15359,N_15283);
nand U15429 (N_15429,N_15233,N_15349);
xor U15430 (N_15430,N_15327,N_15294);
xnor U15431 (N_15431,N_15202,N_15317);
nand U15432 (N_15432,N_15264,N_15204);
xnor U15433 (N_15433,N_15306,N_15345);
nand U15434 (N_15434,N_15243,N_15309);
nor U15435 (N_15435,N_15208,N_15329);
nor U15436 (N_15436,N_15350,N_15228);
nand U15437 (N_15437,N_15271,N_15288);
and U15438 (N_15438,N_15230,N_15203);
and U15439 (N_15439,N_15221,N_15346);
or U15440 (N_15440,N_15232,N_15252);
and U15441 (N_15441,N_15215,N_15239);
nand U15442 (N_15442,N_15281,N_15263);
and U15443 (N_15443,N_15323,N_15301);
and U15444 (N_15444,N_15246,N_15328);
nor U15445 (N_15445,N_15283,N_15254);
and U15446 (N_15446,N_15208,N_15316);
and U15447 (N_15447,N_15272,N_15238);
xnor U15448 (N_15448,N_15356,N_15354);
or U15449 (N_15449,N_15304,N_15268);
nor U15450 (N_15450,N_15299,N_15230);
nor U15451 (N_15451,N_15221,N_15246);
nor U15452 (N_15452,N_15356,N_15200);
nor U15453 (N_15453,N_15267,N_15357);
nor U15454 (N_15454,N_15345,N_15292);
and U15455 (N_15455,N_15321,N_15217);
xnor U15456 (N_15456,N_15265,N_15228);
or U15457 (N_15457,N_15222,N_15334);
nor U15458 (N_15458,N_15251,N_15306);
nor U15459 (N_15459,N_15243,N_15308);
nand U15460 (N_15460,N_15274,N_15287);
nand U15461 (N_15461,N_15310,N_15241);
nor U15462 (N_15462,N_15343,N_15353);
xor U15463 (N_15463,N_15340,N_15255);
nand U15464 (N_15464,N_15275,N_15302);
nor U15465 (N_15465,N_15359,N_15202);
or U15466 (N_15466,N_15344,N_15215);
or U15467 (N_15467,N_15340,N_15244);
xor U15468 (N_15468,N_15220,N_15294);
and U15469 (N_15469,N_15261,N_15315);
and U15470 (N_15470,N_15234,N_15239);
xor U15471 (N_15471,N_15215,N_15217);
or U15472 (N_15472,N_15293,N_15359);
nor U15473 (N_15473,N_15359,N_15239);
nand U15474 (N_15474,N_15311,N_15268);
and U15475 (N_15475,N_15307,N_15349);
or U15476 (N_15476,N_15359,N_15235);
xor U15477 (N_15477,N_15271,N_15319);
xnor U15478 (N_15478,N_15343,N_15339);
xor U15479 (N_15479,N_15250,N_15259);
and U15480 (N_15480,N_15241,N_15346);
and U15481 (N_15481,N_15351,N_15273);
xnor U15482 (N_15482,N_15288,N_15319);
nand U15483 (N_15483,N_15327,N_15344);
nor U15484 (N_15484,N_15305,N_15317);
xnor U15485 (N_15485,N_15257,N_15304);
nand U15486 (N_15486,N_15286,N_15270);
nor U15487 (N_15487,N_15292,N_15265);
xnor U15488 (N_15488,N_15202,N_15282);
or U15489 (N_15489,N_15311,N_15345);
or U15490 (N_15490,N_15286,N_15239);
xor U15491 (N_15491,N_15316,N_15230);
or U15492 (N_15492,N_15313,N_15249);
xnor U15493 (N_15493,N_15254,N_15280);
xor U15494 (N_15494,N_15289,N_15336);
xor U15495 (N_15495,N_15358,N_15311);
xnor U15496 (N_15496,N_15292,N_15351);
nand U15497 (N_15497,N_15238,N_15332);
and U15498 (N_15498,N_15328,N_15353);
or U15499 (N_15499,N_15240,N_15202);
and U15500 (N_15500,N_15295,N_15333);
nor U15501 (N_15501,N_15338,N_15286);
or U15502 (N_15502,N_15313,N_15216);
nand U15503 (N_15503,N_15337,N_15237);
nor U15504 (N_15504,N_15288,N_15235);
nand U15505 (N_15505,N_15317,N_15308);
or U15506 (N_15506,N_15298,N_15306);
and U15507 (N_15507,N_15338,N_15336);
or U15508 (N_15508,N_15234,N_15331);
and U15509 (N_15509,N_15323,N_15234);
and U15510 (N_15510,N_15259,N_15262);
nor U15511 (N_15511,N_15307,N_15244);
nand U15512 (N_15512,N_15276,N_15200);
or U15513 (N_15513,N_15267,N_15240);
or U15514 (N_15514,N_15354,N_15200);
or U15515 (N_15515,N_15321,N_15201);
or U15516 (N_15516,N_15268,N_15239);
or U15517 (N_15517,N_15262,N_15318);
nor U15518 (N_15518,N_15213,N_15313);
and U15519 (N_15519,N_15285,N_15255);
nand U15520 (N_15520,N_15444,N_15366);
xor U15521 (N_15521,N_15416,N_15407);
xor U15522 (N_15522,N_15361,N_15427);
nor U15523 (N_15523,N_15396,N_15389);
xor U15524 (N_15524,N_15469,N_15461);
nor U15525 (N_15525,N_15436,N_15435);
xnor U15526 (N_15526,N_15470,N_15446);
nand U15527 (N_15527,N_15467,N_15500);
nor U15528 (N_15528,N_15372,N_15370);
nand U15529 (N_15529,N_15489,N_15397);
nor U15530 (N_15530,N_15507,N_15501);
nand U15531 (N_15531,N_15494,N_15448);
nand U15532 (N_15532,N_15378,N_15517);
nor U15533 (N_15533,N_15515,N_15443);
nor U15534 (N_15534,N_15504,N_15519);
or U15535 (N_15535,N_15455,N_15360);
or U15536 (N_15536,N_15387,N_15428);
or U15537 (N_15537,N_15404,N_15405);
xor U15538 (N_15538,N_15392,N_15450);
nor U15539 (N_15539,N_15502,N_15367);
nor U15540 (N_15540,N_15365,N_15381);
and U15541 (N_15541,N_15497,N_15481);
nor U15542 (N_15542,N_15373,N_15430);
nand U15543 (N_15543,N_15419,N_15493);
nor U15544 (N_15544,N_15482,N_15496);
and U15545 (N_15545,N_15512,N_15447);
and U15546 (N_15546,N_15433,N_15458);
nor U15547 (N_15547,N_15398,N_15487);
or U15548 (N_15548,N_15383,N_15460);
or U15549 (N_15549,N_15457,N_15362);
and U15550 (N_15550,N_15425,N_15379);
or U15551 (N_15551,N_15498,N_15422);
nor U15552 (N_15552,N_15485,N_15483);
or U15553 (N_15553,N_15380,N_15429);
and U15554 (N_15554,N_15363,N_15424);
and U15555 (N_15555,N_15475,N_15477);
and U15556 (N_15556,N_15393,N_15514);
or U15557 (N_15557,N_15403,N_15472);
xnor U15558 (N_15558,N_15452,N_15402);
and U15559 (N_15559,N_15456,N_15463);
xor U15560 (N_15560,N_15412,N_15386);
xnor U15561 (N_15561,N_15505,N_15449);
xor U15562 (N_15562,N_15484,N_15385);
and U15563 (N_15563,N_15516,N_15462);
nor U15564 (N_15564,N_15390,N_15437);
and U15565 (N_15565,N_15479,N_15391);
nor U15566 (N_15566,N_15395,N_15459);
nand U15567 (N_15567,N_15454,N_15371);
nor U15568 (N_15568,N_15453,N_15369);
or U15569 (N_15569,N_15408,N_15431);
xor U15570 (N_15570,N_15406,N_15480);
xnor U15571 (N_15571,N_15426,N_15432);
and U15572 (N_15572,N_15394,N_15518);
xnor U15573 (N_15573,N_15375,N_15478);
xnor U15574 (N_15574,N_15418,N_15486);
or U15575 (N_15575,N_15468,N_15415);
nor U15576 (N_15576,N_15464,N_15491);
xnor U15577 (N_15577,N_15503,N_15401);
or U15578 (N_15578,N_15364,N_15421);
nand U15579 (N_15579,N_15466,N_15417);
and U15580 (N_15580,N_15411,N_15509);
and U15581 (N_15581,N_15451,N_15409);
nor U15582 (N_15582,N_15476,N_15488);
nor U15583 (N_15583,N_15495,N_15384);
and U15584 (N_15584,N_15473,N_15439);
or U15585 (N_15585,N_15511,N_15382);
or U15586 (N_15586,N_15490,N_15414);
nand U15587 (N_15587,N_15376,N_15471);
or U15588 (N_15588,N_15506,N_15400);
xnor U15589 (N_15589,N_15423,N_15508);
nor U15590 (N_15590,N_15465,N_15413);
nand U15591 (N_15591,N_15377,N_15442);
nand U15592 (N_15592,N_15440,N_15510);
or U15593 (N_15593,N_15368,N_15434);
nand U15594 (N_15594,N_15374,N_15388);
or U15595 (N_15595,N_15492,N_15420);
nor U15596 (N_15596,N_15445,N_15399);
and U15597 (N_15597,N_15410,N_15438);
xnor U15598 (N_15598,N_15474,N_15499);
nor U15599 (N_15599,N_15441,N_15513);
and U15600 (N_15600,N_15505,N_15411);
nand U15601 (N_15601,N_15372,N_15403);
nand U15602 (N_15602,N_15392,N_15513);
or U15603 (N_15603,N_15452,N_15420);
nand U15604 (N_15604,N_15484,N_15487);
nand U15605 (N_15605,N_15422,N_15413);
xnor U15606 (N_15606,N_15407,N_15456);
or U15607 (N_15607,N_15391,N_15425);
xnor U15608 (N_15608,N_15365,N_15508);
or U15609 (N_15609,N_15459,N_15502);
and U15610 (N_15610,N_15482,N_15443);
nand U15611 (N_15611,N_15468,N_15435);
nor U15612 (N_15612,N_15369,N_15409);
or U15613 (N_15613,N_15393,N_15510);
and U15614 (N_15614,N_15492,N_15484);
xor U15615 (N_15615,N_15392,N_15362);
xor U15616 (N_15616,N_15459,N_15454);
and U15617 (N_15617,N_15494,N_15427);
or U15618 (N_15618,N_15379,N_15410);
xnor U15619 (N_15619,N_15420,N_15444);
and U15620 (N_15620,N_15481,N_15438);
xnor U15621 (N_15621,N_15460,N_15472);
nand U15622 (N_15622,N_15466,N_15363);
and U15623 (N_15623,N_15378,N_15473);
nand U15624 (N_15624,N_15494,N_15505);
and U15625 (N_15625,N_15438,N_15466);
and U15626 (N_15626,N_15460,N_15444);
nand U15627 (N_15627,N_15419,N_15416);
and U15628 (N_15628,N_15467,N_15437);
nand U15629 (N_15629,N_15391,N_15424);
xnor U15630 (N_15630,N_15497,N_15511);
or U15631 (N_15631,N_15467,N_15464);
or U15632 (N_15632,N_15487,N_15494);
nand U15633 (N_15633,N_15473,N_15454);
nor U15634 (N_15634,N_15500,N_15402);
nor U15635 (N_15635,N_15366,N_15431);
or U15636 (N_15636,N_15482,N_15480);
xor U15637 (N_15637,N_15432,N_15451);
xnor U15638 (N_15638,N_15398,N_15365);
xnor U15639 (N_15639,N_15435,N_15487);
xor U15640 (N_15640,N_15393,N_15498);
nor U15641 (N_15641,N_15506,N_15479);
nand U15642 (N_15642,N_15486,N_15399);
nand U15643 (N_15643,N_15431,N_15506);
or U15644 (N_15644,N_15363,N_15494);
or U15645 (N_15645,N_15496,N_15417);
or U15646 (N_15646,N_15431,N_15387);
nor U15647 (N_15647,N_15492,N_15460);
or U15648 (N_15648,N_15444,N_15428);
and U15649 (N_15649,N_15450,N_15494);
and U15650 (N_15650,N_15436,N_15434);
and U15651 (N_15651,N_15469,N_15416);
nor U15652 (N_15652,N_15378,N_15370);
and U15653 (N_15653,N_15474,N_15363);
or U15654 (N_15654,N_15499,N_15371);
nor U15655 (N_15655,N_15429,N_15457);
or U15656 (N_15656,N_15431,N_15421);
nand U15657 (N_15657,N_15515,N_15511);
nor U15658 (N_15658,N_15503,N_15462);
and U15659 (N_15659,N_15424,N_15482);
nand U15660 (N_15660,N_15402,N_15394);
nand U15661 (N_15661,N_15456,N_15517);
or U15662 (N_15662,N_15495,N_15471);
nand U15663 (N_15663,N_15477,N_15510);
nand U15664 (N_15664,N_15395,N_15410);
nor U15665 (N_15665,N_15391,N_15392);
and U15666 (N_15666,N_15473,N_15444);
nand U15667 (N_15667,N_15421,N_15448);
and U15668 (N_15668,N_15506,N_15436);
or U15669 (N_15669,N_15511,N_15467);
xnor U15670 (N_15670,N_15420,N_15373);
nor U15671 (N_15671,N_15455,N_15456);
and U15672 (N_15672,N_15452,N_15441);
xnor U15673 (N_15673,N_15401,N_15508);
and U15674 (N_15674,N_15417,N_15419);
or U15675 (N_15675,N_15402,N_15369);
nand U15676 (N_15676,N_15442,N_15445);
or U15677 (N_15677,N_15502,N_15501);
nand U15678 (N_15678,N_15402,N_15479);
nor U15679 (N_15679,N_15395,N_15500);
nor U15680 (N_15680,N_15556,N_15539);
nor U15681 (N_15681,N_15533,N_15550);
nand U15682 (N_15682,N_15527,N_15615);
xnor U15683 (N_15683,N_15626,N_15590);
or U15684 (N_15684,N_15653,N_15596);
and U15685 (N_15685,N_15634,N_15618);
xor U15686 (N_15686,N_15629,N_15553);
xor U15687 (N_15687,N_15620,N_15548);
or U15688 (N_15688,N_15655,N_15595);
or U15689 (N_15689,N_15524,N_15574);
nor U15690 (N_15690,N_15534,N_15611);
xor U15691 (N_15691,N_15635,N_15525);
or U15692 (N_15692,N_15673,N_15630);
nor U15693 (N_15693,N_15564,N_15586);
and U15694 (N_15694,N_15554,N_15555);
or U15695 (N_15695,N_15613,N_15542);
nor U15696 (N_15696,N_15632,N_15601);
nand U15697 (N_15697,N_15521,N_15640);
or U15698 (N_15698,N_15605,N_15562);
and U15699 (N_15699,N_15591,N_15663);
xor U15700 (N_15700,N_15641,N_15565);
nor U15701 (N_15701,N_15650,N_15594);
nor U15702 (N_15702,N_15543,N_15606);
or U15703 (N_15703,N_15649,N_15593);
nand U15704 (N_15704,N_15528,N_15633);
nor U15705 (N_15705,N_15625,N_15537);
nor U15706 (N_15706,N_15599,N_15580);
nor U15707 (N_15707,N_15647,N_15670);
xor U15708 (N_15708,N_15610,N_15566);
and U15709 (N_15709,N_15549,N_15668);
nor U15710 (N_15710,N_15529,N_15675);
xnor U15711 (N_15711,N_15679,N_15569);
xnor U15712 (N_15712,N_15652,N_15667);
xor U15713 (N_15713,N_15531,N_15575);
or U15714 (N_15714,N_15623,N_15608);
xor U15715 (N_15715,N_15617,N_15535);
and U15716 (N_15716,N_15614,N_15631);
nand U15717 (N_15717,N_15622,N_15578);
nand U15718 (N_15718,N_15571,N_15627);
nand U15719 (N_15719,N_15636,N_15609);
and U15720 (N_15720,N_15520,N_15592);
xnor U15721 (N_15721,N_15665,N_15644);
xnor U15722 (N_15722,N_15536,N_15600);
nor U15723 (N_15723,N_15545,N_15648);
and U15724 (N_15724,N_15607,N_15616);
xor U15725 (N_15725,N_15603,N_15589);
and U15726 (N_15726,N_15619,N_15587);
nor U15727 (N_15727,N_15597,N_15658);
nor U15728 (N_15728,N_15678,N_15598);
or U15729 (N_15729,N_15560,N_15544);
or U15730 (N_15730,N_15637,N_15643);
nand U15731 (N_15731,N_15656,N_15538);
and U15732 (N_15732,N_15661,N_15642);
nand U15733 (N_15733,N_15561,N_15577);
nor U15734 (N_15734,N_15551,N_15582);
nand U15735 (N_15735,N_15669,N_15666);
or U15736 (N_15736,N_15530,N_15585);
xnor U15737 (N_15737,N_15638,N_15651);
nor U15738 (N_15738,N_15662,N_15664);
nor U15739 (N_15739,N_15654,N_15570);
xnor U15740 (N_15740,N_15602,N_15558);
nor U15741 (N_15741,N_15628,N_15522);
xor U15742 (N_15742,N_15557,N_15552);
or U15743 (N_15743,N_15676,N_15584);
xnor U15744 (N_15744,N_15604,N_15583);
xor U15745 (N_15745,N_15526,N_15588);
xnor U15746 (N_15746,N_15612,N_15657);
nor U15747 (N_15747,N_15677,N_15671);
or U15748 (N_15748,N_15540,N_15568);
and U15749 (N_15749,N_15672,N_15621);
xor U15750 (N_15750,N_15579,N_15541);
nor U15751 (N_15751,N_15547,N_15546);
or U15752 (N_15752,N_15674,N_15532);
nand U15753 (N_15753,N_15559,N_15563);
nand U15754 (N_15754,N_15572,N_15659);
nand U15755 (N_15755,N_15639,N_15573);
or U15756 (N_15756,N_15567,N_15576);
nand U15757 (N_15757,N_15624,N_15645);
or U15758 (N_15758,N_15660,N_15581);
xor U15759 (N_15759,N_15523,N_15646);
or U15760 (N_15760,N_15623,N_15630);
xnor U15761 (N_15761,N_15543,N_15535);
nand U15762 (N_15762,N_15548,N_15532);
nor U15763 (N_15763,N_15551,N_15526);
nand U15764 (N_15764,N_15616,N_15588);
nand U15765 (N_15765,N_15598,N_15667);
and U15766 (N_15766,N_15552,N_15676);
and U15767 (N_15767,N_15664,N_15563);
or U15768 (N_15768,N_15570,N_15572);
or U15769 (N_15769,N_15612,N_15655);
nor U15770 (N_15770,N_15654,N_15554);
and U15771 (N_15771,N_15589,N_15525);
and U15772 (N_15772,N_15639,N_15592);
and U15773 (N_15773,N_15543,N_15671);
nor U15774 (N_15774,N_15614,N_15625);
xnor U15775 (N_15775,N_15609,N_15520);
or U15776 (N_15776,N_15634,N_15553);
xnor U15777 (N_15777,N_15604,N_15527);
or U15778 (N_15778,N_15534,N_15618);
or U15779 (N_15779,N_15609,N_15540);
and U15780 (N_15780,N_15647,N_15605);
nor U15781 (N_15781,N_15557,N_15631);
nand U15782 (N_15782,N_15607,N_15643);
or U15783 (N_15783,N_15677,N_15672);
nor U15784 (N_15784,N_15574,N_15615);
nor U15785 (N_15785,N_15543,N_15633);
nor U15786 (N_15786,N_15606,N_15669);
nor U15787 (N_15787,N_15677,N_15535);
and U15788 (N_15788,N_15661,N_15618);
or U15789 (N_15789,N_15631,N_15598);
and U15790 (N_15790,N_15581,N_15574);
nor U15791 (N_15791,N_15562,N_15653);
or U15792 (N_15792,N_15636,N_15551);
xnor U15793 (N_15793,N_15550,N_15656);
and U15794 (N_15794,N_15631,N_15613);
nor U15795 (N_15795,N_15606,N_15591);
nor U15796 (N_15796,N_15605,N_15585);
and U15797 (N_15797,N_15547,N_15588);
nor U15798 (N_15798,N_15547,N_15661);
nor U15799 (N_15799,N_15638,N_15621);
and U15800 (N_15800,N_15583,N_15614);
xnor U15801 (N_15801,N_15655,N_15635);
nor U15802 (N_15802,N_15555,N_15598);
nand U15803 (N_15803,N_15651,N_15557);
nand U15804 (N_15804,N_15638,N_15627);
nor U15805 (N_15805,N_15643,N_15520);
xor U15806 (N_15806,N_15550,N_15522);
xnor U15807 (N_15807,N_15661,N_15558);
nand U15808 (N_15808,N_15555,N_15634);
xnor U15809 (N_15809,N_15657,N_15645);
xor U15810 (N_15810,N_15527,N_15667);
nor U15811 (N_15811,N_15524,N_15587);
and U15812 (N_15812,N_15532,N_15554);
nand U15813 (N_15813,N_15677,N_15652);
and U15814 (N_15814,N_15618,N_15647);
xnor U15815 (N_15815,N_15637,N_15630);
and U15816 (N_15816,N_15562,N_15665);
xnor U15817 (N_15817,N_15627,N_15549);
or U15818 (N_15818,N_15527,N_15659);
and U15819 (N_15819,N_15565,N_15580);
nand U15820 (N_15820,N_15650,N_15616);
or U15821 (N_15821,N_15530,N_15539);
xnor U15822 (N_15822,N_15662,N_15560);
nand U15823 (N_15823,N_15546,N_15607);
xor U15824 (N_15824,N_15612,N_15644);
xor U15825 (N_15825,N_15589,N_15567);
nand U15826 (N_15826,N_15542,N_15615);
nand U15827 (N_15827,N_15677,N_15610);
xnor U15828 (N_15828,N_15664,N_15538);
and U15829 (N_15829,N_15528,N_15643);
nand U15830 (N_15830,N_15665,N_15574);
or U15831 (N_15831,N_15552,N_15654);
or U15832 (N_15832,N_15676,N_15657);
xor U15833 (N_15833,N_15552,N_15594);
or U15834 (N_15834,N_15609,N_15591);
nor U15835 (N_15835,N_15573,N_15611);
nand U15836 (N_15836,N_15571,N_15585);
nor U15837 (N_15837,N_15547,N_15669);
and U15838 (N_15838,N_15602,N_15634);
or U15839 (N_15839,N_15618,N_15563);
and U15840 (N_15840,N_15687,N_15701);
nand U15841 (N_15841,N_15697,N_15773);
xor U15842 (N_15842,N_15761,N_15835);
nor U15843 (N_15843,N_15784,N_15832);
nor U15844 (N_15844,N_15819,N_15830);
xnor U15845 (N_15845,N_15804,N_15808);
or U15846 (N_15846,N_15689,N_15831);
xnor U15847 (N_15847,N_15749,N_15682);
xnor U15848 (N_15848,N_15820,N_15745);
nand U15849 (N_15849,N_15792,N_15720);
or U15850 (N_15850,N_15709,N_15801);
nand U15851 (N_15851,N_15695,N_15762);
xnor U15852 (N_15852,N_15726,N_15700);
nor U15853 (N_15853,N_15800,N_15732);
or U15854 (N_15854,N_15767,N_15793);
and U15855 (N_15855,N_15777,N_15719);
or U15856 (N_15856,N_15789,N_15833);
or U15857 (N_15857,N_15818,N_15699);
nor U15858 (N_15858,N_15763,N_15780);
or U15859 (N_15859,N_15730,N_15765);
nor U15860 (N_15860,N_15690,N_15828);
xor U15861 (N_15861,N_15812,N_15686);
and U15862 (N_15862,N_15756,N_15729);
nor U15863 (N_15863,N_15711,N_15814);
and U15864 (N_15864,N_15769,N_15751);
nor U15865 (N_15865,N_15742,N_15684);
xnor U15866 (N_15866,N_15740,N_15781);
nor U15867 (N_15867,N_15685,N_15736);
and U15868 (N_15868,N_15707,N_15787);
xor U15869 (N_15869,N_15794,N_15836);
or U15870 (N_15870,N_15779,N_15776);
xor U15871 (N_15871,N_15731,N_15798);
nand U15872 (N_15872,N_15747,N_15680);
nand U15873 (N_15873,N_15683,N_15741);
or U15874 (N_15874,N_15755,N_15753);
or U15875 (N_15875,N_15771,N_15752);
xnor U15876 (N_15876,N_15691,N_15692);
nor U15877 (N_15877,N_15802,N_15723);
or U15878 (N_15878,N_15764,N_15754);
nor U15879 (N_15879,N_15821,N_15760);
and U15880 (N_15880,N_15746,N_15724);
or U15881 (N_15881,N_15681,N_15688);
or U15882 (N_15882,N_15811,N_15713);
and U15883 (N_15883,N_15768,N_15757);
nand U15884 (N_15884,N_15743,N_15813);
or U15885 (N_15885,N_15807,N_15698);
and U15886 (N_15886,N_15710,N_15778);
or U15887 (N_15887,N_15708,N_15829);
xor U15888 (N_15888,N_15825,N_15737);
xnor U15889 (N_15889,N_15714,N_15744);
and U15890 (N_15890,N_15772,N_15809);
nor U15891 (N_15891,N_15693,N_15803);
or U15892 (N_15892,N_15706,N_15838);
and U15893 (N_15893,N_15790,N_15727);
xor U15894 (N_15894,N_15824,N_15759);
nand U15895 (N_15895,N_15816,N_15786);
and U15896 (N_15896,N_15783,N_15728);
nand U15897 (N_15897,N_15834,N_15817);
nand U15898 (N_15898,N_15827,N_15718);
and U15899 (N_15899,N_15810,N_15775);
nand U15900 (N_15900,N_15822,N_15715);
nand U15901 (N_15901,N_15734,N_15748);
and U15902 (N_15902,N_15717,N_15704);
nor U15903 (N_15903,N_15782,N_15797);
nor U15904 (N_15904,N_15702,N_15739);
or U15905 (N_15905,N_15799,N_15815);
nand U15906 (N_15906,N_15694,N_15722);
nand U15907 (N_15907,N_15712,N_15703);
nand U15908 (N_15908,N_15725,N_15721);
or U15909 (N_15909,N_15788,N_15750);
or U15910 (N_15910,N_15774,N_15770);
xnor U15911 (N_15911,N_15826,N_15733);
xor U15912 (N_15912,N_15796,N_15735);
xnor U15913 (N_15913,N_15806,N_15839);
nor U15914 (N_15914,N_15738,N_15795);
or U15915 (N_15915,N_15805,N_15791);
nand U15916 (N_15916,N_15758,N_15705);
nand U15917 (N_15917,N_15696,N_15837);
nor U15918 (N_15918,N_15823,N_15766);
or U15919 (N_15919,N_15716,N_15785);
and U15920 (N_15920,N_15711,N_15829);
or U15921 (N_15921,N_15729,N_15768);
xnor U15922 (N_15922,N_15750,N_15680);
xnor U15923 (N_15923,N_15817,N_15681);
and U15924 (N_15924,N_15835,N_15762);
nor U15925 (N_15925,N_15714,N_15730);
or U15926 (N_15926,N_15827,N_15716);
and U15927 (N_15927,N_15813,N_15837);
nor U15928 (N_15928,N_15712,N_15830);
or U15929 (N_15929,N_15739,N_15828);
or U15930 (N_15930,N_15745,N_15806);
and U15931 (N_15931,N_15822,N_15728);
xnor U15932 (N_15932,N_15693,N_15703);
nor U15933 (N_15933,N_15762,N_15763);
xor U15934 (N_15934,N_15807,N_15809);
nor U15935 (N_15935,N_15801,N_15794);
nor U15936 (N_15936,N_15688,N_15734);
and U15937 (N_15937,N_15686,N_15720);
or U15938 (N_15938,N_15822,N_15772);
nor U15939 (N_15939,N_15721,N_15699);
xor U15940 (N_15940,N_15697,N_15735);
or U15941 (N_15941,N_15700,N_15749);
nand U15942 (N_15942,N_15764,N_15767);
or U15943 (N_15943,N_15811,N_15766);
nand U15944 (N_15944,N_15801,N_15760);
nor U15945 (N_15945,N_15750,N_15773);
nor U15946 (N_15946,N_15807,N_15818);
nor U15947 (N_15947,N_15753,N_15734);
nor U15948 (N_15948,N_15770,N_15790);
nand U15949 (N_15949,N_15774,N_15735);
nand U15950 (N_15950,N_15701,N_15791);
or U15951 (N_15951,N_15829,N_15682);
nand U15952 (N_15952,N_15782,N_15723);
nand U15953 (N_15953,N_15682,N_15823);
and U15954 (N_15954,N_15791,N_15835);
or U15955 (N_15955,N_15825,N_15694);
nor U15956 (N_15956,N_15681,N_15736);
nand U15957 (N_15957,N_15741,N_15833);
or U15958 (N_15958,N_15792,N_15772);
or U15959 (N_15959,N_15684,N_15776);
nand U15960 (N_15960,N_15693,N_15711);
and U15961 (N_15961,N_15803,N_15769);
and U15962 (N_15962,N_15712,N_15738);
nor U15963 (N_15963,N_15834,N_15777);
and U15964 (N_15964,N_15781,N_15701);
nor U15965 (N_15965,N_15805,N_15681);
and U15966 (N_15966,N_15815,N_15757);
or U15967 (N_15967,N_15706,N_15778);
nor U15968 (N_15968,N_15716,N_15808);
or U15969 (N_15969,N_15815,N_15681);
nor U15970 (N_15970,N_15693,N_15763);
xnor U15971 (N_15971,N_15807,N_15788);
and U15972 (N_15972,N_15830,N_15809);
and U15973 (N_15973,N_15756,N_15696);
and U15974 (N_15974,N_15700,N_15685);
nand U15975 (N_15975,N_15828,N_15686);
xnor U15976 (N_15976,N_15716,N_15756);
or U15977 (N_15977,N_15747,N_15695);
nor U15978 (N_15978,N_15765,N_15745);
xnor U15979 (N_15979,N_15683,N_15753);
and U15980 (N_15980,N_15770,N_15807);
nand U15981 (N_15981,N_15811,N_15711);
and U15982 (N_15982,N_15831,N_15744);
nor U15983 (N_15983,N_15775,N_15704);
xnor U15984 (N_15984,N_15786,N_15805);
nor U15985 (N_15985,N_15768,N_15799);
or U15986 (N_15986,N_15759,N_15728);
and U15987 (N_15987,N_15715,N_15716);
xor U15988 (N_15988,N_15707,N_15769);
nor U15989 (N_15989,N_15739,N_15738);
and U15990 (N_15990,N_15817,N_15714);
nor U15991 (N_15991,N_15704,N_15736);
nand U15992 (N_15992,N_15811,N_15788);
nand U15993 (N_15993,N_15688,N_15699);
nor U15994 (N_15994,N_15727,N_15796);
xor U15995 (N_15995,N_15786,N_15775);
xnor U15996 (N_15996,N_15836,N_15822);
xor U15997 (N_15997,N_15800,N_15762);
nor U15998 (N_15998,N_15822,N_15680);
nor U15999 (N_15999,N_15807,N_15780);
xor U16000 (N_16000,N_15904,N_15876);
nor U16001 (N_16001,N_15841,N_15878);
nand U16002 (N_16002,N_15959,N_15996);
nor U16003 (N_16003,N_15874,N_15997);
xnor U16004 (N_16004,N_15954,N_15879);
xor U16005 (N_16005,N_15858,N_15948);
and U16006 (N_16006,N_15920,N_15905);
and U16007 (N_16007,N_15985,N_15974);
xor U16008 (N_16008,N_15892,N_15960);
nand U16009 (N_16009,N_15932,N_15843);
xor U16010 (N_16010,N_15942,N_15909);
nor U16011 (N_16011,N_15919,N_15943);
xnor U16012 (N_16012,N_15978,N_15946);
xnor U16013 (N_16013,N_15992,N_15889);
nor U16014 (N_16014,N_15986,N_15886);
and U16015 (N_16015,N_15977,N_15928);
or U16016 (N_16016,N_15900,N_15924);
nand U16017 (N_16017,N_15880,N_15933);
xnor U16018 (N_16018,N_15949,N_15870);
xor U16019 (N_16019,N_15911,N_15883);
nand U16020 (N_16020,N_15916,N_15845);
or U16021 (N_16021,N_15939,N_15938);
or U16022 (N_16022,N_15875,N_15903);
or U16023 (N_16023,N_15898,N_15935);
and U16024 (N_16024,N_15910,N_15966);
xor U16025 (N_16025,N_15979,N_15990);
xor U16026 (N_16026,N_15976,N_15941);
xnor U16027 (N_16027,N_15973,N_15930);
nor U16028 (N_16028,N_15860,N_15955);
or U16029 (N_16029,N_15970,N_15871);
xnor U16030 (N_16030,N_15850,N_15840);
xnor U16031 (N_16031,N_15934,N_15906);
or U16032 (N_16032,N_15994,N_15912);
xnor U16033 (N_16033,N_15913,N_15988);
nor U16034 (N_16034,N_15859,N_15854);
or U16035 (N_16035,N_15953,N_15961);
and U16036 (N_16036,N_15915,N_15931);
and U16037 (N_16037,N_15914,N_15866);
and U16038 (N_16038,N_15951,N_15929);
nand U16039 (N_16039,N_15962,N_15851);
nor U16040 (N_16040,N_15944,N_15971);
or U16041 (N_16041,N_15852,N_15921);
or U16042 (N_16042,N_15895,N_15980);
and U16043 (N_16043,N_15918,N_15902);
xnor U16044 (N_16044,N_15957,N_15995);
xnor U16045 (N_16045,N_15862,N_15899);
xnor U16046 (N_16046,N_15847,N_15967);
nand U16047 (N_16047,N_15950,N_15917);
nor U16048 (N_16048,N_15887,N_15881);
nor U16049 (N_16049,N_15873,N_15984);
xnor U16050 (N_16050,N_15877,N_15936);
or U16051 (N_16051,N_15882,N_15945);
nor U16052 (N_16052,N_15947,N_15891);
xor U16053 (N_16053,N_15926,N_15975);
nand U16054 (N_16054,N_15925,N_15861);
nor U16055 (N_16055,N_15867,N_15853);
or U16056 (N_16056,N_15956,N_15963);
xor U16057 (N_16057,N_15999,N_15857);
and U16058 (N_16058,N_15968,N_15922);
nor U16059 (N_16059,N_15849,N_15969);
xnor U16060 (N_16060,N_15964,N_15993);
nor U16061 (N_16061,N_15863,N_15842);
nand U16062 (N_16062,N_15894,N_15848);
nand U16063 (N_16063,N_15885,N_15908);
nand U16064 (N_16064,N_15965,N_15983);
and U16065 (N_16065,N_15856,N_15872);
or U16066 (N_16066,N_15991,N_15972);
and U16067 (N_16067,N_15937,N_15844);
nor U16068 (N_16068,N_15846,N_15958);
nand U16069 (N_16069,N_15864,N_15901);
or U16070 (N_16070,N_15888,N_15927);
xor U16071 (N_16071,N_15890,N_15869);
nand U16072 (N_16072,N_15865,N_15982);
or U16073 (N_16073,N_15884,N_15896);
and U16074 (N_16074,N_15998,N_15987);
and U16075 (N_16075,N_15868,N_15893);
nor U16076 (N_16076,N_15989,N_15907);
and U16077 (N_16077,N_15897,N_15855);
or U16078 (N_16078,N_15981,N_15952);
or U16079 (N_16079,N_15923,N_15940);
or U16080 (N_16080,N_15897,N_15935);
nor U16081 (N_16081,N_15841,N_15945);
xor U16082 (N_16082,N_15908,N_15951);
xnor U16083 (N_16083,N_15925,N_15953);
nor U16084 (N_16084,N_15915,N_15930);
xnor U16085 (N_16085,N_15843,N_15988);
or U16086 (N_16086,N_15864,N_15959);
nor U16087 (N_16087,N_15908,N_15894);
xnor U16088 (N_16088,N_15929,N_15881);
nor U16089 (N_16089,N_15862,N_15960);
nand U16090 (N_16090,N_15900,N_15906);
and U16091 (N_16091,N_15893,N_15926);
nor U16092 (N_16092,N_15967,N_15872);
xor U16093 (N_16093,N_15940,N_15947);
nand U16094 (N_16094,N_15916,N_15847);
xnor U16095 (N_16095,N_15897,N_15959);
xnor U16096 (N_16096,N_15952,N_15856);
and U16097 (N_16097,N_15863,N_15926);
xor U16098 (N_16098,N_15977,N_15949);
or U16099 (N_16099,N_15842,N_15946);
nor U16100 (N_16100,N_15864,N_15861);
nand U16101 (N_16101,N_15989,N_15939);
xnor U16102 (N_16102,N_15958,N_15866);
xnor U16103 (N_16103,N_15908,N_15921);
xnor U16104 (N_16104,N_15988,N_15900);
xor U16105 (N_16105,N_15845,N_15927);
or U16106 (N_16106,N_15901,N_15850);
and U16107 (N_16107,N_15894,N_15980);
nand U16108 (N_16108,N_15968,N_15983);
or U16109 (N_16109,N_15889,N_15947);
xor U16110 (N_16110,N_15902,N_15970);
and U16111 (N_16111,N_15902,N_15876);
xor U16112 (N_16112,N_15926,N_15961);
or U16113 (N_16113,N_15856,N_15847);
nor U16114 (N_16114,N_15940,N_15992);
nor U16115 (N_16115,N_15844,N_15890);
and U16116 (N_16116,N_15915,N_15880);
and U16117 (N_16117,N_15898,N_15866);
nor U16118 (N_16118,N_15975,N_15948);
xnor U16119 (N_16119,N_15960,N_15878);
nor U16120 (N_16120,N_15980,N_15988);
nor U16121 (N_16121,N_15972,N_15884);
xnor U16122 (N_16122,N_15976,N_15856);
nand U16123 (N_16123,N_15917,N_15931);
nand U16124 (N_16124,N_15952,N_15872);
xnor U16125 (N_16125,N_15928,N_15959);
xor U16126 (N_16126,N_15991,N_15869);
nor U16127 (N_16127,N_15884,N_15899);
nor U16128 (N_16128,N_15882,N_15872);
nor U16129 (N_16129,N_15957,N_15900);
nand U16130 (N_16130,N_15885,N_15925);
or U16131 (N_16131,N_15891,N_15961);
or U16132 (N_16132,N_15957,N_15942);
or U16133 (N_16133,N_15978,N_15856);
nand U16134 (N_16134,N_15841,N_15935);
and U16135 (N_16135,N_15933,N_15985);
nor U16136 (N_16136,N_15862,N_15988);
nand U16137 (N_16137,N_15944,N_15966);
xor U16138 (N_16138,N_15950,N_15853);
or U16139 (N_16139,N_15907,N_15986);
and U16140 (N_16140,N_15924,N_15941);
nand U16141 (N_16141,N_15916,N_15981);
nor U16142 (N_16142,N_15919,N_15931);
xor U16143 (N_16143,N_15976,N_15840);
and U16144 (N_16144,N_15985,N_15851);
nor U16145 (N_16145,N_15973,N_15989);
nand U16146 (N_16146,N_15956,N_15901);
nand U16147 (N_16147,N_15850,N_15913);
or U16148 (N_16148,N_15936,N_15955);
or U16149 (N_16149,N_15956,N_15947);
nor U16150 (N_16150,N_15981,N_15911);
nor U16151 (N_16151,N_15872,N_15971);
xor U16152 (N_16152,N_15992,N_15996);
nor U16153 (N_16153,N_15876,N_15956);
or U16154 (N_16154,N_15913,N_15909);
nor U16155 (N_16155,N_15840,N_15953);
xor U16156 (N_16156,N_15854,N_15876);
nand U16157 (N_16157,N_15888,N_15874);
nor U16158 (N_16158,N_15926,N_15956);
and U16159 (N_16159,N_15993,N_15954);
nor U16160 (N_16160,N_16020,N_16027);
or U16161 (N_16161,N_16131,N_16123);
xnor U16162 (N_16162,N_16074,N_16143);
nand U16163 (N_16163,N_16121,N_16099);
xnor U16164 (N_16164,N_16033,N_16073);
nand U16165 (N_16165,N_16114,N_16103);
nand U16166 (N_16166,N_16015,N_16034);
and U16167 (N_16167,N_16079,N_16064);
and U16168 (N_16168,N_16060,N_16000);
nor U16169 (N_16169,N_16050,N_16130);
nand U16170 (N_16170,N_16117,N_16093);
nor U16171 (N_16171,N_16051,N_16148);
nand U16172 (N_16172,N_16001,N_16155);
xor U16173 (N_16173,N_16014,N_16048);
nand U16174 (N_16174,N_16151,N_16030);
nand U16175 (N_16175,N_16055,N_16021);
or U16176 (N_16176,N_16141,N_16107);
nor U16177 (N_16177,N_16044,N_16157);
nor U16178 (N_16178,N_16084,N_16115);
xnor U16179 (N_16179,N_16111,N_16106);
xnor U16180 (N_16180,N_16108,N_16012);
nor U16181 (N_16181,N_16072,N_16126);
nor U16182 (N_16182,N_16152,N_16009);
and U16183 (N_16183,N_16156,N_16004);
and U16184 (N_16184,N_16045,N_16092);
nor U16185 (N_16185,N_16153,N_16023);
or U16186 (N_16186,N_16049,N_16081);
and U16187 (N_16187,N_16005,N_16052);
nor U16188 (N_16188,N_16019,N_16031);
xnor U16189 (N_16189,N_16071,N_16142);
xnor U16190 (N_16190,N_16085,N_16075);
nand U16191 (N_16191,N_16007,N_16042);
nor U16192 (N_16192,N_16083,N_16017);
xor U16193 (N_16193,N_16088,N_16119);
nand U16194 (N_16194,N_16137,N_16102);
or U16195 (N_16195,N_16006,N_16101);
nand U16196 (N_16196,N_16016,N_16035);
and U16197 (N_16197,N_16150,N_16089);
or U16198 (N_16198,N_16100,N_16149);
or U16199 (N_16199,N_16145,N_16138);
nor U16200 (N_16200,N_16080,N_16022);
or U16201 (N_16201,N_16011,N_16109);
or U16202 (N_16202,N_16038,N_16046);
or U16203 (N_16203,N_16037,N_16120);
nand U16204 (N_16204,N_16010,N_16002);
or U16205 (N_16205,N_16139,N_16024);
or U16206 (N_16206,N_16082,N_16062);
nor U16207 (N_16207,N_16122,N_16159);
or U16208 (N_16208,N_16094,N_16118);
nor U16209 (N_16209,N_16066,N_16090);
and U16210 (N_16210,N_16147,N_16032);
xnor U16211 (N_16211,N_16132,N_16029);
and U16212 (N_16212,N_16095,N_16128);
xnor U16213 (N_16213,N_16056,N_16047);
nand U16214 (N_16214,N_16069,N_16036);
or U16215 (N_16215,N_16076,N_16070);
or U16216 (N_16216,N_16065,N_16058);
nor U16217 (N_16217,N_16113,N_16098);
nor U16218 (N_16218,N_16008,N_16144);
or U16219 (N_16219,N_16135,N_16134);
nor U16220 (N_16220,N_16054,N_16061);
xnor U16221 (N_16221,N_16105,N_16091);
xnor U16222 (N_16222,N_16158,N_16028);
nand U16223 (N_16223,N_16125,N_16146);
xnor U16224 (N_16224,N_16043,N_16154);
nor U16225 (N_16225,N_16039,N_16025);
nor U16226 (N_16226,N_16124,N_16133);
xor U16227 (N_16227,N_16040,N_16053);
xor U16228 (N_16228,N_16041,N_16018);
nor U16229 (N_16229,N_16003,N_16068);
and U16230 (N_16230,N_16078,N_16127);
and U16231 (N_16231,N_16110,N_16140);
nor U16232 (N_16232,N_16096,N_16112);
nand U16233 (N_16233,N_16104,N_16057);
or U16234 (N_16234,N_16086,N_16077);
nor U16235 (N_16235,N_16013,N_16136);
nor U16236 (N_16236,N_16097,N_16129);
nor U16237 (N_16237,N_16059,N_16063);
xor U16238 (N_16238,N_16116,N_16067);
nor U16239 (N_16239,N_16026,N_16087);
nor U16240 (N_16240,N_16044,N_16112);
nand U16241 (N_16241,N_16066,N_16109);
xnor U16242 (N_16242,N_16150,N_16155);
xnor U16243 (N_16243,N_16071,N_16011);
or U16244 (N_16244,N_16032,N_16001);
nor U16245 (N_16245,N_16004,N_16141);
nor U16246 (N_16246,N_16118,N_16071);
or U16247 (N_16247,N_16128,N_16064);
xor U16248 (N_16248,N_16086,N_16144);
nand U16249 (N_16249,N_16125,N_16081);
and U16250 (N_16250,N_16062,N_16045);
nor U16251 (N_16251,N_16009,N_16136);
or U16252 (N_16252,N_16006,N_16042);
nor U16253 (N_16253,N_16045,N_16097);
and U16254 (N_16254,N_16055,N_16048);
xnor U16255 (N_16255,N_16000,N_16107);
and U16256 (N_16256,N_16011,N_16043);
xnor U16257 (N_16257,N_16124,N_16114);
and U16258 (N_16258,N_16122,N_16043);
nand U16259 (N_16259,N_16133,N_16080);
and U16260 (N_16260,N_16033,N_16074);
or U16261 (N_16261,N_16045,N_16023);
nand U16262 (N_16262,N_16070,N_16146);
nand U16263 (N_16263,N_16111,N_16047);
nand U16264 (N_16264,N_16052,N_16045);
nand U16265 (N_16265,N_16136,N_16131);
xnor U16266 (N_16266,N_16007,N_16018);
or U16267 (N_16267,N_16086,N_16015);
xnor U16268 (N_16268,N_16137,N_16052);
and U16269 (N_16269,N_16059,N_16035);
xor U16270 (N_16270,N_16099,N_16098);
xor U16271 (N_16271,N_16025,N_16092);
nor U16272 (N_16272,N_16059,N_16001);
and U16273 (N_16273,N_16123,N_16056);
or U16274 (N_16274,N_16025,N_16091);
nand U16275 (N_16275,N_16119,N_16030);
nand U16276 (N_16276,N_16118,N_16153);
and U16277 (N_16277,N_16141,N_16112);
xor U16278 (N_16278,N_16069,N_16087);
and U16279 (N_16279,N_16052,N_16038);
and U16280 (N_16280,N_16036,N_16080);
or U16281 (N_16281,N_16150,N_16093);
nor U16282 (N_16282,N_16067,N_16027);
xor U16283 (N_16283,N_16029,N_16110);
xnor U16284 (N_16284,N_16121,N_16007);
and U16285 (N_16285,N_16039,N_16060);
nor U16286 (N_16286,N_16143,N_16009);
or U16287 (N_16287,N_16001,N_16102);
and U16288 (N_16288,N_16036,N_16046);
xor U16289 (N_16289,N_16045,N_16021);
xnor U16290 (N_16290,N_16039,N_16150);
nand U16291 (N_16291,N_16154,N_16145);
xor U16292 (N_16292,N_16008,N_16111);
and U16293 (N_16293,N_16135,N_16022);
nand U16294 (N_16294,N_16156,N_16018);
or U16295 (N_16295,N_16064,N_16002);
nand U16296 (N_16296,N_16065,N_16158);
or U16297 (N_16297,N_16090,N_16128);
xor U16298 (N_16298,N_16023,N_16075);
nand U16299 (N_16299,N_16010,N_16008);
and U16300 (N_16300,N_16007,N_16005);
or U16301 (N_16301,N_16153,N_16134);
and U16302 (N_16302,N_16017,N_16113);
nor U16303 (N_16303,N_16086,N_16049);
nand U16304 (N_16304,N_16013,N_16123);
nand U16305 (N_16305,N_16140,N_16114);
and U16306 (N_16306,N_16139,N_16029);
nand U16307 (N_16307,N_16051,N_16135);
and U16308 (N_16308,N_16000,N_16141);
xnor U16309 (N_16309,N_16056,N_16119);
nor U16310 (N_16310,N_16081,N_16031);
xor U16311 (N_16311,N_16109,N_16077);
and U16312 (N_16312,N_16080,N_16037);
xor U16313 (N_16313,N_16128,N_16005);
xor U16314 (N_16314,N_16060,N_16120);
xor U16315 (N_16315,N_16155,N_16032);
and U16316 (N_16316,N_16068,N_16005);
and U16317 (N_16317,N_16145,N_16026);
and U16318 (N_16318,N_16100,N_16145);
nand U16319 (N_16319,N_16101,N_16057);
xnor U16320 (N_16320,N_16239,N_16294);
and U16321 (N_16321,N_16272,N_16305);
or U16322 (N_16322,N_16308,N_16309);
nand U16323 (N_16323,N_16303,N_16186);
and U16324 (N_16324,N_16185,N_16285);
nand U16325 (N_16325,N_16189,N_16219);
nand U16326 (N_16326,N_16302,N_16223);
xor U16327 (N_16327,N_16177,N_16298);
nand U16328 (N_16328,N_16292,N_16266);
nor U16329 (N_16329,N_16237,N_16276);
nand U16330 (N_16330,N_16288,N_16280);
nand U16331 (N_16331,N_16233,N_16240);
and U16332 (N_16332,N_16284,N_16174);
and U16333 (N_16333,N_16307,N_16290);
nand U16334 (N_16334,N_16318,N_16163);
and U16335 (N_16335,N_16204,N_16317);
nor U16336 (N_16336,N_16169,N_16254);
or U16337 (N_16337,N_16218,N_16238);
nand U16338 (N_16338,N_16224,N_16214);
or U16339 (N_16339,N_16241,N_16282);
and U16340 (N_16340,N_16226,N_16275);
nor U16341 (N_16341,N_16242,N_16262);
and U16342 (N_16342,N_16197,N_16182);
xor U16343 (N_16343,N_16183,N_16304);
and U16344 (N_16344,N_16230,N_16210);
or U16345 (N_16345,N_16180,N_16217);
and U16346 (N_16346,N_16194,N_16313);
nand U16347 (N_16347,N_16175,N_16221);
nor U16348 (N_16348,N_16289,N_16193);
or U16349 (N_16349,N_16301,N_16206);
nor U16350 (N_16350,N_16190,N_16192);
or U16351 (N_16351,N_16267,N_16273);
or U16352 (N_16352,N_16184,N_16311);
and U16353 (N_16353,N_16249,N_16203);
nor U16354 (N_16354,N_16231,N_16209);
nand U16355 (N_16355,N_16167,N_16283);
xor U16356 (N_16356,N_16235,N_16220);
nand U16357 (N_16357,N_16176,N_16227);
and U16358 (N_16358,N_16168,N_16271);
xnor U16359 (N_16359,N_16312,N_16306);
nand U16360 (N_16360,N_16281,N_16222);
and U16361 (N_16361,N_16314,N_16248);
nor U16362 (N_16362,N_16202,N_16256);
nand U16363 (N_16363,N_16232,N_16161);
nor U16364 (N_16364,N_16244,N_16315);
xnor U16365 (N_16365,N_16251,N_16246);
nand U16366 (N_16366,N_16173,N_16212);
and U16367 (N_16367,N_16236,N_16205);
nor U16368 (N_16368,N_16171,N_16179);
nor U16369 (N_16369,N_16181,N_16234);
or U16370 (N_16370,N_16274,N_16287);
nor U16371 (N_16371,N_16247,N_16293);
or U16372 (N_16372,N_16198,N_16188);
nand U16373 (N_16373,N_16257,N_16208);
or U16374 (N_16374,N_16196,N_16291);
xnor U16375 (N_16375,N_16228,N_16259);
and U16376 (N_16376,N_16178,N_16263);
nand U16377 (N_16377,N_16172,N_16191);
nand U16378 (N_16378,N_16200,N_16162);
xnor U16379 (N_16379,N_16253,N_16300);
xnor U16380 (N_16380,N_16215,N_16299);
and U16381 (N_16381,N_16211,N_16310);
nand U16382 (N_16382,N_16243,N_16195);
and U16383 (N_16383,N_16277,N_16319);
and U16384 (N_16384,N_16160,N_16250);
xnor U16385 (N_16385,N_16165,N_16213);
xnor U16386 (N_16386,N_16225,N_16264);
nand U16387 (N_16387,N_16269,N_16260);
or U16388 (N_16388,N_16270,N_16258);
or U16389 (N_16389,N_16187,N_16216);
and U16390 (N_16390,N_16296,N_16316);
or U16391 (N_16391,N_16207,N_16295);
xor U16392 (N_16392,N_16255,N_16166);
nand U16393 (N_16393,N_16286,N_16268);
nand U16394 (N_16394,N_16199,N_16265);
or U16395 (N_16395,N_16297,N_16245);
or U16396 (N_16396,N_16261,N_16164);
xor U16397 (N_16397,N_16170,N_16279);
xnor U16398 (N_16398,N_16229,N_16252);
or U16399 (N_16399,N_16201,N_16278);
or U16400 (N_16400,N_16289,N_16259);
xor U16401 (N_16401,N_16166,N_16311);
nor U16402 (N_16402,N_16292,N_16175);
nor U16403 (N_16403,N_16172,N_16171);
nand U16404 (N_16404,N_16162,N_16258);
xnor U16405 (N_16405,N_16239,N_16206);
nor U16406 (N_16406,N_16317,N_16276);
nand U16407 (N_16407,N_16188,N_16200);
and U16408 (N_16408,N_16172,N_16257);
xnor U16409 (N_16409,N_16253,N_16274);
or U16410 (N_16410,N_16241,N_16239);
xor U16411 (N_16411,N_16254,N_16296);
and U16412 (N_16412,N_16184,N_16278);
and U16413 (N_16413,N_16214,N_16311);
nand U16414 (N_16414,N_16275,N_16270);
or U16415 (N_16415,N_16296,N_16299);
xnor U16416 (N_16416,N_16218,N_16247);
or U16417 (N_16417,N_16296,N_16291);
nor U16418 (N_16418,N_16288,N_16216);
nand U16419 (N_16419,N_16175,N_16187);
or U16420 (N_16420,N_16177,N_16287);
nand U16421 (N_16421,N_16294,N_16240);
xnor U16422 (N_16422,N_16295,N_16222);
xnor U16423 (N_16423,N_16269,N_16266);
and U16424 (N_16424,N_16219,N_16198);
or U16425 (N_16425,N_16306,N_16181);
nor U16426 (N_16426,N_16317,N_16203);
nor U16427 (N_16427,N_16296,N_16248);
nand U16428 (N_16428,N_16197,N_16178);
nor U16429 (N_16429,N_16297,N_16232);
nor U16430 (N_16430,N_16287,N_16229);
nor U16431 (N_16431,N_16285,N_16160);
or U16432 (N_16432,N_16255,N_16224);
and U16433 (N_16433,N_16258,N_16170);
xor U16434 (N_16434,N_16221,N_16179);
or U16435 (N_16435,N_16289,N_16278);
xor U16436 (N_16436,N_16241,N_16250);
nand U16437 (N_16437,N_16269,N_16254);
or U16438 (N_16438,N_16232,N_16307);
nor U16439 (N_16439,N_16205,N_16183);
xor U16440 (N_16440,N_16242,N_16315);
or U16441 (N_16441,N_16273,N_16226);
nand U16442 (N_16442,N_16214,N_16313);
xor U16443 (N_16443,N_16272,N_16239);
nor U16444 (N_16444,N_16251,N_16279);
nand U16445 (N_16445,N_16164,N_16228);
nand U16446 (N_16446,N_16264,N_16198);
or U16447 (N_16447,N_16257,N_16259);
nand U16448 (N_16448,N_16282,N_16267);
nor U16449 (N_16449,N_16231,N_16264);
nor U16450 (N_16450,N_16208,N_16222);
or U16451 (N_16451,N_16271,N_16282);
xnor U16452 (N_16452,N_16168,N_16229);
nand U16453 (N_16453,N_16222,N_16170);
nand U16454 (N_16454,N_16245,N_16163);
xor U16455 (N_16455,N_16276,N_16164);
and U16456 (N_16456,N_16286,N_16275);
nand U16457 (N_16457,N_16219,N_16217);
nand U16458 (N_16458,N_16263,N_16287);
or U16459 (N_16459,N_16239,N_16269);
nor U16460 (N_16460,N_16264,N_16273);
xnor U16461 (N_16461,N_16214,N_16218);
and U16462 (N_16462,N_16251,N_16309);
or U16463 (N_16463,N_16207,N_16273);
nand U16464 (N_16464,N_16206,N_16316);
xnor U16465 (N_16465,N_16296,N_16288);
nand U16466 (N_16466,N_16288,N_16228);
xor U16467 (N_16467,N_16226,N_16256);
xnor U16468 (N_16468,N_16312,N_16227);
xnor U16469 (N_16469,N_16223,N_16278);
nor U16470 (N_16470,N_16230,N_16308);
xnor U16471 (N_16471,N_16290,N_16246);
nor U16472 (N_16472,N_16183,N_16261);
nand U16473 (N_16473,N_16235,N_16294);
or U16474 (N_16474,N_16295,N_16276);
nor U16475 (N_16475,N_16319,N_16258);
nand U16476 (N_16476,N_16244,N_16245);
or U16477 (N_16477,N_16231,N_16193);
or U16478 (N_16478,N_16235,N_16305);
xor U16479 (N_16479,N_16251,N_16310);
and U16480 (N_16480,N_16388,N_16450);
and U16481 (N_16481,N_16395,N_16375);
or U16482 (N_16482,N_16337,N_16446);
or U16483 (N_16483,N_16336,N_16374);
nand U16484 (N_16484,N_16402,N_16370);
nand U16485 (N_16485,N_16349,N_16438);
and U16486 (N_16486,N_16361,N_16340);
nand U16487 (N_16487,N_16398,N_16386);
or U16488 (N_16488,N_16334,N_16327);
nand U16489 (N_16489,N_16472,N_16382);
or U16490 (N_16490,N_16320,N_16416);
and U16491 (N_16491,N_16444,N_16366);
and U16492 (N_16492,N_16471,N_16476);
nand U16493 (N_16493,N_16325,N_16420);
nand U16494 (N_16494,N_16479,N_16379);
or U16495 (N_16495,N_16335,N_16412);
or U16496 (N_16496,N_16463,N_16469);
nor U16497 (N_16497,N_16397,N_16474);
or U16498 (N_16498,N_16372,N_16356);
or U16499 (N_16499,N_16385,N_16467);
nand U16500 (N_16500,N_16433,N_16451);
nor U16501 (N_16501,N_16363,N_16437);
nand U16502 (N_16502,N_16460,N_16442);
and U16503 (N_16503,N_16464,N_16443);
or U16504 (N_16504,N_16459,N_16404);
nor U16505 (N_16505,N_16411,N_16330);
xor U16506 (N_16506,N_16400,N_16371);
nor U16507 (N_16507,N_16345,N_16415);
and U16508 (N_16508,N_16351,N_16454);
nor U16509 (N_16509,N_16339,N_16458);
or U16510 (N_16510,N_16425,N_16429);
xnor U16511 (N_16511,N_16419,N_16473);
and U16512 (N_16512,N_16417,N_16468);
nor U16513 (N_16513,N_16403,N_16440);
nor U16514 (N_16514,N_16383,N_16405);
and U16515 (N_16515,N_16323,N_16428);
or U16516 (N_16516,N_16427,N_16389);
nor U16517 (N_16517,N_16324,N_16399);
xor U16518 (N_16518,N_16431,N_16392);
and U16519 (N_16519,N_16434,N_16462);
xnor U16520 (N_16520,N_16384,N_16346);
nor U16521 (N_16521,N_16430,N_16461);
nand U16522 (N_16522,N_16341,N_16401);
or U16523 (N_16523,N_16360,N_16477);
nor U16524 (N_16524,N_16377,N_16328);
xnor U16525 (N_16525,N_16435,N_16338);
nor U16526 (N_16526,N_16364,N_16432);
nor U16527 (N_16527,N_16390,N_16391);
nand U16528 (N_16528,N_16453,N_16414);
xnor U16529 (N_16529,N_16466,N_16343);
nor U16530 (N_16530,N_16394,N_16342);
and U16531 (N_16531,N_16322,N_16449);
xnor U16532 (N_16532,N_16457,N_16424);
nor U16533 (N_16533,N_16448,N_16423);
and U16534 (N_16534,N_16354,N_16376);
nand U16535 (N_16535,N_16441,N_16406);
nand U16536 (N_16536,N_16413,N_16378);
nor U16537 (N_16537,N_16465,N_16409);
nor U16538 (N_16538,N_16381,N_16352);
and U16539 (N_16539,N_16353,N_16445);
nor U16540 (N_16540,N_16359,N_16408);
nor U16541 (N_16541,N_16332,N_16365);
nand U16542 (N_16542,N_16367,N_16407);
nand U16543 (N_16543,N_16348,N_16439);
nor U16544 (N_16544,N_16455,N_16393);
xnor U16545 (N_16545,N_16358,N_16426);
nand U16546 (N_16546,N_16410,N_16421);
and U16547 (N_16547,N_16362,N_16396);
xnor U16548 (N_16548,N_16321,N_16478);
and U16549 (N_16549,N_16369,N_16368);
xor U16550 (N_16550,N_16387,N_16326);
nand U16551 (N_16551,N_16347,N_16329);
nor U16552 (N_16552,N_16475,N_16373);
nor U16553 (N_16553,N_16452,N_16357);
nand U16554 (N_16554,N_16418,N_16380);
nor U16555 (N_16555,N_16456,N_16344);
xnor U16556 (N_16556,N_16470,N_16331);
and U16557 (N_16557,N_16355,N_16333);
xor U16558 (N_16558,N_16436,N_16447);
nand U16559 (N_16559,N_16422,N_16350);
and U16560 (N_16560,N_16357,N_16393);
or U16561 (N_16561,N_16476,N_16472);
nand U16562 (N_16562,N_16429,N_16342);
or U16563 (N_16563,N_16360,N_16458);
xor U16564 (N_16564,N_16335,N_16455);
xnor U16565 (N_16565,N_16462,N_16377);
nor U16566 (N_16566,N_16408,N_16379);
and U16567 (N_16567,N_16416,N_16378);
and U16568 (N_16568,N_16421,N_16398);
xnor U16569 (N_16569,N_16416,N_16361);
xnor U16570 (N_16570,N_16325,N_16402);
or U16571 (N_16571,N_16373,N_16338);
xnor U16572 (N_16572,N_16354,N_16339);
nand U16573 (N_16573,N_16405,N_16328);
or U16574 (N_16574,N_16439,N_16354);
nor U16575 (N_16575,N_16335,N_16407);
xnor U16576 (N_16576,N_16325,N_16361);
nor U16577 (N_16577,N_16443,N_16376);
or U16578 (N_16578,N_16456,N_16432);
nor U16579 (N_16579,N_16428,N_16350);
or U16580 (N_16580,N_16384,N_16424);
nor U16581 (N_16581,N_16428,N_16361);
or U16582 (N_16582,N_16324,N_16454);
nor U16583 (N_16583,N_16344,N_16360);
and U16584 (N_16584,N_16331,N_16378);
or U16585 (N_16585,N_16343,N_16321);
xnor U16586 (N_16586,N_16449,N_16425);
and U16587 (N_16587,N_16396,N_16471);
nor U16588 (N_16588,N_16437,N_16401);
xnor U16589 (N_16589,N_16365,N_16460);
nor U16590 (N_16590,N_16327,N_16394);
and U16591 (N_16591,N_16331,N_16384);
or U16592 (N_16592,N_16392,N_16368);
and U16593 (N_16593,N_16387,N_16381);
nand U16594 (N_16594,N_16469,N_16473);
and U16595 (N_16595,N_16455,N_16466);
nor U16596 (N_16596,N_16441,N_16421);
nand U16597 (N_16597,N_16360,N_16419);
or U16598 (N_16598,N_16355,N_16375);
and U16599 (N_16599,N_16446,N_16386);
nor U16600 (N_16600,N_16421,N_16358);
and U16601 (N_16601,N_16419,N_16380);
nand U16602 (N_16602,N_16388,N_16419);
or U16603 (N_16603,N_16372,N_16328);
xor U16604 (N_16604,N_16451,N_16375);
or U16605 (N_16605,N_16398,N_16407);
or U16606 (N_16606,N_16460,N_16415);
or U16607 (N_16607,N_16456,N_16380);
xnor U16608 (N_16608,N_16341,N_16423);
nor U16609 (N_16609,N_16346,N_16347);
nor U16610 (N_16610,N_16478,N_16433);
nand U16611 (N_16611,N_16414,N_16320);
and U16612 (N_16612,N_16428,N_16365);
xnor U16613 (N_16613,N_16347,N_16417);
or U16614 (N_16614,N_16359,N_16380);
and U16615 (N_16615,N_16347,N_16460);
xor U16616 (N_16616,N_16381,N_16441);
and U16617 (N_16617,N_16320,N_16452);
xor U16618 (N_16618,N_16476,N_16383);
nor U16619 (N_16619,N_16418,N_16347);
xor U16620 (N_16620,N_16464,N_16412);
or U16621 (N_16621,N_16436,N_16413);
xor U16622 (N_16622,N_16339,N_16479);
and U16623 (N_16623,N_16421,N_16335);
nand U16624 (N_16624,N_16463,N_16443);
nor U16625 (N_16625,N_16371,N_16337);
or U16626 (N_16626,N_16417,N_16448);
and U16627 (N_16627,N_16399,N_16322);
xor U16628 (N_16628,N_16429,N_16381);
xnor U16629 (N_16629,N_16321,N_16470);
and U16630 (N_16630,N_16426,N_16431);
xnor U16631 (N_16631,N_16462,N_16326);
and U16632 (N_16632,N_16381,N_16434);
nand U16633 (N_16633,N_16331,N_16456);
nand U16634 (N_16634,N_16381,N_16351);
or U16635 (N_16635,N_16454,N_16439);
xor U16636 (N_16636,N_16436,N_16325);
and U16637 (N_16637,N_16330,N_16466);
nand U16638 (N_16638,N_16438,N_16359);
nor U16639 (N_16639,N_16383,N_16464);
nand U16640 (N_16640,N_16494,N_16630);
or U16641 (N_16641,N_16505,N_16486);
nor U16642 (N_16642,N_16536,N_16523);
xor U16643 (N_16643,N_16632,N_16490);
nor U16644 (N_16644,N_16568,N_16508);
nand U16645 (N_16645,N_16579,N_16537);
and U16646 (N_16646,N_16495,N_16620);
nor U16647 (N_16647,N_16542,N_16511);
nand U16648 (N_16648,N_16501,N_16482);
nor U16649 (N_16649,N_16637,N_16598);
or U16650 (N_16650,N_16577,N_16563);
nand U16651 (N_16651,N_16496,N_16565);
nor U16652 (N_16652,N_16625,N_16609);
or U16653 (N_16653,N_16507,N_16531);
xor U16654 (N_16654,N_16610,N_16618);
nand U16655 (N_16655,N_16556,N_16627);
or U16656 (N_16656,N_16533,N_16596);
and U16657 (N_16657,N_16592,N_16607);
or U16658 (N_16658,N_16564,N_16539);
or U16659 (N_16659,N_16639,N_16619);
or U16660 (N_16660,N_16535,N_16510);
nand U16661 (N_16661,N_16498,N_16546);
or U16662 (N_16662,N_16480,N_16540);
nor U16663 (N_16663,N_16597,N_16572);
xnor U16664 (N_16664,N_16558,N_16584);
nand U16665 (N_16665,N_16624,N_16551);
xor U16666 (N_16666,N_16608,N_16541);
or U16667 (N_16667,N_16562,N_16509);
and U16668 (N_16668,N_16599,N_16487);
nand U16669 (N_16669,N_16555,N_16493);
nand U16670 (N_16670,N_16634,N_16524);
or U16671 (N_16671,N_16525,N_16603);
nand U16672 (N_16672,N_16512,N_16553);
and U16673 (N_16673,N_16623,N_16600);
and U16674 (N_16674,N_16491,N_16485);
nor U16675 (N_16675,N_16506,N_16514);
xnor U16676 (N_16676,N_16517,N_16571);
xnor U16677 (N_16677,N_16566,N_16518);
xnor U16678 (N_16678,N_16529,N_16586);
xor U16679 (N_16679,N_16612,N_16628);
nor U16680 (N_16680,N_16595,N_16616);
or U16681 (N_16681,N_16538,N_16549);
and U16682 (N_16682,N_16513,N_16500);
xnor U16683 (N_16683,N_16545,N_16589);
nor U16684 (N_16684,N_16527,N_16578);
nor U16685 (N_16685,N_16483,N_16526);
nor U16686 (N_16686,N_16521,N_16499);
nand U16687 (N_16687,N_16590,N_16534);
or U16688 (N_16688,N_16488,N_16629);
xnor U16689 (N_16689,N_16593,N_16548);
or U16690 (N_16690,N_16583,N_16606);
and U16691 (N_16691,N_16515,N_16638);
and U16692 (N_16692,N_16560,N_16587);
or U16693 (N_16693,N_16503,N_16613);
nand U16694 (N_16694,N_16622,N_16516);
or U16695 (N_16695,N_16615,N_16561);
xor U16696 (N_16696,N_16626,N_16636);
and U16697 (N_16697,N_16481,N_16614);
or U16698 (N_16698,N_16582,N_16573);
xor U16699 (N_16699,N_16575,N_16631);
and U16700 (N_16700,N_16557,N_16497);
nand U16701 (N_16701,N_16504,N_16532);
nor U16702 (N_16702,N_16617,N_16611);
nand U16703 (N_16703,N_16594,N_16552);
xor U16704 (N_16704,N_16570,N_16492);
xnor U16705 (N_16705,N_16519,N_16522);
and U16706 (N_16706,N_16574,N_16559);
or U16707 (N_16707,N_16591,N_16520);
or U16708 (N_16708,N_16605,N_16544);
or U16709 (N_16709,N_16530,N_16621);
nand U16710 (N_16710,N_16567,N_16554);
or U16711 (N_16711,N_16588,N_16581);
nand U16712 (N_16712,N_16547,N_16484);
nor U16713 (N_16713,N_16569,N_16602);
and U16714 (N_16714,N_16604,N_16585);
nor U16715 (N_16715,N_16528,N_16489);
nand U16716 (N_16716,N_16543,N_16550);
and U16717 (N_16717,N_16576,N_16633);
xnor U16718 (N_16718,N_16635,N_16580);
and U16719 (N_16719,N_16502,N_16601);
or U16720 (N_16720,N_16606,N_16491);
xor U16721 (N_16721,N_16571,N_16498);
or U16722 (N_16722,N_16483,N_16597);
nor U16723 (N_16723,N_16540,N_16626);
or U16724 (N_16724,N_16613,N_16481);
and U16725 (N_16725,N_16599,N_16526);
and U16726 (N_16726,N_16617,N_16565);
xor U16727 (N_16727,N_16520,N_16630);
xnor U16728 (N_16728,N_16599,N_16598);
nor U16729 (N_16729,N_16526,N_16629);
or U16730 (N_16730,N_16565,N_16555);
and U16731 (N_16731,N_16627,N_16541);
xnor U16732 (N_16732,N_16568,N_16489);
or U16733 (N_16733,N_16630,N_16580);
nor U16734 (N_16734,N_16542,N_16585);
or U16735 (N_16735,N_16542,N_16573);
nand U16736 (N_16736,N_16617,N_16503);
nor U16737 (N_16737,N_16604,N_16493);
or U16738 (N_16738,N_16487,N_16605);
and U16739 (N_16739,N_16527,N_16576);
nor U16740 (N_16740,N_16606,N_16565);
nor U16741 (N_16741,N_16613,N_16620);
nor U16742 (N_16742,N_16558,N_16516);
nor U16743 (N_16743,N_16627,N_16601);
or U16744 (N_16744,N_16607,N_16517);
nand U16745 (N_16745,N_16563,N_16582);
and U16746 (N_16746,N_16637,N_16633);
and U16747 (N_16747,N_16517,N_16623);
nor U16748 (N_16748,N_16550,N_16594);
nand U16749 (N_16749,N_16509,N_16511);
nor U16750 (N_16750,N_16611,N_16533);
and U16751 (N_16751,N_16601,N_16531);
or U16752 (N_16752,N_16526,N_16630);
nor U16753 (N_16753,N_16622,N_16558);
or U16754 (N_16754,N_16564,N_16560);
or U16755 (N_16755,N_16529,N_16505);
nand U16756 (N_16756,N_16514,N_16541);
and U16757 (N_16757,N_16507,N_16560);
nand U16758 (N_16758,N_16508,N_16625);
nand U16759 (N_16759,N_16501,N_16520);
xor U16760 (N_16760,N_16604,N_16506);
and U16761 (N_16761,N_16626,N_16523);
xnor U16762 (N_16762,N_16613,N_16504);
nand U16763 (N_16763,N_16486,N_16508);
and U16764 (N_16764,N_16501,N_16586);
and U16765 (N_16765,N_16626,N_16571);
nand U16766 (N_16766,N_16497,N_16603);
or U16767 (N_16767,N_16568,N_16556);
nor U16768 (N_16768,N_16609,N_16637);
nor U16769 (N_16769,N_16534,N_16548);
and U16770 (N_16770,N_16565,N_16543);
nand U16771 (N_16771,N_16566,N_16551);
xnor U16772 (N_16772,N_16559,N_16508);
nor U16773 (N_16773,N_16625,N_16530);
nor U16774 (N_16774,N_16572,N_16497);
xnor U16775 (N_16775,N_16569,N_16511);
xor U16776 (N_16776,N_16492,N_16501);
nand U16777 (N_16777,N_16607,N_16632);
nand U16778 (N_16778,N_16590,N_16624);
nand U16779 (N_16779,N_16553,N_16519);
nand U16780 (N_16780,N_16631,N_16486);
xnor U16781 (N_16781,N_16526,N_16578);
xor U16782 (N_16782,N_16480,N_16572);
nor U16783 (N_16783,N_16585,N_16615);
and U16784 (N_16784,N_16622,N_16522);
nor U16785 (N_16785,N_16588,N_16529);
nor U16786 (N_16786,N_16543,N_16522);
nand U16787 (N_16787,N_16585,N_16630);
or U16788 (N_16788,N_16572,N_16518);
or U16789 (N_16789,N_16592,N_16527);
and U16790 (N_16790,N_16556,N_16637);
xor U16791 (N_16791,N_16576,N_16639);
nor U16792 (N_16792,N_16611,N_16590);
nor U16793 (N_16793,N_16595,N_16607);
nor U16794 (N_16794,N_16568,N_16537);
and U16795 (N_16795,N_16638,N_16611);
and U16796 (N_16796,N_16554,N_16581);
and U16797 (N_16797,N_16603,N_16582);
xor U16798 (N_16798,N_16630,N_16609);
nor U16799 (N_16799,N_16560,N_16510);
xnor U16800 (N_16800,N_16683,N_16665);
nor U16801 (N_16801,N_16795,N_16717);
nor U16802 (N_16802,N_16725,N_16744);
and U16803 (N_16803,N_16739,N_16648);
and U16804 (N_16804,N_16712,N_16729);
xnor U16805 (N_16805,N_16760,N_16669);
or U16806 (N_16806,N_16719,N_16799);
xnor U16807 (N_16807,N_16780,N_16640);
xor U16808 (N_16808,N_16714,N_16794);
xnor U16809 (N_16809,N_16778,N_16661);
nor U16810 (N_16810,N_16689,N_16668);
nor U16811 (N_16811,N_16646,N_16641);
or U16812 (N_16812,N_16710,N_16713);
xnor U16813 (N_16813,N_16658,N_16696);
xnor U16814 (N_16814,N_16749,N_16747);
xnor U16815 (N_16815,N_16722,N_16734);
nor U16816 (N_16816,N_16723,N_16738);
and U16817 (N_16817,N_16771,N_16718);
nand U16818 (N_16818,N_16666,N_16781);
xor U16819 (N_16819,N_16774,N_16775);
or U16820 (N_16820,N_16770,N_16787);
and U16821 (N_16821,N_16758,N_16663);
or U16822 (N_16822,N_16692,N_16732);
or U16823 (N_16823,N_16691,N_16773);
nand U16824 (N_16824,N_16730,N_16702);
xor U16825 (N_16825,N_16674,N_16650);
and U16826 (N_16826,N_16755,N_16673);
or U16827 (N_16827,N_16642,N_16728);
and U16828 (N_16828,N_16785,N_16643);
nand U16829 (N_16829,N_16726,N_16733);
nand U16830 (N_16830,N_16687,N_16798);
xnor U16831 (N_16831,N_16660,N_16686);
or U16832 (N_16832,N_16754,N_16703);
xnor U16833 (N_16833,N_16792,N_16784);
nor U16834 (N_16834,N_16685,N_16740);
xnor U16835 (N_16835,N_16779,N_16670);
xnor U16836 (N_16836,N_16705,N_16682);
nand U16837 (N_16837,N_16757,N_16708);
xnor U16838 (N_16838,N_16671,N_16796);
nor U16839 (N_16839,N_16655,N_16777);
nand U16840 (N_16840,N_16743,N_16776);
nand U16841 (N_16841,N_16651,N_16786);
nand U16842 (N_16842,N_16647,N_16644);
and U16843 (N_16843,N_16649,N_16764);
nand U16844 (N_16844,N_16707,N_16791);
nor U16845 (N_16845,N_16720,N_16700);
and U16846 (N_16846,N_16763,N_16761);
xor U16847 (N_16847,N_16762,N_16657);
xor U16848 (N_16848,N_16676,N_16721);
xor U16849 (N_16849,N_16697,N_16767);
xnor U16850 (N_16850,N_16694,N_16790);
and U16851 (N_16851,N_16675,N_16716);
xor U16852 (N_16852,N_16797,N_16709);
nand U16853 (N_16853,N_16772,N_16706);
and U16854 (N_16854,N_16737,N_16698);
xor U16855 (N_16855,N_16736,N_16793);
xnor U16856 (N_16856,N_16677,N_16684);
xor U16857 (N_16857,N_16680,N_16750);
and U16858 (N_16858,N_16765,N_16693);
xnor U16859 (N_16859,N_16667,N_16679);
nand U16860 (N_16860,N_16656,N_16662);
xor U16861 (N_16861,N_16769,N_16768);
nand U16862 (N_16862,N_16664,N_16727);
or U16863 (N_16863,N_16724,N_16659);
or U16864 (N_16864,N_16745,N_16766);
nand U16865 (N_16865,N_16654,N_16715);
nand U16866 (N_16866,N_16681,N_16690);
xnor U16867 (N_16867,N_16782,N_16672);
nor U16868 (N_16868,N_16751,N_16753);
xor U16869 (N_16869,N_16756,N_16731);
nor U16870 (N_16870,N_16704,N_16699);
nand U16871 (N_16871,N_16688,N_16678);
nor U16872 (N_16872,N_16742,N_16653);
and U16873 (N_16873,N_16645,N_16788);
xnor U16874 (N_16874,N_16652,N_16741);
xor U16875 (N_16875,N_16735,N_16695);
xor U16876 (N_16876,N_16789,N_16752);
xor U16877 (N_16877,N_16748,N_16783);
or U16878 (N_16878,N_16746,N_16759);
nor U16879 (N_16879,N_16701,N_16711);
nor U16880 (N_16880,N_16665,N_16661);
xnor U16881 (N_16881,N_16700,N_16788);
nor U16882 (N_16882,N_16700,N_16675);
xnor U16883 (N_16883,N_16798,N_16726);
and U16884 (N_16884,N_16687,N_16666);
nor U16885 (N_16885,N_16734,N_16682);
and U16886 (N_16886,N_16726,N_16760);
nand U16887 (N_16887,N_16662,N_16758);
and U16888 (N_16888,N_16782,N_16773);
nor U16889 (N_16889,N_16685,N_16678);
nand U16890 (N_16890,N_16777,N_16748);
nand U16891 (N_16891,N_16737,N_16674);
nand U16892 (N_16892,N_16711,N_16747);
nand U16893 (N_16893,N_16740,N_16698);
or U16894 (N_16894,N_16668,N_16739);
nor U16895 (N_16895,N_16754,N_16663);
nor U16896 (N_16896,N_16786,N_16679);
and U16897 (N_16897,N_16776,N_16750);
nand U16898 (N_16898,N_16772,N_16671);
and U16899 (N_16899,N_16675,N_16685);
nand U16900 (N_16900,N_16748,N_16672);
nor U16901 (N_16901,N_16703,N_16676);
nand U16902 (N_16902,N_16654,N_16710);
and U16903 (N_16903,N_16751,N_16676);
nor U16904 (N_16904,N_16743,N_16688);
nor U16905 (N_16905,N_16719,N_16723);
nor U16906 (N_16906,N_16712,N_16681);
nand U16907 (N_16907,N_16790,N_16739);
nor U16908 (N_16908,N_16710,N_16762);
nand U16909 (N_16909,N_16650,N_16672);
xor U16910 (N_16910,N_16798,N_16792);
xnor U16911 (N_16911,N_16683,N_16659);
and U16912 (N_16912,N_16753,N_16752);
and U16913 (N_16913,N_16771,N_16773);
nand U16914 (N_16914,N_16702,N_16733);
xor U16915 (N_16915,N_16769,N_16794);
xor U16916 (N_16916,N_16799,N_16716);
and U16917 (N_16917,N_16772,N_16751);
nor U16918 (N_16918,N_16676,N_16643);
nor U16919 (N_16919,N_16744,N_16716);
xor U16920 (N_16920,N_16752,N_16736);
or U16921 (N_16921,N_16671,N_16699);
or U16922 (N_16922,N_16790,N_16753);
nand U16923 (N_16923,N_16787,N_16661);
or U16924 (N_16924,N_16738,N_16666);
nor U16925 (N_16925,N_16705,N_16673);
and U16926 (N_16926,N_16762,N_16769);
nand U16927 (N_16927,N_16692,N_16764);
xnor U16928 (N_16928,N_16740,N_16743);
or U16929 (N_16929,N_16740,N_16656);
or U16930 (N_16930,N_16756,N_16750);
nand U16931 (N_16931,N_16755,N_16789);
and U16932 (N_16932,N_16702,N_16653);
nand U16933 (N_16933,N_16757,N_16776);
xor U16934 (N_16934,N_16794,N_16772);
nor U16935 (N_16935,N_16698,N_16702);
xor U16936 (N_16936,N_16723,N_16696);
and U16937 (N_16937,N_16687,N_16656);
or U16938 (N_16938,N_16792,N_16729);
nand U16939 (N_16939,N_16694,N_16741);
xor U16940 (N_16940,N_16730,N_16796);
xnor U16941 (N_16941,N_16645,N_16770);
nor U16942 (N_16942,N_16720,N_16754);
xnor U16943 (N_16943,N_16671,N_16793);
or U16944 (N_16944,N_16697,N_16789);
nand U16945 (N_16945,N_16708,N_16703);
and U16946 (N_16946,N_16645,N_16674);
xor U16947 (N_16947,N_16761,N_16785);
xnor U16948 (N_16948,N_16670,N_16648);
nor U16949 (N_16949,N_16676,N_16718);
xor U16950 (N_16950,N_16725,N_16799);
or U16951 (N_16951,N_16772,N_16797);
nand U16952 (N_16952,N_16666,N_16712);
or U16953 (N_16953,N_16653,N_16654);
and U16954 (N_16954,N_16785,N_16799);
and U16955 (N_16955,N_16657,N_16688);
xnor U16956 (N_16956,N_16779,N_16690);
or U16957 (N_16957,N_16734,N_16779);
nor U16958 (N_16958,N_16794,N_16789);
and U16959 (N_16959,N_16677,N_16707);
nand U16960 (N_16960,N_16846,N_16896);
nand U16961 (N_16961,N_16932,N_16803);
nor U16962 (N_16962,N_16938,N_16847);
or U16963 (N_16963,N_16941,N_16910);
and U16964 (N_16964,N_16901,N_16810);
nor U16965 (N_16965,N_16857,N_16916);
xor U16966 (N_16966,N_16939,N_16887);
nand U16967 (N_16967,N_16940,N_16871);
or U16968 (N_16968,N_16894,N_16806);
nor U16969 (N_16969,N_16907,N_16861);
or U16970 (N_16970,N_16903,N_16917);
nand U16971 (N_16971,N_16825,N_16912);
nor U16972 (N_16972,N_16851,N_16947);
xor U16973 (N_16973,N_16948,N_16919);
nor U16974 (N_16974,N_16818,N_16937);
and U16975 (N_16975,N_16839,N_16942);
nor U16976 (N_16976,N_16884,N_16935);
nand U16977 (N_16977,N_16908,N_16951);
and U16978 (N_16978,N_16809,N_16930);
xor U16979 (N_16979,N_16911,N_16892);
nand U16980 (N_16980,N_16882,N_16831);
and U16981 (N_16981,N_16922,N_16843);
nor U16982 (N_16982,N_16842,N_16813);
nand U16983 (N_16983,N_16824,N_16891);
nor U16984 (N_16984,N_16817,N_16881);
xnor U16985 (N_16985,N_16864,N_16921);
nor U16986 (N_16986,N_16832,N_16838);
or U16987 (N_16987,N_16858,N_16927);
or U16988 (N_16988,N_16934,N_16954);
nor U16989 (N_16989,N_16853,N_16863);
nor U16990 (N_16990,N_16889,N_16821);
or U16991 (N_16991,N_16867,N_16957);
nand U16992 (N_16992,N_16950,N_16890);
nand U16993 (N_16993,N_16905,N_16829);
and U16994 (N_16994,N_16873,N_16840);
nor U16995 (N_16995,N_16893,N_16897);
nor U16996 (N_16996,N_16915,N_16936);
xor U16997 (N_16997,N_16944,N_16876);
nor U16998 (N_16998,N_16949,N_16906);
xor U16999 (N_16999,N_16868,N_16933);
nand U17000 (N_17000,N_16928,N_16860);
nand U17001 (N_17001,N_16914,N_16913);
nand U17002 (N_17002,N_16946,N_16837);
nor U17003 (N_17003,N_16826,N_16902);
nand U17004 (N_17004,N_16835,N_16811);
and U17005 (N_17005,N_16856,N_16878);
or U17006 (N_17006,N_16959,N_16812);
nor U17007 (N_17007,N_16879,N_16807);
and U17008 (N_17008,N_16816,N_16926);
and U17009 (N_17009,N_16952,N_16841);
and U17010 (N_17010,N_16855,N_16943);
or U17011 (N_17011,N_16850,N_16909);
xnor U17012 (N_17012,N_16869,N_16866);
xnor U17013 (N_17013,N_16845,N_16804);
xor U17014 (N_17014,N_16859,N_16814);
nand U17015 (N_17015,N_16828,N_16888);
and U17016 (N_17016,N_16834,N_16865);
xnor U17017 (N_17017,N_16899,N_16872);
nand U17018 (N_17018,N_16875,N_16808);
or U17019 (N_17019,N_16827,N_16819);
nor U17020 (N_17020,N_16898,N_16802);
or U17021 (N_17021,N_16931,N_16823);
nor U17022 (N_17022,N_16870,N_16958);
and U17023 (N_17023,N_16929,N_16805);
or U17024 (N_17024,N_16925,N_16848);
or U17025 (N_17025,N_16815,N_16874);
xnor U17026 (N_17026,N_16854,N_16945);
and U17027 (N_17027,N_16955,N_16895);
and U17028 (N_17028,N_16920,N_16836);
nor U17029 (N_17029,N_16833,N_16924);
or U17030 (N_17030,N_16923,N_16886);
nand U17031 (N_17031,N_16849,N_16830);
xnor U17032 (N_17032,N_16801,N_16877);
nor U17033 (N_17033,N_16800,N_16885);
nand U17034 (N_17034,N_16862,N_16822);
nor U17035 (N_17035,N_16844,N_16904);
and U17036 (N_17036,N_16900,N_16883);
nor U17037 (N_17037,N_16956,N_16820);
and U17038 (N_17038,N_16953,N_16918);
nand U17039 (N_17039,N_16852,N_16880);
xnor U17040 (N_17040,N_16806,N_16906);
nand U17041 (N_17041,N_16899,N_16853);
and U17042 (N_17042,N_16834,N_16924);
nor U17043 (N_17043,N_16941,N_16857);
nand U17044 (N_17044,N_16815,N_16832);
or U17045 (N_17045,N_16897,N_16832);
nor U17046 (N_17046,N_16830,N_16935);
nor U17047 (N_17047,N_16953,N_16894);
nor U17048 (N_17048,N_16942,N_16909);
xnor U17049 (N_17049,N_16930,N_16917);
nand U17050 (N_17050,N_16809,N_16895);
nor U17051 (N_17051,N_16829,N_16941);
or U17052 (N_17052,N_16856,N_16892);
and U17053 (N_17053,N_16939,N_16894);
nor U17054 (N_17054,N_16821,N_16828);
and U17055 (N_17055,N_16933,N_16903);
xor U17056 (N_17056,N_16836,N_16953);
nand U17057 (N_17057,N_16934,N_16847);
xor U17058 (N_17058,N_16942,N_16841);
nand U17059 (N_17059,N_16831,N_16927);
and U17060 (N_17060,N_16910,N_16950);
nand U17061 (N_17061,N_16816,N_16807);
xnor U17062 (N_17062,N_16821,N_16835);
or U17063 (N_17063,N_16825,N_16803);
nor U17064 (N_17064,N_16836,N_16861);
nor U17065 (N_17065,N_16869,N_16859);
nand U17066 (N_17066,N_16957,N_16918);
nand U17067 (N_17067,N_16929,N_16928);
and U17068 (N_17068,N_16810,N_16812);
nand U17069 (N_17069,N_16944,N_16836);
nor U17070 (N_17070,N_16911,N_16882);
nor U17071 (N_17071,N_16913,N_16816);
xnor U17072 (N_17072,N_16942,N_16834);
nor U17073 (N_17073,N_16856,N_16819);
nor U17074 (N_17074,N_16908,N_16909);
nor U17075 (N_17075,N_16819,N_16829);
nand U17076 (N_17076,N_16810,N_16806);
nand U17077 (N_17077,N_16846,N_16909);
nand U17078 (N_17078,N_16845,N_16802);
and U17079 (N_17079,N_16950,N_16818);
and U17080 (N_17080,N_16844,N_16819);
xor U17081 (N_17081,N_16941,N_16851);
nor U17082 (N_17082,N_16931,N_16946);
and U17083 (N_17083,N_16857,N_16886);
and U17084 (N_17084,N_16821,N_16868);
nand U17085 (N_17085,N_16956,N_16827);
or U17086 (N_17086,N_16921,N_16836);
nand U17087 (N_17087,N_16818,N_16916);
and U17088 (N_17088,N_16934,N_16815);
xnor U17089 (N_17089,N_16806,N_16936);
nand U17090 (N_17090,N_16926,N_16879);
or U17091 (N_17091,N_16901,N_16905);
or U17092 (N_17092,N_16944,N_16805);
and U17093 (N_17093,N_16907,N_16912);
or U17094 (N_17094,N_16852,N_16938);
or U17095 (N_17095,N_16877,N_16931);
nor U17096 (N_17096,N_16903,N_16949);
nand U17097 (N_17097,N_16836,N_16844);
xor U17098 (N_17098,N_16869,N_16940);
nor U17099 (N_17099,N_16856,N_16934);
xnor U17100 (N_17100,N_16939,N_16892);
or U17101 (N_17101,N_16913,N_16836);
xor U17102 (N_17102,N_16932,N_16947);
or U17103 (N_17103,N_16947,N_16890);
and U17104 (N_17104,N_16955,N_16822);
xnor U17105 (N_17105,N_16840,N_16846);
xnor U17106 (N_17106,N_16882,N_16839);
nand U17107 (N_17107,N_16914,N_16812);
nand U17108 (N_17108,N_16890,N_16908);
nor U17109 (N_17109,N_16951,N_16842);
and U17110 (N_17110,N_16894,N_16896);
and U17111 (N_17111,N_16927,N_16892);
nand U17112 (N_17112,N_16833,N_16896);
or U17113 (N_17113,N_16925,N_16808);
nor U17114 (N_17114,N_16837,N_16855);
or U17115 (N_17115,N_16847,N_16820);
and U17116 (N_17116,N_16811,N_16954);
nand U17117 (N_17117,N_16841,N_16868);
nand U17118 (N_17118,N_16931,N_16924);
nor U17119 (N_17119,N_16877,N_16908);
nand U17120 (N_17120,N_16975,N_17094);
xnor U17121 (N_17121,N_16967,N_17069);
and U17122 (N_17122,N_17104,N_17034);
or U17123 (N_17123,N_17042,N_16965);
nor U17124 (N_17124,N_17080,N_16971);
xnor U17125 (N_17125,N_17103,N_17052);
and U17126 (N_17126,N_17028,N_16979);
and U17127 (N_17127,N_17062,N_17043);
xor U17128 (N_17128,N_17089,N_17008);
nand U17129 (N_17129,N_17078,N_17115);
and U17130 (N_17130,N_16999,N_16977);
xor U17131 (N_17131,N_17102,N_16969);
or U17132 (N_17132,N_17095,N_17090);
or U17133 (N_17133,N_17013,N_17076);
nor U17134 (N_17134,N_16982,N_17077);
nand U17135 (N_17135,N_17117,N_17074);
nand U17136 (N_17136,N_17079,N_17018);
nor U17137 (N_17137,N_16980,N_16978);
xnor U17138 (N_17138,N_17075,N_16976);
or U17139 (N_17139,N_16998,N_17057);
or U17140 (N_17140,N_17005,N_17110);
or U17141 (N_17141,N_17007,N_17070);
and U17142 (N_17142,N_16996,N_17055);
and U17143 (N_17143,N_16960,N_16968);
xnor U17144 (N_17144,N_17032,N_17119);
nand U17145 (N_17145,N_17003,N_16985);
nor U17146 (N_17146,N_17108,N_17024);
xnor U17147 (N_17147,N_17009,N_17025);
xor U17148 (N_17148,N_17100,N_17066);
nor U17149 (N_17149,N_16981,N_16984);
xnor U17150 (N_17150,N_17012,N_17002);
nor U17151 (N_17151,N_17093,N_17099);
nand U17152 (N_17152,N_17016,N_17097);
nand U17153 (N_17153,N_16991,N_17082);
nor U17154 (N_17154,N_17050,N_17045);
nand U17155 (N_17155,N_16997,N_17054);
or U17156 (N_17156,N_17088,N_17059);
nand U17157 (N_17157,N_16986,N_17058);
nand U17158 (N_17158,N_17114,N_16983);
nor U17159 (N_17159,N_16992,N_17063);
nand U17160 (N_17160,N_17116,N_17021);
and U17161 (N_17161,N_17048,N_17109);
and U17162 (N_17162,N_17085,N_17030);
nand U17163 (N_17163,N_17001,N_16963);
and U17164 (N_17164,N_17112,N_17113);
nor U17165 (N_17165,N_16964,N_17049);
xor U17166 (N_17166,N_17118,N_17060);
or U17167 (N_17167,N_17111,N_16974);
nor U17168 (N_17168,N_16973,N_17064);
and U17169 (N_17169,N_17096,N_16989);
xor U17170 (N_17170,N_17026,N_17040);
xor U17171 (N_17171,N_17038,N_17047);
nor U17172 (N_17172,N_17061,N_17065);
nor U17173 (N_17173,N_16961,N_17083);
xnor U17174 (N_17174,N_17036,N_17084);
and U17175 (N_17175,N_17041,N_17027);
xor U17176 (N_17176,N_17046,N_17006);
nor U17177 (N_17177,N_16972,N_17073);
nand U17178 (N_17178,N_17051,N_16988);
or U17179 (N_17179,N_16966,N_17014);
nor U17180 (N_17180,N_17044,N_17000);
or U17181 (N_17181,N_17011,N_17010);
or U17182 (N_17182,N_17031,N_17022);
nand U17183 (N_17183,N_16995,N_16970);
and U17184 (N_17184,N_16962,N_17081);
nor U17185 (N_17185,N_17086,N_17004);
nand U17186 (N_17186,N_17098,N_17019);
or U17187 (N_17187,N_16990,N_17092);
or U17188 (N_17188,N_16993,N_17056);
or U17189 (N_17189,N_17017,N_17072);
and U17190 (N_17190,N_17106,N_17101);
nor U17191 (N_17191,N_17037,N_16987);
nand U17192 (N_17192,N_17023,N_17020);
nand U17193 (N_17193,N_17035,N_17039);
nor U17194 (N_17194,N_17087,N_17053);
and U17195 (N_17195,N_17067,N_17105);
or U17196 (N_17196,N_17071,N_17068);
nand U17197 (N_17197,N_17033,N_17091);
or U17198 (N_17198,N_17029,N_16994);
or U17199 (N_17199,N_17107,N_17015);
nor U17200 (N_17200,N_17087,N_16988);
nor U17201 (N_17201,N_16979,N_16968);
xnor U17202 (N_17202,N_16974,N_17014);
nand U17203 (N_17203,N_16976,N_17021);
nand U17204 (N_17204,N_17097,N_17107);
nor U17205 (N_17205,N_17002,N_17113);
xnor U17206 (N_17206,N_16960,N_17043);
or U17207 (N_17207,N_17043,N_16998);
or U17208 (N_17208,N_17078,N_17044);
and U17209 (N_17209,N_17053,N_16985);
nor U17210 (N_17210,N_17117,N_17111);
or U17211 (N_17211,N_17068,N_17075);
nand U17212 (N_17212,N_17053,N_17027);
xor U17213 (N_17213,N_17027,N_17044);
nor U17214 (N_17214,N_17097,N_17020);
xnor U17215 (N_17215,N_16978,N_16964);
and U17216 (N_17216,N_17101,N_17032);
or U17217 (N_17217,N_17068,N_16991);
xnor U17218 (N_17218,N_17113,N_16972);
and U17219 (N_17219,N_17031,N_17089);
nand U17220 (N_17220,N_17110,N_17048);
nor U17221 (N_17221,N_17042,N_17044);
or U17222 (N_17222,N_17002,N_17000);
nand U17223 (N_17223,N_17062,N_17030);
nand U17224 (N_17224,N_17006,N_17095);
and U17225 (N_17225,N_16972,N_16986);
nor U17226 (N_17226,N_16991,N_17030);
xor U17227 (N_17227,N_17084,N_16978);
xor U17228 (N_17228,N_17026,N_17082);
nand U17229 (N_17229,N_17042,N_17007);
or U17230 (N_17230,N_16983,N_17074);
nor U17231 (N_17231,N_17030,N_17033);
or U17232 (N_17232,N_16999,N_17044);
or U17233 (N_17233,N_17038,N_17081);
nor U17234 (N_17234,N_17025,N_17082);
nor U17235 (N_17235,N_16993,N_16969);
nor U17236 (N_17236,N_16994,N_17103);
or U17237 (N_17237,N_17073,N_17086);
nor U17238 (N_17238,N_17034,N_17047);
or U17239 (N_17239,N_17106,N_17111);
or U17240 (N_17240,N_16971,N_17093);
nor U17241 (N_17241,N_17087,N_16992);
xor U17242 (N_17242,N_16984,N_16978);
nand U17243 (N_17243,N_16969,N_17092);
nand U17244 (N_17244,N_17086,N_17068);
or U17245 (N_17245,N_17014,N_17065);
and U17246 (N_17246,N_17112,N_17085);
xor U17247 (N_17247,N_17068,N_17074);
and U17248 (N_17248,N_17102,N_17001);
xor U17249 (N_17249,N_17074,N_17049);
nor U17250 (N_17250,N_17067,N_17057);
or U17251 (N_17251,N_17051,N_17106);
or U17252 (N_17252,N_17116,N_17011);
and U17253 (N_17253,N_17040,N_17074);
and U17254 (N_17254,N_17021,N_16998);
xor U17255 (N_17255,N_16963,N_17069);
nand U17256 (N_17256,N_17011,N_17007);
nor U17257 (N_17257,N_17070,N_17097);
nor U17258 (N_17258,N_17004,N_16960);
or U17259 (N_17259,N_17066,N_16989);
and U17260 (N_17260,N_17050,N_17069);
nand U17261 (N_17261,N_17067,N_16963);
and U17262 (N_17262,N_17067,N_17118);
xnor U17263 (N_17263,N_16993,N_17023);
and U17264 (N_17264,N_17078,N_17028);
nor U17265 (N_17265,N_16966,N_17025);
xor U17266 (N_17266,N_17115,N_16998);
or U17267 (N_17267,N_17051,N_16965);
nand U17268 (N_17268,N_17116,N_17109);
xor U17269 (N_17269,N_17065,N_17005);
and U17270 (N_17270,N_16985,N_17051);
nor U17271 (N_17271,N_17103,N_17090);
or U17272 (N_17272,N_16987,N_17027);
nor U17273 (N_17273,N_16968,N_17024);
nand U17274 (N_17274,N_17106,N_16971);
nand U17275 (N_17275,N_17040,N_17111);
or U17276 (N_17276,N_17058,N_17014);
nor U17277 (N_17277,N_17060,N_17004);
nor U17278 (N_17278,N_17069,N_17014);
xor U17279 (N_17279,N_17080,N_17030);
or U17280 (N_17280,N_17190,N_17161);
nand U17281 (N_17281,N_17150,N_17247);
or U17282 (N_17282,N_17259,N_17145);
and U17283 (N_17283,N_17122,N_17123);
nand U17284 (N_17284,N_17176,N_17239);
or U17285 (N_17285,N_17128,N_17152);
nor U17286 (N_17286,N_17199,N_17255);
nand U17287 (N_17287,N_17157,N_17265);
xnor U17288 (N_17288,N_17207,N_17245);
and U17289 (N_17289,N_17276,N_17253);
or U17290 (N_17290,N_17221,N_17121);
nand U17291 (N_17291,N_17154,N_17146);
nand U17292 (N_17292,N_17162,N_17164);
and U17293 (N_17293,N_17225,N_17129);
nand U17294 (N_17294,N_17256,N_17249);
xnor U17295 (N_17295,N_17126,N_17254);
and U17296 (N_17296,N_17186,N_17266);
and U17297 (N_17297,N_17187,N_17242);
or U17298 (N_17298,N_17173,N_17148);
nor U17299 (N_17299,N_17144,N_17258);
and U17300 (N_17300,N_17216,N_17274);
nand U17301 (N_17301,N_17264,N_17278);
and U17302 (N_17302,N_17175,N_17184);
nor U17303 (N_17303,N_17268,N_17211);
xor U17304 (N_17304,N_17200,N_17260);
nand U17305 (N_17305,N_17214,N_17237);
or U17306 (N_17306,N_17140,N_17203);
xor U17307 (N_17307,N_17205,N_17262);
xnor U17308 (N_17308,N_17182,N_17141);
nand U17309 (N_17309,N_17269,N_17217);
and U17310 (N_17310,N_17236,N_17235);
or U17311 (N_17311,N_17153,N_17189);
nand U17312 (N_17312,N_17196,N_17215);
nand U17313 (N_17313,N_17230,N_17130);
nor U17314 (N_17314,N_17257,N_17136);
or U17315 (N_17315,N_17261,N_17272);
nand U17316 (N_17316,N_17166,N_17243);
and U17317 (N_17317,N_17171,N_17227);
or U17318 (N_17318,N_17270,N_17159);
nand U17319 (N_17319,N_17202,N_17142);
nand U17320 (N_17320,N_17228,N_17151);
or U17321 (N_17321,N_17251,N_17180);
or U17322 (N_17322,N_17223,N_17206);
nor U17323 (N_17323,N_17198,N_17279);
nor U17324 (N_17324,N_17127,N_17133);
nor U17325 (N_17325,N_17135,N_17213);
nand U17326 (N_17326,N_17234,N_17191);
and U17327 (N_17327,N_17158,N_17188);
xor U17328 (N_17328,N_17275,N_17143);
xnor U17329 (N_17329,N_17149,N_17156);
xor U17330 (N_17330,N_17193,N_17177);
and U17331 (N_17331,N_17208,N_17124);
xnor U17332 (N_17332,N_17267,N_17218);
nand U17333 (N_17333,N_17163,N_17168);
or U17334 (N_17334,N_17155,N_17192);
and U17335 (N_17335,N_17212,N_17185);
xnor U17336 (N_17336,N_17160,N_17226);
nand U17337 (N_17337,N_17195,N_17277);
nor U17338 (N_17338,N_17222,N_17170);
xnor U17339 (N_17339,N_17137,N_17139);
nand U17340 (N_17340,N_17120,N_17201);
nor U17341 (N_17341,N_17250,N_17194);
and U17342 (N_17342,N_17131,N_17238);
xor U17343 (N_17343,N_17167,N_17132);
and U17344 (N_17344,N_17183,N_17241);
and U17345 (N_17345,N_17219,N_17233);
or U17346 (N_17346,N_17263,N_17220);
xor U17347 (N_17347,N_17240,N_17248);
or U17348 (N_17348,N_17178,N_17273);
or U17349 (N_17349,N_17165,N_17179);
nor U17350 (N_17350,N_17174,N_17197);
or U17351 (N_17351,N_17231,N_17232);
xnor U17352 (N_17352,N_17147,N_17210);
and U17353 (N_17353,N_17246,N_17134);
nor U17354 (N_17354,N_17125,N_17172);
or U17355 (N_17355,N_17169,N_17252);
or U17356 (N_17356,N_17181,N_17271);
and U17357 (N_17357,N_17224,N_17229);
nand U17358 (N_17358,N_17138,N_17244);
or U17359 (N_17359,N_17204,N_17209);
or U17360 (N_17360,N_17181,N_17273);
nor U17361 (N_17361,N_17195,N_17256);
xnor U17362 (N_17362,N_17267,N_17254);
nor U17363 (N_17363,N_17192,N_17166);
or U17364 (N_17364,N_17276,N_17237);
xor U17365 (N_17365,N_17246,N_17131);
or U17366 (N_17366,N_17127,N_17178);
xnor U17367 (N_17367,N_17209,N_17203);
and U17368 (N_17368,N_17219,N_17165);
xor U17369 (N_17369,N_17234,N_17249);
or U17370 (N_17370,N_17130,N_17164);
and U17371 (N_17371,N_17240,N_17143);
and U17372 (N_17372,N_17251,N_17148);
or U17373 (N_17373,N_17210,N_17187);
xnor U17374 (N_17374,N_17155,N_17169);
nor U17375 (N_17375,N_17147,N_17227);
xnor U17376 (N_17376,N_17279,N_17162);
or U17377 (N_17377,N_17161,N_17162);
and U17378 (N_17378,N_17209,N_17145);
or U17379 (N_17379,N_17141,N_17191);
or U17380 (N_17380,N_17126,N_17139);
or U17381 (N_17381,N_17217,N_17138);
or U17382 (N_17382,N_17197,N_17252);
xnor U17383 (N_17383,N_17157,N_17196);
xnor U17384 (N_17384,N_17177,N_17203);
nand U17385 (N_17385,N_17265,N_17151);
and U17386 (N_17386,N_17161,N_17278);
or U17387 (N_17387,N_17194,N_17142);
or U17388 (N_17388,N_17224,N_17157);
nand U17389 (N_17389,N_17184,N_17176);
nand U17390 (N_17390,N_17271,N_17252);
or U17391 (N_17391,N_17133,N_17199);
and U17392 (N_17392,N_17176,N_17214);
or U17393 (N_17393,N_17250,N_17144);
nand U17394 (N_17394,N_17221,N_17197);
and U17395 (N_17395,N_17178,N_17203);
nor U17396 (N_17396,N_17203,N_17157);
xnor U17397 (N_17397,N_17161,N_17246);
xnor U17398 (N_17398,N_17219,N_17238);
xor U17399 (N_17399,N_17162,N_17247);
and U17400 (N_17400,N_17198,N_17169);
nor U17401 (N_17401,N_17261,N_17230);
xor U17402 (N_17402,N_17134,N_17130);
or U17403 (N_17403,N_17247,N_17165);
xnor U17404 (N_17404,N_17243,N_17210);
nor U17405 (N_17405,N_17237,N_17178);
xnor U17406 (N_17406,N_17258,N_17263);
nor U17407 (N_17407,N_17127,N_17275);
and U17408 (N_17408,N_17243,N_17242);
nor U17409 (N_17409,N_17137,N_17213);
or U17410 (N_17410,N_17178,N_17139);
or U17411 (N_17411,N_17141,N_17271);
or U17412 (N_17412,N_17180,N_17128);
nor U17413 (N_17413,N_17246,N_17127);
nor U17414 (N_17414,N_17133,N_17220);
nor U17415 (N_17415,N_17189,N_17210);
or U17416 (N_17416,N_17247,N_17253);
nand U17417 (N_17417,N_17204,N_17137);
and U17418 (N_17418,N_17274,N_17239);
xnor U17419 (N_17419,N_17250,N_17254);
nor U17420 (N_17420,N_17183,N_17252);
or U17421 (N_17421,N_17232,N_17137);
or U17422 (N_17422,N_17223,N_17134);
nor U17423 (N_17423,N_17143,N_17144);
nor U17424 (N_17424,N_17207,N_17180);
xnor U17425 (N_17425,N_17255,N_17196);
or U17426 (N_17426,N_17174,N_17161);
nor U17427 (N_17427,N_17141,N_17163);
nor U17428 (N_17428,N_17142,N_17275);
or U17429 (N_17429,N_17250,N_17175);
nand U17430 (N_17430,N_17153,N_17165);
and U17431 (N_17431,N_17215,N_17122);
nand U17432 (N_17432,N_17152,N_17241);
xnor U17433 (N_17433,N_17233,N_17144);
or U17434 (N_17434,N_17221,N_17213);
and U17435 (N_17435,N_17196,N_17179);
or U17436 (N_17436,N_17134,N_17244);
nor U17437 (N_17437,N_17249,N_17151);
nor U17438 (N_17438,N_17137,N_17135);
nor U17439 (N_17439,N_17141,N_17244);
xor U17440 (N_17440,N_17401,N_17427);
and U17441 (N_17441,N_17308,N_17322);
or U17442 (N_17442,N_17354,N_17352);
nor U17443 (N_17443,N_17303,N_17312);
xnor U17444 (N_17444,N_17386,N_17346);
nor U17445 (N_17445,N_17324,N_17399);
and U17446 (N_17446,N_17385,N_17311);
and U17447 (N_17447,N_17335,N_17376);
xnor U17448 (N_17448,N_17280,N_17300);
and U17449 (N_17449,N_17287,N_17415);
or U17450 (N_17450,N_17368,N_17298);
xnor U17451 (N_17451,N_17296,N_17323);
and U17452 (N_17452,N_17294,N_17379);
xnor U17453 (N_17453,N_17337,N_17383);
xnor U17454 (N_17454,N_17360,N_17364);
or U17455 (N_17455,N_17299,N_17336);
or U17456 (N_17456,N_17367,N_17378);
nor U17457 (N_17457,N_17351,N_17405);
or U17458 (N_17458,N_17409,N_17431);
or U17459 (N_17459,N_17374,N_17421);
or U17460 (N_17460,N_17332,N_17377);
xnor U17461 (N_17461,N_17398,N_17411);
xnor U17462 (N_17462,N_17406,N_17284);
nand U17463 (N_17463,N_17315,N_17345);
xor U17464 (N_17464,N_17326,N_17305);
nand U17465 (N_17465,N_17433,N_17373);
nor U17466 (N_17466,N_17396,N_17432);
and U17467 (N_17467,N_17316,N_17321);
and U17468 (N_17468,N_17435,N_17416);
nand U17469 (N_17469,N_17304,N_17290);
and U17470 (N_17470,N_17343,N_17387);
and U17471 (N_17471,N_17403,N_17397);
or U17472 (N_17472,N_17342,N_17414);
or U17473 (N_17473,N_17293,N_17281);
and U17474 (N_17474,N_17286,N_17333);
nor U17475 (N_17475,N_17412,N_17301);
or U17476 (N_17476,N_17372,N_17417);
or U17477 (N_17477,N_17370,N_17282);
and U17478 (N_17478,N_17307,N_17359);
nor U17479 (N_17479,N_17283,N_17389);
and U17480 (N_17480,N_17390,N_17327);
and U17481 (N_17481,N_17329,N_17349);
nor U17482 (N_17482,N_17292,N_17402);
and U17483 (N_17483,N_17340,N_17388);
or U17484 (N_17484,N_17381,N_17436);
or U17485 (N_17485,N_17353,N_17361);
and U17486 (N_17486,N_17437,N_17426);
nor U17487 (N_17487,N_17438,N_17369);
and U17488 (N_17488,N_17356,N_17289);
xor U17489 (N_17489,N_17423,N_17428);
or U17490 (N_17490,N_17334,N_17310);
or U17491 (N_17491,N_17341,N_17391);
and U17492 (N_17492,N_17288,N_17328);
nor U17493 (N_17493,N_17400,N_17347);
nand U17494 (N_17494,N_17338,N_17420);
nand U17495 (N_17495,N_17410,N_17358);
nor U17496 (N_17496,N_17407,N_17320);
nand U17497 (N_17497,N_17422,N_17291);
and U17498 (N_17498,N_17309,N_17371);
and U17499 (N_17499,N_17380,N_17319);
nor U17500 (N_17500,N_17419,N_17429);
or U17501 (N_17501,N_17418,N_17393);
or U17502 (N_17502,N_17394,N_17325);
or U17503 (N_17503,N_17285,N_17297);
xnor U17504 (N_17504,N_17365,N_17413);
nand U17505 (N_17505,N_17350,N_17384);
xor U17506 (N_17506,N_17439,N_17317);
nand U17507 (N_17507,N_17408,N_17430);
nand U17508 (N_17508,N_17355,N_17318);
or U17509 (N_17509,N_17392,N_17366);
and U17510 (N_17510,N_17348,N_17395);
nor U17511 (N_17511,N_17295,N_17375);
and U17512 (N_17512,N_17314,N_17357);
nand U17513 (N_17513,N_17306,N_17313);
xor U17514 (N_17514,N_17331,N_17424);
or U17515 (N_17515,N_17404,N_17363);
or U17516 (N_17516,N_17434,N_17330);
or U17517 (N_17517,N_17425,N_17382);
and U17518 (N_17518,N_17339,N_17362);
and U17519 (N_17519,N_17302,N_17344);
nand U17520 (N_17520,N_17394,N_17354);
nor U17521 (N_17521,N_17386,N_17331);
or U17522 (N_17522,N_17409,N_17307);
nor U17523 (N_17523,N_17376,N_17361);
and U17524 (N_17524,N_17364,N_17283);
xnor U17525 (N_17525,N_17408,N_17333);
or U17526 (N_17526,N_17303,N_17434);
nand U17527 (N_17527,N_17411,N_17385);
and U17528 (N_17528,N_17284,N_17301);
nor U17529 (N_17529,N_17320,N_17404);
and U17530 (N_17530,N_17390,N_17299);
xnor U17531 (N_17531,N_17297,N_17366);
nor U17532 (N_17532,N_17436,N_17405);
and U17533 (N_17533,N_17409,N_17281);
nand U17534 (N_17534,N_17393,N_17317);
or U17535 (N_17535,N_17423,N_17396);
nor U17536 (N_17536,N_17382,N_17365);
nor U17537 (N_17537,N_17414,N_17367);
and U17538 (N_17538,N_17286,N_17422);
or U17539 (N_17539,N_17371,N_17416);
and U17540 (N_17540,N_17427,N_17429);
nand U17541 (N_17541,N_17314,N_17419);
and U17542 (N_17542,N_17431,N_17371);
xnor U17543 (N_17543,N_17400,N_17418);
or U17544 (N_17544,N_17283,N_17288);
or U17545 (N_17545,N_17347,N_17361);
and U17546 (N_17546,N_17342,N_17353);
or U17547 (N_17547,N_17438,N_17314);
or U17548 (N_17548,N_17350,N_17424);
and U17549 (N_17549,N_17326,N_17422);
nor U17550 (N_17550,N_17329,N_17285);
nand U17551 (N_17551,N_17423,N_17302);
nand U17552 (N_17552,N_17310,N_17381);
and U17553 (N_17553,N_17309,N_17423);
or U17554 (N_17554,N_17358,N_17392);
nor U17555 (N_17555,N_17368,N_17411);
nor U17556 (N_17556,N_17431,N_17407);
nor U17557 (N_17557,N_17329,N_17370);
nand U17558 (N_17558,N_17323,N_17427);
nor U17559 (N_17559,N_17326,N_17430);
or U17560 (N_17560,N_17297,N_17298);
and U17561 (N_17561,N_17352,N_17342);
nor U17562 (N_17562,N_17328,N_17401);
nand U17563 (N_17563,N_17306,N_17410);
and U17564 (N_17564,N_17308,N_17286);
and U17565 (N_17565,N_17358,N_17426);
nor U17566 (N_17566,N_17336,N_17285);
xor U17567 (N_17567,N_17299,N_17420);
nand U17568 (N_17568,N_17349,N_17309);
or U17569 (N_17569,N_17352,N_17309);
xnor U17570 (N_17570,N_17361,N_17332);
nand U17571 (N_17571,N_17438,N_17296);
or U17572 (N_17572,N_17361,N_17315);
nor U17573 (N_17573,N_17339,N_17288);
and U17574 (N_17574,N_17358,N_17437);
or U17575 (N_17575,N_17377,N_17401);
or U17576 (N_17576,N_17436,N_17357);
xor U17577 (N_17577,N_17387,N_17328);
nand U17578 (N_17578,N_17311,N_17356);
nand U17579 (N_17579,N_17409,N_17315);
xnor U17580 (N_17580,N_17295,N_17314);
nand U17581 (N_17581,N_17403,N_17284);
xnor U17582 (N_17582,N_17343,N_17318);
nand U17583 (N_17583,N_17349,N_17396);
nor U17584 (N_17584,N_17369,N_17346);
or U17585 (N_17585,N_17425,N_17401);
xnor U17586 (N_17586,N_17378,N_17386);
or U17587 (N_17587,N_17424,N_17403);
and U17588 (N_17588,N_17359,N_17289);
xor U17589 (N_17589,N_17331,N_17316);
or U17590 (N_17590,N_17345,N_17316);
nor U17591 (N_17591,N_17384,N_17352);
nor U17592 (N_17592,N_17327,N_17430);
nor U17593 (N_17593,N_17337,N_17394);
xor U17594 (N_17594,N_17382,N_17407);
nor U17595 (N_17595,N_17435,N_17388);
xor U17596 (N_17596,N_17387,N_17411);
nor U17597 (N_17597,N_17346,N_17358);
nand U17598 (N_17598,N_17298,N_17296);
or U17599 (N_17599,N_17401,N_17306);
or U17600 (N_17600,N_17465,N_17587);
nand U17601 (N_17601,N_17535,N_17454);
xor U17602 (N_17602,N_17488,N_17524);
and U17603 (N_17603,N_17474,N_17507);
nand U17604 (N_17604,N_17493,N_17492);
or U17605 (N_17605,N_17545,N_17468);
xnor U17606 (N_17606,N_17484,N_17574);
nor U17607 (N_17607,N_17518,N_17511);
nand U17608 (N_17608,N_17483,N_17499);
nand U17609 (N_17609,N_17544,N_17531);
or U17610 (N_17610,N_17455,N_17522);
and U17611 (N_17611,N_17478,N_17526);
nor U17612 (N_17612,N_17443,N_17501);
nand U17613 (N_17613,N_17538,N_17489);
xor U17614 (N_17614,N_17473,N_17503);
or U17615 (N_17615,N_17521,N_17576);
nor U17616 (N_17616,N_17547,N_17461);
or U17617 (N_17617,N_17516,N_17475);
nor U17618 (N_17618,N_17519,N_17569);
or U17619 (N_17619,N_17497,N_17546);
xnor U17620 (N_17620,N_17567,N_17456);
or U17621 (N_17621,N_17581,N_17565);
or U17622 (N_17622,N_17450,N_17557);
nand U17623 (N_17623,N_17570,N_17527);
or U17624 (N_17624,N_17543,N_17495);
xnor U17625 (N_17625,N_17537,N_17481);
nor U17626 (N_17626,N_17528,N_17476);
and U17627 (N_17627,N_17529,N_17471);
or U17628 (N_17628,N_17560,N_17575);
nand U17629 (N_17629,N_17512,N_17515);
xnor U17630 (N_17630,N_17551,N_17448);
or U17631 (N_17631,N_17564,N_17589);
and U17632 (N_17632,N_17447,N_17556);
nand U17633 (N_17633,N_17485,N_17494);
nand U17634 (N_17634,N_17568,N_17451);
and U17635 (N_17635,N_17580,N_17444);
nand U17636 (N_17636,N_17458,N_17533);
and U17637 (N_17637,N_17536,N_17571);
or U17638 (N_17638,N_17463,N_17597);
nor U17639 (N_17639,N_17464,N_17477);
nor U17640 (N_17640,N_17504,N_17586);
nand U17641 (N_17641,N_17466,N_17442);
xnor U17642 (N_17642,N_17594,N_17452);
nand U17643 (N_17643,N_17561,N_17534);
and U17644 (N_17644,N_17498,N_17505);
nor U17645 (N_17645,N_17530,N_17539);
xnor U17646 (N_17646,N_17592,N_17541);
nor U17647 (N_17647,N_17514,N_17479);
or U17648 (N_17648,N_17508,N_17578);
and U17649 (N_17649,N_17513,N_17453);
and U17650 (N_17650,N_17462,N_17579);
nand U17651 (N_17651,N_17566,N_17506);
or U17652 (N_17652,N_17460,N_17532);
nor U17653 (N_17653,N_17523,N_17525);
nor U17654 (N_17654,N_17596,N_17585);
nand U17655 (N_17655,N_17549,N_17590);
nor U17656 (N_17656,N_17520,N_17552);
or U17657 (N_17657,N_17555,N_17490);
xor U17658 (N_17658,N_17588,N_17553);
and U17659 (N_17659,N_17496,N_17467);
nand U17660 (N_17660,N_17583,N_17449);
nand U17661 (N_17661,N_17480,N_17558);
and U17662 (N_17662,N_17470,N_17469);
or U17663 (N_17663,N_17459,N_17598);
xnor U17664 (N_17664,N_17593,N_17595);
xnor U17665 (N_17665,N_17502,N_17542);
and U17666 (N_17666,N_17487,N_17491);
nor U17667 (N_17667,N_17573,N_17550);
nand U17668 (N_17668,N_17559,N_17540);
and U17669 (N_17669,N_17500,N_17599);
nand U17670 (N_17670,N_17582,N_17584);
nor U17671 (N_17671,N_17554,N_17440);
xnor U17672 (N_17672,N_17441,N_17562);
nand U17673 (N_17673,N_17472,N_17548);
xnor U17674 (N_17674,N_17517,N_17457);
and U17675 (N_17675,N_17572,N_17445);
and U17676 (N_17676,N_17563,N_17591);
nor U17677 (N_17677,N_17510,N_17509);
xor U17678 (N_17678,N_17486,N_17446);
xor U17679 (N_17679,N_17577,N_17482);
xnor U17680 (N_17680,N_17472,N_17594);
nand U17681 (N_17681,N_17508,N_17562);
or U17682 (N_17682,N_17562,N_17463);
nor U17683 (N_17683,N_17491,N_17471);
xnor U17684 (N_17684,N_17547,N_17565);
nor U17685 (N_17685,N_17557,N_17484);
nor U17686 (N_17686,N_17446,N_17451);
or U17687 (N_17687,N_17566,N_17553);
and U17688 (N_17688,N_17595,N_17503);
nand U17689 (N_17689,N_17450,N_17459);
and U17690 (N_17690,N_17589,N_17511);
and U17691 (N_17691,N_17502,N_17494);
xor U17692 (N_17692,N_17555,N_17450);
xor U17693 (N_17693,N_17596,N_17492);
and U17694 (N_17694,N_17445,N_17440);
nor U17695 (N_17695,N_17475,N_17451);
nand U17696 (N_17696,N_17457,N_17497);
and U17697 (N_17697,N_17585,N_17570);
nand U17698 (N_17698,N_17445,N_17444);
xnor U17699 (N_17699,N_17472,N_17484);
or U17700 (N_17700,N_17555,N_17565);
nand U17701 (N_17701,N_17517,N_17553);
nor U17702 (N_17702,N_17574,N_17455);
xnor U17703 (N_17703,N_17440,N_17451);
or U17704 (N_17704,N_17516,N_17539);
and U17705 (N_17705,N_17588,N_17485);
or U17706 (N_17706,N_17516,N_17528);
nand U17707 (N_17707,N_17560,N_17442);
or U17708 (N_17708,N_17566,N_17593);
nor U17709 (N_17709,N_17458,N_17542);
nand U17710 (N_17710,N_17556,N_17501);
and U17711 (N_17711,N_17485,N_17553);
nand U17712 (N_17712,N_17516,N_17444);
xor U17713 (N_17713,N_17544,N_17543);
xnor U17714 (N_17714,N_17497,N_17452);
nand U17715 (N_17715,N_17519,N_17494);
and U17716 (N_17716,N_17587,N_17508);
and U17717 (N_17717,N_17533,N_17506);
or U17718 (N_17718,N_17456,N_17519);
xor U17719 (N_17719,N_17562,N_17502);
nand U17720 (N_17720,N_17536,N_17567);
xnor U17721 (N_17721,N_17467,N_17473);
nand U17722 (N_17722,N_17556,N_17546);
nor U17723 (N_17723,N_17449,N_17462);
nand U17724 (N_17724,N_17588,N_17463);
or U17725 (N_17725,N_17500,N_17565);
nor U17726 (N_17726,N_17582,N_17443);
nor U17727 (N_17727,N_17518,N_17594);
nand U17728 (N_17728,N_17481,N_17568);
xor U17729 (N_17729,N_17499,N_17513);
or U17730 (N_17730,N_17578,N_17559);
and U17731 (N_17731,N_17453,N_17480);
xnor U17732 (N_17732,N_17562,N_17482);
or U17733 (N_17733,N_17527,N_17460);
or U17734 (N_17734,N_17529,N_17452);
nor U17735 (N_17735,N_17463,N_17526);
nand U17736 (N_17736,N_17467,N_17571);
and U17737 (N_17737,N_17495,N_17578);
nand U17738 (N_17738,N_17510,N_17444);
nand U17739 (N_17739,N_17473,N_17484);
xnor U17740 (N_17740,N_17459,N_17455);
or U17741 (N_17741,N_17470,N_17484);
xor U17742 (N_17742,N_17512,N_17547);
nand U17743 (N_17743,N_17544,N_17593);
xor U17744 (N_17744,N_17531,N_17599);
and U17745 (N_17745,N_17565,N_17518);
or U17746 (N_17746,N_17550,N_17459);
and U17747 (N_17747,N_17579,N_17469);
nand U17748 (N_17748,N_17503,N_17457);
nor U17749 (N_17749,N_17440,N_17550);
xor U17750 (N_17750,N_17590,N_17571);
nor U17751 (N_17751,N_17505,N_17523);
nand U17752 (N_17752,N_17491,N_17451);
and U17753 (N_17753,N_17522,N_17584);
nand U17754 (N_17754,N_17516,N_17542);
or U17755 (N_17755,N_17589,N_17486);
nor U17756 (N_17756,N_17569,N_17526);
nor U17757 (N_17757,N_17567,N_17482);
xnor U17758 (N_17758,N_17559,N_17505);
nor U17759 (N_17759,N_17445,N_17551);
and U17760 (N_17760,N_17703,N_17648);
nor U17761 (N_17761,N_17671,N_17737);
xnor U17762 (N_17762,N_17603,N_17616);
and U17763 (N_17763,N_17756,N_17646);
or U17764 (N_17764,N_17684,N_17744);
nand U17765 (N_17765,N_17759,N_17640);
and U17766 (N_17766,N_17696,N_17641);
nand U17767 (N_17767,N_17625,N_17618);
nand U17768 (N_17768,N_17712,N_17733);
xnor U17769 (N_17769,N_17617,N_17729);
nand U17770 (N_17770,N_17693,N_17645);
nand U17771 (N_17771,N_17687,N_17615);
nor U17772 (N_17772,N_17680,N_17723);
or U17773 (N_17773,N_17601,N_17732);
xor U17774 (N_17774,N_17686,N_17678);
nor U17775 (N_17775,N_17716,N_17635);
xnor U17776 (N_17776,N_17690,N_17624);
nand U17777 (N_17777,N_17639,N_17644);
or U17778 (N_17778,N_17629,N_17606);
xnor U17779 (N_17779,N_17630,N_17749);
nor U17780 (N_17780,N_17745,N_17621);
or U17781 (N_17781,N_17655,N_17662);
and U17782 (N_17782,N_17750,N_17682);
or U17783 (N_17783,N_17698,N_17734);
nor U17784 (N_17784,N_17674,N_17642);
xnor U17785 (N_17785,N_17608,N_17620);
xor U17786 (N_17786,N_17746,N_17604);
nor U17787 (N_17787,N_17713,N_17681);
nor U17788 (N_17788,N_17677,N_17637);
and U17789 (N_17789,N_17758,N_17638);
nand U17790 (N_17790,N_17704,N_17720);
or U17791 (N_17791,N_17685,N_17747);
nand U17792 (N_17792,N_17697,N_17705);
or U17793 (N_17793,N_17728,N_17700);
nor U17794 (N_17794,N_17631,N_17632);
xnor U17795 (N_17795,N_17600,N_17722);
xnor U17796 (N_17796,N_17748,N_17725);
nor U17797 (N_17797,N_17717,N_17643);
xor U17798 (N_17798,N_17741,N_17649);
and U17799 (N_17799,N_17730,N_17669);
xnor U17800 (N_17800,N_17663,N_17688);
nand U17801 (N_17801,N_17719,N_17602);
nand U17802 (N_17802,N_17753,N_17679);
nand U17803 (N_17803,N_17752,N_17605);
and U17804 (N_17804,N_17736,N_17726);
or U17805 (N_17805,N_17636,N_17614);
and U17806 (N_17806,N_17709,N_17727);
nand U17807 (N_17807,N_17612,N_17665);
xor U17808 (N_17808,N_17609,N_17658);
nand U17809 (N_17809,N_17659,N_17654);
or U17810 (N_17810,N_17607,N_17743);
or U17811 (N_17811,N_17683,N_17611);
xor U17812 (N_17812,N_17652,N_17622);
nand U17813 (N_17813,N_17626,N_17754);
or U17814 (N_17814,N_17755,N_17657);
nand U17815 (N_17815,N_17708,N_17735);
nand U17816 (N_17816,N_17692,N_17738);
nand U17817 (N_17817,N_17660,N_17647);
or U17818 (N_17818,N_17628,N_17714);
and U17819 (N_17819,N_17691,N_17613);
nand U17820 (N_17820,N_17673,N_17664);
or U17821 (N_17821,N_17751,N_17715);
xnor U17822 (N_17822,N_17670,N_17675);
nand U17823 (N_17823,N_17651,N_17661);
or U17824 (N_17824,N_17731,N_17711);
or U17825 (N_17825,N_17653,N_17672);
or U17826 (N_17826,N_17666,N_17721);
and U17827 (N_17827,N_17656,N_17718);
or U17828 (N_17828,N_17740,N_17650);
xor U17829 (N_17829,N_17667,N_17634);
or U17830 (N_17830,N_17724,N_17706);
and U17831 (N_17831,N_17695,N_17619);
or U17832 (N_17832,N_17757,N_17699);
or U17833 (N_17833,N_17710,N_17627);
nor U17834 (N_17834,N_17707,N_17694);
or U17835 (N_17835,N_17633,N_17676);
nand U17836 (N_17836,N_17668,N_17623);
or U17837 (N_17837,N_17689,N_17610);
xor U17838 (N_17838,N_17742,N_17702);
nand U17839 (N_17839,N_17701,N_17739);
xor U17840 (N_17840,N_17735,N_17733);
xor U17841 (N_17841,N_17749,N_17736);
nor U17842 (N_17842,N_17685,N_17710);
nor U17843 (N_17843,N_17673,N_17624);
and U17844 (N_17844,N_17614,N_17605);
or U17845 (N_17845,N_17675,N_17722);
and U17846 (N_17846,N_17697,N_17726);
and U17847 (N_17847,N_17687,N_17624);
and U17848 (N_17848,N_17717,N_17675);
xor U17849 (N_17849,N_17634,N_17612);
nand U17850 (N_17850,N_17750,N_17621);
xnor U17851 (N_17851,N_17692,N_17627);
xor U17852 (N_17852,N_17729,N_17700);
xor U17853 (N_17853,N_17681,N_17690);
nand U17854 (N_17854,N_17691,N_17728);
and U17855 (N_17855,N_17617,N_17612);
xnor U17856 (N_17856,N_17728,N_17750);
xnor U17857 (N_17857,N_17743,N_17645);
or U17858 (N_17858,N_17731,N_17617);
and U17859 (N_17859,N_17733,N_17605);
or U17860 (N_17860,N_17663,N_17629);
or U17861 (N_17861,N_17635,N_17749);
nand U17862 (N_17862,N_17717,N_17651);
or U17863 (N_17863,N_17622,N_17645);
xor U17864 (N_17864,N_17602,N_17654);
and U17865 (N_17865,N_17668,N_17622);
and U17866 (N_17866,N_17624,N_17620);
nand U17867 (N_17867,N_17638,N_17706);
nor U17868 (N_17868,N_17732,N_17719);
xor U17869 (N_17869,N_17604,N_17654);
and U17870 (N_17870,N_17712,N_17641);
nand U17871 (N_17871,N_17689,N_17708);
xnor U17872 (N_17872,N_17642,N_17742);
nand U17873 (N_17873,N_17659,N_17713);
nor U17874 (N_17874,N_17720,N_17677);
nand U17875 (N_17875,N_17729,N_17607);
nor U17876 (N_17876,N_17607,N_17686);
and U17877 (N_17877,N_17673,N_17705);
or U17878 (N_17878,N_17634,N_17706);
nor U17879 (N_17879,N_17697,N_17625);
nand U17880 (N_17880,N_17622,N_17729);
or U17881 (N_17881,N_17752,N_17632);
nor U17882 (N_17882,N_17743,N_17663);
nor U17883 (N_17883,N_17712,N_17623);
xnor U17884 (N_17884,N_17669,N_17648);
or U17885 (N_17885,N_17611,N_17739);
or U17886 (N_17886,N_17733,N_17682);
xor U17887 (N_17887,N_17701,N_17709);
and U17888 (N_17888,N_17633,N_17689);
xnor U17889 (N_17889,N_17611,N_17684);
and U17890 (N_17890,N_17721,N_17668);
and U17891 (N_17891,N_17624,N_17619);
nand U17892 (N_17892,N_17663,N_17712);
and U17893 (N_17893,N_17705,N_17663);
or U17894 (N_17894,N_17643,N_17736);
or U17895 (N_17895,N_17628,N_17639);
nor U17896 (N_17896,N_17625,N_17680);
nor U17897 (N_17897,N_17625,N_17744);
nor U17898 (N_17898,N_17607,N_17720);
nand U17899 (N_17899,N_17663,N_17754);
and U17900 (N_17900,N_17624,N_17681);
and U17901 (N_17901,N_17619,N_17730);
and U17902 (N_17902,N_17614,N_17704);
and U17903 (N_17903,N_17610,N_17656);
and U17904 (N_17904,N_17737,N_17629);
or U17905 (N_17905,N_17632,N_17714);
nor U17906 (N_17906,N_17720,N_17636);
nand U17907 (N_17907,N_17691,N_17627);
and U17908 (N_17908,N_17719,N_17703);
and U17909 (N_17909,N_17670,N_17695);
and U17910 (N_17910,N_17722,N_17754);
xnor U17911 (N_17911,N_17677,N_17734);
nand U17912 (N_17912,N_17711,N_17697);
or U17913 (N_17913,N_17649,N_17602);
xnor U17914 (N_17914,N_17701,N_17693);
nand U17915 (N_17915,N_17722,N_17743);
xnor U17916 (N_17916,N_17654,N_17664);
and U17917 (N_17917,N_17668,N_17730);
nor U17918 (N_17918,N_17696,N_17684);
or U17919 (N_17919,N_17718,N_17695);
nand U17920 (N_17920,N_17781,N_17908);
xnor U17921 (N_17921,N_17852,N_17892);
or U17922 (N_17922,N_17903,N_17853);
nor U17923 (N_17923,N_17856,N_17810);
nor U17924 (N_17924,N_17907,N_17896);
or U17925 (N_17925,N_17760,N_17769);
and U17926 (N_17926,N_17763,N_17899);
nand U17927 (N_17927,N_17880,N_17799);
or U17928 (N_17928,N_17774,N_17775);
xnor U17929 (N_17929,N_17886,N_17883);
and U17930 (N_17930,N_17788,N_17868);
xor U17931 (N_17931,N_17767,N_17790);
nand U17932 (N_17932,N_17772,N_17794);
nor U17933 (N_17933,N_17806,N_17793);
and U17934 (N_17934,N_17796,N_17834);
xor U17935 (N_17935,N_17818,N_17800);
nor U17936 (N_17936,N_17837,N_17863);
nand U17937 (N_17937,N_17808,N_17839);
nand U17938 (N_17938,N_17885,N_17911);
nor U17939 (N_17939,N_17768,N_17916);
xnor U17940 (N_17940,N_17847,N_17821);
or U17941 (N_17941,N_17840,N_17783);
or U17942 (N_17942,N_17838,N_17872);
nand U17943 (N_17943,N_17813,N_17773);
nand U17944 (N_17944,N_17841,N_17833);
or U17945 (N_17945,N_17902,N_17829);
xnor U17946 (N_17946,N_17785,N_17875);
xor U17947 (N_17947,N_17910,N_17823);
xor U17948 (N_17948,N_17848,N_17845);
nor U17949 (N_17949,N_17913,N_17895);
nor U17950 (N_17950,N_17814,N_17816);
nand U17951 (N_17951,N_17827,N_17844);
nor U17952 (N_17952,N_17897,N_17822);
xor U17953 (N_17953,N_17820,N_17878);
nand U17954 (N_17954,N_17851,N_17807);
and U17955 (N_17955,N_17843,N_17867);
nand U17956 (N_17956,N_17915,N_17854);
nand U17957 (N_17957,N_17792,N_17874);
xnor U17958 (N_17958,N_17906,N_17869);
or U17959 (N_17959,N_17836,N_17779);
or U17960 (N_17960,N_17861,N_17876);
xor U17961 (N_17961,N_17776,N_17797);
xnor U17962 (N_17962,N_17771,N_17761);
and U17963 (N_17963,N_17842,N_17786);
nand U17964 (N_17964,N_17884,N_17909);
and U17965 (N_17965,N_17887,N_17871);
nand U17966 (N_17966,N_17789,N_17804);
nand U17967 (N_17967,N_17798,N_17824);
and U17968 (N_17968,N_17860,N_17855);
or U17969 (N_17969,N_17811,N_17762);
xnor U17970 (N_17970,N_17905,N_17894);
and U17971 (N_17971,N_17826,N_17801);
or U17972 (N_17972,N_17805,N_17901);
nand U17973 (N_17973,N_17914,N_17893);
nor U17974 (N_17974,N_17912,N_17819);
and U17975 (N_17975,N_17770,N_17889);
xnor U17976 (N_17976,N_17780,N_17917);
nand U17977 (N_17977,N_17891,N_17859);
nor U17978 (N_17978,N_17835,N_17803);
nor U17979 (N_17979,N_17898,N_17815);
xnor U17980 (N_17980,N_17825,N_17830);
nor U17981 (N_17981,N_17764,N_17877);
xor U17982 (N_17982,N_17904,N_17802);
nor U17983 (N_17983,N_17866,N_17890);
or U17984 (N_17984,N_17778,N_17873);
nor U17985 (N_17985,N_17812,N_17795);
and U17986 (N_17986,N_17900,N_17865);
nor U17987 (N_17987,N_17787,N_17817);
and U17988 (N_17988,N_17858,N_17782);
xnor U17989 (N_17989,N_17846,N_17882);
nor U17990 (N_17990,N_17850,N_17832);
or U17991 (N_17991,N_17849,N_17888);
nor U17992 (N_17992,N_17777,N_17864);
and U17993 (N_17993,N_17766,N_17791);
nand U17994 (N_17994,N_17809,N_17870);
nand U17995 (N_17995,N_17857,N_17919);
or U17996 (N_17996,N_17831,N_17765);
nor U17997 (N_17997,N_17881,N_17862);
nand U17998 (N_17998,N_17918,N_17784);
xor U17999 (N_17999,N_17828,N_17879);
nand U18000 (N_18000,N_17871,N_17863);
nand U18001 (N_18001,N_17875,N_17908);
nand U18002 (N_18002,N_17798,N_17890);
or U18003 (N_18003,N_17855,N_17795);
and U18004 (N_18004,N_17836,N_17781);
xnor U18005 (N_18005,N_17875,N_17862);
and U18006 (N_18006,N_17855,N_17829);
nand U18007 (N_18007,N_17838,N_17864);
nor U18008 (N_18008,N_17848,N_17861);
nand U18009 (N_18009,N_17783,N_17827);
nor U18010 (N_18010,N_17801,N_17820);
xor U18011 (N_18011,N_17916,N_17770);
and U18012 (N_18012,N_17914,N_17834);
nor U18013 (N_18013,N_17778,N_17890);
nor U18014 (N_18014,N_17862,N_17888);
xor U18015 (N_18015,N_17769,N_17869);
and U18016 (N_18016,N_17867,N_17792);
xnor U18017 (N_18017,N_17897,N_17857);
and U18018 (N_18018,N_17884,N_17863);
xor U18019 (N_18019,N_17910,N_17831);
and U18020 (N_18020,N_17813,N_17892);
nor U18021 (N_18021,N_17790,N_17900);
or U18022 (N_18022,N_17892,N_17910);
or U18023 (N_18023,N_17816,N_17910);
nand U18024 (N_18024,N_17905,N_17875);
nand U18025 (N_18025,N_17869,N_17907);
or U18026 (N_18026,N_17816,N_17872);
and U18027 (N_18027,N_17778,N_17820);
nand U18028 (N_18028,N_17787,N_17915);
nor U18029 (N_18029,N_17836,N_17843);
nand U18030 (N_18030,N_17855,N_17863);
nand U18031 (N_18031,N_17869,N_17879);
or U18032 (N_18032,N_17908,N_17856);
nor U18033 (N_18033,N_17831,N_17855);
or U18034 (N_18034,N_17870,N_17784);
and U18035 (N_18035,N_17762,N_17881);
xor U18036 (N_18036,N_17902,N_17800);
or U18037 (N_18037,N_17804,N_17795);
nor U18038 (N_18038,N_17823,N_17901);
and U18039 (N_18039,N_17823,N_17853);
or U18040 (N_18040,N_17849,N_17875);
nand U18041 (N_18041,N_17900,N_17841);
and U18042 (N_18042,N_17829,N_17828);
or U18043 (N_18043,N_17812,N_17790);
or U18044 (N_18044,N_17767,N_17782);
or U18045 (N_18045,N_17891,N_17787);
nor U18046 (N_18046,N_17834,N_17885);
nor U18047 (N_18047,N_17773,N_17769);
nor U18048 (N_18048,N_17859,N_17767);
xor U18049 (N_18049,N_17807,N_17820);
and U18050 (N_18050,N_17876,N_17859);
nand U18051 (N_18051,N_17839,N_17861);
nor U18052 (N_18052,N_17892,N_17859);
and U18053 (N_18053,N_17894,N_17866);
and U18054 (N_18054,N_17772,N_17805);
nor U18055 (N_18055,N_17798,N_17793);
nand U18056 (N_18056,N_17897,N_17761);
nor U18057 (N_18057,N_17772,N_17878);
or U18058 (N_18058,N_17791,N_17915);
xnor U18059 (N_18059,N_17807,N_17833);
xor U18060 (N_18060,N_17863,N_17780);
and U18061 (N_18061,N_17846,N_17776);
or U18062 (N_18062,N_17826,N_17767);
or U18063 (N_18063,N_17910,N_17884);
nor U18064 (N_18064,N_17872,N_17897);
xnor U18065 (N_18065,N_17904,N_17775);
or U18066 (N_18066,N_17813,N_17862);
nand U18067 (N_18067,N_17882,N_17790);
and U18068 (N_18068,N_17892,N_17845);
nor U18069 (N_18069,N_17875,N_17821);
or U18070 (N_18070,N_17820,N_17854);
nor U18071 (N_18071,N_17857,N_17846);
xor U18072 (N_18072,N_17801,N_17916);
xor U18073 (N_18073,N_17892,N_17908);
or U18074 (N_18074,N_17917,N_17828);
nand U18075 (N_18075,N_17838,N_17801);
nand U18076 (N_18076,N_17767,N_17872);
xor U18077 (N_18077,N_17840,N_17865);
nor U18078 (N_18078,N_17802,N_17846);
and U18079 (N_18079,N_17774,N_17823);
nand U18080 (N_18080,N_17935,N_18020);
nor U18081 (N_18081,N_18002,N_17989);
or U18082 (N_18082,N_18027,N_17965);
nor U18083 (N_18083,N_17944,N_18074);
nand U18084 (N_18084,N_18062,N_17995);
and U18085 (N_18085,N_18075,N_18041);
nand U18086 (N_18086,N_18031,N_18011);
or U18087 (N_18087,N_18036,N_18021);
nand U18088 (N_18088,N_18069,N_17987);
or U18089 (N_18089,N_17959,N_18042);
xor U18090 (N_18090,N_18078,N_18033);
nand U18091 (N_18091,N_17940,N_18000);
nor U18092 (N_18092,N_17977,N_17963);
xor U18093 (N_18093,N_17985,N_17996);
or U18094 (N_18094,N_18015,N_17924);
or U18095 (N_18095,N_18070,N_17973);
nand U18096 (N_18096,N_18073,N_17981);
nand U18097 (N_18097,N_17922,N_17999);
nand U18098 (N_18098,N_17964,N_17950);
xnor U18099 (N_18099,N_17947,N_17983);
or U18100 (N_18100,N_18037,N_17994);
and U18101 (N_18101,N_18049,N_18052);
and U18102 (N_18102,N_18014,N_17957);
xor U18103 (N_18103,N_17980,N_18022);
xor U18104 (N_18104,N_18076,N_18056);
nor U18105 (N_18105,N_17978,N_17945);
nand U18106 (N_18106,N_18030,N_17921);
nor U18107 (N_18107,N_17993,N_18043);
and U18108 (N_18108,N_17953,N_18026);
or U18109 (N_18109,N_17939,N_18006);
xor U18110 (N_18110,N_18072,N_18035);
or U18111 (N_18111,N_18045,N_18009);
nand U18112 (N_18112,N_17969,N_18064);
and U18113 (N_18113,N_18029,N_17920);
nand U18114 (N_18114,N_17982,N_17960);
xnor U18115 (N_18115,N_17984,N_17943);
or U18116 (N_18116,N_18058,N_18051);
nand U18117 (N_18117,N_17933,N_17923);
xnor U18118 (N_18118,N_17928,N_18008);
or U18119 (N_18119,N_18071,N_17949);
nor U18120 (N_18120,N_17942,N_18040);
and U18121 (N_18121,N_18005,N_18010);
xnor U18122 (N_18122,N_18038,N_18077);
nor U18123 (N_18123,N_18061,N_18050);
and U18124 (N_18124,N_17972,N_17974);
and U18125 (N_18125,N_18046,N_17931);
nand U18126 (N_18126,N_17956,N_17970);
nor U18127 (N_18127,N_17979,N_17929);
nor U18128 (N_18128,N_17968,N_18044);
xor U18129 (N_18129,N_18001,N_17990);
or U18130 (N_18130,N_18004,N_17988);
xor U18131 (N_18131,N_18019,N_17948);
nand U18132 (N_18132,N_18079,N_18012);
nor U18133 (N_18133,N_17976,N_17951);
xor U18134 (N_18134,N_17954,N_18028);
nor U18135 (N_18135,N_18024,N_17926);
and U18136 (N_18136,N_17991,N_18053);
nor U18137 (N_18137,N_17955,N_17941);
nand U18138 (N_18138,N_18032,N_17952);
nor U18139 (N_18139,N_18023,N_17946);
and U18140 (N_18140,N_17938,N_17927);
or U18141 (N_18141,N_18039,N_17966);
and U18142 (N_18142,N_17925,N_18059);
nand U18143 (N_18143,N_18047,N_17975);
nor U18144 (N_18144,N_18060,N_17998);
nand U18145 (N_18145,N_18017,N_17986);
or U18146 (N_18146,N_18003,N_18054);
xor U18147 (N_18147,N_17967,N_17958);
xnor U18148 (N_18148,N_17937,N_17930);
nand U18149 (N_18149,N_18048,N_18055);
nor U18150 (N_18150,N_18007,N_18013);
xor U18151 (N_18151,N_17992,N_17961);
nor U18152 (N_18152,N_18057,N_18018);
xor U18153 (N_18153,N_18067,N_18034);
xnor U18154 (N_18154,N_18068,N_18016);
and U18155 (N_18155,N_17936,N_18063);
or U18156 (N_18156,N_17997,N_17932);
nand U18157 (N_18157,N_18066,N_17934);
nor U18158 (N_18158,N_18065,N_17971);
or U18159 (N_18159,N_17962,N_18025);
xor U18160 (N_18160,N_18034,N_18070);
nand U18161 (N_18161,N_18043,N_18012);
nor U18162 (N_18162,N_17983,N_18060);
and U18163 (N_18163,N_17988,N_18052);
nand U18164 (N_18164,N_18033,N_17962);
nand U18165 (N_18165,N_18061,N_17973);
or U18166 (N_18166,N_18038,N_17964);
nand U18167 (N_18167,N_18014,N_17958);
and U18168 (N_18168,N_18010,N_18055);
nor U18169 (N_18169,N_18049,N_17999);
nand U18170 (N_18170,N_18053,N_17992);
nor U18171 (N_18171,N_18063,N_18051);
or U18172 (N_18172,N_17948,N_17935);
xnor U18173 (N_18173,N_18058,N_18075);
or U18174 (N_18174,N_18008,N_18000);
nor U18175 (N_18175,N_18069,N_17979);
and U18176 (N_18176,N_18070,N_17952);
or U18177 (N_18177,N_17985,N_18038);
xor U18178 (N_18178,N_18001,N_18066);
nor U18179 (N_18179,N_17965,N_17974);
or U18180 (N_18180,N_17968,N_18025);
or U18181 (N_18181,N_18031,N_18015);
and U18182 (N_18182,N_17928,N_17953);
and U18183 (N_18183,N_18038,N_18071);
and U18184 (N_18184,N_17971,N_18078);
and U18185 (N_18185,N_17974,N_17934);
or U18186 (N_18186,N_18077,N_18028);
or U18187 (N_18187,N_18019,N_17962);
and U18188 (N_18188,N_17945,N_18059);
and U18189 (N_18189,N_18079,N_17985);
nor U18190 (N_18190,N_17960,N_17950);
nand U18191 (N_18191,N_17941,N_17920);
or U18192 (N_18192,N_18031,N_18027);
or U18193 (N_18193,N_18061,N_17960);
nand U18194 (N_18194,N_18016,N_18001);
xnor U18195 (N_18195,N_18038,N_18061);
and U18196 (N_18196,N_18036,N_17997);
and U18197 (N_18197,N_18006,N_17980);
nand U18198 (N_18198,N_18040,N_18021);
nor U18199 (N_18199,N_17934,N_18042);
nor U18200 (N_18200,N_18053,N_17924);
or U18201 (N_18201,N_18040,N_18071);
or U18202 (N_18202,N_18026,N_17962);
nand U18203 (N_18203,N_18002,N_18026);
nor U18204 (N_18204,N_18038,N_18067);
or U18205 (N_18205,N_18033,N_18019);
xor U18206 (N_18206,N_17939,N_18043);
or U18207 (N_18207,N_17938,N_18059);
or U18208 (N_18208,N_18034,N_18053);
or U18209 (N_18209,N_18051,N_18027);
and U18210 (N_18210,N_17980,N_18005);
and U18211 (N_18211,N_17930,N_18034);
nor U18212 (N_18212,N_17956,N_17920);
and U18213 (N_18213,N_18058,N_17990);
or U18214 (N_18214,N_18070,N_18047);
nor U18215 (N_18215,N_17928,N_18029);
or U18216 (N_18216,N_17921,N_17991);
or U18217 (N_18217,N_17921,N_17957);
and U18218 (N_18218,N_18058,N_17935);
nand U18219 (N_18219,N_17974,N_18038);
nor U18220 (N_18220,N_18020,N_18026);
and U18221 (N_18221,N_17962,N_18045);
and U18222 (N_18222,N_18053,N_18012);
xor U18223 (N_18223,N_18008,N_18051);
or U18224 (N_18224,N_18005,N_18011);
xor U18225 (N_18225,N_17929,N_17993);
xor U18226 (N_18226,N_17994,N_18035);
and U18227 (N_18227,N_18065,N_18030);
nand U18228 (N_18228,N_18020,N_17964);
nor U18229 (N_18229,N_18019,N_18031);
xnor U18230 (N_18230,N_18058,N_18040);
or U18231 (N_18231,N_18058,N_18067);
or U18232 (N_18232,N_18070,N_17925);
or U18233 (N_18233,N_18078,N_17945);
and U18234 (N_18234,N_18048,N_18006);
nand U18235 (N_18235,N_17979,N_17923);
nand U18236 (N_18236,N_18062,N_18022);
and U18237 (N_18237,N_18063,N_17962);
or U18238 (N_18238,N_17936,N_18059);
nor U18239 (N_18239,N_17924,N_18043);
xor U18240 (N_18240,N_18219,N_18093);
and U18241 (N_18241,N_18106,N_18145);
nand U18242 (N_18242,N_18108,N_18177);
or U18243 (N_18243,N_18155,N_18110);
and U18244 (N_18244,N_18089,N_18238);
xnor U18245 (N_18245,N_18109,N_18144);
nor U18246 (N_18246,N_18191,N_18210);
nor U18247 (N_18247,N_18149,N_18084);
or U18248 (N_18248,N_18220,N_18166);
nand U18249 (N_18249,N_18102,N_18209);
or U18250 (N_18250,N_18123,N_18185);
nor U18251 (N_18251,N_18201,N_18232);
nor U18252 (N_18252,N_18234,N_18160);
xnor U18253 (N_18253,N_18130,N_18125);
nand U18254 (N_18254,N_18158,N_18203);
nor U18255 (N_18255,N_18111,N_18099);
and U18256 (N_18256,N_18150,N_18097);
and U18257 (N_18257,N_18200,N_18133);
nand U18258 (N_18258,N_18085,N_18083);
nand U18259 (N_18259,N_18169,N_18206);
or U18260 (N_18260,N_18211,N_18100);
and U18261 (N_18261,N_18204,N_18136);
or U18262 (N_18262,N_18134,N_18222);
nand U18263 (N_18263,N_18187,N_18218);
xor U18264 (N_18264,N_18113,N_18132);
and U18265 (N_18265,N_18140,N_18226);
or U18266 (N_18266,N_18159,N_18216);
or U18267 (N_18267,N_18094,N_18090);
xor U18268 (N_18268,N_18139,N_18175);
or U18269 (N_18269,N_18167,N_18189);
xnor U18270 (N_18270,N_18137,N_18143);
xnor U18271 (N_18271,N_18118,N_18198);
and U18272 (N_18272,N_18184,N_18237);
and U18273 (N_18273,N_18229,N_18212);
nand U18274 (N_18274,N_18117,N_18152);
or U18275 (N_18275,N_18213,N_18195);
nand U18276 (N_18276,N_18171,N_18147);
and U18277 (N_18277,N_18215,N_18225);
or U18278 (N_18278,N_18214,N_18164);
and U18279 (N_18279,N_18179,N_18082);
nor U18280 (N_18280,N_18115,N_18086);
xnor U18281 (N_18281,N_18174,N_18178);
and U18282 (N_18282,N_18230,N_18194);
xor U18283 (N_18283,N_18156,N_18168);
and U18284 (N_18284,N_18221,N_18095);
xnor U18285 (N_18285,N_18188,N_18107);
nor U18286 (N_18286,N_18165,N_18239);
or U18287 (N_18287,N_18173,N_18154);
and U18288 (N_18288,N_18183,N_18129);
nor U18289 (N_18289,N_18148,N_18098);
xor U18290 (N_18290,N_18087,N_18141);
nand U18291 (N_18291,N_18151,N_18190);
nand U18292 (N_18292,N_18199,N_18081);
and U18293 (N_18293,N_18193,N_18236);
nand U18294 (N_18294,N_18224,N_18162);
nor U18295 (N_18295,N_18146,N_18091);
nand U18296 (N_18296,N_18138,N_18207);
xor U18297 (N_18297,N_18126,N_18180);
or U18298 (N_18298,N_18223,N_18202);
xor U18299 (N_18299,N_18172,N_18227);
nand U18300 (N_18300,N_18105,N_18120);
and U18301 (N_18301,N_18142,N_18186);
or U18302 (N_18302,N_18157,N_18235);
or U18303 (N_18303,N_18205,N_18182);
and U18304 (N_18304,N_18128,N_18196);
xor U18305 (N_18305,N_18119,N_18116);
xor U18306 (N_18306,N_18153,N_18103);
or U18307 (N_18307,N_18231,N_18163);
and U18308 (N_18308,N_18192,N_18112);
nor U18309 (N_18309,N_18161,N_18217);
or U18310 (N_18310,N_18233,N_18176);
or U18311 (N_18311,N_18135,N_18197);
nand U18312 (N_18312,N_18131,N_18127);
xnor U18313 (N_18313,N_18124,N_18122);
or U18314 (N_18314,N_18088,N_18080);
or U18315 (N_18315,N_18096,N_18101);
or U18316 (N_18316,N_18170,N_18114);
or U18317 (N_18317,N_18104,N_18092);
nor U18318 (N_18318,N_18121,N_18228);
xnor U18319 (N_18319,N_18181,N_18208);
nand U18320 (N_18320,N_18197,N_18198);
nand U18321 (N_18321,N_18080,N_18234);
or U18322 (N_18322,N_18199,N_18091);
nand U18323 (N_18323,N_18092,N_18183);
and U18324 (N_18324,N_18084,N_18133);
and U18325 (N_18325,N_18226,N_18189);
nor U18326 (N_18326,N_18171,N_18102);
and U18327 (N_18327,N_18206,N_18173);
and U18328 (N_18328,N_18203,N_18194);
nor U18329 (N_18329,N_18118,N_18135);
nand U18330 (N_18330,N_18219,N_18145);
nand U18331 (N_18331,N_18168,N_18192);
or U18332 (N_18332,N_18103,N_18197);
nand U18333 (N_18333,N_18088,N_18101);
or U18334 (N_18334,N_18133,N_18234);
nand U18335 (N_18335,N_18162,N_18152);
and U18336 (N_18336,N_18110,N_18235);
and U18337 (N_18337,N_18210,N_18227);
and U18338 (N_18338,N_18122,N_18123);
nor U18339 (N_18339,N_18151,N_18157);
nand U18340 (N_18340,N_18144,N_18238);
or U18341 (N_18341,N_18133,N_18159);
nor U18342 (N_18342,N_18193,N_18119);
xnor U18343 (N_18343,N_18111,N_18211);
xor U18344 (N_18344,N_18126,N_18119);
nor U18345 (N_18345,N_18143,N_18097);
nand U18346 (N_18346,N_18177,N_18139);
or U18347 (N_18347,N_18107,N_18173);
xnor U18348 (N_18348,N_18172,N_18124);
xnor U18349 (N_18349,N_18202,N_18211);
and U18350 (N_18350,N_18101,N_18178);
xnor U18351 (N_18351,N_18097,N_18121);
nand U18352 (N_18352,N_18092,N_18080);
and U18353 (N_18353,N_18080,N_18082);
xor U18354 (N_18354,N_18230,N_18114);
and U18355 (N_18355,N_18136,N_18112);
xnor U18356 (N_18356,N_18239,N_18164);
or U18357 (N_18357,N_18143,N_18160);
or U18358 (N_18358,N_18201,N_18220);
and U18359 (N_18359,N_18099,N_18121);
and U18360 (N_18360,N_18085,N_18219);
or U18361 (N_18361,N_18199,N_18161);
nand U18362 (N_18362,N_18140,N_18236);
nor U18363 (N_18363,N_18100,N_18112);
or U18364 (N_18364,N_18174,N_18134);
xnor U18365 (N_18365,N_18178,N_18158);
or U18366 (N_18366,N_18186,N_18159);
nand U18367 (N_18367,N_18171,N_18118);
xnor U18368 (N_18368,N_18124,N_18203);
and U18369 (N_18369,N_18217,N_18225);
and U18370 (N_18370,N_18104,N_18210);
or U18371 (N_18371,N_18148,N_18158);
or U18372 (N_18372,N_18168,N_18092);
nor U18373 (N_18373,N_18233,N_18152);
and U18374 (N_18374,N_18082,N_18117);
and U18375 (N_18375,N_18173,N_18143);
nor U18376 (N_18376,N_18107,N_18085);
and U18377 (N_18377,N_18178,N_18156);
xor U18378 (N_18378,N_18139,N_18158);
xor U18379 (N_18379,N_18211,N_18143);
or U18380 (N_18380,N_18146,N_18165);
xor U18381 (N_18381,N_18164,N_18112);
and U18382 (N_18382,N_18092,N_18147);
nand U18383 (N_18383,N_18213,N_18201);
or U18384 (N_18384,N_18217,N_18123);
nor U18385 (N_18385,N_18134,N_18165);
xor U18386 (N_18386,N_18094,N_18231);
nand U18387 (N_18387,N_18130,N_18092);
and U18388 (N_18388,N_18189,N_18166);
nor U18389 (N_18389,N_18086,N_18138);
and U18390 (N_18390,N_18215,N_18239);
nand U18391 (N_18391,N_18149,N_18193);
nor U18392 (N_18392,N_18222,N_18187);
and U18393 (N_18393,N_18084,N_18207);
nor U18394 (N_18394,N_18091,N_18099);
or U18395 (N_18395,N_18236,N_18110);
or U18396 (N_18396,N_18208,N_18172);
xnor U18397 (N_18397,N_18093,N_18225);
or U18398 (N_18398,N_18218,N_18154);
or U18399 (N_18399,N_18081,N_18126);
nor U18400 (N_18400,N_18353,N_18258);
or U18401 (N_18401,N_18327,N_18256);
nor U18402 (N_18402,N_18339,N_18338);
nor U18403 (N_18403,N_18300,N_18269);
xor U18404 (N_18404,N_18303,N_18297);
nand U18405 (N_18405,N_18278,N_18268);
or U18406 (N_18406,N_18249,N_18370);
or U18407 (N_18407,N_18282,N_18326);
or U18408 (N_18408,N_18250,N_18348);
nor U18409 (N_18409,N_18331,N_18379);
nor U18410 (N_18410,N_18289,N_18386);
or U18411 (N_18411,N_18365,N_18354);
xnor U18412 (N_18412,N_18364,N_18349);
or U18413 (N_18413,N_18265,N_18344);
xnor U18414 (N_18414,N_18288,N_18266);
and U18415 (N_18415,N_18387,N_18322);
nor U18416 (N_18416,N_18356,N_18377);
nor U18417 (N_18417,N_18333,N_18281);
nor U18418 (N_18418,N_18395,N_18351);
xor U18419 (N_18419,N_18315,N_18362);
and U18420 (N_18420,N_18367,N_18332);
xnor U18421 (N_18421,N_18350,N_18324);
xnor U18422 (N_18422,N_18318,N_18275);
xor U18423 (N_18423,N_18343,N_18264);
xor U18424 (N_18424,N_18301,N_18399);
nor U18425 (N_18425,N_18299,N_18274);
nor U18426 (N_18426,N_18312,N_18306);
or U18427 (N_18427,N_18316,N_18345);
nor U18428 (N_18428,N_18396,N_18261);
or U18429 (N_18429,N_18311,N_18357);
or U18430 (N_18430,N_18391,N_18393);
or U18431 (N_18431,N_18310,N_18375);
xor U18432 (N_18432,N_18245,N_18241);
or U18433 (N_18433,N_18397,N_18384);
xnor U18434 (N_18434,N_18342,N_18304);
nand U18435 (N_18435,N_18248,N_18291);
and U18436 (N_18436,N_18279,N_18368);
nand U18437 (N_18437,N_18325,N_18293);
and U18438 (N_18438,N_18390,N_18251);
nand U18439 (N_18439,N_18260,N_18321);
nand U18440 (N_18440,N_18270,N_18277);
nor U18441 (N_18441,N_18371,N_18337);
xor U18442 (N_18442,N_18243,N_18313);
xnor U18443 (N_18443,N_18254,N_18244);
xnor U18444 (N_18444,N_18271,N_18330);
nand U18445 (N_18445,N_18374,N_18319);
nor U18446 (N_18446,N_18352,N_18240);
nand U18447 (N_18447,N_18341,N_18314);
nor U18448 (N_18448,N_18292,N_18335);
xor U18449 (N_18449,N_18290,N_18252);
xnor U18450 (N_18450,N_18283,N_18328);
xor U18451 (N_18451,N_18369,N_18347);
or U18452 (N_18452,N_18273,N_18259);
and U18453 (N_18453,N_18296,N_18382);
and U18454 (N_18454,N_18383,N_18320);
and U18455 (N_18455,N_18253,N_18267);
or U18456 (N_18456,N_18360,N_18378);
or U18457 (N_18457,N_18394,N_18363);
or U18458 (N_18458,N_18398,N_18376);
xnor U18459 (N_18459,N_18295,N_18309);
and U18460 (N_18460,N_18246,N_18263);
xnor U18461 (N_18461,N_18247,N_18334);
nand U18462 (N_18462,N_18308,N_18255);
nand U18463 (N_18463,N_18340,N_18329);
or U18464 (N_18464,N_18346,N_18381);
nor U18465 (N_18465,N_18272,N_18294);
xnor U18466 (N_18466,N_18305,N_18359);
or U18467 (N_18467,N_18286,N_18372);
xnor U18468 (N_18468,N_18257,N_18385);
and U18469 (N_18469,N_18284,N_18380);
xor U18470 (N_18470,N_18317,N_18336);
or U18471 (N_18471,N_18287,N_18361);
xor U18472 (N_18472,N_18392,N_18388);
and U18473 (N_18473,N_18307,N_18358);
and U18474 (N_18474,N_18280,N_18276);
nand U18475 (N_18475,N_18262,N_18323);
or U18476 (N_18476,N_18285,N_18355);
and U18477 (N_18477,N_18366,N_18242);
and U18478 (N_18478,N_18302,N_18373);
and U18479 (N_18479,N_18298,N_18389);
xnor U18480 (N_18480,N_18282,N_18300);
or U18481 (N_18481,N_18243,N_18364);
nand U18482 (N_18482,N_18319,N_18329);
nand U18483 (N_18483,N_18309,N_18368);
nand U18484 (N_18484,N_18333,N_18365);
or U18485 (N_18485,N_18345,N_18301);
xnor U18486 (N_18486,N_18316,N_18286);
nand U18487 (N_18487,N_18241,N_18334);
nand U18488 (N_18488,N_18350,N_18273);
and U18489 (N_18489,N_18341,N_18371);
or U18490 (N_18490,N_18382,N_18345);
and U18491 (N_18491,N_18309,N_18364);
nand U18492 (N_18492,N_18310,N_18397);
xor U18493 (N_18493,N_18271,N_18293);
nand U18494 (N_18494,N_18297,N_18301);
and U18495 (N_18495,N_18240,N_18371);
xor U18496 (N_18496,N_18255,N_18298);
xor U18497 (N_18497,N_18253,N_18244);
nand U18498 (N_18498,N_18357,N_18242);
or U18499 (N_18499,N_18378,N_18288);
and U18500 (N_18500,N_18329,N_18333);
or U18501 (N_18501,N_18370,N_18377);
or U18502 (N_18502,N_18361,N_18363);
nor U18503 (N_18503,N_18373,N_18297);
xor U18504 (N_18504,N_18257,N_18368);
nand U18505 (N_18505,N_18357,N_18332);
and U18506 (N_18506,N_18321,N_18369);
xnor U18507 (N_18507,N_18298,N_18327);
nand U18508 (N_18508,N_18364,N_18252);
and U18509 (N_18509,N_18359,N_18321);
or U18510 (N_18510,N_18296,N_18368);
and U18511 (N_18511,N_18252,N_18323);
xnor U18512 (N_18512,N_18320,N_18374);
xor U18513 (N_18513,N_18289,N_18353);
and U18514 (N_18514,N_18254,N_18266);
xor U18515 (N_18515,N_18240,N_18262);
nand U18516 (N_18516,N_18242,N_18331);
or U18517 (N_18517,N_18342,N_18343);
and U18518 (N_18518,N_18320,N_18332);
nand U18519 (N_18519,N_18301,N_18260);
nand U18520 (N_18520,N_18294,N_18326);
nand U18521 (N_18521,N_18324,N_18359);
or U18522 (N_18522,N_18247,N_18270);
and U18523 (N_18523,N_18343,N_18326);
xnor U18524 (N_18524,N_18313,N_18269);
and U18525 (N_18525,N_18314,N_18355);
xor U18526 (N_18526,N_18299,N_18297);
and U18527 (N_18527,N_18383,N_18345);
nor U18528 (N_18528,N_18342,N_18385);
or U18529 (N_18529,N_18292,N_18295);
nor U18530 (N_18530,N_18259,N_18260);
or U18531 (N_18531,N_18319,N_18336);
nand U18532 (N_18532,N_18299,N_18248);
xor U18533 (N_18533,N_18362,N_18309);
and U18534 (N_18534,N_18317,N_18376);
or U18535 (N_18535,N_18355,N_18295);
nand U18536 (N_18536,N_18255,N_18387);
or U18537 (N_18537,N_18364,N_18306);
nand U18538 (N_18538,N_18243,N_18386);
xnor U18539 (N_18539,N_18319,N_18310);
nand U18540 (N_18540,N_18339,N_18351);
nor U18541 (N_18541,N_18287,N_18299);
nor U18542 (N_18542,N_18247,N_18399);
and U18543 (N_18543,N_18253,N_18257);
or U18544 (N_18544,N_18332,N_18373);
and U18545 (N_18545,N_18280,N_18356);
nand U18546 (N_18546,N_18313,N_18271);
nand U18547 (N_18547,N_18356,N_18264);
and U18548 (N_18548,N_18358,N_18249);
nand U18549 (N_18549,N_18314,N_18254);
nand U18550 (N_18550,N_18296,N_18322);
nor U18551 (N_18551,N_18273,N_18244);
nor U18552 (N_18552,N_18369,N_18325);
or U18553 (N_18553,N_18275,N_18297);
and U18554 (N_18554,N_18394,N_18354);
or U18555 (N_18555,N_18308,N_18373);
xor U18556 (N_18556,N_18246,N_18372);
nand U18557 (N_18557,N_18386,N_18399);
nand U18558 (N_18558,N_18306,N_18311);
and U18559 (N_18559,N_18304,N_18325);
xor U18560 (N_18560,N_18410,N_18472);
nand U18561 (N_18561,N_18435,N_18434);
nand U18562 (N_18562,N_18474,N_18408);
nor U18563 (N_18563,N_18527,N_18430);
or U18564 (N_18564,N_18461,N_18510);
and U18565 (N_18565,N_18543,N_18485);
and U18566 (N_18566,N_18419,N_18489);
and U18567 (N_18567,N_18421,N_18509);
xor U18568 (N_18568,N_18450,N_18463);
or U18569 (N_18569,N_18529,N_18401);
or U18570 (N_18570,N_18441,N_18455);
xnor U18571 (N_18571,N_18500,N_18460);
nand U18572 (N_18572,N_18414,N_18512);
or U18573 (N_18573,N_18518,N_18483);
xnor U18574 (N_18574,N_18535,N_18515);
xnor U18575 (N_18575,N_18487,N_18456);
or U18576 (N_18576,N_18537,N_18536);
nor U18577 (N_18577,N_18439,N_18502);
nor U18578 (N_18578,N_18523,N_18406);
and U18579 (N_18579,N_18422,N_18533);
and U18580 (N_18580,N_18544,N_18541);
xnor U18581 (N_18581,N_18548,N_18480);
and U18582 (N_18582,N_18504,N_18442);
nor U18583 (N_18583,N_18492,N_18416);
and U18584 (N_18584,N_18400,N_18545);
and U18585 (N_18585,N_18464,N_18458);
and U18586 (N_18586,N_18433,N_18481);
or U18587 (N_18587,N_18501,N_18443);
nor U18588 (N_18588,N_18553,N_18417);
xor U18589 (N_18589,N_18547,N_18552);
nor U18590 (N_18590,N_18542,N_18484);
and U18591 (N_18591,N_18444,N_18428);
xor U18592 (N_18592,N_18491,N_18412);
or U18593 (N_18593,N_18448,N_18475);
or U18594 (N_18594,N_18521,N_18511);
xnor U18595 (N_18595,N_18415,N_18516);
and U18596 (N_18596,N_18532,N_18452);
or U18597 (N_18597,N_18470,N_18559);
xor U18598 (N_18598,N_18478,N_18497);
xor U18599 (N_18599,N_18438,N_18445);
or U18600 (N_18600,N_18507,N_18498);
xor U18601 (N_18601,N_18505,N_18517);
and U18602 (N_18602,N_18409,N_18457);
nor U18603 (N_18603,N_18465,N_18479);
nand U18604 (N_18604,N_18528,N_18440);
or U18605 (N_18605,N_18437,N_18469);
or U18606 (N_18606,N_18534,N_18432);
or U18607 (N_18607,N_18436,N_18420);
nand U18608 (N_18608,N_18495,N_18524);
nand U18609 (N_18609,N_18519,N_18473);
and U18610 (N_18610,N_18427,N_18467);
and U18611 (N_18611,N_18551,N_18411);
xor U18612 (N_18612,N_18531,N_18538);
and U18613 (N_18613,N_18447,N_18558);
nor U18614 (N_18614,N_18407,N_18468);
nand U18615 (N_18615,N_18555,N_18546);
nor U18616 (N_18616,N_18466,N_18549);
nor U18617 (N_18617,N_18508,N_18493);
nand U18618 (N_18618,N_18506,N_18503);
and U18619 (N_18619,N_18540,N_18418);
nand U18620 (N_18620,N_18404,N_18431);
nand U18621 (N_18621,N_18488,N_18522);
nor U18622 (N_18622,N_18539,N_18471);
nand U18623 (N_18623,N_18423,N_18454);
nor U18624 (N_18624,N_18449,N_18446);
xor U18625 (N_18625,N_18482,N_18490);
nand U18626 (N_18626,N_18462,N_18425);
nand U18627 (N_18627,N_18550,N_18403);
and U18628 (N_18628,N_18496,N_18453);
nor U18629 (N_18629,N_18557,N_18494);
nor U18630 (N_18630,N_18476,N_18477);
nand U18631 (N_18631,N_18556,N_18525);
xor U18632 (N_18632,N_18514,N_18424);
or U18633 (N_18633,N_18413,N_18526);
nor U18634 (N_18634,N_18486,N_18402);
or U18635 (N_18635,N_18520,N_18405);
xor U18636 (N_18636,N_18513,N_18530);
xor U18637 (N_18637,N_18429,N_18459);
nor U18638 (N_18638,N_18554,N_18426);
xnor U18639 (N_18639,N_18451,N_18499);
or U18640 (N_18640,N_18415,N_18437);
or U18641 (N_18641,N_18531,N_18446);
nor U18642 (N_18642,N_18501,N_18539);
xnor U18643 (N_18643,N_18537,N_18466);
nor U18644 (N_18644,N_18444,N_18520);
xor U18645 (N_18645,N_18450,N_18476);
nor U18646 (N_18646,N_18461,N_18401);
or U18647 (N_18647,N_18521,N_18463);
xnor U18648 (N_18648,N_18514,N_18538);
nor U18649 (N_18649,N_18433,N_18413);
nor U18650 (N_18650,N_18505,N_18536);
and U18651 (N_18651,N_18426,N_18462);
xor U18652 (N_18652,N_18441,N_18492);
xor U18653 (N_18653,N_18461,N_18433);
nand U18654 (N_18654,N_18465,N_18502);
xnor U18655 (N_18655,N_18412,N_18533);
xor U18656 (N_18656,N_18493,N_18559);
nor U18657 (N_18657,N_18475,N_18499);
xnor U18658 (N_18658,N_18500,N_18464);
nor U18659 (N_18659,N_18448,N_18467);
xor U18660 (N_18660,N_18505,N_18488);
nand U18661 (N_18661,N_18458,N_18477);
or U18662 (N_18662,N_18484,N_18509);
xnor U18663 (N_18663,N_18467,N_18557);
and U18664 (N_18664,N_18427,N_18457);
or U18665 (N_18665,N_18424,N_18445);
or U18666 (N_18666,N_18422,N_18518);
nand U18667 (N_18667,N_18489,N_18435);
or U18668 (N_18668,N_18547,N_18546);
and U18669 (N_18669,N_18427,N_18468);
or U18670 (N_18670,N_18445,N_18400);
or U18671 (N_18671,N_18489,N_18512);
or U18672 (N_18672,N_18412,N_18546);
and U18673 (N_18673,N_18523,N_18534);
nand U18674 (N_18674,N_18442,N_18425);
and U18675 (N_18675,N_18412,N_18540);
and U18676 (N_18676,N_18556,N_18539);
and U18677 (N_18677,N_18477,N_18507);
and U18678 (N_18678,N_18558,N_18419);
nor U18679 (N_18679,N_18475,N_18456);
or U18680 (N_18680,N_18459,N_18526);
and U18681 (N_18681,N_18439,N_18512);
nor U18682 (N_18682,N_18406,N_18490);
nor U18683 (N_18683,N_18517,N_18403);
nand U18684 (N_18684,N_18418,N_18477);
xor U18685 (N_18685,N_18474,N_18443);
nor U18686 (N_18686,N_18433,N_18555);
xor U18687 (N_18687,N_18466,N_18545);
and U18688 (N_18688,N_18439,N_18416);
nand U18689 (N_18689,N_18495,N_18510);
or U18690 (N_18690,N_18461,N_18418);
nor U18691 (N_18691,N_18414,N_18456);
nand U18692 (N_18692,N_18482,N_18460);
and U18693 (N_18693,N_18535,N_18520);
xnor U18694 (N_18694,N_18543,N_18516);
and U18695 (N_18695,N_18402,N_18555);
nand U18696 (N_18696,N_18481,N_18528);
xor U18697 (N_18697,N_18554,N_18508);
nand U18698 (N_18698,N_18462,N_18448);
xor U18699 (N_18699,N_18401,N_18419);
nor U18700 (N_18700,N_18429,N_18472);
and U18701 (N_18701,N_18408,N_18519);
nand U18702 (N_18702,N_18416,N_18510);
or U18703 (N_18703,N_18548,N_18467);
or U18704 (N_18704,N_18557,N_18525);
or U18705 (N_18705,N_18462,N_18402);
and U18706 (N_18706,N_18406,N_18473);
xnor U18707 (N_18707,N_18549,N_18552);
xor U18708 (N_18708,N_18480,N_18487);
or U18709 (N_18709,N_18482,N_18503);
nand U18710 (N_18710,N_18547,N_18414);
and U18711 (N_18711,N_18496,N_18470);
xor U18712 (N_18712,N_18555,N_18426);
and U18713 (N_18713,N_18553,N_18525);
nor U18714 (N_18714,N_18558,N_18556);
and U18715 (N_18715,N_18479,N_18476);
and U18716 (N_18716,N_18413,N_18441);
xor U18717 (N_18717,N_18533,N_18523);
or U18718 (N_18718,N_18417,N_18521);
or U18719 (N_18719,N_18511,N_18445);
and U18720 (N_18720,N_18573,N_18585);
nor U18721 (N_18721,N_18596,N_18646);
and U18722 (N_18722,N_18595,N_18659);
nor U18723 (N_18723,N_18614,N_18617);
xor U18724 (N_18724,N_18579,N_18578);
or U18725 (N_18725,N_18608,N_18640);
nor U18726 (N_18726,N_18615,N_18582);
nor U18727 (N_18727,N_18671,N_18677);
or U18728 (N_18728,N_18633,N_18672);
or U18729 (N_18729,N_18564,N_18717);
xnor U18730 (N_18730,N_18713,N_18632);
nor U18731 (N_18731,N_18652,N_18698);
xor U18732 (N_18732,N_18570,N_18618);
or U18733 (N_18733,N_18621,N_18651);
or U18734 (N_18734,N_18625,N_18636);
and U18735 (N_18735,N_18681,N_18690);
and U18736 (N_18736,N_18688,N_18656);
or U18737 (N_18737,N_18707,N_18624);
nor U18738 (N_18738,N_18580,N_18657);
or U18739 (N_18739,N_18601,N_18691);
nor U18740 (N_18740,N_18703,N_18712);
or U18741 (N_18741,N_18599,N_18562);
and U18742 (N_18742,N_18714,N_18612);
or U18743 (N_18743,N_18635,N_18631);
and U18744 (N_18744,N_18598,N_18620);
and U18745 (N_18745,N_18699,N_18686);
nand U18746 (N_18746,N_18600,N_18639);
nand U18747 (N_18747,N_18571,N_18708);
and U18748 (N_18748,N_18711,N_18692);
or U18749 (N_18749,N_18649,N_18650);
nand U18750 (N_18750,N_18648,N_18704);
nor U18751 (N_18751,N_18715,N_18643);
or U18752 (N_18752,N_18594,N_18687);
and U18753 (N_18753,N_18623,N_18576);
or U18754 (N_18754,N_18626,N_18697);
or U18755 (N_18755,N_18577,N_18683);
and U18756 (N_18756,N_18709,N_18622);
nor U18757 (N_18757,N_18700,N_18638);
or U18758 (N_18758,N_18675,N_18642);
and U18759 (N_18759,N_18563,N_18592);
nor U18760 (N_18760,N_18565,N_18678);
or U18761 (N_18761,N_18665,N_18607);
nand U18762 (N_18762,N_18566,N_18561);
nand U18763 (N_18763,N_18696,N_18574);
and U18764 (N_18764,N_18597,N_18705);
nor U18765 (N_18765,N_18706,N_18637);
or U18766 (N_18766,N_18567,N_18627);
xnor U18767 (N_18767,N_18611,N_18680);
and U18768 (N_18768,N_18644,N_18604);
nand U18769 (N_18769,N_18682,N_18716);
nor U18770 (N_18770,N_18629,N_18605);
and U18771 (N_18771,N_18662,N_18590);
nor U18772 (N_18772,N_18653,N_18606);
or U18773 (N_18773,N_18718,N_18654);
nor U18774 (N_18774,N_18581,N_18694);
nor U18775 (N_18775,N_18641,N_18695);
xor U18776 (N_18776,N_18668,N_18593);
or U18777 (N_18777,N_18584,N_18591);
nor U18778 (N_18778,N_18586,N_18689);
xnor U18779 (N_18779,N_18702,N_18588);
nand U18780 (N_18780,N_18669,N_18679);
and U18781 (N_18781,N_18670,N_18693);
and U18782 (N_18782,N_18701,N_18674);
xor U18783 (N_18783,N_18569,N_18613);
nor U18784 (N_18784,N_18610,N_18602);
nor U18785 (N_18785,N_18628,N_18673);
and U18786 (N_18786,N_18619,N_18603);
nor U18787 (N_18787,N_18589,N_18710);
xnor U18788 (N_18788,N_18587,N_18685);
and U18789 (N_18789,N_18560,N_18676);
nor U18790 (N_18790,N_18660,N_18575);
and U18791 (N_18791,N_18719,N_18568);
xor U18792 (N_18792,N_18609,N_18572);
nand U18793 (N_18793,N_18661,N_18634);
nand U18794 (N_18794,N_18667,N_18616);
nor U18795 (N_18795,N_18630,N_18655);
and U18796 (N_18796,N_18663,N_18647);
or U18797 (N_18797,N_18666,N_18645);
and U18798 (N_18798,N_18583,N_18684);
xor U18799 (N_18799,N_18658,N_18664);
xor U18800 (N_18800,N_18636,N_18684);
nor U18801 (N_18801,N_18695,N_18667);
xor U18802 (N_18802,N_18632,N_18690);
nor U18803 (N_18803,N_18689,N_18638);
and U18804 (N_18804,N_18657,N_18586);
nand U18805 (N_18805,N_18636,N_18583);
or U18806 (N_18806,N_18573,N_18616);
xnor U18807 (N_18807,N_18604,N_18625);
nor U18808 (N_18808,N_18648,N_18626);
and U18809 (N_18809,N_18615,N_18607);
xnor U18810 (N_18810,N_18679,N_18604);
and U18811 (N_18811,N_18561,N_18685);
nor U18812 (N_18812,N_18587,N_18711);
nor U18813 (N_18813,N_18667,N_18651);
and U18814 (N_18814,N_18602,N_18623);
and U18815 (N_18815,N_18700,N_18672);
nor U18816 (N_18816,N_18615,N_18645);
xnor U18817 (N_18817,N_18654,N_18615);
xor U18818 (N_18818,N_18705,N_18617);
or U18819 (N_18819,N_18574,N_18572);
or U18820 (N_18820,N_18624,N_18573);
nand U18821 (N_18821,N_18694,N_18630);
or U18822 (N_18822,N_18631,N_18680);
nand U18823 (N_18823,N_18648,N_18621);
and U18824 (N_18824,N_18650,N_18657);
or U18825 (N_18825,N_18613,N_18653);
xnor U18826 (N_18826,N_18637,N_18583);
nor U18827 (N_18827,N_18640,N_18592);
nand U18828 (N_18828,N_18585,N_18578);
nand U18829 (N_18829,N_18658,N_18615);
nor U18830 (N_18830,N_18638,N_18715);
xor U18831 (N_18831,N_18672,N_18566);
nor U18832 (N_18832,N_18690,N_18649);
and U18833 (N_18833,N_18596,N_18614);
xnor U18834 (N_18834,N_18564,N_18692);
nand U18835 (N_18835,N_18666,N_18572);
and U18836 (N_18836,N_18575,N_18593);
nand U18837 (N_18837,N_18616,N_18626);
nand U18838 (N_18838,N_18649,N_18708);
nand U18839 (N_18839,N_18610,N_18695);
or U18840 (N_18840,N_18675,N_18589);
xor U18841 (N_18841,N_18597,N_18619);
nor U18842 (N_18842,N_18619,N_18570);
and U18843 (N_18843,N_18643,N_18699);
nor U18844 (N_18844,N_18712,N_18642);
nand U18845 (N_18845,N_18631,N_18693);
and U18846 (N_18846,N_18713,N_18615);
xnor U18847 (N_18847,N_18591,N_18699);
or U18848 (N_18848,N_18691,N_18644);
nand U18849 (N_18849,N_18577,N_18561);
xor U18850 (N_18850,N_18641,N_18719);
nand U18851 (N_18851,N_18617,N_18607);
or U18852 (N_18852,N_18632,N_18665);
nor U18853 (N_18853,N_18585,N_18630);
nor U18854 (N_18854,N_18711,N_18704);
and U18855 (N_18855,N_18659,N_18633);
and U18856 (N_18856,N_18658,N_18567);
nand U18857 (N_18857,N_18699,N_18564);
nor U18858 (N_18858,N_18612,N_18592);
nand U18859 (N_18859,N_18576,N_18691);
nand U18860 (N_18860,N_18711,N_18644);
nor U18861 (N_18861,N_18712,N_18686);
or U18862 (N_18862,N_18602,N_18640);
xor U18863 (N_18863,N_18653,N_18702);
nand U18864 (N_18864,N_18686,N_18683);
and U18865 (N_18865,N_18569,N_18717);
nand U18866 (N_18866,N_18694,N_18597);
nand U18867 (N_18867,N_18582,N_18584);
xor U18868 (N_18868,N_18639,N_18679);
and U18869 (N_18869,N_18665,N_18663);
or U18870 (N_18870,N_18600,N_18666);
or U18871 (N_18871,N_18699,N_18672);
nor U18872 (N_18872,N_18617,N_18621);
nor U18873 (N_18873,N_18591,N_18589);
nand U18874 (N_18874,N_18599,N_18704);
nand U18875 (N_18875,N_18567,N_18660);
nor U18876 (N_18876,N_18633,N_18600);
and U18877 (N_18877,N_18651,N_18716);
or U18878 (N_18878,N_18587,N_18699);
nor U18879 (N_18879,N_18698,N_18564);
nand U18880 (N_18880,N_18854,N_18790);
nand U18881 (N_18881,N_18752,N_18745);
xnor U18882 (N_18882,N_18767,N_18763);
nand U18883 (N_18883,N_18769,N_18877);
or U18884 (N_18884,N_18783,N_18778);
or U18885 (N_18885,N_18787,N_18858);
xor U18886 (N_18886,N_18867,N_18824);
or U18887 (N_18887,N_18782,N_18733);
or U18888 (N_18888,N_18773,N_18802);
nand U18889 (N_18889,N_18764,N_18806);
and U18890 (N_18890,N_18766,N_18746);
xor U18891 (N_18891,N_18727,N_18846);
or U18892 (N_18892,N_18755,N_18871);
and U18893 (N_18893,N_18837,N_18736);
nand U18894 (N_18894,N_18774,N_18722);
and U18895 (N_18895,N_18723,N_18726);
and U18896 (N_18896,N_18855,N_18779);
nand U18897 (N_18897,N_18742,N_18798);
and U18898 (N_18898,N_18864,N_18724);
or U18899 (N_18899,N_18757,N_18804);
nand U18900 (N_18900,N_18777,N_18841);
xnor U18901 (N_18901,N_18720,N_18836);
nor U18902 (N_18902,N_18738,N_18730);
nor U18903 (N_18903,N_18868,N_18833);
xnor U18904 (N_18904,N_18795,N_18750);
and U18905 (N_18905,N_18827,N_18850);
or U18906 (N_18906,N_18849,N_18876);
xor U18907 (N_18907,N_18820,N_18812);
and U18908 (N_18908,N_18759,N_18878);
xnor U18909 (N_18909,N_18776,N_18843);
nor U18910 (N_18910,N_18744,N_18748);
and U18911 (N_18911,N_18751,N_18870);
or U18912 (N_18912,N_18873,N_18734);
nand U18913 (N_18913,N_18740,N_18771);
and U18914 (N_18914,N_18754,N_18851);
nor U18915 (N_18915,N_18753,N_18801);
xor U18916 (N_18916,N_18874,N_18791);
xor U18917 (N_18917,N_18770,N_18829);
xnor U18918 (N_18918,N_18799,N_18793);
nand U18919 (N_18919,N_18807,N_18866);
nor U18920 (N_18920,N_18853,N_18808);
nand U18921 (N_18921,N_18732,N_18844);
nor U18922 (N_18922,N_18784,N_18735);
and U18923 (N_18923,N_18859,N_18749);
nor U18924 (N_18924,N_18794,N_18819);
xor U18925 (N_18925,N_18842,N_18821);
nor U18926 (N_18926,N_18848,N_18743);
nor U18927 (N_18927,N_18813,N_18856);
nand U18928 (N_18928,N_18879,N_18765);
and U18929 (N_18929,N_18810,N_18869);
and U18930 (N_18930,N_18830,N_18756);
xnor U18931 (N_18931,N_18865,N_18863);
nand U18932 (N_18932,N_18805,N_18721);
or U18933 (N_18933,N_18861,N_18835);
and U18934 (N_18934,N_18729,N_18811);
and U18935 (N_18935,N_18741,N_18803);
xnor U18936 (N_18936,N_18831,N_18828);
nand U18937 (N_18937,N_18737,N_18760);
and U18938 (N_18938,N_18809,N_18762);
nand U18939 (N_18939,N_18818,N_18825);
and U18940 (N_18940,N_18775,N_18875);
or U18941 (N_18941,N_18822,N_18747);
xnor U18942 (N_18942,N_18789,N_18786);
nor U18943 (N_18943,N_18768,N_18772);
xnor U18944 (N_18944,N_18728,N_18781);
or U18945 (N_18945,N_18788,N_18832);
nand U18946 (N_18946,N_18796,N_18839);
nand U18947 (N_18947,N_18852,N_18840);
and U18948 (N_18948,N_18857,N_18838);
nor U18949 (N_18949,N_18872,N_18834);
xnor U18950 (N_18950,N_18797,N_18800);
and U18951 (N_18951,N_18862,N_18814);
xor U18952 (N_18952,N_18761,N_18739);
nor U18953 (N_18953,N_18780,N_18845);
and U18954 (N_18954,N_18758,N_18816);
xnor U18955 (N_18955,N_18826,N_18725);
and U18956 (N_18956,N_18731,N_18817);
nand U18957 (N_18957,N_18792,N_18860);
nor U18958 (N_18958,N_18815,N_18823);
or U18959 (N_18959,N_18785,N_18847);
nor U18960 (N_18960,N_18856,N_18849);
and U18961 (N_18961,N_18770,N_18754);
nor U18962 (N_18962,N_18727,N_18775);
and U18963 (N_18963,N_18854,N_18735);
nor U18964 (N_18964,N_18800,N_18877);
xor U18965 (N_18965,N_18752,N_18857);
or U18966 (N_18966,N_18873,N_18780);
and U18967 (N_18967,N_18725,N_18821);
nand U18968 (N_18968,N_18821,N_18780);
nand U18969 (N_18969,N_18741,N_18784);
nor U18970 (N_18970,N_18848,N_18829);
nand U18971 (N_18971,N_18846,N_18837);
nand U18972 (N_18972,N_18826,N_18863);
xor U18973 (N_18973,N_18857,N_18795);
nand U18974 (N_18974,N_18850,N_18840);
or U18975 (N_18975,N_18859,N_18819);
and U18976 (N_18976,N_18803,N_18744);
nor U18977 (N_18977,N_18851,N_18806);
and U18978 (N_18978,N_18799,N_18766);
and U18979 (N_18979,N_18766,N_18789);
xnor U18980 (N_18980,N_18847,N_18738);
nor U18981 (N_18981,N_18756,N_18776);
nand U18982 (N_18982,N_18867,N_18872);
or U18983 (N_18983,N_18726,N_18783);
and U18984 (N_18984,N_18730,N_18833);
or U18985 (N_18985,N_18732,N_18782);
or U18986 (N_18986,N_18782,N_18781);
nand U18987 (N_18987,N_18756,N_18735);
xor U18988 (N_18988,N_18736,N_18755);
xnor U18989 (N_18989,N_18840,N_18739);
nand U18990 (N_18990,N_18829,N_18740);
nand U18991 (N_18991,N_18732,N_18749);
nand U18992 (N_18992,N_18767,N_18776);
nand U18993 (N_18993,N_18812,N_18796);
nand U18994 (N_18994,N_18737,N_18807);
nand U18995 (N_18995,N_18828,N_18780);
nand U18996 (N_18996,N_18802,N_18738);
and U18997 (N_18997,N_18800,N_18737);
and U18998 (N_18998,N_18868,N_18720);
nand U18999 (N_18999,N_18828,N_18754);
nand U19000 (N_19000,N_18852,N_18867);
or U19001 (N_19001,N_18790,N_18762);
or U19002 (N_19002,N_18774,N_18829);
nor U19003 (N_19003,N_18727,N_18754);
nor U19004 (N_19004,N_18869,N_18777);
or U19005 (N_19005,N_18723,N_18829);
or U19006 (N_19006,N_18799,N_18742);
or U19007 (N_19007,N_18748,N_18793);
and U19008 (N_19008,N_18828,N_18776);
nand U19009 (N_19009,N_18863,N_18813);
nand U19010 (N_19010,N_18741,N_18744);
nor U19011 (N_19011,N_18721,N_18770);
or U19012 (N_19012,N_18746,N_18852);
and U19013 (N_19013,N_18803,N_18793);
or U19014 (N_19014,N_18846,N_18743);
nor U19015 (N_19015,N_18724,N_18759);
and U19016 (N_19016,N_18805,N_18825);
xnor U19017 (N_19017,N_18777,N_18871);
xor U19018 (N_19018,N_18832,N_18799);
or U19019 (N_19019,N_18783,N_18801);
and U19020 (N_19020,N_18848,N_18740);
and U19021 (N_19021,N_18791,N_18754);
nor U19022 (N_19022,N_18840,N_18835);
nor U19023 (N_19023,N_18749,N_18775);
nor U19024 (N_19024,N_18760,N_18824);
nor U19025 (N_19025,N_18768,N_18783);
and U19026 (N_19026,N_18824,N_18724);
nor U19027 (N_19027,N_18836,N_18862);
xor U19028 (N_19028,N_18729,N_18789);
xor U19029 (N_19029,N_18846,N_18802);
xor U19030 (N_19030,N_18793,N_18741);
nand U19031 (N_19031,N_18846,N_18870);
xnor U19032 (N_19032,N_18747,N_18859);
xor U19033 (N_19033,N_18853,N_18784);
and U19034 (N_19034,N_18838,N_18877);
nor U19035 (N_19035,N_18779,N_18748);
nor U19036 (N_19036,N_18738,N_18835);
nand U19037 (N_19037,N_18814,N_18844);
nand U19038 (N_19038,N_18735,N_18871);
or U19039 (N_19039,N_18813,N_18817);
nand U19040 (N_19040,N_18915,N_18947);
and U19041 (N_19041,N_18993,N_18889);
and U19042 (N_19042,N_18953,N_18934);
nand U19043 (N_19043,N_18978,N_18894);
nor U19044 (N_19044,N_19016,N_18961);
or U19045 (N_19045,N_18983,N_19018);
nand U19046 (N_19046,N_18922,N_18946);
or U19047 (N_19047,N_18986,N_19019);
or U19048 (N_19048,N_18899,N_19023);
xnor U19049 (N_19049,N_18919,N_18988);
and U19050 (N_19050,N_19009,N_18903);
or U19051 (N_19051,N_18966,N_18973);
or U19052 (N_19052,N_18900,N_18982);
nor U19053 (N_19053,N_18970,N_18932);
and U19054 (N_19054,N_18910,N_18976);
and U19055 (N_19055,N_18908,N_19029);
and U19056 (N_19056,N_18886,N_18942);
xnor U19057 (N_19057,N_18904,N_18995);
xnor U19058 (N_19058,N_18950,N_18989);
xnor U19059 (N_19059,N_18937,N_18911);
nand U19060 (N_19060,N_19003,N_19002);
nand U19061 (N_19061,N_18979,N_18999);
or U19062 (N_19062,N_18955,N_18985);
or U19063 (N_19063,N_18967,N_19021);
xnor U19064 (N_19064,N_18906,N_18883);
and U19065 (N_19065,N_18925,N_19011);
and U19066 (N_19066,N_18944,N_18981);
nor U19067 (N_19067,N_19006,N_19022);
nor U19068 (N_19068,N_18998,N_18948);
nand U19069 (N_19069,N_18939,N_18909);
and U19070 (N_19070,N_18994,N_18980);
nand U19071 (N_19071,N_19035,N_19036);
or U19072 (N_19072,N_18921,N_18969);
xor U19073 (N_19073,N_18987,N_18935);
and U19074 (N_19074,N_18931,N_18996);
or U19075 (N_19075,N_18974,N_18958);
or U19076 (N_19076,N_18963,N_18941);
nor U19077 (N_19077,N_18924,N_18896);
or U19078 (N_19078,N_19027,N_18972);
xor U19079 (N_19079,N_19025,N_18957);
and U19080 (N_19080,N_19033,N_19008);
xnor U19081 (N_19081,N_18907,N_18890);
or U19082 (N_19082,N_18895,N_18905);
and U19083 (N_19083,N_19034,N_18940);
and U19084 (N_19084,N_18949,N_19038);
xnor U19085 (N_19085,N_19001,N_19024);
or U19086 (N_19086,N_18920,N_18990);
nor U19087 (N_19087,N_18891,N_18898);
or U19088 (N_19088,N_18951,N_19017);
nand U19089 (N_19089,N_19032,N_19026);
xor U19090 (N_19090,N_19039,N_18930);
nor U19091 (N_19091,N_18952,N_18887);
and U19092 (N_19092,N_19012,N_18975);
nand U19093 (N_19093,N_18960,N_18897);
nand U19094 (N_19094,N_18926,N_19004);
nand U19095 (N_19095,N_18881,N_18892);
or U19096 (N_19096,N_18914,N_18971);
nor U19097 (N_19097,N_18945,N_19015);
nand U19098 (N_19098,N_18938,N_18933);
nand U19099 (N_19099,N_18928,N_18936);
nor U19100 (N_19100,N_19005,N_18916);
or U19101 (N_19101,N_18913,N_19037);
nand U19102 (N_19102,N_19031,N_19028);
xnor U19103 (N_19103,N_19020,N_18929);
nand U19104 (N_19104,N_18885,N_18962);
nor U19105 (N_19105,N_19014,N_18884);
and U19106 (N_19106,N_18901,N_18991);
and U19107 (N_19107,N_18997,N_18964);
and U19108 (N_19108,N_18954,N_18923);
or U19109 (N_19109,N_18968,N_19030);
nor U19110 (N_19110,N_18918,N_18882);
nand U19111 (N_19111,N_19000,N_18959);
or U19112 (N_19112,N_19013,N_18984);
and U19113 (N_19113,N_18992,N_18943);
and U19114 (N_19114,N_18927,N_18965);
and U19115 (N_19115,N_18977,N_19010);
nor U19116 (N_19116,N_18912,N_18956);
and U19117 (N_19117,N_19007,N_18888);
nand U19118 (N_19118,N_18902,N_18880);
nand U19119 (N_19119,N_18893,N_18917);
and U19120 (N_19120,N_18985,N_18994);
or U19121 (N_19121,N_18968,N_18904);
or U19122 (N_19122,N_18946,N_18889);
xor U19123 (N_19123,N_19031,N_19016);
xor U19124 (N_19124,N_18885,N_19007);
or U19125 (N_19125,N_19007,N_19021);
nor U19126 (N_19126,N_19009,N_19028);
nor U19127 (N_19127,N_18921,N_19013);
and U19128 (N_19128,N_18908,N_18970);
xor U19129 (N_19129,N_19035,N_18920);
xnor U19130 (N_19130,N_18909,N_18972);
xor U19131 (N_19131,N_18914,N_18964);
nand U19132 (N_19132,N_18940,N_18966);
nor U19133 (N_19133,N_19038,N_18974);
and U19134 (N_19134,N_19025,N_18923);
or U19135 (N_19135,N_18901,N_19026);
nor U19136 (N_19136,N_18972,N_18920);
nor U19137 (N_19137,N_19002,N_18933);
nor U19138 (N_19138,N_19012,N_19023);
nand U19139 (N_19139,N_18940,N_18898);
nand U19140 (N_19140,N_18954,N_19000);
nor U19141 (N_19141,N_19011,N_18910);
nor U19142 (N_19142,N_18963,N_18971);
nor U19143 (N_19143,N_19002,N_18999);
nand U19144 (N_19144,N_18970,N_19006);
nand U19145 (N_19145,N_18916,N_18967);
and U19146 (N_19146,N_18997,N_18950);
and U19147 (N_19147,N_18937,N_18951);
nand U19148 (N_19148,N_18885,N_18948);
and U19149 (N_19149,N_18970,N_18894);
xnor U19150 (N_19150,N_19010,N_18985);
nand U19151 (N_19151,N_18988,N_18933);
nand U19152 (N_19152,N_18965,N_18890);
nand U19153 (N_19153,N_18885,N_19030);
nand U19154 (N_19154,N_19002,N_19004);
xor U19155 (N_19155,N_18961,N_19012);
xnor U19156 (N_19156,N_18995,N_19014);
nand U19157 (N_19157,N_18972,N_18989);
and U19158 (N_19158,N_19038,N_18915);
xor U19159 (N_19159,N_18917,N_19037);
nand U19160 (N_19160,N_18919,N_18960);
nand U19161 (N_19161,N_18890,N_19002);
and U19162 (N_19162,N_18969,N_18893);
and U19163 (N_19163,N_18977,N_18940);
and U19164 (N_19164,N_18894,N_19030);
nand U19165 (N_19165,N_19021,N_18965);
nor U19166 (N_19166,N_18905,N_18938);
nand U19167 (N_19167,N_19032,N_19031);
nand U19168 (N_19168,N_19037,N_19006);
nor U19169 (N_19169,N_18979,N_18967);
or U19170 (N_19170,N_18959,N_18914);
nor U19171 (N_19171,N_19033,N_18952);
and U19172 (N_19172,N_18983,N_18907);
or U19173 (N_19173,N_18997,N_19013);
and U19174 (N_19174,N_19002,N_18906);
or U19175 (N_19175,N_18941,N_18971);
nand U19176 (N_19176,N_18958,N_19030);
and U19177 (N_19177,N_18903,N_19014);
xor U19178 (N_19178,N_19012,N_18941);
nor U19179 (N_19179,N_18947,N_19037);
nor U19180 (N_19180,N_18953,N_18986);
xor U19181 (N_19181,N_18911,N_18892);
or U19182 (N_19182,N_18979,N_18968);
nor U19183 (N_19183,N_18988,N_18889);
or U19184 (N_19184,N_18939,N_18916);
nand U19185 (N_19185,N_18929,N_18990);
and U19186 (N_19186,N_18931,N_18990);
or U19187 (N_19187,N_18893,N_18965);
or U19188 (N_19188,N_19036,N_18915);
xor U19189 (N_19189,N_18923,N_19007);
and U19190 (N_19190,N_18928,N_18912);
nand U19191 (N_19191,N_18972,N_19007);
nand U19192 (N_19192,N_18928,N_18965);
nor U19193 (N_19193,N_18914,N_18916);
and U19194 (N_19194,N_18884,N_18883);
nand U19195 (N_19195,N_18993,N_18938);
nor U19196 (N_19196,N_18884,N_18903);
nand U19197 (N_19197,N_19007,N_19037);
and U19198 (N_19198,N_19017,N_18981);
xor U19199 (N_19199,N_18961,N_18977);
nand U19200 (N_19200,N_19040,N_19100);
nor U19201 (N_19201,N_19113,N_19167);
nand U19202 (N_19202,N_19075,N_19140);
or U19203 (N_19203,N_19134,N_19122);
or U19204 (N_19204,N_19138,N_19068);
or U19205 (N_19205,N_19131,N_19045);
and U19206 (N_19206,N_19168,N_19149);
and U19207 (N_19207,N_19185,N_19159);
or U19208 (N_19208,N_19172,N_19106);
xor U19209 (N_19209,N_19057,N_19077);
nand U19210 (N_19210,N_19109,N_19071);
xnor U19211 (N_19211,N_19170,N_19189);
nor U19212 (N_19212,N_19067,N_19151);
xor U19213 (N_19213,N_19053,N_19090);
nand U19214 (N_19214,N_19184,N_19166);
or U19215 (N_19215,N_19093,N_19177);
and U19216 (N_19216,N_19187,N_19086);
nor U19217 (N_19217,N_19130,N_19146);
or U19218 (N_19218,N_19176,N_19137);
xor U19219 (N_19219,N_19144,N_19047);
nor U19220 (N_19220,N_19078,N_19043);
or U19221 (N_19221,N_19169,N_19120);
nor U19222 (N_19222,N_19193,N_19142);
or U19223 (N_19223,N_19083,N_19141);
and U19224 (N_19224,N_19054,N_19076);
and U19225 (N_19225,N_19059,N_19175);
xnor U19226 (N_19226,N_19183,N_19085);
and U19227 (N_19227,N_19095,N_19186);
xor U19228 (N_19228,N_19114,N_19139);
and U19229 (N_19229,N_19181,N_19048);
and U19230 (N_19230,N_19108,N_19060);
nor U19231 (N_19231,N_19165,N_19179);
xnor U19232 (N_19232,N_19042,N_19063);
xnor U19233 (N_19233,N_19133,N_19198);
xnor U19234 (N_19234,N_19056,N_19191);
or U19235 (N_19235,N_19121,N_19074);
nand U19236 (N_19236,N_19157,N_19164);
or U19237 (N_19237,N_19041,N_19194);
xor U19238 (N_19238,N_19088,N_19118);
and U19239 (N_19239,N_19143,N_19046);
nor U19240 (N_19240,N_19092,N_19123);
xnor U19241 (N_19241,N_19190,N_19069);
xnor U19242 (N_19242,N_19188,N_19080);
or U19243 (N_19243,N_19197,N_19104);
xnor U19244 (N_19244,N_19107,N_19097);
nor U19245 (N_19245,N_19150,N_19135);
nand U19246 (N_19246,N_19119,N_19136);
nand U19247 (N_19247,N_19082,N_19062);
or U19248 (N_19248,N_19148,N_19128);
xor U19249 (N_19249,N_19084,N_19125);
or U19250 (N_19250,N_19091,N_19072);
and U19251 (N_19251,N_19099,N_19098);
xnor U19252 (N_19252,N_19180,N_19126);
or U19253 (N_19253,N_19055,N_19105);
nor U19254 (N_19254,N_19089,N_19160);
xor U19255 (N_19255,N_19155,N_19154);
and U19256 (N_19256,N_19182,N_19110);
or U19257 (N_19257,N_19070,N_19049);
and U19258 (N_19258,N_19163,N_19058);
or U19259 (N_19259,N_19147,N_19073);
nand U19260 (N_19260,N_19102,N_19124);
xor U19261 (N_19261,N_19096,N_19195);
and U19262 (N_19262,N_19153,N_19152);
or U19263 (N_19263,N_19129,N_19145);
or U19264 (N_19264,N_19101,N_19052);
nand U19265 (N_19265,N_19103,N_19111);
nand U19266 (N_19266,N_19192,N_19112);
xnor U19267 (N_19267,N_19044,N_19116);
nor U19268 (N_19268,N_19094,N_19065);
nand U19269 (N_19269,N_19174,N_19132);
nand U19270 (N_19270,N_19199,N_19079);
xor U19271 (N_19271,N_19061,N_19050);
xor U19272 (N_19272,N_19171,N_19156);
nand U19273 (N_19273,N_19196,N_19066);
nor U19274 (N_19274,N_19127,N_19064);
and U19275 (N_19275,N_19158,N_19087);
xor U19276 (N_19276,N_19173,N_19178);
nor U19277 (N_19277,N_19051,N_19081);
nand U19278 (N_19278,N_19117,N_19115);
or U19279 (N_19279,N_19162,N_19161);
nand U19280 (N_19280,N_19076,N_19192);
xor U19281 (N_19281,N_19048,N_19094);
nand U19282 (N_19282,N_19064,N_19128);
and U19283 (N_19283,N_19166,N_19068);
nor U19284 (N_19284,N_19105,N_19076);
nor U19285 (N_19285,N_19124,N_19108);
or U19286 (N_19286,N_19122,N_19194);
nand U19287 (N_19287,N_19185,N_19115);
nand U19288 (N_19288,N_19111,N_19074);
nor U19289 (N_19289,N_19081,N_19063);
or U19290 (N_19290,N_19047,N_19145);
nor U19291 (N_19291,N_19162,N_19071);
xor U19292 (N_19292,N_19132,N_19078);
nor U19293 (N_19293,N_19150,N_19095);
nand U19294 (N_19294,N_19152,N_19103);
xor U19295 (N_19295,N_19063,N_19071);
or U19296 (N_19296,N_19194,N_19165);
and U19297 (N_19297,N_19165,N_19055);
and U19298 (N_19298,N_19120,N_19050);
and U19299 (N_19299,N_19144,N_19043);
nor U19300 (N_19300,N_19189,N_19043);
nand U19301 (N_19301,N_19171,N_19133);
xnor U19302 (N_19302,N_19110,N_19085);
xnor U19303 (N_19303,N_19056,N_19071);
and U19304 (N_19304,N_19169,N_19186);
nand U19305 (N_19305,N_19156,N_19041);
nor U19306 (N_19306,N_19156,N_19194);
nand U19307 (N_19307,N_19116,N_19140);
nand U19308 (N_19308,N_19117,N_19175);
or U19309 (N_19309,N_19116,N_19148);
xor U19310 (N_19310,N_19074,N_19041);
nor U19311 (N_19311,N_19182,N_19078);
and U19312 (N_19312,N_19141,N_19171);
or U19313 (N_19313,N_19112,N_19183);
and U19314 (N_19314,N_19139,N_19095);
nand U19315 (N_19315,N_19154,N_19167);
xnor U19316 (N_19316,N_19080,N_19099);
nand U19317 (N_19317,N_19050,N_19066);
xor U19318 (N_19318,N_19084,N_19057);
xnor U19319 (N_19319,N_19158,N_19195);
or U19320 (N_19320,N_19161,N_19085);
or U19321 (N_19321,N_19055,N_19138);
xnor U19322 (N_19322,N_19071,N_19131);
and U19323 (N_19323,N_19162,N_19122);
xnor U19324 (N_19324,N_19070,N_19048);
xor U19325 (N_19325,N_19131,N_19134);
nand U19326 (N_19326,N_19044,N_19167);
nand U19327 (N_19327,N_19097,N_19149);
xnor U19328 (N_19328,N_19167,N_19156);
nand U19329 (N_19329,N_19052,N_19176);
xor U19330 (N_19330,N_19195,N_19191);
nor U19331 (N_19331,N_19184,N_19195);
nor U19332 (N_19332,N_19159,N_19178);
nor U19333 (N_19333,N_19177,N_19074);
and U19334 (N_19334,N_19067,N_19068);
or U19335 (N_19335,N_19185,N_19094);
xor U19336 (N_19336,N_19116,N_19076);
xnor U19337 (N_19337,N_19146,N_19115);
nand U19338 (N_19338,N_19122,N_19177);
nor U19339 (N_19339,N_19129,N_19118);
or U19340 (N_19340,N_19061,N_19073);
xnor U19341 (N_19341,N_19101,N_19051);
nand U19342 (N_19342,N_19051,N_19103);
nand U19343 (N_19343,N_19065,N_19190);
nand U19344 (N_19344,N_19116,N_19061);
or U19345 (N_19345,N_19179,N_19071);
nor U19346 (N_19346,N_19152,N_19140);
or U19347 (N_19347,N_19116,N_19193);
and U19348 (N_19348,N_19051,N_19040);
xnor U19349 (N_19349,N_19128,N_19171);
and U19350 (N_19350,N_19086,N_19113);
nor U19351 (N_19351,N_19150,N_19054);
nor U19352 (N_19352,N_19063,N_19172);
and U19353 (N_19353,N_19175,N_19173);
and U19354 (N_19354,N_19129,N_19070);
xor U19355 (N_19355,N_19190,N_19090);
nor U19356 (N_19356,N_19162,N_19127);
and U19357 (N_19357,N_19160,N_19161);
or U19358 (N_19358,N_19100,N_19130);
nand U19359 (N_19359,N_19098,N_19050);
nor U19360 (N_19360,N_19333,N_19226);
xor U19361 (N_19361,N_19263,N_19326);
xnor U19362 (N_19362,N_19331,N_19337);
xnor U19363 (N_19363,N_19327,N_19213);
and U19364 (N_19364,N_19211,N_19217);
nand U19365 (N_19365,N_19275,N_19303);
nand U19366 (N_19366,N_19352,N_19249);
and U19367 (N_19367,N_19339,N_19235);
nand U19368 (N_19368,N_19287,N_19247);
and U19369 (N_19369,N_19265,N_19210);
and U19370 (N_19370,N_19222,N_19223);
nor U19371 (N_19371,N_19207,N_19302);
xnor U19372 (N_19372,N_19301,N_19271);
xnor U19373 (N_19373,N_19291,N_19262);
or U19374 (N_19374,N_19237,N_19205);
and U19375 (N_19375,N_19225,N_19330);
or U19376 (N_19376,N_19351,N_19261);
and U19377 (N_19377,N_19289,N_19215);
and U19378 (N_19378,N_19206,N_19208);
and U19379 (N_19379,N_19346,N_19347);
or U19380 (N_19380,N_19338,N_19267);
or U19381 (N_19381,N_19232,N_19266);
nor U19382 (N_19382,N_19281,N_19345);
and U19383 (N_19383,N_19328,N_19341);
nand U19384 (N_19384,N_19293,N_19309);
or U19385 (N_19385,N_19238,N_19220);
xor U19386 (N_19386,N_19348,N_19343);
nor U19387 (N_19387,N_19231,N_19219);
or U19388 (N_19388,N_19254,N_19274);
nand U19389 (N_19389,N_19251,N_19212);
or U19390 (N_19390,N_19290,N_19294);
nor U19391 (N_19391,N_19240,N_19233);
and U19392 (N_19392,N_19342,N_19243);
nor U19393 (N_19393,N_19257,N_19307);
nand U19394 (N_19394,N_19319,N_19221);
nand U19395 (N_19395,N_19277,N_19284);
nor U19396 (N_19396,N_19276,N_19236);
xnor U19397 (N_19397,N_19256,N_19259);
nand U19398 (N_19398,N_19248,N_19355);
nor U19399 (N_19399,N_19313,N_19269);
nor U19400 (N_19400,N_19264,N_19308);
nand U19401 (N_19401,N_19353,N_19286);
nor U19402 (N_19402,N_19258,N_19298);
and U19403 (N_19403,N_19239,N_19332);
nor U19404 (N_19404,N_19321,N_19255);
and U19405 (N_19405,N_19200,N_19273);
and U19406 (N_19406,N_19203,N_19299);
or U19407 (N_19407,N_19296,N_19316);
xnor U19408 (N_19408,N_19329,N_19317);
or U19409 (N_19409,N_19312,N_19204);
and U19410 (N_19410,N_19268,N_19280);
nor U19411 (N_19411,N_19202,N_19246);
nor U19412 (N_19412,N_19357,N_19310);
and U19413 (N_19413,N_19209,N_19272);
or U19414 (N_19414,N_19201,N_19349);
nand U19415 (N_19415,N_19283,N_19334);
xnor U19416 (N_19416,N_19336,N_19324);
xor U19417 (N_19417,N_19358,N_19228);
nand U19418 (N_19418,N_19335,N_19241);
xnor U19419 (N_19419,N_19359,N_19216);
nand U19420 (N_19420,N_19305,N_19253);
or U19421 (N_19421,N_19323,N_19344);
and U19422 (N_19422,N_19315,N_19295);
nor U19423 (N_19423,N_19260,N_19320);
nor U19424 (N_19424,N_19229,N_19356);
and U19425 (N_19425,N_19270,N_19292);
or U19426 (N_19426,N_19245,N_19325);
xor U19427 (N_19427,N_19244,N_19288);
nor U19428 (N_19428,N_19230,N_19224);
xnor U19429 (N_19429,N_19279,N_19227);
and U19430 (N_19430,N_19306,N_19311);
or U19431 (N_19431,N_19285,N_19340);
or U19432 (N_19432,N_19350,N_19314);
nand U19433 (N_19433,N_19300,N_19234);
and U19434 (N_19434,N_19297,N_19354);
nor U19435 (N_19435,N_19214,N_19318);
nand U19436 (N_19436,N_19218,N_19322);
or U19437 (N_19437,N_19242,N_19282);
and U19438 (N_19438,N_19252,N_19304);
and U19439 (N_19439,N_19278,N_19250);
nand U19440 (N_19440,N_19310,N_19307);
or U19441 (N_19441,N_19270,N_19326);
nand U19442 (N_19442,N_19306,N_19252);
and U19443 (N_19443,N_19242,N_19257);
or U19444 (N_19444,N_19328,N_19315);
xor U19445 (N_19445,N_19260,N_19296);
or U19446 (N_19446,N_19312,N_19229);
xnor U19447 (N_19447,N_19356,N_19219);
nor U19448 (N_19448,N_19229,N_19347);
xnor U19449 (N_19449,N_19359,N_19243);
nor U19450 (N_19450,N_19283,N_19324);
nor U19451 (N_19451,N_19261,N_19258);
xnor U19452 (N_19452,N_19211,N_19254);
nor U19453 (N_19453,N_19323,N_19319);
xor U19454 (N_19454,N_19357,N_19233);
xnor U19455 (N_19455,N_19351,N_19343);
and U19456 (N_19456,N_19305,N_19205);
or U19457 (N_19457,N_19219,N_19224);
nor U19458 (N_19458,N_19204,N_19314);
nor U19459 (N_19459,N_19276,N_19315);
and U19460 (N_19460,N_19332,N_19229);
xor U19461 (N_19461,N_19308,N_19204);
nand U19462 (N_19462,N_19328,N_19202);
xnor U19463 (N_19463,N_19254,N_19250);
nor U19464 (N_19464,N_19356,N_19288);
nand U19465 (N_19465,N_19312,N_19249);
or U19466 (N_19466,N_19329,N_19324);
or U19467 (N_19467,N_19349,N_19261);
nor U19468 (N_19468,N_19252,N_19315);
and U19469 (N_19469,N_19225,N_19239);
nand U19470 (N_19470,N_19235,N_19317);
nor U19471 (N_19471,N_19227,N_19212);
nor U19472 (N_19472,N_19230,N_19241);
nor U19473 (N_19473,N_19213,N_19267);
nor U19474 (N_19474,N_19211,N_19338);
nor U19475 (N_19475,N_19220,N_19233);
nor U19476 (N_19476,N_19340,N_19224);
nor U19477 (N_19477,N_19320,N_19328);
and U19478 (N_19478,N_19265,N_19231);
nor U19479 (N_19479,N_19254,N_19358);
xor U19480 (N_19480,N_19344,N_19303);
nor U19481 (N_19481,N_19301,N_19308);
nand U19482 (N_19482,N_19282,N_19230);
or U19483 (N_19483,N_19295,N_19343);
or U19484 (N_19484,N_19343,N_19291);
nor U19485 (N_19485,N_19229,N_19355);
and U19486 (N_19486,N_19331,N_19218);
or U19487 (N_19487,N_19331,N_19234);
or U19488 (N_19488,N_19242,N_19226);
xor U19489 (N_19489,N_19264,N_19356);
nand U19490 (N_19490,N_19292,N_19349);
nor U19491 (N_19491,N_19256,N_19218);
nor U19492 (N_19492,N_19264,N_19316);
and U19493 (N_19493,N_19321,N_19211);
nand U19494 (N_19494,N_19239,N_19220);
nand U19495 (N_19495,N_19295,N_19218);
nor U19496 (N_19496,N_19230,N_19345);
xnor U19497 (N_19497,N_19332,N_19303);
nand U19498 (N_19498,N_19222,N_19255);
or U19499 (N_19499,N_19331,N_19247);
or U19500 (N_19500,N_19232,N_19288);
nor U19501 (N_19501,N_19258,N_19349);
xor U19502 (N_19502,N_19283,N_19274);
nand U19503 (N_19503,N_19317,N_19314);
nor U19504 (N_19504,N_19290,N_19309);
or U19505 (N_19505,N_19285,N_19289);
or U19506 (N_19506,N_19333,N_19275);
xnor U19507 (N_19507,N_19260,N_19300);
nand U19508 (N_19508,N_19307,N_19295);
xor U19509 (N_19509,N_19318,N_19312);
xnor U19510 (N_19510,N_19288,N_19315);
nand U19511 (N_19511,N_19274,N_19300);
nor U19512 (N_19512,N_19337,N_19218);
and U19513 (N_19513,N_19204,N_19281);
nor U19514 (N_19514,N_19277,N_19350);
nand U19515 (N_19515,N_19325,N_19252);
or U19516 (N_19516,N_19357,N_19218);
or U19517 (N_19517,N_19338,N_19283);
and U19518 (N_19518,N_19310,N_19305);
or U19519 (N_19519,N_19261,N_19295);
xnor U19520 (N_19520,N_19400,N_19434);
nor U19521 (N_19521,N_19399,N_19392);
nand U19522 (N_19522,N_19456,N_19386);
nor U19523 (N_19523,N_19367,N_19489);
or U19524 (N_19524,N_19490,N_19409);
nand U19525 (N_19525,N_19424,N_19498);
and U19526 (N_19526,N_19503,N_19439);
nor U19527 (N_19527,N_19485,N_19425);
nand U19528 (N_19528,N_19492,N_19507);
or U19529 (N_19529,N_19417,N_19517);
nand U19530 (N_19530,N_19366,N_19422);
xnor U19531 (N_19531,N_19370,N_19446);
and U19532 (N_19532,N_19463,N_19478);
and U19533 (N_19533,N_19459,N_19379);
nand U19534 (N_19534,N_19437,N_19482);
nand U19535 (N_19535,N_19426,N_19442);
or U19536 (N_19536,N_19472,N_19419);
or U19537 (N_19537,N_19408,N_19451);
nand U19538 (N_19538,N_19362,N_19511);
nor U19539 (N_19539,N_19509,N_19397);
nand U19540 (N_19540,N_19469,N_19404);
or U19541 (N_19541,N_19372,N_19443);
nor U19542 (N_19542,N_19371,N_19480);
xor U19543 (N_19543,N_19506,N_19468);
nor U19544 (N_19544,N_19410,N_19405);
or U19545 (N_19545,N_19368,N_19365);
nand U19546 (N_19546,N_19501,N_19448);
or U19547 (N_19547,N_19364,N_19487);
xnor U19548 (N_19548,N_19402,N_19374);
and U19549 (N_19549,N_19396,N_19514);
xor U19550 (N_19550,N_19475,N_19470);
xor U19551 (N_19551,N_19383,N_19429);
and U19552 (N_19552,N_19385,N_19418);
and U19553 (N_19553,N_19462,N_19497);
nor U19554 (N_19554,N_19412,N_19427);
nor U19555 (N_19555,N_19423,N_19416);
xor U19556 (N_19556,N_19414,N_19398);
or U19557 (N_19557,N_19465,N_19493);
xor U19558 (N_19558,N_19496,N_19441);
and U19559 (N_19559,N_19488,N_19458);
xor U19560 (N_19560,N_19403,N_19415);
or U19561 (N_19561,N_19373,N_19519);
nand U19562 (N_19562,N_19432,N_19376);
xor U19563 (N_19563,N_19394,N_19411);
xor U19564 (N_19564,N_19483,N_19481);
or U19565 (N_19565,N_19430,N_19495);
or U19566 (N_19566,N_19395,N_19513);
nand U19567 (N_19567,N_19477,N_19460);
nor U19568 (N_19568,N_19389,N_19484);
and U19569 (N_19569,N_19510,N_19502);
nand U19570 (N_19570,N_19486,N_19491);
xor U19571 (N_19571,N_19406,N_19512);
xnor U19572 (N_19572,N_19466,N_19420);
nand U19573 (N_19573,N_19438,N_19377);
xnor U19574 (N_19574,N_19381,N_19384);
xnor U19575 (N_19575,N_19382,N_19518);
or U19576 (N_19576,N_19457,N_19388);
nor U19577 (N_19577,N_19378,N_19361);
nand U19578 (N_19578,N_19391,N_19444);
nand U19579 (N_19579,N_19433,N_19504);
or U19580 (N_19580,N_19428,N_19369);
xnor U19581 (N_19581,N_19494,N_19516);
xnor U19582 (N_19582,N_19387,N_19499);
nor U19583 (N_19583,N_19452,N_19471);
xnor U19584 (N_19584,N_19407,N_19360);
nor U19585 (N_19585,N_19476,N_19467);
nand U19586 (N_19586,N_19508,N_19375);
and U19587 (N_19587,N_19473,N_19440);
nor U19588 (N_19588,N_19363,N_19455);
nor U19589 (N_19589,N_19500,N_19401);
and U19590 (N_19590,N_19454,N_19447);
nor U19591 (N_19591,N_19449,N_19479);
and U19592 (N_19592,N_19505,N_19461);
nand U19593 (N_19593,N_19515,N_19450);
nor U19594 (N_19594,N_19445,N_19436);
or U19595 (N_19595,N_19464,N_19413);
nand U19596 (N_19596,N_19380,N_19421);
nand U19597 (N_19597,N_19431,N_19474);
xor U19598 (N_19598,N_19435,N_19390);
xnor U19599 (N_19599,N_19393,N_19453);
nor U19600 (N_19600,N_19464,N_19371);
nor U19601 (N_19601,N_19495,N_19409);
or U19602 (N_19602,N_19454,N_19373);
or U19603 (N_19603,N_19435,N_19389);
or U19604 (N_19604,N_19452,N_19472);
nor U19605 (N_19605,N_19459,N_19482);
xor U19606 (N_19606,N_19444,N_19368);
nor U19607 (N_19607,N_19462,N_19466);
or U19608 (N_19608,N_19479,N_19426);
and U19609 (N_19609,N_19427,N_19391);
nand U19610 (N_19610,N_19434,N_19413);
xnor U19611 (N_19611,N_19519,N_19448);
and U19612 (N_19612,N_19473,N_19421);
or U19613 (N_19613,N_19385,N_19518);
or U19614 (N_19614,N_19374,N_19412);
xnor U19615 (N_19615,N_19391,N_19410);
nor U19616 (N_19616,N_19391,N_19429);
nand U19617 (N_19617,N_19472,N_19483);
nor U19618 (N_19618,N_19424,N_19510);
nand U19619 (N_19619,N_19410,N_19477);
and U19620 (N_19620,N_19475,N_19360);
or U19621 (N_19621,N_19426,N_19482);
nor U19622 (N_19622,N_19481,N_19510);
nor U19623 (N_19623,N_19485,N_19364);
nand U19624 (N_19624,N_19473,N_19436);
and U19625 (N_19625,N_19412,N_19415);
nor U19626 (N_19626,N_19491,N_19401);
nor U19627 (N_19627,N_19476,N_19413);
nand U19628 (N_19628,N_19483,N_19404);
xor U19629 (N_19629,N_19384,N_19500);
or U19630 (N_19630,N_19436,N_19371);
nand U19631 (N_19631,N_19464,N_19365);
or U19632 (N_19632,N_19474,N_19366);
xnor U19633 (N_19633,N_19364,N_19432);
xor U19634 (N_19634,N_19459,N_19477);
xor U19635 (N_19635,N_19498,N_19485);
xnor U19636 (N_19636,N_19369,N_19396);
or U19637 (N_19637,N_19370,N_19458);
nand U19638 (N_19638,N_19442,N_19486);
or U19639 (N_19639,N_19434,N_19510);
nand U19640 (N_19640,N_19379,N_19395);
and U19641 (N_19641,N_19437,N_19430);
nor U19642 (N_19642,N_19425,N_19426);
nor U19643 (N_19643,N_19516,N_19375);
nor U19644 (N_19644,N_19516,N_19461);
nand U19645 (N_19645,N_19405,N_19499);
xor U19646 (N_19646,N_19427,N_19404);
nor U19647 (N_19647,N_19390,N_19364);
nand U19648 (N_19648,N_19379,N_19494);
and U19649 (N_19649,N_19458,N_19447);
nand U19650 (N_19650,N_19456,N_19387);
xnor U19651 (N_19651,N_19445,N_19496);
nand U19652 (N_19652,N_19388,N_19484);
nor U19653 (N_19653,N_19492,N_19392);
nor U19654 (N_19654,N_19393,N_19502);
xor U19655 (N_19655,N_19411,N_19422);
nand U19656 (N_19656,N_19489,N_19490);
and U19657 (N_19657,N_19424,N_19434);
or U19658 (N_19658,N_19455,N_19423);
nor U19659 (N_19659,N_19500,N_19462);
or U19660 (N_19660,N_19426,N_19396);
nor U19661 (N_19661,N_19411,N_19496);
and U19662 (N_19662,N_19479,N_19474);
and U19663 (N_19663,N_19363,N_19513);
and U19664 (N_19664,N_19493,N_19518);
and U19665 (N_19665,N_19490,N_19482);
nand U19666 (N_19666,N_19480,N_19379);
nor U19667 (N_19667,N_19452,N_19385);
nor U19668 (N_19668,N_19409,N_19360);
nand U19669 (N_19669,N_19458,N_19361);
or U19670 (N_19670,N_19454,N_19365);
xor U19671 (N_19671,N_19397,N_19488);
xnor U19672 (N_19672,N_19506,N_19483);
and U19673 (N_19673,N_19373,N_19465);
xor U19674 (N_19674,N_19463,N_19392);
xnor U19675 (N_19675,N_19484,N_19433);
and U19676 (N_19676,N_19363,N_19386);
xnor U19677 (N_19677,N_19387,N_19429);
nand U19678 (N_19678,N_19392,N_19470);
nor U19679 (N_19679,N_19418,N_19372);
xnor U19680 (N_19680,N_19609,N_19642);
or U19681 (N_19681,N_19544,N_19570);
xnor U19682 (N_19682,N_19660,N_19628);
nand U19683 (N_19683,N_19526,N_19679);
xor U19684 (N_19684,N_19671,N_19614);
and U19685 (N_19685,N_19595,N_19550);
xnor U19686 (N_19686,N_19599,N_19635);
nand U19687 (N_19687,N_19649,N_19530);
or U19688 (N_19688,N_19668,N_19627);
xnor U19689 (N_19689,N_19541,N_19621);
and U19690 (N_19690,N_19670,N_19655);
or U19691 (N_19691,N_19563,N_19525);
or U19692 (N_19692,N_19528,N_19572);
nand U19693 (N_19693,N_19589,N_19584);
nor U19694 (N_19694,N_19669,N_19607);
xnor U19695 (N_19695,N_19556,N_19667);
nand U19696 (N_19696,N_19664,N_19587);
xor U19697 (N_19697,N_19551,N_19612);
nor U19698 (N_19698,N_19569,N_19663);
and U19699 (N_19699,N_19577,N_19610);
nor U19700 (N_19700,N_19547,N_19677);
xor U19701 (N_19701,N_19586,N_19552);
nand U19702 (N_19702,N_19558,N_19590);
and U19703 (N_19703,N_19532,N_19580);
and U19704 (N_19704,N_19553,N_19606);
xor U19705 (N_19705,N_19542,N_19651);
nor U19706 (N_19706,N_19529,N_19620);
or U19707 (N_19707,N_19576,N_19601);
and U19708 (N_19708,N_19625,N_19661);
nand U19709 (N_19709,N_19629,N_19571);
nor U19710 (N_19710,N_19593,N_19578);
nand U19711 (N_19711,N_19531,N_19662);
nor U19712 (N_19712,N_19656,N_19636);
xnor U19713 (N_19713,N_19592,N_19622);
nand U19714 (N_19714,N_19545,N_19568);
nor U19715 (N_19715,N_19643,N_19579);
or U19716 (N_19716,N_19658,N_19523);
nor U19717 (N_19717,N_19638,N_19646);
or U19718 (N_19718,N_19652,N_19549);
or U19719 (N_19719,N_19522,N_19666);
and U19720 (N_19720,N_19546,N_19650);
or U19721 (N_19721,N_19672,N_19539);
nand U19722 (N_19722,N_19555,N_19585);
nand U19723 (N_19723,N_19534,N_19600);
nor U19724 (N_19724,N_19557,N_19659);
or U19725 (N_19725,N_19560,N_19603);
and U19726 (N_19726,N_19535,N_19648);
xnor U19727 (N_19727,N_19597,N_19573);
xor U19728 (N_19728,N_19675,N_19634);
xnor U19729 (N_19729,N_19617,N_19561);
nor U19730 (N_19730,N_19653,N_19637);
nand U19731 (N_19731,N_19678,N_19524);
or U19732 (N_19732,N_19536,N_19582);
nor U19733 (N_19733,N_19567,N_19583);
nor U19734 (N_19734,N_19538,N_19543);
or U19735 (N_19735,N_19598,N_19574);
and U19736 (N_19736,N_19615,N_19613);
and U19737 (N_19737,N_19564,N_19611);
nand U19738 (N_19738,N_19644,N_19673);
and U19739 (N_19739,N_19565,N_19527);
xnor U19740 (N_19740,N_19631,N_19520);
nor U19741 (N_19741,N_19632,N_19676);
and U19742 (N_19742,N_19581,N_19559);
xnor U19743 (N_19743,N_19575,N_19605);
nand U19744 (N_19744,N_19596,N_19566);
xnor U19745 (N_19745,N_19647,N_19626);
or U19746 (N_19746,N_19616,N_19657);
nand U19747 (N_19747,N_19618,N_19540);
xor U19748 (N_19748,N_19665,N_19562);
xnor U19749 (N_19749,N_19588,N_19623);
nor U19750 (N_19750,N_19537,N_19533);
xor U19751 (N_19751,N_19674,N_19639);
or U19752 (N_19752,N_19641,N_19594);
and U19753 (N_19753,N_19548,N_19591);
and U19754 (N_19754,N_19554,N_19640);
nand U19755 (N_19755,N_19602,N_19608);
nand U19756 (N_19756,N_19633,N_19645);
and U19757 (N_19757,N_19654,N_19604);
or U19758 (N_19758,N_19521,N_19624);
and U19759 (N_19759,N_19619,N_19630);
xnor U19760 (N_19760,N_19589,N_19615);
and U19761 (N_19761,N_19640,N_19590);
xor U19762 (N_19762,N_19622,N_19565);
xnor U19763 (N_19763,N_19675,N_19628);
nor U19764 (N_19764,N_19656,N_19578);
and U19765 (N_19765,N_19608,N_19621);
nor U19766 (N_19766,N_19594,N_19602);
xor U19767 (N_19767,N_19575,N_19600);
and U19768 (N_19768,N_19666,N_19547);
and U19769 (N_19769,N_19643,N_19638);
nor U19770 (N_19770,N_19646,N_19658);
xor U19771 (N_19771,N_19590,N_19530);
xnor U19772 (N_19772,N_19617,N_19596);
nor U19773 (N_19773,N_19668,N_19522);
and U19774 (N_19774,N_19663,N_19556);
nand U19775 (N_19775,N_19522,N_19625);
or U19776 (N_19776,N_19627,N_19648);
nand U19777 (N_19777,N_19529,N_19520);
nor U19778 (N_19778,N_19657,N_19592);
nand U19779 (N_19779,N_19596,N_19616);
nand U19780 (N_19780,N_19618,N_19612);
xor U19781 (N_19781,N_19525,N_19605);
or U19782 (N_19782,N_19592,N_19569);
and U19783 (N_19783,N_19524,N_19590);
xor U19784 (N_19784,N_19561,N_19526);
or U19785 (N_19785,N_19659,N_19538);
xor U19786 (N_19786,N_19581,N_19641);
xnor U19787 (N_19787,N_19604,N_19665);
or U19788 (N_19788,N_19602,N_19626);
xor U19789 (N_19789,N_19578,N_19569);
or U19790 (N_19790,N_19671,N_19613);
or U19791 (N_19791,N_19588,N_19612);
and U19792 (N_19792,N_19609,N_19653);
and U19793 (N_19793,N_19673,N_19539);
or U19794 (N_19794,N_19628,N_19662);
nand U19795 (N_19795,N_19642,N_19649);
or U19796 (N_19796,N_19639,N_19600);
xor U19797 (N_19797,N_19555,N_19672);
nand U19798 (N_19798,N_19547,N_19679);
and U19799 (N_19799,N_19538,N_19530);
xor U19800 (N_19800,N_19662,N_19576);
and U19801 (N_19801,N_19594,N_19605);
nand U19802 (N_19802,N_19599,N_19669);
nor U19803 (N_19803,N_19544,N_19549);
and U19804 (N_19804,N_19591,N_19669);
xnor U19805 (N_19805,N_19539,N_19668);
or U19806 (N_19806,N_19598,N_19639);
xnor U19807 (N_19807,N_19543,N_19602);
or U19808 (N_19808,N_19654,N_19541);
xnor U19809 (N_19809,N_19662,N_19587);
nand U19810 (N_19810,N_19671,N_19622);
nand U19811 (N_19811,N_19521,N_19663);
xor U19812 (N_19812,N_19658,N_19675);
nor U19813 (N_19813,N_19677,N_19564);
nor U19814 (N_19814,N_19608,N_19539);
nor U19815 (N_19815,N_19623,N_19552);
nor U19816 (N_19816,N_19574,N_19625);
nor U19817 (N_19817,N_19524,N_19567);
nand U19818 (N_19818,N_19661,N_19613);
xor U19819 (N_19819,N_19584,N_19559);
xor U19820 (N_19820,N_19611,N_19620);
xnor U19821 (N_19821,N_19539,N_19549);
nor U19822 (N_19822,N_19636,N_19575);
nand U19823 (N_19823,N_19592,N_19526);
xnor U19824 (N_19824,N_19570,N_19524);
nor U19825 (N_19825,N_19594,N_19588);
xnor U19826 (N_19826,N_19535,N_19568);
xnor U19827 (N_19827,N_19637,N_19671);
xor U19828 (N_19828,N_19570,N_19637);
or U19829 (N_19829,N_19653,N_19596);
and U19830 (N_19830,N_19558,N_19583);
nand U19831 (N_19831,N_19609,N_19592);
and U19832 (N_19832,N_19556,N_19610);
and U19833 (N_19833,N_19662,N_19566);
xnor U19834 (N_19834,N_19564,N_19522);
nor U19835 (N_19835,N_19664,N_19636);
or U19836 (N_19836,N_19658,N_19547);
or U19837 (N_19837,N_19621,N_19635);
nor U19838 (N_19838,N_19654,N_19678);
xor U19839 (N_19839,N_19661,N_19566);
or U19840 (N_19840,N_19794,N_19692);
and U19841 (N_19841,N_19836,N_19693);
nand U19842 (N_19842,N_19830,N_19779);
xor U19843 (N_19843,N_19747,N_19742);
or U19844 (N_19844,N_19827,N_19732);
nor U19845 (N_19845,N_19785,N_19786);
xnor U19846 (N_19846,N_19758,N_19705);
nand U19847 (N_19847,N_19690,N_19807);
nand U19848 (N_19848,N_19755,N_19696);
nor U19849 (N_19849,N_19832,N_19804);
nand U19850 (N_19850,N_19806,N_19714);
and U19851 (N_19851,N_19756,N_19688);
nand U19852 (N_19852,N_19760,N_19740);
nor U19853 (N_19853,N_19774,N_19810);
nand U19854 (N_19854,N_19770,N_19728);
or U19855 (N_19855,N_19733,N_19710);
nand U19856 (N_19856,N_19695,N_19821);
or U19857 (N_19857,N_19788,N_19697);
xor U19858 (N_19858,N_19789,N_19777);
and U19859 (N_19859,N_19826,N_19684);
nor U19860 (N_19860,N_19701,N_19681);
xnor U19861 (N_19861,N_19752,N_19730);
xor U19862 (N_19862,N_19817,N_19716);
nand U19863 (N_19863,N_19795,N_19722);
xor U19864 (N_19864,N_19775,N_19725);
nand U19865 (N_19865,N_19825,N_19778);
nand U19866 (N_19866,N_19753,N_19745);
and U19867 (N_19867,N_19709,N_19796);
xnor U19868 (N_19868,N_19811,N_19797);
nor U19869 (N_19869,N_19707,N_19741);
and U19870 (N_19870,N_19835,N_19735);
xor U19871 (N_19871,N_19781,N_19833);
nor U19872 (N_19872,N_19720,N_19772);
nor U19873 (N_19873,N_19689,N_19746);
xor U19874 (N_19874,N_19766,N_19822);
nor U19875 (N_19875,N_19839,N_19762);
or U19876 (N_19876,N_19818,N_19736);
xor U19877 (N_19877,N_19837,N_19767);
xor U19878 (N_19878,N_19769,N_19738);
xnor U19879 (N_19879,N_19792,N_19829);
and U19880 (N_19880,N_19780,N_19704);
nand U19881 (N_19881,N_19803,N_19734);
and U19882 (N_19882,N_19721,N_19828);
nor U19883 (N_19883,N_19823,N_19703);
nor U19884 (N_19884,N_19683,N_19750);
nor U19885 (N_19885,N_19790,N_19754);
nand U19886 (N_19886,N_19751,N_19719);
and U19887 (N_19887,N_19686,N_19765);
and U19888 (N_19888,N_19798,N_19700);
or U19889 (N_19889,N_19706,N_19749);
or U19890 (N_19890,N_19791,N_19834);
xnor U19891 (N_19891,N_19727,N_19799);
and U19892 (N_19892,N_19812,N_19702);
nor U19893 (N_19893,N_19694,N_19711);
and U19894 (N_19894,N_19800,N_19699);
xor U19895 (N_19895,N_19713,N_19723);
and U19896 (N_19896,N_19712,N_19737);
nor U19897 (N_19897,N_19748,N_19813);
and U19898 (N_19898,N_19805,N_19717);
nand U19899 (N_19899,N_19744,N_19831);
nand U19900 (N_19900,N_19764,N_19682);
nand U19901 (N_19901,N_19757,N_19784);
or U19902 (N_19902,N_19708,N_19802);
nor U19903 (N_19903,N_19771,N_19814);
nor U19904 (N_19904,N_19763,N_19687);
nor U19905 (N_19905,N_19726,N_19724);
xor U19906 (N_19906,N_19782,N_19783);
and U19907 (N_19907,N_19808,N_19680);
and U19908 (N_19908,N_19838,N_19820);
or U19909 (N_19909,N_19739,N_19743);
nand U19910 (N_19910,N_19759,N_19801);
or U19911 (N_19911,N_19731,N_19815);
and U19912 (N_19912,N_19718,N_19776);
or U19913 (N_19913,N_19773,N_19816);
or U19914 (N_19914,N_19685,N_19715);
xnor U19915 (N_19915,N_19691,N_19793);
nand U19916 (N_19916,N_19768,N_19787);
and U19917 (N_19917,N_19819,N_19729);
xnor U19918 (N_19918,N_19824,N_19809);
and U19919 (N_19919,N_19761,N_19698);
xnor U19920 (N_19920,N_19725,N_19686);
nand U19921 (N_19921,N_19725,N_19705);
and U19922 (N_19922,N_19790,N_19682);
and U19923 (N_19923,N_19713,N_19773);
nor U19924 (N_19924,N_19796,N_19794);
nand U19925 (N_19925,N_19691,N_19833);
nand U19926 (N_19926,N_19700,N_19805);
or U19927 (N_19927,N_19727,N_19794);
or U19928 (N_19928,N_19740,N_19785);
xor U19929 (N_19929,N_19803,N_19837);
nand U19930 (N_19930,N_19835,N_19718);
nand U19931 (N_19931,N_19816,N_19799);
nand U19932 (N_19932,N_19720,N_19730);
nor U19933 (N_19933,N_19795,N_19784);
and U19934 (N_19934,N_19752,N_19828);
nand U19935 (N_19935,N_19833,N_19820);
xnor U19936 (N_19936,N_19695,N_19785);
or U19937 (N_19937,N_19831,N_19755);
xnor U19938 (N_19938,N_19761,N_19830);
nand U19939 (N_19939,N_19688,N_19711);
and U19940 (N_19940,N_19822,N_19765);
nand U19941 (N_19941,N_19697,N_19759);
nand U19942 (N_19942,N_19833,N_19729);
or U19943 (N_19943,N_19685,N_19719);
nor U19944 (N_19944,N_19770,N_19723);
and U19945 (N_19945,N_19752,N_19744);
and U19946 (N_19946,N_19748,N_19703);
or U19947 (N_19947,N_19742,N_19782);
or U19948 (N_19948,N_19785,N_19832);
or U19949 (N_19949,N_19734,N_19764);
nand U19950 (N_19950,N_19837,N_19799);
nor U19951 (N_19951,N_19804,N_19787);
and U19952 (N_19952,N_19766,N_19812);
xnor U19953 (N_19953,N_19740,N_19732);
xnor U19954 (N_19954,N_19801,N_19839);
and U19955 (N_19955,N_19742,N_19806);
or U19956 (N_19956,N_19763,N_19702);
nand U19957 (N_19957,N_19776,N_19826);
nand U19958 (N_19958,N_19721,N_19742);
nor U19959 (N_19959,N_19753,N_19803);
or U19960 (N_19960,N_19827,N_19770);
nor U19961 (N_19961,N_19741,N_19687);
nor U19962 (N_19962,N_19732,N_19708);
xor U19963 (N_19963,N_19735,N_19817);
and U19964 (N_19964,N_19741,N_19764);
nor U19965 (N_19965,N_19790,N_19809);
and U19966 (N_19966,N_19795,N_19701);
and U19967 (N_19967,N_19739,N_19708);
nand U19968 (N_19968,N_19831,N_19746);
or U19969 (N_19969,N_19714,N_19707);
nand U19970 (N_19970,N_19766,N_19680);
nor U19971 (N_19971,N_19770,N_19708);
nand U19972 (N_19972,N_19805,N_19799);
xnor U19973 (N_19973,N_19772,N_19795);
nor U19974 (N_19974,N_19818,N_19757);
nand U19975 (N_19975,N_19790,N_19804);
and U19976 (N_19976,N_19827,N_19733);
or U19977 (N_19977,N_19725,N_19763);
or U19978 (N_19978,N_19787,N_19775);
xor U19979 (N_19979,N_19726,N_19827);
nand U19980 (N_19980,N_19728,N_19692);
or U19981 (N_19981,N_19700,N_19762);
nor U19982 (N_19982,N_19830,N_19771);
nand U19983 (N_19983,N_19728,N_19805);
nand U19984 (N_19984,N_19696,N_19695);
nand U19985 (N_19985,N_19779,N_19827);
nor U19986 (N_19986,N_19760,N_19697);
or U19987 (N_19987,N_19695,N_19802);
or U19988 (N_19988,N_19817,N_19803);
nor U19989 (N_19989,N_19823,N_19735);
nor U19990 (N_19990,N_19830,N_19768);
and U19991 (N_19991,N_19701,N_19791);
xnor U19992 (N_19992,N_19835,N_19809);
nor U19993 (N_19993,N_19696,N_19828);
or U19994 (N_19994,N_19780,N_19720);
nor U19995 (N_19995,N_19709,N_19743);
xor U19996 (N_19996,N_19814,N_19718);
nand U19997 (N_19997,N_19810,N_19711);
and U19998 (N_19998,N_19710,N_19707);
or U19999 (N_19999,N_19720,N_19718);
nand UO_0 (O_0,N_19869,N_19948);
nor UO_1 (O_1,N_19879,N_19993);
nand UO_2 (O_2,N_19933,N_19911);
or UO_3 (O_3,N_19884,N_19921);
and UO_4 (O_4,N_19875,N_19864);
or UO_5 (O_5,N_19912,N_19891);
and UO_6 (O_6,N_19905,N_19913);
nand UO_7 (O_7,N_19997,N_19872);
or UO_8 (O_8,N_19925,N_19899);
nor UO_9 (O_9,N_19976,N_19845);
xor UO_10 (O_10,N_19862,N_19940);
or UO_11 (O_11,N_19980,N_19945);
or UO_12 (O_12,N_19907,N_19934);
xor UO_13 (O_13,N_19860,N_19944);
nor UO_14 (O_14,N_19906,N_19946);
xor UO_15 (O_15,N_19871,N_19932);
xnor UO_16 (O_16,N_19991,N_19842);
nor UO_17 (O_17,N_19920,N_19941);
xnor UO_18 (O_18,N_19959,N_19895);
nor UO_19 (O_19,N_19865,N_19967);
or UO_20 (O_20,N_19892,N_19840);
xor UO_21 (O_21,N_19953,N_19985);
or UO_22 (O_22,N_19977,N_19935);
or UO_23 (O_23,N_19988,N_19947);
nor UO_24 (O_24,N_19850,N_19973);
nand UO_25 (O_25,N_19958,N_19957);
nor UO_26 (O_26,N_19908,N_19928);
xor UO_27 (O_27,N_19999,N_19943);
or UO_28 (O_28,N_19852,N_19882);
or UO_29 (O_29,N_19883,N_19971);
or UO_30 (O_30,N_19962,N_19982);
xnor UO_31 (O_31,N_19969,N_19848);
nor UO_32 (O_32,N_19990,N_19847);
nor UO_33 (O_33,N_19964,N_19897);
or UO_34 (O_34,N_19841,N_19924);
and UO_35 (O_35,N_19878,N_19995);
xnor UO_36 (O_36,N_19868,N_19874);
nand UO_37 (O_37,N_19896,N_19952);
xor UO_38 (O_38,N_19877,N_19910);
or UO_39 (O_39,N_19949,N_19916);
or UO_40 (O_40,N_19979,N_19965);
xnor UO_41 (O_41,N_19901,N_19903);
xor UO_42 (O_42,N_19900,N_19972);
and UO_43 (O_43,N_19960,N_19849);
nand UO_44 (O_44,N_19996,N_19902);
xor UO_45 (O_45,N_19939,N_19954);
and UO_46 (O_46,N_19894,N_19986);
xnor UO_47 (O_47,N_19987,N_19956);
xnor UO_48 (O_48,N_19994,N_19927);
nor UO_49 (O_49,N_19863,N_19914);
or UO_50 (O_50,N_19930,N_19918);
nand UO_51 (O_51,N_19880,N_19861);
nor UO_52 (O_52,N_19978,N_19876);
xor UO_53 (O_53,N_19858,N_19981);
xnor UO_54 (O_54,N_19983,N_19881);
nand UO_55 (O_55,N_19857,N_19950);
and UO_56 (O_56,N_19856,N_19917);
and UO_57 (O_57,N_19955,N_19938);
or UO_58 (O_58,N_19904,N_19844);
nand UO_59 (O_59,N_19968,N_19888);
nand UO_60 (O_60,N_19889,N_19961);
xnor UO_61 (O_61,N_19998,N_19974);
or UO_62 (O_62,N_19887,N_19923);
nor UO_63 (O_63,N_19984,N_19885);
nor UO_64 (O_64,N_19922,N_19853);
nor UO_65 (O_65,N_19851,N_19929);
or UO_66 (O_66,N_19843,N_19886);
or UO_67 (O_67,N_19942,N_19846);
or UO_68 (O_68,N_19893,N_19951);
or UO_69 (O_69,N_19919,N_19989);
xnor UO_70 (O_70,N_19867,N_19926);
or UO_71 (O_71,N_19859,N_19963);
or UO_72 (O_72,N_19855,N_19890);
nor UO_73 (O_73,N_19909,N_19870);
xor UO_74 (O_74,N_19873,N_19975);
and UO_75 (O_75,N_19915,N_19992);
nand UO_76 (O_76,N_19854,N_19937);
or UO_77 (O_77,N_19936,N_19966);
and UO_78 (O_78,N_19931,N_19898);
xnor UO_79 (O_79,N_19970,N_19866);
nor UO_80 (O_80,N_19949,N_19952);
nor UO_81 (O_81,N_19920,N_19943);
nor UO_82 (O_82,N_19878,N_19869);
xor UO_83 (O_83,N_19882,N_19987);
or UO_84 (O_84,N_19900,N_19866);
nand UO_85 (O_85,N_19843,N_19917);
or UO_86 (O_86,N_19966,N_19991);
xor UO_87 (O_87,N_19986,N_19999);
and UO_88 (O_88,N_19900,N_19860);
nand UO_89 (O_89,N_19898,N_19897);
nor UO_90 (O_90,N_19846,N_19945);
or UO_91 (O_91,N_19999,N_19997);
or UO_92 (O_92,N_19931,N_19997);
nand UO_93 (O_93,N_19937,N_19972);
xor UO_94 (O_94,N_19883,N_19987);
xnor UO_95 (O_95,N_19864,N_19857);
and UO_96 (O_96,N_19946,N_19883);
or UO_97 (O_97,N_19903,N_19843);
and UO_98 (O_98,N_19899,N_19933);
or UO_99 (O_99,N_19915,N_19991);
nand UO_100 (O_100,N_19920,N_19979);
nand UO_101 (O_101,N_19869,N_19997);
and UO_102 (O_102,N_19870,N_19871);
and UO_103 (O_103,N_19973,N_19982);
and UO_104 (O_104,N_19998,N_19853);
or UO_105 (O_105,N_19997,N_19984);
xnor UO_106 (O_106,N_19862,N_19930);
and UO_107 (O_107,N_19986,N_19987);
or UO_108 (O_108,N_19988,N_19924);
nand UO_109 (O_109,N_19861,N_19995);
and UO_110 (O_110,N_19972,N_19925);
or UO_111 (O_111,N_19925,N_19889);
nor UO_112 (O_112,N_19935,N_19930);
xor UO_113 (O_113,N_19983,N_19965);
xor UO_114 (O_114,N_19921,N_19971);
nor UO_115 (O_115,N_19924,N_19914);
xor UO_116 (O_116,N_19987,N_19980);
xnor UO_117 (O_117,N_19943,N_19933);
nor UO_118 (O_118,N_19969,N_19930);
nor UO_119 (O_119,N_19878,N_19843);
nor UO_120 (O_120,N_19916,N_19938);
or UO_121 (O_121,N_19884,N_19984);
nor UO_122 (O_122,N_19881,N_19893);
or UO_123 (O_123,N_19981,N_19893);
and UO_124 (O_124,N_19933,N_19873);
and UO_125 (O_125,N_19898,N_19982);
nor UO_126 (O_126,N_19971,N_19969);
or UO_127 (O_127,N_19904,N_19855);
and UO_128 (O_128,N_19975,N_19869);
xor UO_129 (O_129,N_19871,N_19867);
nand UO_130 (O_130,N_19928,N_19941);
nand UO_131 (O_131,N_19846,N_19870);
or UO_132 (O_132,N_19951,N_19942);
nand UO_133 (O_133,N_19951,N_19918);
nor UO_134 (O_134,N_19998,N_19953);
xnor UO_135 (O_135,N_19998,N_19897);
nor UO_136 (O_136,N_19881,N_19888);
xor UO_137 (O_137,N_19940,N_19840);
nor UO_138 (O_138,N_19882,N_19982);
nor UO_139 (O_139,N_19917,N_19904);
nand UO_140 (O_140,N_19940,N_19904);
nor UO_141 (O_141,N_19917,N_19930);
and UO_142 (O_142,N_19966,N_19987);
or UO_143 (O_143,N_19944,N_19968);
nor UO_144 (O_144,N_19989,N_19903);
nand UO_145 (O_145,N_19924,N_19846);
or UO_146 (O_146,N_19910,N_19993);
and UO_147 (O_147,N_19881,N_19879);
and UO_148 (O_148,N_19857,N_19985);
nor UO_149 (O_149,N_19960,N_19902);
xor UO_150 (O_150,N_19910,N_19866);
nor UO_151 (O_151,N_19946,N_19852);
xnor UO_152 (O_152,N_19856,N_19888);
nand UO_153 (O_153,N_19841,N_19941);
and UO_154 (O_154,N_19898,N_19972);
nor UO_155 (O_155,N_19927,N_19971);
xor UO_156 (O_156,N_19952,N_19943);
xor UO_157 (O_157,N_19915,N_19843);
and UO_158 (O_158,N_19994,N_19919);
nand UO_159 (O_159,N_19870,N_19991);
xor UO_160 (O_160,N_19993,N_19855);
or UO_161 (O_161,N_19841,N_19986);
nor UO_162 (O_162,N_19991,N_19907);
or UO_163 (O_163,N_19912,N_19910);
or UO_164 (O_164,N_19996,N_19976);
nor UO_165 (O_165,N_19904,N_19865);
or UO_166 (O_166,N_19952,N_19951);
nand UO_167 (O_167,N_19942,N_19875);
xor UO_168 (O_168,N_19935,N_19939);
and UO_169 (O_169,N_19931,N_19924);
nand UO_170 (O_170,N_19932,N_19972);
xnor UO_171 (O_171,N_19894,N_19996);
nand UO_172 (O_172,N_19857,N_19956);
nor UO_173 (O_173,N_19901,N_19999);
and UO_174 (O_174,N_19950,N_19840);
nand UO_175 (O_175,N_19844,N_19857);
or UO_176 (O_176,N_19897,N_19940);
and UO_177 (O_177,N_19897,N_19860);
nor UO_178 (O_178,N_19991,N_19932);
or UO_179 (O_179,N_19868,N_19887);
or UO_180 (O_180,N_19960,N_19874);
nor UO_181 (O_181,N_19930,N_19909);
xnor UO_182 (O_182,N_19850,N_19896);
nand UO_183 (O_183,N_19850,N_19976);
nor UO_184 (O_184,N_19869,N_19957);
nand UO_185 (O_185,N_19906,N_19842);
nand UO_186 (O_186,N_19971,N_19854);
nand UO_187 (O_187,N_19843,N_19967);
nor UO_188 (O_188,N_19910,N_19944);
nand UO_189 (O_189,N_19920,N_19859);
or UO_190 (O_190,N_19854,N_19953);
nand UO_191 (O_191,N_19864,N_19989);
nand UO_192 (O_192,N_19977,N_19974);
or UO_193 (O_193,N_19866,N_19865);
nor UO_194 (O_194,N_19940,N_19914);
xnor UO_195 (O_195,N_19928,N_19997);
xor UO_196 (O_196,N_19859,N_19888);
nand UO_197 (O_197,N_19863,N_19956);
nand UO_198 (O_198,N_19922,N_19979);
nor UO_199 (O_199,N_19873,N_19875);
nor UO_200 (O_200,N_19984,N_19881);
xnor UO_201 (O_201,N_19872,N_19903);
and UO_202 (O_202,N_19878,N_19965);
xnor UO_203 (O_203,N_19997,N_19941);
or UO_204 (O_204,N_19934,N_19927);
xnor UO_205 (O_205,N_19869,N_19947);
nand UO_206 (O_206,N_19960,N_19933);
nor UO_207 (O_207,N_19979,N_19905);
xnor UO_208 (O_208,N_19911,N_19841);
xnor UO_209 (O_209,N_19911,N_19949);
nor UO_210 (O_210,N_19878,N_19901);
or UO_211 (O_211,N_19866,N_19877);
xor UO_212 (O_212,N_19861,N_19895);
nand UO_213 (O_213,N_19938,N_19868);
or UO_214 (O_214,N_19857,N_19951);
nand UO_215 (O_215,N_19995,N_19912);
nor UO_216 (O_216,N_19902,N_19853);
nand UO_217 (O_217,N_19844,N_19898);
nor UO_218 (O_218,N_19947,N_19881);
nor UO_219 (O_219,N_19875,N_19904);
xnor UO_220 (O_220,N_19870,N_19917);
and UO_221 (O_221,N_19840,N_19920);
or UO_222 (O_222,N_19948,N_19875);
or UO_223 (O_223,N_19848,N_19883);
nor UO_224 (O_224,N_19936,N_19924);
nor UO_225 (O_225,N_19969,N_19953);
nand UO_226 (O_226,N_19908,N_19965);
or UO_227 (O_227,N_19960,N_19963);
or UO_228 (O_228,N_19951,N_19993);
nor UO_229 (O_229,N_19911,N_19990);
xnor UO_230 (O_230,N_19966,N_19848);
and UO_231 (O_231,N_19931,N_19987);
or UO_232 (O_232,N_19906,N_19900);
nor UO_233 (O_233,N_19928,N_19846);
and UO_234 (O_234,N_19974,N_19851);
and UO_235 (O_235,N_19857,N_19899);
nor UO_236 (O_236,N_19885,N_19922);
nand UO_237 (O_237,N_19840,N_19842);
xnor UO_238 (O_238,N_19866,N_19884);
or UO_239 (O_239,N_19867,N_19891);
nand UO_240 (O_240,N_19942,N_19962);
nor UO_241 (O_241,N_19986,N_19844);
nand UO_242 (O_242,N_19911,N_19979);
or UO_243 (O_243,N_19929,N_19985);
or UO_244 (O_244,N_19923,N_19998);
or UO_245 (O_245,N_19913,N_19975);
nand UO_246 (O_246,N_19889,N_19964);
xor UO_247 (O_247,N_19909,N_19864);
or UO_248 (O_248,N_19844,N_19976);
nand UO_249 (O_249,N_19860,N_19980);
or UO_250 (O_250,N_19937,N_19945);
or UO_251 (O_251,N_19845,N_19841);
xnor UO_252 (O_252,N_19870,N_19916);
nor UO_253 (O_253,N_19963,N_19891);
or UO_254 (O_254,N_19911,N_19973);
xor UO_255 (O_255,N_19946,N_19880);
nor UO_256 (O_256,N_19907,N_19900);
nor UO_257 (O_257,N_19980,N_19918);
xor UO_258 (O_258,N_19905,N_19960);
and UO_259 (O_259,N_19930,N_19855);
nor UO_260 (O_260,N_19977,N_19932);
or UO_261 (O_261,N_19859,N_19981);
and UO_262 (O_262,N_19972,N_19902);
nor UO_263 (O_263,N_19956,N_19860);
nor UO_264 (O_264,N_19853,N_19904);
xnor UO_265 (O_265,N_19879,N_19874);
and UO_266 (O_266,N_19939,N_19878);
nand UO_267 (O_267,N_19972,N_19872);
and UO_268 (O_268,N_19880,N_19912);
or UO_269 (O_269,N_19950,N_19978);
nand UO_270 (O_270,N_19931,N_19890);
nand UO_271 (O_271,N_19990,N_19903);
nand UO_272 (O_272,N_19930,N_19846);
nor UO_273 (O_273,N_19983,N_19935);
xor UO_274 (O_274,N_19858,N_19849);
nand UO_275 (O_275,N_19902,N_19924);
nor UO_276 (O_276,N_19899,N_19843);
or UO_277 (O_277,N_19987,N_19988);
or UO_278 (O_278,N_19864,N_19886);
and UO_279 (O_279,N_19891,N_19970);
xor UO_280 (O_280,N_19952,N_19934);
nand UO_281 (O_281,N_19908,N_19857);
or UO_282 (O_282,N_19850,N_19860);
and UO_283 (O_283,N_19852,N_19870);
or UO_284 (O_284,N_19889,N_19953);
nand UO_285 (O_285,N_19918,N_19947);
xnor UO_286 (O_286,N_19922,N_19889);
and UO_287 (O_287,N_19900,N_19983);
nand UO_288 (O_288,N_19888,N_19905);
nand UO_289 (O_289,N_19994,N_19890);
nor UO_290 (O_290,N_19956,N_19988);
xor UO_291 (O_291,N_19969,N_19995);
xnor UO_292 (O_292,N_19924,N_19933);
and UO_293 (O_293,N_19932,N_19857);
nand UO_294 (O_294,N_19908,N_19979);
nand UO_295 (O_295,N_19913,N_19966);
nor UO_296 (O_296,N_19990,N_19893);
nor UO_297 (O_297,N_19841,N_19943);
nor UO_298 (O_298,N_19959,N_19884);
nor UO_299 (O_299,N_19981,N_19990);
nand UO_300 (O_300,N_19879,N_19975);
nor UO_301 (O_301,N_19896,N_19958);
or UO_302 (O_302,N_19912,N_19990);
nand UO_303 (O_303,N_19879,N_19969);
xnor UO_304 (O_304,N_19843,N_19857);
nor UO_305 (O_305,N_19979,N_19925);
or UO_306 (O_306,N_19969,N_19886);
nor UO_307 (O_307,N_19841,N_19931);
xnor UO_308 (O_308,N_19931,N_19985);
nor UO_309 (O_309,N_19926,N_19915);
xor UO_310 (O_310,N_19867,N_19878);
or UO_311 (O_311,N_19984,N_19861);
nand UO_312 (O_312,N_19883,N_19972);
nor UO_313 (O_313,N_19895,N_19949);
and UO_314 (O_314,N_19953,N_19982);
and UO_315 (O_315,N_19857,N_19926);
nor UO_316 (O_316,N_19979,N_19842);
nor UO_317 (O_317,N_19850,N_19878);
nand UO_318 (O_318,N_19877,N_19914);
xnor UO_319 (O_319,N_19980,N_19888);
nand UO_320 (O_320,N_19991,N_19919);
xor UO_321 (O_321,N_19941,N_19847);
or UO_322 (O_322,N_19986,N_19919);
xnor UO_323 (O_323,N_19897,N_19902);
or UO_324 (O_324,N_19948,N_19909);
xnor UO_325 (O_325,N_19927,N_19881);
nor UO_326 (O_326,N_19961,N_19953);
nor UO_327 (O_327,N_19965,N_19931);
xnor UO_328 (O_328,N_19897,N_19982);
nand UO_329 (O_329,N_19964,N_19965);
or UO_330 (O_330,N_19959,N_19955);
and UO_331 (O_331,N_19918,N_19945);
and UO_332 (O_332,N_19849,N_19879);
or UO_333 (O_333,N_19857,N_19927);
nand UO_334 (O_334,N_19905,N_19942);
nand UO_335 (O_335,N_19845,N_19994);
xnor UO_336 (O_336,N_19917,N_19968);
xnor UO_337 (O_337,N_19981,N_19863);
nor UO_338 (O_338,N_19945,N_19942);
or UO_339 (O_339,N_19924,N_19901);
or UO_340 (O_340,N_19909,N_19973);
nor UO_341 (O_341,N_19915,N_19940);
xnor UO_342 (O_342,N_19960,N_19978);
xor UO_343 (O_343,N_19937,N_19872);
or UO_344 (O_344,N_19913,N_19933);
nand UO_345 (O_345,N_19919,N_19949);
xor UO_346 (O_346,N_19852,N_19949);
xnor UO_347 (O_347,N_19878,N_19913);
and UO_348 (O_348,N_19891,N_19898);
and UO_349 (O_349,N_19892,N_19917);
and UO_350 (O_350,N_19997,N_19911);
or UO_351 (O_351,N_19948,N_19900);
xor UO_352 (O_352,N_19845,N_19897);
xor UO_353 (O_353,N_19918,N_19977);
and UO_354 (O_354,N_19934,N_19851);
nand UO_355 (O_355,N_19990,N_19937);
and UO_356 (O_356,N_19908,N_19877);
and UO_357 (O_357,N_19926,N_19963);
or UO_358 (O_358,N_19919,N_19960);
nand UO_359 (O_359,N_19973,N_19966);
and UO_360 (O_360,N_19866,N_19961);
or UO_361 (O_361,N_19913,N_19962);
nand UO_362 (O_362,N_19858,N_19938);
xnor UO_363 (O_363,N_19863,N_19978);
xor UO_364 (O_364,N_19971,N_19986);
and UO_365 (O_365,N_19925,N_19931);
or UO_366 (O_366,N_19842,N_19951);
or UO_367 (O_367,N_19958,N_19975);
and UO_368 (O_368,N_19880,N_19952);
nor UO_369 (O_369,N_19851,N_19874);
xor UO_370 (O_370,N_19912,N_19993);
and UO_371 (O_371,N_19942,N_19953);
nor UO_372 (O_372,N_19981,N_19876);
and UO_373 (O_373,N_19954,N_19941);
and UO_374 (O_374,N_19910,N_19977);
or UO_375 (O_375,N_19992,N_19965);
nor UO_376 (O_376,N_19860,N_19906);
or UO_377 (O_377,N_19992,N_19859);
and UO_378 (O_378,N_19991,N_19875);
nor UO_379 (O_379,N_19878,N_19873);
nand UO_380 (O_380,N_19934,N_19964);
or UO_381 (O_381,N_19847,N_19999);
nand UO_382 (O_382,N_19897,N_19931);
nor UO_383 (O_383,N_19995,N_19957);
xor UO_384 (O_384,N_19970,N_19864);
nand UO_385 (O_385,N_19928,N_19911);
and UO_386 (O_386,N_19891,N_19853);
nor UO_387 (O_387,N_19926,N_19914);
or UO_388 (O_388,N_19842,N_19878);
nor UO_389 (O_389,N_19910,N_19889);
nor UO_390 (O_390,N_19975,N_19911);
nand UO_391 (O_391,N_19924,N_19872);
and UO_392 (O_392,N_19850,N_19957);
nand UO_393 (O_393,N_19927,N_19952);
nand UO_394 (O_394,N_19950,N_19867);
and UO_395 (O_395,N_19905,N_19884);
xor UO_396 (O_396,N_19998,N_19921);
or UO_397 (O_397,N_19952,N_19907);
nand UO_398 (O_398,N_19953,N_19917);
nor UO_399 (O_399,N_19988,N_19929);
nand UO_400 (O_400,N_19894,N_19911);
nand UO_401 (O_401,N_19873,N_19984);
nor UO_402 (O_402,N_19961,N_19988);
or UO_403 (O_403,N_19878,N_19950);
or UO_404 (O_404,N_19862,N_19907);
or UO_405 (O_405,N_19889,N_19971);
and UO_406 (O_406,N_19900,N_19924);
nor UO_407 (O_407,N_19974,N_19870);
or UO_408 (O_408,N_19905,N_19958);
nor UO_409 (O_409,N_19933,N_19978);
nand UO_410 (O_410,N_19908,N_19937);
nand UO_411 (O_411,N_19924,N_19996);
nor UO_412 (O_412,N_19927,N_19958);
nand UO_413 (O_413,N_19873,N_19974);
nor UO_414 (O_414,N_19919,N_19934);
or UO_415 (O_415,N_19894,N_19944);
or UO_416 (O_416,N_19910,N_19968);
or UO_417 (O_417,N_19933,N_19849);
and UO_418 (O_418,N_19890,N_19851);
and UO_419 (O_419,N_19970,N_19907);
xor UO_420 (O_420,N_19899,N_19993);
nand UO_421 (O_421,N_19840,N_19988);
xnor UO_422 (O_422,N_19900,N_19844);
and UO_423 (O_423,N_19981,N_19849);
nand UO_424 (O_424,N_19856,N_19979);
xor UO_425 (O_425,N_19924,N_19911);
nand UO_426 (O_426,N_19876,N_19902);
xor UO_427 (O_427,N_19858,N_19962);
xnor UO_428 (O_428,N_19980,N_19964);
xor UO_429 (O_429,N_19919,N_19858);
nand UO_430 (O_430,N_19986,N_19888);
nand UO_431 (O_431,N_19918,N_19965);
xnor UO_432 (O_432,N_19884,N_19992);
nand UO_433 (O_433,N_19992,N_19916);
nand UO_434 (O_434,N_19887,N_19906);
or UO_435 (O_435,N_19872,N_19947);
or UO_436 (O_436,N_19948,N_19954);
nor UO_437 (O_437,N_19873,N_19967);
xnor UO_438 (O_438,N_19964,N_19935);
xor UO_439 (O_439,N_19923,N_19900);
or UO_440 (O_440,N_19923,N_19840);
and UO_441 (O_441,N_19977,N_19968);
nor UO_442 (O_442,N_19919,N_19935);
nand UO_443 (O_443,N_19891,N_19906);
and UO_444 (O_444,N_19926,N_19932);
or UO_445 (O_445,N_19927,N_19845);
xor UO_446 (O_446,N_19939,N_19882);
nor UO_447 (O_447,N_19911,N_19940);
or UO_448 (O_448,N_19976,N_19938);
or UO_449 (O_449,N_19944,N_19959);
nand UO_450 (O_450,N_19876,N_19853);
or UO_451 (O_451,N_19913,N_19902);
nor UO_452 (O_452,N_19964,N_19848);
xnor UO_453 (O_453,N_19970,N_19940);
and UO_454 (O_454,N_19943,N_19844);
nor UO_455 (O_455,N_19846,N_19933);
xor UO_456 (O_456,N_19922,N_19919);
xor UO_457 (O_457,N_19905,N_19898);
nand UO_458 (O_458,N_19970,N_19973);
xor UO_459 (O_459,N_19848,N_19938);
nor UO_460 (O_460,N_19861,N_19841);
xnor UO_461 (O_461,N_19945,N_19969);
nor UO_462 (O_462,N_19934,N_19944);
and UO_463 (O_463,N_19880,N_19927);
nand UO_464 (O_464,N_19939,N_19897);
nor UO_465 (O_465,N_19990,N_19989);
nor UO_466 (O_466,N_19849,N_19894);
xor UO_467 (O_467,N_19975,N_19969);
xor UO_468 (O_468,N_19953,N_19996);
xor UO_469 (O_469,N_19909,N_19854);
nor UO_470 (O_470,N_19907,N_19869);
nand UO_471 (O_471,N_19914,N_19891);
xor UO_472 (O_472,N_19943,N_19998);
nor UO_473 (O_473,N_19956,N_19924);
nand UO_474 (O_474,N_19976,N_19979);
nand UO_475 (O_475,N_19883,N_19905);
xnor UO_476 (O_476,N_19942,N_19956);
xor UO_477 (O_477,N_19855,N_19969);
or UO_478 (O_478,N_19991,N_19981);
nor UO_479 (O_479,N_19971,N_19956);
or UO_480 (O_480,N_19980,N_19968);
or UO_481 (O_481,N_19944,N_19943);
nand UO_482 (O_482,N_19945,N_19840);
and UO_483 (O_483,N_19916,N_19953);
nand UO_484 (O_484,N_19961,N_19847);
nand UO_485 (O_485,N_19862,N_19983);
nor UO_486 (O_486,N_19931,N_19920);
and UO_487 (O_487,N_19858,N_19959);
or UO_488 (O_488,N_19985,N_19973);
xor UO_489 (O_489,N_19926,N_19853);
nor UO_490 (O_490,N_19901,N_19943);
nand UO_491 (O_491,N_19965,N_19993);
nand UO_492 (O_492,N_19927,N_19956);
xnor UO_493 (O_493,N_19888,N_19866);
and UO_494 (O_494,N_19871,N_19915);
and UO_495 (O_495,N_19840,N_19876);
nor UO_496 (O_496,N_19861,N_19851);
and UO_497 (O_497,N_19975,N_19988);
or UO_498 (O_498,N_19939,N_19918);
nand UO_499 (O_499,N_19942,N_19887);
and UO_500 (O_500,N_19866,N_19967);
or UO_501 (O_501,N_19895,N_19939);
or UO_502 (O_502,N_19989,N_19893);
xnor UO_503 (O_503,N_19885,N_19959);
nor UO_504 (O_504,N_19935,N_19857);
xnor UO_505 (O_505,N_19845,N_19970);
xor UO_506 (O_506,N_19961,N_19865);
or UO_507 (O_507,N_19947,N_19984);
nor UO_508 (O_508,N_19956,N_19913);
nor UO_509 (O_509,N_19844,N_19963);
and UO_510 (O_510,N_19844,N_19969);
xnor UO_511 (O_511,N_19908,N_19936);
or UO_512 (O_512,N_19849,N_19996);
nor UO_513 (O_513,N_19916,N_19964);
nor UO_514 (O_514,N_19841,N_19948);
or UO_515 (O_515,N_19900,N_19868);
nor UO_516 (O_516,N_19914,N_19987);
nor UO_517 (O_517,N_19869,N_19905);
nor UO_518 (O_518,N_19985,N_19860);
xor UO_519 (O_519,N_19914,N_19841);
nand UO_520 (O_520,N_19902,N_19955);
or UO_521 (O_521,N_19956,N_19874);
nand UO_522 (O_522,N_19938,N_19995);
and UO_523 (O_523,N_19915,N_19897);
nor UO_524 (O_524,N_19892,N_19903);
xnor UO_525 (O_525,N_19858,N_19864);
nor UO_526 (O_526,N_19894,N_19994);
and UO_527 (O_527,N_19958,N_19869);
xnor UO_528 (O_528,N_19847,N_19909);
and UO_529 (O_529,N_19889,N_19843);
xor UO_530 (O_530,N_19986,N_19995);
xor UO_531 (O_531,N_19872,N_19975);
nor UO_532 (O_532,N_19841,N_19900);
nor UO_533 (O_533,N_19866,N_19905);
nand UO_534 (O_534,N_19972,N_19947);
and UO_535 (O_535,N_19906,N_19851);
nor UO_536 (O_536,N_19847,N_19908);
or UO_537 (O_537,N_19984,N_19905);
or UO_538 (O_538,N_19966,N_19952);
nor UO_539 (O_539,N_19896,N_19868);
or UO_540 (O_540,N_19851,N_19873);
nor UO_541 (O_541,N_19860,N_19857);
or UO_542 (O_542,N_19888,N_19966);
nand UO_543 (O_543,N_19878,N_19991);
or UO_544 (O_544,N_19921,N_19893);
xnor UO_545 (O_545,N_19964,N_19878);
or UO_546 (O_546,N_19954,N_19934);
xnor UO_547 (O_547,N_19877,N_19878);
or UO_548 (O_548,N_19896,N_19929);
nor UO_549 (O_549,N_19886,N_19892);
or UO_550 (O_550,N_19968,N_19994);
xnor UO_551 (O_551,N_19916,N_19893);
or UO_552 (O_552,N_19914,N_19921);
and UO_553 (O_553,N_19968,N_19959);
or UO_554 (O_554,N_19968,N_19859);
and UO_555 (O_555,N_19863,N_19905);
nor UO_556 (O_556,N_19925,N_19990);
nand UO_557 (O_557,N_19948,N_19904);
nand UO_558 (O_558,N_19852,N_19969);
or UO_559 (O_559,N_19851,N_19888);
and UO_560 (O_560,N_19869,N_19995);
or UO_561 (O_561,N_19889,N_19892);
nand UO_562 (O_562,N_19926,N_19977);
or UO_563 (O_563,N_19980,N_19978);
nor UO_564 (O_564,N_19843,N_19936);
xor UO_565 (O_565,N_19914,N_19900);
xor UO_566 (O_566,N_19885,N_19850);
nor UO_567 (O_567,N_19971,N_19876);
or UO_568 (O_568,N_19977,N_19964);
nand UO_569 (O_569,N_19982,N_19952);
nor UO_570 (O_570,N_19998,N_19950);
nor UO_571 (O_571,N_19866,N_19927);
nand UO_572 (O_572,N_19857,N_19967);
or UO_573 (O_573,N_19935,N_19955);
nand UO_574 (O_574,N_19898,N_19921);
or UO_575 (O_575,N_19848,N_19962);
or UO_576 (O_576,N_19963,N_19989);
or UO_577 (O_577,N_19924,N_19916);
xnor UO_578 (O_578,N_19987,N_19850);
and UO_579 (O_579,N_19907,N_19958);
and UO_580 (O_580,N_19885,N_19942);
or UO_581 (O_581,N_19877,N_19841);
nand UO_582 (O_582,N_19876,N_19992);
or UO_583 (O_583,N_19853,N_19947);
and UO_584 (O_584,N_19994,N_19854);
xor UO_585 (O_585,N_19913,N_19908);
and UO_586 (O_586,N_19861,N_19928);
nor UO_587 (O_587,N_19987,N_19978);
or UO_588 (O_588,N_19957,N_19883);
and UO_589 (O_589,N_19942,N_19964);
and UO_590 (O_590,N_19980,N_19902);
and UO_591 (O_591,N_19978,N_19961);
and UO_592 (O_592,N_19951,N_19931);
xor UO_593 (O_593,N_19963,N_19882);
and UO_594 (O_594,N_19883,N_19984);
xor UO_595 (O_595,N_19951,N_19905);
or UO_596 (O_596,N_19925,N_19890);
nor UO_597 (O_597,N_19949,N_19930);
and UO_598 (O_598,N_19924,N_19930);
xor UO_599 (O_599,N_19987,N_19985);
xnor UO_600 (O_600,N_19873,N_19858);
or UO_601 (O_601,N_19925,N_19909);
or UO_602 (O_602,N_19917,N_19895);
and UO_603 (O_603,N_19988,N_19979);
nor UO_604 (O_604,N_19949,N_19845);
and UO_605 (O_605,N_19957,N_19848);
nor UO_606 (O_606,N_19965,N_19859);
or UO_607 (O_607,N_19855,N_19976);
nor UO_608 (O_608,N_19861,N_19870);
or UO_609 (O_609,N_19974,N_19918);
nor UO_610 (O_610,N_19844,N_19894);
nor UO_611 (O_611,N_19867,N_19916);
or UO_612 (O_612,N_19886,N_19900);
xor UO_613 (O_613,N_19937,N_19846);
nand UO_614 (O_614,N_19920,N_19843);
xor UO_615 (O_615,N_19930,N_19933);
or UO_616 (O_616,N_19841,N_19853);
nand UO_617 (O_617,N_19939,N_19925);
or UO_618 (O_618,N_19874,N_19932);
or UO_619 (O_619,N_19845,N_19948);
and UO_620 (O_620,N_19902,N_19938);
and UO_621 (O_621,N_19979,N_19846);
xnor UO_622 (O_622,N_19913,N_19972);
or UO_623 (O_623,N_19901,N_19928);
and UO_624 (O_624,N_19905,N_19961);
and UO_625 (O_625,N_19959,N_19881);
nand UO_626 (O_626,N_19910,N_19920);
or UO_627 (O_627,N_19983,N_19856);
or UO_628 (O_628,N_19952,N_19845);
xnor UO_629 (O_629,N_19950,N_19929);
or UO_630 (O_630,N_19977,N_19907);
nor UO_631 (O_631,N_19992,N_19962);
nand UO_632 (O_632,N_19916,N_19929);
nand UO_633 (O_633,N_19870,N_19965);
nor UO_634 (O_634,N_19856,N_19897);
nor UO_635 (O_635,N_19988,N_19875);
and UO_636 (O_636,N_19967,N_19953);
and UO_637 (O_637,N_19914,N_19946);
xnor UO_638 (O_638,N_19923,N_19932);
nand UO_639 (O_639,N_19856,N_19920);
and UO_640 (O_640,N_19996,N_19994);
nor UO_641 (O_641,N_19913,N_19932);
and UO_642 (O_642,N_19992,N_19964);
and UO_643 (O_643,N_19979,N_19904);
nand UO_644 (O_644,N_19906,N_19982);
nand UO_645 (O_645,N_19963,N_19982);
and UO_646 (O_646,N_19939,N_19856);
nor UO_647 (O_647,N_19901,N_19990);
or UO_648 (O_648,N_19982,N_19981);
nor UO_649 (O_649,N_19991,N_19857);
xnor UO_650 (O_650,N_19905,N_19989);
and UO_651 (O_651,N_19866,N_19980);
nand UO_652 (O_652,N_19966,N_19941);
nand UO_653 (O_653,N_19848,N_19852);
or UO_654 (O_654,N_19937,N_19917);
and UO_655 (O_655,N_19926,N_19877);
nand UO_656 (O_656,N_19967,N_19882);
nor UO_657 (O_657,N_19853,N_19996);
xnor UO_658 (O_658,N_19871,N_19983);
or UO_659 (O_659,N_19906,N_19846);
or UO_660 (O_660,N_19877,N_19961);
nor UO_661 (O_661,N_19868,N_19875);
nand UO_662 (O_662,N_19887,N_19895);
and UO_663 (O_663,N_19964,N_19915);
xnor UO_664 (O_664,N_19961,N_19888);
xnor UO_665 (O_665,N_19872,N_19925);
or UO_666 (O_666,N_19980,N_19946);
xnor UO_667 (O_667,N_19886,N_19925);
or UO_668 (O_668,N_19960,N_19943);
and UO_669 (O_669,N_19877,N_19907);
nor UO_670 (O_670,N_19955,N_19900);
nand UO_671 (O_671,N_19942,N_19999);
and UO_672 (O_672,N_19893,N_19908);
nand UO_673 (O_673,N_19926,N_19974);
or UO_674 (O_674,N_19993,N_19930);
nor UO_675 (O_675,N_19852,N_19905);
xor UO_676 (O_676,N_19840,N_19994);
nand UO_677 (O_677,N_19878,N_19870);
or UO_678 (O_678,N_19867,N_19875);
and UO_679 (O_679,N_19845,N_19921);
or UO_680 (O_680,N_19854,N_19855);
and UO_681 (O_681,N_19979,N_19862);
nor UO_682 (O_682,N_19965,N_19844);
nor UO_683 (O_683,N_19999,N_19895);
nor UO_684 (O_684,N_19948,N_19893);
and UO_685 (O_685,N_19945,N_19953);
xor UO_686 (O_686,N_19849,N_19889);
nor UO_687 (O_687,N_19976,N_19954);
nor UO_688 (O_688,N_19893,N_19856);
nand UO_689 (O_689,N_19884,N_19874);
and UO_690 (O_690,N_19957,N_19990);
or UO_691 (O_691,N_19970,N_19948);
and UO_692 (O_692,N_19909,N_19883);
nand UO_693 (O_693,N_19957,N_19926);
xnor UO_694 (O_694,N_19893,N_19918);
and UO_695 (O_695,N_19887,N_19852);
and UO_696 (O_696,N_19902,N_19920);
or UO_697 (O_697,N_19912,N_19974);
and UO_698 (O_698,N_19954,N_19879);
nor UO_699 (O_699,N_19961,N_19871);
or UO_700 (O_700,N_19940,N_19877);
xnor UO_701 (O_701,N_19942,N_19840);
xor UO_702 (O_702,N_19894,N_19862);
and UO_703 (O_703,N_19883,N_19962);
and UO_704 (O_704,N_19866,N_19990);
xor UO_705 (O_705,N_19896,N_19925);
nor UO_706 (O_706,N_19911,N_19843);
nor UO_707 (O_707,N_19918,N_19907);
or UO_708 (O_708,N_19866,N_19954);
nor UO_709 (O_709,N_19918,N_19936);
xnor UO_710 (O_710,N_19959,N_19997);
and UO_711 (O_711,N_19888,N_19949);
or UO_712 (O_712,N_19923,N_19968);
or UO_713 (O_713,N_19845,N_19961);
nand UO_714 (O_714,N_19914,N_19859);
and UO_715 (O_715,N_19944,N_19909);
and UO_716 (O_716,N_19911,N_19913);
or UO_717 (O_717,N_19847,N_19906);
and UO_718 (O_718,N_19958,N_19850);
and UO_719 (O_719,N_19867,N_19855);
xor UO_720 (O_720,N_19993,N_19982);
and UO_721 (O_721,N_19978,N_19848);
nand UO_722 (O_722,N_19980,N_19867);
or UO_723 (O_723,N_19987,N_19892);
or UO_724 (O_724,N_19937,N_19970);
nand UO_725 (O_725,N_19928,N_19878);
nand UO_726 (O_726,N_19906,N_19959);
nand UO_727 (O_727,N_19841,N_19895);
nand UO_728 (O_728,N_19871,N_19862);
nor UO_729 (O_729,N_19841,N_19967);
or UO_730 (O_730,N_19890,N_19963);
nand UO_731 (O_731,N_19847,N_19902);
or UO_732 (O_732,N_19844,N_19957);
nor UO_733 (O_733,N_19978,N_19862);
and UO_734 (O_734,N_19926,N_19879);
and UO_735 (O_735,N_19984,N_19944);
and UO_736 (O_736,N_19920,N_19956);
xor UO_737 (O_737,N_19929,N_19893);
nand UO_738 (O_738,N_19895,N_19953);
or UO_739 (O_739,N_19884,N_19949);
and UO_740 (O_740,N_19928,N_19974);
nor UO_741 (O_741,N_19916,N_19905);
or UO_742 (O_742,N_19930,N_19852);
or UO_743 (O_743,N_19943,N_19868);
xor UO_744 (O_744,N_19992,N_19927);
and UO_745 (O_745,N_19916,N_19897);
nand UO_746 (O_746,N_19847,N_19926);
xnor UO_747 (O_747,N_19938,N_19877);
nor UO_748 (O_748,N_19885,N_19890);
or UO_749 (O_749,N_19844,N_19950);
nand UO_750 (O_750,N_19917,N_19942);
or UO_751 (O_751,N_19893,N_19915);
nor UO_752 (O_752,N_19872,N_19990);
nand UO_753 (O_753,N_19998,N_19941);
and UO_754 (O_754,N_19928,N_19884);
and UO_755 (O_755,N_19898,N_19998);
and UO_756 (O_756,N_19992,N_19980);
nand UO_757 (O_757,N_19844,N_19922);
nand UO_758 (O_758,N_19872,N_19898);
nor UO_759 (O_759,N_19912,N_19881);
or UO_760 (O_760,N_19858,N_19934);
nand UO_761 (O_761,N_19873,N_19888);
nand UO_762 (O_762,N_19929,N_19925);
nand UO_763 (O_763,N_19878,N_19936);
nor UO_764 (O_764,N_19938,N_19919);
and UO_765 (O_765,N_19928,N_19847);
and UO_766 (O_766,N_19978,N_19890);
nand UO_767 (O_767,N_19881,N_19916);
or UO_768 (O_768,N_19987,N_19919);
or UO_769 (O_769,N_19988,N_19937);
and UO_770 (O_770,N_19905,N_19921);
xor UO_771 (O_771,N_19887,N_19938);
and UO_772 (O_772,N_19988,N_19906);
or UO_773 (O_773,N_19938,N_19872);
or UO_774 (O_774,N_19960,N_19840);
or UO_775 (O_775,N_19853,N_19978);
and UO_776 (O_776,N_19969,N_19985);
xnor UO_777 (O_777,N_19872,N_19862);
or UO_778 (O_778,N_19986,N_19857);
nand UO_779 (O_779,N_19968,N_19862);
nand UO_780 (O_780,N_19854,N_19862);
nor UO_781 (O_781,N_19998,N_19883);
and UO_782 (O_782,N_19958,N_19991);
or UO_783 (O_783,N_19902,N_19928);
nor UO_784 (O_784,N_19974,N_19861);
nor UO_785 (O_785,N_19851,N_19867);
or UO_786 (O_786,N_19959,N_19909);
or UO_787 (O_787,N_19876,N_19886);
xor UO_788 (O_788,N_19906,N_19859);
or UO_789 (O_789,N_19994,N_19895);
nand UO_790 (O_790,N_19918,N_19931);
xnor UO_791 (O_791,N_19955,N_19989);
nor UO_792 (O_792,N_19861,N_19912);
or UO_793 (O_793,N_19888,N_19901);
and UO_794 (O_794,N_19995,N_19918);
nand UO_795 (O_795,N_19867,N_19920);
nand UO_796 (O_796,N_19949,N_19982);
and UO_797 (O_797,N_19848,N_19932);
or UO_798 (O_798,N_19997,N_19902);
xnor UO_799 (O_799,N_19975,N_19886);
and UO_800 (O_800,N_19897,N_19847);
and UO_801 (O_801,N_19958,N_19993);
or UO_802 (O_802,N_19926,N_19909);
nand UO_803 (O_803,N_19947,N_19845);
nand UO_804 (O_804,N_19885,N_19930);
nand UO_805 (O_805,N_19897,N_19909);
and UO_806 (O_806,N_19975,N_19963);
or UO_807 (O_807,N_19851,N_19977);
or UO_808 (O_808,N_19952,N_19893);
and UO_809 (O_809,N_19919,N_19854);
xnor UO_810 (O_810,N_19962,N_19894);
or UO_811 (O_811,N_19860,N_19898);
or UO_812 (O_812,N_19887,N_19928);
or UO_813 (O_813,N_19991,N_19859);
nor UO_814 (O_814,N_19844,N_19909);
xnor UO_815 (O_815,N_19994,N_19868);
or UO_816 (O_816,N_19849,N_19980);
nor UO_817 (O_817,N_19942,N_19936);
and UO_818 (O_818,N_19884,N_19964);
nor UO_819 (O_819,N_19912,N_19927);
or UO_820 (O_820,N_19949,N_19886);
and UO_821 (O_821,N_19956,N_19852);
and UO_822 (O_822,N_19910,N_19924);
xnor UO_823 (O_823,N_19851,N_19850);
and UO_824 (O_824,N_19953,N_19903);
nand UO_825 (O_825,N_19860,N_19955);
or UO_826 (O_826,N_19980,N_19887);
nand UO_827 (O_827,N_19894,N_19925);
or UO_828 (O_828,N_19957,N_19977);
nand UO_829 (O_829,N_19874,N_19925);
nand UO_830 (O_830,N_19909,N_19868);
or UO_831 (O_831,N_19897,N_19842);
nor UO_832 (O_832,N_19927,N_19915);
nand UO_833 (O_833,N_19887,N_19940);
nand UO_834 (O_834,N_19909,N_19889);
or UO_835 (O_835,N_19902,N_19973);
nand UO_836 (O_836,N_19908,N_19982);
nand UO_837 (O_837,N_19912,N_19899);
xor UO_838 (O_838,N_19966,N_19870);
and UO_839 (O_839,N_19950,N_19940);
and UO_840 (O_840,N_19911,N_19993);
xnor UO_841 (O_841,N_19892,N_19966);
or UO_842 (O_842,N_19990,N_19867);
xnor UO_843 (O_843,N_19889,N_19868);
or UO_844 (O_844,N_19892,N_19943);
nand UO_845 (O_845,N_19895,N_19910);
or UO_846 (O_846,N_19843,N_19862);
or UO_847 (O_847,N_19982,N_19992);
or UO_848 (O_848,N_19980,N_19894);
or UO_849 (O_849,N_19956,N_19882);
nand UO_850 (O_850,N_19886,N_19941);
and UO_851 (O_851,N_19904,N_19931);
and UO_852 (O_852,N_19955,N_19922);
or UO_853 (O_853,N_19940,N_19959);
and UO_854 (O_854,N_19923,N_19857);
or UO_855 (O_855,N_19898,N_19867);
nor UO_856 (O_856,N_19866,N_19931);
xnor UO_857 (O_857,N_19922,N_19934);
xor UO_858 (O_858,N_19911,N_19942);
nor UO_859 (O_859,N_19860,N_19997);
and UO_860 (O_860,N_19928,N_19852);
nor UO_861 (O_861,N_19910,N_19995);
nand UO_862 (O_862,N_19949,N_19992);
nor UO_863 (O_863,N_19904,N_19888);
and UO_864 (O_864,N_19906,N_19863);
or UO_865 (O_865,N_19858,N_19916);
nand UO_866 (O_866,N_19873,N_19863);
nand UO_867 (O_867,N_19893,N_19896);
nand UO_868 (O_868,N_19941,N_19902);
and UO_869 (O_869,N_19860,N_19981);
and UO_870 (O_870,N_19904,N_19989);
and UO_871 (O_871,N_19929,N_19962);
and UO_872 (O_872,N_19869,N_19976);
nor UO_873 (O_873,N_19853,N_19932);
xor UO_874 (O_874,N_19907,N_19893);
nand UO_875 (O_875,N_19841,N_19860);
and UO_876 (O_876,N_19842,N_19890);
and UO_877 (O_877,N_19994,N_19955);
or UO_878 (O_878,N_19885,N_19961);
and UO_879 (O_879,N_19925,N_19892);
or UO_880 (O_880,N_19991,N_19924);
nand UO_881 (O_881,N_19879,N_19858);
and UO_882 (O_882,N_19912,N_19946);
and UO_883 (O_883,N_19919,N_19860);
xor UO_884 (O_884,N_19970,N_19887);
and UO_885 (O_885,N_19878,N_19917);
nor UO_886 (O_886,N_19954,N_19922);
or UO_887 (O_887,N_19941,N_19913);
nor UO_888 (O_888,N_19968,N_19863);
xnor UO_889 (O_889,N_19956,N_19945);
nand UO_890 (O_890,N_19865,N_19855);
nor UO_891 (O_891,N_19865,N_19868);
and UO_892 (O_892,N_19891,N_19985);
or UO_893 (O_893,N_19971,N_19980);
and UO_894 (O_894,N_19984,N_19869);
and UO_895 (O_895,N_19901,N_19932);
or UO_896 (O_896,N_19904,N_19934);
and UO_897 (O_897,N_19925,N_19904);
xnor UO_898 (O_898,N_19995,N_19873);
or UO_899 (O_899,N_19982,N_19936);
or UO_900 (O_900,N_19921,N_19863);
and UO_901 (O_901,N_19879,N_19844);
nand UO_902 (O_902,N_19940,N_19901);
xor UO_903 (O_903,N_19923,N_19894);
or UO_904 (O_904,N_19877,N_19923);
or UO_905 (O_905,N_19840,N_19878);
nand UO_906 (O_906,N_19891,N_19841);
and UO_907 (O_907,N_19987,N_19941);
or UO_908 (O_908,N_19881,N_19930);
xor UO_909 (O_909,N_19872,N_19876);
and UO_910 (O_910,N_19933,N_19897);
nor UO_911 (O_911,N_19926,N_19900);
nand UO_912 (O_912,N_19931,N_19846);
nand UO_913 (O_913,N_19879,N_19977);
nor UO_914 (O_914,N_19937,N_19966);
nand UO_915 (O_915,N_19864,N_19885);
nand UO_916 (O_916,N_19991,N_19940);
nor UO_917 (O_917,N_19923,N_19949);
nand UO_918 (O_918,N_19977,N_19952);
and UO_919 (O_919,N_19967,N_19983);
and UO_920 (O_920,N_19846,N_19987);
and UO_921 (O_921,N_19875,N_19922);
nor UO_922 (O_922,N_19851,N_19975);
nand UO_923 (O_923,N_19937,N_19965);
xnor UO_924 (O_924,N_19984,N_19973);
or UO_925 (O_925,N_19881,N_19875);
xor UO_926 (O_926,N_19928,N_19959);
and UO_927 (O_927,N_19968,N_19988);
or UO_928 (O_928,N_19883,N_19941);
or UO_929 (O_929,N_19972,N_19894);
or UO_930 (O_930,N_19952,N_19851);
and UO_931 (O_931,N_19955,N_19914);
nor UO_932 (O_932,N_19915,N_19851);
and UO_933 (O_933,N_19961,N_19929);
nand UO_934 (O_934,N_19961,N_19901);
nor UO_935 (O_935,N_19999,N_19983);
nand UO_936 (O_936,N_19883,N_19931);
and UO_937 (O_937,N_19973,N_19933);
nor UO_938 (O_938,N_19926,N_19899);
nand UO_939 (O_939,N_19997,N_19966);
nor UO_940 (O_940,N_19886,N_19848);
or UO_941 (O_941,N_19972,N_19910);
xor UO_942 (O_942,N_19984,N_19909);
xor UO_943 (O_943,N_19868,N_19946);
or UO_944 (O_944,N_19976,N_19910);
nor UO_945 (O_945,N_19905,N_19934);
nand UO_946 (O_946,N_19859,N_19954);
and UO_947 (O_947,N_19937,N_19891);
and UO_948 (O_948,N_19895,N_19966);
xnor UO_949 (O_949,N_19850,N_19903);
nor UO_950 (O_950,N_19870,N_19971);
nand UO_951 (O_951,N_19895,N_19901);
or UO_952 (O_952,N_19883,N_19943);
nand UO_953 (O_953,N_19984,N_19964);
nor UO_954 (O_954,N_19992,N_19939);
or UO_955 (O_955,N_19904,N_19897);
or UO_956 (O_956,N_19919,N_19873);
xnor UO_957 (O_957,N_19916,N_19843);
xnor UO_958 (O_958,N_19914,N_19918);
or UO_959 (O_959,N_19924,N_19994);
and UO_960 (O_960,N_19881,N_19922);
or UO_961 (O_961,N_19953,N_19965);
nand UO_962 (O_962,N_19894,N_19889);
and UO_963 (O_963,N_19847,N_19924);
nand UO_964 (O_964,N_19871,N_19852);
nand UO_965 (O_965,N_19919,N_19962);
nor UO_966 (O_966,N_19968,N_19882);
nor UO_967 (O_967,N_19996,N_19841);
xnor UO_968 (O_968,N_19863,N_19991);
or UO_969 (O_969,N_19904,N_19942);
or UO_970 (O_970,N_19917,N_19869);
or UO_971 (O_971,N_19863,N_19845);
and UO_972 (O_972,N_19953,N_19891);
xnor UO_973 (O_973,N_19874,N_19942);
nor UO_974 (O_974,N_19952,N_19844);
nor UO_975 (O_975,N_19998,N_19874);
or UO_976 (O_976,N_19896,N_19879);
or UO_977 (O_977,N_19862,N_19935);
or UO_978 (O_978,N_19878,N_19907);
nor UO_979 (O_979,N_19900,N_19984);
nand UO_980 (O_980,N_19964,N_19932);
or UO_981 (O_981,N_19950,N_19845);
or UO_982 (O_982,N_19847,N_19940);
xor UO_983 (O_983,N_19979,N_19875);
or UO_984 (O_984,N_19850,N_19894);
xnor UO_985 (O_985,N_19862,N_19941);
and UO_986 (O_986,N_19960,N_19847);
or UO_987 (O_987,N_19971,N_19934);
nand UO_988 (O_988,N_19901,N_19983);
or UO_989 (O_989,N_19987,N_19909);
nor UO_990 (O_990,N_19893,N_19961);
nor UO_991 (O_991,N_19994,N_19902);
nor UO_992 (O_992,N_19879,N_19913);
nor UO_993 (O_993,N_19845,N_19857);
or UO_994 (O_994,N_19867,N_19893);
nor UO_995 (O_995,N_19898,N_19938);
xor UO_996 (O_996,N_19847,N_19966);
or UO_997 (O_997,N_19997,N_19897);
xnor UO_998 (O_998,N_19841,N_19852);
nor UO_999 (O_999,N_19944,N_19961);
xor UO_1000 (O_1000,N_19910,N_19875);
nor UO_1001 (O_1001,N_19855,N_19896);
and UO_1002 (O_1002,N_19892,N_19883);
xor UO_1003 (O_1003,N_19948,N_19850);
nor UO_1004 (O_1004,N_19855,N_19850);
or UO_1005 (O_1005,N_19891,N_19941);
nor UO_1006 (O_1006,N_19852,N_19968);
nor UO_1007 (O_1007,N_19966,N_19970);
or UO_1008 (O_1008,N_19862,N_19891);
or UO_1009 (O_1009,N_19877,N_19919);
nor UO_1010 (O_1010,N_19908,N_19862);
nor UO_1011 (O_1011,N_19968,N_19865);
xnor UO_1012 (O_1012,N_19989,N_19950);
and UO_1013 (O_1013,N_19880,N_19895);
and UO_1014 (O_1014,N_19843,N_19938);
nor UO_1015 (O_1015,N_19861,N_19918);
nand UO_1016 (O_1016,N_19958,N_19892);
nor UO_1017 (O_1017,N_19962,N_19905);
or UO_1018 (O_1018,N_19984,N_19892);
xor UO_1019 (O_1019,N_19988,N_19962);
or UO_1020 (O_1020,N_19970,N_19986);
nand UO_1021 (O_1021,N_19904,N_19846);
nor UO_1022 (O_1022,N_19906,N_19871);
or UO_1023 (O_1023,N_19875,N_19909);
nand UO_1024 (O_1024,N_19971,N_19897);
and UO_1025 (O_1025,N_19845,N_19840);
or UO_1026 (O_1026,N_19894,N_19990);
xnor UO_1027 (O_1027,N_19883,N_19950);
and UO_1028 (O_1028,N_19983,N_19930);
or UO_1029 (O_1029,N_19929,N_19842);
xor UO_1030 (O_1030,N_19967,N_19949);
nand UO_1031 (O_1031,N_19972,N_19960);
or UO_1032 (O_1032,N_19928,N_19972);
nand UO_1033 (O_1033,N_19968,N_19984);
nand UO_1034 (O_1034,N_19888,N_19977);
nand UO_1035 (O_1035,N_19890,N_19937);
nor UO_1036 (O_1036,N_19928,N_19994);
nor UO_1037 (O_1037,N_19842,N_19846);
or UO_1038 (O_1038,N_19919,N_19997);
nor UO_1039 (O_1039,N_19846,N_19934);
nor UO_1040 (O_1040,N_19869,N_19899);
nand UO_1041 (O_1041,N_19984,N_19882);
nor UO_1042 (O_1042,N_19998,N_19848);
xnor UO_1043 (O_1043,N_19976,N_19927);
nor UO_1044 (O_1044,N_19935,N_19982);
nor UO_1045 (O_1045,N_19967,N_19918);
or UO_1046 (O_1046,N_19965,N_19915);
and UO_1047 (O_1047,N_19949,N_19939);
xnor UO_1048 (O_1048,N_19884,N_19932);
or UO_1049 (O_1049,N_19951,N_19995);
xnor UO_1050 (O_1050,N_19848,N_19931);
nor UO_1051 (O_1051,N_19968,N_19876);
nand UO_1052 (O_1052,N_19950,N_19959);
xnor UO_1053 (O_1053,N_19868,N_19918);
nand UO_1054 (O_1054,N_19881,N_19935);
nor UO_1055 (O_1055,N_19849,N_19874);
nor UO_1056 (O_1056,N_19983,N_19917);
xnor UO_1057 (O_1057,N_19909,N_19990);
xor UO_1058 (O_1058,N_19948,N_19977);
and UO_1059 (O_1059,N_19904,N_19872);
or UO_1060 (O_1060,N_19879,N_19851);
or UO_1061 (O_1061,N_19848,N_19903);
xor UO_1062 (O_1062,N_19856,N_19971);
nand UO_1063 (O_1063,N_19859,N_19940);
xnor UO_1064 (O_1064,N_19900,N_19918);
nand UO_1065 (O_1065,N_19955,N_19936);
or UO_1066 (O_1066,N_19933,N_19986);
xor UO_1067 (O_1067,N_19937,N_19870);
or UO_1068 (O_1068,N_19937,N_19989);
nand UO_1069 (O_1069,N_19841,N_19865);
nor UO_1070 (O_1070,N_19989,N_19935);
and UO_1071 (O_1071,N_19992,N_19978);
or UO_1072 (O_1072,N_19882,N_19957);
and UO_1073 (O_1073,N_19929,N_19942);
nand UO_1074 (O_1074,N_19906,N_19926);
xor UO_1075 (O_1075,N_19975,N_19966);
nand UO_1076 (O_1076,N_19990,N_19992);
and UO_1077 (O_1077,N_19992,N_19860);
xnor UO_1078 (O_1078,N_19922,N_19862);
or UO_1079 (O_1079,N_19844,N_19860);
nor UO_1080 (O_1080,N_19850,N_19907);
or UO_1081 (O_1081,N_19962,N_19886);
and UO_1082 (O_1082,N_19977,N_19869);
and UO_1083 (O_1083,N_19959,N_19926);
nand UO_1084 (O_1084,N_19937,N_19895);
xnor UO_1085 (O_1085,N_19961,N_19983);
nor UO_1086 (O_1086,N_19917,N_19975);
xor UO_1087 (O_1087,N_19878,N_19858);
and UO_1088 (O_1088,N_19848,N_19987);
nor UO_1089 (O_1089,N_19890,N_19942);
nor UO_1090 (O_1090,N_19899,N_19879);
nand UO_1091 (O_1091,N_19873,N_19883);
nor UO_1092 (O_1092,N_19949,N_19885);
or UO_1093 (O_1093,N_19896,N_19899);
xnor UO_1094 (O_1094,N_19862,N_19997);
and UO_1095 (O_1095,N_19967,N_19976);
and UO_1096 (O_1096,N_19872,N_19873);
nor UO_1097 (O_1097,N_19874,N_19873);
and UO_1098 (O_1098,N_19938,N_19920);
nand UO_1099 (O_1099,N_19848,N_19959);
nand UO_1100 (O_1100,N_19907,N_19905);
and UO_1101 (O_1101,N_19909,N_19879);
and UO_1102 (O_1102,N_19892,N_19924);
nor UO_1103 (O_1103,N_19954,N_19840);
and UO_1104 (O_1104,N_19895,N_19842);
or UO_1105 (O_1105,N_19916,N_19946);
and UO_1106 (O_1106,N_19997,N_19933);
nand UO_1107 (O_1107,N_19849,N_19938);
nand UO_1108 (O_1108,N_19840,N_19875);
nor UO_1109 (O_1109,N_19907,N_19855);
and UO_1110 (O_1110,N_19942,N_19973);
xor UO_1111 (O_1111,N_19914,N_19880);
nor UO_1112 (O_1112,N_19851,N_19846);
or UO_1113 (O_1113,N_19986,N_19931);
nand UO_1114 (O_1114,N_19922,N_19938);
xnor UO_1115 (O_1115,N_19874,N_19863);
or UO_1116 (O_1116,N_19867,N_19886);
xnor UO_1117 (O_1117,N_19904,N_19941);
nor UO_1118 (O_1118,N_19871,N_19855);
and UO_1119 (O_1119,N_19905,N_19902);
and UO_1120 (O_1120,N_19846,N_19909);
and UO_1121 (O_1121,N_19919,N_19951);
and UO_1122 (O_1122,N_19976,N_19980);
nand UO_1123 (O_1123,N_19935,N_19994);
nor UO_1124 (O_1124,N_19945,N_19978);
and UO_1125 (O_1125,N_19933,N_19972);
and UO_1126 (O_1126,N_19963,N_19959);
nor UO_1127 (O_1127,N_19848,N_19975);
and UO_1128 (O_1128,N_19899,N_19930);
xor UO_1129 (O_1129,N_19985,N_19949);
or UO_1130 (O_1130,N_19857,N_19949);
xor UO_1131 (O_1131,N_19998,N_19859);
xor UO_1132 (O_1132,N_19959,N_19937);
or UO_1133 (O_1133,N_19862,N_19955);
xor UO_1134 (O_1134,N_19946,N_19958);
or UO_1135 (O_1135,N_19857,N_19867);
or UO_1136 (O_1136,N_19873,N_19971);
and UO_1137 (O_1137,N_19974,N_19925);
nand UO_1138 (O_1138,N_19952,N_19875);
or UO_1139 (O_1139,N_19875,N_19978);
nand UO_1140 (O_1140,N_19947,N_19994);
and UO_1141 (O_1141,N_19841,N_19876);
xnor UO_1142 (O_1142,N_19927,N_19889);
nor UO_1143 (O_1143,N_19840,N_19841);
or UO_1144 (O_1144,N_19967,N_19902);
or UO_1145 (O_1145,N_19906,N_19914);
or UO_1146 (O_1146,N_19878,N_19987);
nand UO_1147 (O_1147,N_19894,N_19891);
or UO_1148 (O_1148,N_19938,N_19970);
nand UO_1149 (O_1149,N_19926,N_19886);
and UO_1150 (O_1150,N_19978,N_19850);
xor UO_1151 (O_1151,N_19955,N_19934);
and UO_1152 (O_1152,N_19855,N_19935);
nand UO_1153 (O_1153,N_19879,N_19953);
nand UO_1154 (O_1154,N_19882,N_19884);
xnor UO_1155 (O_1155,N_19925,N_19908);
xnor UO_1156 (O_1156,N_19942,N_19906);
nand UO_1157 (O_1157,N_19937,N_19907);
and UO_1158 (O_1158,N_19963,N_19957);
or UO_1159 (O_1159,N_19952,N_19998);
nand UO_1160 (O_1160,N_19948,N_19844);
and UO_1161 (O_1161,N_19953,N_19988);
xor UO_1162 (O_1162,N_19872,N_19857);
and UO_1163 (O_1163,N_19918,N_19958);
or UO_1164 (O_1164,N_19984,N_19950);
nand UO_1165 (O_1165,N_19949,N_19931);
or UO_1166 (O_1166,N_19858,N_19964);
nor UO_1167 (O_1167,N_19890,N_19974);
or UO_1168 (O_1168,N_19900,N_19964);
xor UO_1169 (O_1169,N_19980,N_19896);
and UO_1170 (O_1170,N_19930,N_19944);
xor UO_1171 (O_1171,N_19868,N_19932);
xnor UO_1172 (O_1172,N_19998,N_19866);
and UO_1173 (O_1173,N_19849,N_19886);
nor UO_1174 (O_1174,N_19873,N_19842);
and UO_1175 (O_1175,N_19852,N_19991);
xnor UO_1176 (O_1176,N_19978,N_19844);
nor UO_1177 (O_1177,N_19927,N_19885);
nand UO_1178 (O_1178,N_19866,N_19939);
nor UO_1179 (O_1179,N_19983,N_19947);
or UO_1180 (O_1180,N_19947,N_19957);
xnor UO_1181 (O_1181,N_19894,N_19993);
and UO_1182 (O_1182,N_19840,N_19844);
xnor UO_1183 (O_1183,N_19917,N_19978);
or UO_1184 (O_1184,N_19927,N_19972);
nor UO_1185 (O_1185,N_19999,N_19877);
or UO_1186 (O_1186,N_19987,N_19864);
xnor UO_1187 (O_1187,N_19869,N_19991);
and UO_1188 (O_1188,N_19849,N_19862);
nand UO_1189 (O_1189,N_19976,N_19981);
and UO_1190 (O_1190,N_19956,N_19843);
or UO_1191 (O_1191,N_19948,N_19924);
nand UO_1192 (O_1192,N_19873,N_19865);
nor UO_1193 (O_1193,N_19925,N_19946);
xor UO_1194 (O_1194,N_19933,N_19945);
nand UO_1195 (O_1195,N_19880,N_19866);
xor UO_1196 (O_1196,N_19852,N_19985);
nand UO_1197 (O_1197,N_19901,N_19951);
nand UO_1198 (O_1198,N_19891,N_19982);
nor UO_1199 (O_1199,N_19994,N_19986);
nand UO_1200 (O_1200,N_19928,N_19982);
and UO_1201 (O_1201,N_19977,N_19962);
or UO_1202 (O_1202,N_19969,N_19891);
and UO_1203 (O_1203,N_19989,N_19889);
nand UO_1204 (O_1204,N_19976,N_19908);
nor UO_1205 (O_1205,N_19994,N_19865);
or UO_1206 (O_1206,N_19878,N_19872);
and UO_1207 (O_1207,N_19940,N_19898);
or UO_1208 (O_1208,N_19921,N_19842);
or UO_1209 (O_1209,N_19855,N_19961);
nand UO_1210 (O_1210,N_19876,N_19955);
and UO_1211 (O_1211,N_19992,N_19909);
and UO_1212 (O_1212,N_19941,N_19898);
or UO_1213 (O_1213,N_19855,N_19903);
xnor UO_1214 (O_1214,N_19929,N_19860);
xnor UO_1215 (O_1215,N_19857,N_19953);
xnor UO_1216 (O_1216,N_19995,N_19970);
or UO_1217 (O_1217,N_19929,N_19849);
nand UO_1218 (O_1218,N_19921,N_19888);
nand UO_1219 (O_1219,N_19975,N_19871);
nand UO_1220 (O_1220,N_19850,N_19941);
nand UO_1221 (O_1221,N_19937,N_19885);
and UO_1222 (O_1222,N_19846,N_19864);
or UO_1223 (O_1223,N_19915,N_19995);
and UO_1224 (O_1224,N_19884,N_19876);
or UO_1225 (O_1225,N_19895,N_19900);
xnor UO_1226 (O_1226,N_19959,N_19912);
or UO_1227 (O_1227,N_19963,N_19885);
and UO_1228 (O_1228,N_19866,N_19947);
nand UO_1229 (O_1229,N_19889,N_19994);
or UO_1230 (O_1230,N_19919,N_19885);
and UO_1231 (O_1231,N_19899,N_19846);
nor UO_1232 (O_1232,N_19941,N_19905);
or UO_1233 (O_1233,N_19861,N_19891);
and UO_1234 (O_1234,N_19897,N_19978);
nand UO_1235 (O_1235,N_19945,N_19985);
xnor UO_1236 (O_1236,N_19991,N_19889);
or UO_1237 (O_1237,N_19938,N_19911);
and UO_1238 (O_1238,N_19900,N_19968);
nand UO_1239 (O_1239,N_19892,N_19995);
or UO_1240 (O_1240,N_19936,N_19893);
nor UO_1241 (O_1241,N_19929,N_19884);
or UO_1242 (O_1242,N_19843,N_19864);
nor UO_1243 (O_1243,N_19858,N_19881);
nor UO_1244 (O_1244,N_19988,N_19880);
xnor UO_1245 (O_1245,N_19880,N_19951);
xor UO_1246 (O_1246,N_19888,N_19889);
and UO_1247 (O_1247,N_19868,N_19880);
or UO_1248 (O_1248,N_19926,N_19936);
xnor UO_1249 (O_1249,N_19996,N_19885);
nand UO_1250 (O_1250,N_19967,N_19952);
or UO_1251 (O_1251,N_19969,N_19927);
xor UO_1252 (O_1252,N_19877,N_19967);
or UO_1253 (O_1253,N_19979,N_19863);
xnor UO_1254 (O_1254,N_19945,N_19889);
xor UO_1255 (O_1255,N_19953,N_19923);
or UO_1256 (O_1256,N_19961,N_19918);
nor UO_1257 (O_1257,N_19865,N_19857);
nor UO_1258 (O_1258,N_19914,N_19898);
nor UO_1259 (O_1259,N_19846,N_19975);
nand UO_1260 (O_1260,N_19856,N_19932);
nand UO_1261 (O_1261,N_19872,N_19851);
nand UO_1262 (O_1262,N_19927,N_19982);
or UO_1263 (O_1263,N_19993,N_19890);
nand UO_1264 (O_1264,N_19938,N_19886);
or UO_1265 (O_1265,N_19876,N_19930);
and UO_1266 (O_1266,N_19905,N_19945);
nand UO_1267 (O_1267,N_19924,N_19849);
and UO_1268 (O_1268,N_19947,N_19961);
nor UO_1269 (O_1269,N_19932,N_19997);
nand UO_1270 (O_1270,N_19900,N_19862);
nand UO_1271 (O_1271,N_19845,N_19904);
and UO_1272 (O_1272,N_19948,N_19950);
xor UO_1273 (O_1273,N_19874,N_19949);
nand UO_1274 (O_1274,N_19853,N_19981);
nor UO_1275 (O_1275,N_19870,N_19929);
nand UO_1276 (O_1276,N_19957,N_19896);
or UO_1277 (O_1277,N_19950,N_19922);
nand UO_1278 (O_1278,N_19930,N_19893);
or UO_1279 (O_1279,N_19863,N_19899);
xor UO_1280 (O_1280,N_19915,N_19901);
xnor UO_1281 (O_1281,N_19960,N_19853);
nor UO_1282 (O_1282,N_19939,N_19987);
nand UO_1283 (O_1283,N_19970,N_19860);
xnor UO_1284 (O_1284,N_19949,N_19968);
or UO_1285 (O_1285,N_19873,N_19936);
or UO_1286 (O_1286,N_19899,N_19979);
nand UO_1287 (O_1287,N_19893,N_19885);
nand UO_1288 (O_1288,N_19938,N_19971);
or UO_1289 (O_1289,N_19948,N_19945);
or UO_1290 (O_1290,N_19841,N_19930);
nand UO_1291 (O_1291,N_19938,N_19928);
xnor UO_1292 (O_1292,N_19905,N_19857);
nand UO_1293 (O_1293,N_19974,N_19920);
nor UO_1294 (O_1294,N_19948,N_19926);
xor UO_1295 (O_1295,N_19963,N_19953);
xor UO_1296 (O_1296,N_19902,N_19848);
nor UO_1297 (O_1297,N_19931,N_19999);
nand UO_1298 (O_1298,N_19992,N_19997);
or UO_1299 (O_1299,N_19878,N_19891);
xor UO_1300 (O_1300,N_19856,N_19935);
or UO_1301 (O_1301,N_19922,N_19966);
xnor UO_1302 (O_1302,N_19843,N_19961);
nor UO_1303 (O_1303,N_19890,N_19840);
and UO_1304 (O_1304,N_19909,N_19962);
and UO_1305 (O_1305,N_19919,N_19883);
and UO_1306 (O_1306,N_19855,N_19945);
or UO_1307 (O_1307,N_19900,N_19898);
nor UO_1308 (O_1308,N_19961,N_19996);
or UO_1309 (O_1309,N_19980,N_19985);
xnor UO_1310 (O_1310,N_19901,N_19853);
nand UO_1311 (O_1311,N_19964,N_19892);
nor UO_1312 (O_1312,N_19853,N_19892);
and UO_1313 (O_1313,N_19880,N_19853);
nand UO_1314 (O_1314,N_19900,N_19922);
xor UO_1315 (O_1315,N_19930,N_19996);
nor UO_1316 (O_1316,N_19939,N_19891);
nand UO_1317 (O_1317,N_19857,N_19913);
or UO_1318 (O_1318,N_19852,N_19899);
nand UO_1319 (O_1319,N_19898,N_19999);
xor UO_1320 (O_1320,N_19861,N_19989);
xor UO_1321 (O_1321,N_19870,N_19851);
nand UO_1322 (O_1322,N_19898,N_19887);
xnor UO_1323 (O_1323,N_19843,N_19879);
and UO_1324 (O_1324,N_19917,N_19952);
xor UO_1325 (O_1325,N_19960,N_19950);
and UO_1326 (O_1326,N_19895,N_19899);
nor UO_1327 (O_1327,N_19846,N_19865);
nor UO_1328 (O_1328,N_19917,N_19925);
xor UO_1329 (O_1329,N_19873,N_19950);
xor UO_1330 (O_1330,N_19854,N_19894);
or UO_1331 (O_1331,N_19887,N_19915);
and UO_1332 (O_1332,N_19987,N_19917);
nand UO_1333 (O_1333,N_19914,N_19853);
or UO_1334 (O_1334,N_19958,N_19874);
or UO_1335 (O_1335,N_19886,N_19915);
nand UO_1336 (O_1336,N_19887,N_19893);
nand UO_1337 (O_1337,N_19954,N_19862);
nand UO_1338 (O_1338,N_19932,N_19954);
xor UO_1339 (O_1339,N_19976,N_19891);
and UO_1340 (O_1340,N_19947,N_19849);
and UO_1341 (O_1341,N_19988,N_19903);
or UO_1342 (O_1342,N_19852,N_19883);
nand UO_1343 (O_1343,N_19843,N_19931);
xor UO_1344 (O_1344,N_19990,N_19987);
nor UO_1345 (O_1345,N_19885,N_19916);
xor UO_1346 (O_1346,N_19889,N_19877);
xor UO_1347 (O_1347,N_19973,N_19901);
nand UO_1348 (O_1348,N_19867,N_19986);
or UO_1349 (O_1349,N_19925,N_19996);
or UO_1350 (O_1350,N_19989,N_19875);
or UO_1351 (O_1351,N_19992,N_19979);
and UO_1352 (O_1352,N_19983,N_19866);
and UO_1353 (O_1353,N_19941,N_19894);
or UO_1354 (O_1354,N_19976,N_19985);
xor UO_1355 (O_1355,N_19916,N_19932);
nand UO_1356 (O_1356,N_19842,N_19915);
and UO_1357 (O_1357,N_19968,N_19898);
and UO_1358 (O_1358,N_19920,N_19891);
nor UO_1359 (O_1359,N_19859,N_19855);
xor UO_1360 (O_1360,N_19978,N_19895);
xnor UO_1361 (O_1361,N_19953,N_19876);
or UO_1362 (O_1362,N_19887,N_19867);
or UO_1363 (O_1363,N_19875,N_19956);
and UO_1364 (O_1364,N_19980,N_19899);
or UO_1365 (O_1365,N_19872,N_19841);
xnor UO_1366 (O_1366,N_19953,N_19885);
or UO_1367 (O_1367,N_19954,N_19875);
nand UO_1368 (O_1368,N_19948,N_19935);
xnor UO_1369 (O_1369,N_19859,N_19890);
xnor UO_1370 (O_1370,N_19933,N_19957);
nor UO_1371 (O_1371,N_19907,N_19927);
and UO_1372 (O_1372,N_19908,N_19881);
xor UO_1373 (O_1373,N_19959,N_19988);
nor UO_1374 (O_1374,N_19904,N_19984);
xor UO_1375 (O_1375,N_19994,N_19978);
and UO_1376 (O_1376,N_19856,N_19962);
and UO_1377 (O_1377,N_19925,N_19898);
nor UO_1378 (O_1378,N_19859,N_19869);
and UO_1379 (O_1379,N_19896,N_19911);
nand UO_1380 (O_1380,N_19913,N_19954);
nand UO_1381 (O_1381,N_19895,N_19845);
and UO_1382 (O_1382,N_19905,N_19885);
and UO_1383 (O_1383,N_19943,N_19882);
and UO_1384 (O_1384,N_19973,N_19917);
or UO_1385 (O_1385,N_19891,N_19875);
nor UO_1386 (O_1386,N_19904,N_19851);
and UO_1387 (O_1387,N_19907,N_19989);
nand UO_1388 (O_1388,N_19876,N_19916);
nor UO_1389 (O_1389,N_19847,N_19840);
xor UO_1390 (O_1390,N_19857,N_19910);
nand UO_1391 (O_1391,N_19844,N_19890);
xnor UO_1392 (O_1392,N_19935,N_19893);
or UO_1393 (O_1393,N_19868,N_19953);
nand UO_1394 (O_1394,N_19939,N_19864);
or UO_1395 (O_1395,N_19912,N_19844);
xnor UO_1396 (O_1396,N_19944,N_19997);
or UO_1397 (O_1397,N_19847,N_19868);
xor UO_1398 (O_1398,N_19981,N_19875);
nor UO_1399 (O_1399,N_19990,N_19855);
xor UO_1400 (O_1400,N_19963,N_19980);
and UO_1401 (O_1401,N_19853,N_19866);
and UO_1402 (O_1402,N_19849,N_19840);
nor UO_1403 (O_1403,N_19891,N_19847);
and UO_1404 (O_1404,N_19968,N_19913);
nand UO_1405 (O_1405,N_19987,N_19890);
nor UO_1406 (O_1406,N_19886,N_19869);
or UO_1407 (O_1407,N_19885,N_19918);
nand UO_1408 (O_1408,N_19878,N_19959);
xnor UO_1409 (O_1409,N_19871,N_19847);
nor UO_1410 (O_1410,N_19982,N_19914);
and UO_1411 (O_1411,N_19993,N_19862);
or UO_1412 (O_1412,N_19941,N_19969);
nor UO_1413 (O_1413,N_19860,N_19908);
nor UO_1414 (O_1414,N_19982,N_19980);
nand UO_1415 (O_1415,N_19891,N_19885);
or UO_1416 (O_1416,N_19935,N_19897);
nor UO_1417 (O_1417,N_19910,N_19901);
and UO_1418 (O_1418,N_19995,N_19885);
xnor UO_1419 (O_1419,N_19904,N_19994);
nor UO_1420 (O_1420,N_19929,N_19902);
nor UO_1421 (O_1421,N_19855,N_19962);
nor UO_1422 (O_1422,N_19973,N_19952);
and UO_1423 (O_1423,N_19886,N_19896);
nor UO_1424 (O_1424,N_19946,N_19927);
or UO_1425 (O_1425,N_19965,N_19852);
nor UO_1426 (O_1426,N_19901,N_19842);
nor UO_1427 (O_1427,N_19985,N_19937);
or UO_1428 (O_1428,N_19920,N_19893);
and UO_1429 (O_1429,N_19897,N_19859);
nor UO_1430 (O_1430,N_19957,N_19928);
or UO_1431 (O_1431,N_19893,N_19890);
nor UO_1432 (O_1432,N_19846,N_19866);
nand UO_1433 (O_1433,N_19946,N_19961);
nor UO_1434 (O_1434,N_19990,N_19885);
nor UO_1435 (O_1435,N_19946,N_19869);
nand UO_1436 (O_1436,N_19934,N_19931);
xor UO_1437 (O_1437,N_19997,N_19948);
and UO_1438 (O_1438,N_19851,N_19964);
nor UO_1439 (O_1439,N_19869,N_19841);
and UO_1440 (O_1440,N_19999,N_19996);
and UO_1441 (O_1441,N_19991,N_19896);
or UO_1442 (O_1442,N_19882,N_19962);
nand UO_1443 (O_1443,N_19912,N_19939);
and UO_1444 (O_1444,N_19999,N_19919);
xnor UO_1445 (O_1445,N_19904,N_19966);
nand UO_1446 (O_1446,N_19895,N_19934);
xor UO_1447 (O_1447,N_19934,N_19871);
xor UO_1448 (O_1448,N_19897,N_19876);
nor UO_1449 (O_1449,N_19888,N_19903);
or UO_1450 (O_1450,N_19994,N_19975);
nor UO_1451 (O_1451,N_19931,N_19845);
nand UO_1452 (O_1452,N_19952,N_19963);
xor UO_1453 (O_1453,N_19887,N_19912);
xnor UO_1454 (O_1454,N_19939,N_19985);
nor UO_1455 (O_1455,N_19948,N_19990);
nor UO_1456 (O_1456,N_19985,N_19910);
xor UO_1457 (O_1457,N_19955,N_19890);
xnor UO_1458 (O_1458,N_19889,N_19860);
nor UO_1459 (O_1459,N_19859,N_19844);
nand UO_1460 (O_1460,N_19953,N_19881);
xor UO_1461 (O_1461,N_19841,N_19887);
nand UO_1462 (O_1462,N_19899,N_19840);
and UO_1463 (O_1463,N_19874,N_19979);
nor UO_1464 (O_1464,N_19888,N_19936);
xnor UO_1465 (O_1465,N_19863,N_19901);
and UO_1466 (O_1466,N_19974,N_19937);
xnor UO_1467 (O_1467,N_19996,N_19880);
or UO_1468 (O_1468,N_19972,N_19922);
xor UO_1469 (O_1469,N_19990,N_19875);
and UO_1470 (O_1470,N_19994,N_19880);
nor UO_1471 (O_1471,N_19980,N_19997);
and UO_1472 (O_1472,N_19887,N_19976);
or UO_1473 (O_1473,N_19849,N_19870);
or UO_1474 (O_1474,N_19977,N_19920);
and UO_1475 (O_1475,N_19980,N_19908);
nor UO_1476 (O_1476,N_19921,N_19841);
nand UO_1477 (O_1477,N_19943,N_19980);
xnor UO_1478 (O_1478,N_19989,N_19858);
nand UO_1479 (O_1479,N_19997,N_19952);
and UO_1480 (O_1480,N_19997,N_19841);
or UO_1481 (O_1481,N_19980,N_19983);
nand UO_1482 (O_1482,N_19990,N_19968);
and UO_1483 (O_1483,N_19868,N_19840);
and UO_1484 (O_1484,N_19965,N_19935);
nand UO_1485 (O_1485,N_19880,N_19845);
nor UO_1486 (O_1486,N_19910,N_19957);
or UO_1487 (O_1487,N_19997,N_19886);
nor UO_1488 (O_1488,N_19869,N_19971);
and UO_1489 (O_1489,N_19975,N_19991);
nand UO_1490 (O_1490,N_19875,N_19953);
xnor UO_1491 (O_1491,N_19971,N_19841);
or UO_1492 (O_1492,N_19864,N_19999);
or UO_1493 (O_1493,N_19906,N_19934);
nor UO_1494 (O_1494,N_19845,N_19843);
nor UO_1495 (O_1495,N_19904,N_19869);
nor UO_1496 (O_1496,N_19991,N_19988);
xor UO_1497 (O_1497,N_19892,N_19907);
xor UO_1498 (O_1498,N_19960,N_19939);
nor UO_1499 (O_1499,N_19857,N_19983);
nor UO_1500 (O_1500,N_19986,N_19998);
or UO_1501 (O_1501,N_19851,N_19947);
xnor UO_1502 (O_1502,N_19986,N_19849);
and UO_1503 (O_1503,N_19921,N_19947);
or UO_1504 (O_1504,N_19960,N_19911);
nand UO_1505 (O_1505,N_19958,N_19911);
nand UO_1506 (O_1506,N_19882,N_19900);
nor UO_1507 (O_1507,N_19991,N_19928);
nor UO_1508 (O_1508,N_19954,N_19855);
or UO_1509 (O_1509,N_19983,N_19852);
or UO_1510 (O_1510,N_19966,N_19873);
nor UO_1511 (O_1511,N_19905,N_19846);
xnor UO_1512 (O_1512,N_19943,N_19860);
or UO_1513 (O_1513,N_19958,N_19844);
nor UO_1514 (O_1514,N_19929,N_19948);
xor UO_1515 (O_1515,N_19880,N_19967);
nand UO_1516 (O_1516,N_19989,N_19970);
or UO_1517 (O_1517,N_19993,N_19937);
and UO_1518 (O_1518,N_19845,N_19858);
nand UO_1519 (O_1519,N_19979,N_19985);
or UO_1520 (O_1520,N_19962,N_19842);
xor UO_1521 (O_1521,N_19954,N_19996);
nor UO_1522 (O_1522,N_19927,N_19894);
and UO_1523 (O_1523,N_19925,N_19994);
nor UO_1524 (O_1524,N_19865,N_19992);
xnor UO_1525 (O_1525,N_19897,N_19950);
xor UO_1526 (O_1526,N_19868,N_19866);
nor UO_1527 (O_1527,N_19936,N_19992);
nor UO_1528 (O_1528,N_19846,N_19940);
nand UO_1529 (O_1529,N_19857,N_19846);
xnor UO_1530 (O_1530,N_19841,N_19939);
nand UO_1531 (O_1531,N_19929,N_19977);
xnor UO_1532 (O_1532,N_19900,N_19887);
or UO_1533 (O_1533,N_19874,N_19872);
nor UO_1534 (O_1534,N_19968,N_19966);
nand UO_1535 (O_1535,N_19867,N_19856);
nor UO_1536 (O_1536,N_19908,N_19843);
and UO_1537 (O_1537,N_19969,N_19944);
xor UO_1538 (O_1538,N_19889,N_19985);
and UO_1539 (O_1539,N_19856,N_19948);
nor UO_1540 (O_1540,N_19875,N_19984);
or UO_1541 (O_1541,N_19907,N_19904);
nand UO_1542 (O_1542,N_19847,N_19971);
xor UO_1543 (O_1543,N_19931,N_19915);
xnor UO_1544 (O_1544,N_19891,N_19907);
and UO_1545 (O_1545,N_19975,N_19957);
nand UO_1546 (O_1546,N_19861,N_19842);
and UO_1547 (O_1547,N_19938,N_19968);
nand UO_1548 (O_1548,N_19960,N_19881);
nor UO_1549 (O_1549,N_19863,N_19960);
or UO_1550 (O_1550,N_19992,N_19885);
nand UO_1551 (O_1551,N_19999,N_19932);
xnor UO_1552 (O_1552,N_19855,N_19941);
nand UO_1553 (O_1553,N_19924,N_19950);
nand UO_1554 (O_1554,N_19862,N_19902);
xor UO_1555 (O_1555,N_19840,N_19948);
or UO_1556 (O_1556,N_19841,N_19855);
and UO_1557 (O_1557,N_19897,N_19949);
xnor UO_1558 (O_1558,N_19912,N_19878);
nor UO_1559 (O_1559,N_19932,N_19900);
nand UO_1560 (O_1560,N_19977,N_19958);
and UO_1561 (O_1561,N_19890,N_19850);
nand UO_1562 (O_1562,N_19848,N_19935);
or UO_1563 (O_1563,N_19945,N_19965);
nor UO_1564 (O_1564,N_19929,N_19933);
xnor UO_1565 (O_1565,N_19912,N_19952);
and UO_1566 (O_1566,N_19852,N_19914);
nand UO_1567 (O_1567,N_19965,N_19956);
nand UO_1568 (O_1568,N_19871,N_19893);
nand UO_1569 (O_1569,N_19861,N_19936);
or UO_1570 (O_1570,N_19998,N_19975);
or UO_1571 (O_1571,N_19889,N_19923);
and UO_1572 (O_1572,N_19967,N_19885);
nor UO_1573 (O_1573,N_19869,N_19872);
or UO_1574 (O_1574,N_19893,N_19987);
and UO_1575 (O_1575,N_19978,N_19951);
nand UO_1576 (O_1576,N_19848,N_19997);
xor UO_1577 (O_1577,N_19941,N_19946);
xnor UO_1578 (O_1578,N_19865,N_19947);
or UO_1579 (O_1579,N_19945,N_19954);
nand UO_1580 (O_1580,N_19912,N_19893);
nor UO_1581 (O_1581,N_19923,N_19926);
nor UO_1582 (O_1582,N_19879,N_19971);
xor UO_1583 (O_1583,N_19848,N_19911);
xor UO_1584 (O_1584,N_19907,N_19887);
nand UO_1585 (O_1585,N_19874,N_19953);
nor UO_1586 (O_1586,N_19943,N_19884);
xor UO_1587 (O_1587,N_19887,N_19926);
nand UO_1588 (O_1588,N_19925,N_19985);
nand UO_1589 (O_1589,N_19910,N_19992);
and UO_1590 (O_1590,N_19846,N_19849);
nand UO_1591 (O_1591,N_19848,N_19925);
nor UO_1592 (O_1592,N_19910,N_19980);
xnor UO_1593 (O_1593,N_19846,N_19863);
and UO_1594 (O_1594,N_19890,N_19867);
nor UO_1595 (O_1595,N_19921,N_19930);
nor UO_1596 (O_1596,N_19988,N_19946);
and UO_1597 (O_1597,N_19937,N_19877);
or UO_1598 (O_1598,N_19856,N_19985);
and UO_1599 (O_1599,N_19972,N_19992);
nor UO_1600 (O_1600,N_19969,N_19845);
and UO_1601 (O_1601,N_19863,N_19923);
nand UO_1602 (O_1602,N_19869,N_19973);
nand UO_1603 (O_1603,N_19869,N_19840);
and UO_1604 (O_1604,N_19934,N_19969);
nand UO_1605 (O_1605,N_19938,N_19952);
and UO_1606 (O_1606,N_19971,N_19892);
or UO_1607 (O_1607,N_19916,N_19866);
and UO_1608 (O_1608,N_19915,N_19942);
and UO_1609 (O_1609,N_19972,N_19884);
nand UO_1610 (O_1610,N_19998,N_19937);
nand UO_1611 (O_1611,N_19961,N_19881);
and UO_1612 (O_1612,N_19890,N_19872);
nand UO_1613 (O_1613,N_19882,N_19942);
nand UO_1614 (O_1614,N_19972,N_19855);
xor UO_1615 (O_1615,N_19966,N_19842);
xor UO_1616 (O_1616,N_19850,N_19960);
nand UO_1617 (O_1617,N_19912,N_19936);
nand UO_1618 (O_1618,N_19939,N_19867);
and UO_1619 (O_1619,N_19910,N_19943);
or UO_1620 (O_1620,N_19899,N_19960);
and UO_1621 (O_1621,N_19868,N_19974);
xnor UO_1622 (O_1622,N_19979,N_19864);
and UO_1623 (O_1623,N_19920,N_19991);
or UO_1624 (O_1624,N_19935,N_19932);
and UO_1625 (O_1625,N_19961,N_19990);
or UO_1626 (O_1626,N_19902,N_19939);
nand UO_1627 (O_1627,N_19859,N_19924);
xor UO_1628 (O_1628,N_19848,N_19890);
nor UO_1629 (O_1629,N_19872,N_19913);
or UO_1630 (O_1630,N_19920,N_19886);
xor UO_1631 (O_1631,N_19859,N_19900);
xnor UO_1632 (O_1632,N_19986,N_19954);
nand UO_1633 (O_1633,N_19863,N_19889);
xor UO_1634 (O_1634,N_19872,N_19950);
nor UO_1635 (O_1635,N_19983,N_19890);
xor UO_1636 (O_1636,N_19895,N_19931);
nand UO_1637 (O_1637,N_19881,N_19919);
or UO_1638 (O_1638,N_19917,N_19859);
nor UO_1639 (O_1639,N_19854,N_19859);
and UO_1640 (O_1640,N_19933,N_19881);
or UO_1641 (O_1641,N_19859,N_19894);
and UO_1642 (O_1642,N_19935,N_19967);
and UO_1643 (O_1643,N_19857,N_19885);
nand UO_1644 (O_1644,N_19938,N_19894);
or UO_1645 (O_1645,N_19963,N_19998);
xnor UO_1646 (O_1646,N_19929,N_19875);
xor UO_1647 (O_1647,N_19846,N_19889);
or UO_1648 (O_1648,N_19866,N_19987);
or UO_1649 (O_1649,N_19958,N_19877);
xnor UO_1650 (O_1650,N_19870,N_19893);
nand UO_1651 (O_1651,N_19869,N_19908);
nand UO_1652 (O_1652,N_19958,N_19995);
and UO_1653 (O_1653,N_19906,N_19841);
or UO_1654 (O_1654,N_19968,N_19855);
and UO_1655 (O_1655,N_19847,N_19907);
xor UO_1656 (O_1656,N_19937,N_19915);
or UO_1657 (O_1657,N_19993,N_19953);
nand UO_1658 (O_1658,N_19959,N_19998);
or UO_1659 (O_1659,N_19854,N_19852);
or UO_1660 (O_1660,N_19924,N_19947);
nor UO_1661 (O_1661,N_19873,N_19891);
xnor UO_1662 (O_1662,N_19938,N_19948);
or UO_1663 (O_1663,N_19955,N_19866);
or UO_1664 (O_1664,N_19929,N_19862);
xor UO_1665 (O_1665,N_19994,N_19903);
and UO_1666 (O_1666,N_19952,N_19840);
or UO_1667 (O_1667,N_19912,N_19851);
or UO_1668 (O_1668,N_19947,N_19855);
or UO_1669 (O_1669,N_19996,N_19857);
nand UO_1670 (O_1670,N_19925,N_19930);
nand UO_1671 (O_1671,N_19863,N_19857);
nor UO_1672 (O_1672,N_19840,N_19885);
xnor UO_1673 (O_1673,N_19840,N_19982);
nor UO_1674 (O_1674,N_19972,N_19844);
or UO_1675 (O_1675,N_19963,N_19872);
or UO_1676 (O_1676,N_19937,N_19860);
and UO_1677 (O_1677,N_19955,N_19874);
or UO_1678 (O_1678,N_19853,N_19921);
xnor UO_1679 (O_1679,N_19994,N_19941);
or UO_1680 (O_1680,N_19983,N_19860);
nand UO_1681 (O_1681,N_19977,N_19856);
and UO_1682 (O_1682,N_19921,N_19997);
nor UO_1683 (O_1683,N_19996,N_19847);
or UO_1684 (O_1684,N_19879,N_19902);
nor UO_1685 (O_1685,N_19844,N_19888);
nor UO_1686 (O_1686,N_19965,N_19948);
nand UO_1687 (O_1687,N_19854,N_19972);
nand UO_1688 (O_1688,N_19950,N_19851);
nor UO_1689 (O_1689,N_19948,N_19855);
nand UO_1690 (O_1690,N_19921,N_19871);
nand UO_1691 (O_1691,N_19874,N_19966);
nor UO_1692 (O_1692,N_19901,N_19936);
nand UO_1693 (O_1693,N_19845,N_19890);
and UO_1694 (O_1694,N_19952,N_19910);
xor UO_1695 (O_1695,N_19852,N_19937);
nand UO_1696 (O_1696,N_19909,N_19892);
or UO_1697 (O_1697,N_19997,N_19938);
and UO_1698 (O_1698,N_19993,N_19960);
nor UO_1699 (O_1699,N_19894,N_19919);
and UO_1700 (O_1700,N_19941,N_19843);
nor UO_1701 (O_1701,N_19847,N_19910);
or UO_1702 (O_1702,N_19974,N_19879);
nor UO_1703 (O_1703,N_19899,N_19858);
or UO_1704 (O_1704,N_19886,N_19928);
or UO_1705 (O_1705,N_19909,N_19977);
or UO_1706 (O_1706,N_19894,N_19987);
nand UO_1707 (O_1707,N_19903,N_19897);
or UO_1708 (O_1708,N_19876,N_19865);
nand UO_1709 (O_1709,N_19914,N_19943);
nor UO_1710 (O_1710,N_19861,N_19875);
or UO_1711 (O_1711,N_19986,N_19989);
and UO_1712 (O_1712,N_19894,N_19885);
xor UO_1713 (O_1713,N_19989,N_19844);
or UO_1714 (O_1714,N_19926,N_19861);
nand UO_1715 (O_1715,N_19988,N_19916);
or UO_1716 (O_1716,N_19911,N_19974);
or UO_1717 (O_1717,N_19840,N_19935);
xor UO_1718 (O_1718,N_19971,N_19904);
nor UO_1719 (O_1719,N_19863,N_19884);
and UO_1720 (O_1720,N_19892,N_19929);
nor UO_1721 (O_1721,N_19873,N_19954);
or UO_1722 (O_1722,N_19894,N_19950);
nand UO_1723 (O_1723,N_19893,N_19996);
or UO_1724 (O_1724,N_19972,N_19911);
nor UO_1725 (O_1725,N_19982,N_19850);
nor UO_1726 (O_1726,N_19975,N_19946);
and UO_1727 (O_1727,N_19973,N_19988);
xor UO_1728 (O_1728,N_19850,N_19889);
or UO_1729 (O_1729,N_19971,N_19910);
or UO_1730 (O_1730,N_19991,N_19974);
nor UO_1731 (O_1731,N_19933,N_19889);
and UO_1732 (O_1732,N_19893,N_19861);
and UO_1733 (O_1733,N_19916,N_19997);
nor UO_1734 (O_1734,N_19900,N_19842);
and UO_1735 (O_1735,N_19985,N_19920);
or UO_1736 (O_1736,N_19872,N_19893);
or UO_1737 (O_1737,N_19986,N_19860);
nand UO_1738 (O_1738,N_19925,N_19883);
or UO_1739 (O_1739,N_19878,N_19970);
and UO_1740 (O_1740,N_19944,N_19908);
and UO_1741 (O_1741,N_19946,N_19955);
nand UO_1742 (O_1742,N_19929,N_19992);
or UO_1743 (O_1743,N_19844,N_19852);
and UO_1744 (O_1744,N_19853,N_19888);
and UO_1745 (O_1745,N_19877,N_19872);
nand UO_1746 (O_1746,N_19867,N_19864);
and UO_1747 (O_1747,N_19997,N_19965);
and UO_1748 (O_1748,N_19987,N_19983);
nand UO_1749 (O_1749,N_19981,N_19886);
xor UO_1750 (O_1750,N_19870,N_19894);
or UO_1751 (O_1751,N_19964,N_19957);
nor UO_1752 (O_1752,N_19896,N_19856);
xor UO_1753 (O_1753,N_19882,N_19867);
xnor UO_1754 (O_1754,N_19938,N_19864);
nor UO_1755 (O_1755,N_19999,N_19883);
and UO_1756 (O_1756,N_19985,N_19868);
and UO_1757 (O_1757,N_19904,N_19914);
and UO_1758 (O_1758,N_19872,N_19905);
and UO_1759 (O_1759,N_19903,N_19885);
or UO_1760 (O_1760,N_19884,N_19926);
nand UO_1761 (O_1761,N_19854,N_19905);
and UO_1762 (O_1762,N_19990,N_19924);
and UO_1763 (O_1763,N_19865,N_19987);
xnor UO_1764 (O_1764,N_19937,N_19874);
and UO_1765 (O_1765,N_19896,N_19984);
and UO_1766 (O_1766,N_19850,N_19848);
and UO_1767 (O_1767,N_19909,N_19933);
xor UO_1768 (O_1768,N_19985,N_19918);
nand UO_1769 (O_1769,N_19924,N_19855);
xnor UO_1770 (O_1770,N_19940,N_19955);
nor UO_1771 (O_1771,N_19916,N_19908);
nor UO_1772 (O_1772,N_19883,N_19940);
and UO_1773 (O_1773,N_19845,N_19867);
or UO_1774 (O_1774,N_19840,N_19922);
and UO_1775 (O_1775,N_19966,N_19900);
and UO_1776 (O_1776,N_19997,N_19878);
and UO_1777 (O_1777,N_19963,N_19981);
and UO_1778 (O_1778,N_19882,N_19935);
or UO_1779 (O_1779,N_19975,N_19842);
nor UO_1780 (O_1780,N_19877,N_19959);
nor UO_1781 (O_1781,N_19976,N_19943);
and UO_1782 (O_1782,N_19949,N_19855);
or UO_1783 (O_1783,N_19984,N_19902);
xnor UO_1784 (O_1784,N_19945,N_19892);
nand UO_1785 (O_1785,N_19947,N_19857);
or UO_1786 (O_1786,N_19974,N_19936);
nand UO_1787 (O_1787,N_19928,N_19851);
nor UO_1788 (O_1788,N_19997,N_19893);
nor UO_1789 (O_1789,N_19986,N_19930);
and UO_1790 (O_1790,N_19939,N_19969);
nand UO_1791 (O_1791,N_19977,N_19972);
and UO_1792 (O_1792,N_19945,N_19896);
and UO_1793 (O_1793,N_19902,N_19900);
and UO_1794 (O_1794,N_19928,N_19931);
and UO_1795 (O_1795,N_19975,N_19849);
xor UO_1796 (O_1796,N_19975,N_19876);
nand UO_1797 (O_1797,N_19919,N_19937);
nor UO_1798 (O_1798,N_19953,N_19845);
and UO_1799 (O_1799,N_19968,N_19987);
nor UO_1800 (O_1800,N_19923,N_19954);
and UO_1801 (O_1801,N_19867,N_19997);
and UO_1802 (O_1802,N_19971,N_19885);
or UO_1803 (O_1803,N_19894,N_19953);
and UO_1804 (O_1804,N_19886,N_19947);
nand UO_1805 (O_1805,N_19907,N_19879);
nand UO_1806 (O_1806,N_19943,N_19956);
and UO_1807 (O_1807,N_19910,N_19898);
or UO_1808 (O_1808,N_19868,N_19951);
and UO_1809 (O_1809,N_19906,N_19950);
and UO_1810 (O_1810,N_19990,N_19900);
nand UO_1811 (O_1811,N_19857,N_19940);
and UO_1812 (O_1812,N_19934,N_19909);
or UO_1813 (O_1813,N_19907,N_19965);
nand UO_1814 (O_1814,N_19995,N_19883);
nand UO_1815 (O_1815,N_19979,N_19916);
nand UO_1816 (O_1816,N_19937,N_19936);
nor UO_1817 (O_1817,N_19965,N_19846);
xor UO_1818 (O_1818,N_19903,N_19910);
nand UO_1819 (O_1819,N_19902,N_19859);
and UO_1820 (O_1820,N_19860,N_19960);
and UO_1821 (O_1821,N_19915,N_19993);
or UO_1822 (O_1822,N_19868,N_19960);
nand UO_1823 (O_1823,N_19919,N_19976);
nor UO_1824 (O_1824,N_19964,N_19847);
and UO_1825 (O_1825,N_19899,N_19939);
nand UO_1826 (O_1826,N_19960,N_19931);
nand UO_1827 (O_1827,N_19879,N_19951);
and UO_1828 (O_1828,N_19846,N_19898);
and UO_1829 (O_1829,N_19914,N_19854);
nor UO_1830 (O_1830,N_19860,N_19968);
nand UO_1831 (O_1831,N_19847,N_19983);
and UO_1832 (O_1832,N_19903,N_19914);
and UO_1833 (O_1833,N_19979,N_19941);
nor UO_1834 (O_1834,N_19901,N_19972);
and UO_1835 (O_1835,N_19982,N_19861);
nand UO_1836 (O_1836,N_19923,N_19947);
xor UO_1837 (O_1837,N_19964,N_19983);
nand UO_1838 (O_1838,N_19952,N_19941);
xor UO_1839 (O_1839,N_19925,N_19948);
xnor UO_1840 (O_1840,N_19999,N_19909);
xnor UO_1841 (O_1841,N_19895,N_19875);
and UO_1842 (O_1842,N_19925,N_19916);
nand UO_1843 (O_1843,N_19958,N_19988);
nand UO_1844 (O_1844,N_19870,N_19855);
xnor UO_1845 (O_1845,N_19911,N_19915);
xnor UO_1846 (O_1846,N_19872,N_19916);
or UO_1847 (O_1847,N_19905,N_19975);
or UO_1848 (O_1848,N_19842,N_19905);
and UO_1849 (O_1849,N_19842,N_19942);
nand UO_1850 (O_1850,N_19905,N_19966);
xnor UO_1851 (O_1851,N_19880,N_19968);
or UO_1852 (O_1852,N_19894,N_19978);
nor UO_1853 (O_1853,N_19999,N_19885);
xor UO_1854 (O_1854,N_19945,N_19964);
or UO_1855 (O_1855,N_19988,N_19989);
xnor UO_1856 (O_1856,N_19859,N_19989);
or UO_1857 (O_1857,N_19859,N_19858);
nand UO_1858 (O_1858,N_19953,N_19947);
nor UO_1859 (O_1859,N_19935,N_19843);
nand UO_1860 (O_1860,N_19945,N_19906);
nand UO_1861 (O_1861,N_19862,N_19911);
or UO_1862 (O_1862,N_19841,N_19927);
nor UO_1863 (O_1863,N_19916,N_19896);
or UO_1864 (O_1864,N_19989,N_19862);
and UO_1865 (O_1865,N_19913,N_19986);
and UO_1866 (O_1866,N_19924,N_19881);
xnor UO_1867 (O_1867,N_19965,N_19995);
nor UO_1868 (O_1868,N_19917,N_19882);
or UO_1869 (O_1869,N_19908,N_19870);
nor UO_1870 (O_1870,N_19888,N_19940);
and UO_1871 (O_1871,N_19907,N_19872);
xor UO_1872 (O_1872,N_19863,N_19973);
and UO_1873 (O_1873,N_19846,N_19960);
nor UO_1874 (O_1874,N_19911,N_19878);
xor UO_1875 (O_1875,N_19875,N_19890);
xor UO_1876 (O_1876,N_19953,N_19867);
xor UO_1877 (O_1877,N_19865,N_19946);
or UO_1878 (O_1878,N_19850,N_19988);
nand UO_1879 (O_1879,N_19895,N_19891);
or UO_1880 (O_1880,N_19997,N_19863);
and UO_1881 (O_1881,N_19962,N_19891);
and UO_1882 (O_1882,N_19840,N_19973);
and UO_1883 (O_1883,N_19882,N_19911);
and UO_1884 (O_1884,N_19840,N_19850);
and UO_1885 (O_1885,N_19896,N_19955);
nand UO_1886 (O_1886,N_19958,N_19914);
or UO_1887 (O_1887,N_19842,N_19907);
nor UO_1888 (O_1888,N_19847,N_19899);
nand UO_1889 (O_1889,N_19977,N_19893);
nand UO_1890 (O_1890,N_19929,N_19963);
or UO_1891 (O_1891,N_19907,N_19994);
nor UO_1892 (O_1892,N_19951,N_19897);
nor UO_1893 (O_1893,N_19954,N_19918);
and UO_1894 (O_1894,N_19966,N_19903);
xnor UO_1895 (O_1895,N_19966,N_19972);
or UO_1896 (O_1896,N_19921,N_19948);
or UO_1897 (O_1897,N_19859,N_19925);
nand UO_1898 (O_1898,N_19847,N_19890);
xnor UO_1899 (O_1899,N_19857,N_19915);
xnor UO_1900 (O_1900,N_19993,N_19845);
nor UO_1901 (O_1901,N_19917,N_19862);
xor UO_1902 (O_1902,N_19909,N_19914);
xnor UO_1903 (O_1903,N_19886,N_19884);
or UO_1904 (O_1904,N_19981,N_19881);
nor UO_1905 (O_1905,N_19977,N_19970);
xor UO_1906 (O_1906,N_19873,N_19885);
or UO_1907 (O_1907,N_19895,N_19866);
nand UO_1908 (O_1908,N_19955,N_19873);
nand UO_1909 (O_1909,N_19923,N_19927);
nand UO_1910 (O_1910,N_19858,N_19893);
and UO_1911 (O_1911,N_19908,N_19872);
or UO_1912 (O_1912,N_19923,N_19991);
or UO_1913 (O_1913,N_19891,N_19966);
or UO_1914 (O_1914,N_19922,N_19920);
nor UO_1915 (O_1915,N_19860,N_19963);
nand UO_1916 (O_1916,N_19858,N_19986);
nor UO_1917 (O_1917,N_19984,N_19982);
or UO_1918 (O_1918,N_19934,N_19960);
nand UO_1919 (O_1919,N_19980,N_19909);
xor UO_1920 (O_1920,N_19943,N_19964);
nand UO_1921 (O_1921,N_19948,N_19889);
nand UO_1922 (O_1922,N_19973,N_19956);
xor UO_1923 (O_1923,N_19841,N_19897);
xor UO_1924 (O_1924,N_19873,N_19968);
or UO_1925 (O_1925,N_19909,N_19904);
xnor UO_1926 (O_1926,N_19882,N_19973);
xor UO_1927 (O_1927,N_19852,N_19923);
and UO_1928 (O_1928,N_19858,N_19930);
and UO_1929 (O_1929,N_19861,N_19947);
xor UO_1930 (O_1930,N_19926,N_19871);
or UO_1931 (O_1931,N_19963,N_19855);
xor UO_1932 (O_1932,N_19951,N_19845);
and UO_1933 (O_1933,N_19956,N_19961);
and UO_1934 (O_1934,N_19961,N_19906);
xnor UO_1935 (O_1935,N_19874,N_19928);
xnor UO_1936 (O_1936,N_19930,N_19963);
xnor UO_1937 (O_1937,N_19876,N_19877);
and UO_1938 (O_1938,N_19949,N_19975);
xor UO_1939 (O_1939,N_19925,N_19910);
nand UO_1940 (O_1940,N_19938,N_19925);
nor UO_1941 (O_1941,N_19883,N_19869);
or UO_1942 (O_1942,N_19863,N_19858);
nand UO_1943 (O_1943,N_19856,N_19902);
nor UO_1944 (O_1944,N_19979,N_19948);
xnor UO_1945 (O_1945,N_19895,N_19985);
and UO_1946 (O_1946,N_19875,N_19943);
and UO_1947 (O_1947,N_19917,N_19950);
xor UO_1948 (O_1948,N_19840,N_19944);
or UO_1949 (O_1949,N_19909,N_19932);
nand UO_1950 (O_1950,N_19936,N_19849);
or UO_1951 (O_1951,N_19865,N_19988);
nand UO_1952 (O_1952,N_19898,N_19974);
nand UO_1953 (O_1953,N_19984,N_19914);
or UO_1954 (O_1954,N_19933,N_19883);
nand UO_1955 (O_1955,N_19900,N_19929);
nor UO_1956 (O_1956,N_19864,N_19949);
nand UO_1957 (O_1957,N_19854,N_19991);
xor UO_1958 (O_1958,N_19855,N_19980);
or UO_1959 (O_1959,N_19995,N_19900);
or UO_1960 (O_1960,N_19976,N_19914);
xnor UO_1961 (O_1961,N_19966,N_19879);
nand UO_1962 (O_1962,N_19932,N_19933);
or UO_1963 (O_1963,N_19877,N_19945);
and UO_1964 (O_1964,N_19945,N_19870);
xnor UO_1965 (O_1965,N_19963,N_19896);
nand UO_1966 (O_1966,N_19904,N_19893);
and UO_1967 (O_1967,N_19946,N_19888);
and UO_1968 (O_1968,N_19840,N_19993);
xor UO_1969 (O_1969,N_19915,N_19883);
or UO_1970 (O_1970,N_19910,N_19882);
nand UO_1971 (O_1971,N_19901,N_19891);
and UO_1972 (O_1972,N_19940,N_19909);
xnor UO_1973 (O_1973,N_19928,N_19888);
or UO_1974 (O_1974,N_19994,N_19951);
nor UO_1975 (O_1975,N_19921,N_19999);
nor UO_1976 (O_1976,N_19993,N_19887);
xnor UO_1977 (O_1977,N_19883,N_19842);
or UO_1978 (O_1978,N_19875,N_19933);
nand UO_1979 (O_1979,N_19905,N_19861);
or UO_1980 (O_1980,N_19934,N_19850);
nand UO_1981 (O_1981,N_19920,N_19864);
nor UO_1982 (O_1982,N_19959,N_19996);
nand UO_1983 (O_1983,N_19915,N_19921);
nand UO_1984 (O_1984,N_19885,N_19842);
and UO_1985 (O_1985,N_19925,N_19877);
and UO_1986 (O_1986,N_19986,N_19886);
xnor UO_1987 (O_1987,N_19880,N_19884);
nor UO_1988 (O_1988,N_19879,N_19845);
nand UO_1989 (O_1989,N_19904,N_19895);
nand UO_1990 (O_1990,N_19907,N_19886);
nor UO_1991 (O_1991,N_19980,N_19869);
nor UO_1992 (O_1992,N_19914,N_19862);
or UO_1993 (O_1993,N_19985,N_19983);
or UO_1994 (O_1994,N_19848,N_19910);
and UO_1995 (O_1995,N_19855,N_19995);
nor UO_1996 (O_1996,N_19970,N_19877);
nor UO_1997 (O_1997,N_19955,N_19843);
nor UO_1998 (O_1998,N_19846,N_19994);
and UO_1999 (O_1999,N_19989,N_19968);
and UO_2000 (O_2000,N_19882,N_19940);
and UO_2001 (O_2001,N_19928,N_19943);
xnor UO_2002 (O_2002,N_19933,N_19871);
and UO_2003 (O_2003,N_19999,N_19995);
nand UO_2004 (O_2004,N_19952,N_19959);
nand UO_2005 (O_2005,N_19896,N_19932);
xnor UO_2006 (O_2006,N_19963,N_19866);
and UO_2007 (O_2007,N_19983,N_19926);
nand UO_2008 (O_2008,N_19987,N_19870);
and UO_2009 (O_2009,N_19870,N_19915);
and UO_2010 (O_2010,N_19973,N_19878);
or UO_2011 (O_2011,N_19886,N_19902);
nand UO_2012 (O_2012,N_19989,N_19947);
xor UO_2013 (O_2013,N_19968,N_19995);
nand UO_2014 (O_2014,N_19971,N_19915);
nor UO_2015 (O_2015,N_19878,N_19967);
nand UO_2016 (O_2016,N_19853,N_19859);
nor UO_2017 (O_2017,N_19879,N_19998);
and UO_2018 (O_2018,N_19955,N_19879);
nor UO_2019 (O_2019,N_19885,N_19901);
xnor UO_2020 (O_2020,N_19964,N_19978);
and UO_2021 (O_2021,N_19936,N_19885);
nor UO_2022 (O_2022,N_19964,N_19855);
and UO_2023 (O_2023,N_19915,N_19970);
and UO_2024 (O_2024,N_19874,N_19901);
nor UO_2025 (O_2025,N_19956,N_19947);
and UO_2026 (O_2026,N_19952,N_19931);
nand UO_2027 (O_2027,N_19918,N_19906);
xor UO_2028 (O_2028,N_19946,N_19954);
or UO_2029 (O_2029,N_19941,N_19870);
xor UO_2030 (O_2030,N_19896,N_19917);
or UO_2031 (O_2031,N_19976,N_19957);
and UO_2032 (O_2032,N_19876,N_19903);
xnor UO_2033 (O_2033,N_19934,N_19961);
xnor UO_2034 (O_2034,N_19924,N_19851);
nor UO_2035 (O_2035,N_19912,N_19869);
and UO_2036 (O_2036,N_19998,N_19871);
and UO_2037 (O_2037,N_19937,N_19921);
nor UO_2038 (O_2038,N_19948,N_19883);
or UO_2039 (O_2039,N_19944,N_19925);
or UO_2040 (O_2040,N_19970,N_19913);
xnor UO_2041 (O_2041,N_19973,N_19997);
nand UO_2042 (O_2042,N_19910,N_19904);
and UO_2043 (O_2043,N_19956,N_19976);
nor UO_2044 (O_2044,N_19987,N_19977);
and UO_2045 (O_2045,N_19982,N_19918);
nand UO_2046 (O_2046,N_19990,N_19869);
xor UO_2047 (O_2047,N_19928,N_19965);
nand UO_2048 (O_2048,N_19950,N_19985);
xor UO_2049 (O_2049,N_19879,N_19920);
nor UO_2050 (O_2050,N_19932,N_19880);
nand UO_2051 (O_2051,N_19873,N_19887);
or UO_2052 (O_2052,N_19853,N_19845);
or UO_2053 (O_2053,N_19978,N_19885);
nand UO_2054 (O_2054,N_19863,N_19867);
xnor UO_2055 (O_2055,N_19967,N_19933);
nor UO_2056 (O_2056,N_19859,N_19995);
nor UO_2057 (O_2057,N_19964,N_19905);
or UO_2058 (O_2058,N_19881,N_19995);
and UO_2059 (O_2059,N_19974,N_19947);
nor UO_2060 (O_2060,N_19995,N_19939);
and UO_2061 (O_2061,N_19975,N_19856);
or UO_2062 (O_2062,N_19846,N_19848);
xnor UO_2063 (O_2063,N_19967,N_19961);
xnor UO_2064 (O_2064,N_19850,N_19880);
xnor UO_2065 (O_2065,N_19882,N_19868);
nand UO_2066 (O_2066,N_19932,N_19891);
nand UO_2067 (O_2067,N_19854,N_19943);
and UO_2068 (O_2068,N_19994,N_19873);
xor UO_2069 (O_2069,N_19887,N_19880);
nand UO_2070 (O_2070,N_19932,N_19915);
nand UO_2071 (O_2071,N_19997,N_19880);
xnor UO_2072 (O_2072,N_19970,N_19875);
xor UO_2073 (O_2073,N_19977,N_19913);
nand UO_2074 (O_2074,N_19843,N_19898);
nor UO_2075 (O_2075,N_19925,N_19858);
or UO_2076 (O_2076,N_19945,N_19880);
and UO_2077 (O_2077,N_19967,N_19962);
nor UO_2078 (O_2078,N_19851,N_19882);
xor UO_2079 (O_2079,N_19962,N_19980);
and UO_2080 (O_2080,N_19973,N_19894);
xor UO_2081 (O_2081,N_19948,N_19930);
nand UO_2082 (O_2082,N_19894,N_19883);
and UO_2083 (O_2083,N_19862,N_19895);
or UO_2084 (O_2084,N_19901,N_19846);
nand UO_2085 (O_2085,N_19986,N_19908);
nand UO_2086 (O_2086,N_19987,N_19975);
xnor UO_2087 (O_2087,N_19932,N_19961);
nor UO_2088 (O_2088,N_19941,N_19881);
xnor UO_2089 (O_2089,N_19882,N_19856);
nand UO_2090 (O_2090,N_19899,N_19881);
nand UO_2091 (O_2091,N_19956,N_19958);
xor UO_2092 (O_2092,N_19967,N_19929);
nor UO_2093 (O_2093,N_19902,N_19935);
and UO_2094 (O_2094,N_19854,N_19902);
nor UO_2095 (O_2095,N_19958,N_19934);
xor UO_2096 (O_2096,N_19979,N_19896);
or UO_2097 (O_2097,N_19978,N_19866);
and UO_2098 (O_2098,N_19931,N_19932);
nor UO_2099 (O_2099,N_19917,N_19875);
nor UO_2100 (O_2100,N_19861,N_19844);
nor UO_2101 (O_2101,N_19907,N_19908);
nor UO_2102 (O_2102,N_19880,N_19885);
xor UO_2103 (O_2103,N_19980,N_19907);
or UO_2104 (O_2104,N_19946,N_19976);
nand UO_2105 (O_2105,N_19937,N_19909);
nor UO_2106 (O_2106,N_19926,N_19868);
or UO_2107 (O_2107,N_19984,N_19920);
or UO_2108 (O_2108,N_19970,N_19996);
nor UO_2109 (O_2109,N_19984,N_19985);
xor UO_2110 (O_2110,N_19898,N_19961);
nand UO_2111 (O_2111,N_19939,N_19857);
xor UO_2112 (O_2112,N_19946,N_19967);
xnor UO_2113 (O_2113,N_19927,N_19864);
and UO_2114 (O_2114,N_19938,N_19850);
nand UO_2115 (O_2115,N_19998,N_19888);
nor UO_2116 (O_2116,N_19903,N_19907);
nand UO_2117 (O_2117,N_19936,N_19875);
and UO_2118 (O_2118,N_19977,N_19898);
and UO_2119 (O_2119,N_19972,N_19976);
nor UO_2120 (O_2120,N_19924,N_19862);
nand UO_2121 (O_2121,N_19898,N_19920);
nand UO_2122 (O_2122,N_19998,N_19924);
nand UO_2123 (O_2123,N_19944,N_19926);
nor UO_2124 (O_2124,N_19860,N_19842);
xor UO_2125 (O_2125,N_19888,N_19854);
nor UO_2126 (O_2126,N_19872,N_19991);
or UO_2127 (O_2127,N_19996,N_19940);
or UO_2128 (O_2128,N_19992,N_19855);
xnor UO_2129 (O_2129,N_19874,N_19898);
and UO_2130 (O_2130,N_19970,N_19850);
nor UO_2131 (O_2131,N_19902,N_19863);
nor UO_2132 (O_2132,N_19892,N_19970);
nand UO_2133 (O_2133,N_19949,N_19850);
nor UO_2134 (O_2134,N_19868,N_19849);
nand UO_2135 (O_2135,N_19850,N_19857);
or UO_2136 (O_2136,N_19970,N_19857);
xor UO_2137 (O_2137,N_19940,N_19975);
nand UO_2138 (O_2138,N_19957,N_19955);
xor UO_2139 (O_2139,N_19995,N_19961);
nor UO_2140 (O_2140,N_19943,N_19919);
nand UO_2141 (O_2141,N_19947,N_19883);
or UO_2142 (O_2142,N_19970,N_19972);
or UO_2143 (O_2143,N_19947,N_19962);
xnor UO_2144 (O_2144,N_19889,N_19957);
or UO_2145 (O_2145,N_19915,N_19880);
nand UO_2146 (O_2146,N_19959,N_19932);
and UO_2147 (O_2147,N_19973,N_19977);
nand UO_2148 (O_2148,N_19921,N_19846);
and UO_2149 (O_2149,N_19964,N_19966);
xor UO_2150 (O_2150,N_19840,N_19854);
xnor UO_2151 (O_2151,N_19876,N_19962);
and UO_2152 (O_2152,N_19859,N_19929);
or UO_2153 (O_2153,N_19858,N_19936);
nand UO_2154 (O_2154,N_19908,N_19992);
or UO_2155 (O_2155,N_19840,N_19888);
and UO_2156 (O_2156,N_19956,N_19873);
or UO_2157 (O_2157,N_19983,N_19845);
or UO_2158 (O_2158,N_19962,N_19986);
or UO_2159 (O_2159,N_19862,N_19886);
or UO_2160 (O_2160,N_19928,N_19868);
or UO_2161 (O_2161,N_19924,N_19976);
xor UO_2162 (O_2162,N_19938,N_19890);
and UO_2163 (O_2163,N_19989,N_19845);
or UO_2164 (O_2164,N_19900,N_19852);
xnor UO_2165 (O_2165,N_19934,N_19897);
and UO_2166 (O_2166,N_19861,N_19899);
nand UO_2167 (O_2167,N_19974,N_19962);
nor UO_2168 (O_2168,N_19897,N_19986);
nor UO_2169 (O_2169,N_19872,N_19846);
or UO_2170 (O_2170,N_19917,N_19866);
nand UO_2171 (O_2171,N_19886,N_19983);
or UO_2172 (O_2172,N_19966,N_19897);
xor UO_2173 (O_2173,N_19840,N_19898);
or UO_2174 (O_2174,N_19857,N_19870);
nand UO_2175 (O_2175,N_19845,N_19971);
xnor UO_2176 (O_2176,N_19975,N_19968);
nand UO_2177 (O_2177,N_19938,N_19942);
nor UO_2178 (O_2178,N_19862,N_19998);
and UO_2179 (O_2179,N_19897,N_19862);
nand UO_2180 (O_2180,N_19931,N_19917);
nand UO_2181 (O_2181,N_19989,N_19908);
and UO_2182 (O_2182,N_19864,N_19921);
nor UO_2183 (O_2183,N_19919,N_19907);
or UO_2184 (O_2184,N_19921,N_19844);
or UO_2185 (O_2185,N_19951,N_19977);
xor UO_2186 (O_2186,N_19905,N_19841);
xnor UO_2187 (O_2187,N_19860,N_19848);
nor UO_2188 (O_2188,N_19974,N_19940);
nor UO_2189 (O_2189,N_19869,N_19898);
nor UO_2190 (O_2190,N_19990,N_19860);
and UO_2191 (O_2191,N_19881,N_19911);
nor UO_2192 (O_2192,N_19931,N_19963);
or UO_2193 (O_2193,N_19928,N_19950);
and UO_2194 (O_2194,N_19884,N_19923);
xnor UO_2195 (O_2195,N_19921,N_19897);
nand UO_2196 (O_2196,N_19854,N_19986);
nand UO_2197 (O_2197,N_19978,N_19984);
nor UO_2198 (O_2198,N_19870,N_19895);
xnor UO_2199 (O_2199,N_19866,N_19923);
or UO_2200 (O_2200,N_19916,N_19855);
xnor UO_2201 (O_2201,N_19892,N_19951);
or UO_2202 (O_2202,N_19919,N_19936);
or UO_2203 (O_2203,N_19855,N_19944);
or UO_2204 (O_2204,N_19883,N_19994);
and UO_2205 (O_2205,N_19890,N_19907);
xnor UO_2206 (O_2206,N_19855,N_19900);
xor UO_2207 (O_2207,N_19964,N_19990);
nor UO_2208 (O_2208,N_19976,N_19874);
nor UO_2209 (O_2209,N_19920,N_19992);
xnor UO_2210 (O_2210,N_19907,N_19985);
nor UO_2211 (O_2211,N_19914,N_19849);
and UO_2212 (O_2212,N_19872,N_19894);
nor UO_2213 (O_2213,N_19843,N_19998);
nand UO_2214 (O_2214,N_19953,N_19921);
or UO_2215 (O_2215,N_19922,N_19861);
xor UO_2216 (O_2216,N_19919,N_19845);
xor UO_2217 (O_2217,N_19983,N_19986);
and UO_2218 (O_2218,N_19994,N_19945);
and UO_2219 (O_2219,N_19843,N_19984);
or UO_2220 (O_2220,N_19907,N_19978);
nor UO_2221 (O_2221,N_19860,N_19852);
nand UO_2222 (O_2222,N_19953,N_19968);
nand UO_2223 (O_2223,N_19943,N_19859);
xnor UO_2224 (O_2224,N_19931,N_19886);
or UO_2225 (O_2225,N_19936,N_19988);
or UO_2226 (O_2226,N_19856,N_19914);
or UO_2227 (O_2227,N_19871,N_19981);
or UO_2228 (O_2228,N_19986,N_19958);
nor UO_2229 (O_2229,N_19957,N_19936);
nand UO_2230 (O_2230,N_19912,N_19872);
and UO_2231 (O_2231,N_19852,N_19864);
xor UO_2232 (O_2232,N_19844,N_19966);
and UO_2233 (O_2233,N_19846,N_19894);
nand UO_2234 (O_2234,N_19880,N_19858);
or UO_2235 (O_2235,N_19961,N_19974);
or UO_2236 (O_2236,N_19965,N_19865);
xnor UO_2237 (O_2237,N_19892,N_19877);
or UO_2238 (O_2238,N_19872,N_19852);
and UO_2239 (O_2239,N_19851,N_19982);
or UO_2240 (O_2240,N_19853,N_19991);
or UO_2241 (O_2241,N_19967,N_19943);
xor UO_2242 (O_2242,N_19891,N_19950);
nor UO_2243 (O_2243,N_19866,N_19855);
xor UO_2244 (O_2244,N_19847,N_19954);
or UO_2245 (O_2245,N_19949,N_19918);
and UO_2246 (O_2246,N_19945,N_19921);
nand UO_2247 (O_2247,N_19989,N_19884);
nand UO_2248 (O_2248,N_19876,N_19932);
or UO_2249 (O_2249,N_19901,N_19979);
nand UO_2250 (O_2250,N_19902,N_19916);
nand UO_2251 (O_2251,N_19938,N_19915);
nor UO_2252 (O_2252,N_19924,N_19907);
and UO_2253 (O_2253,N_19879,N_19904);
or UO_2254 (O_2254,N_19933,N_19904);
xor UO_2255 (O_2255,N_19877,N_19888);
or UO_2256 (O_2256,N_19972,N_19948);
nand UO_2257 (O_2257,N_19868,N_19854);
nand UO_2258 (O_2258,N_19914,N_19993);
nor UO_2259 (O_2259,N_19984,N_19998);
and UO_2260 (O_2260,N_19900,N_19979);
xnor UO_2261 (O_2261,N_19902,N_19885);
nor UO_2262 (O_2262,N_19928,N_19963);
and UO_2263 (O_2263,N_19950,N_19987);
nand UO_2264 (O_2264,N_19902,N_19869);
nand UO_2265 (O_2265,N_19938,N_19950);
nor UO_2266 (O_2266,N_19872,N_19977);
and UO_2267 (O_2267,N_19946,N_19970);
nand UO_2268 (O_2268,N_19913,N_19877);
nor UO_2269 (O_2269,N_19869,N_19918);
or UO_2270 (O_2270,N_19911,N_19910);
xor UO_2271 (O_2271,N_19882,N_19977);
nand UO_2272 (O_2272,N_19976,N_19878);
or UO_2273 (O_2273,N_19983,N_19897);
nand UO_2274 (O_2274,N_19881,N_19992);
xor UO_2275 (O_2275,N_19984,N_19986);
nand UO_2276 (O_2276,N_19958,N_19880);
nor UO_2277 (O_2277,N_19873,N_19868);
nor UO_2278 (O_2278,N_19983,N_19848);
nor UO_2279 (O_2279,N_19991,N_19841);
or UO_2280 (O_2280,N_19947,N_19980);
xnor UO_2281 (O_2281,N_19940,N_19947);
and UO_2282 (O_2282,N_19846,N_19860);
or UO_2283 (O_2283,N_19909,N_19946);
nand UO_2284 (O_2284,N_19976,N_19865);
nand UO_2285 (O_2285,N_19932,N_19989);
nor UO_2286 (O_2286,N_19924,N_19926);
nand UO_2287 (O_2287,N_19943,N_19924);
or UO_2288 (O_2288,N_19934,N_19984);
nor UO_2289 (O_2289,N_19897,N_19963);
or UO_2290 (O_2290,N_19934,N_19923);
nand UO_2291 (O_2291,N_19950,N_19991);
nor UO_2292 (O_2292,N_19882,N_19848);
nor UO_2293 (O_2293,N_19870,N_19942);
nand UO_2294 (O_2294,N_19963,N_19888);
xnor UO_2295 (O_2295,N_19961,N_19954);
nand UO_2296 (O_2296,N_19893,N_19857);
and UO_2297 (O_2297,N_19862,N_19846);
xor UO_2298 (O_2298,N_19983,N_19877);
and UO_2299 (O_2299,N_19971,N_19866);
nor UO_2300 (O_2300,N_19858,N_19943);
or UO_2301 (O_2301,N_19908,N_19957);
xnor UO_2302 (O_2302,N_19923,N_19933);
or UO_2303 (O_2303,N_19864,N_19942);
xnor UO_2304 (O_2304,N_19985,N_19874);
xnor UO_2305 (O_2305,N_19888,N_19978);
and UO_2306 (O_2306,N_19970,N_19904);
or UO_2307 (O_2307,N_19945,N_19939);
and UO_2308 (O_2308,N_19895,N_19916);
nand UO_2309 (O_2309,N_19918,N_19848);
nor UO_2310 (O_2310,N_19941,N_19880);
and UO_2311 (O_2311,N_19913,N_19990);
nand UO_2312 (O_2312,N_19962,N_19859);
nor UO_2313 (O_2313,N_19898,N_19875);
nand UO_2314 (O_2314,N_19865,N_19958);
xor UO_2315 (O_2315,N_19904,N_19999);
and UO_2316 (O_2316,N_19891,N_19849);
xor UO_2317 (O_2317,N_19922,N_19952);
nand UO_2318 (O_2318,N_19875,N_19865);
or UO_2319 (O_2319,N_19990,N_19996);
nor UO_2320 (O_2320,N_19986,N_19974);
xor UO_2321 (O_2321,N_19903,N_19900);
and UO_2322 (O_2322,N_19876,N_19871);
xor UO_2323 (O_2323,N_19846,N_19840);
nand UO_2324 (O_2324,N_19893,N_19913);
or UO_2325 (O_2325,N_19965,N_19858);
and UO_2326 (O_2326,N_19983,N_19870);
or UO_2327 (O_2327,N_19840,N_19987);
and UO_2328 (O_2328,N_19938,N_19880);
xor UO_2329 (O_2329,N_19932,N_19973);
and UO_2330 (O_2330,N_19929,N_19909);
xor UO_2331 (O_2331,N_19972,N_19866);
nand UO_2332 (O_2332,N_19875,N_19849);
or UO_2333 (O_2333,N_19859,N_19935);
nand UO_2334 (O_2334,N_19966,N_19893);
xor UO_2335 (O_2335,N_19907,N_19858);
nand UO_2336 (O_2336,N_19997,N_19935);
nor UO_2337 (O_2337,N_19917,N_19954);
or UO_2338 (O_2338,N_19860,N_19989);
nor UO_2339 (O_2339,N_19930,N_19945);
or UO_2340 (O_2340,N_19978,N_19966);
xnor UO_2341 (O_2341,N_19848,N_19900);
xor UO_2342 (O_2342,N_19917,N_19855);
and UO_2343 (O_2343,N_19914,N_19878);
or UO_2344 (O_2344,N_19885,N_19939);
nor UO_2345 (O_2345,N_19907,N_19921);
and UO_2346 (O_2346,N_19917,N_19865);
nand UO_2347 (O_2347,N_19914,N_19968);
or UO_2348 (O_2348,N_19842,N_19938);
xnor UO_2349 (O_2349,N_19863,N_19970);
and UO_2350 (O_2350,N_19881,N_19847);
nor UO_2351 (O_2351,N_19958,N_19891);
or UO_2352 (O_2352,N_19903,N_19995);
xor UO_2353 (O_2353,N_19961,N_19844);
and UO_2354 (O_2354,N_19853,N_19930);
nor UO_2355 (O_2355,N_19905,N_19919);
nand UO_2356 (O_2356,N_19994,N_19912);
xnor UO_2357 (O_2357,N_19904,N_19951);
nand UO_2358 (O_2358,N_19900,N_19997);
xor UO_2359 (O_2359,N_19891,N_19946);
xnor UO_2360 (O_2360,N_19863,N_19861);
nand UO_2361 (O_2361,N_19997,N_19957);
xnor UO_2362 (O_2362,N_19911,N_19873);
nor UO_2363 (O_2363,N_19956,N_19872);
nand UO_2364 (O_2364,N_19891,N_19856);
and UO_2365 (O_2365,N_19972,N_19870);
nor UO_2366 (O_2366,N_19987,N_19982);
or UO_2367 (O_2367,N_19951,N_19933);
xor UO_2368 (O_2368,N_19892,N_19869);
and UO_2369 (O_2369,N_19957,N_19935);
nor UO_2370 (O_2370,N_19858,N_19944);
nor UO_2371 (O_2371,N_19864,N_19888);
nand UO_2372 (O_2372,N_19865,N_19859);
and UO_2373 (O_2373,N_19909,N_19905);
and UO_2374 (O_2374,N_19872,N_19892);
or UO_2375 (O_2375,N_19852,N_19845);
and UO_2376 (O_2376,N_19919,N_19990);
xnor UO_2377 (O_2377,N_19990,N_19897);
nor UO_2378 (O_2378,N_19860,N_19971);
and UO_2379 (O_2379,N_19890,N_19920);
or UO_2380 (O_2380,N_19906,N_19998);
and UO_2381 (O_2381,N_19850,N_19979);
or UO_2382 (O_2382,N_19922,N_19982);
or UO_2383 (O_2383,N_19917,N_19912);
nor UO_2384 (O_2384,N_19866,N_19959);
nor UO_2385 (O_2385,N_19898,N_19948);
xnor UO_2386 (O_2386,N_19873,N_19903);
nand UO_2387 (O_2387,N_19957,N_19969);
nand UO_2388 (O_2388,N_19900,N_19946);
and UO_2389 (O_2389,N_19973,N_19929);
and UO_2390 (O_2390,N_19926,N_19956);
and UO_2391 (O_2391,N_19990,N_19857);
or UO_2392 (O_2392,N_19972,N_19908);
and UO_2393 (O_2393,N_19983,N_19996);
xor UO_2394 (O_2394,N_19903,N_19896);
and UO_2395 (O_2395,N_19968,N_19982);
nor UO_2396 (O_2396,N_19841,N_19848);
nor UO_2397 (O_2397,N_19897,N_19953);
nand UO_2398 (O_2398,N_19867,N_19951);
or UO_2399 (O_2399,N_19972,N_19936);
or UO_2400 (O_2400,N_19972,N_19915);
nand UO_2401 (O_2401,N_19976,N_19929);
xnor UO_2402 (O_2402,N_19852,N_19846);
or UO_2403 (O_2403,N_19971,N_19970);
xor UO_2404 (O_2404,N_19934,N_19860);
xor UO_2405 (O_2405,N_19901,N_19933);
nor UO_2406 (O_2406,N_19899,N_19981);
nand UO_2407 (O_2407,N_19926,N_19993);
and UO_2408 (O_2408,N_19954,N_19979);
nand UO_2409 (O_2409,N_19842,N_19903);
and UO_2410 (O_2410,N_19871,N_19992);
nand UO_2411 (O_2411,N_19901,N_19868);
or UO_2412 (O_2412,N_19972,N_19892);
xnor UO_2413 (O_2413,N_19868,N_19895);
and UO_2414 (O_2414,N_19905,N_19959);
and UO_2415 (O_2415,N_19897,N_19993);
and UO_2416 (O_2416,N_19893,N_19964);
or UO_2417 (O_2417,N_19857,N_19877);
nor UO_2418 (O_2418,N_19980,N_19950);
or UO_2419 (O_2419,N_19928,N_19975);
nand UO_2420 (O_2420,N_19933,N_19995);
xor UO_2421 (O_2421,N_19934,N_19936);
nand UO_2422 (O_2422,N_19967,N_19874);
nand UO_2423 (O_2423,N_19947,N_19894);
nand UO_2424 (O_2424,N_19901,N_19921);
xor UO_2425 (O_2425,N_19919,N_19850);
and UO_2426 (O_2426,N_19878,N_19924);
and UO_2427 (O_2427,N_19944,N_19958);
nand UO_2428 (O_2428,N_19980,N_19939);
or UO_2429 (O_2429,N_19912,N_19997);
xor UO_2430 (O_2430,N_19869,N_19922);
or UO_2431 (O_2431,N_19967,N_19855);
and UO_2432 (O_2432,N_19981,N_19971);
xnor UO_2433 (O_2433,N_19920,N_19869);
xnor UO_2434 (O_2434,N_19912,N_19934);
xor UO_2435 (O_2435,N_19957,N_19872);
and UO_2436 (O_2436,N_19927,N_19888);
nand UO_2437 (O_2437,N_19934,N_19945);
and UO_2438 (O_2438,N_19947,N_19909);
xor UO_2439 (O_2439,N_19998,N_19961);
xnor UO_2440 (O_2440,N_19937,N_19896);
xor UO_2441 (O_2441,N_19841,N_19987);
or UO_2442 (O_2442,N_19965,N_19982);
or UO_2443 (O_2443,N_19955,N_19971);
or UO_2444 (O_2444,N_19899,N_19946);
or UO_2445 (O_2445,N_19881,N_19921);
and UO_2446 (O_2446,N_19922,N_19944);
nand UO_2447 (O_2447,N_19920,N_19955);
nor UO_2448 (O_2448,N_19864,N_19910);
or UO_2449 (O_2449,N_19879,N_19937);
nand UO_2450 (O_2450,N_19929,N_19940);
xnor UO_2451 (O_2451,N_19937,N_19886);
nor UO_2452 (O_2452,N_19867,N_19959);
nor UO_2453 (O_2453,N_19926,N_19870);
xnor UO_2454 (O_2454,N_19987,N_19895);
or UO_2455 (O_2455,N_19868,N_19937);
nand UO_2456 (O_2456,N_19924,N_19987);
nor UO_2457 (O_2457,N_19981,N_19915);
and UO_2458 (O_2458,N_19840,N_19919);
nor UO_2459 (O_2459,N_19856,N_19943);
nor UO_2460 (O_2460,N_19957,N_19855);
nor UO_2461 (O_2461,N_19964,N_19881);
or UO_2462 (O_2462,N_19849,N_19899);
nand UO_2463 (O_2463,N_19899,N_19997);
nor UO_2464 (O_2464,N_19971,N_19976);
and UO_2465 (O_2465,N_19992,N_19856);
or UO_2466 (O_2466,N_19988,N_19982);
nor UO_2467 (O_2467,N_19884,N_19897);
and UO_2468 (O_2468,N_19840,N_19965);
nor UO_2469 (O_2469,N_19938,N_19974);
xor UO_2470 (O_2470,N_19943,N_19886);
nand UO_2471 (O_2471,N_19879,N_19924);
nor UO_2472 (O_2472,N_19942,N_19988);
nor UO_2473 (O_2473,N_19922,N_19857);
xnor UO_2474 (O_2474,N_19946,N_19903);
xnor UO_2475 (O_2475,N_19925,N_19867);
or UO_2476 (O_2476,N_19903,N_19951);
or UO_2477 (O_2477,N_19909,N_19882);
or UO_2478 (O_2478,N_19984,N_19990);
nand UO_2479 (O_2479,N_19881,N_19901);
nor UO_2480 (O_2480,N_19901,N_19905);
or UO_2481 (O_2481,N_19957,N_19843);
nor UO_2482 (O_2482,N_19867,N_19860);
or UO_2483 (O_2483,N_19841,N_19883);
nor UO_2484 (O_2484,N_19877,N_19902);
nor UO_2485 (O_2485,N_19958,N_19894);
nand UO_2486 (O_2486,N_19932,N_19886);
xnor UO_2487 (O_2487,N_19977,N_19853);
nor UO_2488 (O_2488,N_19898,N_19924);
nor UO_2489 (O_2489,N_19969,N_19913);
xor UO_2490 (O_2490,N_19844,N_19964);
or UO_2491 (O_2491,N_19851,N_19936);
or UO_2492 (O_2492,N_19850,N_19929);
xnor UO_2493 (O_2493,N_19859,N_19967);
nor UO_2494 (O_2494,N_19865,N_19878);
nand UO_2495 (O_2495,N_19998,N_19892);
or UO_2496 (O_2496,N_19917,N_19848);
nand UO_2497 (O_2497,N_19900,N_19870);
and UO_2498 (O_2498,N_19879,N_19964);
xnor UO_2499 (O_2499,N_19840,N_19979);
endmodule