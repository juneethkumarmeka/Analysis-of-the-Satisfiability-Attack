module basic_2000_20000_2500_40_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_987,In_1600);
and U1 (N_1,In_1383,In_863);
nor U2 (N_2,In_754,In_1252);
nor U3 (N_3,In_832,In_361);
nor U4 (N_4,In_216,In_242);
nor U5 (N_5,In_1615,In_59);
nand U6 (N_6,In_110,In_1121);
nand U7 (N_7,In_1443,In_427);
nand U8 (N_8,In_667,In_606);
nor U9 (N_9,In_1965,In_683);
nor U10 (N_10,In_1424,In_707);
or U11 (N_11,In_120,In_1685);
nand U12 (N_12,In_1039,In_390);
or U13 (N_13,In_353,In_946);
or U14 (N_14,In_1516,In_1502);
or U15 (N_15,In_652,In_1228);
and U16 (N_16,In_664,In_457);
and U17 (N_17,In_1710,In_1298);
nand U18 (N_18,In_116,In_200);
or U19 (N_19,In_1647,In_849);
nand U20 (N_20,In_1519,In_875);
or U21 (N_21,In_412,In_223);
and U22 (N_22,In_1003,In_1489);
and U23 (N_23,In_1782,In_1898);
nor U24 (N_24,In_592,In_1990);
and U25 (N_25,In_90,In_382);
and U26 (N_26,In_559,In_705);
nor U27 (N_27,In_1587,In_1896);
or U28 (N_28,In_1353,In_1620);
nand U29 (N_29,In_1104,In_1708);
and U30 (N_30,In_338,In_1068);
and U31 (N_31,In_1037,In_1688);
and U32 (N_32,In_481,In_1787);
and U33 (N_33,In_1726,In_609);
nor U34 (N_34,In_1011,In_1741);
nand U35 (N_35,In_1404,In_9);
nand U36 (N_36,In_1805,In_1700);
nor U37 (N_37,In_929,In_607);
and U38 (N_38,In_1016,In_1450);
nor U39 (N_39,In_1374,In_253);
xor U40 (N_40,In_1268,In_673);
nand U41 (N_41,In_969,In_1638);
and U42 (N_42,In_750,In_1105);
nand U43 (N_43,In_1999,In_2);
xnor U44 (N_44,In_307,In_380);
nand U45 (N_45,In_212,In_1528);
nor U46 (N_46,In_1623,In_636);
nand U47 (N_47,In_171,In_1000);
and U48 (N_48,In_1265,In_260);
or U49 (N_49,In_1259,In_1818);
and U50 (N_50,In_419,In_1789);
nand U51 (N_51,In_1996,In_1807);
nor U52 (N_52,In_947,In_1276);
nand U53 (N_53,In_348,In_240);
nand U54 (N_54,In_1018,In_1695);
nand U55 (N_55,In_1233,In_1526);
nand U56 (N_56,In_550,In_1014);
xor U57 (N_57,In_1618,In_290);
and U58 (N_58,In_1307,In_1510);
and U59 (N_59,In_689,In_88);
xnor U60 (N_60,In_60,In_524);
nand U61 (N_61,In_439,In_1044);
or U62 (N_62,In_53,In_594);
and U63 (N_63,In_1888,In_1961);
or U64 (N_64,In_1690,In_1495);
nor U65 (N_65,In_1270,In_1207);
or U66 (N_66,In_157,In_639);
or U67 (N_67,In_858,In_85);
and U68 (N_68,In_87,In_1798);
xor U69 (N_69,In_796,In_1670);
and U70 (N_70,In_1354,In_1114);
xnor U71 (N_71,In_505,In_1950);
or U72 (N_72,In_1477,In_275);
and U73 (N_73,In_1702,In_710);
and U74 (N_74,In_1186,In_1271);
and U75 (N_75,In_1141,In_1028);
nand U76 (N_76,In_167,In_440);
or U77 (N_77,In_1226,In_1345);
and U78 (N_78,In_1181,In_437);
nor U79 (N_79,In_1476,In_1802);
or U80 (N_80,In_1127,In_230);
or U81 (N_81,In_1760,In_1753);
nor U82 (N_82,In_1209,In_410);
or U83 (N_83,In_807,In_991);
or U84 (N_84,In_5,In_1573);
nand U85 (N_85,In_158,In_1064);
or U86 (N_86,In_1664,In_776);
or U87 (N_87,In_1929,In_458);
xor U88 (N_88,In_601,In_590);
nor U89 (N_89,In_1848,In_1933);
nor U90 (N_90,In_70,In_1159);
nand U91 (N_91,In_852,In_1656);
nand U92 (N_92,In_700,In_1998);
xnor U93 (N_93,In_441,In_1019);
nand U94 (N_94,In_1578,In_1692);
nor U95 (N_95,In_715,In_300);
nand U96 (N_96,In_864,In_1429);
xnor U97 (N_97,In_1743,In_224);
nor U98 (N_98,In_487,In_722);
xnor U99 (N_99,In_247,In_808);
and U100 (N_100,In_1053,In_674);
and U101 (N_101,In_266,In_1512);
and U102 (N_102,In_998,In_1568);
or U103 (N_103,In_217,In_638);
and U104 (N_104,In_714,In_1934);
and U105 (N_105,In_1938,In_1561);
or U106 (N_106,In_650,In_264);
or U107 (N_107,In_1917,In_297);
nand U108 (N_108,In_857,In_1111);
xnor U109 (N_109,In_469,In_571);
and U110 (N_110,In_949,In_67);
nor U111 (N_111,In_399,In_976);
xnor U112 (N_112,In_301,In_1310);
nand U113 (N_113,In_201,In_1800);
or U114 (N_114,In_740,In_1732);
xor U115 (N_115,In_1140,In_1080);
or U116 (N_116,In_890,In_1508);
xor U117 (N_117,In_1976,In_1660);
nor U118 (N_118,In_1543,In_344);
nand U119 (N_119,In_1597,In_1804);
or U120 (N_120,In_691,In_826);
nor U121 (N_121,In_599,In_385);
xnor U122 (N_122,In_1791,In_396);
nand U123 (N_123,In_726,In_1914);
nor U124 (N_124,In_234,In_1054);
nor U125 (N_125,In_1055,In_416);
xor U126 (N_126,In_83,In_1645);
and U127 (N_127,In_1427,In_1029);
and U128 (N_128,In_1306,In_1672);
nor U129 (N_129,In_869,In_267);
xnor U130 (N_130,In_403,In_731);
nor U131 (N_131,In_827,In_66);
xnor U132 (N_132,In_28,In_1750);
nor U133 (N_133,In_1870,In_921);
nor U134 (N_134,In_377,In_1363);
nor U135 (N_135,In_1110,In_1714);
nand U136 (N_136,In_1634,In_1815);
or U137 (N_137,In_1862,In_136);
and U138 (N_138,In_716,In_1567);
nor U139 (N_139,In_447,In_884);
or U140 (N_140,In_501,In_1416);
and U141 (N_141,In_149,In_1122);
and U142 (N_142,In_1986,In_1684);
xor U143 (N_143,In_842,In_521);
nor U144 (N_144,In_1774,In_617);
and U145 (N_145,In_367,In_55);
or U146 (N_146,In_54,In_384);
nor U147 (N_147,In_865,In_1903);
xnor U148 (N_148,In_549,In_1352);
and U149 (N_149,In_1553,In_958);
nand U150 (N_150,In_1440,In_333);
nor U151 (N_151,In_156,In_186);
nor U152 (N_152,In_678,In_231);
and U153 (N_153,In_1267,In_1148);
and U154 (N_154,In_308,In_1407);
or U155 (N_155,In_1892,In_1409);
nor U156 (N_156,In_1949,In_96);
nand U157 (N_157,In_1058,In_355);
nor U158 (N_158,In_1803,In_1844);
nor U159 (N_159,In_1169,In_1861);
and U160 (N_160,In_572,In_850);
nand U161 (N_161,In_1160,In_533);
xnor U162 (N_162,In_1269,In_1913);
and U163 (N_163,In_1355,In_1012);
and U164 (N_164,In_520,In_1017);
or U165 (N_165,In_288,In_916);
xnor U166 (N_166,In_1668,In_1577);
nor U167 (N_167,In_983,In_1653);
xnor U168 (N_168,In_1386,In_1663);
nand U169 (N_169,In_641,In_1439);
or U170 (N_170,In_1706,In_1241);
nand U171 (N_171,In_1430,In_368);
and U172 (N_172,In_925,In_1799);
and U173 (N_173,In_1935,In_1924);
and U174 (N_174,In_1651,In_509);
or U175 (N_175,In_1921,In_515);
xnor U176 (N_176,In_1304,In_672);
nor U177 (N_177,In_1829,In_6);
and U178 (N_178,In_35,In_174);
nand U179 (N_179,In_1387,In_1682);
xor U180 (N_180,In_107,In_1824);
or U181 (N_181,In_1371,In_1562);
nor U182 (N_182,In_123,In_33);
xnor U183 (N_183,In_1605,In_1649);
xor U184 (N_184,In_510,In_119);
or U185 (N_185,In_1112,In_398);
xor U186 (N_186,In_1052,In_1904);
xor U187 (N_187,In_1812,In_1822);
nand U188 (N_188,In_257,In_767);
and U189 (N_189,In_1835,In_241);
nand U190 (N_190,In_213,In_283);
nor U191 (N_191,In_1957,In_1853);
nand U192 (N_192,In_1324,In_1274);
or U193 (N_193,In_1225,In_1863);
nor U194 (N_194,In_887,In_1214);
and U195 (N_195,In_1166,In_1249);
and U196 (N_196,In_1780,In_1788);
or U197 (N_197,In_1722,In_1070);
nor U198 (N_198,In_1444,In_1588);
and U199 (N_199,In_774,In_1085);
xor U200 (N_200,In_1885,In_1833);
xnor U201 (N_201,In_584,In_880);
or U202 (N_202,In_1981,In_1593);
and U203 (N_203,In_114,In_1057);
and U204 (N_204,In_1704,In_434);
xnor U205 (N_205,In_331,In_777);
or U206 (N_206,In_1453,In_284);
nor U207 (N_207,In_159,In_340);
nand U208 (N_208,In_1224,In_728);
and U209 (N_209,In_1980,In_661);
and U210 (N_210,In_719,In_1479);
nor U211 (N_211,In_866,In_1051);
and U212 (N_212,In_304,In_751);
or U213 (N_213,In_1256,In_1627);
xnor U214 (N_214,In_687,In_578);
or U215 (N_215,In_815,In_313);
and U216 (N_216,In_369,In_1624);
nand U217 (N_217,In_124,In_554);
and U218 (N_218,In_1317,In_975);
nor U219 (N_219,In_1579,In_506);
nand U220 (N_220,In_604,In_907);
nor U221 (N_221,In_1107,In_688);
or U222 (N_222,In_812,In_321);
xnor U223 (N_223,In_1125,In_249);
nor U224 (N_224,In_536,In_932);
or U225 (N_225,In_670,In_915);
xor U226 (N_226,In_1100,In_1841);
xor U227 (N_227,In_937,In_1185);
nor U228 (N_228,In_1446,In_855);
or U229 (N_229,In_188,In_10);
nand U230 (N_230,In_1161,In_897);
or U231 (N_231,In_955,In_1556);
and U232 (N_232,In_644,In_1487);
nand U233 (N_233,In_694,In_820);
xnor U234 (N_234,In_1022,In_1557);
nand U235 (N_235,In_530,In_1323);
and U236 (N_236,In_1779,In_16);
or U237 (N_237,In_588,In_324);
xnor U238 (N_238,In_675,In_1088);
nand U239 (N_239,In_111,In_1548);
and U240 (N_240,In_773,In_1007);
nand U241 (N_241,In_1534,In_893);
and U242 (N_242,In_359,In_1197);
xnor U243 (N_243,In_580,In_1683);
and U244 (N_244,In_1717,In_1958);
xnor U245 (N_245,In_135,In_1840);
nor U246 (N_246,In_453,In_273);
xor U247 (N_247,In_172,In_127);
and U248 (N_248,In_1408,In_1425);
nand U249 (N_249,In_1852,In_31);
or U250 (N_250,In_1314,In_1813);
xor U251 (N_251,In_128,In_1368);
or U252 (N_252,In_1358,In_1308);
nand U253 (N_253,In_1655,In_951);
xnor U254 (N_254,In_1351,In_1689);
xor U255 (N_255,In_1074,In_1203);
or U256 (N_256,In_1817,In_1388);
nand U257 (N_257,In_1941,In_1895);
nand U258 (N_258,In_423,In_1631);
xnor U259 (N_259,In_495,In_1246);
and U260 (N_260,In_1887,In_1846);
nor U261 (N_261,In_115,In_473);
and U262 (N_262,In_1406,In_931);
or U263 (N_263,In_1983,In_593);
nor U264 (N_264,In_362,In_1766);
and U265 (N_265,In_965,In_1189);
xnor U266 (N_266,In_1486,In_1756);
nor U267 (N_267,In_323,In_248);
xnor U268 (N_268,In_1609,In_972);
and U269 (N_269,In_1994,In_1943);
or U270 (N_270,In_997,In_1681);
nor U271 (N_271,In_1469,In_30);
nor U272 (N_272,In_1454,In_1637);
and U273 (N_273,In_547,In_1737);
nand U274 (N_274,In_737,In_763);
or U275 (N_275,In_328,In_494);
xor U276 (N_276,In_529,In_1966);
xor U277 (N_277,In_435,In_1466);
or U278 (N_278,In_134,In_1715);
nor U279 (N_279,In_103,In_744);
or U280 (N_280,In_1176,In_1213);
nor U281 (N_281,In_252,In_225);
nand U282 (N_282,In_195,In_97);
and U283 (N_283,In_1874,In_1217);
xor U284 (N_284,In_303,In_392);
nand U285 (N_285,In_904,In_493);
or U286 (N_286,In_924,In_1020);
xor U287 (N_287,In_1826,In_1092);
or U288 (N_288,In_1626,In_1296);
nand U289 (N_289,In_51,In_838);
nor U290 (N_290,In_513,In_204);
nor U291 (N_291,In_1385,In_839);
nand U292 (N_292,In_235,In_1939);
or U293 (N_293,In_130,In_671);
and U294 (N_294,In_424,In_197);
xnor U295 (N_295,In_980,In_229);
and U296 (N_296,In_490,In_479);
nand U297 (N_297,In_1883,In_1922);
and U298 (N_298,In_243,In_1101);
nor U299 (N_299,In_1135,In_851);
or U300 (N_300,In_1792,In_1518);
nor U301 (N_301,In_1832,In_1794);
and U302 (N_302,In_208,In_1097);
nor U303 (N_303,In_1108,In_1030);
or U304 (N_304,In_1035,In_100);
and U305 (N_305,In_1928,In_1083);
nand U306 (N_306,In_787,In_995);
or U307 (N_307,In_1738,In_1496);
xnor U308 (N_308,In_553,In_1202);
and U309 (N_309,In_141,In_206);
nor U310 (N_310,In_786,In_1628);
nor U311 (N_311,In_486,In_364);
and U312 (N_312,In_1109,In_1441);
and U313 (N_313,In_163,In_1574);
and U314 (N_314,In_1311,In_1032);
xor U315 (N_315,In_1698,In_1396);
and U316 (N_316,In_795,In_560);
and U317 (N_317,In_1549,In_1900);
nor U318 (N_318,In_1081,In_1381);
xnor U319 (N_319,In_1184,In_745);
or U320 (N_320,In_1725,In_676);
xor U321 (N_321,In_61,In_1625);
and U322 (N_322,In_270,In_1608);
nand U323 (N_323,In_1232,In_346);
or U324 (N_324,In_293,In_155);
nor U325 (N_325,In_1350,In_1857);
or U326 (N_326,In_271,In_1544);
xnor U327 (N_327,In_1115,In_1819);
xnor U328 (N_328,In_1820,In_436);
or U329 (N_329,In_1586,In_1468);
xnor U330 (N_330,In_1517,In_1773);
or U331 (N_331,In_657,In_358);
and U332 (N_332,In_1010,In_17);
nor U333 (N_333,In_1560,In_142);
or U334 (N_334,In_1705,In_36);
xor U335 (N_335,In_1691,In_342);
nand U336 (N_336,In_1342,In_394);
xor U337 (N_337,In_1258,In_106);
nand U338 (N_338,In_939,In_189);
nand U339 (N_339,In_1179,In_1402);
xnor U340 (N_340,In_1757,In_1514);
and U341 (N_341,In_508,In_1398);
and U342 (N_342,In_1130,In_1944);
nand U343 (N_343,In_1940,In_977);
or U344 (N_344,In_666,In_1090);
or U345 (N_345,In_1891,In_1931);
xnor U346 (N_346,In_1361,In_782);
and U347 (N_347,In_899,In_605);
or U348 (N_348,In_905,In_1808);
xnor U349 (N_349,In_175,In_268);
or U350 (N_350,In_56,In_1783);
or U351 (N_351,In_811,In_1978);
xnor U352 (N_352,In_1971,In_1004);
nand U353 (N_353,In_1372,In_181);
xnor U354 (N_354,In_86,In_1373);
and U355 (N_355,In_772,In_1239);
nor U356 (N_356,In_545,In_1294);
or U357 (N_357,In_72,In_1318);
nor U358 (N_358,In_118,In_1893);
nand U359 (N_359,In_214,In_713);
and U360 (N_360,In_1945,In_1814);
nor U361 (N_361,In_1410,In_1733);
or U362 (N_362,In_1635,In_1867);
nand U363 (N_363,In_1460,In_1591);
nand U364 (N_364,In_761,In_1763);
or U365 (N_365,In_1098,In_1751);
xor U366 (N_366,In_129,In_121);
xnor U367 (N_367,In_665,In_1703);
xnor U368 (N_368,In_1828,In_298);
xnor U369 (N_369,In_1134,In_57);
nand U370 (N_370,In_280,In_352);
and U371 (N_371,In_25,In_563);
and U372 (N_372,In_1330,In_1218);
nand U373 (N_373,In_1995,In_1065);
and U374 (N_374,In_1089,In_988);
nand U375 (N_375,In_1724,In_809);
and U376 (N_376,In_282,In_37);
or U377 (N_377,In_34,In_612);
or U378 (N_378,In_783,In_1834);
and U379 (N_379,In_1009,In_372);
nor U380 (N_380,In_1143,In_1932);
xor U381 (N_381,In_27,In_1126);
nor U382 (N_382,In_860,In_1227);
or U383 (N_383,In_443,In_1333);
and U384 (N_384,In_1947,In_1005);
nand U385 (N_385,In_464,In_1752);
xnor U386 (N_386,In_642,In_959);
xnor U387 (N_387,In_1997,In_351);
and U388 (N_388,In_1580,In_994);
and U389 (N_389,In_1912,In_1901);
xor U390 (N_390,In_519,In_1216);
nand U391 (N_391,In_75,In_1585);
and U392 (N_392,In_1073,In_228);
nor U393 (N_393,In_1366,In_1419);
nand U394 (N_394,In_1379,In_244);
nand U395 (N_395,In_1478,In_828);
xor U396 (N_396,In_927,In_255);
nand U397 (N_397,In_758,In_32);
nand U398 (N_398,In_1540,In_373);
nor U399 (N_399,In_1347,In_272);
or U400 (N_400,In_1831,In_1927);
nand U401 (N_401,In_1699,In_68);
nand U402 (N_402,In_1719,In_1493);
xnor U403 (N_403,In_913,In_1375);
xor U404 (N_404,In_1335,In_859);
nand U405 (N_405,In_1583,In_942);
and U406 (N_406,In_566,In_1889);
or U407 (N_407,In_697,In_1288);
nor U408 (N_408,In_526,In_64);
and U409 (N_409,In_576,In_42);
and U410 (N_410,In_289,In_325);
and U411 (N_411,In_393,In_1069);
and U412 (N_412,In_1281,In_1162);
and U413 (N_413,In_548,In_1842);
or U414 (N_414,In_837,In_1973);
nor U415 (N_415,In_917,In_349);
nand U416 (N_416,In_381,In_404);
nor U417 (N_417,In_1930,In_628);
or U418 (N_418,In_1915,In_844);
nand U419 (N_419,In_1102,In_1328);
and U420 (N_420,In_1292,In_1124);
nand U421 (N_421,In_581,In_356);
nand U422 (N_422,In_1155,In_226);
or U423 (N_423,In_693,In_1067);
and U424 (N_424,In_662,In_1576);
and U425 (N_425,In_1401,In_1856);
nand U426 (N_426,In_1295,In_1303);
nand U427 (N_427,In_1911,In_1535);
xor U428 (N_428,In_1395,In_1721);
xor U429 (N_429,In_885,In_993);
nor U430 (N_430,In_339,In_1793);
or U431 (N_431,In_1880,In_1641);
nor U432 (N_432,In_113,In_1598);
nand U433 (N_433,In_749,In_1488);
and U434 (N_434,In_1536,In_1322);
nand U435 (N_435,In_1445,In_1767);
and U436 (N_436,In_418,In_296);
nor U437 (N_437,In_1150,In_698);
nor U438 (N_438,In_1123,In_621);
nor U439 (N_439,In_1099,In_1128);
xor U440 (N_440,In_684,In_1761);
nand U441 (N_441,In_1456,In_1886);
and U442 (N_442,In_1437,In_1190);
xor U443 (N_443,In_140,In_92);
nand U444 (N_444,In_1152,In_194);
or U445 (N_445,In_1899,In_1312);
nand U446 (N_446,In_1119,In_1242);
and U447 (N_447,In_81,In_173);
xor U448 (N_448,In_1622,In_825);
and U449 (N_449,In_1118,In_1484);
and U450 (N_450,In_1279,In_1718);
nand U451 (N_451,In_1147,In_953);
or U452 (N_452,In_1969,In_1093);
xnor U453 (N_453,In_1707,In_971);
xnor U454 (N_454,In_202,In_1254);
or U455 (N_455,In_1428,In_1277);
nor U456 (N_456,In_1731,In_836);
xor U457 (N_457,In_1376,In_190);
and U458 (N_458,In_798,In_867);
or U459 (N_459,In_1075,In_537);
nand U460 (N_460,In_912,In_1513);
or U461 (N_461,In_968,In_829);
and U462 (N_462,In_1500,In_1747);
or U463 (N_463,In_1063,In_1);
nand U464 (N_464,In_1422,In_791);
nand U465 (N_465,In_1275,In_1195);
or U466 (N_466,In_889,In_1606);
nand U467 (N_467,In_1178,In_841);
nor U468 (N_468,In_1391,In_1905);
nand U469 (N_469,In_1056,In_1979);
and U470 (N_470,In_1529,In_1730);
or U471 (N_471,In_1417,In_1483);
nand U472 (N_472,In_164,In_327);
nand U473 (N_473,In_507,In_870);
and U474 (N_474,In_1613,In_1248);
nand U475 (N_475,In_265,In_1482);
nor U476 (N_476,In_898,In_1956);
xor U477 (N_477,In_653,In_1229);
and U478 (N_478,In_360,In_861);
xnor U479 (N_479,In_1530,In_191);
and U480 (N_480,In_285,In_278);
or U481 (N_481,In_1764,In_1790);
and U482 (N_482,In_309,In_775);
xor U483 (N_483,In_1953,In_236);
nand U484 (N_484,In_1827,In_1984);
nor U485 (N_485,In_1091,In_451);
and U486 (N_486,In_1157,In_1411);
or U487 (N_487,In_770,In_1182);
xor U488 (N_488,In_1985,In_1629);
or U489 (N_489,In_1769,In_1854);
and U490 (N_490,In_794,In_1555);
nor U491 (N_491,In_1902,In_945);
xor U492 (N_492,In_1955,In_538);
and U493 (N_493,In_1532,In_161);
nor U494 (N_494,In_1652,In_19);
and U495 (N_495,In_835,In_422);
nand U496 (N_496,In_718,In_1859);
or U497 (N_497,In_375,In_540);
xnor U498 (N_498,In_1015,In_1866);
and U499 (N_499,In_1192,In_502);
nor U500 (N_500,In_198,N_475);
xnor U501 (N_501,N_173,N_102);
and U502 (N_502,N_235,In_944);
and U503 (N_503,In_1238,In_562);
nand U504 (N_504,N_110,N_177);
nand U505 (N_505,In_1972,In_1423);
and U506 (N_506,In_1650,In_822);
and U507 (N_507,In_1079,In_922);
xor U508 (N_508,N_402,N_129);
or U509 (N_509,N_489,In_1964);
xor U510 (N_510,In_1537,In_967);
and U511 (N_511,In_238,N_331);
and U512 (N_512,In_222,In_63);
nor U513 (N_513,In_1282,In_1785);
or U514 (N_514,In_1414,In_785);
or U515 (N_515,N_450,N_35);
xor U516 (N_516,In_1748,N_395);
nand U517 (N_517,In_748,N_77);
and U518 (N_518,In_281,N_435);
or U519 (N_519,In_251,In_908);
and U520 (N_520,In_735,N_262);
and U521 (N_521,In_543,N_307);
nor U522 (N_522,In_1616,N_399);
and U523 (N_523,N_100,In_1736);
or U524 (N_524,In_523,N_445);
xnor U525 (N_525,In_1204,In_534);
nand U526 (N_526,N_281,In_1611);
or U527 (N_527,In_1849,N_82);
or U528 (N_528,In_1462,In_1435);
xor U529 (N_529,In_1264,In_299);
nor U530 (N_530,In_1369,In_1084);
or U531 (N_531,In_894,In_1951);
and U532 (N_532,N_300,In_677);
or U533 (N_533,In_466,N_265);
nor U534 (N_534,In_1260,In_1448);
and U535 (N_535,In_431,In_1836);
nand U536 (N_536,In_65,In_1472);
xnor U537 (N_537,In_500,N_389);
and U538 (N_538,N_492,N_104);
or U539 (N_539,N_38,In_1338);
xnor U540 (N_540,In_21,N_365);
nand U541 (N_541,In_1559,In_615);
nand U542 (N_542,N_280,In_1405);
or U543 (N_543,In_1806,In_635);
and U544 (N_544,N_387,In_525);
nor U545 (N_545,N_473,In_91);
and U546 (N_546,In_909,In_648);
and U547 (N_547,In_472,N_125);
nand U548 (N_548,In_1042,N_459);
or U549 (N_549,N_205,In_1033);
and U550 (N_550,N_369,In_1049);
nand U551 (N_551,In_1072,In_1470);
nand U552 (N_552,In_611,N_426);
nand U553 (N_553,In_415,In_646);
xnor U554 (N_554,In_1390,In_1610);
or U555 (N_555,N_67,N_170);
nand U556 (N_556,In_527,In_1727);
nor U557 (N_557,N_135,In_778);
nand U558 (N_558,In_319,In_357);
nand U559 (N_559,In_765,In_986);
and U560 (N_560,N_119,In_444);
and U561 (N_561,In_582,In_169);
nand U562 (N_562,In_1603,In_354);
nor U563 (N_563,In_1309,N_403);
and U564 (N_564,N_5,In_1076);
or U565 (N_565,In_1475,In_420);
and U566 (N_566,In_261,In_1050);
nand U567 (N_567,In_1146,In_1302);
nor U568 (N_568,In_1382,N_449);
or U569 (N_569,N_360,N_305);
xor U570 (N_570,N_417,N_491);
nand U571 (N_571,In_1299,N_226);
and U572 (N_572,In_1397,In_317);
xnor U573 (N_573,N_284,In_608);
nand U574 (N_574,In_1673,In_1937);
or U575 (N_575,In_1250,N_263);
or U576 (N_576,In_1293,In_1908);
or U577 (N_577,N_33,N_26);
xnor U578 (N_578,N_471,N_164);
nand U579 (N_579,N_467,In_1116);
nand U580 (N_580,In_1952,N_255);
nor U581 (N_581,In_177,In_1661);
or U582 (N_582,In_1926,In_144);
nand U583 (N_583,In_8,N_422);
or U584 (N_584,In_433,N_394);
nor U585 (N_585,In_491,In_269);
or U586 (N_586,In_779,In_1851);
nand U587 (N_587,In_1208,In_879);
xnor U588 (N_588,N_409,N_434);
xnor U589 (N_589,In_1008,In_414);
and U590 (N_590,N_487,In_1421);
xnor U591 (N_591,N_151,N_314);
and U592 (N_592,In_1023,N_220);
or U593 (N_593,N_27,In_211);
nor U594 (N_594,N_57,In_1156);
nand U595 (N_595,In_1522,In_442);
xor U596 (N_596,In_73,In_948);
and U597 (N_597,In_183,In_1062);
or U598 (N_598,N_222,In_1301);
nor U599 (N_599,N_105,In_759);
xor U600 (N_600,In_1346,In_151);
nor U601 (N_601,In_1236,In_1403);
nand U602 (N_602,In_125,N_165);
nor U603 (N_603,N_115,In_1701);
nor U604 (N_604,In_848,N_29);
nand U605 (N_605,In_600,In_1497);
and U606 (N_606,N_283,In_1458);
nor U607 (N_607,N_246,In_854);
and U608 (N_608,In_834,N_248);
nand U609 (N_609,In_1400,In_48);
and U610 (N_610,In_330,In_1570);
nand U611 (N_611,N_109,In_58);
and U612 (N_612,In_148,In_564);
nand U613 (N_613,N_329,In_89);
and U614 (N_614,N_32,In_645);
and U615 (N_615,In_425,In_131);
xor U616 (N_616,In_692,In_363);
nor U617 (N_617,In_1321,In_1523);
or U618 (N_618,In_1918,N_204);
xor U619 (N_619,N_452,N_215);
nand U620 (N_620,In_1153,In_143);
nor U621 (N_621,N_159,In_999);
or U622 (N_622,In_101,In_93);
xnor U623 (N_623,N_495,N_274);
nand U624 (N_624,In_803,In_1433);
nand U625 (N_625,In_411,In_1671);
nor U626 (N_626,N_140,In_910);
xnor U627 (N_627,In_877,In_1261);
and U628 (N_628,In_1639,In_920);
or U629 (N_629,In_1873,In_1272);
and U630 (N_630,In_789,In_1078);
or U631 (N_631,N_146,In_1735);
nand U632 (N_632,In_957,N_406);
and U633 (N_633,In_1975,In_535);
or U634 (N_634,N_355,N_9);
nor U635 (N_635,In_314,In_1558);
or U636 (N_636,In_1511,In_518);
or U637 (N_637,N_128,N_260);
nand U638 (N_638,N_138,In_1545);
nor U639 (N_639,In_1463,In_1554);
xnor U640 (N_640,In_1744,N_377);
and U641 (N_641,N_212,In_237);
nor U642 (N_642,In_753,In_911);
nor U643 (N_643,In_934,N_267);
nand U644 (N_644,In_426,In_1480);
or U645 (N_645,In_1196,N_55);
nor U646 (N_646,In_277,N_181);
nand U647 (N_647,N_113,In_663);
nor U648 (N_648,In_1621,N_424);
and U649 (N_649,In_488,In_165);
nand U650 (N_650,In_77,In_484);
nand U651 (N_651,In_1337,In_1709);
or U652 (N_652,N_197,In_1129);
nand U653 (N_653,In_717,In_591);
or U654 (N_654,In_504,In_1452);
xnor U655 (N_655,In_489,In_1170);
nor U656 (N_656,In_1847,N_7);
or U657 (N_657,In_417,In_557);
and U658 (N_658,In_448,In_1739);
nor U659 (N_659,In_596,N_418);
xnor U660 (N_660,In_366,In_1038);
or U661 (N_661,In_764,In_542);
nor U662 (N_662,In_896,N_133);
nor U663 (N_663,N_12,In_445);
nand U664 (N_664,N_86,In_1855);
and U665 (N_665,In_1320,N_218);
and U666 (N_666,In_1644,In_651);
nand U667 (N_667,In_1315,In_45);
and U668 (N_668,In_1954,In_1755);
xor U669 (N_669,N_167,In_810);
xor U670 (N_670,In_145,N_321);
xor U671 (N_671,In_84,In_1602);
or U672 (N_672,In_246,In_485);
nand U673 (N_673,In_193,In_1158);
nand U674 (N_674,In_1640,In_1262);
and U675 (N_675,In_614,N_122);
xnor U676 (N_676,In_1716,N_60);
and U677 (N_677,N_14,N_397);
nand U678 (N_678,In_792,In_29);
nor U679 (N_679,N_411,In_79);
xor U680 (N_680,N_393,In_1669);
nand U681 (N_681,N_400,In_1244);
nor U682 (N_682,In_1823,In_819);
nor U683 (N_683,In_1890,N_462);
nand U684 (N_684,In_960,In_814);
and U685 (N_685,In_474,In_1749);
and U686 (N_686,In_1442,N_311);
nor U687 (N_687,In_632,In_1499);
or U688 (N_688,In_26,In_1464);
xnor U689 (N_689,In_1031,N_392);
nor U690 (N_690,N_493,In_1491);
and U691 (N_691,In_3,In_23);
nand U692 (N_692,In_205,In_1285);
or U693 (N_693,N_175,In_874);
and U694 (N_694,In_409,N_290);
xor U695 (N_695,In_1284,In_1498);
or U696 (N_696,In_685,In_402);
nor U697 (N_697,In_345,In_1667);
and U698 (N_698,In_556,In_1910);
and U699 (N_699,N_116,In_1786);
or U700 (N_700,N_323,In_568);
nor U701 (N_701,In_483,In_455);
xnor U702 (N_702,N_455,In_391);
or U703 (N_703,N_120,In_1237);
and U704 (N_704,In_1509,In_732);
nand U705 (N_705,N_453,In_480);
and U706 (N_706,In_613,In_199);
nor U707 (N_707,In_432,N_474);
nor U708 (N_708,In_681,In_1654);
or U709 (N_709,In_256,In_12);
xnor U710 (N_710,In_170,In_1230);
and U711 (N_711,N_276,N_420);
and U712 (N_712,In_1521,In_1047);
or U713 (N_713,In_1365,N_324);
or U714 (N_714,N_66,N_47);
xnor U715 (N_715,In_736,N_22);
xor U716 (N_716,N_132,N_483);
nor U717 (N_717,In_813,N_421);
or U718 (N_718,In_1925,N_21);
and U719 (N_719,In_406,In_1220);
nor U720 (N_720,In_741,N_432);
nand U721 (N_721,In_1370,In_1538);
nand U722 (N_722,In_69,In_847);
and U723 (N_723,In_1746,In_1377);
xor U724 (N_724,In_1393,N_101);
nand U725 (N_725,In_326,In_82);
nand U726 (N_726,In_1106,In_1503);
nor U727 (N_727,N_64,In_1843);
nor U728 (N_728,In_1201,N_240);
nor U729 (N_729,In_933,In_712);
nand U730 (N_730,N_210,In_311);
or U731 (N_731,In_647,In_147);
nand U732 (N_732,In_1006,N_349);
or U733 (N_733,In_1758,In_477);
nor U734 (N_734,N_20,In_1686);
nand U735 (N_735,N_43,In_781);
nor U736 (N_736,In_626,In_1977);
xor U737 (N_737,In_1520,In_1564);
and U738 (N_738,In_1187,In_1103);
or U739 (N_739,N_154,N_370);
and U740 (N_740,N_79,N_4);
nand U741 (N_741,In_292,In_603);
nand U742 (N_742,In_1617,In_1046);
and U743 (N_743,In_430,In_139);
nor U744 (N_744,In_1633,N_443);
or U745 (N_745,N_117,N_419);
nor U746 (N_746,In_1343,N_341);
nor U747 (N_747,In_1599,N_490);
xnor U748 (N_748,N_390,In_831);
nor U749 (N_749,In_1871,N_476);
or U750 (N_750,N_145,In_1959);
and U751 (N_751,N_427,In_76);
nor U752 (N_752,In_1876,N_373);
xnor U753 (N_753,In_13,In_219);
nor U754 (N_754,N_158,In_962);
nand U755 (N_755,In_168,N_96);
and U756 (N_756,N_106,In_1041);
nor U757 (N_757,N_81,In_1694);
and U758 (N_758,In_1257,In_1332);
or U759 (N_759,In_1131,N_203);
nor U760 (N_760,In_1210,In_496);
nor U761 (N_761,N_224,N_184);
xor U762 (N_762,In_370,N_383);
or U763 (N_763,In_1485,In_956);
or U764 (N_764,In_514,In_727);
nand U765 (N_765,In_1198,In_1970);
and U766 (N_766,N_404,In_701);
nand U767 (N_767,In_1678,In_337);
nor U768 (N_768,In_914,N_316);
xnor U769 (N_769,In_963,In_1745);
or U770 (N_770,In_1795,N_206);
or U771 (N_771,In_1604,In_1086);
nand U772 (N_772,In_964,In_895);
and U773 (N_773,In_1581,In_1974);
and U774 (N_774,In_1167,In_1313);
nor U775 (N_775,In_471,N_258);
nor U776 (N_776,N_454,N_249);
nor U777 (N_777,N_195,N_36);
nor U778 (N_778,In_133,In_274);
nand U779 (N_779,In_1461,In_365);
nand U780 (N_780,N_189,In_1027);
xor U781 (N_781,In_371,In_1601);
nor U782 (N_782,In_1572,In_1471);
nor U783 (N_783,N_478,In_1331);
xor U784 (N_784,In_1360,In_192);
nor U785 (N_785,In_1988,In_1325);
xnor U786 (N_786,N_352,In_1142);
or U787 (N_787,N_13,N_130);
and U788 (N_788,N_148,In_1326);
nand U789 (N_789,In_1154,N_437);
nor U790 (N_790,In_322,N_353);
or U791 (N_791,In_709,In_871);
or U792 (N_792,In_1546,In_146);
nand U793 (N_793,In_1096,N_208);
or U794 (N_794,N_58,In_649);
and U795 (N_795,In_1247,In_1223);
or U796 (N_796,In_512,In_1066);
xor U797 (N_797,In_1253,N_484);
or U798 (N_798,In_1729,N_259);
and U799 (N_799,In_1594,In_579);
xor U800 (N_800,N_465,In_1431);
nand U801 (N_801,In_633,In_1273);
and U802 (N_802,In_1838,In_180);
or U803 (N_803,In_941,N_303);
xor U804 (N_804,In_1222,In_1742);
and U805 (N_805,N_63,N_481);
and U806 (N_806,In_1596,In_619);
and U807 (N_807,N_90,In_379);
xor U808 (N_808,In_1942,In_295);
and U809 (N_809,N_375,In_232);
or U810 (N_810,In_50,N_335);
and U811 (N_811,In_881,N_433);
or U812 (N_812,In_1438,In_1340);
or U813 (N_813,In_724,In_1992);
and U814 (N_814,N_198,In_872);
nand U815 (N_815,In_1881,N_34);
xnor U816 (N_816,In_551,In_1920);
nor U817 (N_817,In_1566,In_821);
xor U818 (N_818,N_350,In_970);
and U819 (N_819,N_76,In_258);
nand U820 (N_820,In_492,N_23);
or U821 (N_821,N_144,In_766);
or U822 (N_822,In_62,N_28);
xor U823 (N_823,In_930,N_108);
or U824 (N_824,N_322,N_74);
nand U825 (N_825,In_1864,In_996);
xor U826 (N_826,In_1850,In_1188);
nor U827 (N_827,N_152,In_1199);
nor U828 (N_828,In_658,N_85);
nand U829 (N_829,In_1378,N_30);
nor U830 (N_830,In_886,In_1643);
xor U831 (N_831,In_1447,In_1095);
xor U832 (N_832,N_163,In_1542);
or U833 (N_833,In_294,In_1993);
and U834 (N_834,N_338,In_47);
or U835 (N_835,In_1240,In_1171);
nand U836 (N_836,N_61,N_87);
xnor U837 (N_837,N_201,In_1021);
nor U838 (N_838,In_1563,In_460);
xor U839 (N_839,In_1525,In_408);
nand U840 (N_840,In_900,N_447);
and U841 (N_841,In_1286,In_610);
and U842 (N_842,In_306,N_488);
and U843 (N_843,In_1389,In_15);
nor U844 (N_844,In_1193,In_978);
xnor U845 (N_845,N_269,N_71);
xnor U846 (N_846,In_1575,In_739);
xor U847 (N_847,In_1329,In_876);
and U848 (N_848,In_1459,N_200);
nor U849 (N_849,In_1420,In_74);
xor U850 (N_850,N_232,In_630);
nand U851 (N_851,N_84,In_723);
xnor U852 (N_852,N_112,In_1963);
and U853 (N_853,In_992,In_1865);
nand U854 (N_854,In_928,In_721);
and U855 (N_855,In_1434,In_1962);
nand U856 (N_856,N_41,In_350);
nand U857 (N_857,In_623,In_511);
xor U858 (N_858,In_1412,In_499);
or U859 (N_859,N_213,In_162);
xnor U860 (N_860,N_40,In_1235);
xnor U861 (N_861,In_892,In_1144);
nor U862 (N_862,In_574,In_4);
nor U863 (N_863,In_310,In_1163);
or U864 (N_864,In_585,In_388);
nor U865 (N_865,In_833,In_1426);
nor U866 (N_866,N_251,In_220);
and U867 (N_867,N_73,N_415);
or U868 (N_868,N_187,N_241);
nand U869 (N_869,In_806,In_720);
nand U870 (N_870,N_194,In_1845);
nor U871 (N_871,N_374,In_315);
or U872 (N_872,N_48,N_451);
nand U873 (N_873,N_219,In_1215);
or U874 (N_874,N_306,N_252);
or U875 (N_875,In_817,In_138);
nand U876 (N_876,N_8,N_428);
xor U877 (N_877,N_209,In_711);
xor U878 (N_878,In_498,In_577);
and U879 (N_879,In_215,In_329);
xnor U880 (N_880,N_380,In_1712);
and U881 (N_881,N_367,N_223);
or U882 (N_882,In_1968,In_1592);
nor U883 (N_883,In_1380,In_1149);
xnor U884 (N_884,N_239,In_598);
and U885 (N_885,N_257,In_686);
nand U886 (N_886,In_1860,N_327);
or U887 (N_887,In_1524,In_974);
xnor U888 (N_888,N_359,In_824);
nand U889 (N_889,In_1136,N_401);
nand U890 (N_890,In_1287,In_102);
nor U891 (N_891,N_330,In_696);
xnor U892 (N_892,In_1194,In_233);
nor U893 (N_893,N_356,In_631);
nand U894 (N_894,N_339,N_149);
and U895 (N_895,N_17,N_391);
nand U896 (N_896,In_1636,In_1251);
nand U897 (N_897,In_522,In_291);
and U898 (N_898,In_1344,In_1728);
nor U899 (N_899,N_264,In_1263);
and U900 (N_900,In_262,N_441);
nor U901 (N_901,In_1674,In_1289);
xor U902 (N_902,N_289,In_1474);
nand U903 (N_903,N_270,In_160);
xnor U904 (N_904,N_313,In_1987);
nand U905 (N_905,In_1457,N_310);
and U906 (N_906,In_1394,In_966);
or U907 (N_907,In_901,In_575);
or U908 (N_908,N_93,N_279);
or U909 (N_909,In_1765,N_496);
or U910 (N_910,In_756,In_428);
nand U911 (N_911,In_210,In_137);
nor U912 (N_912,In_1657,N_134);
and U913 (N_913,In_1936,In_1771);
or U914 (N_914,In_1697,In_1013);
nor U915 (N_915,N_221,N_340);
nand U916 (N_916,In_98,In_954);
and U917 (N_917,In_1117,In_528);
xor U918 (N_918,N_344,In_18);
nor U919 (N_919,In_706,N_89);
or U920 (N_920,In_1025,In_1077);
xor U921 (N_921,In_1589,In_1177);
nor U922 (N_922,N_413,In_347);
nor U923 (N_923,N_328,In_1245);
and U924 (N_924,In_738,In_1630);
and U925 (N_925,N_103,In_482);
and U926 (N_926,In_452,In_71);
or U927 (N_927,In_1168,N_436);
and U928 (N_928,N_245,In_1801);
nor U929 (N_929,In_1339,N_111);
nand U930 (N_930,N_461,N_282);
or U931 (N_931,N_302,N_498);
or U932 (N_932,N_72,In_1872);
nand U933 (N_933,In_1280,In_943);
nor U934 (N_934,In_429,In_1877);
nor U935 (N_935,In_558,N_179);
xor U936 (N_936,N_153,N_225);
nor U937 (N_937,In_784,N_334);
and U938 (N_938,N_59,N_31);
nand U939 (N_939,In_627,N_287);
nor U940 (N_940,In_1504,In_1255);
xor U941 (N_941,In_105,N_333);
and U942 (N_942,In_1451,N_286);
nor U943 (N_943,In_853,In_679);
or U944 (N_944,In_1659,In_1291);
or U945 (N_945,N_155,In_1948);
and U946 (N_946,In_1002,N_10);
or U947 (N_947,In_1492,In_1666);
nor U948 (N_948,In_656,In_449);
xor U949 (N_949,N_298,In_760);
and U950 (N_950,In_771,In_1060);
and U951 (N_951,N_114,N_444);
and U952 (N_952,In_1481,In_263);
xor U953 (N_953,In_407,N_168);
xor U954 (N_954,N_256,In_539);
xnor U955 (N_955,In_1206,In_816);
and U956 (N_956,In_386,In_622);
xor U957 (N_957,In_182,In_276);
nand U958 (N_958,In_1145,In_1221);
nand U959 (N_959,In_830,In_209);
xor U960 (N_960,N_143,In_804);
or U961 (N_961,In_989,In_919);
nand U962 (N_962,In_132,N_188);
nor U963 (N_963,N_336,In_517);
nand U964 (N_964,In_940,N_49);
and U965 (N_965,N_142,N_273);
xor U966 (N_966,N_361,In_1319);
and U967 (N_967,N_382,In_1283);
and U968 (N_968,In_1467,N_15);
nor U969 (N_969,N_458,N_343);
or U970 (N_970,In_625,N_396);
and U971 (N_971,In_1026,In_1582);
or U972 (N_972,In_655,In_587);
nand U973 (N_973,In_1205,In_1696);
xnor U974 (N_974,N_342,N_141);
or U975 (N_975,In_1810,In_573);
xor U976 (N_976,In_769,In_39);
and U977 (N_977,In_112,N_65);
or U978 (N_978,In_1642,In_680);
and U979 (N_979,In_1071,In_1436);
and U980 (N_980,In_126,N_479);
nor U981 (N_981,In_1036,N_364);
nand U982 (N_982,N_440,In_799);
nor U983 (N_983,In_595,N_278);
and U984 (N_984,N_243,N_25);
nor U985 (N_985,In_1139,N_44);
and U986 (N_986,N_228,N_160);
nand U987 (N_987,N_231,In_629);
xor U988 (N_988,N_39,In_746);
xor U989 (N_989,In_1830,In_1713);
xor U990 (N_990,N_381,N_412);
xnor U991 (N_991,In_1759,In_1527);
nand U992 (N_992,In_973,In_1392);
or U993 (N_993,In_1212,In_923);
nand U994 (N_994,In_602,N_192);
or U995 (N_995,In_1113,N_161);
nor U996 (N_996,N_95,In_1569);
nor U997 (N_997,N_174,In_873);
and U998 (N_998,In_207,In_99);
xnor U999 (N_999,N_236,In_318);
nand U1000 (N_1000,In_1781,N_169);
xnor U1001 (N_1001,In_788,N_176);
xnor U1002 (N_1002,N_946,In_383);
nor U1003 (N_1003,N_660,N_667);
and U1004 (N_1004,In_708,In_654);
and U1005 (N_1005,N_357,In_902);
nand U1006 (N_1006,N_557,In_104);
nor U1007 (N_1007,N_559,N_237);
or U1008 (N_1008,In_1183,In_843);
and U1009 (N_1009,In_730,N_199);
nand U1010 (N_1010,N_882,N_11);
or U1011 (N_1011,N_191,N_740);
nand U1012 (N_1012,N_940,N_362);
nand U1013 (N_1013,N_701,In_109);
nor U1014 (N_1014,N_836,N_351);
and U1015 (N_1015,N_577,In_704);
and U1016 (N_1016,N_91,N_150);
or U1017 (N_1017,N_196,N_319);
and U1018 (N_1018,N_642,In_400);
nor U1019 (N_1019,N_876,In_316);
xnor U1020 (N_1020,In_1231,N_960);
nand U1021 (N_1021,N_707,In_555);
or U1022 (N_1022,N_871,In_1165);
nor U1023 (N_1023,N_630,N_309);
and U1024 (N_1024,N_299,N_677);
and U1025 (N_1025,In_1675,N_885);
nand U1026 (N_1026,In_1180,N_234);
nand U1027 (N_1027,In_1878,N_570);
nand U1028 (N_1028,N_738,N_728);
nand U1029 (N_1029,N_875,N_581);
and U1030 (N_1030,N_632,N_556);
and U1031 (N_1031,N_366,In_1906);
nor U1032 (N_1032,N_229,In_725);
nor U1033 (N_1033,N_729,N_767);
nand U1034 (N_1034,N_514,In_1676);
or U1035 (N_1035,N_587,N_318);
xor U1036 (N_1036,In_395,N_725);
nand U1037 (N_1037,N_681,N_16);
nand U1038 (N_1038,In_985,N_346);
xnor U1039 (N_1039,N_863,N_752);
xor U1040 (N_1040,N_994,N_665);
xnor U1041 (N_1041,N_442,N_80);
and U1042 (N_1042,In_1191,N_506);
nor U1043 (N_1043,In_793,N_526);
xor U1044 (N_1044,N_523,In_185);
and U1045 (N_1045,In_1679,In_374);
xnor U1046 (N_1046,In_461,N_663);
xor U1047 (N_1047,N_860,N_136);
nor U1048 (N_1048,N_908,In_1219);
nand U1049 (N_1049,N_868,N_574);
nor U1050 (N_1050,In_387,N_470);
xnor U1051 (N_1051,N_690,N_631);
nand U1052 (N_1052,N_430,In_454);
or U1053 (N_1053,N_596,N_796);
nor U1054 (N_1054,N_710,N_572);
xnor U1055 (N_1055,In_1590,N_656);
nand U1056 (N_1056,N_233,In_1837);
and U1057 (N_1057,N_547,N_997);
nand U1058 (N_1058,In_532,N_627);
or U1059 (N_1059,In_1809,N_705);
xnor U1060 (N_1060,In_78,N_861);
nand U1061 (N_1061,N_943,N_919);
or U1062 (N_1062,In_961,In_570);
or U1063 (N_1063,N_758,N_671);
nor U1064 (N_1064,N_745,In_43);
xor U1065 (N_1065,N_765,In_1839);
xnor U1066 (N_1066,N_985,N_654);
or U1067 (N_1067,N_583,N_819);
or U1068 (N_1068,In_561,In_1882);
xnor U1069 (N_1069,N_612,N_884);
or U1070 (N_1070,In_38,N_854);
nand U1071 (N_1071,N_977,N_46);
and U1072 (N_1072,N_504,N_757);
or U1073 (N_1073,N_803,N_981);
nand U1074 (N_1074,N_576,N_931);
nand U1075 (N_1075,N_984,In_862);
and U1076 (N_1076,N_408,In_1797);
nand U1077 (N_1077,N_768,N_794);
nand U1078 (N_1078,In_755,In_888);
and U1079 (N_1079,In_11,N_680);
xor U1080 (N_1080,In_1506,N_567);
or U1081 (N_1081,N_550,N_247);
or U1082 (N_1082,N_737,N_802);
xor U1083 (N_1083,In_546,N_840);
xor U1084 (N_1084,In_153,N_524);
nor U1085 (N_1085,N_730,N_388);
and U1086 (N_1086,In_245,In_1415);
xnor U1087 (N_1087,In_312,In_336);
nor U1088 (N_1088,N_895,N_988);
and U1089 (N_1089,N_987,In_1300);
or U1090 (N_1090,N_512,In_1151);
and U1091 (N_1091,N_598,In_1687);
nand U1092 (N_1092,N_2,N_78);
nor U1093 (N_1093,In_1680,In_1336);
and U1094 (N_1094,In_378,N_719);
nand U1095 (N_1095,In_221,N_94);
or U1096 (N_1096,In_150,N_800);
nand U1097 (N_1097,N_894,In_1138);
nor U1098 (N_1098,In_1367,N_634);
nor U1099 (N_1099,N_372,N_762);
nand U1100 (N_1100,N_976,In_1174);
or U1101 (N_1101,N_963,N_472);
nor U1102 (N_1102,N_996,In_589);
or U1103 (N_1103,In_1754,In_768);
xor U1104 (N_1104,N_633,N_964);
xor U1105 (N_1105,In_845,N_121);
or U1106 (N_1106,N_614,N_909);
and U1107 (N_1107,N_957,N_805);
xor U1108 (N_1108,N_3,N_593);
or U1109 (N_1109,In_475,In_1334);
nor U1110 (N_1110,N_549,N_589);
or U1111 (N_1111,N_972,N_563);
nand U1112 (N_1112,In_790,In_1677);
nand U1113 (N_1113,In_1584,N_953);
and U1114 (N_1114,N_621,N_410);
nor U1115 (N_1115,N_786,N_670);
xnor U1116 (N_1116,N_922,N_851);
xor U1117 (N_1117,N_658,In_891);
nor U1118 (N_1118,In_20,N_613);
nand U1119 (N_1119,N_217,N_918);
or U1120 (N_1120,N_804,N_688);
nand U1121 (N_1121,In_936,N_254);
and U1122 (N_1122,N_485,N_822);
and U1123 (N_1123,N_749,N_466);
nor U1124 (N_1124,N_775,N_691);
and U1125 (N_1125,N_590,In_1327);
nor U1126 (N_1126,N_689,N_682);
nand U1127 (N_1127,N_571,In_1648);
or U1128 (N_1128,N_672,In_467);
xor U1129 (N_1129,N_891,N_68);
or U1130 (N_1130,N_182,N_864);
nand U1131 (N_1131,N_358,In_1043);
nor U1132 (N_1132,N_952,N_288);
nor U1133 (N_1133,N_275,N_354);
xor U1134 (N_1134,N_522,N_605);
nor U1135 (N_1135,In_801,N_501);
xor U1136 (N_1136,N_635,N_123);
nor U1137 (N_1137,In_1825,N_521);
nor U1138 (N_1138,In_94,In_1034);
nor U1139 (N_1139,In_1665,In_1541);
nand U1140 (N_1140,N_639,N_325);
or U1141 (N_1141,N_558,N_912);
or U1142 (N_1142,In_1061,N_900);
and U1143 (N_1143,In_1982,N_540);
nor U1144 (N_1144,N_890,N_833);
or U1145 (N_1145,In_227,N_845);
nand U1146 (N_1146,N_772,N_544);
xnor U1147 (N_1147,N_457,N_754);
and U1148 (N_1148,N_995,N_675);
nand U1149 (N_1149,N_292,In_397);
or U1150 (N_1150,N_883,In_332);
nor U1151 (N_1151,In_1539,In_1432);
nor U1152 (N_1152,In_1364,N_867);
or U1153 (N_1153,In_1723,N_42);
or U1154 (N_1154,N_830,N_185);
nor U1155 (N_1155,N_539,N_733);
nor U1156 (N_1156,N_892,In_463);
xor U1157 (N_1157,N_56,In_660);
xor U1158 (N_1158,N_178,N_546);
nand U1159 (N_1159,N_849,In_950);
and U1160 (N_1160,N_156,N_520);
nand U1161 (N_1161,N_835,N_676);
nor U1162 (N_1162,In_938,N_817);
and U1163 (N_1163,In_1356,In_179);
nor U1164 (N_1164,In_1960,In_1515);
xnor U1165 (N_1165,N_643,N_950);
nand U1166 (N_1166,In_935,N_131);
xnor U1167 (N_1167,N_207,N_368);
nand U1168 (N_1168,In_187,N_425);
nor U1169 (N_1169,N_935,N_238);
and U1170 (N_1170,N_304,In_1897);
nand U1171 (N_1171,In_80,In_1418);
nor U1172 (N_1172,N_899,In_1505);
or U1173 (N_1173,N_893,In_1413);
or U1174 (N_1174,N_617,N_575);
xnor U1175 (N_1175,In_450,N_527);
nor U1176 (N_1176,N_948,N_717);
xnor U1177 (N_1177,N_536,In_1341);
nand U1178 (N_1178,In_438,N_770);
and U1179 (N_1179,N_75,N_959);
nor U1180 (N_1180,N_456,N_916);
nor U1181 (N_1181,In_1349,N_715);
xnor U1182 (N_1182,In_1473,In_1919);
or U1183 (N_1183,N_748,In_41);
nand U1184 (N_1184,In_1362,In_178);
xnor U1185 (N_1185,N_315,In_1646);
nand U1186 (N_1186,In_456,N_933);
or U1187 (N_1187,N_647,N_934);
xnor U1188 (N_1188,N_743,In_1720);
xnor U1189 (N_1189,N_271,N_911);
nand U1190 (N_1190,N_983,N_921);
or U1191 (N_1191,N_846,N_573);
nand U1192 (N_1192,N_242,N_664);
nor U1193 (N_1193,In_1711,N_505);
or U1194 (N_1194,N_162,N_961);
or U1195 (N_1195,N_942,In_1024);
or U1196 (N_1196,In_152,N_702);
or U1197 (N_1197,In_1133,N_568);
xor U1198 (N_1198,N_620,In_1619);
or U1199 (N_1199,N_530,In_868);
nand U1200 (N_1200,N_820,N_734);
or U1201 (N_1201,N_180,N_808);
and U1202 (N_1202,N_70,N_301);
nand U1203 (N_1203,N_930,N_166);
and U1204 (N_1204,N_69,N_713);
nand U1205 (N_1205,In_343,N_517);
xor U1206 (N_1206,N_732,In_1278);
and U1207 (N_1207,In_49,N_494);
or U1208 (N_1208,N_525,N_293);
nor U1209 (N_1209,In_1465,N_756);
nand U1210 (N_1210,In_1909,N_986);
xor U1211 (N_1211,In_7,In_544);
nand U1212 (N_1212,N_692,N_782);
nand U1213 (N_1213,In_446,In_878);
nand U1214 (N_1214,N_739,N_543);
xor U1215 (N_1215,N_929,In_95);
nor U1216 (N_1216,N_463,N_807);
nand U1217 (N_1217,N_889,N_761);
xor U1218 (N_1218,N_312,N_880);
nand U1219 (N_1219,N_781,N_566);
nor U1220 (N_1220,N_975,In_567);
nor U1221 (N_1221,N_460,In_1164);
nand U1222 (N_1222,In_1777,In_1316);
or U1223 (N_1223,N_939,N_641);
nand U1224 (N_1224,In_1211,N_597);
nand U1225 (N_1225,In_659,In_1501);
xor U1226 (N_1226,In_1132,N_956);
or U1227 (N_1227,N_727,In_1455);
and U1228 (N_1228,N_515,N_50);
xnor U1229 (N_1229,In_802,N_53);
or U1230 (N_1230,N_619,N_962);
nor U1231 (N_1231,In_46,In_1768);
nor U1232 (N_1232,N_423,N_780);
and U1233 (N_1233,In_286,N_838);
and U1234 (N_1234,In_1547,In_1297);
nand U1235 (N_1235,N_541,N_858);
xnor U1236 (N_1236,N_777,N_947);
or U1237 (N_1237,N_706,N_850);
xor U1238 (N_1238,N_230,N_98);
or U1239 (N_1239,N_771,N_897);
nor U1240 (N_1240,N_628,N_764);
nand U1241 (N_1241,N_62,In_1595);
or U1242 (N_1242,In_1531,In_503);
or U1243 (N_1243,In_1533,In_952);
and U1244 (N_1244,In_982,N_595);
nand U1245 (N_1245,N_945,N_801);
or U1246 (N_1246,N_712,N_827);
or U1247 (N_1247,N_296,In_1879);
nor U1248 (N_1248,In_1778,In_176);
or U1249 (N_1249,N_971,N_936);
or U1250 (N_1250,N_915,N_266);
nor U1251 (N_1251,In_846,In_462);
nand U1252 (N_1252,N_295,N_1);
xnor U1253 (N_1253,N_439,N_704);
xor U1254 (N_1254,N_924,N_659);
or U1255 (N_1255,In_184,In_690);
nor U1256 (N_1256,N_797,In_335);
or U1257 (N_1257,In_918,N_464);
xnor U1258 (N_1258,N_839,N_652);
nor U1259 (N_1259,N_385,In_1048);
nand U1260 (N_1260,In_1552,In_583);
xnor U1261 (N_1261,In_742,N_651);
nor U1262 (N_1262,In_1449,N_966);
xor U1263 (N_1263,In_1045,N_186);
nor U1264 (N_1264,N_773,N_949);
nor U1265 (N_1265,N_308,N_347);
nor U1266 (N_1266,N_431,N_793);
nor U1267 (N_1267,N_999,N_855);
and U1268 (N_1268,N_856,N_332);
xor U1269 (N_1269,N_500,In_682);
nor U1270 (N_1270,N_52,In_856);
nand U1271 (N_1271,In_1305,N_906);
and U1272 (N_1272,N_511,N_967);
and U1273 (N_1273,N_973,N_611);
nand U1274 (N_1274,N_363,N_227);
or U1275 (N_1275,N_508,In_218);
xnor U1276 (N_1276,N_533,In_702);
xnor U1277 (N_1277,N_811,N_602);
nand U1278 (N_1278,N_716,N_684);
xnor U1279 (N_1279,In_44,N_553);
nand U1280 (N_1280,N_560,N_244);
or U1281 (N_1281,N_37,N_790);
and U1282 (N_1282,N_731,In_1082);
nor U1283 (N_1283,N_376,N_700);
nand U1284 (N_1284,N_905,N_584);
xor U1285 (N_1285,N_594,N_0);
nand U1286 (N_1286,In_1734,N_592);
nor U1287 (N_1287,N_147,N_193);
nand U1288 (N_1288,In_1348,N_545);
and U1289 (N_1289,In_620,In_984);
and U1290 (N_1290,In_376,In_734);
or U1291 (N_1291,In_1565,In_1868);
or U1292 (N_1292,N_591,N_958);
xnor U1293 (N_1293,N_898,N_720);
or U1294 (N_1294,In_1607,N_297);
nand U1295 (N_1295,In_1740,N_416);
xnor U1296 (N_1296,N_923,N_92);
or U1297 (N_1297,In_643,In_305);
nor U1298 (N_1298,N_644,In_695);
or U1299 (N_1299,In_476,N_853);
nor U1300 (N_1300,N_814,In_405);
or U1301 (N_1301,In_1175,In_459);
or U1302 (N_1302,N_653,N_751);
nor U1303 (N_1303,N_928,In_1776);
nand U1304 (N_1304,N_862,N_879);
or U1305 (N_1305,N_607,N_171);
and U1306 (N_1306,N_914,In_478);
nor U1307 (N_1307,In_40,In_1923);
nor U1308 (N_1308,N_991,N_414);
and U1309 (N_1309,In_1243,N_588);
or U1310 (N_1310,N_857,N_623);
nor U1311 (N_1311,N_784,In_729);
xor U1312 (N_1312,N_534,N_873);
or U1313 (N_1313,In_341,N_379);
and U1314 (N_1314,N_645,In_0);
nand U1315 (N_1315,In_52,N_429);
or U1316 (N_1316,N_859,N_678);
xnor U1317 (N_1317,N_139,In_108);
or U1318 (N_1318,N_448,N_726);
xor U1319 (N_1319,N_778,N_917);
nand U1320 (N_1320,N_649,N_552);
or U1321 (N_1321,In_1989,In_1173);
or U1322 (N_1322,N_721,In_1770);
nor U1323 (N_1323,N_708,N_696);
or U1324 (N_1324,N_982,In_762);
and U1325 (N_1325,N_97,N_637);
xnor U1326 (N_1326,In_1612,In_703);
nand U1327 (N_1327,N_766,N_990);
nand U1328 (N_1328,In_1550,N_565);
xnor U1329 (N_1329,N_735,N_887);
nand U1330 (N_1330,N_600,N_190);
xor U1331 (N_1331,N_842,N_736);
xor U1332 (N_1332,In_259,In_389);
or U1333 (N_1333,N_913,N_538);
xnor U1334 (N_1334,In_250,N_268);
nor U1335 (N_1335,N_674,N_686);
and U1336 (N_1336,In_597,N_211);
nand U1337 (N_1337,In_1357,N_548);
xor U1338 (N_1338,In_1384,N_798);
nand U1339 (N_1339,N_697,N_769);
and U1340 (N_1340,N_841,N_137);
xor U1341 (N_1341,N_723,In_1290);
or U1342 (N_1342,N_468,N_486);
or U1343 (N_1343,In_823,N_699);
and U1344 (N_1344,In_1858,In_1916);
nand U1345 (N_1345,N_679,In_565);
or U1346 (N_1346,N_992,N_562);
or U1347 (N_1347,N_750,N_795);
nand U1348 (N_1348,N_818,N_789);
or U1349 (N_1349,N_202,N_384);
xnor U1350 (N_1350,N_126,N_722);
and U1351 (N_1351,N_469,N_847);
xnor U1352 (N_1352,N_657,N_989);
nand U1353 (N_1353,In_1137,N_510);
or U1354 (N_1354,N_622,N_54);
xor U1355 (N_1355,N_519,N_926);
and U1356 (N_1356,N_941,In_1991);
or U1357 (N_1357,In_1894,N_760);
or U1358 (N_1358,In_634,N_127);
and U1359 (N_1359,In_401,N_446);
or U1360 (N_1360,N_499,In_203);
xor U1361 (N_1361,N_809,N_601);
nor U1362 (N_1362,N_993,N_998);
nand U1363 (N_1363,In_800,In_1087);
xnor U1364 (N_1364,N_834,In_1875);
nand U1365 (N_1365,N_865,N_172);
nand U1366 (N_1366,N_610,In_470);
and U1367 (N_1367,N_604,N_537);
xor U1368 (N_1368,N_714,In_1359);
nor U1369 (N_1369,N_874,N_901);
xor U1370 (N_1370,N_759,N_407);
nor U1371 (N_1371,N_683,N_616);
and U1372 (N_1372,N_650,In_24);
nand U1373 (N_1373,N_693,In_780);
nor U1374 (N_1374,In_1772,In_840);
or U1375 (N_1375,N_955,In_117);
and U1376 (N_1376,In_1399,N_638);
and U1377 (N_1377,N_744,N_18);
or U1378 (N_1378,N_685,N_636);
and U1379 (N_1379,N_107,In_1172);
or U1380 (N_1380,In_883,N_640);
nand U1381 (N_1381,N_477,N_261);
xor U1382 (N_1382,In_254,In_154);
xnor U1383 (N_1383,In_743,In_1869);
and U1384 (N_1384,N_816,N_45);
xnor U1385 (N_1385,N_666,N_815);
and U1386 (N_1386,N_497,In_624);
nor U1387 (N_1387,N_599,N_618);
nand U1388 (N_1388,N_535,N_348);
xor U1389 (N_1389,In_1494,In_757);
nor U1390 (N_1390,In_279,N_969);
and U1391 (N_1391,N_954,In_586);
and U1392 (N_1392,In_465,N_19);
or U1393 (N_1393,N_24,N_746);
and U1394 (N_1394,N_832,N_799);
nor U1395 (N_1395,N_779,N_774);
nor U1396 (N_1396,N_509,In_1507);
nand U1397 (N_1397,N_157,N_337);
and U1398 (N_1398,N_903,In_1693);
xor U1399 (N_1399,N_886,N_551);
or U1400 (N_1400,N_648,N_405);
or U1401 (N_1401,N_965,N_698);
nand U1402 (N_1402,N_531,In_14);
and U1403 (N_1403,N_371,In_1632);
nor U1404 (N_1404,N_277,In_287);
nand U1405 (N_1405,In_1784,In_122);
and U1406 (N_1406,In_334,In_1884);
xnor U1407 (N_1407,N_582,N_763);
or U1408 (N_1408,N_844,N_831);
nor U1409 (N_1409,N_979,N_386);
xnor U1410 (N_1410,N_944,N_585);
nor U1411 (N_1411,N_787,In_1571);
nor U1412 (N_1412,In_1551,N_99);
and U1413 (N_1413,N_829,N_561);
nand U1414 (N_1414,N_978,N_951);
nor U1415 (N_1415,N_980,In_752);
nand U1416 (N_1416,N_272,In_640);
and U1417 (N_1417,N_826,N_253);
nand U1418 (N_1418,N_555,In_239);
nor U1419 (N_1419,N_124,N_669);
or U1420 (N_1420,In_320,N_542);
nand U1421 (N_1421,N_378,N_866);
xor U1422 (N_1422,In_541,N_937);
nand U1423 (N_1423,N_848,In_1266);
nand U1424 (N_1424,N_83,N_755);
nor U1425 (N_1425,In_981,N_872);
xnor U1426 (N_1426,In_468,N_825);
nor U1427 (N_1427,N_516,N_662);
nand U1428 (N_1428,In_979,In_1200);
nand U1429 (N_1429,N_294,N_564);
or U1430 (N_1430,N_938,N_503);
or U1431 (N_1431,N_927,N_285);
and U1432 (N_1432,In_805,N_974);
or U1433 (N_1433,N_896,N_877);
xor U1434 (N_1434,N_824,N_709);
or U1435 (N_1435,N_606,N_788);
nand U1436 (N_1436,In_616,N_673);
or U1437 (N_1437,In_1967,In_413);
nor U1438 (N_1438,In_22,N_502);
or U1439 (N_1439,In_747,In_906);
xor U1440 (N_1440,In_618,N_88);
or U1441 (N_1441,In_1762,In_516);
or U1442 (N_1442,N_806,N_747);
or U1443 (N_1443,In_1001,N_532);
nand U1444 (N_1444,N_742,In_196);
or U1445 (N_1445,In_1662,N_625);
nand U1446 (N_1446,N_783,N_326);
nor U1447 (N_1447,N_580,In_421);
nand U1448 (N_1448,N_785,N_813);
and U1449 (N_1449,In_1490,N_608);
nor U1450 (N_1450,N_925,In_1059);
and U1451 (N_1451,N_480,N_317);
nand U1452 (N_1452,In_669,N_518);
nor U1453 (N_1453,In_818,N_554);
nand U1454 (N_1454,N_646,In_1946);
xor U1455 (N_1455,In_531,In_1816);
nand U1456 (N_1456,N_823,N_843);
or U1457 (N_1457,In_903,N_624);
and U1458 (N_1458,N_703,N_920);
xor U1459 (N_1459,N_216,In_1811);
and U1460 (N_1460,N_852,N_694);
nor U1461 (N_1461,N_881,N_661);
and U1462 (N_1462,N_741,N_250);
nor U1463 (N_1463,In_1907,N_51);
or U1464 (N_1464,N_291,N_615);
nand U1465 (N_1465,N_320,N_6);
xor U1466 (N_1466,N_655,N_812);
xor U1467 (N_1467,N_724,In_497);
and U1468 (N_1468,N_668,N_482);
nand U1469 (N_1469,N_569,N_837);
nor U1470 (N_1470,In_668,N_910);
nor U1471 (N_1471,N_687,In_1796);
or U1472 (N_1472,N_578,N_513);
xnor U1473 (N_1473,N_695,In_699);
or U1474 (N_1474,N_711,N_603);
nor U1475 (N_1475,In_990,N_529);
nand U1476 (N_1476,In_926,N_902);
nand U1477 (N_1477,In_1234,N_753);
nand U1478 (N_1478,In_552,N_792);
or U1479 (N_1479,N_345,In_569);
and U1480 (N_1480,N_398,N_904);
or U1481 (N_1481,N_609,N_888);
nand U1482 (N_1482,N_810,N_791);
nor U1483 (N_1483,N_528,In_166);
and U1484 (N_1484,In_637,N_821);
nor U1485 (N_1485,In_882,In_1040);
and U1486 (N_1486,In_1775,N_626);
nor U1487 (N_1487,In_733,In_1120);
and U1488 (N_1488,In_797,In_302);
and U1489 (N_1489,N_869,N_776);
nand U1490 (N_1490,In_1821,N_932);
nand U1491 (N_1491,In_1658,N_968);
xor U1492 (N_1492,N_579,N_870);
and U1493 (N_1493,N_907,N_878);
nor U1494 (N_1494,N_214,In_1094);
xor U1495 (N_1495,N_718,N_507);
or U1496 (N_1496,N_629,N_586);
and U1497 (N_1497,N_118,N_828);
or U1498 (N_1498,N_183,In_1614);
xor U1499 (N_1499,N_970,N_438);
xor U1500 (N_1500,N_1486,N_1345);
xnor U1501 (N_1501,N_1427,N_1296);
nand U1502 (N_1502,N_1022,N_1484);
nor U1503 (N_1503,N_1147,N_1247);
and U1504 (N_1504,N_1050,N_1242);
xnor U1505 (N_1505,N_1420,N_1160);
and U1506 (N_1506,N_1360,N_1034);
and U1507 (N_1507,N_1409,N_1112);
xor U1508 (N_1508,N_1304,N_1004);
and U1509 (N_1509,N_1488,N_1104);
and U1510 (N_1510,N_1070,N_1415);
xor U1511 (N_1511,N_1211,N_1074);
nand U1512 (N_1512,N_1191,N_1081);
or U1513 (N_1513,N_1079,N_1480);
or U1514 (N_1514,N_1161,N_1435);
xnor U1515 (N_1515,N_1390,N_1493);
nand U1516 (N_1516,N_1338,N_1349);
or U1517 (N_1517,N_1392,N_1008);
xor U1518 (N_1518,N_1019,N_1379);
or U1519 (N_1519,N_1496,N_1295);
nand U1520 (N_1520,N_1031,N_1416);
or U1521 (N_1521,N_1120,N_1389);
nand U1522 (N_1522,N_1264,N_1281);
nor U1523 (N_1523,N_1271,N_1422);
and U1524 (N_1524,N_1378,N_1298);
and U1525 (N_1525,N_1197,N_1046);
xor U1526 (N_1526,N_1066,N_1325);
nor U1527 (N_1527,N_1470,N_1413);
nor U1528 (N_1528,N_1340,N_1241);
xnor U1529 (N_1529,N_1218,N_1494);
nor U1530 (N_1530,N_1381,N_1425);
nor U1531 (N_1531,N_1274,N_1351);
or U1532 (N_1532,N_1092,N_1491);
and U1533 (N_1533,N_1370,N_1439);
and U1534 (N_1534,N_1299,N_1164);
nor U1535 (N_1535,N_1387,N_1430);
or U1536 (N_1536,N_1321,N_1253);
or U1537 (N_1537,N_1169,N_1256);
xor U1538 (N_1538,N_1414,N_1015);
or U1539 (N_1539,N_1216,N_1097);
nand U1540 (N_1540,N_1053,N_1106);
and U1541 (N_1541,N_1438,N_1399);
xnor U1542 (N_1542,N_1385,N_1442);
and U1543 (N_1543,N_1145,N_1018);
nand U1544 (N_1544,N_1263,N_1189);
and U1545 (N_1545,N_1013,N_1434);
and U1546 (N_1546,N_1003,N_1306);
and U1547 (N_1547,N_1344,N_1005);
nor U1548 (N_1548,N_1375,N_1071);
nand U1549 (N_1549,N_1251,N_1115);
nor U1550 (N_1550,N_1465,N_1291);
or U1551 (N_1551,N_1431,N_1463);
nand U1552 (N_1552,N_1180,N_1236);
and U1553 (N_1553,N_1178,N_1181);
xnor U1554 (N_1554,N_1286,N_1101);
and U1555 (N_1555,N_1208,N_1064);
nand U1556 (N_1556,N_1275,N_1453);
and U1557 (N_1557,N_1045,N_1175);
xnor U1558 (N_1558,N_1123,N_1204);
nor U1559 (N_1559,N_1130,N_1094);
xnor U1560 (N_1560,N_1300,N_1258);
or U1561 (N_1561,N_1010,N_1479);
and U1562 (N_1562,N_1358,N_1400);
or U1563 (N_1563,N_1449,N_1477);
nor U1564 (N_1564,N_1394,N_1002);
nand U1565 (N_1565,N_1380,N_1355);
or U1566 (N_1566,N_1194,N_1309);
nand U1567 (N_1567,N_1121,N_1026);
xor U1568 (N_1568,N_1052,N_1265);
and U1569 (N_1569,N_1199,N_1012);
nor U1570 (N_1570,N_1095,N_1323);
or U1571 (N_1571,N_1047,N_1077);
nand U1572 (N_1572,N_1224,N_1410);
nor U1573 (N_1573,N_1317,N_1198);
or U1574 (N_1574,N_1332,N_1156);
xor U1575 (N_1575,N_1343,N_1455);
or U1576 (N_1576,N_1452,N_1411);
xor U1577 (N_1577,N_1244,N_1214);
nor U1578 (N_1578,N_1327,N_1170);
nor U1579 (N_1579,N_1049,N_1469);
or U1580 (N_1580,N_1402,N_1267);
and U1581 (N_1581,N_1361,N_1372);
nand U1582 (N_1582,N_1011,N_1226);
and U1583 (N_1583,N_1280,N_1168);
and U1584 (N_1584,N_1472,N_1294);
and U1585 (N_1585,N_1466,N_1030);
nor U1586 (N_1586,N_1468,N_1292);
and U1587 (N_1587,N_1122,N_1137);
or U1588 (N_1588,N_1219,N_1276);
and U1589 (N_1589,N_1210,N_1157);
nand U1590 (N_1590,N_1404,N_1179);
or U1591 (N_1591,N_1406,N_1068);
or U1592 (N_1592,N_1350,N_1405);
nor U1593 (N_1593,N_1313,N_1141);
and U1594 (N_1594,N_1132,N_1129);
xnor U1595 (N_1595,N_1475,N_1329);
or U1596 (N_1596,N_1090,N_1273);
nand U1597 (N_1597,N_1039,N_1305);
nor U1598 (N_1598,N_1205,N_1100);
or U1599 (N_1599,N_1203,N_1188);
xor U1600 (N_1600,N_1110,N_1445);
and U1601 (N_1601,N_1383,N_1467);
and U1602 (N_1602,N_1352,N_1283);
or U1603 (N_1603,N_1202,N_1301);
nand U1604 (N_1604,N_1419,N_1240);
and U1605 (N_1605,N_1232,N_1474);
or U1606 (N_1606,N_1159,N_1221);
or U1607 (N_1607,N_1213,N_1073);
nor U1608 (N_1608,N_1368,N_1333);
and U1609 (N_1609,N_1348,N_1084);
and U1610 (N_1610,N_1393,N_1423);
xor U1611 (N_1611,N_1401,N_1353);
and U1612 (N_1612,N_1143,N_1284);
or U1613 (N_1613,N_1458,N_1040);
nand U1614 (N_1614,N_1408,N_1036);
nand U1615 (N_1615,N_1109,N_1282);
and U1616 (N_1616,N_1476,N_1193);
nand U1617 (N_1617,N_1376,N_1089);
nor U1618 (N_1618,N_1029,N_1293);
nor U1619 (N_1619,N_1302,N_1076);
and U1620 (N_1620,N_1136,N_1154);
nor U1621 (N_1621,N_1262,N_1055);
nand U1622 (N_1622,N_1007,N_1058);
and U1623 (N_1623,N_1020,N_1139);
and U1624 (N_1624,N_1266,N_1043);
or U1625 (N_1625,N_1478,N_1080);
and U1626 (N_1626,N_1142,N_1063);
and U1627 (N_1627,N_1364,N_1146);
and U1628 (N_1628,N_1495,N_1217);
nor U1629 (N_1629,N_1114,N_1057);
nor U1630 (N_1630,N_1354,N_1497);
xnor U1631 (N_1631,N_1174,N_1303);
nor U1632 (N_1632,N_1127,N_1314);
xor U1633 (N_1633,N_1326,N_1315);
and U1634 (N_1634,N_1421,N_1287);
nor U1635 (N_1635,N_1395,N_1085);
nand U1636 (N_1636,N_1492,N_1021);
nor U1637 (N_1637,N_1482,N_1065);
xor U1638 (N_1638,N_1148,N_1384);
and U1639 (N_1639,N_1183,N_1185);
nor U1640 (N_1640,N_1386,N_1102);
nor U1641 (N_1641,N_1254,N_1398);
or U1642 (N_1642,N_1206,N_1324);
nand U1643 (N_1643,N_1374,N_1172);
nand U1644 (N_1644,N_1086,N_1196);
and U1645 (N_1645,N_1319,N_1418);
nor U1646 (N_1646,N_1245,N_1075);
nand U1647 (N_1647,N_1403,N_1116);
nand U1648 (N_1648,N_1464,N_1243);
nand U1649 (N_1649,N_1187,N_1330);
nor U1650 (N_1650,N_1457,N_1190);
and U1651 (N_1651,N_1429,N_1083);
xor U1652 (N_1652,N_1288,N_1237);
nand U1653 (N_1653,N_1006,N_1252);
and U1654 (N_1654,N_1437,N_1220);
xor U1655 (N_1655,N_1072,N_1270);
nor U1656 (N_1656,N_1487,N_1250);
xor U1657 (N_1657,N_1407,N_1311);
or U1658 (N_1658,N_1391,N_1268);
nand U1659 (N_1659,N_1186,N_1082);
or U1660 (N_1660,N_1347,N_1239);
or U1661 (N_1661,N_1272,N_1054);
or U1662 (N_1662,N_1150,N_1337);
xnor U1663 (N_1663,N_1209,N_1499);
and U1664 (N_1664,N_1451,N_1339);
nand U1665 (N_1665,N_1357,N_1182);
nor U1666 (N_1666,N_1126,N_1087);
nand U1667 (N_1667,N_1341,N_1259);
and U1668 (N_1668,N_1336,N_1234);
nand U1669 (N_1669,N_1207,N_1447);
nor U1670 (N_1670,N_1215,N_1155);
and U1671 (N_1671,N_1162,N_1278);
nor U1672 (N_1672,N_1227,N_1119);
xor U1673 (N_1673,N_1098,N_1125);
nand U1674 (N_1674,N_1277,N_1362);
and U1675 (N_1675,N_1246,N_1257);
and U1676 (N_1676,N_1223,N_1108);
or U1677 (N_1677,N_1165,N_1366);
xnor U1678 (N_1678,N_1025,N_1322);
and U1679 (N_1679,N_1307,N_1105);
or U1680 (N_1680,N_1099,N_1044);
nand U1681 (N_1681,N_1056,N_1001);
or U1682 (N_1682,N_1062,N_1334);
nor U1683 (N_1683,N_1113,N_1436);
xnor U1684 (N_1684,N_1200,N_1225);
nand U1685 (N_1685,N_1363,N_1235);
or U1686 (N_1686,N_1038,N_1201);
and U1687 (N_1687,N_1483,N_1035);
nand U1688 (N_1688,N_1342,N_1152);
xor U1689 (N_1689,N_1177,N_1433);
xnor U1690 (N_1690,N_1171,N_1233);
nor U1691 (N_1691,N_1255,N_1229);
nand U1692 (N_1692,N_1091,N_1489);
and U1693 (N_1693,N_1444,N_1000);
xor U1694 (N_1694,N_1412,N_1228);
or U1695 (N_1695,N_1118,N_1377);
or U1696 (N_1696,N_1397,N_1184);
nor U1697 (N_1697,N_1249,N_1440);
nand U1698 (N_1698,N_1331,N_1135);
or U1699 (N_1699,N_1051,N_1033);
nor U1700 (N_1700,N_1212,N_1424);
and U1701 (N_1701,N_1310,N_1285);
nor U1702 (N_1702,N_1260,N_1432);
and U1703 (N_1703,N_1060,N_1153);
and U1704 (N_1704,N_1023,N_1490);
and U1705 (N_1705,N_1149,N_1382);
or U1706 (N_1706,N_1318,N_1037);
or U1707 (N_1707,N_1163,N_1454);
nand U1708 (N_1708,N_1059,N_1048);
or U1709 (N_1709,N_1096,N_1328);
xnor U1710 (N_1710,N_1238,N_1473);
xor U1711 (N_1711,N_1151,N_1441);
nor U1712 (N_1712,N_1450,N_1131);
and U1713 (N_1713,N_1230,N_1428);
xor U1714 (N_1714,N_1088,N_1396);
nand U1715 (N_1715,N_1456,N_1461);
xor U1716 (N_1716,N_1371,N_1027);
xnor U1717 (N_1717,N_1297,N_1167);
xnor U1718 (N_1718,N_1192,N_1014);
or U1719 (N_1719,N_1369,N_1173);
and U1720 (N_1720,N_1176,N_1009);
nand U1721 (N_1721,N_1446,N_1359);
or U1722 (N_1722,N_1356,N_1061);
nor U1723 (N_1723,N_1290,N_1269);
xnor U1724 (N_1724,N_1367,N_1024);
nand U1725 (N_1725,N_1388,N_1093);
nand U1726 (N_1726,N_1248,N_1158);
nand U1727 (N_1727,N_1448,N_1316);
and U1728 (N_1728,N_1417,N_1471);
or U1729 (N_1729,N_1134,N_1138);
or U1730 (N_1730,N_1078,N_1460);
or U1731 (N_1731,N_1289,N_1462);
nand U1732 (N_1732,N_1308,N_1426);
nor U1733 (N_1733,N_1144,N_1498);
xor U1734 (N_1734,N_1111,N_1231);
nor U1735 (N_1735,N_1222,N_1133);
nor U1736 (N_1736,N_1067,N_1195);
nand U1737 (N_1737,N_1459,N_1103);
or U1738 (N_1738,N_1124,N_1481);
and U1739 (N_1739,N_1041,N_1028);
nand U1740 (N_1740,N_1107,N_1117);
and U1741 (N_1741,N_1365,N_1312);
nand U1742 (N_1742,N_1373,N_1279);
nor U1743 (N_1743,N_1261,N_1166);
xor U1744 (N_1744,N_1032,N_1016);
and U1745 (N_1745,N_1320,N_1017);
or U1746 (N_1746,N_1346,N_1140);
nor U1747 (N_1747,N_1335,N_1042);
xor U1748 (N_1748,N_1128,N_1485);
nor U1749 (N_1749,N_1443,N_1069);
or U1750 (N_1750,N_1277,N_1297);
or U1751 (N_1751,N_1272,N_1298);
nor U1752 (N_1752,N_1401,N_1093);
nor U1753 (N_1753,N_1010,N_1490);
and U1754 (N_1754,N_1153,N_1355);
and U1755 (N_1755,N_1161,N_1486);
or U1756 (N_1756,N_1015,N_1310);
nand U1757 (N_1757,N_1458,N_1323);
or U1758 (N_1758,N_1385,N_1479);
nand U1759 (N_1759,N_1314,N_1372);
nand U1760 (N_1760,N_1311,N_1216);
or U1761 (N_1761,N_1307,N_1179);
xnor U1762 (N_1762,N_1050,N_1173);
xor U1763 (N_1763,N_1233,N_1026);
and U1764 (N_1764,N_1135,N_1041);
nand U1765 (N_1765,N_1060,N_1321);
nor U1766 (N_1766,N_1217,N_1334);
and U1767 (N_1767,N_1408,N_1108);
nand U1768 (N_1768,N_1203,N_1436);
xor U1769 (N_1769,N_1169,N_1292);
or U1770 (N_1770,N_1457,N_1248);
or U1771 (N_1771,N_1443,N_1140);
nor U1772 (N_1772,N_1361,N_1010);
or U1773 (N_1773,N_1429,N_1248);
nand U1774 (N_1774,N_1015,N_1020);
nand U1775 (N_1775,N_1012,N_1370);
or U1776 (N_1776,N_1141,N_1101);
and U1777 (N_1777,N_1211,N_1418);
and U1778 (N_1778,N_1040,N_1180);
xnor U1779 (N_1779,N_1413,N_1479);
or U1780 (N_1780,N_1033,N_1134);
xor U1781 (N_1781,N_1243,N_1341);
xnor U1782 (N_1782,N_1223,N_1267);
nor U1783 (N_1783,N_1474,N_1091);
and U1784 (N_1784,N_1296,N_1033);
or U1785 (N_1785,N_1248,N_1237);
and U1786 (N_1786,N_1126,N_1270);
xnor U1787 (N_1787,N_1443,N_1257);
nor U1788 (N_1788,N_1495,N_1299);
and U1789 (N_1789,N_1015,N_1410);
and U1790 (N_1790,N_1098,N_1407);
or U1791 (N_1791,N_1390,N_1336);
nand U1792 (N_1792,N_1260,N_1118);
nand U1793 (N_1793,N_1455,N_1267);
nor U1794 (N_1794,N_1001,N_1248);
or U1795 (N_1795,N_1026,N_1103);
xor U1796 (N_1796,N_1356,N_1206);
xor U1797 (N_1797,N_1411,N_1289);
nand U1798 (N_1798,N_1187,N_1263);
or U1799 (N_1799,N_1216,N_1371);
xnor U1800 (N_1800,N_1473,N_1329);
nor U1801 (N_1801,N_1125,N_1414);
nor U1802 (N_1802,N_1453,N_1365);
or U1803 (N_1803,N_1076,N_1073);
xor U1804 (N_1804,N_1102,N_1157);
nand U1805 (N_1805,N_1112,N_1090);
and U1806 (N_1806,N_1021,N_1137);
nor U1807 (N_1807,N_1229,N_1160);
or U1808 (N_1808,N_1063,N_1272);
nand U1809 (N_1809,N_1317,N_1107);
and U1810 (N_1810,N_1478,N_1276);
xnor U1811 (N_1811,N_1091,N_1193);
or U1812 (N_1812,N_1032,N_1024);
xnor U1813 (N_1813,N_1151,N_1236);
or U1814 (N_1814,N_1258,N_1495);
or U1815 (N_1815,N_1257,N_1333);
nor U1816 (N_1816,N_1110,N_1468);
nor U1817 (N_1817,N_1058,N_1408);
xnor U1818 (N_1818,N_1370,N_1396);
xor U1819 (N_1819,N_1335,N_1048);
or U1820 (N_1820,N_1281,N_1105);
xor U1821 (N_1821,N_1258,N_1358);
nand U1822 (N_1822,N_1446,N_1235);
and U1823 (N_1823,N_1494,N_1245);
xnor U1824 (N_1824,N_1286,N_1483);
and U1825 (N_1825,N_1196,N_1377);
and U1826 (N_1826,N_1470,N_1134);
and U1827 (N_1827,N_1158,N_1476);
or U1828 (N_1828,N_1495,N_1126);
or U1829 (N_1829,N_1257,N_1345);
or U1830 (N_1830,N_1079,N_1335);
nor U1831 (N_1831,N_1029,N_1406);
or U1832 (N_1832,N_1307,N_1084);
and U1833 (N_1833,N_1031,N_1360);
and U1834 (N_1834,N_1128,N_1071);
nand U1835 (N_1835,N_1050,N_1193);
or U1836 (N_1836,N_1019,N_1274);
and U1837 (N_1837,N_1230,N_1470);
xor U1838 (N_1838,N_1227,N_1012);
nor U1839 (N_1839,N_1347,N_1266);
or U1840 (N_1840,N_1385,N_1382);
nor U1841 (N_1841,N_1068,N_1420);
nor U1842 (N_1842,N_1092,N_1471);
and U1843 (N_1843,N_1460,N_1175);
or U1844 (N_1844,N_1255,N_1410);
and U1845 (N_1845,N_1007,N_1207);
nand U1846 (N_1846,N_1267,N_1082);
or U1847 (N_1847,N_1094,N_1229);
or U1848 (N_1848,N_1416,N_1030);
and U1849 (N_1849,N_1021,N_1092);
nor U1850 (N_1850,N_1396,N_1393);
xor U1851 (N_1851,N_1009,N_1251);
nand U1852 (N_1852,N_1106,N_1225);
xor U1853 (N_1853,N_1305,N_1337);
or U1854 (N_1854,N_1040,N_1158);
nand U1855 (N_1855,N_1310,N_1099);
xor U1856 (N_1856,N_1141,N_1483);
or U1857 (N_1857,N_1217,N_1390);
or U1858 (N_1858,N_1366,N_1326);
or U1859 (N_1859,N_1277,N_1084);
nor U1860 (N_1860,N_1232,N_1166);
nand U1861 (N_1861,N_1435,N_1004);
or U1862 (N_1862,N_1235,N_1115);
nand U1863 (N_1863,N_1454,N_1438);
xnor U1864 (N_1864,N_1127,N_1273);
or U1865 (N_1865,N_1082,N_1278);
nand U1866 (N_1866,N_1228,N_1342);
or U1867 (N_1867,N_1019,N_1188);
nand U1868 (N_1868,N_1175,N_1453);
xnor U1869 (N_1869,N_1245,N_1120);
and U1870 (N_1870,N_1198,N_1020);
and U1871 (N_1871,N_1366,N_1426);
nand U1872 (N_1872,N_1377,N_1481);
and U1873 (N_1873,N_1049,N_1338);
and U1874 (N_1874,N_1480,N_1246);
or U1875 (N_1875,N_1444,N_1331);
nor U1876 (N_1876,N_1448,N_1420);
or U1877 (N_1877,N_1300,N_1356);
or U1878 (N_1878,N_1337,N_1005);
and U1879 (N_1879,N_1434,N_1237);
xnor U1880 (N_1880,N_1008,N_1313);
nand U1881 (N_1881,N_1265,N_1430);
nand U1882 (N_1882,N_1274,N_1185);
nand U1883 (N_1883,N_1302,N_1113);
and U1884 (N_1884,N_1167,N_1396);
nor U1885 (N_1885,N_1129,N_1083);
nand U1886 (N_1886,N_1128,N_1273);
and U1887 (N_1887,N_1384,N_1359);
and U1888 (N_1888,N_1150,N_1236);
and U1889 (N_1889,N_1299,N_1134);
nor U1890 (N_1890,N_1189,N_1156);
or U1891 (N_1891,N_1074,N_1259);
or U1892 (N_1892,N_1214,N_1474);
nor U1893 (N_1893,N_1370,N_1175);
nor U1894 (N_1894,N_1431,N_1200);
or U1895 (N_1895,N_1158,N_1308);
and U1896 (N_1896,N_1471,N_1359);
or U1897 (N_1897,N_1348,N_1077);
or U1898 (N_1898,N_1104,N_1478);
nor U1899 (N_1899,N_1066,N_1005);
nand U1900 (N_1900,N_1006,N_1026);
and U1901 (N_1901,N_1484,N_1222);
nand U1902 (N_1902,N_1110,N_1181);
or U1903 (N_1903,N_1292,N_1175);
and U1904 (N_1904,N_1118,N_1069);
nand U1905 (N_1905,N_1129,N_1176);
nor U1906 (N_1906,N_1418,N_1195);
or U1907 (N_1907,N_1288,N_1474);
nand U1908 (N_1908,N_1200,N_1451);
and U1909 (N_1909,N_1273,N_1120);
nand U1910 (N_1910,N_1338,N_1284);
and U1911 (N_1911,N_1292,N_1465);
or U1912 (N_1912,N_1102,N_1116);
nor U1913 (N_1913,N_1289,N_1387);
nand U1914 (N_1914,N_1331,N_1039);
nand U1915 (N_1915,N_1050,N_1062);
nand U1916 (N_1916,N_1244,N_1414);
xnor U1917 (N_1917,N_1252,N_1175);
nor U1918 (N_1918,N_1022,N_1252);
nand U1919 (N_1919,N_1282,N_1217);
xnor U1920 (N_1920,N_1138,N_1191);
nand U1921 (N_1921,N_1419,N_1364);
nor U1922 (N_1922,N_1023,N_1440);
nor U1923 (N_1923,N_1208,N_1301);
and U1924 (N_1924,N_1264,N_1106);
xor U1925 (N_1925,N_1499,N_1472);
and U1926 (N_1926,N_1199,N_1079);
nor U1927 (N_1927,N_1330,N_1348);
xnor U1928 (N_1928,N_1427,N_1328);
nor U1929 (N_1929,N_1389,N_1069);
nor U1930 (N_1930,N_1447,N_1406);
nor U1931 (N_1931,N_1110,N_1130);
nand U1932 (N_1932,N_1397,N_1432);
nor U1933 (N_1933,N_1133,N_1431);
or U1934 (N_1934,N_1353,N_1146);
and U1935 (N_1935,N_1476,N_1404);
or U1936 (N_1936,N_1153,N_1484);
or U1937 (N_1937,N_1311,N_1053);
or U1938 (N_1938,N_1481,N_1345);
and U1939 (N_1939,N_1225,N_1346);
nor U1940 (N_1940,N_1216,N_1491);
nand U1941 (N_1941,N_1176,N_1462);
nor U1942 (N_1942,N_1137,N_1058);
or U1943 (N_1943,N_1360,N_1444);
or U1944 (N_1944,N_1487,N_1205);
nand U1945 (N_1945,N_1433,N_1277);
nor U1946 (N_1946,N_1479,N_1407);
xnor U1947 (N_1947,N_1186,N_1045);
and U1948 (N_1948,N_1186,N_1236);
nand U1949 (N_1949,N_1004,N_1097);
xnor U1950 (N_1950,N_1235,N_1069);
and U1951 (N_1951,N_1490,N_1210);
nand U1952 (N_1952,N_1482,N_1002);
nand U1953 (N_1953,N_1429,N_1162);
xnor U1954 (N_1954,N_1493,N_1079);
and U1955 (N_1955,N_1451,N_1064);
nand U1956 (N_1956,N_1132,N_1352);
or U1957 (N_1957,N_1102,N_1091);
or U1958 (N_1958,N_1068,N_1176);
nand U1959 (N_1959,N_1027,N_1325);
or U1960 (N_1960,N_1099,N_1320);
or U1961 (N_1961,N_1385,N_1402);
xor U1962 (N_1962,N_1461,N_1155);
and U1963 (N_1963,N_1374,N_1307);
nand U1964 (N_1964,N_1094,N_1054);
xnor U1965 (N_1965,N_1211,N_1468);
and U1966 (N_1966,N_1078,N_1114);
or U1967 (N_1967,N_1090,N_1380);
nand U1968 (N_1968,N_1380,N_1207);
nand U1969 (N_1969,N_1102,N_1380);
or U1970 (N_1970,N_1114,N_1382);
or U1971 (N_1971,N_1008,N_1306);
nand U1972 (N_1972,N_1078,N_1159);
nand U1973 (N_1973,N_1006,N_1496);
nand U1974 (N_1974,N_1330,N_1239);
nand U1975 (N_1975,N_1181,N_1303);
nor U1976 (N_1976,N_1319,N_1123);
or U1977 (N_1977,N_1239,N_1232);
xor U1978 (N_1978,N_1317,N_1256);
or U1979 (N_1979,N_1018,N_1156);
xnor U1980 (N_1980,N_1476,N_1114);
nor U1981 (N_1981,N_1056,N_1242);
nor U1982 (N_1982,N_1467,N_1410);
nor U1983 (N_1983,N_1115,N_1029);
nand U1984 (N_1984,N_1040,N_1287);
or U1985 (N_1985,N_1029,N_1118);
xor U1986 (N_1986,N_1415,N_1138);
nand U1987 (N_1987,N_1286,N_1099);
xor U1988 (N_1988,N_1392,N_1370);
xor U1989 (N_1989,N_1414,N_1195);
nor U1990 (N_1990,N_1155,N_1402);
and U1991 (N_1991,N_1439,N_1476);
nor U1992 (N_1992,N_1171,N_1324);
or U1993 (N_1993,N_1258,N_1031);
nand U1994 (N_1994,N_1409,N_1214);
nand U1995 (N_1995,N_1040,N_1465);
nor U1996 (N_1996,N_1115,N_1051);
nor U1997 (N_1997,N_1343,N_1038);
or U1998 (N_1998,N_1154,N_1098);
nor U1999 (N_1999,N_1488,N_1420);
nor U2000 (N_2000,N_1528,N_1733);
or U2001 (N_2001,N_1636,N_1756);
nand U2002 (N_2002,N_1899,N_1639);
or U2003 (N_2003,N_1894,N_1778);
or U2004 (N_2004,N_1923,N_1822);
nand U2005 (N_2005,N_1637,N_1737);
or U2006 (N_2006,N_1764,N_1663);
xnor U2007 (N_2007,N_1978,N_1754);
or U2008 (N_2008,N_1815,N_1510);
nand U2009 (N_2009,N_1695,N_1929);
nand U2010 (N_2010,N_1890,N_1846);
and U2011 (N_2011,N_1717,N_1839);
or U2012 (N_2012,N_1776,N_1877);
or U2013 (N_2013,N_1755,N_1950);
and U2014 (N_2014,N_1848,N_1644);
xor U2015 (N_2015,N_1675,N_1579);
or U2016 (N_2016,N_1531,N_1607);
xnor U2017 (N_2017,N_1593,N_1605);
nand U2018 (N_2018,N_1986,N_1585);
nor U2019 (N_2019,N_1862,N_1603);
or U2020 (N_2020,N_1614,N_1803);
xnor U2021 (N_2021,N_1845,N_1727);
nand U2022 (N_2022,N_1601,N_1565);
or U2023 (N_2023,N_1933,N_1627);
xor U2024 (N_2024,N_1806,N_1811);
nor U2025 (N_2025,N_1854,N_1504);
xnor U2026 (N_2026,N_1514,N_1560);
or U2027 (N_2027,N_1793,N_1685);
and U2028 (N_2028,N_1796,N_1789);
and U2029 (N_2029,N_1936,N_1613);
or U2030 (N_2030,N_1974,N_1958);
nand U2031 (N_2031,N_1692,N_1887);
xor U2032 (N_2032,N_1716,N_1645);
or U2033 (N_2033,N_1745,N_1784);
or U2034 (N_2034,N_1729,N_1930);
xnor U2035 (N_2035,N_1909,N_1970);
nor U2036 (N_2036,N_1892,N_1828);
nand U2037 (N_2037,N_1766,N_1819);
xnor U2038 (N_2038,N_1797,N_1689);
and U2039 (N_2039,N_1505,N_1698);
xor U2040 (N_2040,N_1691,N_1515);
nand U2041 (N_2041,N_1699,N_1836);
and U2042 (N_2042,N_1540,N_1643);
nand U2043 (N_2043,N_1667,N_1773);
or U2044 (N_2044,N_1992,N_1997);
or U2045 (N_2045,N_1654,N_1906);
xnor U2046 (N_2046,N_1511,N_1999);
xnor U2047 (N_2047,N_1652,N_1704);
and U2048 (N_2048,N_1810,N_1650);
xor U2049 (N_2049,N_1620,N_1577);
nor U2050 (N_2050,N_1640,N_1509);
xor U2051 (N_2051,N_1934,N_1517);
nor U2052 (N_2052,N_1533,N_1713);
or U2053 (N_2053,N_1963,N_1611);
and U2054 (N_2054,N_1855,N_1673);
nor U2055 (N_2055,N_1911,N_1995);
nor U2056 (N_2056,N_1834,N_1990);
or U2057 (N_2057,N_1825,N_1738);
nand U2058 (N_2058,N_1569,N_1946);
nand U2059 (N_2059,N_1922,N_1628);
xor U2060 (N_2060,N_1649,N_1941);
nor U2061 (N_2061,N_1897,N_1655);
or U2062 (N_2062,N_1696,N_1521);
nor U2063 (N_2063,N_1966,N_1881);
nor U2064 (N_2064,N_1910,N_1570);
nor U2065 (N_2065,N_1982,N_1872);
nand U2066 (N_2066,N_1953,N_1981);
nand U2067 (N_2067,N_1747,N_1952);
and U2068 (N_2068,N_1954,N_1718);
xnor U2069 (N_2069,N_1840,N_1775);
xnor U2070 (N_2070,N_1571,N_1534);
or U2071 (N_2071,N_1888,N_1710);
nand U2072 (N_2072,N_1817,N_1705);
or U2073 (N_2073,N_1557,N_1731);
or U2074 (N_2074,N_1693,N_1683);
or U2075 (N_2075,N_1641,N_1939);
and U2076 (N_2076,N_1559,N_1860);
nand U2077 (N_2077,N_1634,N_1724);
and U2078 (N_2078,N_1891,N_1626);
nor U2079 (N_2079,N_1588,N_1556);
nand U2080 (N_2080,N_1612,N_1753);
nand U2081 (N_2081,N_1550,N_1546);
and U2082 (N_2082,N_1824,N_1771);
or U2083 (N_2083,N_1945,N_1538);
nor U2084 (N_2084,N_1527,N_1545);
nand U2085 (N_2085,N_1554,N_1656);
nor U2086 (N_2086,N_1568,N_1779);
xor U2087 (N_2087,N_1838,N_1786);
or U2088 (N_2088,N_1595,N_1969);
nand U2089 (N_2089,N_1617,N_1622);
nand U2090 (N_2090,N_1761,N_1799);
nor U2091 (N_2091,N_1908,N_1980);
or U2092 (N_2092,N_1916,N_1851);
and U2093 (N_2093,N_1878,N_1508);
nand U2094 (N_2094,N_1935,N_1742);
nor U2095 (N_2095,N_1991,N_1985);
nor U2096 (N_2096,N_1587,N_1657);
nand U2097 (N_2097,N_1940,N_1760);
nand U2098 (N_2098,N_1706,N_1833);
nor U2099 (N_2099,N_1998,N_1555);
xnor U2100 (N_2100,N_1676,N_1751);
and U2101 (N_2101,N_1948,N_1541);
and U2102 (N_2102,N_1807,N_1506);
and U2103 (N_2103,N_1821,N_1873);
xor U2104 (N_2104,N_1700,N_1616);
and U2105 (N_2105,N_1904,N_1519);
and U2106 (N_2106,N_1726,N_1516);
or U2107 (N_2107,N_1635,N_1594);
and U2108 (N_2108,N_1841,N_1621);
and U2109 (N_2109,N_1648,N_1863);
or U2110 (N_2110,N_1866,N_1827);
nand U2111 (N_2111,N_1791,N_1837);
nand U2112 (N_2112,N_1679,N_1677);
xor U2113 (N_2113,N_1502,N_1987);
or U2114 (N_2114,N_1578,N_1767);
nor U2115 (N_2115,N_1665,N_1943);
and U2116 (N_2116,N_1591,N_1900);
nand U2117 (N_2117,N_1927,N_1674);
and U2118 (N_2118,N_1883,N_1542);
or U2119 (N_2119,N_1740,N_1915);
nor U2120 (N_2120,N_1592,N_1814);
nor U2121 (N_2121,N_1563,N_1709);
or U2122 (N_2122,N_1507,N_1772);
xor U2123 (N_2123,N_1720,N_1602);
xnor U2124 (N_2124,N_1867,N_1905);
or U2125 (N_2125,N_1886,N_1765);
and U2126 (N_2126,N_1971,N_1875);
and U2127 (N_2127,N_1794,N_1730);
nor U2128 (N_2128,N_1926,N_1746);
xor U2129 (N_2129,N_1896,N_1660);
and U2130 (N_2130,N_1711,N_1543);
xnor U2131 (N_2131,N_1748,N_1993);
or U2132 (N_2132,N_1647,N_1670);
nand U2133 (N_2133,N_1889,N_1879);
and U2134 (N_2134,N_1532,N_1813);
and U2135 (N_2135,N_1526,N_1816);
or U2136 (N_2136,N_1523,N_1962);
nand U2137 (N_2137,N_1633,N_1801);
or U2138 (N_2138,N_1610,N_1805);
nand U2139 (N_2139,N_1979,N_1763);
and U2140 (N_2140,N_1947,N_1653);
xnor U2141 (N_2141,N_1880,N_1820);
nor U2142 (N_2142,N_1608,N_1988);
xor U2143 (N_2143,N_1576,N_1931);
nand U2144 (N_2144,N_1960,N_1818);
nor U2145 (N_2145,N_1580,N_1809);
nor U2146 (N_2146,N_1938,N_1917);
nor U2147 (N_2147,N_1712,N_1549);
xnor U2148 (N_2148,N_1924,N_1902);
or U2149 (N_2149,N_1949,N_1512);
nand U2150 (N_2150,N_1996,N_1732);
nor U2151 (N_2151,N_1690,N_1800);
and U2152 (N_2152,N_1882,N_1672);
xor U2153 (N_2153,N_1823,N_1812);
xnor U2154 (N_2154,N_1625,N_1537);
and U2155 (N_2155,N_1604,N_1918);
xnor U2156 (N_2156,N_1629,N_1965);
nor U2157 (N_2157,N_1937,N_1664);
and U2158 (N_2158,N_1544,N_1669);
or U2159 (N_2159,N_1661,N_1869);
nand U2160 (N_2160,N_1864,N_1868);
or U2161 (N_2161,N_1852,N_1619);
nor U2162 (N_2162,N_1826,N_1686);
and U2163 (N_2163,N_1850,N_1770);
xnor U2164 (N_2164,N_1758,N_1702);
xor U2165 (N_2165,N_1522,N_1623);
or U2166 (N_2166,N_1944,N_1870);
xor U2167 (N_2167,N_1553,N_1694);
nand U2168 (N_2168,N_1638,N_1972);
or U2169 (N_2169,N_1893,N_1903);
and U2170 (N_2170,N_1624,N_1808);
and U2171 (N_2171,N_1600,N_1662);
and U2172 (N_2172,N_1795,N_1697);
xor U2173 (N_2173,N_1501,N_1725);
or U2174 (N_2174,N_1874,N_1843);
and U2175 (N_2175,N_1581,N_1895);
nor U2176 (N_2176,N_1583,N_1562);
nand U2177 (N_2177,N_1928,N_1994);
or U2178 (N_2178,N_1914,N_1885);
nor U2179 (N_2179,N_1925,N_1658);
or U2180 (N_2180,N_1983,N_1682);
xnor U2181 (N_2181,N_1856,N_1567);
or U2182 (N_2182,N_1500,N_1844);
and U2183 (N_2183,N_1574,N_1535);
and U2184 (N_2184,N_1707,N_1921);
and U2185 (N_2185,N_1884,N_1596);
xnor U2186 (N_2186,N_1520,N_1989);
nand U2187 (N_2187,N_1932,N_1642);
nand U2188 (N_2188,N_1714,N_1715);
xnor U2189 (N_2189,N_1744,N_1781);
xor U2190 (N_2190,N_1842,N_1802);
nor U2191 (N_2191,N_1831,N_1736);
and U2192 (N_2192,N_1548,N_1762);
nor U2193 (N_2193,N_1804,N_1798);
or U2194 (N_2194,N_1721,N_1768);
nand U2195 (N_2195,N_1680,N_1835);
xor U2196 (N_2196,N_1750,N_1968);
xnor U2197 (N_2197,N_1792,N_1566);
nor U2198 (N_2198,N_1630,N_1572);
nand U2199 (N_2199,N_1849,N_1539);
or U2200 (N_2200,N_1774,N_1956);
nor U2201 (N_2201,N_1898,N_1876);
xnor U2202 (N_2202,N_1728,N_1919);
or U2203 (N_2203,N_1973,N_1769);
or U2204 (N_2204,N_1759,N_1787);
xor U2205 (N_2205,N_1651,N_1959);
nand U2206 (N_2206,N_1708,N_1551);
and U2207 (N_2207,N_1598,N_1552);
or U2208 (N_2208,N_1782,N_1536);
nor U2209 (N_2209,N_1861,N_1865);
nor U2210 (N_2210,N_1920,N_1967);
nand U2211 (N_2211,N_1688,N_1857);
xnor U2212 (N_2212,N_1951,N_1942);
nor U2213 (N_2213,N_1599,N_1561);
nor U2214 (N_2214,N_1703,N_1907);
xnor U2215 (N_2215,N_1547,N_1777);
or U2216 (N_2216,N_1859,N_1735);
nor U2217 (N_2217,N_1739,N_1913);
xnor U2218 (N_2218,N_1977,N_1575);
nor U2219 (N_2219,N_1976,N_1785);
xnor U2220 (N_2220,N_1830,N_1632);
and U2221 (N_2221,N_1668,N_1590);
xor U2222 (N_2222,N_1788,N_1757);
or U2223 (N_2223,N_1722,N_1701);
xnor U2224 (N_2224,N_1558,N_1573);
nand U2225 (N_2225,N_1961,N_1752);
or U2226 (N_2226,N_1871,N_1687);
or U2227 (N_2227,N_1586,N_1678);
and U2228 (N_2228,N_1790,N_1564);
nand U2229 (N_2229,N_1666,N_1524);
and U2230 (N_2230,N_1530,N_1529);
xor U2231 (N_2231,N_1584,N_1681);
nand U2232 (N_2232,N_1597,N_1525);
nand U2233 (N_2233,N_1741,N_1615);
or U2234 (N_2234,N_1780,N_1858);
xor U2235 (N_2235,N_1912,N_1853);
or U2236 (N_2236,N_1955,N_1901);
nand U2237 (N_2237,N_1829,N_1719);
and U2238 (N_2238,N_1618,N_1723);
nor U2239 (N_2239,N_1659,N_1503);
xor U2240 (N_2240,N_1518,N_1749);
or U2241 (N_2241,N_1513,N_1646);
xor U2242 (N_2242,N_1783,N_1957);
xor U2243 (N_2243,N_1631,N_1606);
and U2244 (N_2244,N_1684,N_1671);
nand U2245 (N_2245,N_1975,N_1734);
nor U2246 (N_2246,N_1609,N_1832);
nor U2247 (N_2247,N_1743,N_1847);
and U2248 (N_2248,N_1589,N_1964);
and U2249 (N_2249,N_1984,N_1582);
nand U2250 (N_2250,N_1940,N_1886);
and U2251 (N_2251,N_1715,N_1760);
nor U2252 (N_2252,N_1902,N_1763);
or U2253 (N_2253,N_1778,N_1871);
xnor U2254 (N_2254,N_1775,N_1830);
nor U2255 (N_2255,N_1960,N_1763);
xnor U2256 (N_2256,N_1651,N_1523);
nand U2257 (N_2257,N_1596,N_1732);
xnor U2258 (N_2258,N_1672,N_1999);
xor U2259 (N_2259,N_1987,N_1917);
and U2260 (N_2260,N_1613,N_1788);
nand U2261 (N_2261,N_1832,N_1589);
or U2262 (N_2262,N_1842,N_1677);
nor U2263 (N_2263,N_1944,N_1838);
nor U2264 (N_2264,N_1691,N_1891);
xnor U2265 (N_2265,N_1907,N_1870);
and U2266 (N_2266,N_1715,N_1792);
or U2267 (N_2267,N_1937,N_1870);
nor U2268 (N_2268,N_1623,N_1526);
nand U2269 (N_2269,N_1706,N_1889);
xnor U2270 (N_2270,N_1668,N_1766);
nand U2271 (N_2271,N_1569,N_1761);
nand U2272 (N_2272,N_1812,N_1642);
nor U2273 (N_2273,N_1523,N_1950);
nand U2274 (N_2274,N_1966,N_1935);
nor U2275 (N_2275,N_1853,N_1840);
xnor U2276 (N_2276,N_1572,N_1688);
and U2277 (N_2277,N_1672,N_1638);
and U2278 (N_2278,N_1807,N_1711);
and U2279 (N_2279,N_1982,N_1765);
xor U2280 (N_2280,N_1522,N_1838);
and U2281 (N_2281,N_1682,N_1754);
or U2282 (N_2282,N_1707,N_1893);
xnor U2283 (N_2283,N_1824,N_1898);
nand U2284 (N_2284,N_1755,N_1612);
nand U2285 (N_2285,N_1637,N_1544);
nor U2286 (N_2286,N_1694,N_1621);
and U2287 (N_2287,N_1741,N_1793);
nand U2288 (N_2288,N_1530,N_1808);
nand U2289 (N_2289,N_1901,N_1961);
nand U2290 (N_2290,N_1964,N_1863);
xnor U2291 (N_2291,N_1687,N_1873);
nor U2292 (N_2292,N_1514,N_1528);
xor U2293 (N_2293,N_1827,N_1906);
or U2294 (N_2294,N_1737,N_1719);
and U2295 (N_2295,N_1786,N_1861);
xor U2296 (N_2296,N_1766,N_1999);
or U2297 (N_2297,N_1716,N_1531);
nand U2298 (N_2298,N_1673,N_1704);
xnor U2299 (N_2299,N_1693,N_1577);
nand U2300 (N_2300,N_1538,N_1794);
or U2301 (N_2301,N_1608,N_1613);
nor U2302 (N_2302,N_1579,N_1711);
nor U2303 (N_2303,N_1741,N_1764);
nor U2304 (N_2304,N_1841,N_1707);
or U2305 (N_2305,N_1521,N_1918);
and U2306 (N_2306,N_1738,N_1505);
and U2307 (N_2307,N_1633,N_1814);
or U2308 (N_2308,N_1924,N_1910);
and U2309 (N_2309,N_1979,N_1778);
nand U2310 (N_2310,N_1944,N_1575);
or U2311 (N_2311,N_1728,N_1940);
nand U2312 (N_2312,N_1575,N_1775);
nand U2313 (N_2313,N_1720,N_1862);
and U2314 (N_2314,N_1801,N_1789);
nor U2315 (N_2315,N_1545,N_1974);
nand U2316 (N_2316,N_1993,N_1902);
or U2317 (N_2317,N_1730,N_1868);
xnor U2318 (N_2318,N_1889,N_1563);
or U2319 (N_2319,N_1689,N_1887);
nand U2320 (N_2320,N_1733,N_1862);
nor U2321 (N_2321,N_1794,N_1622);
nand U2322 (N_2322,N_1841,N_1719);
xor U2323 (N_2323,N_1504,N_1685);
xnor U2324 (N_2324,N_1832,N_1508);
nand U2325 (N_2325,N_1656,N_1564);
or U2326 (N_2326,N_1509,N_1902);
nor U2327 (N_2327,N_1835,N_1553);
xor U2328 (N_2328,N_1954,N_1608);
xnor U2329 (N_2329,N_1529,N_1822);
nor U2330 (N_2330,N_1890,N_1529);
nand U2331 (N_2331,N_1607,N_1759);
nand U2332 (N_2332,N_1990,N_1672);
nor U2333 (N_2333,N_1630,N_1932);
nand U2334 (N_2334,N_1801,N_1781);
and U2335 (N_2335,N_1544,N_1722);
or U2336 (N_2336,N_1666,N_1808);
and U2337 (N_2337,N_1962,N_1578);
or U2338 (N_2338,N_1945,N_1990);
xnor U2339 (N_2339,N_1797,N_1820);
and U2340 (N_2340,N_1980,N_1830);
xor U2341 (N_2341,N_1767,N_1641);
nor U2342 (N_2342,N_1947,N_1546);
nand U2343 (N_2343,N_1591,N_1882);
nor U2344 (N_2344,N_1776,N_1505);
xnor U2345 (N_2345,N_1783,N_1916);
xor U2346 (N_2346,N_1966,N_1704);
xor U2347 (N_2347,N_1674,N_1588);
nand U2348 (N_2348,N_1550,N_1602);
nor U2349 (N_2349,N_1776,N_1821);
xnor U2350 (N_2350,N_1816,N_1703);
or U2351 (N_2351,N_1555,N_1972);
or U2352 (N_2352,N_1647,N_1611);
nand U2353 (N_2353,N_1646,N_1888);
xor U2354 (N_2354,N_1811,N_1772);
or U2355 (N_2355,N_1581,N_1639);
nor U2356 (N_2356,N_1858,N_1530);
and U2357 (N_2357,N_1717,N_1974);
nand U2358 (N_2358,N_1533,N_1786);
nand U2359 (N_2359,N_1625,N_1735);
or U2360 (N_2360,N_1709,N_1791);
xor U2361 (N_2361,N_1667,N_1940);
nand U2362 (N_2362,N_1792,N_1764);
nand U2363 (N_2363,N_1551,N_1711);
or U2364 (N_2364,N_1791,N_1773);
nor U2365 (N_2365,N_1843,N_1993);
nor U2366 (N_2366,N_1869,N_1901);
nand U2367 (N_2367,N_1974,N_1836);
xor U2368 (N_2368,N_1920,N_1501);
and U2369 (N_2369,N_1887,N_1617);
nor U2370 (N_2370,N_1991,N_1640);
xnor U2371 (N_2371,N_1586,N_1852);
nand U2372 (N_2372,N_1896,N_1893);
nand U2373 (N_2373,N_1945,N_1819);
nand U2374 (N_2374,N_1718,N_1959);
xnor U2375 (N_2375,N_1943,N_1538);
nand U2376 (N_2376,N_1920,N_1900);
nand U2377 (N_2377,N_1680,N_1714);
nor U2378 (N_2378,N_1821,N_1630);
nand U2379 (N_2379,N_1564,N_1829);
and U2380 (N_2380,N_1605,N_1732);
nand U2381 (N_2381,N_1796,N_1851);
nand U2382 (N_2382,N_1528,N_1817);
xnor U2383 (N_2383,N_1770,N_1745);
xnor U2384 (N_2384,N_1666,N_1972);
and U2385 (N_2385,N_1703,N_1807);
nand U2386 (N_2386,N_1609,N_1847);
nor U2387 (N_2387,N_1975,N_1917);
or U2388 (N_2388,N_1912,N_1589);
nand U2389 (N_2389,N_1621,N_1810);
xnor U2390 (N_2390,N_1569,N_1895);
nor U2391 (N_2391,N_1958,N_1747);
or U2392 (N_2392,N_1579,N_1859);
and U2393 (N_2393,N_1590,N_1665);
nand U2394 (N_2394,N_1701,N_1576);
nor U2395 (N_2395,N_1834,N_1974);
nand U2396 (N_2396,N_1713,N_1852);
and U2397 (N_2397,N_1995,N_1699);
or U2398 (N_2398,N_1880,N_1956);
or U2399 (N_2399,N_1855,N_1716);
and U2400 (N_2400,N_1671,N_1508);
nand U2401 (N_2401,N_1547,N_1515);
or U2402 (N_2402,N_1876,N_1703);
or U2403 (N_2403,N_1924,N_1747);
nand U2404 (N_2404,N_1572,N_1574);
or U2405 (N_2405,N_1523,N_1964);
or U2406 (N_2406,N_1631,N_1685);
or U2407 (N_2407,N_1972,N_1777);
or U2408 (N_2408,N_1627,N_1918);
xor U2409 (N_2409,N_1801,N_1953);
nor U2410 (N_2410,N_1687,N_1945);
xnor U2411 (N_2411,N_1918,N_1911);
xor U2412 (N_2412,N_1977,N_1991);
xnor U2413 (N_2413,N_1628,N_1800);
and U2414 (N_2414,N_1894,N_1861);
and U2415 (N_2415,N_1715,N_1654);
and U2416 (N_2416,N_1502,N_1870);
nor U2417 (N_2417,N_1807,N_1989);
xor U2418 (N_2418,N_1503,N_1648);
or U2419 (N_2419,N_1746,N_1773);
xnor U2420 (N_2420,N_1907,N_1669);
nand U2421 (N_2421,N_1533,N_1993);
or U2422 (N_2422,N_1698,N_1631);
nor U2423 (N_2423,N_1888,N_1739);
nor U2424 (N_2424,N_1948,N_1572);
and U2425 (N_2425,N_1760,N_1888);
xnor U2426 (N_2426,N_1905,N_1943);
or U2427 (N_2427,N_1970,N_1943);
and U2428 (N_2428,N_1834,N_1545);
nor U2429 (N_2429,N_1774,N_1699);
or U2430 (N_2430,N_1550,N_1957);
xnor U2431 (N_2431,N_1822,N_1953);
nor U2432 (N_2432,N_1902,N_1703);
or U2433 (N_2433,N_1564,N_1928);
or U2434 (N_2434,N_1535,N_1548);
and U2435 (N_2435,N_1544,N_1801);
or U2436 (N_2436,N_1698,N_1515);
or U2437 (N_2437,N_1809,N_1955);
and U2438 (N_2438,N_1604,N_1804);
and U2439 (N_2439,N_1550,N_1655);
nor U2440 (N_2440,N_1766,N_1784);
or U2441 (N_2441,N_1703,N_1794);
nor U2442 (N_2442,N_1887,N_1851);
and U2443 (N_2443,N_1957,N_1794);
or U2444 (N_2444,N_1976,N_1613);
or U2445 (N_2445,N_1689,N_1928);
or U2446 (N_2446,N_1811,N_1906);
xnor U2447 (N_2447,N_1582,N_1754);
or U2448 (N_2448,N_1555,N_1515);
nand U2449 (N_2449,N_1516,N_1899);
nor U2450 (N_2450,N_1641,N_1655);
and U2451 (N_2451,N_1692,N_1701);
nand U2452 (N_2452,N_1723,N_1952);
nor U2453 (N_2453,N_1602,N_1704);
xor U2454 (N_2454,N_1875,N_1598);
or U2455 (N_2455,N_1990,N_1771);
nand U2456 (N_2456,N_1689,N_1959);
nand U2457 (N_2457,N_1839,N_1699);
and U2458 (N_2458,N_1542,N_1961);
and U2459 (N_2459,N_1555,N_1967);
xor U2460 (N_2460,N_1819,N_1799);
nand U2461 (N_2461,N_1890,N_1929);
nor U2462 (N_2462,N_1817,N_1978);
and U2463 (N_2463,N_1856,N_1776);
or U2464 (N_2464,N_1910,N_1802);
nor U2465 (N_2465,N_1759,N_1961);
or U2466 (N_2466,N_1631,N_1753);
nor U2467 (N_2467,N_1740,N_1500);
and U2468 (N_2468,N_1645,N_1859);
nor U2469 (N_2469,N_1553,N_1866);
nor U2470 (N_2470,N_1858,N_1720);
nand U2471 (N_2471,N_1872,N_1503);
nor U2472 (N_2472,N_1830,N_1984);
or U2473 (N_2473,N_1804,N_1521);
nor U2474 (N_2474,N_1817,N_1902);
and U2475 (N_2475,N_1864,N_1730);
nor U2476 (N_2476,N_1815,N_1891);
nand U2477 (N_2477,N_1515,N_1510);
nor U2478 (N_2478,N_1521,N_1720);
and U2479 (N_2479,N_1605,N_1862);
or U2480 (N_2480,N_1700,N_1620);
nand U2481 (N_2481,N_1542,N_1762);
or U2482 (N_2482,N_1729,N_1625);
xnor U2483 (N_2483,N_1551,N_1944);
and U2484 (N_2484,N_1916,N_1778);
nand U2485 (N_2485,N_1531,N_1807);
and U2486 (N_2486,N_1769,N_1884);
nor U2487 (N_2487,N_1756,N_1972);
xor U2488 (N_2488,N_1866,N_1731);
nand U2489 (N_2489,N_1873,N_1886);
and U2490 (N_2490,N_1532,N_1756);
nor U2491 (N_2491,N_1703,N_1741);
xor U2492 (N_2492,N_1530,N_1727);
nor U2493 (N_2493,N_1727,N_1980);
xor U2494 (N_2494,N_1825,N_1969);
xor U2495 (N_2495,N_1582,N_1824);
nor U2496 (N_2496,N_1786,N_1870);
nor U2497 (N_2497,N_1501,N_1560);
or U2498 (N_2498,N_1855,N_1743);
nor U2499 (N_2499,N_1741,N_1623);
nand U2500 (N_2500,N_2158,N_2318);
xnor U2501 (N_2501,N_2303,N_2136);
xor U2502 (N_2502,N_2164,N_2347);
nand U2503 (N_2503,N_2448,N_2041);
nor U2504 (N_2504,N_2371,N_2001);
nor U2505 (N_2505,N_2081,N_2422);
and U2506 (N_2506,N_2152,N_2431);
nand U2507 (N_2507,N_2178,N_2101);
or U2508 (N_2508,N_2295,N_2102);
nor U2509 (N_2509,N_2380,N_2486);
or U2510 (N_2510,N_2415,N_2378);
and U2511 (N_2511,N_2266,N_2096);
or U2512 (N_2512,N_2079,N_2269);
nor U2513 (N_2513,N_2206,N_2416);
nor U2514 (N_2514,N_2302,N_2449);
xor U2515 (N_2515,N_2377,N_2012);
or U2516 (N_2516,N_2032,N_2019);
or U2517 (N_2517,N_2260,N_2381);
and U2518 (N_2518,N_2350,N_2367);
nor U2519 (N_2519,N_2296,N_2224);
nor U2520 (N_2520,N_2157,N_2087);
xor U2521 (N_2521,N_2268,N_2360);
nand U2522 (N_2522,N_2006,N_2361);
nand U2523 (N_2523,N_2015,N_2300);
nor U2524 (N_2524,N_2163,N_2310);
or U2525 (N_2525,N_2290,N_2446);
or U2526 (N_2526,N_2483,N_2423);
and U2527 (N_2527,N_2090,N_2430);
nor U2528 (N_2528,N_2344,N_2452);
or U2529 (N_2529,N_2281,N_2166);
nor U2530 (N_2530,N_2043,N_2459);
and U2531 (N_2531,N_2306,N_2405);
or U2532 (N_2532,N_2257,N_2485);
xor U2533 (N_2533,N_2258,N_2141);
nor U2534 (N_2534,N_2403,N_2146);
nand U2535 (N_2535,N_2017,N_2174);
nor U2536 (N_2536,N_2467,N_2180);
or U2537 (N_2537,N_2330,N_2168);
nand U2538 (N_2538,N_2011,N_2428);
or U2539 (N_2539,N_2433,N_2481);
nor U2540 (N_2540,N_2442,N_2341);
and U2541 (N_2541,N_2273,N_2272);
or U2542 (N_2542,N_2456,N_2349);
nand U2543 (N_2543,N_2143,N_2264);
or U2544 (N_2544,N_2196,N_2280);
nor U2545 (N_2545,N_2394,N_2155);
nor U2546 (N_2546,N_2248,N_2104);
or U2547 (N_2547,N_2319,N_2128);
nand U2548 (N_2548,N_2308,N_2169);
xnor U2549 (N_2549,N_2094,N_2470);
xor U2550 (N_2550,N_2228,N_2355);
and U2551 (N_2551,N_2004,N_2005);
nand U2552 (N_2552,N_2251,N_2261);
xor U2553 (N_2553,N_2401,N_2109);
nand U2554 (N_2554,N_2199,N_2255);
nand U2555 (N_2555,N_2425,N_2201);
nand U2556 (N_2556,N_2484,N_2133);
nor U2557 (N_2557,N_2082,N_2029);
xor U2558 (N_2558,N_2322,N_2444);
or U2559 (N_2559,N_2490,N_2263);
and U2560 (N_2560,N_2131,N_2333);
and U2561 (N_2561,N_2307,N_2020);
and U2562 (N_2562,N_2114,N_2050);
xor U2563 (N_2563,N_2217,N_2348);
or U2564 (N_2564,N_2439,N_2288);
xnor U2565 (N_2565,N_2235,N_2031);
nand U2566 (N_2566,N_2060,N_2223);
nor U2567 (N_2567,N_2135,N_2399);
or U2568 (N_2568,N_2250,N_2113);
nand U2569 (N_2569,N_2071,N_2085);
xnor U2570 (N_2570,N_2398,N_2480);
xor U2571 (N_2571,N_2025,N_2320);
or U2572 (N_2572,N_2154,N_2412);
xor U2573 (N_2573,N_2373,N_2216);
xor U2574 (N_2574,N_2495,N_2191);
xor U2575 (N_2575,N_2215,N_2368);
nor U2576 (N_2576,N_2353,N_2345);
and U2577 (N_2577,N_2427,N_2222);
nand U2578 (N_2578,N_2179,N_2325);
nand U2579 (N_2579,N_2065,N_2159);
and U2580 (N_2580,N_2498,N_2241);
and U2581 (N_2581,N_2124,N_2386);
and U2582 (N_2582,N_2331,N_2336);
nand U2583 (N_2583,N_2132,N_2332);
or U2584 (N_2584,N_2406,N_2384);
nor U2585 (N_2585,N_2207,N_2026);
nand U2586 (N_2586,N_2342,N_2461);
nand U2587 (N_2587,N_2095,N_2013);
and U2588 (N_2588,N_2238,N_2002);
and U2589 (N_2589,N_2186,N_2089);
nand U2590 (N_2590,N_2148,N_2183);
nor U2591 (N_2591,N_2172,N_2057);
or U2592 (N_2592,N_2462,N_2203);
xor U2593 (N_2593,N_2229,N_2334);
xnor U2594 (N_2594,N_2056,N_2118);
and U2595 (N_2595,N_2083,N_2441);
xor U2596 (N_2596,N_2115,N_2225);
and U2597 (N_2597,N_2497,N_2291);
nor U2598 (N_2598,N_2039,N_2070);
nand U2599 (N_2599,N_2458,N_2077);
and U2600 (N_2600,N_2468,N_2010);
or U2601 (N_2601,N_2088,N_2016);
and U2602 (N_2602,N_2123,N_2033);
nor U2603 (N_2603,N_2297,N_2121);
nor U2604 (N_2604,N_2080,N_2093);
nand U2605 (N_2605,N_2364,N_2335);
or U2606 (N_2606,N_2282,N_2022);
xnor U2607 (N_2607,N_2482,N_2054);
or U2608 (N_2608,N_2438,N_2034);
xnor U2609 (N_2609,N_2429,N_2110);
nor U2610 (N_2610,N_2214,N_2219);
and U2611 (N_2611,N_2202,N_2383);
or U2612 (N_2612,N_2313,N_2091);
xor U2613 (N_2613,N_2086,N_2359);
nor U2614 (N_2614,N_2126,N_2193);
or U2615 (N_2615,N_2052,N_2173);
or U2616 (N_2616,N_2245,N_2063);
nor U2617 (N_2617,N_2287,N_2140);
nor U2618 (N_2618,N_2242,N_2098);
nor U2619 (N_2619,N_2137,N_2471);
nor U2620 (N_2620,N_2233,N_2189);
or U2621 (N_2621,N_2315,N_2419);
or U2622 (N_2622,N_2387,N_2473);
or U2623 (N_2623,N_2460,N_2030);
and U2624 (N_2624,N_2323,N_2413);
nor U2625 (N_2625,N_2477,N_2418);
nand U2626 (N_2626,N_2144,N_2036);
xnor U2627 (N_2627,N_2312,N_2211);
nand U2628 (N_2628,N_2254,N_2227);
nand U2629 (N_2629,N_2329,N_2494);
and U2630 (N_2630,N_2309,N_2119);
xnor U2631 (N_2631,N_2125,N_2177);
nand U2632 (N_2632,N_2393,N_2051);
nor U2633 (N_2633,N_2145,N_2165);
nor U2634 (N_2634,N_2479,N_2321);
or U2635 (N_2635,N_2221,N_2392);
and U2636 (N_2636,N_2058,N_2437);
nor U2637 (N_2637,N_2424,N_2075);
nor U2638 (N_2638,N_2105,N_2374);
nor U2639 (N_2639,N_2084,N_2338);
nor U2640 (N_2640,N_2073,N_2003);
nor U2641 (N_2641,N_2408,N_2175);
nand U2642 (N_2642,N_2220,N_2390);
nand U2643 (N_2643,N_2234,N_2443);
xnor U2644 (N_2644,N_2259,N_2018);
xnor U2645 (N_2645,N_2324,N_2407);
or U2646 (N_2646,N_2038,N_2369);
nor U2647 (N_2647,N_2314,N_2044);
xor U2648 (N_2648,N_2279,N_2277);
nand U2649 (N_2649,N_2362,N_2357);
nor U2650 (N_2650,N_2046,N_2187);
or U2651 (N_2651,N_2205,N_2055);
and U2652 (N_2652,N_2372,N_2346);
xnor U2653 (N_2653,N_2311,N_2301);
xor U2654 (N_2654,N_2226,N_2100);
and U2655 (N_2655,N_2466,N_2354);
xor U2656 (N_2656,N_2487,N_2198);
and U2657 (N_2657,N_2370,N_2240);
and U2658 (N_2658,N_2385,N_2162);
nor U2659 (N_2659,N_2210,N_2435);
nor U2660 (N_2660,N_2108,N_2270);
nand U2661 (N_2661,N_2213,N_2363);
xnor U2662 (N_2662,N_2375,N_2286);
nor U2663 (N_2663,N_2298,N_2097);
nand U2664 (N_2664,N_2299,N_2129);
or U2665 (N_2665,N_2285,N_2496);
and U2666 (N_2666,N_2457,N_2293);
xor U2667 (N_2667,N_2000,N_2142);
nand U2668 (N_2668,N_2171,N_2426);
xnor U2669 (N_2669,N_2014,N_2305);
xor U2670 (N_2670,N_2064,N_2023);
or U2671 (N_2671,N_2184,N_2409);
xor U2672 (N_2672,N_2289,N_2062);
xnor U2673 (N_2673,N_2404,N_2436);
xor U2674 (N_2674,N_2116,N_2474);
or U2675 (N_2675,N_2076,N_2343);
nand U2676 (N_2676,N_2068,N_2134);
xor U2677 (N_2677,N_2472,N_2351);
nand U2678 (N_2678,N_2249,N_2190);
nand U2679 (N_2679,N_2037,N_2489);
xnor U2680 (N_2680,N_2035,N_2476);
nor U2681 (N_2681,N_2265,N_2061);
nand U2682 (N_2682,N_2067,N_2192);
or U2683 (N_2683,N_2453,N_2161);
and U2684 (N_2684,N_2316,N_2130);
nor U2685 (N_2685,N_2111,N_2493);
nor U2686 (N_2686,N_2440,N_2465);
and U2687 (N_2687,N_2278,N_2147);
or U2688 (N_2688,N_2139,N_2151);
and U2689 (N_2689,N_2382,N_2150);
or U2690 (N_2690,N_2042,N_2231);
nand U2691 (N_2691,N_2262,N_2391);
and U2692 (N_2692,N_2078,N_2317);
xor U2693 (N_2693,N_2209,N_2117);
or U2694 (N_2694,N_2247,N_2092);
or U2695 (N_2695,N_2195,N_2112);
nor U2696 (N_2696,N_2007,N_2421);
and U2697 (N_2697,N_2120,N_2284);
xor U2698 (N_2698,N_2358,N_2454);
nor U2699 (N_2699,N_2417,N_2397);
nor U2700 (N_2700,N_2246,N_2045);
nand U2701 (N_2701,N_2326,N_2138);
xnor U2702 (N_2702,N_2200,N_2072);
and U2703 (N_2703,N_2339,N_2182);
nand U2704 (N_2704,N_2066,N_2244);
and U2705 (N_2705,N_2283,N_2432);
nand U2706 (N_2706,N_2376,N_2069);
and U2707 (N_2707,N_2469,N_2450);
xnor U2708 (N_2708,N_2356,N_2451);
xnor U2709 (N_2709,N_2176,N_2181);
nand U2710 (N_2710,N_2271,N_2239);
nor U2711 (N_2711,N_2153,N_2021);
or U2712 (N_2712,N_2099,N_2294);
nand U2713 (N_2713,N_2107,N_2388);
xnor U2714 (N_2714,N_2028,N_2160);
and U2715 (N_2715,N_2366,N_2127);
or U2716 (N_2716,N_2274,N_2414);
or U2717 (N_2717,N_2024,N_2243);
nand U2718 (N_2718,N_2395,N_2420);
xnor U2719 (N_2719,N_2047,N_2252);
and U2720 (N_2720,N_2237,N_2411);
or U2721 (N_2721,N_2156,N_2267);
nand U2722 (N_2722,N_2204,N_2027);
xnor U2723 (N_2723,N_2304,N_2389);
xnor U2724 (N_2724,N_2103,N_2253);
and U2725 (N_2725,N_2276,N_2122);
nand U2726 (N_2726,N_2464,N_2410);
xnor U2727 (N_2727,N_2048,N_2230);
and U2728 (N_2728,N_2167,N_2059);
nor U2729 (N_2729,N_2492,N_2491);
or U2730 (N_2730,N_2396,N_2188);
and U2731 (N_2731,N_2434,N_2379);
nor U2732 (N_2732,N_2340,N_2455);
and U2733 (N_2733,N_2402,N_2212);
or U2734 (N_2734,N_2365,N_2208);
and U2735 (N_2735,N_2218,N_2049);
and U2736 (N_2736,N_2040,N_2499);
nand U2737 (N_2737,N_2327,N_2236);
or U2738 (N_2738,N_2009,N_2488);
and U2739 (N_2739,N_2463,N_2475);
nand U2740 (N_2740,N_2328,N_2337);
and U2741 (N_2741,N_2170,N_2149);
xnor U2742 (N_2742,N_2275,N_2106);
nand U2743 (N_2743,N_2053,N_2352);
xor U2744 (N_2744,N_2232,N_2074);
and U2745 (N_2745,N_2400,N_2194);
nand U2746 (N_2746,N_2008,N_2447);
nor U2747 (N_2747,N_2292,N_2185);
or U2748 (N_2748,N_2445,N_2478);
xor U2749 (N_2749,N_2256,N_2197);
xnor U2750 (N_2750,N_2179,N_2449);
nand U2751 (N_2751,N_2432,N_2041);
nor U2752 (N_2752,N_2195,N_2410);
nand U2753 (N_2753,N_2411,N_2399);
and U2754 (N_2754,N_2330,N_2122);
nor U2755 (N_2755,N_2302,N_2384);
and U2756 (N_2756,N_2316,N_2336);
nor U2757 (N_2757,N_2399,N_2118);
and U2758 (N_2758,N_2192,N_2130);
nand U2759 (N_2759,N_2330,N_2470);
and U2760 (N_2760,N_2325,N_2187);
or U2761 (N_2761,N_2424,N_2464);
or U2762 (N_2762,N_2463,N_2451);
and U2763 (N_2763,N_2454,N_2322);
nor U2764 (N_2764,N_2128,N_2276);
xor U2765 (N_2765,N_2036,N_2465);
nand U2766 (N_2766,N_2150,N_2375);
nand U2767 (N_2767,N_2187,N_2139);
xnor U2768 (N_2768,N_2382,N_2421);
nor U2769 (N_2769,N_2466,N_2344);
nand U2770 (N_2770,N_2008,N_2082);
or U2771 (N_2771,N_2281,N_2245);
or U2772 (N_2772,N_2415,N_2028);
nand U2773 (N_2773,N_2253,N_2248);
or U2774 (N_2774,N_2289,N_2406);
nor U2775 (N_2775,N_2040,N_2304);
xor U2776 (N_2776,N_2296,N_2002);
nand U2777 (N_2777,N_2411,N_2046);
nand U2778 (N_2778,N_2222,N_2002);
or U2779 (N_2779,N_2376,N_2280);
nand U2780 (N_2780,N_2293,N_2267);
and U2781 (N_2781,N_2183,N_2479);
and U2782 (N_2782,N_2103,N_2066);
and U2783 (N_2783,N_2276,N_2147);
nand U2784 (N_2784,N_2299,N_2347);
or U2785 (N_2785,N_2016,N_2106);
or U2786 (N_2786,N_2053,N_2322);
xnor U2787 (N_2787,N_2250,N_2173);
and U2788 (N_2788,N_2430,N_2307);
and U2789 (N_2789,N_2238,N_2246);
or U2790 (N_2790,N_2436,N_2217);
nand U2791 (N_2791,N_2330,N_2484);
nor U2792 (N_2792,N_2399,N_2288);
nor U2793 (N_2793,N_2025,N_2324);
nand U2794 (N_2794,N_2164,N_2018);
nand U2795 (N_2795,N_2248,N_2415);
and U2796 (N_2796,N_2190,N_2403);
xnor U2797 (N_2797,N_2071,N_2133);
and U2798 (N_2798,N_2141,N_2091);
or U2799 (N_2799,N_2331,N_2129);
or U2800 (N_2800,N_2376,N_2091);
nand U2801 (N_2801,N_2318,N_2359);
or U2802 (N_2802,N_2060,N_2472);
and U2803 (N_2803,N_2052,N_2408);
nor U2804 (N_2804,N_2440,N_2463);
or U2805 (N_2805,N_2092,N_2010);
nand U2806 (N_2806,N_2343,N_2253);
xnor U2807 (N_2807,N_2491,N_2074);
or U2808 (N_2808,N_2493,N_2350);
or U2809 (N_2809,N_2203,N_2049);
nand U2810 (N_2810,N_2438,N_2121);
or U2811 (N_2811,N_2481,N_2465);
xnor U2812 (N_2812,N_2056,N_2124);
xor U2813 (N_2813,N_2439,N_2398);
xor U2814 (N_2814,N_2113,N_2066);
xnor U2815 (N_2815,N_2175,N_2469);
or U2816 (N_2816,N_2200,N_2287);
and U2817 (N_2817,N_2046,N_2040);
xnor U2818 (N_2818,N_2145,N_2255);
and U2819 (N_2819,N_2053,N_2429);
nand U2820 (N_2820,N_2425,N_2393);
nor U2821 (N_2821,N_2166,N_2088);
xnor U2822 (N_2822,N_2344,N_2208);
and U2823 (N_2823,N_2467,N_2490);
nand U2824 (N_2824,N_2000,N_2359);
or U2825 (N_2825,N_2455,N_2315);
nor U2826 (N_2826,N_2197,N_2470);
xnor U2827 (N_2827,N_2460,N_2238);
nor U2828 (N_2828,N_2316,N_2344);
xor U2829 (N_2829,N_2263,N_2151);
or U2830 (N_2830,N_2220,N_2208);
nor U2831 (N_2831,N_2442,N_2104);
nand U2832 (N_2832,N_2431,N_2202);
nand U2833 (N_2833,N_2060,N_2101);
nand U2834 (N_2834,N_2324,N_2365);
xnor U2835 (N_2835,N_2194,N_2037);
and U2836 (N_2836,N_2481,N_2081);
nor U2837 (N_2837,N_2236,N_2362);
and U2838 (N_2838,N_2219,N_2423);
and U2839 (N_2839,N_2220,N_2145);
and U2840 (N_2840,N_2478,N_2321);
nor U2841 (N_2841,N_2123,N_2339);
nand U2842 (N_2842,N_2406,N_2261);
nand U2843 (N_2843,N_2023,N_2145);
or U2844 (N_2844,N_2336,N_2091);
xor U2845 (N_2845,N_2004,N_2240);
nand U2846 (N_2846,N_2450,N_2202);
or U2847 (N_2847,N_2163,N_2450);
and U2848 (N_2848,N_2410,N_2324);
nand U2849 (N_2849,N_2389,N_2069);
nand U2850 (N_2850,N_2084,N_2391);
or U2851 (N_2851,N_2259,N_2082);
nand U2852 (N_2852,N_2244,N_2241);
xor U2853 (N_2853,N_2111,N_2205);
nor U2854 (N_2854,N_2412,N_2275);
nor U2855 (N_2855,N_2439,N_2176);
nand U2856 (N_2856,N_2376,N_2105);
or U2857 (N_2857,N_2394,N_2401);
nand U2858 (N_2858,N_2380,N_2433);
or U2859 (N_2859,N_2091,N_2449);
xor U2860 (N_2860,N_2373,N_2111);
or U2861 (N_2861,N_2147,N_2218);
or U2862 (N_2862,N_2029,N_2352);
xnor U2863 (N_2863,N_2453,N_2325);
and U2864 (N_2864,N_2358,N_2478);
nand U2865 (N_2865,N_2487,N_2482);
xnor U2866 (N_2866,N_2013,N_2408);
nor U2867 (N_2867,N_2448,N_2031);
and U2868 (N_2868,N_2024,N_2460);
and U2869 (N_2869,N_2190,N_2340);
xor U2870 (N_2870,N_2004,N_2426);
nor U2871 (N_2871,N_2145,N_2094);
xor U2872 (N_2872,N_2442,N_2455);
nand U2873 (N_2873,N_2093,N_2467);
and U2874 (N_2874,N_2222,N_2071);
nor U2875 (N_2875,N_2188,N_2217);
nand U2876 (N_2876,N_2189,N_2004);
and U2877 (N_2877,N_2167,N_2317);
nor U2878 (N_2878,N_2493,N_2186);
or U2879 (N_2879,N_2197,N_2391);
nor U2880 (N_2880,N_2220,N_2060);
and U2881 (N_2881,N_2431,N_2295);
nor U2882 (N_2882,N_2038,N_2456);
nor U2883 (N_2883,N_2375,N_2332);
xnor U2884 (N_2884,N_2426,N_2438);
xnor U2885 (N_2885,N_2096,N_2348);
nor U2886 (N_2886,N_2486,N_2478);
nand U2887 (N_2887,N_2489,N_2348);
nand U2888 (N_2888,N_2496,N_2319);
xor U2889 (N_2889,N_2406,N_2114);
nor U2890 (N_2890,N_2361,N_2327);
nor U2891 (N_2891,N_2460,N_2154);
nand U2892 (N_2892,N_2197,N_2338);
nand U2893 (N_2893,N_2107,N_2159);
or U2894 (N_2894,N_2282,N_2075);
or U2895 (N_2895,N_2133,N_2129);
or U2896 (N_2896,N_2069,N_2090);
nand U2897 (N_2897,N_2061,N_2100);
nand U2898 (N_2898,N_2364,N_2331);
nor U2899 (N_2899,N_2400,N_2113);
nand U2900 (N_2900,N_2201,N_2310);
nand U2901 (N_2901,N_2328,N_2048);
or U2902 (N_2902,N_2437,N_2029);
and U2903 (N_2903,N_2433,N_2136);
xnor U2904 (N_2904,N_2051,N_2342);
and U2905 (N_2905,N_2479,N_2021);
and U2906 (N_2906,N_2352,N_2010);
and U2907 (N_2907,N_2346,N_2051);
or U2908 (N_2908,N_2491,N_2035);
or U2909 (N_2909,N_2349,N_2185);
xnor U2910 (N_2910,N_2465,N_2410);
nand U2911 (N_2911,N_2114,N_2020);
xor U2912 (N_2912,N_2261,N_2041);
and U2913 (N_2913,N_2493,N_2282);
and U2914 (N_2914,N_2355,N_2459);
and U2915 (N_2915,N_2452,N_2434);
xnor U2916 (N_2916,N_2158,N_2227);
nor U2917 (N_2917,N_2311,N_2381);
nor U2918 (N_2918,N_2216,N_2133);
xor U2919 (N_2919,N_2009,N_2241);
xor U2920 (N_2920,N_2039,N_2233);
nor U2921 (N_2921,N_2468,N_2236);
or U2922 (N_2922,N_2287,N_2214);
nand U2923 (N_2923,N_2207,N_2425);
xnor U2924 (N_2924,N_2071,N_2092);
nor U2925 (N_2925,N_2188,N_2196);
nor U2926 (N_2926,N_2418,N_2271);
nor U2927 (N_2927,N_2126,N_2408);
and U2928 (N_2928,N_2147,N_2389);
nand U2929 (N_2929,N_2204,N_2041);
nor U2930 (N_2930,N_2278,N_2377);
nand U2931 (N_2931,N_2171,N_2150);
nor U2932 (N_2932,N_2009,N_2282);
or U2933 (N_2933,N_2283,N_2195);
nor U2934 (N_2934,N_2009,N_2162);
nor U2935 (N_2935,N_2222,N_2112);
and U2936 (N_2936,N_2321,N_2489);
xnor U2937 (N_2937,N_2174,N_2202);
nor U2938 (N_2938,N_2260,N_2368);
nor U2939 (N_2939,N_2129,N_2385);
nand U2940 (N_2940,N_2118,N_2062);
nor U2941 (N_2941,N_2424,N_2139);
or U2942 (N_2942,N_2199,N_2016);
nand U2943 (N_2943,N_2440,N_2473);
nor U2944 (N_2944,N_2485,N_2083);
nand U2945 (N_2945,N_2160,N_2198);
or U2946 (N_2946,N_2317,N_2289);
nor U2947 (N_2947,N_2318,N_2066);
nor U2948 (N_2948,N_2276,N_2423);
and U2949 (N_2949,N_2221,N_2449);
nand U2950 (N_2950,N_2072,N_2013);
or U2951 (N_2951,N_2040,N_2001);
xnor U2952 (N_2952,N_2335,N_2432);
and U2953 (N_2953,N_2258,N_2465);
xor U2954 (N_2954,N_2082,N_2207);
nand U2955 (N_2955,N_2293,N_2327);
xor U2956 (N_2956,N_2461,N_2284);
or U2957 (N_2957,N_2102,N_2376);
nor U2958 (N_2958,N_2418,N_2333);
and U2959 (N_2959,N_2466,N_2379);
nand U2960 (N_2960,N_2358,N_2198);
nor U2961 (N_2961,N_2392,N_2343);
or U2962 (N_2962,N_2195,N_2197);
xor U2963 (N_2963,N_2113,N_2158);
xor U2964 (N_2964,N_2325,N_2348);
xor U2965 (N_2965,N_2407,N_2461);
or U2966 (N_2966,N_2064,N_2460);
xor U2967 (N_2967,N_2362,N_2400);
and U2968 (N_2968,N_2024,N_2233);
or U2969 (N_2969,N_2311,N_2141);
and U2970 (N_2970,N_2313,N_2323);
nand U2971 (N_2971,N_2051,N_2101);
nor U2972 (N_2972,N_2334,N_2218);
nand U2973 (N_2973,N_2212,N_2268);
and U2974 (N_2974,N_2004,N_2448);
xnor U2975 (N_2975,N_2428,N_2101);
nor U2976 (N_2976,N_2003,N_2229);
nor U2977 (N_2977,N_2453,N_2272);
nand U2978 (N_2978,N_2225,N_2039);
xnor U2979 (N_2979,N_2417,N_2005);
nor U2980 (N_2980,N_2211,N_2411);
nand U2981 (N_2981,N_2221,N_2123);
nor U2982 (N_2982,N_2000,N_2057);
or U2983 (N_2983,N_2431,N_2200);
and U2984 (N_2984,N_2335,N_2338);
and U2985 (N_2985,N_2348,N_2043);
xor U2986 (N_2986,N_2273,N_2091);
and U2987 (N_2987,N_2325,N_2226);
and U2988 (N_2988,N_2495,N_2000);
and U2989 (N_2989,N_2488,N_2189);
or U2990 (N_2990,N_2021,N_2067);
nand U2991 (N_2991,N_2308,N_2071);
nor U2992 (N_2992,N_2232,N_2278);
xor U2993 (N_2993,N_2060,N_2156);
and U2994 (N_2994,N_2201,N_2301);
nor U2995 (N_2995,N_2491,N_2118);
or U2996 (N_2996,N_2242,N_2458);
or U2997 (N_2997,N_2115,N_2143);
or U2998 (N_2998,N_2186,N_2149);
and U2999 (N_2999,N_2042,N_2282);
or U3000 (N_3000,N_2572,N_2605);
nor U3001 (N_3001,N_2684,N_2922);
nor U3002 (N_3002,N_2784,N_2722);
nor U3003 (N_3003,N_2614,N_2942);
or U3004 (N_3004,N_2851,N_2612);
xnor U3005 (N_3005,N_2693,N_2850);
and U3006 (N_3006,N_2628,N_2621);
or U3007 (N_3007,N_2772,N_2787);
nor U3008 (N_3008,N_2582,N_2640);
or U3009 (N_3009,N_2530,N_2747);
or U3010 (N_3010,N_2812,N_2541);
xnor U3011 (N_3011,N_2689,N_2741);
and U3012 (N_3012,N_2529,N_2798);
nor U3013 (N_3013,N_2597,N_2762);
nor U3014 (N_3014,N_2910,N_2944);
nor U3015 (N_3015,N_2828,N_2859);
nand U3016 (N_3016,N_2526,N_2724);
xor U3017 (N_3017,N_2646,N_2679);
nand U3018 (N_3018,N_2977,N_2583);
nand U3019 (N_3019,N_2979,N_2745);
xor U3020 (N_3020,N_2904,N_2706);
nand U3021 (N_3021,N_2815,N_2600);
nand U3022 (N_3022,N_2726,N_2575);
and U3023 (N_3023,N_2748,N_2734);
or U3024 (N_3024,N_2873,N_2554);
nand U3025 (N_3025,N_2644,N_2766);
and U3026 (N_3026,N_2622,N_2744);
and U3027 (N_3027,N_2842,N_2522);
nand U3028 (N_3028,N_2774,N_2682);
and U3029 (N_3029,N_2611,N_2671);
nor U3030 (N_3030,N_2545,N_2581);
nor U3031 (N_3031,N_2564,N_2585);
xor U3032 (N_3032,N_2567,N_2672);
or U3033 (N_3033,N_2801,N_2932);
xnor U3034 (N_3034,N_2771,N_2565);
and U3035 (N_3035,N_2894,N_2691);
nand U3036 (N_3036,N_2651,N_2685);
or U3037 (N_3037,N_2764,N_2665);
nand U3038 (N_3038,N_2916,N_2725);
nor U3039 (N_3039,N_2702,N_2900);
nor U3040 (N_3040,N_2843,N_2811);
xor U3041 (N_3041,N_2964,N_2837);
nor U3042 (N_3042,N_2559,N_2946);
and U3043 (N_3043,N_2561,N_2872);
nand U3044 (N_3044,N_2666,N_2729);
and U3045 (N_3045,N_2603,N_2550);
xnor U3046 (N_3046,N_2958,N_2524);
nor U3047 (N_3047,N_2794,N_2905);
or U3048 (N_3048,N_2928,N_2678);
nor U3049 (N_3049,N_2997,N_2508);
nand U3050 (N_3050,N_2710,N_2949);
nor U3051 (N_3051,N_2841,N_2765);
and U3052 (N_3052,N_2985,N_2831);
nand U3053 (N_3053,N_2505,N_2819);
xnor U3054 (N_3054,N_2845,N_2566);
nor U3055 (N_3055,N_2519,N_2950);
nor U3056 (N_3056,N_2832,N_2971);
and U3057 (N_3057,N_2589,N_2986);
nor U3058 (N_3058,N_2601,N_2968);
or U3059 (N_3059,N_2763,N_2624);
and U3060 (N_3060,N_2629,N_2535);
and U3061 (N_3061,N_2556,N_2770);
and U3062 (N_3062,N_2929,N_2675);
and U3063 (N_3063,N_2827,N_2750);
nand U3064 (N_3064,N_2551,N_2751);
and U3065 (N_3065,N_2733,N_2876);
nand U3066 (N_3066,N_2547,N_2890);
or U3067 (N_3067,N_2538,N_2783);
and U3068 (N_3068,N_2793,N_2777);
and U3069 (N_3069,N_2925,N_2506);
or U3070 (N_3070,N_2604,N_2655);
or U3071 (N_3071,N_2715,N_2808);
and U3072 (N_3072,N_2934,N_2716);
nand U3073 (N_3073,N_2849,N_2947);
nand U3074 (N_3074,N_2713,N_2768);
or U3075 (N_3075,N_2643,N_2857);
xor U3076 (N_3076,N_2983,N_2563);
nor U3077 (N_3077,N_2534,N_2790);
nand U3078 (N_3078,N_2630,N_2926);
nor U3079 (N_3079,N_2825,N_2659);
nor U3080 (N_3080,N_2860,N_2939);
and U3081 (N_3081,N_2711,N_2924);
and U3082 (N_3082,N_2754,N_2776);
nor U3083 (N_3083,N_2502,N_2573);
or U3084 (N_3084,N_2952,N_2978);
and U3085 (N_3085,N_2806,N_2697);
nand U3086 (N_3086,N_2858,N_2680);
xnor U3087 (N_3087,N_2528,N_2999);
xnor U3088 (N_3088,N_2855,N_2636);
or U3089 (N_3089,N_2536,N_2609);
xnor U3090 (N_3090,N_2778,N_2627);
nand U3091 (N_3091,N_2795,N_2881);
and U3092 (N_3092,N_2661,N_2769);
nor U3093 (N_3093,N_2595,N_2759);
xnor U3094 (N_3094,N_2948,N_2513);
xnor U3095 (N_3095,N_2911,N_2560);
nand U3096 (N_3096,N_2512,N_2633);
and U3097 (N_3097,N_2515,N_2995);
or U3098 (N_3098,N_2520,N_2931);
and U3099 (N_3099,N_2521,N_2791);
or U3100 (N_3100,N_2623,N_2533);
nand U3101 (N_3101,N_2617,N_2730);
nor U3102 (N_3102,N_2935,N_2915);
or U3103 (N_3103,N_2933,N_2940);
nand U3104 (N_3104,N_2829,N_2917);
or U3105 (N_3105,N_2509,N_2516);
nand U3106 (N_3106,N_2525,N_2818);
and U3107 (N_3107,N_2886,N_2518);
nor U3108 (N_3108,N_2960,N_2688);
nand U3109 (N_3109,N_2738,N_2957);
or U3110 (N_3110,N_2606,N_2782);
nor U3111 (N_3111,N_2714,N_2761);
or U3112 (N_3112,N_2820,N_2891);
nor U3113 (N_3113,N_2638,N_2861);
nand U3114 (N_3114,N_2781,N_2826);
xor U3115 (N_3115,N_2898,N_2871);
nand U3116 (N_3116,N_2709,N_2959);
or U3117 (N_3117,N_2830,N_2936);
nand U3118 (N_3118,N_2591,N_2718);
and U3119 (N_3119,N_2846,N_2896);
or U3120 (N_3120,N_2884,N_2681);
nand U3121 (N_3121,N_2874,N_2882);
xor U3122 (N_3122,N_2887,N_2993);
xor U3123 (N_3123,N_2531,N_2792);
nor U3124 (N_3124,N_2739,N_2988);
nand U3125 (N_3125,N_2517,N_2954);
nor U3126 (N_3126,N_2727,N_2635);
xnor U3127 (N_3127,N_2821,N_2523);
and U3128 (N_3128,N_2692,N_2892);
xor U3129 (N_3129,N_2967,N_2943);
nand U3130 (N_3130,N_2824,N_2704);
xnor U3131 (N_3131,N_2568,N_2945);
and U3132 (N_3132,N_2695,N_2642);
or U3133 (N_3133,N_2576,N_2987);
xor U3134 (N_3134,N_2866,N_2619);
or U3135 (N_3135,N_2880,N_2719);
nand U3136 (N_3136,N_2863,N_2869);
and U3137 (N_3137,N_2833,N_2594);
xor U3138 (N_3138,N_2854,N_2558);
nor U3139 (N_3139,N_2970,N_2647);
nand U3140 (N_3140,N_2598,N_2779);
and U3141 (N_3141,N_2639,N_2885);
xnor U3142 (N_3142,N_2804,N_2834);
xor U3143 (N_3143,N_2701,N_2656);
nor U3144 (N_3144,N_2599,N_2789);
nor U3145 (N_3145,N_2879,N_2590);
nand U3146 (N_3146,N_2717,N_2721);
and U3147 (N_3147,N_2735,N_2813);
xor U3148 (N_3148,N_2549,N_2749);
or U3149 (N_3149,N_2976,N_2963);
nor U3150 (N_3150,N_2580,N_2546);
nand U3151 (N_3151,N_2975,N_2980);
and U3152 (N_3152,N_2542,N_2705);
and U3153 (N_3153,N_2908,N_2839);
and U3154 (N_3154,N_2562,N_2867);
or U3155 (N_3155,N_2994,N_2920);
and U3156 (N_3156,N_2586,N_2670);
nor U3157 (N_3157,N_2631,N_2912);
nand U3158 (N_3158,N_2927,N_2760);
nand U3159 (N_3159,N_2785,N_2951);
xor U3160 (N_3160,N_2676,N_2532);
or U3161 (N_3161,N_2955,N_2501);
nor U3162 (N_3162,N_2660,N_2981);
or U3163 (N_3163,N_2853,N_2903);
or U3164 (N_3164,N_2972,N_2984);
xor U3165 (N_3165,N_2543,N_2864);
and U3166 (N_3166,N_2658,N_2579);
nand U3167 (N_3167,N_2596,N_2708);
nor U3168 (N_3168,N_2991,N_2607);
or U3169 (N_3169,N_2743,N_2992);
xor U3170 (N_3170,N_2620,N_2956);
or U3171 (N_3171,N_2897,N_2878);
or U3172 (N_3172,N_2786,N_2856);
nor U3173 (N_3173,N_2756,N_2736);
xor U3174 (N_3174,N_2544,N_2757);
or U3175 (N_3175,N_2571,N_2775);
nor U3176 (N_3176,N_2966,N_2577);
or U3177 (N_3177,N_2570,N_2650);
nand U3178 (N_3178,N_2937,N_2998);
nand U3179 (N_3179,N_2667,N_2652);
nor U3180 (N_3180,N_2755,N_2796);
and U3181 (N_3181,N_2803,N_2847);
xor U3182 (N_3182,N_2923,N_2625);
or U3183 (N_3183,N_2870,N_2868);
or U3184 (N_3184,N_2973,N_2921);
nand U3185 (N_3185,N_2780,N_2626);
xnor U3186 (N_3186,N_2669,N_2698);
or U3187 (N_3187,N_2608,N_2840);
nor U3188 (N_3188,N_2817,N_2503);
xnor U3189 (N_3189,N_2810,N_2555);
nor U3190 (N_3190,N_2888,N_2587);
or U3191 (N_3191,N_2694,N_2909);
nor U3192 (N_3192,N_2664,N_2742);
nand U3193 (N_3193,N_2862,N_2537);
nand U3194 (N_3194,N_2737,N_2654);
nor U3195 (N_3195,N_2641,N_2674);
nor U3196 (N_3196,N_2877,N_2875);
xor U3197 (N_3197,N_2703,N_2696);
or U3198 (N_3198,N_2602,N_2690);
nor U3199 (N_3199,N_2953,N_2919);
nor U3200 (N_3200,N_2788,N_2634);
and U3201 (N_3201,N_2961,N_2901);
and U3202 (N_3202,N_2663,N_2700);
or U3203 (N_3203,N_2557,N_2809);
or U3204 (N_3204,N_2699,N_2800);
xnor U3205 (N_3205,N_2574,N_2687);
or U3206 (N_3206,N_2707,N_2814);
xor U3207 (N_3207,N_2527,N_2773);
or U3208 (N_3208,N_2836,N_2511);
xnor U3209 (N_3209,N_2504,N_2712);
nand U3210 (N_3210,N_2822,N_2683);
and U3211 (N_3211,N_2752,N_2962);
nand U3212 (N_3212,N_2510,N_2982);
nor U3213 (N_3213,N_2720,N_2838);
or U3214 (N_3214,N_2500,N_2740);
nor U3215 (N_3215,N_2823,N_2974);
nand U3216 (N_3216,N_2649,N_2632);
xor U3217 (N_3217,N_2723,N_2507);
nor U3218 (N_3218,N_2889,N_2799);
xor U3219 (N_3219,N_2797,N_2677);
xnor U3220 (N_3220,N_2673,N_2802);
nor U3221 (N_3221,N_2969,N_2835);
and U3222 (N_3222,N_2615,N_2569);
xnor U3223 (N_3223,N_2514,N_2645);
nand U3224 (N_3224,N_2552,N_2657);
xnor U3225 (N_3225,N_2731,N_2805);
nor U3226 (N_3226,N_2893,N_2852);
nand U3227 (N_3227,N_2637,N_2807);
nand U3228 (N_3228,N_2618,N_2653);
nand U3229 (N_3229,N_2914,N_2767);
xnor U3230 (N_3230,N_2592,N_2686);
and U3231 (N_3231,N_2906,N_2553);
or U3232 (N_3232,N_2930,N_2588);
nor U3233 (N_3233,N_2593,N_2753);
and U3234 (N_3234,N_2907,N_2728);
nand U3235 (N_3235,N_2918,N_2913);
nor U3236 (N_3236,N_2539,N_2989);
or U3237 (N_3237,N_2668,N_2662);
nor U3238 (N_3238,N_2844,N_2648);
and U3239 (N_3239,N_2899,N_2816);
and U3240 (N_3240,N_2616,N_2540);
and U3241 (N_3241,N_2584,N_2613);
nand U3242 (N_3242,N_2865,N_2758);
xnor U3243 (N_3243,N_2848,N_2578);
or U3244 (N_3244,N_2895,N_2938);
and U3245 (N_3245,N_2996,N_2965);
or U3246 (N_3246,N_2902,N_2746);
nand U3247 (N_3247,N_2990,N_2732);
nor U3248 (N_3248,N_2941,N_2610);
xor U3249 (N_3249,N_2548,N_2883);
nor U3250 (N_3250,N_2868,N_2664);
or U3251 (N_3251,N_2554,N_2834);
or U3252 (N_3252,N_2508,N_2991);
and U3253 (N_3253,N_2665,N_2705);
or U3254 (N_3254,N_2882,N_2957);
nand U3255 (N_3255,N_2974,N_2790);
and U3256 (N_3256,N_2853,N_2547);
nor U3257 (N_3257,N_2625,N_2771);
and U3258 (N_3258,N_2615,N_2589);
nand U3259 (N_3259,N_2704,N_2724);
and U3260 (N_3260,N_2703,N_2791);
xor U3261 (N_3261,N_2634,N_2822);
xor U3262 (N_3262,N_2931,N_2797);
nand U3263 (N_3263,N_2544,N_2533);
xor U3264 (N_3264,N_2652,N_2686);
nand U3265 (N_3265,N_2566,N_2592);
and U3266 (N_3266,N_2541,N_2932);
nor U3267 (N_3267,N_2835,N_2573);
xnor U3268 (N_3268,N_2835,N_2826);
nand U3269 (N_3269,N_2884,N_2583);
or U3270 (N_3270,N_2814,N_2775);
nor U3271 (N_3271,N_2778,N_2506);
nor U3272 (N_3272,N_2690,N_2687);
nand U3273 (N_3273,N_2996,N_2679);
nor U3274 (N_3274,N_2649,N_2672);
xnor U3275 (N_3275,N_2966,N_2923);
nand U3276 (N_3276,N_2740,N_2968);
nor U3277 (N_3277,N_2585,N_2732);
nor U3278 (N_3278,N_2911,N_2732);
or U3279 (N_3279,N_2645,N_2810);
xnor U3280 (N_3280,N_2867,N_2558);
or U3281 (N_3281,N_2853,N_2627);
xor U3282 (N_3282,N_2882,N_2774);
or U3283 (N_3283,N_2586,N_2760);
nor U3284 (N_3284,N_2922,N_2845);
nor U3285 (N_3285,N_2976,N_2915);
xor U3286 (N_3286,N_2775,N_2605);
xnor U3287 (N_3287,N_2571,N_2934);
or U3288 (N_3288,N_2749,N_2826);
and U3289 (N_3289,N_2726,N_2647);
nand U3290 (N_3290,N_2748,N_2636);
or U3291 (N_3291,N_2703,N_2986);
and U3292 (N_3292,N_2576,N_2791);
xnor U3293 (N_3293,N_2933,N_2592);
nand U3294 (N_3294,N_2849,N_2510);
xnor U3295 (N_3295,N_2633,N_2648);
xnor U3296 (N_3296,N_2717,N_2639);
xnor U3297 (N_3297,N_2911,N_2738);
nor U3298 (N_3298,N_2877,N_2737);
and U3299 (N_3299,N_2517,N_2850);
nand U3300 (N_3300,N_2524,N_2918);
nor U3301 (N_3301,N_2643,N_2848);
nand U3302 (N_3302,N_2910,N_2695);
and U3303 (N_3303,N_2936,N_2941);
nand U3304 (N_3304,N_2624,N_2659);
nor U3305 (N_3305,N_2677,N_2996);
nor U3306 (N_3306,N_2590,N_2515);
xor U3307 (N_3307,N_2561,N_2951);
xnor U3308 (N_3308,N_2827,N_2672);
or U3309 (N_3309,N_2951,N_2835);
nand U3310 (N_3310,N_2804,N_2525);
nor U3311 (N_3311,N_2577,N_2710);
xor U3312 (N_3312,N_2978,N_2660);
or U3313 (N_3313,N_2909,N_2762);
nand U3314 (N_3314,N_2602,N_2540);
or U3315 (N_3315,N_2800,N_2919);
and U3316 (N_3316,N_2947,N_2550);
nand U3317 (N_3317,N_2769,N_2662);
or U3318 (N_3318,N_2916,N_2544);
nand U3319 (N_3319,N_2721,N_2827);
nor U3320 (N_3320,N_2797,N_2602);
nor U3321 (N_3321,N_2888,N_2725);
or U3322 (N_3322,N_2905,N_2568);
nor U3323 (N_3323,N_2604,N_2700);
and U3324 (N_3324,N_2515,N_2736);
and U3325 (N_3325,N_2778,N_2690);
nor U3326 (N_3326,N_2910,N_2735);
and U3327 (N_3327,N_2971,N_2741);
and U3328 (N_3328,N_2973,N_2592);
nor U3329 (N_3329,N_2714,N_2929);
nand U3330 (N_3330,N_2918,N_2737);
or U3331 (N_3331,N_2576,N_2525);
or U3332 (N_3332,N_2774,N_2786);
xnor U3333 (N_3333,N_2630,N_2894);
or U3334 (N_3334,N_2615,N_2997);
and U3335 (N_3335,N_2541,N_2875);
or U3336 (N_3336,N_2996,N_2514);
nand U3337 (N_3337,N_2598,N_2839);
nand U3338 (N_3338,N_2847,N_2899);
or U3339 (N_3339,N_2912,N_2856);
nor U3340 (N_3340,N_2501,N_2720);
nand U3341 (N_3341,N_2924,N_2647);
and U3342 (N_3342,N_2639,N_2525);
nor U3343 (N_3343,N_2770,N_2718);
or U3344 (N_3344,N_2701,N_2549);
or U3345 (N_3345,N_2632,N_2637);
nor U3346 (N_3346,N_2890,N_2856);
xor U3347 (N_3347,N_2743,N_2969);
or U3348 (N_3348,N_2754,N_2779);
or U3349 (N_3349,N_2670,N_2641);
or U3350 (N_3350,N_2847,N_2859);
xnor U3351 (N_3351,N_2586,N_2777);
nor U3352 (N_3352,N_2739,N_2816);
and U3353 (N_3353,N_2603,N_2913);
and U3354 (N_3354,N_2548,N_2738);
and U3355 (N_3355,N_2839,N_2818);
nand U3356 (N_3356,N_2563,N_2671);
or U3357 (N_3357,N_2823,N_2770);
xor U3358 (N_3358,N_2791,N_2674);
xor U3359 (N_3359,N_2622,N_2578);
and U3360 (N_3360,N_2882,N_2513);
and U3361 (N_3361,N_2948,N_2989);
and U3362 (N_3362,N_2551,N_2711);
or U3363 (N_3363,N_2509,N_2730);
nand U3364 (N_3364,N_2663,N_2952);
xor U3365 (N_3365,N_2999,N_2897);
nor U3366 (N_3366,N_2619,N_2521);
nor U3367 (N_3367,N_2988,N_2516);
and U3368 (N_3368,N_2713,N_2896);
xor U3369 (N_3369,N_2755,N_2820);
xnor U3370 (N_3370,N_2626,N_2976);
xor U3371 (N_3371,N_2779,N_2955);
or U3372 (N_3372,N_2968,N_2759);
and U3373 (N_3373,N_2849,N_2526);
xor U3374 (N_3374,N_2658,N_2709);
xor U3375 (N_3375,N_2841,N_2863);
nand U3376 (N_3376,N_2747,N_2548);
nand U3377 (N_3377,N_2993,N_2876);
or U3378 (N_3378,N_2947,N_2539);
or U3379 (N_3379,N_2531,N_2789);
xnor U3380 (N_3380,N_2750,N_2860);
xnor U3381 (N_3381,N_2603,N_2543);
xor U3382 (N_3382,N_2530,N_2820);
and U3383 (N_3383,N_2671,N_2642);
xnor U3384 (N_3384,N_2845,N_2826);
nand U3385 (N_3385,N_2962,N_2822);
nand U3386 (N_3386,N_2617,N_2565);
or U3387 (N_3387,N_2547,N_2533);
or U3388 (N_3388,N_2649,N_2668);
and U3389 (N_3389,N_2579,N_2777);
nand U3390 (N_3390,N_2885,N_2897);
xor U3391 (N_3391,N_2994,N_2530);
nand U3392 (N_3392,N_2923,N_2874);
or U3393 (N_3393,N_2731,N_2733);
nand U3394 (N_3394,N_2724,N_2766);
xnor U3395 (N_3395,N_2520,N_2626);
or U3396 (N_3396,N_2979,N_2865);
nor U3397 (N_3397,N_2823,N_2666);
or U3398 (N_3398,N_2549,N_2752);
or U3399 (N_3399,N_2983,N_2595);
xnor U3400 (N_3400,N_2662,N_2712);
nor U3401 (N_3401,N_2870,N_2822);
xnor U3402 (N_3402,N_2586,N_2689);
xnor U3403 (N_3403,N_2916,N_2507);
nor U3404 (N_3404,N_2631,N_2675);
or U3405 (N_3405,N_2794,N_2688);
xor U3406 (N_3406,N_2959,N_2778);
xor U3407 (N_3407,N_2891,N_2543);
nor U3408 (N_3408,N_2844,N_2854);
nand U3409 (N_3409,N_2595,N_2658);
nor U3410 (N_3410,N_2952,N_2800);
or U3411 (N_3411,N_2853,N_2852);
nand U3412 (N_3412,N_2604,N_2971);
nand U3413 (N_3413,N_2619,N_2860);
nand U3414 (N_3414,N_2827,N_2640);
nand U3415 (N_3415,N_2625,N_2905);
xnor U3416 (N_3416,N_2804,N_2545);
or U3417 (N_3417,N_2878,N_2832);
nand U3418 (N_3418,N_2802,N_2901);
and U3419 (N_3419,N_2526,N_2612);
or U3420 (N_3420,N_2783,N_2516);
nor U3421 (N_3421,N_2676,N_2735);
xnor U3422 (N_3422,N_2595,N_2744);
or U3423 (N_3423,N_2954,N_2811);
nand U3424 (N_3424,N_2671,N_2851);
nor U3425 (N_3425,N_2705,N_2937);
or U3426 (N_3426,N_2836,N_2919);
nor U3427 (N_3427,N_2868,N_2698);
nand U3428 (N_3428,N_2802,N_2510);
and U3429 (N_3429,N_2779,N_2821);
xor U3430 (N_3430,N_2620,N_2944);
or U3431 (N_3431,N_2502,N_2537);
nand U3432 (N_3432,N_2665,N_2734);
or U3433 (N_3433,N_2982,N_2969);
and U3434 (N_3434,N_2784,N_2965);
nor U3435 (N_3435,N_2664,N_2884);
xnor U3436 (N_3436,N_2942,N_2788);
and U3437 (N_3437,N_2764,N_2596);
nand U3438 (N_3438,N_2664,N_2829);
and U3439 (N_3439,N_2613,N_2746);
nand U3440 (N_3440,N_2660,N_2949);
nor U3441 (N_3441,N_2680,N_2542);
nand U3442 (N_3442,N_2830,N_2565);
xnor U3443 (N_3443,N_2540,N_2950);
nand U3444 (N_3444,N_2630,N_2539);
or U3445 (N_3445,N_2607,N_2902);
or U3446 (N_3446,N_2559,N_2553);
xnor U3447 (N_3447,N_2810,N_2997);
xnor U3448 (N_3448,N_2763,N_2724);
nand U3449 (N_3449,N_2822,N_2565);
xnor U3450 (N_3450,N_2875,N_2672);
nor U3451 (N_3451,N_2916,N_2747);
nor U3452 (N_3452,N_2726,N_2739);
nor U3453 (N_3453,N_2690,N_2603);
xor U3454 (N_3454,N_2577,N_2597);
xor U3455 (N_3455,N_2968,N_2702);
and U3456 (N_3456,N_2639,N_2612);
nand U3457 (N_3457,N_2715,N_2871);
and U3458 (N_3458,N_2704,N_2680);
nand U3459 (N_3459,N_2604,N_2958);
or U3460 (N_3460,N_2708,N_2795);
xnor U3461 (N_3461,N_2547,N_2910);
or U3462 (N_3462,N_2576,N_2786);
xnor U3463 (N_3463,N_2762,N_2514);
or U3464 (N_3464,N_2974,N_2840);
or U3465 (N_3465,N_2823,N_2568);
nor U3466 (N_3466,N_2946,N_2702);
nand U3467 (N_3467,N_2696,N_2739);
xnor U3468 (N_3468,N_2643,N_2908);
xor U3469 (N_3469,N_2859,N_2580);
nand U3470 (N_3470,N_2822,N_2685);
or U3471 (N_3471,N_2661,N_2986);
nand U3472 (N_3472,N_2511,N_2556);
nand U3473 (N_3473,N_2734,N_2746);
xnor U3474 (N_3474,N_2905,N_2633);
nand U3475 (N_3475,N_2730,N_2511);
xnor U3476 (N_3476,N_2892,N_2929);
nand U3477 (N_3477,N_2771,N_2983);
xor U3478 (N_3478,N_2895,N_2914);
xor U3479 (N_3479,N_2734,N_2975);
nand U3480 (N_3480,N_2880,N_2962);
nor U3481 (N_3481,N_2760,N_2996);
and U3482 (N_3482,N_2849,N_2592);
xor U3483 (N_3483,N_2526,N_2952);
nand U3484 (N_3484,N_2634,N_2766);
nand U3485 (N_3485,N_2559,N_2584);
and U3486 (N_3486,N_2835,N_2552);
and U3487 (N_3487,N_2955,N_2823);
nand U3488 (N_3488,N_2676,N_2941);
and U3489 (N_3489,N_2551,N_2813);
nor U3490 (N_3490,N_2549,N_2793);
or U3491 (N_3491,N_2878,N_2646);
and U3492 (N_3492,N_2637,N_2514);
xnor U3493 (N_3493,N_2915,N_2535);
and U3494 (N_3494,N_2693,N_2964);
and U3495 (N_3495,N_2719,N_2986);
nand U3496 (N_3496,N_2655,N_2621);
nor U3497 (N_3497,N_2957,N_2697);
nand U3498 (N_3498,N_2909,N_2579);
xnor U3499 (N_3499,N_2542,N_2959);
nor U3500 (N_3500,N_3297,N_3283);
and U3501 (N_3501,N_3489,N_3309);
and U3502 (N_3502,N_3437,N_3161);
xnor U3503 (N_3503,N_3118,N_3075);
nand U3504 (N_3504,N_3197,N_3009);
or U3505 (N_3505,N_3200,N_3185);
or U3506 (N_3506,N_3040,N_3452);
nor U3507 (N_3507,N_3443,N_3416);
nand U3508 (N_3508,N_3227,N_3268);
or U3509 (N_3509,N_3417,N_3481);
nor U3510 (N_3510,N_3070,N_3491);
nor U3511 (N_3511,N_3105,N_3289);
or U3512 (N_3512,N_3005,N_3327);
xor U3513 (N_3513,N_3486,N_3001);
and U3514 (N_3514,N_3298,N_3037);
nand U3515 (N_3515,N_3494,N_3454);
or U3516 (N_3516,N_3103,N_3072);
or U3517 (N_3517,N_3435,N_3313);
nor U3518 (N_3518,N_3145,N_3134);
or U3519 (N_3519,N_3461,N_3484);
xnor U3520 (N_3520,N_3176,N_3074);
and U3521 (N_3521,N_3191,N_3036);
and U3522 (N_3522,N_3476,N_3352);
and U3523 (N_3523,N_3066,N_3394);
nand U3524 (N_3524,N_3446,N_3162);
nand U3525 (N_3525,N_3468,N_3333);
or U3526 (N_3526,N_3159,N_3376);
and U3527 (N_3527,N_3223,N_3255);
nor U3528 (N_3528,N_3382,N_3234);
nor U3529 (N_3529,N_3131,N_3373);
nor U3530 (N_3530,N_3083,N_3323);
xor U3531 (N_3531,N_3369,N_3477);
xnor U3532 (N_3532,N_3100,N_3206);
nor U3533 (N_3533,N_3194,N_3364);
nand U3534 (N_3534,N_3222,N_3095);
nor U3535 (N_3535,N_3168,N_3160);
xor U3536 (N_3536,N_3346,N_3294);
nor U3537 (N_3537,N_3123,N_3456);
or U3538 (N_3538,N_3071,N_3004);
and U3539 (N_3539,N_3126,N_3007);
nor U3540 (N_3540,N_3235,N_3102);
or U3541 (N_3541,N_3473,N_3339);
nand U3542 (N_3542,N_3342,N_3141);
xnor U3543 (N_3543,N_3124,N_3460);
nand U3544 (N_3544,N_3020,N_3090);
nand U3545 (N_3545,N_3219,N_3244);
nand U3546 (N_3546,N_3198,N_3390);
nor U3547 (N_3547,N_3371,N_3202);
nor U3548 (N_3548,N_3434,N_3326);
or U3549 (N_3549,N_3081,N_3467);
or U3550 (N_3550,N_3142,N_3015);
xnor U3551 (N_3551,N_3034,N_3117);
xor U3552 (N_3552,N_3455,N_3174);
nor U3553 (N_3553,N_3453,N_3366);
xor U3554 (N_3554,N_3210,N_3496);
and U3555 (N_3555,N_3096,N_3308);
xor U3556 (N_3556,N_3125,N_3431);
xor U3557 (N_3557,N_3304,N_3155);
and U3558 (N_3558,N_3393,N_3183);
or U3559 (N_3559,N_3248,N_3225);
and U3560 (N_3560,N_3285,N_3064);
and U3561 (N_3561,N_3139,N_3377);
nor U3562 (N_3562,N_3426,N_3493);
nand U3563 (N_3563,N_3316,N_3432);
or U3564 (N_3564,N_3166,N_3330);
nor U3565 (N_3565,N_3447,N_3212);
and U3566 (N_3566,N_3048,N_3173);
and U3567 (N_3567,N_3345,N_3024);
or U3568 (N_3568,N_3153,N_3088);
xnor U3569 (N_3569,N_3193,N_3119);
or U3570 (N_3570,N_3211,N_3314);
and U3571 (N_3571,N_3457,N_3281);
nand U3572 (N_3572,N_3082,N_3495);
nand U3573 (N_3573,N_3329,N_3472);
nand U3574 (N_3574,N_3488,N_3355);
nor U3575 (N_3575,N_3278,N_3325);
and U3576 (N_3576,N_3053,N_3092);
nor U3577 (N_3577,N_3152,N_3184);
or U3578 (N_3578,N_3063,N_3420);
nor U3579 (N_3579,N_3343,N_3470);
and U3580 (N_3580,N_3121,N_3334);
nand U3581 (N_3581,N_3052,N_3413);
nand U3582 (N_3582,N_3016,N_3143);
xnor U3583 (N_3583,N_3207,N_3291);
and U3584 (N_3584,N_3035,N_3350);
nand U3585 (N_3585,N_3190,N_3362);
and U3586 (N_3586,N_3384,N_3242);
nor U3587 (N_3587,N_3101,N_3490);
nand U3588 (N_3588,N_3012,N_3406);
xnor U3589 (N_3589,N_3295,N_3165);
or U3590 (N_3590,N_3111,N_3208);
xor U3591 (N_3591,N_3499,N_3412);
or U3592 (N_3592,N_3353,N_3232);
and U3593 (N_3593,N_3263,N_3360);
or U3594 (N_3594,N_3032,N_3010);
xor U3595 (N_3595,N_3337,N_3019);
xnor U3596 (N_3596,N_3429,N_3449);
xnor U3597 (N_3597,N_3370,N_3475);
or U3598 (N_3598,N_3149,N_3469);
nor U3599 (N_3599,N_3196,N_3240);
nand U3600 (N_3600,N_3167,N_3367);
xnor U3601 (N_3601,N_3182,N_3013);
and U3602 (N_3602,N_3324,N_3265);
or U3603 (N_3603,N_3471,N_3112);
nand U3604 (N_3604,N_3279,N_3109);
nor U3605 (N_3605,N_3135,N_3409);
nand U3606 (N_3606,N_3444,N_3419);
nand U3607 (N_3607,N_3215,N_3178);
and U3608 (N_3608,N_3114,N_3361);
and U3609 (N_3609,N_3132,N_3328);
or U3610 (N_3610,N_3104,N_3485);
xnor U3611 (N_3611,N_3459,N_3395);
xnor U3612 (N_3612,N_3249,N_3405);
nand U3613 (N_3613,N_3136,N_3230);
and U3614 (N_3614,N_3372,N_3347);
or U3615 (N_3615,N_3307,N_3106);
nor U3616 (N_3616,N_3008,N_3340);
xnor U3617 (N_3617,N_3170,N_3236);
nand U3618 (N_3618,N_3042,N_3478);
nand U3619 (N_3619,N_3127,N_3050);
nand U3620 (N_3620,N_3055,N_3389);
or U3621 (N_3621,N_3058,N_3256);
and U3622 (N_3622,N_3480,N_3401);
xor U3623 (N_3623,N_3262,N_3287);
and U3624 (N_3624,N_3217,N_3421);
xnor U3625 (N_3625,N_3116,N_3415);
xnor U3626 (N_3626,N_3445,N_3466);
xor U3627 (N_3627,N_3128,N_3451);
or U3628 (N_3628,N_3154,N_3302);
nor U3629 (N_3629,N_3483,N_3332);
and U3630 (N_3630,N_3220,N_3077);
and U3631 (N_3631,N_3296,N_3321);
and U3632 (N_3632,N_3006,N_3271);
xor U3633 (N_3633,N_3274,N_3425);
xnor U3634 (N_3634,N_3311,N_3423);
nor U3635 (N_3635,N_3356,N_3348);
nand U3636 (N_3636,N_3051,N_3046);
nor U3637 (N_3637,N_3336,N_3041);
xor U3638 (N_3638,N_3204,N_3043);
or U3639 (N_3639,N_3318,N_3427);
nand U3640 (N_3640,N_3438,N_3363);
nand U3641 (N_3641,N_3085,N_3442);
or U3642 (N_3642,N_3171,N_3031);
nand U3643 (N_3643,N_3086,N_3110);
and U3644 (N_3644,N_3186,N_3250);
xor U3645 (N_3645,N_3246,N_3293);
and U3646 (N_3646,N_3054,N_3224);
or U3647 (N_3647,N_3306,N_3441);
xor U3648 (N_3648,N_3270,N_3078);
nor U3649 (N_3649,N_3399,N_3463);
and U3650 (N_3650,N_3277,N_3322);
or U3651 (N_3651,N_3267,N_3238);
and U3652 (N_3652,N_3216,N_3241);
and U3653 (N_3653,N_3060,N_3286);
nand U3654 (N_3654,N_3418,N_3315);
nand U3655 (N_3655,N_3014,N_3331);
xor U3656 (N_3656,N_3381,N_3099);
and U3657 (N_3657,N_3002,N_3436);
and U3658 (N_3658,N_3253,N_3069);
xnor U3659 (N_3659,N_3156,N_3059);
nand U3660 (N_3660,N_3138,N_3402);
or U3661 (N_3661,N_3301,N_3079);
xnor U3662 (N_3662,N_3404,N_3122);
nand U3663 (N_3663,N_3067,N_3312);
nor U3664 (N_3664,N_3094,N_3179);
and U3665 (N_3665,N_3218,N_3027);
nor U3666 (N_3666,N_3057,N_3018);
or U3667 (N_3667,N_3247,N_3221);
or U3668 (N_3668,N_3113,N_3140);
nor U3669 (N_3669,N_3093,N_3084);
nand U3670 (N_3670,N_3497,N_3269);
nand U3671 (N_3671,N_3319,N_3407);
nor U3672 (N_3672,N_3341,N_3189);
or U3673 (N_3673,N_3017,N_3396);
nor U3674 (N_3674,N_3080,N_3158);
xor U3675 (N_3675,N_3275,N_3310);
and U3676 (N_3676,N_3282,N_3129);
nor U3677 (N_3677,N_3033,N_3264);
xor U3678 (N_3678,N_3428,N_3440);
nand U3679 (N_3679,N_3335,N_3172);
xnor U3680 (N_3680,N_3192,N_3414);
or U3681 (N_3681,N_3378,N_3025);
and U3682 (N_3682,N_3147,N_3028);
xnor U3683 (N_3683,N_3021,N_3379);
or U3684 (N_3684,N_3231,N_3030);
nand U3685 (N_3685,N_3261,N_3115);
nor U3686 (N_3686,N_3003,N_3365);
nor U3687 (N_3687,N_3357,N_3492);
nand U3688 (N_3688,N_3462,N_3380);
and U3689 (N_3689,N_3266,N_3000);
or U3690 (N_3690,N_3068,N_3400);
nand U3691 (N_3691,N_3257,N_3011);
or U3692 (N_3692,N_3398,N_3252);
nor U3693 (N_3693,N_3303,N_3273);
nor U3694 (N_3694,N_3087,N_3047);
nor U3695 (N_3695,N_3146,N_3214);
or U3696 (N_3696,N_3076,N_3203);
nand U3697 (N_3697,N_3272,N_3243);
or U3698 (N_3698,N_3107,N_3359);
xnor U3699 (N_3699,N_3169,N_3098);
nand U3700 (N_3700,N_3299,N_3305);
and U3701 (N_3701,N_3338,N_3411);
or U3702 (N_3702,N_3391,N_3387);
xnor U3703 (N_3703,N_3038,N_3392);
or U3704 (N_3704,N_3164,N_3022);
nor U3705 (N_3705,N_3430,N_3276);
nand U3706 (N_3706,N_3233,N_3280);
xnor U3707 (N_3707,N_3245,N_3199);
nor U3708 (N_3708,N_3150,N_3288);
and U3709 (N_3709,N_3151,N_3130);
nand U3710 (N_3710,N_3422,N_3201);
nor U3711 (N_3711,N_3259,N_3097);
nand U3712 (N_3712,N_3292,N_3195);
or U3713 (N_3713,N_3354,N_3408);
nor U3714 (N_3714,N_3385,N_3209);
nor U3715 (N_3715,N_3450,N_3175);
nor U3716 (N_3716,N_3045,N_3320);
xnor U3717 (N_3717,N_3482,N_3251);
nor U3718 (N_3718,N_3061,N_3375);
and U3719 (N_3719,N_3374,N_3237);
or U3720 (N_3720,N_3205,N_3023);
nand U3721 (N_3721,N_3073,N_3163);
nor U3722 (N_3722,N_3133,N_3029);
or U3723 (N_3723,N_3228,N_3187);
nor U3724 (N_3724,N_3464,N_3039);
xnor U3725 (N_3725,N_3226,N_3344);
or U3726 (N_3726,N_3383,N_3397);
or U3727 (N_3727,N_3108,N_3358);
and U3728 (N_3728,N_3410,N_3181);
nor U3729 (N_3729,N_3284,N_3089);
and U3730 (N_3730,N_3177,N_3424);
and U3731 (N_3731,N_3062,N_3300);
nor U3732 (N_3732,N_3465,N_3229);
or U3733 (N_3733,N_3188,N_3044);
and U3734 (N_3734,N_3479,N_3474);
or U3735 (N_3735,N_3388,N_3458);
nor U3736 (N_3736,N_3448,N_3351);
xnor U3737 (N_3737,N_3433,N_3258);
nor U3738 (N_3738,N_3239,N_3403);
nor U3739 (N_3739,N_3065,N_3260);
and U3740 (N_3740,N_3290,N_3213);
nand U3741 (N_3741,N_3120,N_3137);
nor U3742 (N_3742,N_3368,N_3439);
xor U3743 (N_3743,N_3317,N_3157);
nor U3744 (N_3744,N_3056,N_3026);
xnor U3745 (N_3745,N_3049,N_3349);
nand U3746 (N_3746,N_3144,N_3498);
nand U3747 (N_3747,N_3148,N_3180);
or U3748 (N_3748,N_3386,N_3487);
nor U3749 (N_3749,N_3091,N_3254);
nand U3750 (N_3750,N_3263,N_3102);
nor U3751 (N_3751,N_3269,N_3248);
xnor U3752 (N_3752,N_3123,N_3448);
and U3753 (N_3753,N_3127,N_3297);
nor U3754 (N_3754,N_3367,N_3297);
xor U3755 (N_3755,N_3228,N_3215);
nor U3756 (N_3756,N_3441,N_3071);
and U3757 (N_3757,N_3446,N_3004);
xnor U3758 (N_3758,N_3386,N_3255);
nor U3759 (N_3759,N_3178,N_3281);
nor U3760 (N_3760,N_3143,N_3167);
or U3761 (N_3761,N_3473,N_3272);
nor U3762 (N_3762,N_3463,N_3280);
or U3763 (N_3763,N_3242,N_3019);
nor U3764 (N_3764,N_3031,N_3246);
nand U3765 (N_3765,N_3339,N_3245);
and U3766 (N_3766,N_3109,N_3114);
and U3767 (N_3767,N_3351,N_3494);
and U3768 (N_3768,N_3117,N_3484);
xnor U3769 (N_3769,N_3211,N_3016);
or U3770 (N_3770,N_3303,N_3118);
and U3771 (N_3771,N_3288,N_3208);
nand U3772 (N_3772,N_3331,N_3199);
and U3773 (N_3773,N_3471,N_3350);
nand U3774 (N_3774,N_3340,N_3479);
nand U3775 (N_3775,N_3398,N_3312);
xor U3776 (N_3776,N_3377,N_3470);
xor U3777 (N_3777,N_3188,N_3107);
xor U3778 (N_3778,N_3125,N_3277);
and U3779 (N_3779,N_3076,N_3245);
nor U3780 (N_3780,N_3080,N_3462);
nand U3781 (N_3781,N_3067,N_3417);
and U3782 (N_3782,N_3054,N_3418);
and U3783 (N_3783,N_3346,N_3075);
or U3784 (N_3784,N_3152,N_3361);
or U3785 (N_3785,N_3191,N_3272);
nand U3786 (N_3786,N_3147,N_3053);
xor U3787 (N_3787,N_3114,N_3177);
nor U3788 (N_3788,N_3314,N_3173);
and U3789 (N_3789,N_3042,N_3065);
xor U3790 (N_3790,N_3283,N_3303);
nand U3791 (N_3791,N_3318,N_3363);
or U3792 (N_3792,N_3365,N_3403);
or U3793 (N_3793,N_3116,N_3108);
nor U3794 (N_3794,N_3263,N_3028);
xnor U3795 (N_3795,N_3051,N_3407);
nor U3796 (N_3796,N_3036,N_3487);
nand U3797 (N_3797,N_3469,N_3074);
and U3798 (N_3798,N_3021,N_3182);
nor U3799 (N_3799,N_3238,N_3446);
or U3800 (N_3800,N_3157,N_3427);
or U3801 (N_3801,N_3146,N_3077);
xor U3802 (N_3802,N_3031,N_3390);
and U3803 (N_3803,N_3295,N_3496);
xor U3804 (N_3804,N_3344,N_3062);
nand U3805 (N_3805,N_3146,N_3200);
or U3806 (N_3806,N_3491,N_3221);
and U3807 (N_3807,N_3410,N_3381);
or U3808 (N_3808,N_3282,N_3227);
xnor U3809 (N_3809,N_3374,N_3045);
or U3810 (N_3810,N_3287,N_3306);
nand U3811 (N_3811,N_3354,N_3431);
nor U3812 (N_3812,N_3043,N_3409);
and U3813 (N_3813,N_3223,N_3098);
or U3814 (N_3814,N_3328,N_3489);
nand U3815 (N_3815,N_3074,N_3044);
or U3816 (N_3816,N_3157,N_3221);
nand U3817 (N_3817,N_3471,N_3068);
or U3818 (N_3818,N_3394,N_3271);
or U3819 (N_3819,N_3078,N_3241);
or U3820 (N_3820,N_3110,N_3129);
nor U3821 (N_3821,N_3211,N_3067);
or U3822 (N_3822,N_3146,N_3073);
nor U3823 (N_3823,N_3170,N_3496);
or U3824 (N_3824,N_3205,N_3333);
or U3825 (N_3825,N_3464,N_3251);
or U3826 (N_3826,N_3394,N_3023);
nand U3827 (N_3827,N_3298,N_3244);
or U3828 (N_3828,N_3223,N_3014);
xnor U3829 (N_3829,N_3210,N_3408);
or U3830 (N_3830,N_3495,N_3452);
and U3831 (N_3831,N_3385,N_3448);
xor U3832 (N_3832,N_3136,N_3130);
nand U3833 (N_3833,N_3305,N_3282);
or U3834 (N_3834,N_3227,N_3358);
or U3835 (N_3835,N_3172,N_3011);
xor U3836 (N_3836,N_3404,N_3322);
nor U3837 (N_3837,N_3085,N_3268);
nor U3838 (N_3838,N_3162,N_3277);
and U3839 (N_3839,N_3146,N_3403);
nor U3840 (N_3840,N_3140,N_3498);
xor U3841 (N_3841,N_3274,N_3101);
nor U3842 (N_3842,N_3169,N_3192);
xnor U3843 (N_3843,N_3207,N_3404);
nor U3844 (N_3844,N_3269,N_3481);
or U3845 (N_3845,N_3246,N_3140);
nor U3846 (N_3846,N_3068,N_3409);
xnor U3847 (N_3847,N_3196,N_3471);
and U3848 (N_3848,N_3459,N_3212);
nand U3849 (N_3849,N_3476,N_3362);
and U3850 (N_3850,N_3131,N_3101);
and U3851 (N_3851,N_3238,N_3179);
or U3852 (N_3852,N_3068,N_3075);
or U3853 (N_3853,N_3135,N_3279);
or U3854 (N_3854,N_3147,N_3272);
or U3855 (N_3855,N_3197,N_3005);
and U3856 (N_3856,N_3293,N_3055);
or U3857 (N_3857,N_3491,N_3342);
or U3858 (N_3858,N_3090,N_3255);
xnor U3859 (N_3859,N_3371,N_3415);
nor U3860 (N_3860,N_3430,N_3303);
nor U3861 (N_3861,N_3090,N_3342);
nor U3862 (N_3862,N_3184,N_3146);
or U3863 (N_3863,N_3341,N_3014);
xnor U3864 (N_3864,N_3003,N_3088);
and U3865 (N_3865,N_3381,N_3032);
or U3866 (N_3866,N_3100,N_3457);
or U3867 (N_3867,N_3139,N_3254);
nand U3868 (N_3868,N_3153,N_3481);
nand U3869 (N_3869,N_3270,N_3286);
nor U3870 (N_3870,N_3018,N_3206);
nor U3871 (N_3871,N_3009,N_3288);
xnor U3872 (N_3872,N_3325,N_3405);
nor U3873 (N_3873,N_3097,N_3061);
nor U3874 (N_3874,N_3106,N_3271);
nor U3875 (N_3875,N_3336,N_3391);
and U3876 (N_3876,N_3492,N_3254);
and U3877 (N_3877,N_3351,N_3110);
nand U3878 (N_3878,N_3313,N_3311);
and U3879 (N_3879,N_3097,N_3225);
xnor U3880 (N_3880,N_3100,N_3111);
nor U3881 (N_3881,N_3468,N_3126);
and U3882 (N_3882,N_3080,N_3320);
or U3883 (N_3883,N_3339,N_3048);
nor U3884 (N_3884,N_3251,N_3024);
nor U3885 (N_3885,N_3020,N_3143);
xor U3886 (N_3886,N_3110,N_3032);
or U3887 (N_3887,N_3268,N_3396);
nand U3888 (N_3888,N_3447,N_3073);
xnor U3889 (N_3889,N_3123,N_3435);
or U3890 (N_3890,N_3366,N_3450);
and U3891 (N_3891,N_3373,N_3064);
and U3892 (N_3892,N_3234,N_3227);
or U3893 (N_3893,N_3318,N_3230);
xor U3894 (N_3894,N_3136,N_3064);
xor U3895 (N_3895,N_3401,N_3082);
nand U3896 (N_3896,N_3400,N_3293);
or U3897 (N_3897,N_3102,N_3462);
and U3898 (N_3898,N_3367,N_3332);
nand U3899 (N_3899,N_3129,N_3017);
nand U3900 (N_3900,N_3166,N_3404);
nor U3901 (N_3901,N_3001,N_3442);
and U3902 (N_3902,N_3109,N_3250);
and U3903 (N_3903,N_3040,N_3030);
nor U3904 (N_3904,N_3028,N_3347);
nand U3905 (N_3905,N_3157,N_3393);
nor U3906 (N_3906,N_3468,N_3263);
nand U3907 (N_3907,N_3393,N_3402);
nor U3908 (N_3908,N_3452,N_3256);
or U3909 (N_3909,N_3193,N_3194);
nor U3910 (N_3910,N_3328,N_3338);
and U3911 (N_3911,N_3233,N_3176);
xor U3912 (N_3912,N_3088,N_3360);
xor U3913 (N_3913,N_3394,N_3337);
nor U3914 (N_3914,N_3498,N_3198);
or U3915 (N_3915,N_3176,N_3054);
xor U3916 (N_3916,N_3381,N_3175);
and U3917 (N_3917,N_3382,N_3057);
nor U3918 (N_3918,N_3347,N_3393);
nor U3919 (N_3919,N_3430,N_3337);
nor U3920 (N_3920,N_3160,N_3180);
nor U3921 (N_3921,N_3242,N_3317);
xnor U3922 (N_3922,N_3107,N_3117);
nand U3923 (N_3923,N_3142,N_3382);
and U3924 (N_3924,N_3160,N_3120);
nand U3925 (N_3925,N_3174,N_3075);
nand U3926 (N_3926,N_3136,N_3094);
or U3927 (N_3927,N_3440,N_3350);
nand U3928 (N_3928,N_3295,N_3101);
xnor U3929 (N_3929,N_3226,N_3463);
nand U3930 (N_3930,N_3266,N_3075);
xor U3931 (N_3931,N_3339,N_3301);
nor U3932 (N_3932,N_3128,N_3483);
nand U3933 (N_3933,N_3343,N_3324);
nor U3934 (N_3934,N_3403,N_3199);
nand U3935 (N_3935,N_3043,N_3116);
nor U3936 (N_3936,N_3202,N_3249);
or U3937 (N_3937,N_3479,N_3112);
nand U3938 (N_3938,N_3220,N_3483);
nor U3939 (N_3939,N_3062,N_3044);
nor U3940 (N_3940,N_3185,N_3391);
or U3941 (N_3941,N_3085,N_3080);
or U3942 (N_3942,N_3013,N_3472);
and U3943 (N_3943,N_3221,N_3301);
or U3944 (N_3944,N_3438,N_3334);
and U3945 (N_3945,N_3304,N_3024);
xnor U3946 (N_3946,N_3322,N_3315);
or U3947 (N_3947,N_3339,N_3246);
or U3948 (N_3948,N_3144,N_3092);
or U3949 (N_3949,N_3183,N_3332);
and U3950 (N_3950,N_3365,N_3148);
or U3951 (N_3951,N_3040,N_3331);
and U3952 (N_3952,N_3408,N_3273);
and U3953 (N_3953,N_3231,N_3223);
nor U3954 (N_3954,N_3322,N_3445);
xnor U3955 (N_3955,N_3487,N_3309);
xor U3956 (N_3956,N_3480,N_3315);
nor U3957 (N_3957,N_3051,N_3394);
and U3958 (N_3958,N_3143,N_3390);
nand U3959 (N_3959,N_3243,N_3138);
nand U3960 (N_3960,N_3021,N_3197);
and U3961 (N_3961,N_3326,N_3365);
nor U3962 (N_3962,N_3040,N_3202);
nand U3963 (N_3963,N_3211,N_3104);
nor U3964 (N_3964,N_3154,N_3265);
nand U3965 (N_3965,N_3306,N_3362);
and U3966 (N_3966,N_3305,N_3120);
nand U3967 (N_3967,N_3055,N_3274);
or U3968 (N_3968,N_3472,N_3321);
and U3969 (N_3969,N_3168,N_3232);
and U3970 (N_3970,N_3309,N_3285);
nor U3971 (N_3971,N_3104,N_3433);
nand U3972 (N_3972,N_3123,N_3296);
and U3973 (N_3973,N_3129,N_3332);
nor U3974 (N_3974,N_3320,N_3156);
nor U3975 (N_3975,N_3007,N_3275);
xnor U3976 (N_3976,N_3138,N_3489);
nor U3977 (N_3977,N_3017,N_3487);
or U3978 (N_3978,N_3026,N_3498);
xnor U3979 (N_3979,N_3048,N_3486);
nand U3980 (N_3980,N_3279,N_3219);
nand U3981 (N_3981,N_3482,N_3197);
and U3982 (N_3982,N_3230,N_3465);
nand U3983 (N_3983,N_3179,N_3125);
or U3984 (N_3984,N_3213,N_3149);
and U3985 (N_3985,N_3138,N_3210);
and U3986 (N_3986,N_3144,N_3392);
xor U3987 (N_3987,N_3386,N_3154);
xnor U3988 (N_3988,N_3010,N_3066);
or U3989 (N_3989,N_3159,N_3210);
nor U3990 (N_3990,N_3093,N_3255);
xnor U3991 (N_3991,N_3228,N_3051);
and U3992 (N_3992,N_3018,N_3377);
or U3993 (N_3993,N_3415,N_3127);
nor U3994 (N_3994,N_3115,N_3370);
xnor U3995 (N_3995,N_3440,N_3491);
xor U3996 (N_3996,N_3089,N_3288);
and U3997 (N_3997,N_3165,N_3252);
or U3998 (N_3998,N_3319,N_3028);
nor U3999 (N_3999,N_3353,N_3409);
and U4000 (N_4000,N_3544,N_3842);
nor U4001 (N_4001,N_3634,N_3723);
nand U4002 (N_4002,N_3504,N_3779);
and U4003 (N_4003,N_3730,N_3569);
nor U4004 (N_4004,N_3680,N_3515);
or U4005 (N_4005,N_3759,N_3951);
xor U4006 (N_4006,N_3732,N_3564);
nand U4007 (N_4007,N_3839,N_3667);
nor U4008 (N_4008,N_3882,N_3994);
nand U4009 (N_4009,N_3674,N_3586);
or U4010 (N_4010,N_3860,N_3834);
or U4011 (N_4011,N_3760,N_3969);
and U4012 (N_4012,N_3602,N_3992);
and U4013 (N_4013,N_3867,N_3506);
nand U4014 (N_4014,N_3687,N_3814);
nand U4015 (N_4015,N_3733,N_3510);
nor U4016 (N_4016,N_3875,N_3995);
or U4017 (N_4017,N_3750,N_3600);
nor U4018 (N_4018,N_3530,N_3826);
nand U4019 (N_4019,N_3933,N_3686);
and U4020 (N_4020,N_3974,N_3986);
or U4021 (N_4021,N_3924,N_3631);
nand U4022 (N_4022,N_3589,N_3554);
nand U4023 (N_4023,N_3528,N_3784);
xor U4024 (N_4024,N_3726,N_3583);
xnor U4025 (N_4025,N_3688,N_3908);
nand U4026 (N_4026,N_3755,N_3537);
or U4027 (N_4027,N_3563,N_3907);
and U4028 (N_4028,N_3889,N_3597);
nor U4029 (N_4029,N_3659,N_3695);
nand U4030 (N_4030,N_3997,N_3522);
and U4031 (N_4031,N_3518,N_3640);
or U4032 (N_4032,N_3658,N_3941);
and U4033 (N_4033,N_3541,N_3558);
nand U4034 (N_4034,N_3998,N_3523);
or U4035 (N_4035,N_3970,N_3845);
and U4036 (N_4036,N_3502,N_3877);
nand U4037 (N_4037,N_3521,N_3802);
or U4038 (N_4038,N_3722,N_3618);
nor U4039 (N_4039,N_3513,N_3989);
xor U4040 (N_4040,N_3773,N_3632);
nand U4041 (N_4041,N_3570,N_3592);
nor U4042 (N_4042,N_3936,N_3988);
nand U4043 (N_4043,N_3792,N_3711);
nand U4044 (N_4044,N_3847,N_3712);
or U4045 (N_4045,N_3525,N_3800);
nor U4046 (N_4046,N_3973,N_3991);
xor U4047 (N_4047,N_3543,N_3761);
and U4048 (N_4048,N_3756,N_3971);
nand U4049 (N_4049,N_3946,N_3888);
and U4050 (N_4050,N_3682,N_3966);
or U4051 (N_4051,N_3607,N_3580);
and U4052 (N_4052,N_3938,N_3813);
and U4053 (N_4053,N_3823,N_3816);
xor U4054 (N_4054,N_3654,N_3780);
and U4055 (N_4055,N_3928,N_3944);
xor U4056 (N_4056,N_3857,N_3613);
nand U4057 (N_4057,N_3996,N_3771);
nand U4058 (N_4058,N_3782,N_3850);
xnor U4059 (N_4059,N_3657,N_3736);
nand U4060 (N_4060,N_3767,N_3638);
xor U4061 (N_4061,N_3603,N_3836);
nor U4062 (N_4062,N_3651,N_3702);
and U4063 (N_4063,N_3934,N_3808);
or U4064 (N_4064,N_3681,N_3775);
nand U4065 (N_4065,N_3999,N_3669);
or U4066 (N_4066,N_3844,N_3552);
and U4067 (N_4067,N_3633,N_3748);
or U4068 (N_4068,N_3747,N_3980);
nand U4069 (N_4069,N_3822,N_3833);
nand U4070 (N_4070,N_3962,N_3954);
nor U4071 (N_4071,N_3741,N_3567);
or U4072 (N_4072,N_3656,N_3621);
xnor U4073 (N_4073,N_3508,N_3745);
or U4074 (N_4074,N_3935,N_3894);
xor U4075 (N_4075,N_3627,N_3519);
or U4076 (N_4076,N_3864,N_3720);
nand U4077 (N_4077,N_3619,N_3719);
or U4078 (N_4078,N_3555,N_3550);
nor U4079 (N_4079,N_3809,N_3795);
nor U4080 (N_4080,N_3866,N_3620);
or U4081 (N_4081,N_3704,N_3899);
or U4082 (N_4082,N_3628,N_3914);
xnor U4083 (N_4083,N_3653,N_3781);
and U4084 (N_4084,N_3961,N_3650);
nand U4085 (N_4085,N_3874,N_3769);
xnor U4086 (N_4086,N_3548,N_3922);
xnor U4087 (N_4087,N_3953,N_3965);
nor U4088 (N_4088,N_3824,N_3786);
or U4089 (N_4089,N_3500,N_3666);
and U4090 (N_4090,N_3531,N_3787);
and U4091 (N_4091,N_3957,N_3766);
nor U4092 (N_4092,N_3673,N_3642);
and U4093 (N_4093,N_3643,N_3940);
nor U4094 (N_4094,N_3532,N_3731);
or U4095 (N_4095,N_3807,N_3849);
or U4096 (N_4096,N_3566,N_3876);
nor U4097 (N_4097,N_3887,N_3920);
or U4098 (N_4098,N_3827,N_3828);
or U4099 (N_4099,N_3945,N_3838);
nand U4100 (N_4100,N_3739,N_3599);
and U4101 (N_4101,N_3605,N_3872);
or U4102 (N_4102,N_3978,N_3890);
or U4103 (N_4103,N_3705,N_3676);
xnor U4104 (N_4104,N_3573,N_3757);
nor U4105 (N_4105,N_3709,N_3830);
nand U4106 (N_4106,N_3865,N_3959);
xnor U4107 (N_4107,N_3539,N_3509);
or U4108 (N_4108,N_3810,N_3851);
nand U4109 (N_4109,N_3511,N_3536);
xor U4110 (N_4110,N_3843,N_3790);
or U4111 (N_4111,N_3579,N_3852);
and U4112 (N_4112,N_3683,N_3987);
and U4113 (N_4113,N_3776,N_3762);
xnor U4114 (N_4114,N_3937,N_3801);
nand U4115 (N_4115,N_3979,N_3854);
and U4116 (N_4116,N_3902,N_3685);
or U4117 (N_4117,N_3553,N_3734);
nand U4118 (N_4118,N_3785,N_3846);
nor U4119 (N_4119,N_3529,N_3533);
xor U4120 (N_4120,N_3968,N_3811);
and U4121 (N_4121,N_3738,N_3770);
nor U4122 (N_4122,N_3869,N_3626);
nand U4123 (N_4123,N_3881,N_3871);
and U4124 (N_4124,N_3630,N_3975);
nor U4125 (N_4125,N_3942,N_3926);
xnor U4126 (N_4126,N_3715,N_3601);
and U4127 (N_4127,N_3527,N_3943);
or U4128 (N_4128,N_3691,N_3963);
nor U4129 (N_4129,N_3636,N_3909);
nand U4130 (N_4130,N_3831,N_3868);
or U4131 (N_4131,N_3571,N_3708);
nand U4132 (N_4132,N_3557,N_3742);
or U4133 (N_4133,N_3644,N_3598);
and U4134 (N_4134,N_3516,N_3675);
nand U4135 (N_4135,N_3964,N_3724);
nor U4136 (N_4136,N_3829,N_3665);
nand U4137 (N_4137,N_3624,N_3743);
nand U4138 (N_4138,N_3900,N_3614);
nor U4139 (N_4139,N_3870,N_3660);
and U4140 (N_4140,N_3594,N_3616);
and U4141 (N_4141,N_3604,N_3668);
nand U4142 (N_4142,N_3958,N_3955);
and U4143 (N_4143,N_3905,N_3950);
and U4144 (N_4144,N_3803,N_3841);
nand U4145 (N_4145,N_3568,N_3983);
and U4146 (N_4146,N_3639,N_3910);
nand U4147 (N_4147,N_3575,N_3777);
and U4148 (N_4148,N_3679,N_3812);
xnor U4149 (N_4149,N_3820,N_3556);
or U4150 (N_4150,N_3699,N_3728);
or U4151 (N_4151,N_3538,N_3512);
or U4152 (N_4152,N_3805,N_3751);
nand U4153 (N_4153,N_3577,N_3898);
nand U4154 (N_4154,N_3774,N_3815);
nor U4155 (N_4155,N_3821,N_3949);
or U4156 (N_4156,N_3609,N_3591);
xor U4157 (N_4157,N_3918,N_3892);
or U4158 (N_4158,N_3697,N_3896);
nor U4159 (N_4159,N_3520,N_3694);
or U4160 (N_4160,N_3749,N_3939);
and U4161 (N_4161,N_3878,N_3646);
nand U4162 (N_4162,N_3572,N_3648);
nor U4163 (N_4163,N_3585,N_3982);
and U4164 (N_4164,N_3678,N_3819);
or U4165 (N_4165,N_3588,N_3990);
or U4166 (N_4166,N_3562,N_3976);
or U4167 (N_4167,N_3623,N_3696);
or U4168 (N_4168,N_3617,N_3647);
or U4169 (N_4169,N_3606,N_3740);
and U4170 (N_4170,N_3885,N_3891);
xor U4171 (N_4171,N_3789,N_3690);
xnor U4172 (N_4172,N_3880,N_3952);
nand U4173 (N_4173,N_3545,N_3977);
and U4174 (N_4174,N_3535,N_3858);
nand U4175 (N_4175,N_3684,N_3758);
and U4176 (N_4176,N_3707,N_3817);
nand U4177 (N_4177,N_3848,N_3931);
nand U4178 (N_4178,N_3596,N_3714);
and U4179 (N_4179,N_3993,N_3517);
xor U4180 (N_4180,N_3559,N_3972);
nor U4181 (N_4181,N_3663,N_3825);
and U4182 (N_4182,N_3895,N_3547);
or U4183 (N_4183,N_3718,N_3855);
nor U4184 (N_4184,N_3911,N_3625);
xor U4185 (N_4185,N_3540,N_3706);
or U4186 (N_4186,N_3692,N_3655);
nor U4187 (N_4187,N_3716,N_3611);
nand U4188 (N_4188,N_3754,N_3729);
nand U4189 (N_4189,N_3664,N_3542);
nand U4190 (N_4190,N_3797,N_3689);
nand U4191 (N_4191,N_3915,N_3565);
and U4192 (N_4192,N_3985,N_3590);
or U4193 (N_4193,N_3727,N_3710);
and U4194 (N_4194,N_3641,N_3917);
nor U4195 (N_4195,N_3788,N_3549);
or U4196 (N_4196,N_3859,N_3622);
and U4197 (N_4197,N_3765,N_3514);
or U4198 (N_4198,N_3507,N_3981);
xor U4199 (N_4199,N_3832,N_3735);
nand U4200 (N_4200,N_3561,N_3753);
nor U4201 (N_4201,N_3574,N_3906);
or U4202 (N_4202,N_3778,N_3593);
xnor U4203 (N_4203,N_3582,N_3652);
or U4204 (N_4204,N_3903,N_3879);
nand U4205 (N_4205,N_3921,N_3923);
nand U4206 (N_4206,N_3635,N_3752);
and U4207 (N_4207,N_3534,N_3893);
and U4208 (N_4208,N_3798,N_3956);
or U4209 (N_4209,N_3737,N_3744);
or U4210 (N_4210,N_3862,N_3560);
or U4211 (N_4211,N_3932,N_3856);
nand U4212 (N_4212,N_3904,N_3698);
or U4213 (N_4213,N_3581,N_3693);
nor U4214 (N_4214,N_3818,N_3610);
xor U4215 (N_4215,N_3806,N_3840);
xor U4216 (N_4216,N_3746,N_3677);
or U4217 (N_4217,N_3883,N_3612);
xnor U4218 (N_4218,N_3967,N_3662);
xnor U4219 (N_4219,N_3948,N_3764);
nand U4220 (N_4220,N_3637,N_3873);
nand U4221 (N_4221,N_3670,N_3629);
xnor U4222 (N_4222,N_3721,N_3947);
nor U4223 (N_4223,N_3700,N_3595);
or U4224 (N_4224,N_3701,N_3526);
and U4225 (N_4225,N_3863,N_3927);
nor U4226 (N_4226,N_3799,N_3661);
xor U4227 (N_4227,N_3703,N_3837);
and U4228 (N_4228,N_3960,N_3768);
nor U4229 (N_4229,N_3649,N_3717);
nor U4230 (N_4230,N_3804,N_3913);
xor U4231 (N_4231,N_3587,N_3793);
or U4232 (N_4232,N_3725,N_3897);
xnor U4233 (N_4233,N_3546,N_3901);
xor U4234 (N_4234,N_3853,N_3884);
or U4235 (N_4235,N_3794,N_3916);
nand U4236 (N_4236,N_3929,N_3835);
nand U4237 (N_4237,N_3505,N_3551);
and U4238 (N_4238,N_3608,N_3919);
and U4239 (N_4239,N_3796,N_3671);
xor U4240 (N_4240,N_3713,N_3503);
nand U4241 (N_4241,N_3672,N_3615);
and U4242 (N_4242,N_3772,N_3925);
or U4243 (N_4243,N_3984,N_3861);
nand U4244 (N_4244,N_3645,N_3783);
and U4245 (N_4245,N_3763,N_3791);
xor U4246 (N_4246,N_3501,N_3576);
and U4247 (N_4247,N_3912,N_3578);
and U4248 (N_4248,N_3930,N_3886);
nor U4249 (N_4249,N_3584,N_3524);
nor U4250 (N_4250,N_3747,N_3570);
nor U4251 (N_4251,N_3678,N_3890);
and U4252 (N_4252,N_3577,N_3701);
or U4253 (N_4253,N_3531,N_3919);
and U4254 (N_4254,N_3725,N_3886);
xor U4255 (N_4255,N_3851,N_3749);
nor U4256 (N_4256,N_3953,N_3723);
xnor U4257 (N_4257,N_3779,N_3920);
or U4258 (N_4258,N_3586,N_3856);
nand U4259 (N_4259,N_3505,N_3681);
or U4260 (N_4260,N_3863,N_3843);
nand U4261 (N_4261,N_3985,N_3622);
or U4262 (N_4262,N_3924,N_3509);
nor U4263 (N_4263,N_3870,N_3631);
nand U4264 (N_4264,N_3652,N_3956);
or U4265 (N_4265,N_3843,N_3524);
xor U4266 (N_4266,N_3660,N_3524);
or U4267 (N_4267,N_3860,N_3822);
xor U4268 (N_4268,N_3563,N_3844);
nor U4269 (N_4269,N_3565,N_3886);
and U4270 (N_4270,N_3799,N_3591);
and U4271 (N_4271,N_3542,N_3788);
or U4272 (N_4272,N_3602,N_3764);
nor U4273 (N_4273,N_3896,N_3647);
xor U4274 (N_4274,N_3892,N_3882);
nand U4275 (N_4275,N_3825,N_3567);
nand U4276 (N_4276,N_3634,N_3867);
xor U4277 (N_4277,N_3538,N_3605);
nand U4278 (N_4278,N_3924,N_3522);
and U4279 (N_4279,N_3800,N_3809);
nand U4280 (N_4280,N_3621,N_3835);
xnor U4281 (N_4281,N_3964,N_3524);
nor U4282 (N_4282,N_3987,N_3900);
and U4283 (N_4283,N_3651,N_3677);
nand U4284 (N_4284,N_3757,N_3639);
xnor U4285 (N_4285,N_3525,N_3662);
nand U4286 (N_4286,N_3689,N_3722);
xnor U4287 (N_4287,N_3929,N_3523);
and U4288 (N_4288,N_3753,N_3885);
nand U4289 (N_4289,N_3560,N_3537);
xor U4290 (N_4290,N_3572,N_3581);
nor U4291 (N_4291,N_3600,N_3766);
or U4292 (N_4292,N_3894,N_3600);
and U4293 (N_4293,N_3524,N_3655);
nor U4294 (N_4294,N_3892,N_3834);
nor U4295 (N_4295,N_3782,N_3962);
nor U4296 (N_4296,N_3598,N_3870);
xnor U4297 (N_4297,N_3720,N_3639);
xnor U4298 (N_4298,N_3662,N_3601);
nand U4299 (N_4299,N_3568,N_3884);
xnor U4300 (N_4300,N_3647,N_3616);
and U4301 (N_4301,N_3503,N_3703);
nor U4302 (N_4302,N_3845,N_3786);
nor U4303 (N_4303,N_3893,N_3673);
xnor U4304 (N_4304,N_3913,N_3945);
or U4305 (N_4305,N_3739,N_3950);
and U4306 (N_4306,N_3764,N_3963);
nand U4307 (N_4307,N_3760,N_3656);
xor U4308 (N_4308,N_3529,N_3972);
nor U4309 (N_4309,N_3878,N_3689);
xnor U4310 (N_4310,N_3524,N_3513);
nand U4311 (N_4311,N_3739,N_3572);
xnor U4312 (N_4312,N_3578,N_3854);
nand U4313 (N_4313,N_3603,N_3725);
nand U4314 (N_4314,N_3534,N_3793);
nand U4315 (N_4315,N_3643,N_3813);
xor U4316 (N_4316,N_3523,N_3601);
nor U4317 (N_4317,N_3679,N_3810);
nand U4318 (N_4318,N_3611,N_3653);
and U4319 (N_4319,N_3834,N_3890);
xnor U4320 (N_4320,N_3709,N_3867);
nor U4321 (N_4321,N_3787,N_3778);
and U4322 (N_4322,N_3966,N_3990);
or U4323 (N_4323,N_3814,N_3559);
and U4324 (N_4324,N_3521,N_3792);
and U4325 (N_4325,N_3867,N_3659);
and U4326 (N_4326,N_3927,N_3866);
and U4327 (N_4327,N_3582,N_3632);
or U4328 (N_4328,N_3895,N_3584);
or U4329 (N_4329,N_3598,N_3851);
or U4330 (N_4330,N_3643,N_3907);
and U4331 (N_4331,N_3718,N_3620);
or U4332 (N_4332,N_3967,N_3663);
nor U4333 (N_4333,N_3851,N_3669);
xor U4334 (N_4334,N_3852,N_3679);
nand U4335 (N_4335,N_3591,N_3665);
nor U4336 (N_4336,N_3572,N_3540);
and U4337 (N_4337,N_3817,N_3893);
xor U4338 (N_4338,N_3671,N_3602);
xnor U4339 (N_4339,N_3832,N_3865);
or U4340 (N_4340,N_3523,N_3948);
and U4341 (N_4341,N_3996,N_3981);
xor U4342 (N_4342,N_3598,N_3712);
and U4343 (N_4343,N_3830,N_3665);
nand U4344 (N_4344,N_3671,N_3620);
or U4345 (N_4345,N_3859,N_3721);
nand U4346 (N_4346,N_3900,N_3689);
nand U4347 (N_4347,N_3701,N_3841);
nand U4348 (N_4348,N_3803,N_3920);
nand U4349 (N_4349,N_3576,N_3702);
or U4350 (N_4350,N_3658,N_3625);
and U4351 (N_4351,N_3557,N_3779);
and U4352 (N_4352,N_3943,N_3958);
xor U4353 (N_4353,N_3810,N_3709);
or U4354 (N_4354,N_3831,N_3662);
or U4355 (N_4355,N_3565,N_3510);
nand U4356 (N_4356,N_3558,N_3652);
and U4357 (N_4357,N_3670,N_3518);
xnor U4358 (N_4358,N_3988,N_3915);
xnor U4359 (N_4359,N_3768,N_3778);
and U4360 (N_4360,N_3508,N_3814);
and U4361 (N_4361,N_3750,N_3955);
nor U4362 (N_4362,N_3624,N_3787);
xnor U4363 (N_4363,N_3611,N_3609);
and U4364 (N_4364,N_3651,N_3850);
or U4365 (N_4365,N_3585,N_3875);
or U4366 (N_4366,N_3840,N_3554);
and U4367 (N_4367,N_3981,N_3573);
and U4368 (N_4368,N_3883,N_3789);
xnor U4369 (N_4369,N_3741,N_3943);
and U4370 (N_4370,N_3586,N_3532);
nand U4371 (N_4371,N_3903,N_3712);
or U4372 (N_4372,N_3567,N_3881);
xor U4373 (N_4373,N_3844,N_3654);
or U4374 (N_4374,N_3816,N_3594);
nor U4375 (N_4375,N_3511,N_3931);
nand U4376 (N_4376,N_3850,N_3711);
nand U4377 (N_4377,N_3888,N_3681);
nand U4378 (N_4378,N_3614,N_3513);
xor U4379 (N_4379,N_3684,N_3975);
xnor U4380 (N_4380,N_3723,N_3614);
nor U4381 (N_4381,N_3911,N_3721);
xnor U4382 (N_4382,N_3692,N_3779);
xor U4383 (N_4383,N_3574,N_3684);
nor U4384 (N_4384,N_3847,N_3600);
nor U4385 (N_4385,N_3713,N_3875);
and U4386 (N_4386,N_3920,N_3552);
xnor U4387 (N_4387,N_3702,N_3927);
or U4388 (N_4388,N_3878,N_3877);
and U4389 (N_4389,N_3932,N_3870);
xor U4390 (N_4390,N_3861,N_3729);
nor U4391 (N_4391,N_3521,N_3691);
or U4392 (N_4392,N_3790,N_3993);
or U4393 (N_4393,N_3984,N_3633);
xnor U4394 (N_4394,N_3935,N_3596);
nor U4395 (N_4395,N_3816,N_3727);
or U4396 (N_4396,N_3911,N_3537);
or U4397 (N_4397,N_3950,N_3789);
xor U4398 (N_4398,N_3676,N_3562);
nor U4399 (N_4399,N_3560,N_3647);
nor U4400 (N_4400,N_3568,N_3688);
xnor U4401 (N_4401,N_3743,N_3748);
xor U4402 (N_4402,N_3694,N_3722);
nand U4403 (N_4403,N_3621,N_3521);
or U4404 (N_4404,N_3603,N_3579);
and U4405 (N_4405,N_3855,N_3609);
or U4406 (N_4406,N_3508,N_3936);
xor U4407 (N_4407,N_3641,N_3833);
nor U4408 (N_4408,N_3906,N_3957);
or U4409 (N_4409,N_3923,N_3615);
nand U4410 (N_4410,N_3926,N_3582);
or U4411 (N_4411,N_3826,N_3672);
xor U4412 (N_4412,N_3592,N_3891);
nand U4413 (N_4413,N_3639,N_3932);
nand U4414 (N_4414,N_3785,N_3537);
and U4415 (N_4415,N_3642,N_3555);
and U4416 (N_4416,N_3501,N_3709);
and U4417 (N_4417,N_3957,N_3673);
nand U4418 (N_4418,N_3955,N_3582);
nand U4419 (N_4419,N_3756,N_3516);
and U4420 (N_4420,N_3653,N_3657);
xor U4421 (N_4421,N_3963,N_3794);
nor U4422 (N_4422,N_3946,N_3812);
nor U4423 (N_4423,N_3736,N_3902);
nand U4424 (N_4424,N_3798,N_3790);
nor U4425 (N_4425,N_3512,N_3824);
nand U4426 (N_4426,N_3671,N_3570);
and U4427 (N_4427,N_3818,N_3554);
or U4428 (N_4428,N_3716,N_3651);
and U4429 (N_4429,N_3611,N_3789);
and U4430 (N_4430,N_3746,N_3618);
nand U4431 (N_4431,N_3595,N_3979);
nand U4432 (N_4432,N_3891,N_3849);
or U4433 (N_4433,N_3787,N_3897);
nand U4434 (N_4434,N_3985,N_3621);
nor U4435 (N_4435,N_3974,N_3930);
nor U4436 (N_4436,N_3528,N_3770);
and U4437 (N_4437,N_3800,N_3817);
or U4438 (N_4438,N_3973,N_3933);
nand U4439 (N_4439,N_3762,N_3533);
nand U4440 (N_4440,N_3726,N_3590);
and U4441 (N_4441,N_3522,N_3885);
or U4442 (N_4442,N_3620,N_3795);
and U4443 (N_4443,N_3602,N_3692);
or U4444 (N_4444,N_3776,N_3863);
or U4445 (N_4445,N_3808,N_3993);
and U4446 (N_4446,N_3924,N_3589);
nor U4447 (N_4447,N_3935,N_3743);
and U4448 (N_4448,N_3733,N_3682);
nor U4449 (N_4449,N_3865,N_3798);
nor U4450 (N_4450,N_3871,N_3653);
nor U4451 (N_4451,N_3688,N_3608);
nand U4452 (N_4452,N_3841,N_3966);
nor U4453 (N_4453,N_3688,N_3749);
xnor U4454 (N_4454,N_3523,N_3812);
nor U4455 (N_4455,N_3557,N_3751);
xor U4456 (N_4456,N_3986,N_3570);
nand U4457 (N_4457,N_3707,N_3560);
or U4458 (N_4458,N_3767,N_3688);
xnor U4459 (N_4459,N_3827,N_3631);
or U4460 (N_4460,N_3720,N_3525);
nand U4461 (N_4461,N_3641,N_3730);
nor U4462 (N_4462,N_3565,N_3827);
nand U4463 (N_4463,N_3787,N_3665);
and U4464 (N_4464,N_3730,N_3713);
nor U4465 (N_4465,N_3537,N_3702);
nor U4466 (N_4466,N_3529,N_3524);
nor U4467 (N_4467,N_3631,N_3603);
nand U4468 (N_4468,N_3856,N_3890);
xor U4469 (N_4469,N_3981,N_3794);
nor U4470 (N_4470,N_3727,N_3824);
xor U4471 (N_4471,N_3574,N_3760);
and U4472 (N_4472,N_3606,N_3883);
nor U4473 (N_4473,N_3826,N_3852);
or U4474 (N_4474,N_3992,N_3779);
nand U4475 (N_4475,N_3991,N_3948);
nand U4476 (N_4476,N_3886,N_3512);
and U4477 (N_4477,N_3696,N_3683);
nand U4478 (N_4478,N_3919,N_3610);
xnor U4479 (N_4479,N_3809,N_3791);
or U4480 (N_4480,N_3823,N_3618);
nand U4481 (N_4481,N_3606,N_3841);
or U4482 (N_4482,N_3940,N_3830);
xor U4483 (N_4483,N_3570,N_3544);
xnor U4484 (N_4484,N_3995,N_3910);
or U4485 (N_4485,N_3904,N_3586);
nand U4486 (N_4486,N_3880,N_3933);
or U4487 (N_4487,N_3914,N_3734);
nor U4488 (N_4488,N_3928,N_3876);
nand U4489 (N_4489,N_3945,N_3749);
or U4490 (N_4490,N_3917,N_3744);
or U4491 (N_4491,N_3571,N_3888);
or U4492 (N_4492,N_3883,N_3611);
nand U4493 (N_4493,N_3612,N_3500);
or U4494 (N_4494,N_3634,N_3915);
xor U4495 (N_4495,N_3604,N_3536);
nor U4496 (N_4496,N_3679,N_3859);
nand U4497 (N_4497,N_3674,N_3861);
nand U4498 (N_4498,N_3954,N_3884);
or U4499 (N_4499,N_3828,N_3576);
nor U4500 (N_4500,N_4371,N_4466);
xor U4501 (N_4501,N_4127,N_4388);
and U4502 (N_4502,N_4032,N_4031);
nor U4503 (N_4503,N_4039,N_4397);
xor U4504 (N_4504,N_4427,N_4376);
and U4505 (N_4505,N_4047,N_4152);
or U4506 (N_4506,N_4210,N_4363);
nor U4507 (N_4507,N_4000,N_4366);
nand U4508 (N_4508,N_4062,N_4431);
nand U4509 (N_4509,N_4475,N_4453);
xor U4510 (N_4510,N_4183,N_4214);
and U4511 (N_4511,N_4356,N_4184);
and U4512 (N_4512,N_4104,N_4156);
xnor U4513 (N_4513,N_4211,N_4041);
nand U4514 (N_4514,N_4442,N_4498);
nand U4515 (N_4515,N_4300,N_4418);
xnor U4516 (N_4516,N_4150,N_4235);
and U4517 (N_4517,N_4261,N_4415);
nor U4518 (N_4518,N_4058,N_4155);
nor U4519 (N_4519,N_4111,N_4189);
nand U4520 (N_4520,N_4249,N_4128);
and U4521 (N_4521,N_4484,N_4190);
nor U4522 (N_4522,N_4030,N_4268);
xnor U4523 (N_4523,N_4055,N_4180);
and U4524 (N_4524,N_4382,N_4037);
nand U4525 (N_4525,N_4368,N_4277);
nor U4526 (N_4526,N_4467,N_4434);
nor U4527 (N_4527,N_4452,N_4425);
or U4528 (N_4528,N_4009,N_4213);
xor U4529 (N_4529,N_4491,N_4384);
nand U4530 (N_4530,N_4473,N_4309);
xor U4531 (N_4531,N_4424,N_4135);
xnor U4532 (N_4532,N_4114,N_4094);
and U4533 (N_4533,N_4014,N_4308);
or U4534 (N_4534,N_4153,N_4499);
nor U4535 (N_4535,N_4051,N_4092);
or U4536 (N_4536,N_4050,N_4107);
or U4537 (N_4537,N_4400,N_4218);
nor U4538 (N_4538,N_4004,N_4337);
nand U4539 (N_4539,N_4341,N_4066);
xor U4540 (N_4540,N_4089,N_4237);
or U4541 (N_4541,N_4377,N_4318);
and U4542 (N_4542,N_4271,N_4296);
nor U4543 (N_4543,N_4082,N_4239);
nand U4544 (N_4544,N_4008,N_4285);
xor U4545 (N_4545,N_4305,N_4005);
nor U4546 (N_4546,N_4310,N_4487);
or U4547 (N_4547,N_4421,N_4206);
nand U4548 (N_4548,N_4345,N_4049);
nand U4549 (N_4549,N_4381,N_4294);
or U4550 (N_4550,N_4406,N_4228);
or U4551 (N_4551,N_4486,N_4369);
xor U4552 (N_4552,N_4247,N_4125);
nor U4553 (N_4553,N_4358,N_4284);
or U4554 (N_4554,N_4026,N_4459);
and U4555 (N_4555,N_4441,N_4251);
nand U4556 (N_4556,N_4478,N_4387);
nand U4557 (N_4557,N_4359,N_4367);
nor U4558 (N_4558,N_4464,N_4013);
nand U4559 (N_4559,N_4056,N_4455);
and U4560 (N_4560,N_4236,N_4410);
or U4561 (N_4561,N_4469,N_4343);
or U4562 (N_4562,N_4462,N_4091);
xnor U4563 (N_4563,N_4053,N_4188);
nor U4564 (N_4564,N_4465,N_4182);
or U4565 (N_4565,N_4109,N_4169);
nor U4566 (N_4566,N_4196,N_4163);
nor U4567 (N_4567,N_4390,N_4302);
and U4568 (N_4568,N_4223,N_4186);
nor U4569 (N_4569,N_4413,N_4185);
or U4570 (N_4570,N_4042,N_4395);
xnor U4571 (N_4571,N_4170,N_4048);
or U4572 (N_4572,N_4205,N_4342);
nor U4573 (N_4573,N_4322,N_4244);
and U4574 (N_4574,N_4178,N_4181);
xnor U4575 (N_4575,N_4079,N_4429);
and U4576 (N_4576,N_4283,N_4315);
xor U4577 (N_4577,N_4176,N_4379);
nor U4578 (N_4578,N_4269,N_4179);
and U4579 (N_4579,N_4344,N_4138);
nor U4580 (N_4580,N_4207,N_4099);
nand U4581 (N_4581,N_4088,N_4033);
or U4582 (N_4582,N_4142,N_4312);
xnor U4583 (N_4583,N_4298,N_4102);
nor U4584 (N_4584,N_4383,N_4215);
nor U4585 (N_4585,N_4291,N_4451);
or U4586 (N_4586,N_4131,N_4497);
xnor U4587 (N_4587,N_4490,N_4168);
xor U4588 (N_4588,N_4350,N_4242);
nand U4589 (N_4589,N_4157,N_4398);
xnor U4590 (N_4590,N_4392,N_4192);
nand U4591 (N_4591,N_4311,N_4015);
and U4592 (N_4592,N_4077,N_4220);
nor U4593 (N_4593,N_4252,N_4304);
nand U4594 (N_4594,N_4248,N_4069);
and U4595 (N_4595,N_4165,N_4212);
xnor U4596 (N_4596,N_4450,N_4065);
nand U4597 (N_4597,N_4333,N_4208);
or U4598 (N_4598,N_4454,N_4297);
nor U4599 (N_4599,N_4468,N_4231);
and U4600 (N_4600,N_4007,N_4044);
nand U4601 (N_4601,N_4265,N_4103);
or U4602 (N_4602,N_4476,N_4159);
nand U4603 (N_4603,N_4115,N_4054);
or U4604 (N_4604,N_4448,N_4154);
and U4605 (N_4605,N_4279,N_4480);
and U4606 (N_4606,N_4313,N_4361);
and U4607 (N_4607,N_4199,N_4141);
xor U4608 (N_4608,N_4360,N_4443);
and U4609 (N_4609,N_4263,N_4105);
xor U4610 (N_4610,N_4430,N_4391);
nor U4611 (N_4611,N_4362,N_4060);
xnor U4612 (N_4612,N_4234,N_4130);
nand U4613 (N_4613,N_4003,N_4258);
nor U4614 (N_4614,N_4243,N_4164);
nand U4615 (N_4615,N_4422,N_4238);
or U4616 (N_4616,N_4194,N_4028);
nand U4617 (N_4617,N_4106,N_4137);
nor U4618 (N_4618,N_4162,N_4483);
and U4619 (N_4619,N_4113,N_4002);
nor U4620 (N_4620,N_4017,N_4436);
and U4621 (N_4621,N_4299,N_4426);
xor U4622 (N_4622,N_4193,N_4319);
xnor U4623 (N_4623,N_4016,N_4257);
and U4624 (N_4624,N_4440,N_4120);
nor U4625 (N_4625,N_4229,N_4045);
nor U4626 (N_4626,N_4063,N_4064);
nor U4627 (N_4627,N_4197,N_4394);
nand U4628 (N_4628,N_4078,N_4292);
nand U4629 (N_4629,N_4389,N_4290);
nor U4630 (N_4630,N_4428,N_4352);
xnor U4631 (N_4631,N_4320,N_4432);
or U4632 (N_4632,N_4123,N_4472);
or U4633 (N_4633,N_4357,N_4256);
and U4634 (N_4634,N_4110,N_4331);
nand U4635 (N_4635,N_4101,N_4353);
xnor U4636 (N_4636,N_4334,N_4492);
or U4637 (N_4637,N_4083,N_4272);
xor U4638 (N_4638,N_4171,N_4340);
or U4639 (N_4639,N_4372,N_4346);
xnor U4640 (N_4640,N_4405,N_4494);
nor U4641 (N_4641,N_4276,N_4253);
or U4642 (N_4642,N_4219,N_4403);
and U4643 (N_4643,N_4006,N_4489);
xnor U4644 (N_4644,N_4386,N_4022);
or U4645 (N_4645,N_4108,N_4437);
nand U4646 (N_4646,N_4295,N_4025);
xor U4647 (N_4647,N_4187,N_4250);
and U4648 (N_4648,N_4275,N_4330);
nor U4649 (N_4649,N_4457,N_4332);
and U4650 (N_4650,N_4325,N_4323);
xnor U4651 (N_4651,N_4148,N_4393);
nor U4652 (N_4652,N_4221,N_4074);
nand U4653 (N_4653,N_4118,N_4446);
nand U4654 (N_4654,N_4241,N_4495);
xnor U4655 (N_4655,N_4160,N_4399);
or U4656 (N_4656,N_4433,N_4067);
or U4657 (N_4657,N_4378,N_4195);
and U4658 (N_4658,N_4059,N_4226);
nor U4659 (N_4659,N_4012,N_4177);
xor U4660 (N_4660,N_4493,N_4460);
and U4661 (N_4661,N_4317,N_4336);
and U4662 (N_4662,N_4282,N_4068);
nand U4663 (N_4663,N_4321,N_4412);
or U4664 (N_4664,N_4408,N_4174);
nand U4665 (N_4665,N_4140,N_4380);
or U4666 (N_4666,N_4349,N_4175);
nand U4667 (N_4667,N_4146,N_4096);
or U4668 (N_4668,N_4144,N_4365);
or U4669 (N_4669,N_4445,N_4095);
or U4670 (N_4670,N_4435,N_4203);
and U4671 (N_4671,N_4011,N_4348);
or U4672 (N_4672,N_4129,N_4139);
and U4673 (N_4673,N_4266,N_4073);
xor U4674 (N_4674,N_4409,N_4071);
and U4675 (N_4675,N_4347,N_4301);
and U4676 (N_4676,N_4246,N_4200);
or U4677 (N_4677,N_4136,N_4438);
nor U4678 (N_4678,N_4364,N_4018);
or U4679 (N_4679,N_4419,N_4477);
xnor U4680 (N_4680,N_4072,N_4307);
xor U4681 (N_4681,N_4270,N_4474);
or U4682 (N_4682,N_4161,N_4401);
nor U4683 (N_4683,N_4267,N_4151);
nor U4684 (N_4684,N_4233,N_4209);
or U4685 (N_4685,N_4149,N_4134);
nand U4686 (N_4686,N_4339,N_4335);
xor U4687 (N_4687,N_4122,N_4133);
or U4688 (N_4688,N_4034,N_4230);
nand U4689 (N_4689,N_4070,N_4288);
nand U4690 (N_4690,N_4173,N_4293);
or U4691 (N_4691,N_4046,N_4204);
or U4692 (N_4692,N_4076,N_4191);
nand U4693 (N_4693,N_4198,N_4132);
or U4694 (N_4694,N_4402,N_4264);
nand U4695 (N_4695,N_4479,N_4040);
xor U4696 (N_4696,N_4035,N_4222);
xor U4697 (N_4697,N_4314,N_4444);
nor U4698 (N_4698,N_4057,N_4216);
and U4699 (N_4699,N_4225,N_4355);
or U4700 (N_4700,N_4087,N_4100);
nor U4701 (N_4701,N_4326,N_4485);
nor U4702 (N_4702,N_4481,N_4232);
xnor U4703 (N_4703,N_4385,N_4396);
nor U4704 (N_4704,N_4423,N_4254);
nor U4705 (N_4705,N_4463,N_4021);
nand U4706 (N_4706,N_4496,N_4081);
nand U4707 (N_4707,N_4374,N_4027);
and U4708 (N_4708,N_4217,N_4086);
nor U4709 (N_4709,N_4407,N_4224);
nand U4710 (N_4710,N_4080,N_4201);
and U4711 (N_4711,N_4098,N_4471);
xor U4712 (N_4712,N_4354,N_4166);
xnor U4713 (N_4713,N_4488,N_4351);
nor U4714 (N_4714,N_4167,N_4019);
xor U4715 (N_4715,N_4172,N_4416);
nand U4716 (N_4716,N_4280,N_4143);
nor U4717 (N_4717,N_4090,N_4112);
xnor U4718 (N_4718,N_4278,N_4255);
or U4719 (N_4719,N_4119,N_4411);
or U4720 (N_4720,N_4001,N_4202);
or U4721 (N_4721,N_4117,N_4449);
nand U4722 (N_4722,N_4158,N_4482);
nand U4723 (N_4723,N_4262,N_4327);
nand U4724 (N_4724,N_4097,N_4287);
xor U4725 (N_4725,N_4328,N_4145);
or U4726 (N_4726,N_4324,N_4259);
nor U4727 (N_4727,N_4085,N_4052);
or U4728 (N_4728,N_4456,N_4329);
or U4729 (N_4729,N_4036,N_4020);
nor U4730 (N_4730,N_4370,N_4286);
nand U4731 (N_4731,N_4075,N_4375);
xor U4732 (N_4732,N_4439,N_4470);
or U4733 (N_4733,N_4338,N_4024);
nand U4734 (N_4734,N_4240,N_4414);
xor U4735 (N_4735,N_4116,N_4274);
and U4736 (N_4736,N_4061,N_4126);
nand U4737 (N_4737,N_4043,N_4084);
nand U4738 (N_4738,N_4093,N_4260);
and U4739 (N_4739,N_4461,N_4447);
xnor U4740 (N_4740,N_4147,N_4029);
xor U4741 (N_4741,N_4373,N_4124);
nand U4742 (N_4742,N_4245,N_4316);
xnor U4743 (N_4743,N_4010,N_4273);
xor U4744 (N_4744,N_4303,N_4404);
nand U4745 (N_4745,N_4038,N_4306);
xnor U4746 (N_4746,N_4281,N_4417);
xor U4747 (N_4747,N_4420,N_4289);
xnor U4748 (N_4748,N_4227,N_4023);
or U4749 (N_4749,N_4458,N_4121);
and U4750 (N_4750,N_4114,N_4269);
and U4751 (N_4751,N_4113,N_4448);
or U4752 (N_4752,N_4296,N_4320);
and U4753 (N_4753,N_4354,N_4407);
nor U4754 (N_4754,N_4267,N_4436);
or U4755 (N_4755,N_4460,N_4237);
nand U4756 (N_4756,N_4419,N_4426);
or U4757 (N_4757,N_4081,N_4326);
or U4758 (N_4758,N_4498,N_4199);
nand U4759 (N_4759,N_4103,N_4400);
nand U4760 (N_4760,N_4122,N_4492);
or U4761 (N_4761,N_4214,N_4052);
and U4762 (N_4762,N_4194,N_4460);
and U4763 (N_4763,N_4157,N_4325);
or U4764 (N_4764,N_4478,N_4037);
or U4765 (N_4765,N_4452,N_4193);
nor U4766 (N_4766,N_4194,N_4382);
and U4767 (N_4767,N_4199,N_4198);
nor U4768 (N_4768,N_4296,N_4356);
nor U4769 (N_4769,N_4070,N_4158);
nand U4770 (N_4770,N_4267,N_4441);
nand U4771 (N_4771,N_4337,N_4051);
nand U4772 (N_4772,N_4055,N_4104);
xnor U4773 (N_4773,N_4037,N_4191);
nand U4774 (N_4774,N_4091,N_4417);
xor U4775 (N_4775,N_4040,N_4172);
nor U4776 (N_4776,N_4027,N_4110);
or U4777 (N_4777,N_4114,N_4264);
nor U4778 (N_4778,N_4136,N_4355);
nor U4779 (N_4779,N_4152,N_4498);
or U4780 (N_4780,N_4167,N_4297);
nand U4781 (N_4781,N_4239,N_4277);
nand U4782 (N_4782,N_4255,N_4486);
xor U4783 (N_4783,N_4498,N_4188);
xnor U4784 (N_4784,N_4418,N_4132);
and U4785 (N_4785,N_4330,N_4040);
and U4786 (N_4786,N_4268,N_4415);
or U4787 (N_4787,N_4036,N_4012);
xnor U4788 (N_4788,N_4025,N_4019);
nor U4789 (N_4789,N_4100,N_4463);
nor U4790 (N_4790,N_4257,N_4260);
nor U4791 (N_4791,N_4143,N_4457);
xor U4792 (N_4792,N_4053,N_4397);
nand U4793 (N_4793,N_4367,N_4075);
nor U4794 (N_4794,N_4420,N_4115);
nor U4795 (N_4795,N_4033,N_4424);
or U4796 (N_4796,N_4071,N_4173);
nand U4797 (N_4797,N_4329,N_4250);
xor U4798 (N_4798,N_4082,N_4144);
nor U4799 (N_4799,N_4029,N_4096);
and U4800 (N_4800,N_4412,N_4319);
nand U4801 (N_4801,N_4284,N_4422);
nor U4802 (N_4802,N_4324,N_4186);
nor U4803 (N_4803,N_4240,N_4423);
or U4804 (N_4804,N_4458,N_4085);
xor U4805 (N_4805,N_4254,N_4455);
or U4806 (N_4806,N_4085,N_4373);
or U4807 (N_4807,N_4115,N_4422);
xnor U4808 (N_4808,N_4406,N_4331);
and U4809 (N_4809,N_4226,N_4372);
xor U4810 (N_4810,N_4191,N_4166);
and U4811 (N_4811,N_4384,N_4024);
or U4812 (N_4812,N_4064,N_4005);
and U4813 (N_4813,N_4427,N_4308);
and U4814 (N_4814,N_4094,N_4241);
xnor U4815 (N_4815,N_4440,N_4313);
or U4816 (N_4816,N_4227,N_4190);
and U4817 (N_4817,N_4116,N_4276);
nor U4818 (N_4818,N_4478,N_4494);
nor U4819 (N_4819,N_4017,N_4360);
nor U4820 (N_4820,N_4017,N_4021);
or U4821 (N_4821,N_4419,N_4464);
and U4822 (N_4822,N_4120,N_4100);
nand U4823 (N_4823,N_4021,N_4496);
or U4824 (N_4824,N_4438,N_4183);
and U4825 (N_4825,N_4367,N_4274);
xor U4826 (N_4826,N_4357,N_4098);
nor U4827 (N_4827,N_4067,N_4097);
nor U4828 (N_4828,N_4458,N_4177);
nor U4829 (N_4829,N_4311,N_4076);
and U4830 (N_4830,N_4237,N_4061);
and U4831 (N_4831,N_4229,N_4089);
or U4832 (N_4832,N_4063,N_4238);
xnor U4833 (N_4833,N_4237,N_4385);
nor U4834 (N_4834,N_4145,N_4402);
nor U4835 (N_4835,N_4321,N_4314);
and U4836 (N_4836,N_4445,N_4196);
xor U4837 (N_4837,N_4336,N_4275);
nand U4838 (N_4838,N_4247,N_4337);
or U4839 (N_4839,N_4383,N_4085);
xnor U4840 (N_4840,N_4176,N_4486);
xor U4841 (N_4841,N_4291,N_4288);
nand U4842 (N_4842,N_4192,N_4342);
and U4843 (N_4843,N_4457,N_4364);
or U4844 (N_4844,N_4319,N_4468);
xor U4845 (N_4845,N_4254,N_4475);
nand U4846 (N_4846,N_4102,N_4461);
xnor U4847 (N_4847,N_4157,N_4271);
nand U4848 (N_4848,N_4180,N_4006);
xnor U4849 (N_4849,N_4280,N_4355);
xor U4850 (N_4850,N_4347,N_4317);
nor U4851 (N_4851,N_4092,N_4259);
xnor U4852 (N_4852,N_4228,N_4304);
xnor U4853 (N_4853,N_4161,N_4286);
nor U4854 (N_4854,N_4088,N_4384);
nor U4855 (N_4855,N_4116,N_4038);
nor U4856 (N_4856,N_4293,N_4163);
and U4857 (N_4857,N_4342,N_4173);
nor U4858 (N_4858,N_4027,N_4433);
nand U4859 (N_4859,N_4264,N_4113);
xnor U4860 (N_4860,N_4302,N_4243);
and U4861 (N_4861,N_4277,N_4305);
nand U4862 (N_4862,N_4034,N_4373);
nand U4863 (N_4863,N_4456,N_4014);
nand U4864 (N_4864,N_4202,N_4427);
xnor U4865 (N_4865,N_4442,N_4458);
and U4866 (N_4866,N_4444,N_4440);
nand U4867 (N_4867,N_4089,N_4256);
or U4868 (N_4868,N_4022,N_4338);
nor U4869 (N_4869,N_4208,N_4290);
or U4870 (N_4870,N_4133,N_4456);
xnor U4871 (N_4871,N_4296,N_4383);
nor U4872 (N_4872,N_4396,N_4235);
or U4873 (N_4873,N_4082,N_4494);
nor U4874 (N_4874,N_4327,N_4303);
nand U4875 (N_4875,N_4471,N_4019);
nand U4876 (N_4876,N_4317,N_4389);
or U4877 (N_4877,N_4289,N_4179);
nor U4878 (N_4878,N_4245,N_4494);
or U4879 (N_4879,N_4292,N_4355);
xnor U4880 (N_4880,N_4349,N_4014);
nand U4881 (N_4881,N_4380,N_4288);
nor U4882 (N_4882,N_4304,N_4309);
nand U4883 (N_4883,N_4410,N_4370);
or U4884 (N_4884,N_4161,N_4115);
nor U4885 (N_4885,N_4467,N_4431);
nor U4886 (N_4886,N_4495,N_4374);
xnor U4887 (N_4887,N_4185,N_4368);
xor U4888 (N_4888,N_4417,N_4374);
and U4889 (N_4889,N_4352,N_4164);
or U4890 (N_4890,N_4163,N_4381);
and U4891 (N_4891,N_4065,N_4096);
and U4892 (N_4892,N_4092,N_4056);
and U4893 (N_4893,N_4392,N_4110);
and U4894 (N_4894,N_4353,N_4146);
nor U4895 (N_4895,N_4493,N_4188);
and U4896 (N_4896,N_4343,N_4227);
xor U4897 (N_4897,N_4209,N_4337);
or U4898 (N_4898,N_4325,N_4068);
xor U4899 (N_4899,N_4444,N_4352);
or U4900 (N_4900,N_4015,N_4439);
xnor U4901 (N_4901,N_4494,N_4262);
xnor U4902 (N_4902,N_4156,N_4283);
and U4903 (N_4903,N_4234,N_4070);
xnor U4904 (N_4904,N_4392,N_4218);
nor U4905 (N_4905,N_4035,N_4125);
xnor U4906 (N_4906,N_4440,N_4079);
nor U4907 (N_4907,N_4296,N_4456);
nand U4908 (N_4908,N_4195,N_4328);
nand U4909 (N_4909,N_4181,N_4187);
xnor U4910 (N_4910,N_4248,N_4196);
xor U4911 (N_4911,N_4084,N_4374);
nor U4912 (N_4912,N_4315,N_4290);
nor U4913 (N_4913,N_4459,N_4132);
and U4914 (N_4914,N_4119,N_4090);
nand U4915 (N_4915,N_4378,N_4403);
nand U4916 (N_4916,N_4439,N_4168);
xnor U4917 (N_4917,N_4486,N_4245);
and U4918 (N_4918,N_4057,N_4305);
nor U4919 (N_4919,N_4132,N_4247);
nor U4920 (N_4920,N_4221,N_4063);
xor U4921 (N_4921,N_4064,N_4210);
and U4922 (N_4922,N_4068,N_4368);
and U4923 (N_4923,N_4324,N_4340);
nand U4924 (N_4924,N_4146,N_4428);
xor U4925 (N_4925,N_4415,N_4342);
and U4926 (N_4926,N_4361,N_4293);
xnor U4927 (N_4927,N_4470,N_4233);
nand U4928 (N_4928,N_4243,N_4258);
nand U4929 (N_4929,N_4102,N_4320);
xor U4930 (N_4930,N_4037,N_4232);
xor U4931 (N_4931,N_4278,N_4409);
nand U4932 (N_4932,N_4290,N_4472);
nor U4933 (N_4933,N_4359,N_4184);
nor U4934 (N_4934,N_4264,N_4247);
xnor U4935 (N_4935,N_4297,N_4194);
nand U4936 (N_4936,N_4028,N_4320);
xor U4937 (N_4937,N_4278,N_4288);
and U4938 (N_4938,N_4162,N_4300);
xor U4939 (N_4939,N_4235,N_4169);
nand U4940 (N_4940,N_4163,N_4090);
and U4941 (N_4941,N_4274,N_4057);
and U4942 (N_4942,N_4343,N_4198);
or U4943 (N_4943,N_4080,N_4183);
xnor U4944 (N_4944,N_4460,N_4461);
nand U4945 (N_4945,N_4004,N_4388);
nand U4946 (N_4946,N_4084,N_4147);
nand U4947 (N_4947,N_4316,N_4028);
xor U4948 (N_4948,N_4483,N_4415);
and U4949 (N_4949,N_4162,N_4161);
nor U4950 (N_4950,N_4338,N_4242);
xnor U4951 (N_4951,N_4089,N_4161);
xor U4952 (N_4952,N_4025,N_4207);
xor U4953 (N_4953,N_4393,N_4328);
and U4954 (N_4954,N_4140,N_4374);
nand U4955 (N_4955,N_4468,N_4218);
nand U4956 (N_4956,N_4181,N_4228);
and U4957 (N_4957,N_4246,N_4465);
nand U4958 (N_4958,N_4184,N_4288);
xor U4959 (N_4959,N_4017,N_4498);
and U4960 (N_4960,N_4489,N_4447);
xnor U4961 (N_4961,N_4414,N_4102);
nand U4962 (N_4962,N_4142,N_4073);
and U4963 (N_4963,N_4263,N_4040);
nor U4964 (N_4964,N_4494,N_4113);
and U4965 (N_4965,N_4496,N_4274);
xnor U4966 (N_4966,N_4214,N_4054);
xor U4967 (N_4967,N_4047,N_4393);
and U4968 (N_4968,N_4339,N_4480);
nand U4969 (N_4969,N_4340,N_4301);
or U4970 (N_4970,N_4026,N_4090);
and U4971 (N_4971,N_4197,N_4375);
nor U4972 (N_4972,N_4465,N_4219);
xor U4973 (N_4973,N_4328,N_4155);
nor U4974 (N_4974,N_4031,N_4291);
xnor U4975 (N_4975,N_4442,N_4491);
nor U4976 (N_4976,N_4263,N_4084);
or U4977 (N_4977,N_4133,N_4275);
xor U4978 (N_4978,N_4496,N_4225);
nor U4979 (N_4979,N_4422,N_4435);
nand U4980 (N_4980,N_4430,N_4036);
nor U4981 (N_4981,N_4297,N_4121);
xor U4982 (N_4982,N_4216,N_4236);
and U4983 (N_4983,N_4398,N_4064);
nand U4984 (N_4984,N_4361,N_4222);
xor U4985 (N_4985,N_4006,N_4307);
or U4986 (N_4986,N_4347,N_4121);
xnor U4987 (N_4987,N_4130,N_4434);
xor U4988 (N_4988,N_4457,N_4136);
or U4989 (N_4989,N_4258,N_4231);
xor U4990 (N_4990,N_4230,N_4040);
nor U4991 (N_4991,N_4385,N_4019);
or U4992 (N_4992,N_4495,N_4454);
or U4993 (N_4993,N_4344,N_4168);
xor U4994 (N_4994,N_4081,N_4431);
and U4995 (N_4995,N_4133,N_4189);
or U4996 (N_4996,N_4488,N_4090);
and U4997 (N_4997,N_4145,N_4015);
xnor U4998 (N_4998,N_4205,N_4337);
or U4999 (N_4999,N_4015,N_4233);
and U5000 (N_5000,N_4559,N_4790);
nor U5001 (N_5001,N_4900,N_4763);
nand U5002 (N_5002,N_4549,N_4817);
and U5003 (N_5003,N_4750,N_4862);
or U5004 (N_5004,N_4886,N_4820);
nor U5005 (N_5005,N_4717,N_4765);
nor U5006 (N_5006,N_4773,N_4595);
and U5007 (N_5007,N_4753,N_4636);
and U5008 (N_5008,N_4921,N_4913);
or U5009 (N_5009,N_4929,N_4819);
or U5010 (N_5010,N_4632,N_4940);
xor U5011 (N_5011,N_4836,N_4698);
or U5012 (N_5012,N_4527,N_4740);
and U5013 (N_5013,N_4749,N_4580);
or U5014 (N_5014,N_4708,N_4659);
xor U5015 (N_5015,N_4991,N_4537);
and U5016 (N_5016,N_4509,N_4788);
xor U5017 (N_5017,N_4898,N_4722);
nor U5018 (N_5018,N_4782,N_4506);
xnor U5019 (N_5019,N_4615,N_4744);
or U5020 (N_5020,N_4590,N_4955);
or U5021 (N_5021,N_4700,N_4910);
nor U5022 (N_5022,N_4508,N_4642);
nor U5023 (N_5023,N_4503,N_4643);
nor U5024 (N_5024,N_4973,N_4847);
nand U5025 (N_5025,N_4675,N_4604);
nor U5026 (N_5026,N_4649,N_4626);
or U5027 (N_5027,N_4568,N_4715);
or U5028 (N_5028,N_4769,N_4889);
nor U5029 (N_5029,N_4582,N_4644);
nand U5030 (N_5030,N_4860,N_4827);
nand U5031 (N_5031,N_4645,N_4752);
xor U5032 (N_5032,N_4767,N_4745);
or U5033 (N_5033,N_4545,N_4881);
and U5034 (N_5034,N_4528,N_4606);
or U5035 (N_5035,N_4883,N_4896);
and U5036 (N_5036,N_4637,N_4928);
xor U5037 (N_5037,N_4917,N_4760);
and U5038 (N_5038,N_4989,N_4920);
or U5039 (N_5039,N_4579,N_4899);
xnor U5040 (N_5040,N_4676,N_4914);
or U5041 (N_5041,N_4796,N_4625);
nor U5042 (N_5042,N_4840,N_4671);
nor U5043 (N_5043,N_4532,N_4747);
nand U5044 (N_5044,N_4791,N_4813);
or U5045 (N_5045,N_4842,N_4657);
xnor U5046 (N_5046,N_4775,N_4570);
nand U5047 (N_5047,N_4967,N_4833);
or U5048 (N_5048,N_4610,N_4622);
nand U5049 (N_5049,N_4500,N_4895);
nor U5050 (N_5050,N_4810,N_4678);
xnor U5051 (N_5051,N_4866,N_4964);
nand U5052 (N_5052,N_4739,N_4864);
xor U5053 (N_5053,N_4779,N_4507);
xnor U5054 (N_5054,N_4607,N_4903);
nand U5055 (N_5055,N_4547,N_4924);
nand U5056 (N_5056,N_4660,N_4858);
and U5057 (N_5057,N_4541,N_4669);
or U5058 (N_5058,N_4902,N_4670);
or U5059 (N_5059,N_4618,N_4523);
xor U5060 (N_5060,N_4915,N_4834);
nor U5061 (N_5061,N_4647,N_4719);
or U5062 (N_5062,N_4540,N_4832);
nand U5063 (N_5063,N_4727,N_4963);
or U5064 (N_5064,N_4887,N_4987);
and U5065 (N_5065,N_4846,N_4777);
and U5066 (N_5066,N_4873,N_4728);
nand U5067 (N_5067,N_4706,N_4758);
and U5068 (N_5068,N_4733,N_4783);
xnor U5069 (N_5069,N_4677,N_4894);
nor U5070 (N_5070,N_4529,N_4923);
nor U5071 (N_5071,N_4612,N_4795);
nand U5072 (N_5072,N_4705,N_4623);
and U5073 (N_5073,N_4861,N_4982);
nand U5074 (N_5074,N_4553,N_4720);
nand U5075 (N_5075,N_4950,N_4613);
or U5076 (N_5076,N_4845,N_4619);
and U5077 (N_5077,N_4598,N_4871);
or U5078 (N_5078,N_4919,N_4609);
or U5079 (N_5079,N_4661,N_4682);
nor U5080 (N_5080,N_4550,N_4966);
xnor U5081 (N_5081,N_4614,N_4511);
and U5082 (N_5082,N_4904,N_4837);
nor U5083 (N_5083,N_4811,N_4936);
and U5084 (N_5084,N_4759,N_4555);
or U5085 (N_5085,N_4948,N_4748);
and U5086 (N_5086,N_4780,N_4674);
nand U5087 (N_5087,N_4852,N_4631);
nor U5088 (N_5088,N_4673,N_4692);
or U5089 (N_5089,N_4627,N_4712);
nand U5090 (N_5090,N_4875,N_4854);
and U5091 (N_5091,N_4867,N_4986);
nand U5092 (N_5092,N_4792,N_4907);
or U5093 (N_5093,N_4561,N_4960);
nor U5094 (N_5094,N_4856,N_4865);
and U5095 (N_5095,N_4571,N_4514);
nand U5096 (N_5096,N_4971,N_4602);
nor U5097 (N_5097,N_4818,N_4738);
xnor U5098 (N_5098,N_4761,N_4906);
nand U5099 (N_5099,N_4957,N_4958);
and U5100 (N_5100,N_4892,N_4962);
nand U5101 (N_5101,N_4799,N_4648);
xor U5102 (N_5102,N_4774,N_4624);
or U5103 (N_5103,N_4513,N_4668);
nor U5104 (N_5104,N_4735,N_4869);
xor U5105 (N_5105,N_4821,N_4686);
or U5106 (N_5106,N_4901,N_4713);
or U5107 (N_5107,N_4594,N_4781);
or U5108 (N_5108,N_4600,N_4583);
and U5109 (N_5109,N_4880,N_4651);
or U5110 (N_5110,N_4517,N_4567);
or U5111 (N_5111,N_4605,N_4656);
xor U5112 (N_5112,N_4542,N_4650);
xor U5113 (N_5113,N_4951,N_4578);
xor U5114 (N_5114,N_4998,N_4634);
and U5115 (N_5115,N_4938,N_4592);
nor U5116 (N_5116,N_4538,N_4793);
nor U5117 (N_5117,N_4990,N_4731);
or U5118 (N_5118,N_4853,N_4638);
nand U5119 (N_5119,N_4771,N_4979);
and U5120 (N_5120,N_4839,N_4888);
and U5121 (N_5121,N_4680,N_4672);
xor U5122 (N_5122,N_4726,N_4601);
nor U5123 (N_5123,N_4653,N_4701);
nor U5124 (N_5124,N_4943,N_4874);
or U5125 (N_5125,N_4803,N_4911);
and U5126 (N_5126,N_4710,N_4746);
and U5127 (N_5127,N_4596,N_4522);
and U5128 (N_5128,N_4597,N_4518);
xor U5129 (N_5129,N_4806,N_4737);
or U5130 (N_5130,N_4654,N_4932);
or U5131 (N_5131,N_4718,N_4812);
xor U5132 (N_5132,N_4961,N_4972);
nor U5133 (N_5133,N_4665,N_4893);
and U5134 (N_5134,N_4617,N_4693);
or U5135 (N_5135,N_4611,N_4997);
xnor U5136 (N_5136,N_4877,N_4531);
nand U5137 (N_5137,N_4694,N_4732);
nor U5138 (N_5138,N_4663,N_4729);
and U5139 (N_5139,N_4699,N_4723);
nor U5140 (N_5140,N_4848,N_4976);
or U5141 (N_5141,N_4849,N_4558);
or U5142 (N_5142,N_4794,N_4530);
or U5143 (N_5143,N_4863,N_4784);
nor U5144 (N_5144,N_4563,N_4786);
nand U5145 (N_5145,N_4802,N_4996);
and U5146 (N_5146,N_4640,N_4879);
xor U5147 (N_5147,N_4515,N_4776);
or U5148 (N_5148,N_4945,N_4741);
nor U5149 (N_5149,N_4985,N_4838);
nor U5150 (N_5150,N_4709,N_4743);
or U5151 (N_5151,N_4825,N_4721);
or U5152 (N_5152,N_4516,N_4603);
and U5153 (N_5153,N_4933,N_4939);
and U5154 (N_5154,N_4608,N_4574);
or U5155 (N_5155,N_4683,N_4897);
nand U5156 (N_5156,N_4978,N_4655);
xnor U5157 (N_5157,N_4981,N_4843);
or U5158 (N_5158,N_4687,N_4857);
nor U5159 (N_5159,N_4844,N_4725);
nand U5160 (N_5160,N_4912,N_4808);
nand U5161 (N_5161,N_4593,N_4512);
or U5162 (N_5162,N_4918,N_4556);
xnor U5163 (N_5163,N_4539,N_4931);
or U5164 (N_5164,N_4646,N_4535);
or U5165 (N_5165,N_4789,N_4804);
and U5166 (N_5166,N_4543,N_4526);
and U5167 (N_5167,N_4942,N_4787);
or U5168 (N_5168,N_4551,N_4946);
xor U5169 (N_5169,N_4850,N_4711);
nand U5170 (N_5170,N_4505,N_4975);
or U5171 (N_5171,N_4520,N_4934);
nand U5172 (N_5172,N_4628,N_4702);
xor U5173 (N_5173,N_4641,N_4560);
xnor U5174 (N_5174,N_4952,N_4956);
xnor U5175 (N_5175,N_4968,N_4587);
nor U5176 (N_5176,N_4635,N_4691);
nand U5177 (N_5177,N_4965,N_4800);
nor U5178 (N_5178,N_4916,N_4616);
or U5179 (N_5179,N_4681,N_4754);
xnor U5180 (N_5180,N_4935,N_4974);
xnor U5181 (N_5181,N_4766,N_4954);
xnor U5182 (N_5182,N_4872,N_4855);
nand U5183 (N_5183,N_4891,N_4851);
nor U5184 (N_5184,N_4992,N_4562);
nor U5185 (N_5185,N_4772,N_4707);
nor U5186 (N_5186,N_4629,N_4947);
xor U5187 (N_5187,N_4521,N_4519);
and U5188 (N_5188,N_4984,N_4764);
and U5189 (N_5189,N_4565,N_4566);
nand U5190 (N_5190,N_4977,N_4824);
and U5191 (N_5191,N_4770,N_4585);
xnor U5192 (N_5192,N_4575,N_4930);
nand U5193 (N_5193,N_4652,N_4878);
or U5194 (N_5194,N_4502,N_4639);
xnor U5195 (N_5195,N_4621,N_4664);
and U5196 (N_5196,N_4548,N_4905);
xor U5197 (N_5197,N_4801,N_4988);
and U5198 (N_5198,N_4533,N_4809);
and U5199 (N_5199,N_4969,N_4742);
nor U5200 (N_5200,N_4949,N_4830);
or U5201 (N_5201,N_4785,N_4696);
nand U5202 (N_5202,N_4983,N_4501);
or U5203 (N_5203,N_4994,N_4884);
nor U5204 (N_5204,N_4666,N_4730);
nor U5205 (N_5205,N_4734,N_4584);
xor U5206 (N_5206,N_4885,N_4546);
nand U5207 (N_5207,N_4630,N_4536);
nor U5208 (N_5208,N_4633,N_4822);
nor U5209 (N_5209,N_4510,N_4577);
or U5210 (N_5210,N_4525,N_4980);
xor U5211 (N_5211,N_4581,N_4882);
and U5212 (N_5212,N_4870,N_4589);
or U5213 (N_5213,N_4755,N_4757);
nor U5214 (N_5214,N_4925,N_4534);
or U5215 (N_5215,N_4922,N_4953);
nand U5216 (N_5216,N_4684,N_4591);
or U5217 (N_5217,N_4576,N_4564);
or U5218 (N_5218,N_4814,N_4805);
and U5219 (N_5219,N_4679,N_4995);
xor U5220 (N_5220,N_4937,N_4724);
or U5221 (N_5221,N_4797,N_4552);
and U5222 (N_5222,N_4890,N_4970);
and U5223 (N_5223,N_4544,N_4662);
nand U5224 (N_5224,N_4999,N_4572);
xor U5225 (N_5225,N_4714,N_4751);
nand U5226 (N_5226,N_4815,N_4756);
or U5227 (N_5227,N_4959,N_4944);
or U5228 (N_5228,N_4826,N_4689);
and U5229 (N_5229,N_4835,N_4716);
nor U5230 (N_5230,N_4690,N_4504);
nand U5231 (N_5231,N_4941,N_4778);
and U5232 (N_5232,N_4697,N_4569);
or U5233 (N_5233,N_4688,N_4859);
and U5234 (N_5234,N_4828,N_4736);
and U5235 (N_5235,N_4762,N_4807);
xnor U5236 (N_5236,N_4831,N_4667);
or U5237 (N_5237,N_4841,N_4993);
xnor U5238 (N_5238,N_4703,N_4620);
nand U5239 (N_5239,N_4876,N_4816);
xnor U5240 (N_5240,N_4658,N_4768);
xor U5241 (N_5241,N_4557,N_4524);
or U5242 (N_5242,N_4685,N_4704);
and U5243 (N_5243,N_4927,N_4909);
nand U5244 (N_5244,N_4823,N_4554);
and U5245 (N_5245,N_4868,N_4926);
xor U5246 (N_5246,N_4695,N_4829);
xnor U5247 (N_5247,N_4586,N_4588);
nand U5248 (N_5248,N_4908,N_4599);
and U5249 (N_5249,N_4798,N_4573);
nor U5250 (N_5250,N_4567,N_4844);
nand U5251 (N_5251,N_4985,N_4955);
nand U5252 (N_5252,N_4794,N_4821);
or U5253 (N_5253,N_4990,N_4650);
xor U5254 (N_5254,N_4992,N_4863);
or U5255 (N_5255,N_4690,N_4845);
xnor U5256 (N_5256,N_4848,N_4739);
nand U5257 (N_5257,N_4840,N_4611);
or U5258 (N_5258,N_4882,N_4906);
nor U5259 (N_5259,N_4733,N_4862);
or U5260 (N_5260,N_4940,N_4742);
nor U5261 (N_5261,N_4548,N_4981);
xnor U5262 (N_5262,N_4770,N_4703);
xor U5263 (N_5263,N_4724,N_4528);
xor U5264 (N_5264,N_4856,N_4530);
nor U5265 (N_5265,N_4532,N_4599);
or U5266 (N_5266,N_4570,N_4969);
nor U5267 (N_5267,N_4601,N_4503);
nor U5268 (N_5268,N_4940,N_4993);
and U5269 (N_5269,N_4803,N_4951);
and U5270 (N_5270,N_4969,N_4582);
nor U5271 (N_5271,N_4579,N_4872);
xor U5272 (N_5272,N_4898,N_4573);
nor U5273 (N_5273,N_4681,N_4730);
nand U5274 (N_5274,N_4905,N_4809);
nor U5275 (N_5275,N_4898,N_4864);
and U5276 (N_5276,N_4978,N_4749);
nor U5277 (N_5277,N_4732,N_4597);
or U5278 (N_5278,N_4886,N_4589);
and U5279 (N_5279,N_4635,N_4846);
and U5280 (N_5280,N_4957,N_4654);
or U5281 (N_5281,N_4751,N_4788);
xnor U5282 (N_5282,N_4547,N_4549);
or U5283 (N_5283,N_4714,N_4669);
and U5284 (N_5284,N_4733,N_4889);
nor U5285 (N_5285,N_4665,N_4542);
or U5286 (N_5286,N_4505,N_4892);
nor U5287 (N_5287,N_4768,N_4596);
nor U5288 (N_5288,N_4644,N_4872);
xnor U5289 (N_5289,N_4592,N_4957);
xor U5290 (N_5290,N_4974,N_4918);
nand U5291 (N_5291,N_4855,N_4920);
and U5292 (N_5292,N_4775,N_4589);
nor U5293 (N_5293,N_4562,N_4647);
nor U5294 (N_5294,N_4682,N_4698);
and U5295 (N_5295,N_4882,N_4515);
xnor U5296 (N_5296,N_4517,N_4768);
xor U5297 (N_5297,N_4543,N_4975);
and U5298 (N_5298,N_4600,N_4925);
or U5299 (N_5299,N_4815,N_4553);
xor U5300 (N_5300,N_4794,N_4993);
nor U5301 (N_5301,N_4700,N_4541);
and U5302 (N_5302,N_4612,N_4669);
nor U5303 (N_5303,N_4768,N_4776);
nand U5304 (N_5304,N_4691,N_4555);
nand U5305 (N_5305,N_4518,N_4619);
and U5306 (N_5306,N_4795,N_4595);
or U5307 (N_5307,N_4532,N_4896);
nand U5308 (N_5308,N_4528,N_4943);
nor U5309 (N_5309,N_4684,N_4998);
nor U5310 (N_5310,N_4599,N_4922);
nand U5311 (N_5311,N_4570,N_4679);
nand U5312 (N_5312,N_4876,N_4520);
xor U5313 (N_5313,N_4902,N_4983);
or U5314 (N_5314,N_4627,N_4937);
xnor U5315 (N_5315,N_4861,N_4780);
xnor U5316 (N_5316,N_4917,N_4912);
nor U5317 (N_5317,N_4742,N_4597);
or U5318 (N_5318,N_4764,N_4876);
nand U5319 (N_5319,N_4985,N_4630);
nor U5320 (N_5320,N_4699,N_4858);
xor U5321 (N_5321,N_4509,N_4999);
xor U5322 (N_5322,N_4592,N_4634);
or U5323 (N_5323,N_4541,N_4920);
or U5324 (N_5324,N_4935,N_4581);
nand U5325 (N_5325,N_4998,N_4502);
xnor U5326 (N_5326,N_4566,N_4641);
xor U5327 (N_5327,N_4996,N_4606);
and U5328 (N_5328,N_4803,N_4960);
or U5329 (N_5329,N_4672,N_4546);
xnor U5330 (N_5330,N_4879,N_4772);
or U5331 (N_5331,N_4552,N_4915);
nand U5332 (N_5332,N_4879,N_4877);
xnor U5333 (N_5333,N_4719,N_4661);
and U5334 (N_5334,N_4535,N_4558);
and U5335 (N_5335,N_4655,N_4941);
nor U5336 (N_5336,N_4856,N_4521);
or U5337 (N_5337,N_4693,N_4886);
xor U5338 (N_5338,N_4811,N_4560);
nand U5339 (N_5339,N_4610,N_4963);
and U5340 (N_5340,N_4858,N_4860);
and U5341 (N_5341,N_4948,N_4818);
xnor U5342 (N_5342,N_4993,N_4578);
xor U5343 (N_5343,N_4593,N_4996);
nor U5344 (N_5344,N_4943,N_4844);
nand U5345 (N_5345,N_4815,N_4863);
or U5346 (N_5346,N_4665,N_4990);
and U5347 (N_5347,N_4584,N_4748);
and U5348 (N_5348,N_4941,N_4806);
nor U5349 (N_5349,N_4782,N_4614);
xnor U5350 (N_5350,N_4613,N_4933);
and U5351 (N_5351,N_4593,N_4829);
xor U5352 (N_5352,N_4567,N_4959);
or U5353 (N_5353,N_4593,N_4680);
nand U5354 (N_5354,N_4880,N_4524);
nand U5355 (N_5355,N_4936,N_4652);
nor U5356 (N_5356,N_4680,N_4562);
or U5357 (N_5357,N_4655,N_4885);
nor U5358 (N_5358,N_4858,N_4822);
and U5359 (N_5359,N_4864,N_4809);
nand U5360 (N_5360,N_4979,N_4878);
and U5361 (N_5361,N_4615,N_4966);
and U5362 (N_5362,N_4898,N_4688);
xnor U5363 (N_5363,N_4736,N_4752);
or U5364 (N_5364,N_4598,N_4511);
and U5365 (N_5365,N_4872,N_4817);
and U5366 (N_5366,N_4934,N_4547);
nand U5367 (N_5367,N_4751,N_4505);
nand U5368 (N_5368,N_4891,N_4932);
nor U5369 (N_5369,N_4513,N_4585);
xnor U5370 (N_5370,N_4927,N_4570);
xnor U5371 (N_5371,N_4858,N_4730);
nand U5372 (N_5372,N_4738,N_4929);
and U5373 (N_5373,N_4522,N_4905);
and U5374 (N_5374,N_4691,N_4610);
nand U5375 (N_5375,N_4849,N_4715);
nand U5376 (N_5376,N_4810,N_4515);
nand U5377 (N_5377,N_4839,N_4891);
xor U5378 (N_5378,N_4828,N_4811);
or U5379 (N_5379,N_4685,N_4654);
or U5380 (N_5380,N_4514,N_4970);
nor U5381 (N_5381,N_4785,N_4743);
nand U5382 (N_5382,N_4660,N_4671);
nand U5383 (N_5383,N_4517,N_4722);
xnor U5384 (N_5384,N_4872,N_4958);
xor U5385 (N_5385,N_4681,N_4580);
nand U5386 (N_5386,N_4585,N_4540);
nand U5387 (N_5387,N_4952,N_4796);
and U5388 (N_5388,N_4716,N_4713);
and U5389 (N_5389,N_4899,N_4948);
or U5390 (N_5390,N_4704,N_4925);
or U5391 (N_5391,N_4859,N_4594);
or U5392 (N_5392,N_4925,N_4920);
and U5393 (N_5393,N_4638,N_4747);
or U5394 (N_5394,N_4703,N_4951);
xor U5395 (N_5395,N_4641,N_4777);
nor U5396 (N_5396,N_4684,N_4649);
xor U5397 (N_5397,N_4603,N_4756);
and U5398 (N_5398,N_4839,N_4613);
nand U5399 (N_5399,N_4570,N_4852);
nand U5400 (N_5400,N_4731,N_4796);
or U5401 (N_5401,N_4590,N_4750);
xor U5402 (N_5402,N_4938,N_4969);
or U5403 (N_5403,N_4523,N_4616);
xnor U5404 (N_5404,N_4692,N_4691);
xor U5405 (N_5405,N_4890,N_4569);
xnor U5406 (N_5406,N_4917,N_4741);
or U5407 (N_5407,N_4569,N_4688);
nor U5408 (N_5408,N_4693,N_4677);
nand U5409 (N_5409,N_4671,N_4685);
xnor U5410 (N_5410,N_4879,N_4517);
xnor U5411 (N_5411,N_4873,N_4511);
xor U5412 (N_5412,N_4809,N_4675);
nand U5413 (N_5413,N_4924,N_4847);
nand U5414 (N_5414,N_4790,N_4932);
nand U5415 (N_5415,N_4556,N_4514);
and U5416 (N_5416,N_4807,N_4811);
nand U5417 (N_5417,N_4839,N_4571);
and U5418 (N_5418,N_4926,N_4812);
or U5419 (N_5419,N_4543,N_4705);
or U5420 (N_5420,N_4536,N_4705);
and U5421 (N_5421,N_4971,N_4686);
nand U5422 (N_5422,N_4950,N_4697);
or U5423 (N_5423,N_4990,N_4645);
nor U5424 (N_5424,N_4510,N_4742);
or U5425 (N_5425,N_4972,N_4674);
or U5426 (N_5426,N_4530,N_4595);
and U5427 (N_5427,N_4649,N_4777);
or U5428 (N_5428,N_4841,N_4614);
or U5429 (N_5429,N_4659,N_4694);
nand U5430 (N_5430,N_4974,N_4568);
nand U5431 (N_5431,N_4727,N_4742);
or U5432 (N_5432,N_4571,N_4610);
nor U5433 (N_5433,N_4611,N_4534);
xnor U5434 (N_5434,N_4931,N_4966);
xnor U5435 (N_5435,N_4987,N_4698);
or U5436 (N_5436,N_4712,N_4674);
or U5437 (N_5437,N_4625,N_4526);
and U5438 (N_5438,N_4819,N_4716);
nor U5439 (N_5439,N_4740,N_4855);
xnor U5440 (N_5440,N_4585,N_4978);
or U5441 (N_5441,N_4944,N_4618);
or U5442 (N_5442,N_4757,N_4750);
or U5443 (N_5443,N_4708,N_4917);
nand U5444 (N_5444,N_4876,N_4812);
and U5445 (N_5445,N_4945,N_4513);
xor U5446 (N_5446,N_4777,N_4686);
nand U5447 (N_5447,N_4820,N_4784);
or U5448 (N_5448,N_4728,N_4982);
or U5449 (N_5449,N_4786,N_4581);
nand U5450 (N_5450,N_4587,N_4815);
and U5451 (N_5451,N_4822,N_4790);
nand U5452 (N_5452,N_4536,N_4718);
xnor U5453 (N_5453,N_4726,N_4675);
xnor U5454 (N_5454,N_4935,N_4882);
or U5455 (N_5455,N_4599,N_4802);
or U5456 (N_5456,N_4600,N_4684);
or U5457 (N_5457,N_4798,N_4847);
nand U5458 (N_5458,N_4534,N_4911);
xor U5459 (N_5459,N_4786,N_4748);
xnor U5460 (N_5460,N_4989,N_4908);
and U5461 (N_5461,N_4660,N_4623);
or U5462 (N_5462,N_4728,N_4824);
or U5463 (N_5463,N_4760,N_4803);
nand U5464 (N_5464,N_4940,N_4680);
xnor U5465 (N_5465,N_4912,N_4892);
and U5466 (N_5466,N_4552,N_4870);
or U5467 (N_5467,N_4691,N_4505);
nor U5468 (N_5468,N_4645,N_4670);
nand U5469 (N_5469,N_4689,N_4949);
xnor U5470 (N_5470,N_4853,N_4867);
or U5471 (N_5471,N_4716,N_4540);
xnor U5472 (N_5472,N_4859,N_4623);
nand U5473 (N_5473,N_4634,N_4923);
or U5474 (N_5474,N_4634,N_4551);
and U5475 (N_5475,N_4673,N_4925);
or U5476 (N_5476,N_4669,N_4967);
and U5477 (N_5477,N_4761,N_4856);
xor U5478 (N_5478,N_4722,N_4602);
nor U5479 (N_5479,N_4537,N_4653);
or U5480 (N_5480,N_4715,N_4825);
nor U5481 (N_5481,N_4913,N_4780);
nor U5482 (N_5482,N_4705,N_4563);
nand U5483 (N_5483,N_4668,N_4643);
xor U5484 (N_5484,N_4615,N_4753);
nor U5485 (N_5485,N_4892,N_4934);
nand U5486 (N_5486,N_4605,N_4942);
xor U5487 (N_5487,N_4690,N_4689);
and U5488 (N_5488,N_4722,N_4663);
nand U5489 (N_5489,N_4659,N_4638);
nor U5490 (N_5490,N_4758,N_4934);
nand U5491 (N_5491,N_4627,N_4912);
nor U5492 (N_5492,N_4944,N_4811);
nor U5493 (N_5493,N_4768,N_4993);
and U5494 (N_5494,N_4936,N_4921);
and U5495 (N_5495,N_4789,N_4916);
nand U5496 (N_5496,N_4596,N_4713);
nand U5497 (N_5497,N_4569,N_4766);
nand U5498 (N_5498,N_4653,N_4924);
nand U5499 (N_5499,N_4931,N_4719);
nor U5500 (N_5500,N_5318,N_5109);
and U5501 (N_5501,N_5315,N_5173);
or U5502 (N_5502,N_5160,N_5395);
and U5503 (N_5503,N_5489,N_5473);
or U5504 (N_5504,N_5348,N_5198);
or U5505 (N_5505,N_5096,N_5210);
and U5506 (N_5506,N_5457,N_5108);
and U5507 (N_5507,N_5064,N_5036);
and U5508 (N_5508,N_5446,N_5261);
xor U5509 (N_5509,N_5305,N_5155);
or U5510 (N_5510,N_5434,N_5491);
xor U5511 (N_5511,N_5167,N_5450);
nor U5512 (N_5512,N_5307,N_5146);
or U5513 (N_5513,N_5381,N_5005);
nand U5514 (N_5514,N_5007,N_5361);
or U5515 (N_5515,N_5199,N_5245);
nor U5516 (N_5516,N_5394,N_5497);
nand U5517 (N_5517,N_5372,N_5006);
and U5518 (N_5518,N_5013,N_5015);
or U5519 (N_5519,N_5073,N_5387);
nor U5520 (N_5520,N_5045,N_5367);
and U5521 (N_5521,N_5057,N_5465);
and U5522 (N_5522,N_5162,N_5448);
or U5523 (N_5523,N_5113,N_5299);
and U5524 (N_5524,N_5243,N_5257);
or U5525 (N_5525,N_5140,N_5370);
or U5526 (N_5526,N_5084,N_5055);
and U5527 (N_5527,N_5314,N_5070);
and U5528 (N_5528,N_5355,N_5079);
nor U5529 (N_5529,N_5075,N_5402);
nor U5530 (N_5530,N_5228,N_5260);
nor U5531 (N_5531,N_5266,N_5408);
and U5532 (N_5532,N_5470,N_5241);
xor U5533 (N_5533,N_5046,N_5293);
and U5534 (N_5534,N_5360,N_5253);
or U5535 (N_5535,N_5347,N_5327);
nand U5536 (N_5536,N_5111,N_5127);
and U5537 (N_5537,N_5164,N_5191);
and U5538 (N_5538,N_5175,N_5100);
or U5539 (N_5539,N_5004,N_5330);
and U5540 (N_5540,N_5214,N_5068);
and U5541 (N_5541,N_5296,N_5066);
nor U5542 (N_5542,N_5389,N_5422);
and U5543 (N_5543,N_5376,N_5391);
xnor U5544 (N_5544,N_5051,N_5308);
nor U5545 (N_5545,N_5209,N_5067);
and U5546 (N_5546,N_5291,N_5374);
and U5547 (N_5547,N_5365,N_5223);
nor U5548 (N_5548,N_5440,N_5144);
and U5549 (N_5549,N_5282,N_5125);
and U5550 (N_5550,N_5041,N_5375);
and U5551 (N_5551,N_5346,N_5369);
nand U5552 (N_5552,N_5479,N_5499);
and U5553 (N_5553,N_5044,N_5280);
and U5554 (N_5554,N_5474,N_5487);
or U5555 (N_5555,N_5224,N_5244);
nor U5556 (N_5556,N_5435,N_5317);
xnor U5557 (N_5557,N_5380,N_5432);
xnor U5558 (N_5558,N_5195,N_5252);
or U5559 (N_5559,N_5377,N_5212);
xnor U5560 (N_5560,N_5178,N_5285);
xor U5561 (N_5561,N_5269,N_5093);
nand U5562 (N_5562,N_5256,N_5115);
xor U5563 (N_5563,N_5171,N_5414);
and U5564 (N_5564,N_5398,N_5083);
nor U5565 (N_5565,N_5400,N_5258);
and U5566 (N_5566,N_5443,N_5119);
nand U5567 (N_5567,N_5233,N_5095);
and U5568 (N_5568,N_5149,N_5021);
nor U5569 (N_5569,N_5238,N_5011);
xor U5570 (N_5570,N_5213,N_5039);
and U5571 (N_5571,N_5366,N_5251);
or U5572 (N_5572,N_5081,N_5118);
and U5573 (N_5573,N_5439,N_5458);
nand U5574 (N_5574,N_5193,N_5215);
or U5575 (N_5575,N_5186,N_5284);
nor U5576 (N_5576,N_5419,N_5472);
xor U5577 (N_5577,N_5185,N_5000);
xnor U5578 (N_5578,N_5102,N_5122);
nor U5579 (N_5579,N_5010,N_5271);
nor U5580 (N_5580,N_5025,N_5071);
and U5581 (N_5581,N_5183,N_5493);
nand U5582 (N_5582,N_5478,N_5364);
and U5583 (N_5583,N_5147,N_5231);
or U5584 (N_5584,N_5054,N_5342);
nand U5585 (N_5585,N_5056,N_5080);
xnor U5586 (N_5586,N_5311,N_5328);
nor U5587 (N_5587,N_5386,N_5012);
nand U5588 (N_5588,N_5325,N_5496);
or U5589 (N_5589,N_5246,N_5301);
or U5590 (N_5590,N_5161,N_5272);
or U5591 (N_5591,N_5456,N_5129);
and U5592 (N_5592,N_5468,N_5047);
and U5593 (N_5593,N_5123,N_5292);
or U5594 (N_5594,N_5481,N_5034);
or U5595 (N_5595,N_5403,N_5385);
xnor U5596 (N_5596,N_5249,N_5437);
and U5597 (N_5597,N_5156,N_5431);
and U5598 (N_5598,N_5485,N_5321);
xor U5599 (N_5599,N_5262,N_5480);
and U5600 (N_5600,N_5237,N_5275);
or U5601 (N_5601,N_5154,N_5225);
and U5602 (N_5602,N_5462,N_5059);
nand U5603 (N_5603,N_5410,N_5356);
or U5604 (N_5604,N_5232,N_5274);
nor U5605 (N_5605,N_5104,N_5494);
nand U5606 (N_5606,N_5357,N_5428);
nand U5607 (N_5607,N_5211,N_5363);
nand U5608 (N_5608,N_5368,N_5290);
or U5609 (N_5609,N_5433,N_5124);
nand U5610 (N_5610,N_5131,N_5240);
xor U5611 (N_5611,N_5338,N_5078);
or U5612 (N_5612,N_5018,N_5168);
nand U5613 (N_5613,N_5393,N_5416);
nor U5614 (N_5614,N_5032,N_5189);
xnor U5615 (N_5615,N_5302,N_5312);
and U5616 (N_5616,N_5340,N_5294);
nor U5617 (N_5617,N_5201,N_5184);
xor U5618 (N_5618,N_5441,N_5415);
nor U5619 (N_5619,N_5339,N_5017);
xnor U5620 (N_5620,N_5390,N_5316);
nand U5621 (N_5621,N_5172,N_5498);
xor U5622 (N_5622,N_5138,N_5306);
nand U5623 (N_5623,N_5424,N_5062);
nor U5624 (N_5624,N_5061,N_5300);
or U5625 (N_5625,N_5313,N_5076);
xor U5626 (N_5626,N_5409,N_5087);
nand U5627 (N_5627,N_5336,N_5278);
nor U5628 (N_5628,N_5188,N_5023);
xor U5629 (N_5629,N_5074,N_5341);
nor U5630 (N_5630,N_5002,N_5333);
or U5631 (N_5631,N_5203,N_5418);
nand U5632 (N_5632,N_5382,N_5235);
nand U5633 (N_5633,N_5334,N_5157);
nor U5634 (N_5634,N_5326,N_5159);
and U5635 (N_5635,N_5177,N_5412);
and U5636 (N_5636,N_5452,N_5362);
nand U5637 (N_5637,N_5350,N_5106);
nand U5638 (N_5638,N_5137,N_5298);
and U5639 (N_5639,N_5098,N_5353);
or U5640 (N_5640,N_5090,N_5322);
xnor U5641 (N_5641,N_5222,N_5247);
nor U5642 (N_5642,N_5145,N_5092);
and U5643 (N_5643,N_5024,N_5219);
nand U5644 (N_5644,N_5218,N_5482);
xnor U5645 (N_5645,N_5273,N_5085);
nor U5646 (N_5646,N_5009,N_5063);
nor U5647 (N_5647,N_5058,N_5270);
and U5648 (N_5648,N_5351,N_5229);
xnor U5649 (N_5649,N_5417,N_5304);
or U5650 (N_5650,N_5152,N_5451);
xnor U5651 (N_5651,N_5476,N_5181);
or U5652 (N_5652,N_5279,N_5148);
nor U5653 (N_5653,N_5069,N_5319);
or U5654 (N_5654,N_5128,N_5254);
nand U5655 (N_5655,N_5220,N_5028);
nand U5656 (N_5656,N_5411,N_5495);
and U5657 (N_5657,N_5116,N_5475);
nor U5658 (N_5658,N_5107,N_5259);
or U5659 (N_5659,N_5197,N_5421);
nor U5660 (N_5660,N_5423,N_5255);
xor U5661 (N_5661,N_5329,N_5179);
or U5662 (N_5662,N_5141,N_5099);
and U5663 (N_5663,N_5460,N_5471);
and U5664 (N_5664,N_5158,N_5442);
nor U5665 (N_5665,N_5163,N_5035);
xor U5666 (N_5666,N_5429,N_5425);
or U5667 (N_5667,N_5042,N_5407);
xnor U5668 (N_5668,N_5345,N_5287);
nand U5669 (N_5669,N_5072,N_5038);
xor U5670 (N_5670,N_5089,N_5276);
nand U5671 (N_5671,N_5033,N_5444);
nand U5672 (N_5672,N_5052,N_5192);
nor U5673 (N_5673,N_5404,N_5295);
or U5674 (N_5674,N_5281,N_5453);
xor U5675 (N_5675,N_5121,N_5239);
and U5676 (N_5676,N_5050,N_5112);
nand U5677 (N_5677,N_5088,N_5170);
and U5678 (N_5678,N_5413,N_5135);
nor U5679 (N_5679,N_5320,N_5323);
and U5680 (N_5680,N_5268,N_5484);
or U5681 (N_5681,N_5030,N_5001);
nor U5682 (N_5682,N_5477,N_5016);
nor U5683 (N_5683,N_5397,N_5142);
xor U5684 (N_5684,N_5343,N_5399);
nor U5685 (N_5685,N_5031,N_5008);
and U5686 (N_5686,N_5267,N_5082);
nor U5687 (N_5687,N_5026,N_5406);
nand U5688 (N_5688,N_5277,N_5352);
nand U5689 (N_5689,N_5027,N_5483);
xnor U5690 (N_5690,N_5150,N_5205);
and U5691 (N_5691,N_5176,N_5234);
and U5692 (N_5692,N_5335,N_5396);
nor U5693 (N_5693,N_5060,N_5447);
xnor U5694 (N_5694,N_5126,N_5392);
xnor U5695 (N_5695,N_5182,N_5003);
nor U5696 (N_5696,N_5194,N_5488);
xor U5697 (N_5697,N_5384,N_5469);
or U5698 (N_5698,N_5286,N_5166);
nand U5699 (N_5699,N_5371,N_5133);
and U5700 (N_5700,N_5200,N_5297);
nand U5701 (N_5701,N_5130,N_5101);
nor U5702 (N_5702,N_5226,N_5303);
nand U5703 (N_5703,N_5065,N_5486);
and U5704 (N_5704,N_5454,N_5337);
nand U5705 (N_5705,N_5180,N_5077);
xnor U5706 (N_5706,N_5204,N_5086);
or U5707 (N_5707,N_5029,N_5132);
or U5708 (N_5708,N_5105,N_5037);
xor U5709 (N_5709,N_5221,N_5464);
or U5710 (N_5710,N_5436,N_5236);
and U5711 (N_5711,N_5227,N_5378);
xor U5712 (N_5712,N_5459,N_5331);
or U5713 (N_5713,N_5383,N_5165);
or U5714 (N_5714,N_5427,N_5216);
or U5715 (N_5715,N_5139,N_5354);
or U5716 (N_5716,N_5208,N_5401);
or U5717 (N_5717,N_5053,N_5187);
and U5718 (N_5718,N_5388,N_5094);
nor U5719 (N_5719,N_5445,N_5289);
nand U5720 (N_5720,N_5438,N_5430);
or U5721 (N_5721,N_5169,N_5020);
or U5722 (N_5722,N_5202,N_5190);
and U5723 (N_5723,N_5151,N_5206);
nand U5724 (N_5724,N_5091,N_5120);
nor U5725 (N_5725,N_5019,N_5426);
nor U5726 (N_5726,N_5373,N_5490);
xnor U5727 (N_5727,N_5461,N_5349);
nor U5728 (N_5728,N_5040,N_5359);
or U5729 (N_5729,N_5463,N_5455);
xnor U5730 (N_5730,N_5136,N_5310);
or U5731 (N_5731,N_5022,N_5114);
nor U5732 (N_5732,N_5492,N_5049);
nand U5733 (N_5733,N_5324,N_5309);
xnor U5734 (N_5734,N_5358,N_5143);
or U5735 (N_5735,N_5153,N_5117);
nand U5736 (N_5736,N_5230,N_5014);
xor U5737 (N_5737,N_5097,N_5420);
nand U5738 (N_5738,N_5265,N_5344);
and U5739 (N_5739,N_5110,N_5048);
or U5740 (N_5740,N_5134,N_5288);
or U5741 (N_5741,N_5248,N_5207);
xor U5742 (N_5742,N_5217,N_5242);
or U5743 (N_5743,N_5263,N_5103);
xnor U5744 (N_5744,N_5449,N_5405);
xor U5745 (N_5745,N_5043,N_5466);
or U5746 (N_5746,N_5250,N_5379);
or U5747 (N_5747,N_5174,N_5332);
nor U5748 (N_5748,N_5196,N_5467);
nand U5749 (N_5749,N_5264,N_5283);
nor U5750 (N_5750,N_5493,N_5396);
xor U5751 (N_5751,N_5157,N_5203);
and U5752 (N_5752,N_5437,N_5354);
xnor U5753 (N_5753,N_5116,N_5210);
nor U5754 (N_5754,N_5392,N_5337);
and U5755 (N_5755,N_5075,N_5022);
nor U5756 (N_5756,N_5058,N_5100);
xor U5757 (N_5757,N_5244,N_5411);
nand U5758 (N_5758,N_5073,N_5100);
xnor U5759 (N_5759,N_5195,N_5224);
and U5760 (N_5760,N_5219,N_5175);
xor U5761 (N_5761,N_5204,N_5241);
and U5762 (N_5762,N_5102,N_5039);
xnor U5763 (N_5763,N_5265,N_5078);
nand U5764 (N_5764,N_5434,N_5094);
and U5765 (N_5765,N_5019,N_5450);
nand U5766 (N_5766,N_5340,N_5178);
or U5767 (N_5767,N_5078,N_5093);
and U5768 (N_5768,N_5157,N_5400);
nand U5769 (N_5769,N_5477,N_5110);
nor U5770 (N_5770,N_5131,N_5350);
xor U5771 (N_5771,N_5118,N_5062);
or U5772 (N_5772,N_5095,N_5317);
or U5773 (N_5773,N_5034,N_5376);
or U5774 (N_5774,N_5483,N_5176);
or U5775 (N_5775,N_5411,N_5357);
nand U5776 (N_5776,N_5283,N_5059);
nor U5777 (N_5777,N_5075,N_5316);
xnor U5778 (N_5778,N_5074,N_5024);
nor U5779 (N_5779,N_5243,N_5156);
xor U5780 (N_5780,N_5462,N_5354);
xor U5781 (N_5781,N_5276,N_5040);
nand U5782 (N_5782,N_5320,N_5439);
nand U5783 (N_5783,N_5129,N_5068);
nand U5784 (N_5784,N_5034,N_5497);
nor U5785 (N_5785,N_5414,N_5080);
or U5786 (N_5786,N_5283,N_5048);
or U5787 (N_5787,N_5165,N_5337);
and U5788 (N_5788,N_5299,N_5051);
xnor U5789 (N_5789,N_5367,N_5423);
and U5790 (N_5790,N_5027,N_5374);
or U5791 (N_5791,N_5469,N_5284);
nor U5792 (N_5792,N_5146,N_5362);
or U5793 (N_5793,N_5373,N_5439);
and U5794 (N_5794,N_5440,N_5047);
xor U5795 (N_5795,N_5306,N_5213);
or U5796 (N_5796,N_5196,N_5173);
or U5797 (N_5797,N_5340,N_5292);
nand U5798 (N_5798,N_5036,N_5073);
or U5799 (N_5799,N_5489,N_5287);
nand U5800 (N_5800,N_5290,N_5227);
or U5801 (N_5801,N_5358,N_5428);
nand U5802 (N_5802,N_5336,N_5236);
xnor U5803 (N_5803,N_5469,N_5169);
nand U5804 (N_5804,N_5235,N_5282);
nand U5805 (N_5805,N_5316,N_5066);
and U5806 (N_5806,N_5099,N_5046);
nand U5807 (N_5807,N_5148,N_5357);
nor U5808 (N_5808,N_5365,N_5477);
xnor U5809 (N_5809,N_5135,N_5120);
or U5810 (N_5810,N_5272,N_5212);
nor U5811 (N_5811,N_5398,N_5145);
and U5812 (N_5812,N_5046,N_5082);
nor U5813 (N_5813,N_5010,N_5311);
xor U5814 (N_5814,N_5388,N_5466);
nor U5815 (N_5815,N_5462,N_5142);
and U5816 (N_5816,N_5111,N_5420);
and U5817 (N_5817,N_5263,N_5001);
and U5818 (N_5818,N_5431,N_5247);
or U5819 (N_5819,N_5417,N_5338);
nand U5820 (N_5820,N_5170,N_5149);
and U5821 (N_5821,N_5164,N_5248);
and U5822 (N_5822,N_5391,N_5434);
and U5823 (N_5823,N_5212,N_5348);
or U5824 (N_5824,N_5126,N_5186);
and U5825 (N_5825,N_5057,N_5110);
nor U5826 (N_5826,N_5156,N_5323);
nor U5827 (N_5827,N_5205,N_5472);
or U5828 (N_5828,N_5476,N_5164);
nand U5829 (N_5829,N_5294,N_5016);
nor U5830 (N_5830,N_5296,N_5362);
xor U5831 (N_5831,N_5232,N_5196);
nand U5832 (N_5832,N_5050,N_5293);
xnor U5833 (N_5833,N_5243,N_5492);
nand U5834 (N_5834,N_5417,N_5347);
nand U5835 (N_5835,N_5043,N_5163);
and U5836 (N_5836,N_5236,N_5166);
or U5837 (N_5837,N_5322,N_5005);
xor U5838 (N_5838,N_5220,N_5256);
nand U5839 (N_5839,N_5010,N_5497);
and U5840 (N_5840,N_5104,N_5201);
nor U5841 (N_5841,N_5075,N_5412);
and U5842 (N_5842,N_5017,N_5196);
and U5843 (N_5843,N_5090,N_5303);
nand U5844 (N_5844,N_5018,N_5485);
xor U5845 (N_5845,N_5188,N_5250);
and U5846 (N_5846,N_5306,N_5161);
nor U5847 (N_5847,N_5411,N_5498);
and U5848 (N_5848,N_5396,N_5009);
and U5849 (N_5849,N_5459,N_5116);
xnor U5850 (N_5850,N_5220,N_5311);
xnor U5851 (N_5851,N_5126,N_5447);
or U5852 (N_5852,N_5381,N_5191);
or U5853 (N_5853,N_5056,N_5110);
or U5854 (N_5854,N_5368,N_5074);
xnor U5855 (N_5855,N_5460,N_5097);
or U5856 (N_5856,N_5452,N_5261);
nand U5857 (N_5857,N_5418,N_5131);
or U5858 (N_5858,N_5188,N_5291);
and U5859 (N_5859,N_5455,N_5365);
nor U5860 (N_5860,N_5416,N_5241);
and U5861 (N_5861,N_5165,N_5308);
nor U5862 (N_5862,N_5006,N_5316);
nand U5863 (N_5863,N_5290,N_5452);
xnor U5864 (N_5864,N_5137,N_5184);
nor U5865 (N_5865,N_5214,N_5350);
and U5866 (N_5866,N_5480,N_5491);
nor U5867 (N_5867,N_5025,N_5233);
nand U5868 (N_5868,N_5325,N_5307);
nor U5869 (N_5869,N_5074,N_5124);
xor U5870 (N_5870,N_5099,N_5020);
or U5871 (N_5871,N_5357,N_5057);
and U5872 (N_5872,N_5370,N_5212);
and U5873 (N_5873,N_5196,N_5238);
xnor U5874 (N_5874,N_5032,N_5326);
nor U5875 (N_5875,N_5441,N_5114);
xor U5876 (N_5876,N_5147,N_5019);
nor U5877 (N_5877,N_5024,N_5156);
nor U5878 (N_5878,N_5448,N_5263);
or U5879 (N_5879,N_5186,N_5313);
or U5880 (N_5880,N_5475,N_5253);
and U5881 (N_5881,N_5040,N_5080);
nor U5882 (N_5882,N_5402,N_5116);
xor U5883 (N_5883,N_5334,N_5457);
or U5884 (N_5884,N_5061,N_5104);
or U5885 (N_5885,N_5448,N_5315);
nand U5886 (N_5886,N_5172,N_5301);
or U5887 (N_5887,N_5054,N_5413);
nand U5888 (N_5888,N_5172,N_5246);
xor U5889 (N_5889,N_5249,N_5264);
nand U5890 (N_5890,N_5476,N_5479);
xnor U5891 (N_5891,N_5280,N_5497);
nor U5892 (N_5892,N_5475,N_5034);
xor U5893 (N_5893,N_5054,N_5326);
nor U5894 (N_5894,N_5081,N_5498);
nand U5895 (N_5895,N_5377,N_5069);
and U5896 (N_5896,N_5211,N_5415);
nand U5897 (N_5897,N_5415,N_5188);
nor U5898 (N_5898,N_5007,N_5121);
nor U5899 (N_5899,N_5199,N_5456);
nand U5900 (N_5900,N_5405,N_5073);
xnor U5901 (N_5901,N_5012,N_5335);
xnor U5902 (N_5902,N_5387,N_5412);
nor U5903 (N_5903,N_5051,N_5147);
xnor U5904 (N_5904,N_5415,N_5072);
xor U5905 (N_5905,N_5237,N_5101);
nand U5906 (N_5906,N_5172,N_5354);
or U5907 (N_5907,N_5360,N_5225);
or U5908 (N_5908,N_5260,N_5458);
nor U5909 (N_5909,N_5096,N_5031);
and U5910 (N_5910,N_5475,N_5381);
nor U5911 (N_5911,N_5372,N_5385);
or U5912 (N_5912,N_5068,N_5321);
xor U5913 (N_5913,N_5241,N_5497);
xnor U5914 (N_5914,N_5132,N_5404);
xor U5915 (N_5915,N_5216,N_5335);
nand U5916 (N_5916,N_5346,N_5349);
nand U5917 (N_5917,N_5354,N_5332);
or U5918 (N_5918,N_5466,N_5014);
and U5919 (N_5919,N_5103,N_5405);
nor U5920 (N_5920,N_5186,N_5256);
nand U5921 (N_5921,N_5093,N_5227);
or U5922 (N_5922,N_5178,N_5379);
nor U5923 (N_5923,N_5447,N_5014);
nor U5924 (N_5924,N_5120,N_5090);
nor U5925 (N_5925,N_5172,N_5382);
xnor U5926 (N_5926,N_5076,N_5469);
and U5927 (N_5927,N_5171,N_5146);
and U5928 (N_5928,N_5340,N_5009);
nand U5929 (N_5929,N_5360,N_5389);
nor U5930 (N_5930,N_5185,N_5240);
and U5931 (N_5931,N_5453,N_5179);
nand U5932 (N_5932,N_5240,N_5241);
or U5933 (N_5933,N_5450,N_5408);
nand U5934 (N_5934,N_5304,N_5292);
nand U5935 (N_5935,N_5045,N_5217);
or U5936 (N_5936,N_5264,N_5484);
nor U5937 (N_5937,N_5098,N_5004);
and U5938 (N_5938,N_5126,N_5011);
nor U5939 (N_5939,N_5135,N_5000);
or U5940 (N_5940,N_5167,N_5345);
nor U5941 (N_5941,N_5110,N_5079);
or U5942 (N_5942,N_5431,N_5135);
nor U5943 (N_5943,N_5418,N_5262);
xor U5944 (N_5944,N_5303,N_5023);
nor U5945 (N_5945,N_5117,N_5497);
nand U5946 (N_5946,N_5496,N_5151);
xor U5947 (N_5947,N_5366,N_5014);
or U5948 (N_5948,N_5455,N_5287);
or U5949 (N_5949,N_5424,N_5331);
xor U5950 (N_5950,N_5005,N_5175);
nor U5951 (N_5951,N_5292,N_5425);
or U5952 (N_5952,N_5170,N_5429);
or U5953 (N_5953,N_5147,N_5105);
xnor U5954 (N_5954,N_5419,N_5001);
nand U5955 (N_5955,N_5092,N_5322);
nor U5956 (N_5956,N_5235,N_5189);
or U5957 (N_5957,N_5213,N_5076);
xnor U5958 (N_5958,N_5223,N_5428);
nand U5959 (N_5959,N_5242,N_5305);
or U5960 (N_5960,N_5345,N_5153);
nand U5961 (N_5961,N_5127,N_5208);
nor U5962 (N_5962,N_5129,N_5069);
xor U5963 (N_5963,N_5001,N_5235);
and U5964 (N_5964,N_5221,N_5029);
xnor U5965 (N_5965,N_5207,N_5345);
nor U5966 (N_5966,N_5067,N_5235);
and U5967 (N_5967,N_5093,N_5083);
xor U5968 (N_5968,N_5371,N_5184);
and U5969 (N_5969,N_5149,N_5271);
and U5970 (N_5970,N_5200,N_5010);
and U5971 (N_5971,N_5070,N_5233);
or U5972 (N_5972,N_5352,N_5275);
or U5973 (N_5973,N_5432,N_5415);
xor U5974 (N_5974,N_5463,N_5468);
and U5975 (N_5975,N_5108,N_5274);
nor U5976 (N_5976,N_5139,N_5172);
nand U5977 (N_5977,N_5113,N_5037);
nand U5978 (N_5978,N_5021,N_5235);
or U5979 (N_5979,N_5382,N_5044);
xor U5980 (N_5980,N_5465,N_5482);
or U5981 (N_5981,N_5124,N_5226);
and U5982 (N_5982,N_5492,N_5225);
and U5983 (N_5983,N_5321,N_5472);
nand U5984 (N_5984,N_5107,N_5385);
and U5985 (N_5985,N_5023,N_5267);
xor U5986 (N_5986,N_5486,N_5442);
or U5987 (N_5987,N_5168,N_5442);
nor U5988 (N_5988,N_5129,N_5066);
nand U5989 (N_5989,N_5214,N_5207);
and U5990 (N_5990,N_5149,N_5294);
xnor U5991 (N_5991,N_5335,N_5341);
or U5992 (N_5992,N_5281,N_5296);
xor U5993 (N_5993,N_5378,N_5042);
nor U5994 (N_5994,N_5025,N_5086);
xor U5995 (N_5995,N_5431,N_5359);
nand U5996 (N_5996,N_5020,N_5000);
and U5997 (N_5997,N_5428,N_5464);
nand U5998 (N_5998,N_5421,N_5209);
xnor U5999 (N_5999,N_5165,N_5192);
xnor U6000 (N_6000,N_5773,N_5598);
and U6001 (N_6001,N_5814,N_5659);
or U6002 (N_6002,N_5990,N_5944);
and U6003 (N_6003,N_5749,N_5796);
nand U6004 (N_6004,N_5599,N_5913);
xor U6005 (N_6005,N_5508,N_5987);
and U6006 (N_6006,N_5891,N_5689);
nor U6007 (N_6007,N_5756,N_5866);
or U6008 (N_6008,N_5658,N_5713);
or U6009 (N_6009,N_5730,N_5981);
and U6010 (N_6010,N_5742,N_5646);
or U6011 (N_6011,N_5989,N_5668);
xnor U6012 (N_6012,N_5531,N_5558);
and U6013 (N_6013,N_5760,N_5771);
and U6014 (N_6014,N_5840,N_5665);
or U6015 (N_6015,N_5770,N_5863);
or U6016 (N_6016,N_5833,N_5893);
nand U6017 (N_6017,N_5739,N_5754);
and U6018 (N_6018,N_5504,N_5575);
and U6019 (N_6019,N_5560,N_5864);
or U6020 (N_6020,N_5835,N_5696);
nand U6021 (N_6021,N_5523,N_5663);
and U6022 (N_6022,N_5967,N_5830);
xor U6023 (N_6023,N_5505,N_5831);
nand U6024 (N_6024,N_5842,N_5611);
nand U6025 (N_6025,N_5861,N_5769);
and U6026 (N_6026,N_5795,N_5894);
nor U6027 (N_6027,N_5594,N_5675);
or U6028 (N_6028,N_5532,N_5536);
nor U6029 (N_6029,N_5927,N_5743);
or U6030 (N_6030,N_5964,N_5746);
nand U6031 (N_6031,N_5661,N_5731);
or U6032 (N_6032,N_5841,N_5709);
xor U6033 (N_6033,N_5670,N_5682);
and U6034 (N_6034,N_5774,N_5643);
or U6035 (N_6035,N_5512,N_5867);
nand U6036 (N_6036,N_5541,N_5984);
xor U6037 (N_6037,N_5951,N_5895);
xnor U6038 (N_6038,N_5591,N_5823);
xor U6039 (N_6039,N_5566,N_5919);
nor U6040 (N_6040,N_5603,N_5715);
nor U6041 (N_6041,N_5677,N_5684);
nor U6042 (N_6042,N_5667,N_5537);
or U6043 (N_6043,N_5828,N_5524);
and U6044 (N_6044,N_5642,N_5681);
or U6045 (N_6045,N_5688,N_5705);
nand U6046 (N_6046,N_5819,N_5837);
nand U6047 (N_6047,N_5971,N_5717);
nand U6048 (N_6048,N_5551,N_5865);
nand U6049 (N_6049,N_5776,N_5953);
and U6050 (N_6050,N_5857,N_5647);
and U6051 (N_6051,N_5683,N_5935);
and U6052 (N_6052,N_5763,N_5539);
and U6053 (N_6053,N_5938,N_5645);
nor U6054 (N_6054,N_5534,N_5936);
nand U6055 (N_6055,N_5597,N_5888);
or U6056 (N_6056,N_5982,N_5615);
and U6057 (N_6057,N_5641,N_5593);
and U6058 (N_6058,N_5966,N_5884);
xnor U6059 (N_6059,N_5589,N_5801);
nand U6060 (N_6060,N_5565,N_5847);
nor U6061 (N_6061,N_5587,N_5772);
xnor U6062 (N_6062,N_5979,N_5764);
nand U6063 (N_6063,N_5704,N_5970);
xnor U6064 (N_6064,N_5555,N_5529);
or U6065 (N_6065,N_5744,N_5917);
nor U6066 (N_6066,N_5693,N_5502);
nor U6067 (N_6067,N_5650,N_5716);
nor U6068 (N_6068,N_5903,N_5997);
or U6069 (N_6069,N_5880,N_5602);
or U6070 (N_6070,N_5649,N_5520);
nor U6071 (N_6071,N_5718,N_5952);
or U6072 (N_6072,N_5526,N_5872);
nand U6073 (N_6073,N_5859,N_5563);
nand U6074 (N_6074,N_5925,N_5932);
nand U6075 (N_6075,N_5889,N_5994);
or U6076 (N_6076,N_5877,N_5965);
xor U6077 (N_6077,N_5825,N_5584);
or U6078 (N_6078,N_5768,N_5573);
and U6079 (N_6079,N_5692,N_5777);
and U6080 (N_6080,N_5601,N_5609);
nor U6081 (N_6081,N_5588,N_5695);
nor U6082 (N_6082,N_5900,N_5781);
xnor U6083 (N_6083,N_5562,N_5910);
xnor U6084 (N_6084,N_5660,N_5701);
nor U6085 (N_6085,N_5912,N_5923);
xnor U6086 (N_6086,N_5875,N_5654);
nor U6087 (N_6087,N_5921,N_5725);
or U6088 (N_6088,N_5623,N_5829);
or U6089 (N_6089,N_5871,N_5977);
nor U6090 (N_6090,N_5518,N_5862);
nand U6091 (N_6091,N_5904,N_5758);
nor U6092 (N_6092,N_5726,N_5976);
xnor U6093 (N_6093,N_5519,N_5902);
nand U6094 (N_6094,N_5707,N_5652);
xnor U6095 (N_6095,N_5712,N_5873);
and U6096 (N_6096,N_5636,N_5515);
nand U6097 (N_6097,N_5991,N_5920);
or U6098 (N_6098,N_5530,N_5929);
and U6099 (N_6099,N_5897,N_5736);
nor U6100 (N_6100,N_5685,N_5948);
and U6101 (N_6101,N_5996,N_5974);
xor U6102 (N_6102,N_5915,N_5583);
and U6103 (N_6103,N_5782,N_5644);
nand U6104 (N_6104,N_5800,N_5896);
nor U6105 (N_6105,N_5568,N_5784);
nor U6106 (N_6106,N_5822,N_5592);
or U6107 (N_6107,N_5501,N_5885);
xnor U6108 (N_6108,N_5590,N_5687);
nor U6109 (N_6109,N_5559,N_5552);
and U6110 (N_6110,N_5824,N_5627);
or U6111 (N_6111,N_5582,N_5890);
or U6112 (N_6112,N_5748,N_5905);
xor U6113 (N_6113,N_5613,N_5858);
and U6114 (N_6114,N_5918,N_5954);
xnor U6115 (N_6115,N_5617,N_5561);
and U6116 (N_6116,N_5878,N_5516);
xnor U6117 (N_6117,N_5803,N_5507);
nor U6118 (N_6118,N_5631,N_5755);
nor U6119 (N_6119,N_5616,N_5943);
and U6120 (N_6120,N_5852,N_5995);
and U6121 (N_6121,N_5849,N_5999);
and U6122 (N_6122,N_5564,N_5838);
or U6123 (N_6123,N_5664,N_5678);
and U6124 (N_6124,N_5699,N_5815);
nand U6125 (N_6125,N_5789,N_5901);
and U6126 (N_6126,N_5785,N_5899);
nor U6127 (N_6127,N_5757,N_5503);
nand U6128 (N_6128,N_5549,N_5998);
and U6129 (N_6129,N_5850,N_5939);
or U6130 (N_6130,N_5596,N_5848);
xor U6131 (N_6131,N_5805,N_5811);
nand U6132 (N_6132,N_5972,N_5787);
or U6133 (N_6133,N_5914,N_5691);
xnor U6134 (N_6134,N_5703,N_5628);
xor U6135 (N_6135,N_5832,N_5876);
xor U6136 (N_6136,N_5638,N_5506);
and U6137 (N_6137,N_5942,N_5543);
nor U6138 (N_6138,N_5514,N_5607);
nor U6139 (N_6139,N_5922,N_5765);
and U6140 (N_6140,N_5633,N_5723);
xor U6141 (N_6141,N_5606,N_5540);
xnor U6142 (N_6142,N_5629,N_5874);
or U6143 (N_6143,N_5993,N_5957);
xnor U6144 (N_6144,N_5724,N_5686);
nor U6145 (N_6145,N_5992,N_5916);
and U6146 (N_6146,N_5797,N_5786);
or U6147 (N_6147,N_5557,N_5887);
nand U6148 (N_6148,N_5567,N_5535);
nor U6149 (N_6149,N_5585,N_5522);
and U6150 (N_6150,N_5752,N_5767);
and U6151 (N_6151,N_5793,N_5856);
nand U6152 (N_6152,N_5794,N_5818);
and U6153 (N_6153,N_5595,N_5745);
nor U6154 (N_6154,N_5930,N_5986);
nand U6155 (N_6155,N_5580,N_5812);
and U6156 (N_6156,N_5721,N_5816);
nor U6157 (N_6157,N_5853,N_5985);
and U6158 (N_6158,N_5546,N_5554);
nor U6159 (N_6159,N_5751,N_5621);
and U6160 (N_6160,N_5517,N_5711);
xor U6161 (N_6161,N_5578,N_5836);
xnor U6162 (N_6162,N_5651,N_5740);
xnor U6163 (N_6163,N_5955,N_5655);
nand U6164 (N_6164,N_5733,N_5624);
xnor U6165 (N_6165,N_5720,N_5612);
xnor U6166 (N_6166,N_5576,N_5706);
nor U6167 (N_6167,N_5750,N_5639);
or U6168 (N_6168,N_5734,N_5924);
nand U6169 (N_6169,N_5538,N_5940);
and U6170 (N_6170,N_5732,N_5779);
or U6171 (N_6171,N_5956,N_5934);
xnor U6172 (N_6172,N_5574,N_5525);
or U6173 (N_6173,N_5988,N_5572);
or U6174 (N_6174,N_5958,N_5571);
nor U6175 (N_6175,N_5653,N_5635);
xor U6176 (N_6176,N_5963,N_5926);
and U6177 (N_6177,N_5845,N_5962);
nand U6178 (N_6178,N_5556,N_5969);
and U6179 (N_6179,N_5809,N_5820);
nand U6180 (N_6180,N_5855,N_5545);
nor U6181 (N_6181,N_5759,N_5608);
nand U6182 (N_6182,N_5610,N_5806);
or U6183 (N_6183,N_5719,N_5834);
nor U6184 (N_6184,N_5960,N_5947);
nand U6185 (N_6185,N_5911,N_5618);
or U6186 (N_6186,N_5778,N_5860);
xor U6187 (N_6187,N_5622,N_5700);
xnor U6188 (N_6188,N_5714,N_5528);
or U6189 (N_6189,N_5509,N_5933);
nor U6190 (N_6190,N_5799,N_5737);
and U6191 (N_6191,N_5791,N_5702);
nor U6192 (N_6192,N_5586,N_5780);
nor U6193 (N_6193,N_5679,N_5980);
and U6194 (N_6194,N_5600,N_5634);
nand U6195 (N_6195,N_5883,N_5881);
nand U6196 (N_6196,N_5698,N_5500);
xnor U6197 (N_6197,N_5729,N_5843);
xnor U6198 (N_6198,N_5513,N_5738);
and U6199 (N_6199,N_5727,N_5978);
and U6200 (N_6200,N_5869,N_5908);
xnor U6201 (N_6201,N_5625,N_5827);
nor U6202 (N_6202,N_5808,N_5846);
or U6203 (N_6203,N_5975,N_5868);
nor U6204 (N_6204,N_5640,N_5870);
or U6205 (N_6205,N_5882,N_5804);
nor U6206 (N_6206,N_5968,N_5762);
nand U6207 (N_6207,N_5826,N_5662);
xor U6208 (N_6208,N_5983,N_5569);
nand U6209 (N_6209,N_5619,N_5673);
xor U6210 (N_6210,N_5550,N_5510);
and U6211 (N_6211,N_5632,N_5680);
and U6212 (N_6212,N_5614,N_5937);
xor U6213 (N_6213,N_5527,N_5690);
nor U6214 (N_6214,N_5810,N_5669);
and U6215 (N_6215,N_5898,N_5626);
xnor U6216 (N_6216,N_5839,N_5931);
nand U6217 (N_6217,N_5722,N_5959);
and U6218 (N_6218,N_5656,N_5973);
or U6219 (N_6219,N_5945,N_5821);
xnor U6220 (N_6220,N_5544,N_5604);
and U6221 (N_6221,N_5676,N_5542);
and U6222 (N_6222,N_5844,N_5671);
xnor U6223 (N_6223,N_5946,N_5728);
or U6224 (N_6224,N_5708,N_5788);
or U6225 (N_6225,N_5941,N_5694);
or U6226 (N_6226,N_5766,N_5548);
or U6227 (N_6227,N_5851,N_5892);
nand U6228 (N_6228,N_5741,N_5521);
xnor U6229 (N_6229,N_5672,N_5637);
nand U6230 (N_6230,N_5854,N_5906);
and U6231 (N_6231,N_5783,N_5547);
xor U6232 (N_6232,N_5674,N_5886);
and U6233 (N_6233,N_5735,N_5533);
nand U6234 (N_6234,N_5697,N_5710);
nand U6235 (N_6235,N_5907,N_5657);
xor U6236 (N_6236,N_5511,N_5802);
nand U6237 (N_6237,N_5630,N_5605);
or U6238 (N_6238,N_5798,N_5950);
xor U6239 (N_6239,N_5648,N_5775);
and U6240 (N_6240,N_5753,N_5961);
and U6241 (N_6241,N_5928,N_5807);
nand U6242 (N_6242,N_5909,N_5581);
nand U6243 (N_6243,N_5817,N_5579);
xor U6244 (N_6244,N_5620,N_5879);
nand U6245 (N_6245,N_5790,N_5570);
nor U6246 (N_6246,N_5792,N_5553);
nand U6247 (N_6247,N_5577,N_5747);
or U6248 (N_6248,N_5761,N_5666);
xnor U6249 (N_6249,N_5813,N_5949);
nand U6250 (N_6250,N_5821,N_5841);
nor U6251 (N_6251,N_5755,N_5653);
and U6252 (N_6252,N_5794,N_5579);
or U6253 (N_6253,N_5899,N_5879);
nand U6254 (N_6254,N_5677,N_5598);
nor U6255 (N_6255,N_5715,N_5527);
or U6256 (N_6256,N_5831,N_5526);
and U6257 (N_6257,N_5574,N_5621);
xor U6258 (N_6258,N_5741,N_5961);
nor U6259 (N_6259,N_5912,N_5991);
and U6260 (N_6260,N_5976,N_5730);
nand U6261 (N_6261,N_5866,N_5788);
or U6262 (N_6262,N_5898,N_5868);
nor U6263 (N_6263,N_5587,N_5506);
xnor U6264 (N_6264,N_5586,N_5999);
xnor U6265 (N_6265,N_5586,N_5587);
or U6266 (N_6266,N_5991,N_5763);
and U6267 (N_6267,N_5566,N_5862);
or U6268 (N_6268,N_5630,N_5829);
and U6269 (N_6269,N_5639,N_5983);
nor U6270 (N_6270,N_5914,N_5836);
nand U6271 (N_6271,N_5953,N_5843);
nor U6272 (N_6272,N_5600,N_5934);
nand U6273 (N_6273,N_5734,N_5723);
nand U6274 (N_6274,N_5913,N_5504);
nor U6275 (N_6275,N_5511,N_5588);
nand U6276 (N_6276,N_5725,N_5624);
xor U6277 (N_6277,N_5694,N_5619);
and U6278 (N_6278,N_5884,N_5817);
nor U6279 (N_6279,N_5849,N_5859);
xor U6280 (N_6280,N_5779,N_5555);
xor U6281 (N_6281,N_5646,N_5897);
xor U6282 (N_6282,N_5658,N_5876);
nor U6283 (N_6283,N_5953,N_5614);
and U6284 (N_6284,N_5948,N_5967);
xor U6285 (N_6285,N_5629,N_5962);
and U6286 (N_6286,N_5672,N_5734);
nor U6287 (N_6287,N_5706,N_5626);
xnor U6288 (N_6288,N_5554,N_5927);
xnor U6289 (N_6289,N_5980,N_5600);
and U6290 (N_6290,N_5713,N_5564);
xor U6291 (N_6291,N_5730,N_5584);
xnor U6292 (N_6292,N_5939,N_5844);
and U6293 (N_6293,N_5822,N_5914);
nand U6294 (N_6294,N_5865,N_5507);
nand U6295 (N_6295,N_5948,N_5934);
nand U6296 (N_6296,N_5797,N_5678);
xor U6297 (N_6297,N_5550,N_5698);
xnor U6298 (N_6298,N_5831,N_5813);
xnor U6299 (N_6299,N_5500,N_5614);
nand U6300 (N_6300,N_5970,N_5820);
nor U6301 (N_6301,N_5664,N_5540);
and U6302 (N_6302,N_5777,N_5698);
nor U6303 (N_6303,N_5750,N_5972);
or U6304 (N_6304,N_5580,N_5603);
nand U6305 (N_6305,N_5944,N_5926);
xor U6306 (N_6306,N_5555,N_5616);
and U6307 (N_6307,N_5762,N_5862);
xor U6308 (N_6308,N_5581,N_5699);
nand U6309 (N_6309,N_5698,N_5679);
nor U6310 (N_6310,N_5874,N_5795);
nor U6311 (N_6311,N_5884,N_5641);
or U6312 (N_6312,N_5751,N_5744);
and U6313 (N_6313,N_5896,N_5517);
nand U6314 (N_6314,N_5949,N_5802);
nand U6315 (N_6315,N_5580,N_5792);
nor U6316 (N_6316,N_5960,N_5761);
or U6317 (N_6317,N_5803,N_5996);
xnor U6318 (N_6318,N_5819,N_5723);
or U6319 (N_6319,N_5621,N_5925);
or U6320 (N_6320,N_5603,N_5698);
and U6321 (N_6321,N_5625,N_5832);
or U6322 (N_6322,N_5870,N_5772);
and U6323 (N_6323,N_5861,N_5521);
nor U6324 (N_6324,N_5911,N_5951);
nor U6325 (N_6325,N_5780,N_5867);
and U6326 (N_6326,N_5763,N_5837);
xor U6327 (N_6327,N_5592,N_5511);
nand U6328 (N_6328,N_5639,N_5636);
nand U6329 (N_6329,N_5743,N_5944);
nand U6330 (N_6330,N_5985,N_5565);
or U6331 (N_6331,N_5757,N_5838);
nand U6332 (N_6332,N_5770,N_5673);
xor U6333 (N_6333,N_5915,N_5958);
nand U6334 (N_6334,N_5638,N_5538);
xnor U6335 (N_6335,N_5827,N_5991);
and U6336 (N_6336,N_5815,N_5647);
xor U6337 (N_6337,N_5933,N_5928);
nor U6338 (N_6338,N_5604,N_5783);
and U6339 (N_6339,N_5907,N_5542);
or U6340 (N_6340,N_5778,N_5701);
nand U6341 (N_6341,N_5800,N_5879);
nor U6342 (N_6342,N_5943,N_5879);
or U6343 (N_6343,N_5851,N_5771);
or U6344 (N_6344,N_5789,N_5814);
nor U6345 (N_6345,N_5659,N_5885);
nor U6346 (N_6346,N_5884,N_5600);
xor U6347 (N_6347,N_5694,N_5625);
nor U6348 (N_6348,N_5863,N_5946);
xnor U6349 (N_6349,N_5905,N_5601);
and U6350 (N_6350,N_5798,N_5776);
and U6351 (N_6351,N_5975,N_5854);
and U6352 (N_6352,N_5635,N_5706);
and U6353 (N_6353,N_5508,N_5700);
nor U6354 (N_6354,N_5786,N_5785);
nor U6355 (N_6355,N_5732,N_5586);
nor U6356 (N_6356,N_5508,N_5701);
or U6357 (N_6357,N_5670,N_5539);
xor U6358 (N_6358,N_5827,N_5980);
nand U6359 (N_6359,N_5963,N_5805);
or U6360 (N_6360,N_5743,N_5792);
nor U6361 (N_6361,N_5784,N_5598);
nor U6362 (N_6362,N_5926,N_5537);
or U6363 (N_6363,N_5870,N_5530);
or U6364 (N_6364,N_5958,N_5795);
or U6365 (N_6365,N_5554,N_5585);
or U6366 (N_6366,N_5680,N_5625);
xor U6367 (N_6367,N_5910,N_5896);
xor U6368 (N_6368,N_5843,N_5929);
xnor U6369 (N_6369,N_5777,N_5682);
and U6370 (N_6370,N_5633,N_5931);
and U6371 (N_6371,N_5745,N_5843);
nand U6372 (N_6372,N_5515,N_5528);
and U6373 (N_6373,N_5815,N_5619);
and U6374 (N_6374,N_5518,N_5914);
or U6375 (N_6375,N_5589,N_5955);
or U6376 (N_6376,N_5938,N_5540);
xor U6377 (N_6377,N_5511,N_5864);
xor U6378 (N_6378,N_5506,N_5925);
nor U6379 (N_6379,N_5832,N_5508);
xnor U6380 (N_6380,N_5553,N_5925);
or U6381 (N_6381,N_5996,N_5550);
nand U6382 (N_6382,N_5610,N_5900);
nor U6383 (N_6383,N_5948,N_5896);
xor U6384 (N_6384,N_5569,N_5615);
nand U6385 (N_6385,N_5693,N_5611);
nand U6386 (N_6386,N_5635,N_5997);
and U6387 (N_6387,N_5573,N_5837);
nor U6388 (N_6388,N_5859,N_5911);
xnor U6389 (N_6389,N_5660,N_5551);
nand U6390 (N_6390,N_5988,N_5866);
xor U6391 (N_6391,N_5834,N_5760);
xnor U6392 (N_6392,N_5588,N_5856);
and U6393 (N_6393,N_5708,N_5799);
xor U6394 (N_6394,N_5677,N_5997);
or U6395 (N_6395,N_5566,N_5504);
xor U6396 (N_6396,N_5610,N_5523);
nor U6397 (N_6397,N_5529,N_5848);
nand U6398 (N_6398,N_5715,N_5690);
nand U6399 (N_6399,N_5761,N_5600);
xor U6400 (N_6400,N_5639,N_5856);
nor U6401 (N_6401,N_5509,N_5786);
xnor U6402 (N_6402,N_5521,N_5571);
or U6403 (N_6403,N_5685,N_5520);
xor U6404 (N_6404,N_5738,N_5781);
and U6405 (N_6405,N_5685,N_5940);
and U6406 (N_6406,N_5923,N_5614);
nor U6407 (N_6407,N_5918,N_5519);
nor U6408 (N_6408,N_5735,N_5933);
nand U6409 (N_6409,N_5964,N_5906);
xor U6410 (N_6410,N_5582,N_5748);
or U6411 (N_6411,N_5663,N_5993);
nand U6412 (N_6412,N_5509,N_5807);
nor U6413 (N_6413,N_5657,N_5872);
nor U6414 (N_6414,N_5711,N_5595);
or U6415 (N_6415,N_5874,N_5920);
nor U6416 (N_6416,N_5680,N_5738);
and U6417 (N_6417,N_5717,N_5547);
and U6418 (N_6418,N_5922,N_5658);
nor U6419 (N_6419,N_5798,N_5953);
or U6420 (N_6420,N_5541,N_5887);
nand U6421 (N_6421,N_5649,N_5875);
and U6422 (N_6422,N_5532,N_5824);
nand U6423 (N_6423,N_5785,N_5553);
xor U6424 (N_6424,N_5603,N_5539);
xnor U6425 (N_6425,N_5925,N_5682);
nand U6426 (N_6426,N_5935,N_5781);
xnor U6427 (N_6427,N_5914,N_5636);
nand U6428 (N_6428,N_5866,N_5641);
xor U6429 (N_6429,N_5816,N_5937);
or U6430 (N_6430,N_5689,N_5537);
nor U6431 (N_6431,N_5870,N_5865);
xnor U6432 (N_6432,N_5690,N_5863);
or U6433 (N_6433,N_5532,N_5747);
xor U6434 (N_6434,N_5753,N_5630);
and U6435 (N_6435,N_5553,N_5653);
and U6436 (N_6436,N_5740,N_5726);
nand U6437 (N_6437,N_5947,N_5799);
and U6438 (N_6438,N_5517,N_5557);
or U6439 (N_6439,N_5604,N_5601);
nor U6440 (N_6440,N_5921,N_5981);
nor U6441 (N_6441,N_5972,N_5886);
nor U6442 (N_6442,N_5586,N_5930);
nand U6443 (N_6443,N_5646,N_5564);
or U6444 (N_6444,N_5933,N_5564);
nor U6445 (N_6445,N_5522,N_5518);
xnor U6446 (N_6446,N_5871,N_5924);
nand U6447 (N_6447,N_5609,N_5762);
nor U6448 (N_6448,N_5927,N_5842);
or U6449 (N_6449,N_5725,N_5922);
or U6450 (N_6450,N_5949,N_5933);
and U6451 (N_6451,N_5898,N_5766);
or U6452 (N_6452,N_5643,N_5955);
nand U6453 (N_6453,N_5709,N_5683);
xnor U6454 (N_6454,N_5940,N_5827);
nand U6455 (N_6455,N_5588,N_5840);
xnor U6456 (N_6456,N_5820,N_5684);
nor U6457 (N_6457,N_5594,N_5633);
and U6458 (N_6458,N_5689,N_5653);
nand U6459 (N_6459,N_5727,N_5706);
nand U6460 (N_6460,N_5788,N_5626);
xnor U6461 (N_6461,N_5505,N_5554);
nor U6462 (N_6462,N_5574,N_5784);
nand U6463 (N_6463,N_5736,N_5918);
and U6464 (N_6464,N_5873,N_5741);
nand U6465 (N_6465,N_5724,N_5715);
nand U6466 (N_6466,N_5677,N_5939);
nor U6467 (N_6467,N_5882,N_5958);
xnor U6468 (N_6468,N_5653,N_5800);
nor U6469 (N_6469,N_5552,N_5971);
nor U6470 (N_6470,N_5780,N_5894);
xnor U6471 (N_6471,N_5862,N_5683);
or U6472 (N_6472,N_5963,N_5607);
and U6473 (N_6473,N_5998,N_5745);
or U6474 (N_6474,N_5964,N_5977);
xor U6475 (N_6475,N_5595,N_5791);
nand U6476 (N_6476,N_5575,N_5841);
and U6477 (N_6477,N_5933,N_5969);
xor U6478 (N_6478,N_5533,N_5722);
nand U6479 (N_6479,N_5625,N_5843);
or U6480 (N_6480,N_5719,N_5677);
xnor U6481 (N_6481,N_5701,N_5517);
nor U6482 (N_6482,N_5884,N_5697);
nand U6483 (N_6483,N_5640,N_5647);
nand U6484 (N_6484,N_5739,N_5704);
nor U6485 (N_6485,N_5711,N_5587);
nand U6486 (N_6486,N_5957,N_5750);
xor U6487 (N_6487,N_5970,N_5702);
nor U6488 (N_6488,N_5864,N_5721);
nor U6489 (N_6489,N_5804,N_5705);
or U6490 (N_6490,N_5764,N_5834);
nor U6491 (N_6491,N_5648,N_5713);
nand U6492 (N_6492,N_5716,N_5692);
nor U6493 (N_6493,N_5921,N_5582);
and U6494 (N_6494,N_5881,N_5564);
or U6495 (N_6495,N_5526,N_5736);
nand U6496 (N_6496,N_5662,N_5586);
nand U6497 (N_6497,N_5812,N_5925);
or U6498 (N_6498,N_5952,N_5604);
nor U6499 (N_6499,N_5990,N_5637);
and U6500 (N_6500,N_6041,N_6177);
nand U6501 (N_6501,N_6308,N_6231);
nor U6502 (N_6502,N_6380,N_6346);
and U6503 (N_6503,N_6127,N_6182);
nor U6504 (N_6504,N_6357,N_6165);
xnor U6505 (N_6505,N_6312,N_6491);
or U6506 (N_6506,N_6303,N_6112);
nand U6507 (N_6507,N_6394,N_6190);
or U6508 (N_6508,N_6474,N_6063);
and U6509 (N_6509,N_6245,N_6388);
nor U6510 (N_6510,N_6289,N_6338);
xor U6511 (N_6511,N_6123,N_6233);
xnor U6512 (N_6512,N_6129,N_6049);
xnor U6513 (N_6513,N_6438,N_6444);
xor U6514 (N_6514,N_6017,N_6087);
xor U6515 (N_6515,N_6354,N_6408);
nand U6516 (N_6516,N_6158,N_6478);
or U6517 (N_6517,N_6159,N_6028);
xnor U6518 (N_6518,N_6389,N_6430);
nand U6519 (N_6519,N_6323,N_6442);
nand U6520 (N_6520,N_6268,N_6241);
or U6521 (N_6521,N_6193,N_6180);
nor U6522 (N_6522,N_6196,N_6113);
nand U6523 (N_6523,N_6061,N_6476);
nor U6524 (N_6524,N_6092,N_6284);
nand U6525 (N_6525,N_6181,N_6214);
nor U6526 (N_6526,N_6424,N_6014);
xnor U6527 (N_6527,N_6269,N_6333);
nand U6528 (N_6528,N_6296,N_6316);
or U6529 (N_6529,N_6151,N_6257);
or U6530 (N_6530,N_6213,N_6383);
and U6531 (N_6531,N_6232,N_6201);
nand U6532 (N_6532,N_6155,N_6412);
and U6533 (N_6533,N_6216,N_6465);
and U6534 (N_6534,N_6433,N_6314);
or U6535 (N_6535,N_6162,N_6148);
nor U6536 (N_6536,N_6105,N_6337);
nand U6537 (N_6537,N_6342,N_6076);
nand U6538 (N_6538,N_6089,N_6117);
xor U6539 (N_6539,N_6208,N_6276);
nor U6540 (N_6540,N_6485,N_6139);
xor U6541 (N_6541,N_6223,N_6083);
nand U6542 (N_6542,N_6043,N_6425);
or U6543 (N_6543,N_6418,N_6225);
and U6544 (N_6544,N_6115,N_6149);
or U6545 (N_6545,N_6362,N_6184);
and U6546 (N_6546,N_6179,N_6070);
xor U6547 (N_6547,N_6454,N_6126);
nor U6548 (N_6548,N_6174,N_6237);
nand U6549 (N_6549,N_6494,N_6359);
or U6550 (N_6550,N_6283,N_6248);
nand U6551 (N_6551,N_6470,N_6456);
nor U6552 (N_6552,N_6263,N_6172);
xnor U6553 (N_6553,N_6031,N_6288);
xor U6554 (N_6554,N_6138,N_6277);
xnor U6555 (N_6555,N_6422,N_6447);
xor U6556 (N_6556,N_6479,N_6004);
xnor U6557 (N_6557,N_6038,N_6492);
or U6558 (N_6558,N_6067,N_6009);
or U6559 (N_6559,N_6496,N_6020);
or U6560 (N_6560,N_6265,N_6091);
nand U6561 (N_6561,N_6484,N_6417);
or U6562 (N_6562,N_6152,N_6207);
nand U6563 (N_6563,N_6315,N_6219);
nor U6564 (N_6564,N_6355,N_6464);
nand U6565 (N_6565,N_6431,N_6317);
xnor U6566 (N_6566,N_6301,N_6048);
and U6567 (N_6567,N_6185,N_6254);
and U6568 (N_6568,N_6104,N_6025);
nand U6569 (N_6569,N_6064,N_6399);
and U6570 (N_6570,N_6015,N_6285);
nand U6571 (N_6571,N_6351,N_6490);
and U6572 (N_6572,N_6413,N_6081);
nor U6573 (N_6573,N_6475,N_6403);
nor U6574 (N_6574,N_6239,N_6000);
xor U6575 (N_6575,N_6090,N_6255);
or U6576 (N_6576,N_6221,N_6347);
or U6577 (N_6577,N_6194,N_6421);
nor U6578 (N_6578,N_6037,N_6175);
or U6579 (N_6579,N_6075,N_6411);
and U6580 (N_6580,N_6209,N_6183);
xor U6581 (N_6581,N_6393,N_6125);
nand U6582 (N_6582,N_6116,N_6471);
nor U6583 (N_6583,N_6198,N_6261);
nand U6584 (N_6584,N_6450,N_6376);
xor U6585 (N_6585,N_6143,N_6085);
xnor U6586 (N_6586,N_6032,N_6266);
or U6587 (N_6587,N_6186,N_6170);
or U6588 (N_6588,N_6229,N_6097);
xor U6589 (N_6589,N_6121,N_6311);
and U6590 (N_6590,N_6042,N_6488);
nor U6591 (N_6591,N_6205,N_6047);
and U6592 (N_6592,N_6345,N_6272);
and U6593 (N_6593,N_6462,N_6106);
or U6594 (N_6594,N_6396,N_6487);
nand U6595 (N_6595,N_6497,N_6260);
nor U6596 (N_6596,N_6005,N_6280);
nor U6597 (N_6597,N_6379,N_6279);
nor U6598 (N_6598,N_6189,N_6271);
nand U6599 (N_6599,N_6324,N_6459);
nor U6600 (N_6600,N_6019,N_6378);
nor U6601 (N_6601,N_6176,N_6350);
xnor U6602 (N_6602,N_6060,N_6332);
nor U6603 (N_6603,N_6247,N_6074);
nor U6604 (N_6604,N_6377,N_6195);
xor U6605 (N_6605,N_6486,N_6415);
xnor U6606 (N_6606,N_6131,N_6251);
nand U6607 (N_6607,N_6055,N_6086);
nand U6608 (N_6608,N_6443,N_6307);
nor U6609 (N_6609,N_6453,N_6199);
or U6610 (N_6610,N_6050,N_6319);
or U6611 (N_6611,N_6304,N_6358);
and U6612 (N_6612,N_6361,N_6080);
xnor U6613 (N_6613,N_6145,N_6321);
and U6614 (N_6614,N_6278,N_6156);
or U6615 (N_6615,N_6458,N_6437);
and U6616 (N_6616,N_6427,N_6439);
nor U6617 (N_6617,N_6066,N_6018);
or U6618 (N_6618,N_6253,N_6419);
nand U6619 (N_6619,N_6264,N_6382);
and U6620 (N_6620,N_6367,N_6107);
nand U6621 (N_6621,N_6056,N_6483);
or U6622 (N_6622,N_6460,N_6398);
or U6623 (N_6623,N_6287,N_6065);
and U6624 (N_6624,N_6495,N_6226);
nand U6625 (N_6625,N_6130,N_6188);
xor U6626 (N_6626,N_6078,N_6243);
nand U6627 (N_6627,N_6275,N_6046);
and U6628 (N_6628,N_6472,N_6344);
xnor U6629 (N_6629,N_6204,N_6309);
nand U6630 (N_6630,N_6365,N_6372);
xnor U6631 (N_6631,N_6256,N_6348);
xnor U6632 (N_6632,N_6059,N_6469);
nand U6633 (N_6633,N_6168,N_6405);
nand U6634 (N_6634,N_6318,N_6095);
or U6635 (N_6635,N_6390,N_6200);
nand U6636 (N_6636,N_6136,N_6498);
xnor U6637 (N_6637,N_6132,N_6334);
nor U6638 (N_6638,N_6142,N_6157);
nand U6639 (N_6639,N_6210,N_6206);
nor U6640 (N_6640,N_6300,N_6119);
and U6641 (N_6641,N_6202,N_6429);
nand U6642 (N_6642,N_6400,N_6294);
xnor U6643 (N_6643,N_6036,N_6002);
nor U6644 (N_6644,N_6466,N_6313);
nor U6645 (N_6645,N_6178,N_6027);
nand U6646 (N_6646,N_6054,N_6402);
xor U6647 (N_6647,N_6051,N_6169);
and U6648 (N_6648,N_6161,N_6094);
nand U6649 (N_6649,N_6297,N_6022);
nand U6650 (N_6650,N_6299,N_6270);
and U6651 (N_6651,N_6135,N_6440);
or U6652 (N_6652,N_6305,N_6404);
nand U6653 (N_6653,N_6432,N_6336);
and U6654 (N_6654,N_6326,N_6325);
and U6655 (N_6655,N_6102,N_6024);
xor U6656 (N_6656,N_6217,N_6473);
nor U6657 (N_6657,N_6410,N_6455);
or U6658 (N_6658,N_6363,N_6381);
nand U6659 (N_6659,N_6212,N_6310);
nor U6660 (N_6660,N_6197,N_6370);
xnor U6661 (N_6661,N_6101,N_6230);
nor U6662 (N_6662,N_6008,N_6369);
xor U6663 (N_6663,N_6220,N_6100);
nor U6664 (N_6664,N_6108,N_6082);
nand U6665 (N_6665,N_6493,N_6006);
and U6666 (N_6666,N_6349,N_6250);
or U6667 (N_6667,N_6273,N_6103);
and U6668 (N_6668,N_6098,N_6441);
and U6669 (N_6669,N_6238,N_6353);
nor U6670 (N_6670,N_6084,N_6397);
nand U6671 (N_6671,N_6290,N_6029);
nand U6672 (N_6672,N_6069,N_6331);
xnor U6673 (N_6673,N_6033,N_6409);
nand U6674 (N_6674,N_6384,N_6414);
xnor U6675 (N_6675,N_6445,N_6057);
nor U6676 (N_6676,N_6030,N_6224);
xor U6677 (N_6677,N_6096,N_6463);
or U6678 (N_6678,N_6118,N_6420);
nand U6679 (N_6679,N_6352,N_6449);
or U6680 (N_6680,N_6001,N_6244);
nand U6681 (N_6681,N_6286,N_6302);
xor U6682 (N_6682,N_6298,N_6062);
or U6683 (N_6683,N_6407,N_6235);
nor U6684 (N_6684,N_6045,N_6053);
or U6685 (N_6685,N_6386,N_6335);
xor U6686 (N_6686,N_6281,N_6146);
nor U6687 (N_6687,N_6150,N_6052);
nand U6688 (N_6688,N_6147,N_6023);
xor U6689 (N_6689,N_6140,N_6114);
xor U6690 (N_6690,N_6236,N_6187);
and U6691 (N_6691,N_6434,N_6395);
and U6692 (N_6692,N_6044,N_6154);
nand U6693 (N_6693,N_6435,N_6259);
nand U6694 (N_6694,N_6026,N_6093);
nor U6695 (N_6695,N_6039,N_6013);
nor U6696 (N_6696,N_6252,N_6203);
and U6697 (N_6697,N_6191,N_6468);
nand U6698 (N_6698,N_6481,N_6356);
or U6699 (N_6699,N_6457,N_6166);
nand U6700 (N_6700,N_6436,N_6291);
nor U6701 (N_6701,N_6160,N_6282);
nand U6702 (N_6702,N_6482,N_6122);
xor U6703 (N_6703,N_6320,N_6423);
nand U6704 (N_6704,N_6164,N_6489);
xnor U6705 (N_6705,N_6133,N_6262);
xor U6706 (N_6706,N_6499,N_6099);
nand U6707 (N_6707,N_6153,N_6034);
nor U6708 (N_6708,N_6144,N_6218);
or U6709 (N_6709,N_6467,N_6035);
nand U6710 (N_6710,N_6012,N_6452);
nand U6711 (N_6711,N_6364,N_6448);
and U6712 (N_6712,N_6293,N_6339);
xor U6713 (N_6713,N_6343,N_6330);
and U6714 (N_6714,N_6374,N_6451);
nor U6715 (N_6715,N_6240,N_6109);
and U6716 (N_6716,N_6021,N_6171);
xnor U6717 (N_6717,N_6228,N_6058);
nand U6718 (N_6718,N_6274,N_6167);
nor U6719 (N_6719,N_6068,N_6387);
nand U6720 (N_6720,N_6480,N_6360);
nor U6721 (N_6721,N_6192,N_6322);
nand U6722 (N_6722,N_6428,N_6371);
nand U6723 (N_6723,N_6227,N_6088);
and U6724 (N_6724,N_6215,N_6375);
or U6725 (N_6725,N_6329,N_6391);
xor U6726 (N_6726,N_6340,N_6267);
and U6727 (N_6727,N_6292,N_6173);
nor U6728 (N_6728,N_6120,N_6392);
xor U6729 (N_6729,N_6234,N_6401);
nor U6730 (N_6730,N_6072,N_6306);
xor U6731 (N_6731,N_6137,N_6295);
xor U6732 (N_6732,N_6011,N_6461);
or U6733 (N_6733,N_6368,N_6328);
and U6734 (N_6734,N_6327,N_6073);
or U6735 (N_6735,N_6222,N_6124);
or U6736 (N_6736,N_6077,N_6446);
xnor U6737 (N_6737,N_6010,N_6110);
nor U6738 (N_6738,N_6040,N_6341);
or U6739 (N_6739,N_6141,N_6079);
xnor U6740 (N_6740,N_6242,N_6016);
nand U6741 (N_6741,N_6246,N_6134);
nor U6742 (N_6742,N_6406,N_6163);
and U6743 (N_6743,N_6366,N_6007);
or U6744 (N_6744,N_6111,N_6258);
nor U6745 (N_6745,N_6373,N_6385);
or U6746 (N_6746,N_6211,N_6416);
xor U6747 (N_6747,N_6426,N_6003);
xnor U6748 (N_6748,N_6477,N_6249);
and U6749 (N_6749,N_6128,N_6071);
nand U6750 (N_6750,N_6353,N_6279);
and U6751 (N_6751,N_6479,N_6227);
nand U6752 (N_6752,N_6299,N_6444);
or U6753 (N_6753,N_6332,N_6002);
nand U6754 (N_6754,N_6408,N_6436);
nor U6755 (N_6755,N_6153,N_6285);
and U6756 (N_6756,N_6199,N_6265);
or U6757 (N_6757,N_6446,N_6390);
nor U6758 (N_6758,N_6244,N_6352);
xnor U6759 (N_6759,N_6222,N_6397);
xor U6760 (N_6760,N_6437,N_6040);
and U6761 (N_6761,N_6318,N_6084);
and U6762 (N_6762,N_6464,N_6472);
xor U6763 (N_6763,N_6154,N_6056);
xnor U6764 (N_6764,N_6348,N_6361);
nor U6765 (N_6765,N_6366,N_6348);
xnor U6766 (N_6766,N_6460,N_6284);
xnor U6767 (N_6767,N_6325,N_6491);
or U6768 (N_6768,N_6278,N_6123);
and U6769 (N_6769,N_6150,N_6138);
nand U6770 (N_6770,N_6001,N_6260);
nor U6771 (N_6771,N_6193,N_6430);
nand U6772 (N_6772,N_6136,N_6231);
nand U6773 (N_6773,N_6456,N_6154);
nor U6774 (N_6774,N_6025,N_6080);
nor U6775 (N_6775,N_6372,N_6212);
xor U6776 (N_6776,N_6081,N_6234);
xnor U6777 (N_6777,N_6047,N_6285);
and U6778 (N_6778,N_6354,N_6056);
xnor U6779 (N_6779,N_6039,N_6148);
xnor U6780 (N_6780,N_6464,N_6017);
or U6781 (N_6781,N_6346,N_6399);
xnor U6782 (N_6782,N_6479,N_6371);
nor U6783 (N_6783,N_6437,N_6464);
nand U6784 (N_6784,N_6244,N_6008);
and U6785 (N_6785,N_6331,N_6240);
or U6786 (N_6786,N_6113,N_6180);
and U6787 (N_6787,N_6217,N_6372);
nor U6788 (N_6788,N_6380,N_6461);
xnor U6789 (N_6789,N_6458,N_6176);
or U6790 (N_6790,N_6273,N_6357);
and U6791 (N_6791,N_6327,N_6024);
nor U6792 (N_6792,N_6229,N_6359);
xnor U6793 (N_6793,N_6351,N_6156);
and U6794 (N_6794,N_6056,N_6319);
xnor U6795 (N_6795,N_6192,N_6318);
or U6796 (N_6796,N_6215,N_6454);
xnor U6797 (N_6797,N_6382,N_6149);
nand U6798 (N_6798,N_6066,N_6335);
nor U6799 (N_6799,N_6197,N_6302);
nand U6800 (N_6800,N_6080,N_6217);
and U6801 (N_6801,N_6490,N_6379);
nand U6802 (N_6802,N_6051,N_6195);
or U6803 (N_6803,N_6301,N_6069);
nor U6804 (N_6804,N_6279,N_6207);
or U6805 (N_6805,N_6437,N_6492);
or U6806 (N_6806,N_6164,N_6157);
and U6807 (N_6807,N_6028,N_6339);
xor U6808 (N_6808,N_6477,N_6371);
nor U6809 (N_6809,N_6499,N_6009);
and U6810 (N_6810,N_6048,N_6070);
nand U6811 (N_6811,N_6029,N_6054);
nor U6812 (N_6812,N_6117,N_6397);
or U6813 (N_6813,N_6464,N_6240);
or U6814 (N_6814,N_6028,N_6286);
or U6815 (N_6815,N_6293,N_6443);
and U6816 (N_6816,N_6318,N_6294);
or U6817 (N_6817,N_6023,N_6220);
nor U6818 (N_6818,N_6291,N_6267);
xor U6819 (N_6819,N_6369,N_6281);
and U6820 (N_6820,N_6180,N_6458);
and U6821 (N_6821,N_6382,N_6410);
and U6822 (N_6822,N_6066,N_6111);
or U6823 (N_6823,N_6210,N_6228);
nor U6824 (N_6824,N_6183,N_6480);
nor U6825 (N_6825,N_6186,N_6271);
nand U6826 (N_6826,N_6422,N_6178);
xnor U6827 (N_6827,N_6272,N_6316);
and U6828 (N_6828,N_6458,N_6358);
and U6829 (N_6829,N_6182,N_6227);
nand U6830 (N_6830,N_6322,N_6142);
nand U6831 (N_6831,N_6436,N_6287);
nor U6832 (N_6832,N_6472,N_6409);
nor U6833 (N_6833,N_6077,N_6107);
nand U6834 (N_6834,N_6207,N_6433);
or U6835 (N_6835,N_6340,N_6311);
and U6836 (N_6836,N_6090,N_6096);
or U6837 (N_6837,N_6360,N_6258);
xnor U6838 (N_6838,N_6237,N_6390);
or U6839 (N_6839,N_6005,N_6282);
and U6840 (N_6840,N_6405,N_6154);
nand U6841 (N_6841,N_6013,N_6331);
nand U6842 (N_6842,N_6406,N_6442);
xor U6843 (N_6843,N_6077,N_6335);
nand U6844 (N_6844,N_6188,N_6236);
nand U6845 (N_6845,N_6102,N_6275);
or U6846 (N_6846,N_6326,N_6110);
nand U6847 (N_6847,N_6335,N_6268);
xnor U6848 (N_6848,N_6102,N_6422);
and U6849 (N_6849,N_6136,N_6333);
and U6850 (N_6850,N_6307,N_6451);
nand U6851 (N_6851,N_6272,N_6101);
nand U6852 (N_6852,N_6065,N_6265);
or U6853 (N_6853,N_6111,N_6354);
xor U6854 (N_6854,N_6306,N_6019);
and U6855 (N_6855,N_6032,N_6352);
nand U6856 (N_6856,N_6356,N_6136);
and U6857 (N_6857,N_6209,N_6327);
nand U6858 (N_6858,N_6043,N_6181);
or U6859 (N_6859,N_6332,N_6134);
nand U6860 (N_6860,N_6398,N_6353);
nand U6861 (N_6861,N_6179,N_6225);
nand U6862 (N_6862,N_6300,N_6388);
and U6863 (N_6863,N_6236,N_6329);
xnor U6864 (N_6864,N_6321,N_6107);
xnor U6865 (N_6865,N_6309,N_6092);
xnor U6866 (N_6866,N_6183,N_6483);
or U6867 (N_6867,N_6283,N_6190);
and U6868 (N_6868,N_6418,N_6056);
or U6869 (N_6869,N_6119,N_6105);
or U6870 (N_6870,N_6435,N_6395);
and U6871 (N_6871,N_6172,N_6026);
xor U6872 (N_6872,N_6256,N_6115);
and U6873 (N_6873,N_6133,N_6013);
and U6874 (N_6874,N_6333,N_6190);
and U6875 (N_6875,N_6271,N_6372);
or U6876 (N_6876,N_6274,N_6472);
xnor U6877 (N_6877,N_6145,N_6369);
nand U6878 (N_6878,N_6221,N_6203);
xnor U6879 (N_6879,N_6393,N_6264);
or U6880 (N_6880,N_6126,N_6476);
nor U6881 (N_6881,N_6405,N_6355);
or U6882 (N_6882,N_6301,N_6055);
nor U6883 (N_6883,N_6368,N_6354);
nand U6884 (N_6884,N_6009,N_6043);
nor U6885 (N_6885,N_6130,N_6238);
nor U6886 (N_6886,N_6251,N_6221);
nand U6887 (N_6887,N_6015,N_6314);
and U6888 (N_6888,N_6014,N_6052);
nand U6889 (N_6889,N_6013,N_6089);
nand U6890 (N_6890,N_6209,N_6301);
xor U6891 (N_6891,N_6279,N_6419);
nor U6892 (N_6892,N_6225,N_6242);
or U6893 (N_6893,N_6381,N_6334);
nor U6894 (N_6894,N_6035,N_6444);
xnor U6895 (N_6895,N_6147,N_6446);
or U6896 (N_6896,N_6330,N_6423);
xor U6897 (N_6897,N_6034,N_6167);
xnor U6898 (N_6898,N_6213,N_6271);
nor U6899 (N_6899,N_6118,N_6404);
xor U6900 (N_6900,N_6255,N_6389);
xor U6901 (N_6901,N_6428,N_6193);
or U6902 (N_6902,N_6065,N_6091);
nor U6903 (N_6903,N_6196,N_6449);
nand U6904 (N_6904,N_6284,N_6183);
and U6905 (N_6905,N_6099,N_6149);
xnor U6906 (N_6906,N_6323,N_6171);
or U6907 (N_6907,N_6417,N_6234);
and U6908 (N_6908,N_6450,N_6023);
and U6909 (N_6909,N_6396,N_6313);
xnor U6910 (N_6910,N_6110,N_6201);
xor U6911 (N_6911,N_6131,N_6201);
xor U6912 (N_6912,N_6193,N_6490);
nand U6913 (N_6913,N_6149,N_6102);
nand U6914 (N_6914,N_6154,N_6252);
or U6915 (N_6915,N_6054,N_6310);
nor U6916 (N_6916,N_6145,N_6214);
nor U6917 (N_6917,N_6168,N_6199);
xnor U6918 (N_6918,N_6112,N_6409);
nor U6919 (N_6919,N_6485,N_6476);
or U6920 (N_6920,N_6442,N_6423);
xnor U6921 (N_6921,N_6044,N_6220);
nor U6922 (N_6922,N_6468,N_6424);
or U6923 (N_6923,N_6065,N_6388);
or U6924 (N_6924,N_6002,N_6194);
xnor U6925 (N_6925,N_6031,N_6386);
or U6926 (N_6926,N_6073,N_6395);
or U6927 (N_6927,N_6426,N_6102);
or U6928 (N_6928,N_6348,N_6338);
xor U6929 (N_6929,N_6374,N_6182);
or U6930 (N_6930,N_6186,N_6220);
and U6931 (N_6931,N_6214,N_6123);
and U6932 (N_6932,N_6086,N_6373);
nor U6933 (N_6933,N_6304,N_6103);
xnor U6934 (N_6934,N_6427,N_6031);
nor U6935 (N_6935,N_6199,N_6478);
and U6936 (N_6936,N_6157,N_6369);
nor U6937 (N_6937,N_6323,N_6082);
nand U6938 (N_6938,N_6076,N_6386);
and U6939 (N_6939,N_6281,N_6115);
nor U6940 (N_6940,N_6183,N_6217);
and U6941 (N_6941,N_6026,N_6028);
nand U6942 (N_6942,N_6237,N_6439);
xnor U6943 (N_6943,N_6428,N_6341);
or U6944 (N_6944,N_6169,N_6211);
and U6945 (N_6945,N_6472,N_6186);
xnor U6946 (N_6946,N_6246,N_6048);
and U6947 (N_6947,N_6340,N_6208);
nand U6948 (N_6948,N_6129,N_6304);
nand U6949 (N_6949,N_6279,N_6335);
xor U6950 (N_6950,N_6136,N_6266);
and U6951 (N_6951,N_6014,N_6200);
and U6952 (N_6952,N_6296,N_6447);
nand U6953 (N_6953,N_6235,N_6300);
nor U6954 (N_6954,N_6074,N_6443);
or U6955 (N_6955,N_6055,N_6337);
nand U6956 (N_6956,N_6450,N_6420);
nand U6957 (N_6957,N_6499,N_6401);
nor U6958 (N_6958,N_6254,N_6051);
xnor U6959 (N_6959,N_6240,N_6077);
xnor U6960 (N_6960,N_6040,N_6201);
nand U6961 (N_6961,N_6030,N_6256);
xnor U6962 (N_6962,N_6226,N_6028);
nand U6963 (N_6963,N_6003,N_6205);
xnor U6964 (N_6964,N_6002,N_6150);
and U6965 (N_6965,N_6303,N_6174);
nor U6966 (N_6966,N_6339,N_6203);
nor U6967 (N_6967,N_6281,N_6062);
or U6968 (N_6968,N_6324,N_6232);
and U6969 (N_6969,N_6145,N_6051);
or U6970 (N_6970,N_6269,N_6030);
or U6971 (N_6971,N_6182,N_6296);
nor U6972 (N_6972,N_6433,N_6132);
or U6973 (N_6973,N_6339,N_6291);
xnor U6974 (N_6974,N_6432,N_6115);
xor U6975 (N_6975,N_6270,N_6410);
nand U6976 (N_6976,N_6042,N_6082);
xor U6977 (N_6977,N_6492,N_6052);
or U6978 (N_6978,N_6465,N_6415);
nand U6979 (N_6979,N_6342,N_6146);
nor U6980 (N_6980,N_6069,N_6286);
nand U6981 (N_6981,N_6421,N_6264);
and U6982 (N_6982,N_6093,N_6259);
nor U6983 (N_6983,N_6343,N_6470);
or U6984 (N_6984,N_6082,N_6448);
or U6985 (N_6985,N_6163,N_6381);
xor U6986 (N_6986,N_6416,N_6235);
nand U6987 (N_6987,N_6229,N_6417);
or U6988 (N_6988,N_6388,N_6169);
and U6989 (N_6989,N_6133,N_6102);
or U6990 (N_6990,N_6212,N_6421);
and U6991 (N_6991,N_6365,N_6333);
nand U6992 (N_6992,N_6207,N_6055);
xor U6993 (N_6993,N_6330,N_6123);
xor U6994 (N_6994,N_6143,N_6392);
and U6995 (N_6995,N_6192,N_6211);
nand U6996 (N_6996,N_6000,N_6088);
or U6997 (N_6997,N_6499,N_6295);
nor U6998 (N_6998,N_6419,N_6210);
nand U6999 (N_6999,N_6350,N_6299);
xor U7000 (N_7000,N_6805,N_6792);
xor U7001 (N_7001,N_6841,N_6583);
nand U7002 (N_7002,N_6548,N_6505);
or U7003 (N_7003,N_6634,N_6659);
or U7004 (N_7004,N_6594,N_6749);
nor U7005 (N_7005,N_6531,N_6510);
nor U7006 (N_7006,N_6507,N_6798);
xnor U7007 (N_7007,N_6752,N_6557);
or U7008 (N_7008,N_6588,N_6703);
and U7009 (N_7009,N_6830,N_6866);
and U7010 (N_7010,N_6738,N_6618);
or U7011 (N_7011,N_6886,N_6576);
nand U7012 (N_7012,N_6808,N_6916);
or U7013 (N_7013,N_6532,N_6791);
xnor U7014 (N_7014,N_6735,N_6893);
nor U7015 (N_7015,N_6944,N_6683);
or U7016 (N_7016,N_6556,N_6905);
nand U7017 (N_7017,N_6954,N_6697);
nor U7018 (N_7018,N_6915,N_6607);
xor U7019 (N_7019,N_6904,N_6721);
xnor U7020 (N_7020,N_6845,N_6843);
or U7021 (N_7021,N_6834,N_6722);
or U7022 (N_7022,N_6636,N_6629);
or U7023 (N_7023,N_6577,N_6995);
nor U7024 (N_7024,N_6760,N_6914);
or U7025 (N_7025,N_6651,N_6641);
and U7026 (N_7026,N_6762,N_6533);
nor U7027 (N_7027,N_6779,N_6974);
nor U7028 (N_7028,N_6997,N_6820);
nor U7029 (N_7029,N_6906,N_6608);
nand U7030 (N_7030,N_6564,N_6580);
xnor U7031 (N_7031,N_6940,N_6751);
nand U7032 (N_7032,N_6931,N_6787);
nand U7033 (N_7033,N_6840,N_6935);
or U7034 (N_7034,N_6753,N_6927);
nor U7035 (N_7035,N_6536,N_6986);
and U7036 (N_7036,N_6695,N_6611);
nand U7037 (N_7037,N_6797,N_6965);
xor U7038 (N_7038,N_6569,N_6833);
and U7039 (N_7039,N_6793,N_6736);
nand U7040 (N_7040,N_6534,N_6757);
or U7041 (N_7041,N_6850,N_6975);
or U7042 (N_7042,N_6624,N_6827);
nand U7043 (N_7043,N_6657,N_6910);
nor U7044 (N_7044,N_6939,N_6720);
nor U7045 (N_7045,N_6933,N_6889);
nor U7046 (N_7046,N_6780,N_6597);
xor U7047 (N_7047,N_6920,N_6728);
nor U7048 (N_7048,N_6957,N_6691);
xor U7049 (N_7049,N_6922,N_6984);
and U7050 (N_7050,N_6681,N_6772);
xnor U7051 (N_7051,N_6699,N_6966);
xor U7052 (N_7052,N_6616,N_6578);
nand U7053 (N_7053,N_6924,N_6590);
nor U7054 (N_7054,N_6609,N_6891);
nor U7055 (N_7055,N_6782,N_6712);
xor U7056 (N_7056,N_6842,N_6989);
xor U7057 (N_7057,N_6513,N_6917);
xor U7058 (N_7058,N_6709,N_6731);
and U7059 (N_7059,N_6803,N_6542);
nand U7060 (N_7060,N_6835,N_6558);
xor U7061 (N_7061,N_6667,N_6584);
or U7062 (N_7062,N_6852,N_6888);
and U7063 (N_7063,N_6781,N_6956);
nor U7064 (N_7064,N_6998,N_6932);
nand U7065 (N_7065,N_6826,N_6620);
nor U7066 (N_7066,N_6586,N_6612);
and U7067 (N_7067,N_6867,N_6689);
xnor U7068 (N_7068,N_6639,N_6959);
nand U7069 (N_7069,N_6719,N_6662);
and U7070 (N_7070,N_6815,N_6605);
nor U7071 (N_7071,N_6771,N_6885);
nor U7072 (N_7072,N_6770,N_6761);
nor U7073 (N_7073,N_6766,N_6972);
xor U7074 (N_7074,N_6942,N_6633);
xor U7075 (N_7075,N_6784,N_6894);
or U7076 (N_7076,N_6858,N_6664);
xnor U7077 (N_7077,N_6809,N_6623);
and U7078 (N_7078,N_6860,N_6692);
or U7079 (N_7079,N_6748,N_6816);
and U7080 (N_7080,N_6747,N_6796);
nor U7081 (N_7081,N_6515,N_6979);
and U7082 (N_7082,N_6746,N_6890);
nand U7083 (N_7083,N_6951,N_6551);
nor U7084 (N_7084,N_6876,N_6754);
and U7085 (N_7085,N_6582,N_6530);
or U7086 (N_7086,N_6725,N_6824);
and U7087 (N_7087,N_6865,N_6898);
nor U7088 (N_7088,N_6658,N_6861);
and U7089 (N_7089,N_6648,N_6755);
nand U7090 (N_7090,N_6879,N_6678);
xnor U7091 (N_7091,N_6570,N_6896);
nor U7092 (N_7092,N_6560,N_6643);
nand U7093 (N_7093,N_6717,N_6537);
xor U7094 (N_7094,N_6546,N_6887);
xnor U7095 (N_7095,N_6656,N_6870);
and U7096 (N_7096,N_6819,N_6601);
and U7097 (N_7097,N_6644,N_6529);
nor U7098 (N_7098,N_6660,N_6615);
xor U7099 (N_7099,N_6523,N_6701);
or U7100 (N_7100,N_6929,N_6535);
nor U7101 (N_7101,N_6555,N_6540);
and U7102 (N_7102,N_6527,N_6726);
nor U7103 (N_7103,N_6925,N_6948);
nand U7104 (N_7104,N_6964,N_6987);
nor U7105 (N_7105,N_6848,N_6702);
nor U7106 (N_7106,N_6985,N_6983);
or U7107 (N_7107,N_6742,N_6961);
or U7108 (N_7108,N_6778,N_6617);
and U7109 (N_7109,N_6730,N_6967);
or U7110 (N_7110,N_6705,N_6642);
or U7111 (N_7111,N_6875,N_6621);
and U7112 (N_7112,N_6574,N_6996);
and U7113 (N_7113,N_6677,N_6775);
or U7114 (N_7114,N_6562,N_6599);
xnor U7115 (N_7115,N_6631,N_6550);
nand U7116 (N_7116,N_6650,N_6579);
xnor U7117 (N_7117,N_6941,N_6517);
nor U7118 (N_7118,N_6810,N_6963);
nor U7119 (N_7119,N_6874,N_6718);
xnor U7120 (N_7120,N_6990,N_6706);
nand U7121 (N_7121,N_6665,N_6981);
and U7122 (N_7122,N_6679,N_6575);
nor U7123 (N_7123,N_6958,N_6856);
nor U7124 (N_7124,N_6902,N_6673);
nand U7125 (N_7125,N_6592,N_6831);
or U7126 (N_7126,N_6855,N_6669);
and U7127 (N_7127,N_6559,N_6571);
or U7128 (N_7128,N_6758,N_6945);
or U7129 (N_7129,N_6960,N_6980);
and U7130 (N_7130,N_6812,N_6973);
or U7131 (N_7131,N_6813,N_6976);
or U7132 (N_7132,N_6610,N_6847);
nor U7133 (N_7133,N_6955,N_6614);
xor U7134 (N_7134,N_6817,N_6968);
nor U7135 (N_7135,N_6868,N_6788);
or U7136 (N_7136,N_6506,N_6789);
nor U7137 (N_7137,N_6880,N_6918);
nor U7138 (N_7138,N_6926,N_6737);
and U7139 (N_7139,N_6518,N_6892);
xnor U7140 (N_7140,N_6829,N_6999);
or U7141 (N_7141,N_6707,N_6836);
xnor U7142 (N_7142,N_6794,N_6934);
xor U7143 (N_7143,N_6991,N_6774);
nand U7144 (N_7144,N_6741,N_6723);
or U7145 (N_7145,N_6943,N_6837);
and U7146 (N_7146,N_6923,N_6688);
and U7147 (N_7147,N_6994,N_6652);
xnor U7148 (N_7148,N_6849,N_6514);
or U7149 (N_7149,N_6853,N_6978);
and U7150 (N_7150,N_6696,N_6949);
nand U7151 (N_7151,N_6568,N_6710);
nand U7152 (N_7152,N_6711,N_6521);
xnor U7153 (N_7153,N_6786,N_6937);
xnor U7154 (N_7154,N_6676,N_6606);
or U7155 (N_7155,N_6903,N_6862);
nor U7156 (N_7156,N_6502,N_6524);
or U7157 (N_7157,N_6908,N_6638);
or U7158 (N_7158,N_6553,N_6622);
nor U7159 (N_7159,N_6732,N_6763);
nand U7160 (N_7160,N_6971,N_6508);
and U7161 (N_7161,N_6544,N_6743);
or U7162 (N_7162,N_6635,N_6729);
nand U7163 (N_7163,N_6704,N_6988);
and U7164 (N_7164,N_6807,N_6670);
xnor U7165 (N_7165,N_6854,N_6977);
nand U7166 (N_7166,N_6646,N_6897);
or U7167 (N_7167,N_6613,N_6566);
and U7168 (N_7168,N_6627,N_6993);
xor U7169 (N_7169,N_6538,N_6581);
or U7170 (N_7170,N_6733,N_6859);
nand U7171 (N_7171,N_6822,N_6572);
xor U7172 (N_7172,N_6804,N_6686);
and U7173 (N_7173,N_6698,N_6844);
nor U7174 (N_7174,N_6913,N_6509);
xnor U7175 (N_7175,N_6640,N_6565);
or U7176 (N_7176,N_6500,N_6992);
or U7177 (N_7177,N_6773,N_6519);
xor U7178 (N_7178,N_6846,N_6740);
nand U7179 (N_7179,N_6928,N_6541);
or U7180 (N_7180,N_6596,N_6525);
nand U7181 (N_7181,N_6573,N_6600);
or U7182 (N_7182,N_6839,N_6739);
and U7183 (N_7183,N_6632,N_6595);
nor U7184 (N_7184,N_6953,N_6900);
nand U7185 (N_7185,N_6593,N_6828);
and U7186 (N_7186,N_6547,N_6589);
or U7187 (N_7187,N_6895,N_6666);
nor U7188 (N_7188,N_6759,N_6806);
nor U7189 (N_7189,N_6511,N_6545);
nand U7190 (N_7190,N_6869,N_6838);
nor U7191 (N_7191,N_6832,N_6554);
nor U7192 (N_7192,N_6795,N_6653);
nor U7193 (N_7193,N_6938,N_6682);
and U7194 (N_7194,N_6672,N_6715);
and U7195 (N_7195,N_6619,N_6982);
nor U7196 (N_7196,N_6814,N_6700);
nand U7197 (N_7197,N_6713,N_6800);
or U7198 (N_7198,N_6877,N_6745);
xor U7199 (N_7199,N_6790,N_6921);
and U7200 (N_7200,N_6919,N_6539);
xnor U7201 (N_7201,N_6684,N_6750);
nand U7202 (N_7202,N_6777,N_6716);
xor U7203 (N_7203,N_6825,N_6675);
and U7204 (N_7204,N_6645,N_6690);
xnor U7205 (N_7205,N_6783,N_6680);
nand U7206 (N_7206,N_6785,N_6907);
xor U7207 (N_7207,N_6901,N_6857);
and U7208 (N_7208,N_6663,N_6734);
and U7209 (N_7209,N_6637,N_6911);
or U7210 (N_7210,N_6687,N_6563);
and U7211 (N_7211,N_6764,N_6811);
xor U7212 (N_7212,N_6881,N_6899);
xor U7213 (N_7213,N_6501,N_6912);
xnor U7214 (N_7214,N_6661,N_6882);
and U7215 (N_7215,N_6604,N_6685);
nor U7216 (N_7216,N_6872,N_6946);
and U7217 (N_7217,N_6674,N_6516);
nand U7218 (N_7218,N_6543,N_6668);
nand U7219 (N_7219,N_6503,N_6756);
nand U7220 (N_7220,N_6909,N_6823);
xnor U7221 (N_7221,N_6873,N_6724);
nor U7222 (N_7222,N_6930,N_6818);
xnor U7223 (N_7223,N_6522,N_6799);
nand U7224 (N_7224,N_6727,N_6626);
and U7225 (N_7225,N_6694,N_6768);
or U7226 (N_7226,N_6628,N_6567);
nand U7227 (N_7227,N_6671,N_6655);
or U7228 (N_7228,N_6630,N_6647);
xnor U7229 (N_7229,N_6871,N_6821);
and U7230 (N_7230,N_6962,N_6625);
xor U7231 (N_7231,N_6765,N_6649);
nand U7232 (N_7232,N_6654,N_6602);
nand U7233 (N_7233,N_6802,N_6950);
nor U7234 (N_7234,N_6520,N_6512);
or U7235 (N_7235,N_6776,N_6526);
nor U7236 (N_7236,N_6744,N_6598);
nor U7237 (N_7237,N_6603,N_6883);
nand U7238 (N_7238,N_6936,N_6801);
nand U7239 (N_7239,N_6561,N_6714);
xor U7240 (N_7240,N_6851,N_6693);
nand U7241 (N_7241,N_6767,N_6947);
nor U7242 (N_7242,N_6587,N_6504);
and U7243 (N_7243,N_6549,N_6708);
nand U7244 (N_7244,N_6878,N_6591);
nand U7245 (N_7245,N_6552,N_6969);
nor U7246 (N_7246,N_6863,N_6952);
nand U7247 (N_7247,N_6585,N_6970);
nor U7248 (N_7248,N_6769,N_6528);
xnor U7249 (N_7249,N_6864,N_6884);
xnor U7250 (N_7250,N_6756,N_6812);
and U7251 (N_7251,N_6524,N_6662);
xor U7252 (N_7252,N_6535,N_6526);
nor U7253 (N_7253,N_6515,N_6626);
xnor U7254 (N_7254,N_6527,N_6720);
nor U7255 (N_7255,N_6506,N_6990);
and U7256 (N_7256,N_6803,N_6779);
and U7257 (N_7257,N_6834,N_6707);
xnor U7258 (N_7258,N_6954,N_6925);
or U7259 (N_7259,N_6655,N_6738);
nor U7260 (N_7260,N_6833,N_6551);
nand U7261 (N_7261,N_6621,N_6598);
xnor U7262 (N_7262,N_6517,N_6976);
and U7263 (N_7263,N_6718,N_6985);
or U7264 (N_7264,N_6784,N_6852);
nand U7265 (N_7265,N_6839,N_6958);
xnor U7266 (N_7266,N_6752,N_6842);
xor U7267 (N_7267,N_6716,N_6957);
nand U7268 (N_7268,N_6552,N_6860);
xor U7269 (N_7269,N_6592,N_6679);
nor U7270 (N_7270,N_6930,N_6781);
or U7271 (N_7271,N_6570,N_6909);
and U7272 (N_7272,N_6547,N_6848);
nand U7273 (N_7273,N_6786,N_6866);
nor U7274 (N_7274,N_6866,N_6624);
or U7275 (N_7275,N_6727,N_6894);
xor U7276 (N_7276,N_6736,N_6569);
nor U7277 (N_7277,N_6544,N_6954);
xnor U7278 (N_7278,N_6804,N_6671);
nor U7279 (N_7279,N_6570,N_6821);
and U7280 (N_7280,N_6990,N_6952);
xor U7281 (N_7281,N_6533,N_6821);
nand U7282 (N_7282,N_6993,N_6837);
xnor U7283 (N_7283,N_6591,N_6585);
nor U7284 (N_7284,N_6633,N_6673);
nor U7285 (N_7285,N_6631,N_6861);
or U7286 (N_7286,N_6923,N_6844);
xnor U7287 (N_7287,N_6805,N_6625);
nor U7288 (N_7288,N_6826,N_6518);
and U7289 (N_7289,N_6944,N_6941);
or U7290 (N_7290,N_6516,N_6910);
or U7291 (N_7291,N_6807,N_6554);
xor U7292 (N_7292,N_6982,N_6770);
xnor U7293 (N_7293,N_6674,N_6871);
and U7294 (N_7294,N_6745,N_6843);
xor U7295 (N_7295,N_6982,N_6895);
and U7296 (N_7296,N_6830,N_6724);
nand U7297 (N_7297,N_6634,N_6966);
xor U7298 (N_7298,N_6645,N_6879);
or U7299 (N_7299,N_6518,N_6616);
nand U7300 (N_7300,N_6743,N_6511);
xnor U7301 (N_7301,N_6826,N_6554);
and U7302 (N_7302,N_6958,N_6930);
nor U7303 (N_7303,N_6673,N_6519);
nor U7304 (N_7304,N_6975,N_6764);
nor U7305 (N_7305,N_6879,N_6546);
xnor U7306 (N_7306,N_6934,N_6918);
nand U7307 (N_7307,N_6751,N_6733);
or U7308 (N_7308,N_6897,N_6606);
nor U7309 (N_7309,N_6741,N_6658);
nor U7310 (N_7310,N_6765,N_6530);
and U7311 (N_7311,N_6706,N_6861);
nand U7312 (N_7312,N_6642,N_6963);
or U7313 (N_7313,N_6875,N_6943);
and U7314 (N_7314,N_6920,N_6801);
xor U7315 (N_7315,N_6862,N_6873);
and U7316 (N_7316,N_6559,N_6871);
or U7317 (N_7317,N_6765,N_6720);
or U7318 (N_7318,N_6723,N_6780);
and U7319 (N_7319,N_6877,N_6953);
and U7320 (N_7320,N_6600,N_6554);
nor U7321 (N_7321,N_6530,N_6588);
and U7322 (N_7322,N_6811,N_6591);
nand U7323 (N_7323,N_6745,N_6524);
xor U7324 (N_7324,N_6801,N_6652);
and U7325 (N_7325,N_6815,N_6560);
nand U7326 (N_7326,N_6825,N_6676);
and U7327 (N_7327,N_6509,N_6688);
nor U7328 (N_7328,N_6987,N_6902);
nand U7329 (N_7329,N_6941,N_6804);
nor U7330 (N_7330,N_6814,N_6997);
nand U7331 (N_7331,N_6815,N_6859);
xnor U7332 (N_7332,N_6665,N_6925);
nor U7333 (N_7333,N_6993,N_6804);
nor U7334 (N_7334,N_6615,N_6650);
nor U7335 (N_7335,N_6797,N_6633);
nor U7336 (N_7336,N_6672,N_6589);
and U7337 (N_7337,N_6825,N_6682);
and U7338 (N_7338,N_6748,N_6864);
and U7339 (N_7339,N_6719,N_6553);
nor U7340 (N_7340,N_6891,N_6872);
nor U7341 (N_7341,N_6527,N_6535);
nand U7342 (N_7342,N_6527,N_6941);
nor U7343 (N_7343,N_6629,N_6727);
or U7344 (N_7344,N_6729,N_6971);
nor U7345 (N_7345,N_6623,N_6731);
nand U7346 (N_7346,N_6927,N_6969);
xor U7347 (N_7347,N_6561,N_6509);
and U7348 (N_7348,N_6902,N_6543);
and U7349 (N_7349,N_6701,N_6510);
nand U7350 (N_7350,N_6561,N_6758);
nand U7351 (N_7351,N_6594,N_6581);
xnor U7352 (N_7352,N_6514,N_6917);
and U7353 (N_7353,N_6865,N_6509);
or U7354 (N_7354,N_6900,N_6955);
or U7355 (N_7355,N_6738,N_6894);
xnor U7356 (N_7356,N_6739,N_6933);
nand U7357 (N_7357,N_6544,N_6706);
and U7358 (N_7358,N_6565,N_6730);
nand U7359 (N_7359,N_6789,N_6866);
and U7360 (N_7360,N_6820,N_6756);
xor U7361 (N_7361,N_6840,N_6633);
nand U7362 (N_7362,N_6810,N_6506);
or U7363 (N_7363,N_6901,N_6536);
nand U7364 (N_7364,N_6662,N_6800);
and U7365 (N_7365,N_6785,N_6776);
and U7366 (N_7366,N_6604,N_6599);
xor U7367 (N_7367,N_6864,N_6615);
or U7368 (N_7368,N_6713,N_6870);
and U7369 (N_7369,N_6700,N_6568);
and U7370 (N_7370,N_6760,N_6530);
and U7371 (N_7371,N_6919,N_6735);
xor U7372 (N_7372,N_6831,N_6840);
xnor U7373 (N_7373,N_6624,N_6819);
nand U7374 (N_7374,N_6913,N_6948);
and U7375 (N_7375,N_6537,N_6749);
nand U7376 (N_7376,N_6527,N_6891);
nor U7377 (N_7377,N_6616,N_6530);
or U7378 (N_7378,N_6762,N_6692);
or U7379 (N_7379,N_6604,N_6876);
and U7380 (N_7380,N_6793,N_6544);
and U7381 (N_7381,N_6707,N_6525);
xor U7382 (N_7382,N_6936,N_6508);
xor U7383 (N_7383,N_6615,N_6666);
and U7384 (N_7384,N_6985,N_6541);
or U7385 (N_7385,N_6628,N_6996);
xor U7386 (N_7386,N_6518,N_6756);
and U7387 (N_7387,N_6510,N_6629);
and U7388 (N_7388,N_6963,N_6705);
nand U7389 (N_7389,N_6671,N_6688);
xor U7390 (N_7390,N_6833,N_6912);
or U7391 (N_7391,N_6766,N_6784);
nor U7392 (N_7392,N_6960,N_6635);
nor U7393 (N_7393,N_6679,N_6644);
nand U7394 (N_7394,N_6792,N_6958);
or U7395 (N_7395,N_6701,N_6663);
xor U7396 (N_7396,N_6924,N_6943);
nand U7397 (N_7397,N_6965,N_6520);
nand U7398 (N_7398,N_6908,N_6940);
or U7399 (N_7399,N_6986,N_6522);
or U7400 (N_7400,N_6547,N_6817);
xor U7401 (N_7401,N_6752,N_6652);
and U7402 (N_7402,N_6856,N_6825);
and U7403 (N_7403,N_6809,N_6958);
or U7404 (N_7404,N_6595,N_6801);
and U7405 (N_7405,N_6856,N_6812);
nand U7406 (N_7406,N_6551,N_6811);
nand U7407 (N_7407,N_6637,N_6688);
nor U7408 (N_7408,N_6713,N_6685);
nor U7409 (N_7409,N_6925,N_6801);
nor U7410 (N_7410,N_6835,N_6633);
nor U7411 (N_7411,N_6900,N_6628);
nor U7412 (N_7412,N_6780,N_6979);
or U7413 (N_7413,N_6911,N_6627);
nand U7414 (N_7414,N_6791,N_6629);
xor U7415 (N_7415,N_6958,N_6890);
nor U7416 (N_7416,N_6594,N_6683);
nor U7417 (N_7417,N_6545,N_6924);
or U7418 (N_7418,N_6830,N_6799);
nand U7419 (N_7419,N_6929,N_6840);
and U7420 (N_7420,N_6900,N_6712);
and U7421 (N_7421,N_6553,N_6748);
xor U7422 (N_7422,N_6953,N_6898);
and U7423 (N_7423,N_6658,N_6724);
or U7424 (N_7424,N_6787,N_6797);
nor U7425 (N_7425,N_6754,N_6584);
or U7426 (N_7426,N_6504,N_6868);
nand U7427 (N_7427,N_6993,N_6924);
nor U7428 (N_7428,N_6611,N_6824);
xor U7429 (N_7429,N_6652,N_6535);
nand U7430 (N_7430,N_6879,N_6538);
and U7431 (N_7431,N_6770,N_6851);
or U7432 (N_7432,N_6837,N_6529);
nor U7433 (N_7433,N_6775,N_6560);
xnor U7434 (N_7434,N_6821,N_6597);
or U7435 (N_7435,N_6685,N_6839);
nand U7436 (N_7436,N_6589,N_6978);
nor U7437 (N_7437,N_6624,N_6983);
nand U7438 (N_7438,N_6535,N_6543);
nand U7439 (N_7439,N_6743,N_6947);
nand U7440 (N_7440,N_6855,N_6872);
nand U7441 (N_7441,N_6978,N_6719);
and U7442 (N_7442,N_6788,N_6937);
nand U7443 (N_7443,N_6585,N_6871);
xor U7444 (N_7444,N_6702,N_6852);
and U7445 (N_7445,N_6897,N_6766);
or U7446 (N_7446,N_6816,N_6513);
nand U7447 (N_7447,N_6706,N_6899);
and U7448 (N_7448,N_6753,N_6669);
nand U7449 (N_7449,N_6514,N_6958);
nor U7450 (N_7450,N_6956,N_6728);
nor U7451 (N_7451,N_6603,N_6833);
or U7452 (N_7452,N_6944,N_6737);
nand U7453 (N_7453,N_6622,N_6826);
or U7454 (N_7454,N_6733,N_6787);
xnor U7455 (N_7455,N_6902,N_6733);
and U7456 (N_7456,N_6764,N_6831);
xor U7457 (N_7457,N_6525,N_6640);
nor U7458 (N_7458,N_6678,N_6712);
and U7459 (N_7459,N_6729,N_6693);
nand U7460 (N_7460,N_6825,N_6795);
nor U7461 (N_7461,N_6673,N_6977);
nand U7462 (N_7462,N_6974,N_6595);
or U7463 (N_7463,N_6512,N_6633);
nand U7464 (N_7464,N_6713,N_6933);
and U7465 (N_7465,N_6673,N_6663);
nand U7466 (N_7466,N_6791,N_6887);
or U7467 (N_7467,N_6501,N_6745);
nand U7468 (N_7468,N_6581,N_6615);
nor U7469 (N_7469,N_6592,N_6529);
nand U7470 (N_7470,N_6634,N_6711);
xor U7471 (N_7471,N_6898,N_6774);
nor U7472 (N_7472,N_6630,N_6785);
nor U7473 (N_7473,N_6909,N_6505);
nor U7474 (N_7474,N_6554,N_6783);
xnor U7475 (N_7475,N_6584,N_6890);
xnor U7476 (N_7476,N_6771,N_6615);
and U7477 (N_7477,N_6822,N_6543);
or U7478 (N_7478,N_6897,N_6927);
nand U7479 (N_7479,N_6854,N_6567);
and U7480 (N_7480,N_6573,N_6895);
or U7481 (N_7481,N_6817,N_6915);
nor U7482 (N_7482,N_6537,N_6775);
xor U7483 (N_7483,N_6780,N_6940);
xnor U7484 (N_7484,N_6702,N_6584);
nor U7485 (N_7485,N_6753,N_6748);
xor U7486 (N_7486,N_6929,N_6761);
nand U7487 (N_7487,N_6552,N_6631);
and U7488 (N_7488,N_6706,N_6963);
nand U7489 (N_7489,N_6538,N_6803);
nand U7490 (N_7490,N_6595,N_6970);
and U7491 (N_7491,N_6803,N_6948);
nor U7492 (N_7492,N_6940,N_6905);
nor U7493 (N_7493,N_6591,N_6798);
nand U7494 (N_7494,N_6706,N_6773);
and U7495 (N_7495,N_6666,N_6843);
or U7496 (N_7496,N_6847,N_6950);
xnor U7497 (N_7497,N_6650,N_6706);
and U7498 (N_7498,N_6820,N_6981);
or U7499 (N_7499,N_6987,N_6681);
and U7500 (N_7500,N_7043,N_7085);
and U7501 (N_7501,N_7236,N_7037);
nand U7502 (N_7502,N_7081,N_7016);
xor U7503 (N_7503,N_7278,N_7414);
xnor U7504 (N_7504,N_7339,N_7411);
and U7505 (N_7505,N_7231,N_7045);
nor U7506 (N_7506,N_7393,N_7413);
and U7507 (N_7507,N_7398,N_7395);
or U7508 (N_7508,N_7267,N_7362);
nor U7509 (N_7509,N_7464,N_7367);
nor U7510 (N_7510,N_7214,N_7299);
and U7511 (N_7511,N_7477,N_7342);
xnor U7512 (N_7512,N_7080,N_7283);
or U7513 (N_7513,N_7489,N_7087);
nor U7514 (N_7514,N_7116,N_7486);
and U7515 (N_7515,N_7293,N_7124);
nor U7516 (N_7516,N_7239,N_7454);
and U7517 (N_7517,N_7114,N_7424);
or U7518 (N_7518,N_7130,N_7333);
nand U7519 (N_7519,N_7257,N_7325);
xor U7520 (N_7520,N_7444,N_7034);
or U7521 (N_7521,N_7328,N_7296);
nand U7522 (N_7522,N_7136,N_7370);
nand U7523 (N_7523,N_7379,N_7055);
or U7524 (N_7524,N_7023,N_7190);
xnor U7525 (N_7525,N_7436,N_7264);
or U7526 (N_7526,N_7331,N_7015);
nand U7527 (N_7527,N_7295,N_7374);
nor U7528 (N_7528,N_7117,N_7448);
and U7529 (N_7529,N_7074,N_7188);
or U7530 (N_7530,N_7173,N_7334);
nor U7531 (N_7531,N_7323,N_7242);
and U7532 (N_7532,N_7307,N_7397);
or U7533 (N_7533,N_7460,N_7490);
and U7534 (N_7534,N_7306,N_7327);
or U7535 (N_7535,N_7010,N_7450);
nand U7536 (N_7536,N_7275,N_7462);
xor U7537 (N_7537,N_7389,N_7358);
and U7538 (N_7538,N_7258,N_7388);
nand U7539 (N_7539,N_7059,N_7083);
xnor U7540 (N_7540,N_7135,N_7259);
xnor U7541 (N_7541,N_7063,N_7143);
nor U7542 (N_7542,N_7218,N_7468);
and U7543 (N_7543,N_7058,N_7423);
and U7544 (N_7544,N_7113,N_7256);
or U7545 (N_7545,N_7095,N_7394);
nand U7546 (N_7546,N_7147,N_7409);
xor U7547 (N_7547,N_7240,N_7150);
and U7548 (N_7548,N_7309,N_7392);
and U7549 (N_7549,N_7094,N_7496);
nor U7550 (N_7550,N_7338,N_7335);
or U7551 (N_7551,N_7207,N_7181);
or U7552 (N_7552,N_7452,N_7006);
nand U7553 (N_7553,N_7065,N_7024);
and U7554 (N_7554,N_7433,N_7429);
nor U7555 (N_7555,N_7203,N_7385);
nor U7556 (N_7556,N_7050,N_7132);
nand U7557 (N_7557,N_7090,N_7194);
or U7558 (N_7558,N_7282,N_7220);
nor U7559 (N_7559,N_7463,N_7202);
or U7560 (N_7560,N_7269,N_7241);
and U7561 (N_7561,N_7435,N_7300);
or U7562 (N_7562,N_7175,N_7308);
nor U7563 (N_7563,N_7329,N_7156);
nor U7564 (N_7564,N_7073,N_7162);
nor U7565 (N_7565,N_7018,N_7227);
nand U7566 (N_7566,N_7245,N_7062);
and U7567 (N_7567,N_7349,N_7281);
and U7568 (N_7568,N_7209,N_7115);
or U7569 (N_7569,N_7294,N_7426);
nand U7570 (N_7570,N_7012,N_7330);
and U7571 (N_7571,N_7149,N_7487);
and U7572 (N_7572,N_7292,N_7076);
or U7573 (N_7573,N_7110,N_7304);
nand U7574 (N_7574,N_7211,N_7048);
or U7575 (N_7575,N_7177,N_7105);
and U7576 (N_7576,N_7079,N_7298);
xnor U7577 (N_7577,N_7100,N_7266);
nor U7578 (N_7578,N_7461,N_7287);
xor U7579 (N_7579,N_7051,N_7163);
xnor U7580 (N_7580,N_7263,N_7168);
and U7581 (N_7581,N_7431,N_7320);
and U7582 (N_7582,N_7021,N_7366);
and U7583 (N_7583,N_7088,N_7072);
nor U7584 (N_7584,N_7430,N_7495);
nand U7585 (N_7585,N_7302,N_7321);
xor U7586 (N_7586,N_7291,N_7446);
nand U7587 (N_7587,N_7474,N_7102);
nor U7588 (N_7588,N_7099,N_7467);
xor U7589 (N_7589,N_7000,N_7224);
nand U7590 (N_7590,N_7142,N_7332);
nor U7591 (N_7591,N_7442,N_7170);
xor U7592 (N_7592,N_7390,N_7164);
and U7593 (N_7593,N_7376,N_7032);
nor U7594 (N_7594,N_7399,N_7350);
nor U7595 (N_7595,N_7415,N_7199);
nor U7596 (N_7596,N_7345,N_7122);
nor U7597 (N_7597,N_7315,N_7494);
and U7598 (N_7598,N_7420,N_7035);
nor U7599 (N_7599,N_7009,N_7054);
or U7600 (N_7600,N_7128,N_7185);
xor U7601 (N_7601,N_7033,N_7145);
or U7602 (N_7602,N_7456,N_7191);
xor U7603 (N_7603,N_7425,N_7377);
nand U7604 (N_7604,N_7449,N_7255);
xor U7605 (N_7605,N_7372,N_7225);
nand U7606 (N_7606,N_7089,N_7466);
or U7607 (N_7607,N_7071,N_7198);
xnor U7608 (N_7608,N_7246,N_7101);
or U7609 (N_7609,N_7154,N_7223);
and U7610 (N_7610,N_7221,N_7052);
nor U7611 (N_7611,N_7410,N_7028);
or U7612 (N_7612,N_7406,N_7151);
nor U7613 (N_7613,N_7493,N_7165);
and U7614 (N_7614,N_7363,N_7003);
xnor U7615 (N_7615,N_7251,N_7235);
or U7616 (N_7616,N_7407,N_7382);
and U7617 (N_7617,N_7457,N_7280);
and U7618 (N_7618,N_7137,N_7357);
or U7619 (N_7619,N_7230,N_7371);
nor U7620 (N_7620,N_7445,N_7391);
or U7621 (N_7621,N_7111,N_7289);
and U7622 (N_7622,N_7483,N_7437);
and U7623 (N_7623,N_7014,N_7030);
nand U7624 (N_7624,N_7476,N_7131);
nand U7625 (N_7625,N_7238,N_7479);
nor U7626 (N_7626,N_7498,N_7305);
and U7627 (N_7627,N_7405,N_7475);
and U7628 (N_7628,N_7134,N_7482);
or U7629 (N_7629,N_7008,N_7233);
or U7630 (N_7630,N_7152,N_7078);
xnor U7631 (N_7631,N_7272,N_7419);
xnor U7632 (N_7632,N_7216,N_7084);
or U7633 (N_7633,N_7192,N_7208);
and U7634 (N_7634,N_7253,N_7344);
nand U7635 (N_7635,N_7180,N_7140);
nor U7636 (N_7636,N_7061,N_7096);
or U7637 (N_7637,N_7481,N_7262);
and U7638 (N_7638,N_7318,N_7404);
or U7639 (N_7639,N_7109,N_7271);
and U7640 (N_7640,N_7066,N_7206);
nor U7641 (N_7641,N_7019,N_7228);
xnor U7642 (N_7642,N_7260,N_7127);
or U7643 (N_7643,N_7057,N_7148);
nor U7644 (N_7644,N_7249,N_7270);
xnor U7645 (N_7645,N_7416,N_7120);
nor U7646 (N_7646,N_7056,N_7312);
nand U7647 (N_7647,N_7020,N_7107);
nor U7648 (N_7648,N_7011,N_7176);
or U7649 (N_7649,N_7195,N_7441);
and U7650 (N_7650,N_7121,N_7252);
nand U7651 (N_7651,N_7352,N_7166);
and U7652 (N_7652,N_7284,N_7417);
or U7653 (N_7653,N_7119,N_7069);
and U7654 (N_7654,N_7356,N_7403);
nand U7655 (N_7655,N_7067,N_7364);
and U7656 (N_7656,N_7244,N_7314);
nor U7657 (N_7657,N_7365,N_7285);
xnor U7658 (N_7658,N_7402,N_7027);
nand U7659 (N_7659,N_7039,N_7373);
or U7660 (N_7660,N_7106,N_7215);
xnor U7661 (N_7661,N_7005,N_7155);
nand U7662 (N_7662,N_7104,N_7288);
xor U7663 (N_7663,N_7485,N_7488);
or U7664 (N_7664,N_7210,N_7053);
nor U7665 (N_7665,N_7369,N_7108);
and U7666 (N_7666,N_7025,N_7179);
or U7667 (N_7667,N_7473,N_7455);
and U7668 (N_7668,N_7311,N_7301);
or U7669 (N_7669,N_7212,N_7491);
nor U7670 (N_7670,N_7360,N_7205);
xor U7671 (N_7671,N_7217,N_7348);
xnor U7672 (N_7672,N_7182,N_7459);
nor U7673 (N_7673,N_7219,N_7492);
or U7674 (N_7674,N_7343,N_7093);
or U7675 (N_7675,N_7297,N_7091);
and U7676 (N_7676,N_7167,N_7480);
nand U7677 (N_7677,N_7317,N_7268);
or U7678 (N_7678,N_7157,N_7123);
or U7679 (N_7679,N_7396,N_7361);
or U7680 (N_7680,N_7153,N_7324);
or U7681 (N_7681,N_7077,N_7243);
and U7682 (N_7682,N_7286,N_7026);
or U7683 (N_7683,N_7440,N_7041);
and U7684 (N_7684,N_7354,N_7322);
or U7685 (N_7685,N_7200,N_7353);
and U7686 (N_7686,N_7472,N_7387);
nor U7687 (N_7687,N_7141,N_7499);
xnor U7688 (N_7688,N_7346,N_7378);
xor U7689 (N_7689,N_7375,N_7160);
nand U7690 (N_7690,N_7447,N_7384);
xnor U7691 (N_7691,N_7196,N_7277);
nand U7692 (N_7692,N_7158,N_7336);
and U7693 (N_7693,N_7412,N_7193);
or U7694 (N_7694,N_7174,N_7001);
and U7695 (N_7695,N_7098,N_7383);
or U7696 (N_7696,N_7274,N_7443);
or U7697 (N_7697,N_7234,N_7161);
nand U7698 (N_7698,N_7310,N_7082);
nand U7699 (N_7699,N_7178,N_7290);
nor U7700 (N_7700,N_7359,N_7368);
nor U7701 (N_7701,N_7451,N_7261);
and U7702 (N_7702,N_7478,N_7184);
nand U7703 (N_7703,N_7421,N_7250);
and U7704 (N_7704,N_7031,N_7002);
nor U7705 (N_7705,N_7386,N_7171);
or U7706 (N_7706,N_7438,N_7213);
nand U7707 (N_7707,N_7279,N_7380);
nand U7708 (N_7708,N_7340,N_7118);
xnor U7709 (N_7709,N_7484,N_7139);
nand U7710 (N_7710,N_7319,N_7273);
or U7711 (N_7711,N_7418,N_7347);
nand U7712 (N_7712,N_7470,N_7204);
nor U7713 (N_7713,N_7038,N_7036);
nor U7714 (N_7714,N_7432,N_7408);
xor U7715 (N_7715,N_7400,N_7017);
xor U7716 (N_7716,N_7047,N_7497);
nor U7717 (N_7717,N_7042,N_7044);
xnor U7718 (N_7718,N_7427,N_7060);
nor U7719 (N_7719,N_7049,N_7326);
or U7720 (N_7720,N_7125,N_7068);
or U7721 (N_7721,N_7265,N_7381);
nand U7722 (N_7722,N_7428,N_7422);
nor U7723 (N_7723,N_7013,N_7126);
or U7724 (N_7724,N_7189,N_7197);
or U7725 (N_7725,N_7401,N_7133);
or U7726 (N_7726,N_7112,N_7351);
or U7727 (N_7727,N_7471,N_7159);
nand U7728 (N_7728,N_7458,N_7186);
or U7729 (N_7729,N_7146,N_7169);
or U7730 (N_7730,N_7434,N_7465);
xor U7731 (N_7731,N_7313,N_7247);
nand U7732 (N_7732,N_7183,N_7237);
and U7733 (N_7733,N_7004,N_7144);
xor U7734 (N_7734,N_7064,N_7232);
and U7735 (N_7735,N_7248,N_7040);
xnor U7736 (N_7736,N_7276,N_7254);
xnor U7737 (N_7737,N_7453,N_7229);
nor U7738 (N_7738,N_7103,N_7138);
nor U7739 (N_7739,N_7355,N_7129);
nor U7740 (N_7740,N_7172,N_7086);
nor U7741 (N_7741,N_7029,N_7022);
and U7742 (N_7742,N_7201,N_7226);
and U7743 (N_7743,N_7222,N_7092);
xor U7744 (N_7744,N_7046,N_7341);
xnor U7745 (N_7745,N_7070,N_7187);
or U7746 (N_7746,N_7337,N_7439);
and U7747 (N_7747,N_7097,N_7007);
xnor U7748 (N_7748,N_7075,N_7303);
xor U7749 (N_7749,N_7316,N_7469);
nor U7750 (N_7750,N_7144,N_7146);
nand U7751 (N_7751,N_7015,N_7387);
or U7752 (N_7752,N_7064,N_7424);
xor U7753 (N_7753,N_7327,N_7055);
xor U7754 (N_7754,N_7448,N_7197);
nor U7755 (N_7755,N_7436,N_7358);
and U7756 (N_7756,N_7349,N_7457);
and U7757 (N_7757,N_7260,N_7183);
nand U7758 (N_7758,N_7459,N_7005);
or U7759 (N_7759,N_7214,N_7439);
or U7760 (N_7760,N_7482,N_7194);
nor U7761 (N_7761,N_7275,N_7078);
nand U7762 (N_7762,N_7161,N_7318);
nor U7763 (N_7763,N_7318,N_7385);
or U7764 (N_7764,N_7038,N_7029);
nor U7765 (N_7765,N_7100,N_7352);
and U7766 (N_7766,N_7321,N_7240);
nor U7767 (N_7767,N_7089,N_7259);
nand U7768 (N_7768,N_7345,N_7063);
nor U7769 (N_7769,N_7228,N_7232);
xnor U7770 (N_7770,N_7317,N_7004);
xnor U7771 (N_7771,N_7231,N_7171);
xor U7772 (N_7772,N_7265,N_7118);
nand U7773 (N_7773,N_7387,N_7066);
nor U7774 (N_7774,N_7298,N_7044);
nand U7775 (N_7775,N_7352,N_7015);
and U7776 (N_7776,N_7240,N_7260);
or U7777 (N_7777,N_7308,N_7273);
and U7778 (N_7778,N_7153,N_7140);
nand U7779 (N_7779,N_7139,N_7440);
nand U7780 (N_7780,N_7027,N_7096);
and U7781 (N_7781,N_7458,N_7112);
or U7782 (N_7782,N_7182,N_7427);
or U7783 (N_7783,N_7342,N_7381);
nor U7784 (N_7784,N_7261,N_7183);
xnor U7785 (N_7785,N_7183,N_7469);
xor U7786 (N_7786,N_7020,N_7222);
and U7787 (N_7787,N_7266,N_7149);
and U7788 (N_7788,N_7414,N_7434);
and U7789 (N_7789,N_7210,N_7206);
nor U7790 (N_7790,N_7476,N_7419);
or U7791 (N_7791,N_7139,N_7236);
xor U7792 (N_7792,N_7133,N_7419);
xnor U7793 (N_7793,N_7044,N_7419);
or U7794 (N_7794,N_7460,N_7149);
and U7795 (N_7795,N_7193,N_7028);
nand U7796 (N_7796,N_7148,N_7083);
nor U7797 (N_7797,N_7273,N_7136);
nor U7798 (N_7798,N_7003,N_7161);
nor U7799 (N_7799,N_7255,N_7095);
nor U7800 (N_7800,N_7278,N_7271);
and U7801 (N_7801,N_7005,N_7216);
nor U7802 (N_7802,N_7032,N_7242);
and U7803 (N_7803,N_7015,N_7283);
xnor U7804 (N_7804,N_7167,N_7450);
nor U7805 (N_7805,N_7419,N_7409);
nor U7806 (N_7806,N_7433,N_7304);
nor U7807 (N_7807,N_7139,N_7060);
nor U7808 (N_7808,N_7303,N_7465);
or U7809 (N_7809,N_7009,N_7364);
and U7810 (N_7810,N_7443,N_7137);
xor U7811 (N_7811,N_7076,N_7004);
nand U7812 (N_7812,N_7420,N_7307);
and U7813 (N_7813,N_7424,N_7152);
nor U7814 (N_7814,N_7006,N_7062);
xor U7815 (N_7815,N_7214,N_7126);
and U7816 (N_7816,N_7446,N_7148);
nor U7817 (N_7817,N_7111,N_7358);
nor U7818 (N_7818,N_7225,N_7492);
xnor U7819 (N_7819,N_7183,N_7057);
and U7820 (N_7820,N_7134,N_7005);
nand U7821 (N_7821,N_7264,N_7437);
or U7822 (N_7822,N_7278,N_7242);
nand U7823 (N_7823,N_7466,N_7219);
and U7824 (N_7824,N_7122,N_7172);
nor U7825 (N_7825,N_7191,N_7098);
nor U7826 (N_7826,N_7123,N_7320);
nor U7827 (N_7827,N_7231,N_7464);
or U7828 (N_7828,N_7281,N_7144);
or U7829 (N_7829,N_7090,N_7433);
or U7830 (N_7830,N_7161,N_7420);
xor U7831 (N_7831,N_7443,N_7159);
nor U7832 (N_7832,N_7052,N_7407);
nand U7833 (N_7833,N_7054,N_7216);
and U7834 (N_7834,N_7121,N_7221);
xor U7835 (N_7835,N_7078,N_7493);
nand U7836 (N_7836,N_7073,N_7093);
and U7837 (N_7837,N_7328,N_7126);
xnor U7838 (N_7838,N_7081,N_7423);
nand U7839 (N_7839,N_7442,N_7466);
or U7840 (N_7840,N_7289,N_7467);
nand U7841 (N_7841,N_7145,N_7419);
or U7842 (N_7842,N_7274,N_7277);
or U7843 (N_7843,N_7318,N_7377);
and U7844 (N_7844,N_7189,N_7232);
or U7845 (N_7845,N_7190,N_7201);
and U7846 (N_7846,N_7490,N_7218);
nor U7847 (N_7847,N_7041,N_7012);
and U7848 (N_7848,N_7291,N_7090);
xnor U7849 (N_7849,N_7103,N_7404);
and U7850 (N_7850,N_7291,N_7404);
and U7851 (N_7851,N_7252,N_7294);
and U7852 (N_7852,N_7067,N_7182);
nor U7853 (N_7853,N_7151,N_7127);
nand U7854 (N_7854,N_7324,N_7231);
nand U7855 (N_7855,N_7348,N_7225);
and U7856 (N_7856,N_7428,N_7008);
nor U7857 (N_7857,N_7049,N_7367);
and U7858 (N_7858,N_7291,N_7443);
or U7859 (N_7859,N_7167,N_7093);
and U7860 (N_7860,N_7267,N_7458);
nand U7861 (N_7861,N_7287,N_7412);
or U7862 (N_7862,N_7449,N_7455);
xor U7863 (N_7863,N_7088,N_7213);
or U7864 (N_7864,N_7044,N_7201);
nor U7865 (N_7865,N_7165,N_7499);
nor U7866 (N_7866,N_7315,N_7354);
xor U7867 (N_7867,N_7110,N_7368);
nor U7868 (N_7868,N_7213,N_7339);
or U7869 (N_7869,N_7257,N_7002);
or U7870 (N_7870,N_7029,N_7229);
and U7871 (N_7871,N_7468,N_7331);
and U7872 (N_7872,N_7071,N_7049);
nand U7873 (N_7873,N_7036,N_7065);
xnor U7874 (N_7874,N_7326,N_7039);
nor U7875 (N_7875,N_7081,N_7355);
nor U7876 (N_7876,N_7350,N_7022);
or U7877 (N_7877,N_7125,N_7237);
or U7878 (N_7878,N_7162,N_7161);
nor U7879 (N_7879,N_7156,N_7039);
nand U7880 (N_7880,N_7242,N_7193);
or U7881 (N_7881,N_7410,N_7302);
xor U7882 (N_7882,N_7412,N_7327);
or U7883 (N_7883,N_7048,N_7107);
nand U7884 (N_7884,N_7427,N_7281);
nor U7885 (N_7885,N_7171,N_7346);
and U7886 (N_7886,N_7053,N_7147);
and U7887 (N_7887,N_7296,N_7242);
xor U7888 (N_7888,N_7168,N_7259);
xnor U7889 (N_7889,N_7364,N_7083);
nor U7890 (N_7890,N_7163,N_7085);
nor U7891 (N_7891,N_7302,N_7003);
nand U7892 (N_7892,N_7169,N_7057);
and U7893 (N_7893,N_7465,N_7015);
and U7894 (N_7894,N_7403,N_7305);
nor U7895 (N_7895,N_7006,N_7282);
nor U7896 (N_7896,N_7047,N_7333);
xor U7897 (N_7897,N_7295,N_7225);
and U7898 (N_7898,N_7320,N_7124);
or U7899 (N_7899,N_7432,N_7165);
xor U7900 (N_7900,N_7313,N_7284);
nand U7901 (N_7901,N_7279,N_7163);
nor U7902 (N_7902,N_7035,N_7312);
nand U7903 (N_7903,N_7149,N_7089);
or U7904 (N_7904,N_7089,N_7465);
xor U7905 (N_7905,N_7152,N_7361);
or U7906 (N_7906,N_7435,N_7431);
or U7907 (N_7907,N_7419,N_7295);
nor U7908 (N_7908,N_7133,N_7335);
or U7909 (N_7909,N_7240,N_7136);
and U7910 (N_7910,N_7374,N_7410);
and U7911 (N_7911,N_7045,N_7188);
nand U7912 (N_7912,N_7466,N_7498);
or U7913 (N_7913,N_7486,N_7131);
or U7914 (N_7914,N_7414,N_7181);
nand U7915 (N_7915,N_7457,N_7444);
or U7916 (N_7916,N_7200,N_7126);
nand U7917 (N_7917,N_7224,N_7240);
xnor U7918 (N_7918,N_7390,N_7187);
xnor U7919 (N_7919,N_7268,N_7314);
xnor U7920 (N_7920,N_7442,N_7116);
nand U7921 (N_7921,N_7004,N_7219);
nand U7922 (N_7922,N_7338,N_7183);
xnor U7923 (N_7923,N_7289,N_7424);
and U7924 (N_7924,N_7284,N_7001);
or U7925 (N_7925,N_7051,N_7371);
xnor U7926 (N_7926,N_7096,N_7236);
nor U7927 (N_7927,N_7303,N_7219);
and U7928 (N_7928,N_7048,N_7121);
and U7929 (N_7929,N_7431,N_7050);
and U7930 (N_7930,N_7231,N_7077);
xnor U7931 (N_7931,N_7018,N_7393);
xor U7932 (N_7932,N_7487,N_7103);
xor U7933 (N_7933,N_7415,N_7427);
or U7934 (N_7934,N_7487,N_7244);
xnor U7935 (N_7935,N_7477,N_7173);
and U7936 (N_7936,N_7213,N_7222);
or U7937 (N_7937,N_7403,N_7139);
nor U7938 (N_7938,N_7157,N_7446);
nand U7939 (N_7939,N_7408,N_7219);
nor U7940 (N_7940,N_7242,N_7158);
nand U7941 (N_7941,N_7386,N_7367);
nor U7942 (N_7942,N_7307,N_7283);
nor U7943 (N_7943,N_7150,N_7280);
nand U7944 (N_7944,N_7380,N_7361);
nand U7945 (N_7945,N_7149,N_7290);
nor U7946 (N_7946,N_7272,N_7184);
nor U7947 (N_7947,N_7124,N_7083);
nand U7948 (N_7948,N_7045,N_7428);
and U7949 (N_7949,N_7336,N_7311);
and U7950 (N_7950,N_7216,N_7205);
nor U7951 (N_7951,N_7138,N_7209);
and U7952 (N_7952,N_7201,N_7451);
nor U7953 (N_7953,N_7219,N_7092);
or U7954 (N_7954,N_7052,N_7147);
and U7955 (N_7955,N_7455,N_7250);
or U7956 (N_7956,N_7136,N_7481);
nand U7957 (N_7957,N_7296,N_7194);
nor U7958 (N_7958,N_7300,N_7332);
or U7959 (N_7959,N_7187,N_7416);
nand U7960 (N_7960,N_7206,N_7301);
nand U7961 (N_7961,N_7466,N_7333);
and U7962 (N_7962,N_7350,N_7301);
and U7963 (N_7963,N_7355,N_7190);
and U7964 (N_7964,N_7364,N_7443);
nand U7965 (N_7965,N_7410,N_7226);
and U7966 (N_7966,N_7390,N_7042);
nand U7967 (N_7967,N_7268,N_7194);
and U7968 (N_7968,N_7478,N_7017);
nand U7969 (N_7969,N_7243,N_7010);
xnor U7970 (N_7970,N_7354,N_7083);
and U7971 (N_7971,N_7482,N_7427);
xnor U7972 (N_7972,N_7223,N_7395);
xor U7973 (N_7973,N_7497,N_7338);
and U7974 (N_7974,N_7484,N_7470);
nor U7975 (N_7975,N_7488,N_7204);
or U7976 (N_7976,N_7425,N_7355);
and U7977 (N_7977,N_7375,N_7096);
or U7978 (N_7978,N_7300,N_7074);
xnor U7979 (N_7979,N_7496,N_7075);
nand U7980 (N_7980,N_7465,N_7429);
and U7981 (N_7981,N_7261,N_7056);
and U7982 (N_7982,N_7175,N_7050);
nor U7983 (N_7983,N_7144,N_7332);
xor U7984 (N_7984,N_7227,N_7207);
and U7985 (N_7985,N_7047,N_7002);
or U7986 (N_7986,N_7016,N_7222);
or U7987 (N_7987,N_7498,N_7270);
and U7988 (N_7988,N_7487,N_7186);
nor U7989 (N_7989,N_7276,N_7423);
nor U7990 (N_7990,N_7324,N_7086);
xnor U7991 (N_7991,N_7111,N_7412);
or U7992 (N_7992,N_7442,N_7316);
and U7993 (N_7993,N_7186,N_7462);
xnor U7994 (N_7994,N_7380,N_7302);
nand U7995 (N_7995,N_7379,N_7411);
xor U7996 (N_7996,N_7113,N_7146);
nor U7997 (N_7997,N_7105,N_7206);
nor U7998 (N_7998,N_7160,N_7411);
xnor U7999 (N_7999,N_7395,N_7421);
nand U8000 (N_8000,N_7666,N_7589);
or U8001 (N_8001,N_7555,N_7635);
or U8002 (N_8002,N_7580,N_7551);
and U8003 (N_8003,N_7526,N_7821);
nand U8004 (N_8004,N_7889,N_7958);
xor U8005 (N_8005,N_7938,N_7664);
xor U8006 (N_8006,N_7903,N_7592);
nor U8007 (N_8007,N_7944,N_7516);
and U8008 (N_8008,N_7887,N_7886);
nor U8009 (N_8009,N_7630,N_7934);
or U8010 (N_8010,N_7579,N_7713);
nand U8011 (N_8011,N_7734,N_7679);
and U8012 (N_8012,N_7930,N_7646);
nand U8013 (N_8013,N_7918,N_7988);
xnor U8014 (N_8014,N_7833,N_7613);
nor U8015 (N_8015,N_7770,N_7917);
nand U8016 (N_8016,N_7844,N_7543);
and U8017 (N_8017,N_7858,N_7537);
or U8018 (N_8018,N_7552,N_7692);
and U8019 (N_8019,N_7603,N_7900);
or U8020 (N_8020,N_7622,N_7849);
nand U8021 (N_8021,N_7504,N_7688);
xor U8022 (N_8022,N_7800,N_7760);
nand U8023 (N_8023,N_7861,N_7680);
nor U8024 (N_8024,N_7864,N_7890);
nand U8025 (N_8025,N_7865,N_7932);
nand U8026 (N_8026,N_7607,N_7984);
nand U8027 (N_8027,N_7573,N_7556);
and U8028 (N_8028,N_7792,N_7565);
or U8029 (N_8029,N_7617,N_7740);
nor U8030 (N_8030,N_7819,N_7969);
xnor U8031 (N_8031,N_7924,N_7732);
nor U8032 (N_8032,N_7651,N_7633);
and U8033 (N_8033,N_7527,N_7851);
or U8034 (N_8034,N_7914,N_7721);
or U8035 (N_8035,N_7758,N_7827);
nor U8036 (N_8036,N_7710,N_7654);
and U8037 (N_8037,N_7789,N_7605);
or U8038 (N_8038,N_7545,N_7701);
and U8039 (N_8039,N_7649,N_7708);
nor U8040 (N_8040,N_7853,N_7945);
xnor U8041 (N_8041,N_7542,N_7793);
and U8042 (N_8042,N_7553,N_7567);
and U8043 (N_8043,N_7765,N_7790);
and U8044 (N_8044,N_7648,N_7628);
nor U8045 (N_8045,N_7523,N_7756);
nor U8046 (N_8046,N_7686,N_7593);
nand U8047 (N_8047,N_7882,N_7875);
or U8048 (N_8048,N_7586,N_7959);
nand U8049 (N_8049,N_7824,N_7677);
xor U8050 (N_8050,N_7750,N_7813);
nand U8051 (N_8051,N_7702,N_7775);
or U8052 (N_8052,N_7684,N_7743);
and U8053 (N_8053,N_7695,N_7896);
or U8054 (N_8054,N_7836,N_7643);
nor U8055 (N_8055,N_7698,N_7870);
nor U8056 (N_8056,N_7948,N_7538);
nand U8057 (N_8057,N_7672,N_7647);
nor U8058 (N_8058,N_7957,N_7976);
nor U8059 (N_8059,N_7719,N_7835);
xor U8060 (N_8060,N_7610,N_7518);
nand U8061 (N_8061,N_7894,N_7727);
nand U8062 (N_8062,N_7621,N_7971);
nor U8063 (N_8063,N_7967,N_7891);
nor U8064 (N_8064,N_7557,N_7787);
or U8065 (N_8065,N_7631,N_7590);
and U8066 (N_8066,N_7954,N_7587);
or U8067 (N_8067,N_7657,N_7892);
nand U8068 (N_8068,N_7873,N_7700);
or U8069 (N_8069,N_7685,N_7525);
and U8070 (N_8070,N_7987,N_7970);
nand U8071 (N_8071,N_7846,N_7842);
xor U8072 (N_8072,N_7747,N_7604);
xnor U8073 (N_8073,N_7759,N_7913);
xnor U8074 (N_8074,N_7895,N_7857);
nand U8075 (N_8075,N_7639,N_7779);
and U8076 (N_8076,N_7642,N_7659);
xor U8077 (N_8077,N_7634,N_7752);
xnor U8078 (N_8078,N_7572,N_7781);
xnor U8079 (N_8079,N_7978,N_7583);
nor U8080 (N_8080,N_7733,N_7626);
xnor U8081 (N_8081,N_7806,N_7506);
and U8082 (N_8082,N_7753,N_7581);
xnor U8083 (N_8083,N_7505,N_7645);
and U8084 (N_8084,N_7986,N_7673);
and U8085 (N_8085,N_7530,N_7600);
nor U8086 (N_8086,N_7879,N_7609);
nor U8087 (N_8087,N_7612,N_7766);
and U8088 (N_8088,N_7711,N_7939);
and U8089 (N_8089,N_7785,N_7755);
nand U8090 (N_8090,N_7624,N_7832);
or U8091 (N_8091,N_7736,N_7783);
or U8092 (N_8092,N_7859,N_7797);
nor U8093 (N_8093,N_7535,N_7510);
or U8094 (N_8094,N_7818,N_7746);
nor U8095 (N_8095,N_7638,N_7714);
and U8096 (N_8096,N_7597,N_7578);
xor U8097 (N_8097,N_7730,N_7905);
xor U8098 (N_8098,N_7860,N_7962);
xor U8099 (N_8099,N_7830,N_7801);
xnor U8100 (N_8100,N_7863,N_7855);
xor U8101 (N_8101,N_7568,N_7623);
or U8102 (N_8102,N_7802,N_7554);
nor U8103 (N_8103,N_7804,N_7699);
or U8104 (N_8104,N_7653,N_7739);
xor U8105 (N_8105,N_7868,N_7769);
or U8106 (N_8106,N_7803,N_7807);
nand U8107 (N_8107,N_7942,N_7697);
xnor U8108 (N_8108,N_7614,N_7540);
or U8109 (N_8109,N_7663,N_7536);
nand U8110 (N_8110,N_7876,N_7534);
or U8111 (N_8111,N_7595,N_7520);
xor U8112 (N_8112,N_7532,N_7784);
nor U8113 (N_8113,N_7549,N_7704);
xor U8114 (N_8114,N_7512,N_7943);
nor U8115 (N_8115,N_7715,N_7897);
and U8116 (N_8116,N_7656,N_7675);
or U8117 (N_8117,N_7550,N_7539);
nor U8118 (N_8118,N_7795,N_7931);
or U8119 (N_8119,N_7618,N_7788);
nor U8120 (N_8120,N_7662,N_7823);
nand U8121 (N_8121,N_7757,N_7817);
nand U8122 (N_8122,N_7687,N_7723);
nand U8123 (N_8123,N_7754,N_7718);
nor U8124 (N_8124,N_7762,N_7862);
and U8125 (N_8125,N_7564,N_7991);
and U8126 (N_8126,N_7728,N_7773);
xnor U8127 (N_8127,N_7794,N_7652);
or U8128 (N_8128,N_7840,N_7919);
nor U8129 (N_8129,N_7611,N_7776);
nand U8130 (N_8130,N_7852,N_7927);
xnor U8131 (N_8131,N_7737,N_7764);
xor U8132 (N_8132,N_7601,N_7906);
and U8133 (N_8133,N_7502,N_7972);
xnor U8134 (N_8134,N_7899,N_7831);
nand U8135 (N_8135,N_7509,N_7582);
nor U8136 (N_8136,N_7636,N_7742);
nand U8137 (N_8137,N_7848,N_7528);
and U8138 (N_8138,N_7508,N_7867);
and U8139 (N_8139,N_7820,N_7637);
nand U8140 (N_8140,N_7885,N_7616);
nor U8141 (N_8141,N_7731,N_7955);
nor U8142 (N_8142,N_7751,N_7625);
and U8143 (N_8143,N_7901,N_7920);
nor U8144 (N_8144,N_7808,N_7606);
and U8145 (N_8145,N_7850,N_7812);
xnor U8146 (N_8146,N_7997,N_7544);
or U8147 (N_8147,N_7996,N_7741);
xor U8148 (N_8148,N_7980,N_7669);
and U8149 (N_8149,N_7993,N_7771);
nand U8150 (N_8150,N_7947,N_7574);
nand U8151 (N_8151,N_7712,N_7560);
nor U8152 (N_8152,N_7777,N_7569);
and U8153 (N_8153,N_7585,N_7854);
xnor U8154 (N_8154,N_7524,N_7627);
nor U8155 (N_8155,N_7973,N_7898);
xor U8156 (N_8156,N_7881,N_7620);
xor U8157 (N_8157,N_7866,N_7665);
nand U8158 (N_8158,N_7904,N_7547);
or U8159 (N_8159,N_7640,N_7632);
and U8160 (N_8160,N_7845,N_7834);
nor U8161 (N_8161,N_7811,N_7884);
or U8162 (N_8162,N_7791,N_7933);
xor U8163 (N_8163,N_7722,N_7594);
and U8164 (N_8164,N_7735,N_7989);
and U8165 (N_8165,N_7936,N_7909);
or U8166 (N_8166,N_7968,N_7922);
and U8167 (N_8167,N_7888,N_7575);
nor U8168 (N_8168,N_7816,N_7966);
xor U8169 (N_8169,N_7563,N_7694);
nand U8170 (N_8170,N_7650,N_7546);
nand U8171 (N_8171,N_7979,N_7916);
or U8172 (N_8172,N_7559,N_7990);
and U8173 (N_8173,N_7706,N_7562);
xor U8174 (N_8174,N_7577,N_7682);
or U8175 (N_8175,N_7693,N_7681);
nor U8176 (N_8176,N_7829,N_7500);
or U8177 (N_8177,N_7963,N_7629);
or U8178 (N_8178,N_7619,N_7641);
nor U8179 (N_8179,N_7515,N_7782);
xor U8180 (N_8180,N_7923,N_7951);
or U8181 (N_8181,N_7522,N_7725);
or U8182 (N_8182,N_7588,N_7602);
nand U8183 (N_8183,N_7940,N_7511);
and U8184 (N_8184,N_7707,N_7982);
nor U8185 (N_8185,N_7571,N_7696);
nand U8186 (N_8186,N_7961,N_7946);
xor U8187 (N_8187,N_7912,N_7837);
nand U8188 (N_8188,N_7763,N_7599);
nand U8189 (N_8189,N_7822,N_7745);
nor U8190 (N_8190,N_7883,N_7877);
nand U8191 (N_8191,N_7683,N_7902);
or U8192 (N_8192,N_7615,N_7507);
nor U8193 (N_8193,N_7558,N_7774);
xor U8194 (N_8194,N_7928,N_7810);
or U8195 (N_8195,N_7908,N_7720);
nand U8196 (N_8196,N_7570,N_7964);
xor U8197 (N_8197,N_7977,N_7729);
or U8198 (N_8198,N_7874,N_7514);
or U8199 (N_8199,N_7778,N_7748);
nand U8200 (N_8200,N_7780,N_7644);
nand U8201 (N_8201,N_7691,N_7838);
xnor U8202 (N_8202,N_7953,N_7591);
nor U8203 (N_8203,N_7965,N_7952);
nor U8204 (N_8204,N_7999,N_7660);
or U8205 (N_8205,N_7561,N_7880);
and U8206 (N_8206,N_7925,N_7926);
xnor U8207 (N_8207,N_7950,N_7761);
or U8208 (N_8208,N_7975,N_7661);
or U8209 (N_8209,N_7671,N_7533);
or U8210 (N_8210,N_7655,N_7893);
nand U8211 (N_8211,N_7847,N_7798);
and U8212 (N_8212,N_7872,N_7856);
nand U8213 (N_8213,N_7738,N_7839);
and U8214 (N_8214,N_7717,N_7541);
and U8215 (N_8215,N_7871,N_7981);
or U8216 (N_8216,N_7517,N_7674);
or U8217 (N_8217,N_7983,N_7676);
xnor U8218 (N_8218,N_7513,N_7548);
nand U8219 (N_8219,N_7941,N_7658);
nor U8220 (N_8220,N_7814,N_7935);
or U8221 (N_8221,N_7670,N_7786);
nor U8222 (N_8222,N_7869,N_7843);
nor U8223 (N_8223,N_7910,N_7678);
and U8224 (N_8224,N_7521,N_7907);
xnor U8225 (N_8225,N_7703,N_7668);
and U8226 (N_8226,N_7998,N_7503);
nor U8227 (N_8227,N_7841,N_7915);
xor U8228 (N_8228,N_7690,N_7825);
nand U8229 (N_8229,N_7911,N_7576);
or U8230 (N_8230,N_7768,N_7985);
and U8231 (N_8231,N_7584,N_7878);
nand U8232 (N_8232,N_7598,N_7501);
nand U8233 (N_8233,N_7809,N_7705);
xor U8234 (N_8234,N_7974,N_7744);
xnor U8235 (N_8235,N_7608,N_7772);
or U8236 (N_8236,N_7716,N_7767);
nand U8237 (N_8237,N_7596,N_7709);
xnor U8238 (N_8238,N_7667,N_7956);
or U8239 (N_8239,N_7724,N_7726);
nand U8240 (N_8240,N_7929,N_7529);
or U8241 (N_8241,N_7796,N_7828);
xor U8242 (N_8242,N_7992,N_7519);
nor U8243 (N_8243,N_7921,N_7815);
nor U8244 (N_8244,N_7949,N_7826);
xnor U8245 (N_8245,N_7566,N_7994);
or U8246 (N_8246,N_7799,N_7749);
and U8247 (N_8247,N_7960,N_7805);
nor U8248 (N_8248,N_7937,N_7531);
and U8249 (N_8249,N_7995,N_7689);
or U8250 (N_8250,N_7780,N_7808);
xor U8251 (N_8251,N_7703,N_7763);
nand U8252 (N_8252,N_7828,N_7676);
or U8253 (N_8253,N_7637,N_7555);
and U8254 (N_8254,N_7562,N_7669);
nor U8255 (N_8255,N_7642,N_7616);
nand U8256 (N_8256,N_7868,N_7537);
or U8257 (N_8257,N_7605,N_7710);
nor U8258 (N_8258,N_7785,N_7972);
xnor U8259 (N_8259,N_7903,N_7612);
nand U8260 (N_8260,N_7756,N_7721);
nand U8261 (N_8261,N_7785,N_7893);
nand U8262 (N_8262,N_7778,N_7630);
xnor U8263 (N_8263,N_7500,N_7632);
nand U8264 (N_8264,N_7615,N_7917);
nand U8265 (N_8265,N_7825,N_7797);
nand U8266 (N_8266,N_7930,N_7823);
or U8267 (N_8267,N_7795,N_7594);
or U8268 (N_8268,N_7573,N_7528);
or U8269 (N_8269,N_7913,N_7823);
and U8270 (N_8270,N_7724,N_7745);
nor U8271 (N_8271,N_7669,N_7769);
xnor U8272 (N_8272,N_7511,N_7705);
xor U8273 (N_8273,N_7636,N_7786);
and U8274 (N_8274,N_7677,N_7822);
and U8275 (N_8275,N_7513,N_7924);
nor U8276 (N_8276,N_7526,N_7733);
or U8277 (N_8277,N_7946,N_7854);
xnor U8278 (N_8278,N_7706,N_7817);
or U8279 (N_8279,N_7530,N_7639);
nor U8280 (N_8280,N_7911,N_7698);
nor U8281 (N_8281,N_7655,N_7771);
nor U8282 (N_8282,N_7811,N_7882);
or U8283 (N_8283,N_7843,N_7857);
nor U8284 (N_8284,N_7582,N_7955);
nor U8285 (N_8285,N_7960,N_7840);
nor U8286 (N_8286,N_7916,N_7941);
nor U8287 (N_8287,N_7832,N_7791);
nor U8288 (N_8288,N_7773,N_7648);
or U8289 (N_8289,N_7553,N_7814);
nor U8290 (N_8290,N_7785,N_7617);
nor U8291 (N_8291,N_7766,N_7961);
nor U8292 (N_8292,N_7595,N_7627);
nor U8293 (N_8293,N_7861,N_7988);
or U8294 (N_8294,N_7500,N_7555);
nor U8295 (N_8295,N_7956,N_7844);
or U8296 (N_8296,N_7644,N_7940);
xor U8297 (N_8297,N_7772,N_7814);
or U8298 (N_8298,N_7872,N_7706);
or U8299 (N_8299,N_7998,N_7619);
and U8300 (N_8300,N_7553,N_7929);
or U8301 (N_8301,N_7924,N_7955);
nand U8302 (N_8302,N_7993,N_7535);
xnor U8303 (N_8303,N_7535,N_7944);
or U8304 (N_8304,N_7719,N_7520);
nand U8305 (N_8305,N_7532,N_7757);
nand U8306 (N_8306,N_7844,N_7944);
xor U8307 (N_8307,N_7845,N_7542);
or U8308 (N_8308,N_7778,N_7851);
and U8309 (N_8309,N_7825,N_7576);
or U8310 (N_8310,N_7891,N_7838);
and U8311 (N_8311,N_7953,N_7512);
nor U8312 (N_8312,N_7628,N_7629);
nand U8313 (N_8313,N_7879,N_7952);
xor U8314 (N_8314,N_7704,N_7571);
or U8315 (N_8315,N_7868,N_7827);
nor U8316 (N_8316,N_7994,N_7607);
nor U8317 (N_8317,N_7536,N_7593);
nand U8318 (N_8318,N_7911,N_7506);
and U8319 (N_8319,N_7545,N_7900);
xnor U8320 (N_8320,N_7563,N_7550);
nand U8321 (N_8321,N_7690,N_7772);
nor U8322 (N_8322,N_7953,N_7560);
or U8323 (N_8323,N_7715,N_7769);
and U8324 (N_8324,N_7870,N_7725);
and U8325 (N_8325,N_7758,N_7800);
nand U8326 (N_8326,N_7734,N_7979);
nor U8327 (N_8327,N_7522,N_7877);
xnor U8328 (N_8328,N_7747,N_7938);
nand U8329 (N_8329,N_7897,N_7717);
xnor U8330 (N_8330,N_7757,N_7916);
xnor U8331 (N_8331,N_7591,N_7608);
and U8332 (N_8332,N_7547,N_7872);
or U8333 (N_8333,N_7581,N_7674);
and U8334 (N_8334,N_7719,N_7954);
nand U8335 (N_8335,N_7997,N_7808);
xor U8336 (N_8336,N_7941,N_7938);
xnor U8337 (N_8337,N_7661,N_7797);
and U8338 (N_8338,N_7813,N_7903);
or U8339 (N_8339,N_7871,N_7937);
nand U8340 (N_8340,N_7816,N_7879);
nand U8341 (N_8341,N_7746,N_7709);
nor U8342 (N_8342,N_7869,N_7891);
nor U8343 (N_8343,N_7555,N_7841);
and U8344 (N_8344,N_7782,N_7959);
or U8345 (N_8345,N_7968,N_7668);
nand U8346 (N_8346,N_7981,N_7796);
nor U8347 (N_8347,N_7504,N_7860);
nor U8348 (N_8348,N_7527,N_7836);
and U8349 (N_8349,N_7974,N_7536);
xnor U8350 (N_8350,N_7595,N_7710);
and U8351 (N_8351,N_7762,N_7865);
and U8352 (N_8352,N_7972,N_7597);
nor U8353 (N_8353,N_7548,N_7503);
nand U8354 (N_8354,N_7842,N_7966);
and U8355 (N_8355,N_7767,N_7904);
nor U8356 (N_8356,N_7903,N_7655);
nand U8357 (N_8357,N_7866,N_7702);
xnor U8358 (N_8358,N_7804,N_7818);
or U8359 (N_8359,N_7685,N_7607);
xnor U8360 (N_8360,N_7900,N_7547);
nor U8361 (N_8361,N_7636,N_7750);
or U8362 (N_8362,N_7682,N_7698);
xnor U8363 (N_8363,N_7887,N_7572);
xor U8364 (N_8364,N_7971,N_7700);
xnor U8365 (N_8365,N_7622,N_7880);
nor U8366 (N_8366,N_7910,N_7514);
nand U8367 (N_8367,N_7974,N_7755);
nand U8368 (N_8368,N_7782,N_7555);
nor U8369 (N_8369,N_7709,N_7790);
nand U8370 (N_8370,N_7726,N_7892);
or U8371 (N_8371,N_7683,N_7613);
nor U8372 (N_8372,N_7720,N_7851);
and U8373 (N_8373,N_7690,N_7591);
and U8374 (N_8374,N_7517,N_7890);
and U8375 (N_8375,N_7635,N_7986);
or U8376 (N_8376,N_7531,N_7580);
and U8377 (N_8377,N_7741,N_7674);
nand U8378 (N_8378,N_7739,N_7787);
or U8379 (N_8379,N_7503,N_7854);
or U8380 (N_8380,N_7935,N_7905);
or U8381 (N_8381,N_7886,N_7873);
nand U8382 (N_8382,N_7556,N_7654);
nor U8383 (N_8383,N_7875,N_7751);
and U8384 (N_8384,N_7532,N_7597);
xnor U8385 (N_8385,N_7528,N_7561);
or U8386 (N_8386,N_7935,N_7960);
and U8387 (N_8387,N_7637,N_7734);
and U8388 (N_8388,N_7707,N_7632);
or U8389 (N_8389,N_7710,N_7676);
nor U8390 (N_8390,N_7749,N_7821);
or U8391 (N_8391,N_7808,N_7822);
nand U8392 (N_8392,N_7797,N_7673);
nand U8393 (N_8393,N_7625,N_7777);
and U8394 (N_8394,N_7847,N_7756);
and U8395 (N_8395,N_7842,N_7533);
nor U8396 (N_8396,N_7781,N_7897);
and U8397 (N_8397,N_7807,N_7699);
or U8398 (N_8398,N_7825,N_7919);
xnor U8399 (N_8399,N_7809,N_7738);
xnor U8400 (N_8400,N_7727,N_7956);
or U8401 (N_8401,N_7948,N_7519);
nand U8402 (N_8402,N_7635,N_7579);
or U8403 (N_8403,N_7592,N_7999);
nor U8404 (N_8404,N_7917,N_7687);
and U8405 (N_8405,N_7547,N_7536);
nor U8406 (N_8406,N_7620,N_7543);
and U8407 (N_8407,N_7952,N_7815);
or U8408 (N_8408,N_7797,N_7516);
and U8409 (N_8409,N_7650,N_7958);
and U8410 (N_8410,N_7987,N_7763);
nor U8411 (N_8411,N_7921,N_7760);
and U8412 (N_8412,N_7962,N_7540);
nand U8413 (N_8413,N_7944,N_7756);
xor U8414 (N_8414,N_7623,N_7927);
xnor U8415 (N_8415,N_7988,N_7694);
xnor U8416 (N_8416,N_7655,N_7613);
xnor U8417 (N_8417,N_7772,N_7776);
nand U8418 (N_8418,N_7606,N_7877);
nor U8419 (N_8419,N_7949,N_7723);
and U8420 (N_8420,N_7888,N_7671);
xor U8421 (N_8421,N_7772,N_7774);
nor U8422 (N_8422,N_7638,N_7603);
and U8423 (N_8423,N_7874,N_7820);
nand U8424 (N_8424,N_7613,N_7941);
nor U8425 (N_8425,N_7888,N_7694);
and U8426 (N_8426,N_7607,N_7962);
nand U8427 (N_8427,N_7832,N_7595);
and U8428 (N_8428,N_7968,N_7817);
and U8429 (N_8429,N_7633,N_7659);
or U8430 (N_8430,N_7839,N_7865);
and U8431 (N_8431,N_7580,N_7590);
xor U8432 (N_8432,N_7761,N_7993);
nor U8433 (N_8433,N_7982,N_7840);
and U8434 (N_8434,N_7576,N_7804);
xor U8435 (N_8435,N_7670,N_7796);
nor U8436 (N_8436,N_7731,N_7515);
nor U8437 (N_8437,N_7623,N_7634);
nor U8438 (N_8438,N_7759,N_7664);
or U8439 (N_8439,N_7607,N_7843);
xnor U8440 (N_8440,N_7635,N_7895);
and U8441 (N_8441,N_7861,N_7974);
nor U8442 (N_8442,N_7644,N_7961);
and U8443 (N_8443,N_7957,N_7978);
xor U8444 (N_8444,N_7610,N_7691);
nand U8445 (N_8445,N_7820,N_7950);
or U8446 (N_8446,N_7893,N_7963);
and U8447 (N_8447,N_7840,N_7894);
or U8448 (N_8448,N_7520,N_7839);
and U8449 (N_8449,N_7804,N_7859);
xor U8450 (N_8450,N_7841,N_7633);
nor U8451 (N_8451,N_7556,N_7781);
xor U8452 (N_8452,N_7960,N_7986);
and U8453 (N_8453,N_7685,N_7552);
xor U8454 (N_8454,N_7672,N_7669);
or U8455 (N_8455,N_7940,N_7538);
and U8456 (N_8456,N_7573,N_7585);
and U8457 (N_8457,N_7872,N_7588);
xnor U8458 (N_8458,N_7938,N_7927);
and U8459 (N_8459,N_7924,N_7592);
nand U8460 (N_8460,N_7837,N_7981);
nand U8461 (N_8461,N_7906,N_7991);
xor U8462 (N_8462,N_7734,N_7840);
nand U8463 (N_8463,N_7816,N_7839);
nor U8464 (N_8464,N_7660,N_7545);
nand U8465 (N_8465,N_7921,N_7750);
nand U8466 (N_8466,N_7645,N_7916);
nor U8467 (N_8467,N_7577,N_7870);
and U8468 (N_8468,N_7741,N_7525);
xnor U8469 (N_8469,N_7639,N_7861);
xnor U8470 (N_8470,N_7625,N_7977);
and U8471 (N_8471,N_7816,N_7678);
xor U8472 (N_8472,N_7691,N_7665);
nor U8473 (N_8473,N_7579,N_7969);
and U8474 (N_8474,N_7847,N_7517);
nand U8475 (N_8475,N_7979,N_7678);
or U8476 (N_8476,N_7594,N_7713);
nand U8477 (N_8477,N_7542,N_7824);
nor U8478 (N_8478,N_7711,N_7573);
xor U8479 (N_8479,N_7873,N_7876);
nor U8480 (N_8480,N_7840,N_7836);
nor U8481 (N_8481,N_7574,N_7913);
xnor U8482 (N_8482,N_7926,N_7574);
or U8483 (N_8483,N_7730,N_7771);
nand U8484 (N_8484,N_7701,N_7828);
or U8485 (N_8485,N_7830,N_7885);
nor U8486 (N_8486,N_7871,N_7664);
or U8487 (N_8487,N_7570,N_7638);
nor U8488 (N_8488,N_7623,N_7775);
or U8489 (N_8489,N_7534,N_7674);
or U8490 (N_8490,N_7502,N_7943);
or U8491 (N_8491,N_7734,N_7685);
nor U8492 (N_8492,N_7814,N_7848);
nor U8493 (N_8493,N_7750,N_7936);
and U8494 (N_8494,N_7970,N_7800);
nand U8495 (N_8495,N_7885,N_7935);
or U8496 (N_8496,N_7992,N_7640);
nand U8497 (N_8497,N_7804,N_7539);
or U8498 (N_8498,N_7561,N_7598);
xnor U8499 (N_8499,N_7991,N_7751);
nand U8500 (N_8500,N_8482,N_8097);
and U8501 (N_8501,N_8091,N_8352);
and U8502 (N_8502,N_8227,N_8100);
xnor U8503 (N_8503,N_8449,N_8036);
xor U8504 (N_8504,N_8178,N_8072);
nand U8505 (N_8505,N_8346,N_8007);
nand U8506 (N_8506,N_8275,N_8447);
xor U8507 (N_8507,N_8414,N_8307);
and U8508 (N_8508,N_8089,N_8380);
or U8509 (N_8509,N_8134,N_8005);
nor U8510 (N_8510,N_8325,N_8437);
xnor U8511 (N_8511,N_8137,N_8408);
xor U8512 (N_8512,N_8110,N_8080);
xnor U8513 (N_8513,N_8396,N_8105);
nand U8514 (N_8514,N_8493,N_8245);
or U8515 (N_8515,N_8282,N_8364);
and U8516 (N_8516,N_8290,N_8451);
xnor U8517 (N_8517,N_8088,N_8019);
nand U8518 (N_8518,N_8454,N_8153);
and U8519 (N_8519,N_8341,N_8361);
xor U8520 (N_8520,N_8104,N_8018);
or U8521 (N_8521,N_8369,N_8326);
and U8522 (N_8522,N_8429,N_8147);
nor U8523 (N_8523,N_8377,N_8405);
or U8524 (N_8524,N_8498,N_8061);
or U8525 (N_8525,N_8191,N_8495);
or U8526 (N_8526,N_8442,N_8185);
xor U8527 (N_8527,N_8141,N_8001);
and U8528 (N_8528,N_8192,N_8206);
and U8529 (N_8529,N_8169,N_8268);
xnor U8530 (N_8530,N_8479,N_8472);
or U8531 (N_8531,N_8054,N_8453);
nor U8532 (N_8532,N_8024,N_8310);
nor U8533 (N_8533,N_8401,N_8195);
or U8534 (N_8534,N_8148,N_8271);
or U8535 (N_8535,N_8238,N_8004);
nand U8536 (N_8536,N_8120,N_8203);
or U8537 (N_8537,N_8150,N_8108);
nand U8538 (N_8538,N_8304,N_8035);
xor U8539 (N_8539,N_8095,N_8286);
nand U8540 (N_8540,N_8127,N_8022);
and U8541 (N_8541,N_8086,N_8115);
nand U8542 (N_8542,N_8237,N_8450);
or U8543 (N_8543,N_8174,N_8478);
xnor U8544 (N_8544,N_8042,N_8388);
and U8545 (N_8545,N_8164,N_8317);
nor U8546 (N_8546,N_8189,N_8138);
xnor U8547 (N_8547,N_8400,N_8183);
nand U8548 (N_8548,N_8101,N_8374);
xor U8549 (N_8549,N_8404,N_8426);
xnor U8550 (N_8550,N_8161,N_8443);
nand U8551 (N_8551,N_8053,N_8213);
xor U8552 (N_8552,N_8210,N_8470);
and U8553 (N_8553,N_8198,N_8133);
or U8554 (N_8554,N_8013,N_8335);
xnor U8555 (N_8555,N_8340,N_8242);
and U8556 (N_8556,N_8157,N_8209);
and U8557 (N_8557,N_8152,N_8350);
and U8558 (N_8558,N_8177,N_8219);
or U8559 (N_8559,N_8234,N_8247);
xnor U8560 (N_8560,N_8395,N_8240);
nand U8561 (N_8561,N_8006,N_8455);
and U8562 (N_8562,N_8309,N_8277);
nor U8563 (N_8563,N_8318,N_8154);
nor U8564 (N_8564,N_8311,N_8412);
or U8565 (N_8565,N_8246,N_8265);
nor U8566 (N_8566,N_8465,N_8038);
nand U8567 (N_8567,N_8354,N_8236);
or U8568 (N_8568,N_8250,N_8471);
xnor U8569 (N_8569,N_8003,N_8109);
xnor U8570 (N_8570,N_8376,N_8029);
or U8571 (N_8571,N_8272,N_8140);
nor U8572 (N_8572,N_8348,N_8468);
nand U8573 (N_8573,N_8264,N_8356);
xor U8574 (N_8574,N_8253,N_8079);
xnor U8575 (N_8575,N_8313,N_8216);
xnor U8576 (N_8576,N_8016,N_8288);
nor U8577 (N_8577,N_8474,N_8049);
nand U8578 (N_8578,N_8440,N_8333);
and U8579 (N_8579,N_8263,N_8258);
xnor U8580 (N_8580,N_8343,N_8139);
and U8581 (N_8581,N_8428,N_8349);
nand U8582 (N_8582,N_8324,N_8360);
xor U8583 (N_8583,N_8459,N_8394);
nand U8584 (N_8584,N_8251,N_8181);
and U8585 (N_8585,N_8381,N_8136);
and U8586 (N_8586,N_8112,N_8302);
xnor U8587 (N_8587,N_8332,N_8048);
and U8588 (N_8588,N_8480,N_8156);
xor U8589 (N_8589,N_8289,N_8434);
and U8590 (N_8590,N_8345,N_8039);
nand U8591 (N_8591,N_8030,N_8166);
or U8592 (N_8592,N_8175,N_8241);
and U8593 (N_8593,N_8432,N_8403);
nand U8594 (N_8594,N_8366,N_8045);
and U8595 (N_8595,N_8491,N_8121);
nor U8596 (N_8596,N_8303,N_8477);
nor U8597 (N_8597,N_8425,N_8033);
and U8598 (N_8598,N_8260,N_8344);
or U8599 (N_8599,N_8050,N_8383);
nand U8600 (N_8600,N_8301,N_8017);
nor U8601 (N_8601,N_8458,N_8365);
or U8602 (N_8602,N_8194,N_8489);
xnor U8603 (N_8603,N_8457,N_8043);
and U8604 (N_8604,N_8116,N_8363);
nand U8605 (N_8605,N_8207,N_8314);
nand U8606 (N_8606,N_8410,N_8222);
and U8607 (N_8607,N_8020,N_8230);
xnor U8608 (N_8608,N_8438,N_8028);
nor U8609 (N_8609,N_8186,N_8398);
xnor U8610 (N_8610,N_8235,N_8145);
nor U8611 (N_8611,N_8308,N_8293);
or U8612 (N_8612,N_8228,N_8098);
nor U8613 (N_8613,N_8391,N_8102);
nand U8614 (N_8614,N_8339,N_8372);
xnor U8615 (N_8615,N_8155,N_8467);
xor U8616 (N_8616,N_8399,N_8062);
or U8617 (N_8617,N_8362,N_8044);
and U8618 (N_8618,N_8023,N_8131);
xnor U8619 (N_8619,N_8221,N_8052);
nand U8620 (N_8620,N_8402,N_8461);
xor U8621 (N_8621,N_8421,N_8492);
or U8622 (N_8622,N_8010,N_8009);
and U8623 (N_8623,N_8046,N_8032);
nor U8624 (N_8624,N_8123,N_8473);
or U8625 (N_8625,N_8446,N_8456);
or U8626 (N_8626,N_8083,N_8323);
nor U8627 (N_8627,N_8070,N_8069);
or U8628 (N_8628,N_8182,N_8170);
nor U8629 (N_8629,N_8433,N_8488);
nor U8630 (N_8630,N_8390,N_8199);
xor U8631 (N_8631,N_8188,N_8357);
nor U8632 (N_8632,N_8312,N_8129);
xnor U8633 (N_8633,N_8321,N_8034);
or U8634 (N_8634,N_8196,N_8485);
nor U8635 (N_8635,N_8081,N_8090);
or U8636 (N_8636,N_8233,N_8217);
and U8637 (N_8637,N_8201,N_8111);
nand U8638 (N_8638,N_8370,N_8299);
nor U8639 (N_8639,N_8397,N_8142);
nand U8640 (N_8640,N_8291,N_8214);
nand U8641 (N_8641,N_8296,N_8287);
nand U8642 (N_8642,N_8257,N_8096);
xor U8643 (N_8643,N_8071,N_8292);
or U8644 (N_8644,N_8204,N_8160);
xnor U8645 (N_8645,N_8243,N_8068);
xor U8646 (N_8646,N_8334,N_8278);
nor U8647 (N_8647,N_8322,N_8436);
or U8648 (N_8648,N_8078,N_8176);
nor U8649 (N_8649,N_8063,N_8431);
nand U8650 (N_8650,N_8211,N_8040);
nor U8651 (N_8651,N_8371,N_8144);
or U8652 (N_8652,N_8392,N_8294);
nand U8653 (N_8653,N_8143,N_8122);
nor U8654 (N_8654,N_8416,N_8439);
and U8655 (N_8655,N_8419,N_8220);
nor U8656 (N_8656,N_8167,N_8355);
nor U8657 (N_8657,N_8226,N_8021);
nand U8658 (N_8658,N_8256,N_8190);
nor U8659 (N_8659,N_8358,N_8469);
nor U8660 (N_8660,N_8295,N_8171);
and U8661 (N_8661,N_8205,N_8483);
xnor U8662 (N_8662,N_8087,N_8389);
and U8663 (N_8663,N_8427,N_8276);
nor U8664 (N_8664,N_8151,N_8387);
nand U8665 (N_8665,N_8342,N_8094);
nor U8666 (N_8666,N_8417,N_8497);
nor U8667 (N_8667,N_8119,N_8012);
and U8668 (N_8668,N_8014,N_8306);
or U8669 (N_8669,N_8279,N_8285);
or U8670 (N_8670,N_8172,N_8281);
or U8671 (N_8671,N_8064,N_8117);
nor U8672 (N_8672,N_8329,N_8353);
xor U8673 (N_8673,N_8315,N_8411);
or U8674 (N_8674,N_8487,N_8375);
nand U8675 (N_8675,N_8011,N_8280);
nor U8676 (N_8676,N_8008,N_8331);
or U8677 (N_8677,N_8422,N_8202);
nand U8678 (N_8678,N_8464,N_8481);
xor U8679 (N_8679,N_8269,N_8475);
nand U8680 (N_8680,N_8093,N_8259);
or U8681 (N_8681,N_8225,N_8056);
xnor U8682 (N_8682,N_8074,N_8076);
nor U8683 (N_8683,N_8073,N_8415);
and U8684 (N_8684,N_8430,N_8359);
or U8685 (N_8685,N_8420,N_8179);
and U8686 (N_8686,N_8298,N_8300);
and U8687 (N_8687,N_8320,N_8476);
or U8688 (N_8688,N_8158,N_8239);
nand U8689 (N_8689,N_8124,N_8099);
nand U8690 (N_8690,N_8060,N_8319);
and U8691 (N_8691,N_8379,N_8067);
or U8692 (N_8692,N_8327,N_8406);
nand U8693 (N_8693,N_8031,N_8218);
nor U8694 (N_8694,N_8163,N_8173);
nand U8695 (N_8695,N_8103,N_8025);
and U8696 (N_8696,N_8180,N_8384);
or U8697 (N_8697,N_8229,N_8126);
nand U8698 (N_8698,N_8284,N_8146);
xnor U8699 (N_8699,N_8149,N_8418);
or U8700 (N_8700,N_8215,N_8462);
nand U8701 (N_8701,N_8162,N_8082);
and U8702 (N_8702,N_8441,N_8484);
nand U8703 (N_8703,N_8385,N_8165);
xnor U8704 (N_8704,N_8424,N_8249);
and U8705 (N_8705,N_8107,N_8125);
nand U8706 (N_8706,N_8435,N_8494);
or U8707 (N_8707,N_8486,N_8338);
xnor U8708 (N_8708,N_8084,N_8267);
nor U8709 (N_8709,N_8496,N_8077);
or U8710 (N_8710,N_8026,N_8466);
and U8711 (N_8711,N_8197,N_8055);
nand U8712 (N_8712,N_8407,N_8114);
or U8713 (N_8713,N_8445,N_8106);
and U8714 (N_8714,N_8460,N_8231);
xor U8715 (N_8715,N_8452,N_8409);
xnor U8716 (N_8716,N_8297,N_8118);
xor U8717 (N_8717,N_8368,N_8305);
xor U8718 (N_8718,N_8037,N_8330);
or U8719 (N_8719,N_8248,N_8200);
nand U8720 (N_8720,N_8041,N_8252);
and U8721 (N_8721,N_8393,N_8351);
or U8722 (N_8722,N_8373,N_8232);
xor U8723 (N_8723,N_8413,N_8386);
xor U8724 (N_8724,N_8128,N_8187);
or U8725 (N_8725,N_8132,N_8075);
xnor U8726 (N_8726,N_8254,N_8316);
or U8727 (N_8727,N_8244,N_8367);
xor U8728 (N_8728,N_8270,N_8448);
xor U8729 (N_8729,N_8159,N_8261);
nand U8730 (N_8730,N_8057,N_8212);
or U8731 (N_8731,N_8423,N_8223);
nand U8732 (N_8732,N_8047,N_8273);
or U8733 (N_8733,N_8000,N_8347);
or U8734 (N_8734,N_8224,N_8337);
or U8735 (N_8735,N_8262,N_8130);
or U8736 (N_8736,N_8184,N_8085);
and U8737 (N_8737,N_8193,N_8168);
or U8738 (N_8738,N_8027,N_8002);
or U8739 (N_8739,N_8382,N_8328);
or U8740 (N_8740,N_8266,N_8092);
nand U8741 (N_8741,N_8015,N_8499);
nor U8742 (N_8742,N_8444,N_8066);
and U8743 (N_8743,N_8255,N_8059);
or U8744 (N_8744,N_8058,N_8463);
xnor U8745 (N_8745,N_8274,N_8283);
nand U8746 (N_8746,N_8113,N_8135);
or U8747 (N_8747,N_8490,N_8051);
nor U8748 (N_8748,N_8378,N_8208);
and U8749 (N_8749,N_8065,N_8336);
or U8750 (N_8750,N_8185,N_8256);
or U8751 (N_8751,N_8434,N_8396);
and U8752 (N_8752,N_8322,N_8218);
nor U8753 (N_8753,N_8081,N_8082);
nor U8754 (N_8754,N_8400,N_8020);
nand U8755 (N_8755,N_8429,N_8073);
xnor U8756 (N_8756,N_8298,N_8185);
and U8757 (N_8757,N_8457,N_8353);
and U8758 (N_8758,N_8475,N_8267);
xor U8759 (N_8759,N_8308,N_8411);
xnor U8760 (N_8760,N_8226,N_8041);
or U8761 (N_8761,N_8499,N_8331);
nor U8762 (N_8762,N_8290,N_8024);
and U8763 (N_8763,N_8128,N_8191);
xnor U8764 (N_8764,N_8425,N_8364);
nor U8765 (N_8765,N_8171,N_8157);
xnor U8766 (N_8766,N_8066,N_8206);
xor U8767 (N_8767,N_8136,N_8181);
nor U8768 (N_8768,N_8401,N_8205);
xor U8769 (N_8769,N_8449,N_8171);
xnor U8770 (N_8770,N_8477,N_8308);
and U8771 (N_8771,N_8082,N_8445);
and U8772 (N_8772,N_8273,N_8017);
and U8773 (N_8773,N_8260,N_8466);
or U8774 (N_8774,N_8182,N_8044);
and U8775 (N_8775,N_8459,N_8478);
nor U8776 (N_8776,N_8363,N_8377);
and U8777 (N_8777,N_8421,N_8287);
nor U8778 (N_8778,N_8454,N_8177);
nor U8779 (N_8779,N_8011,N_8054);
xnor U8780 (N_8780,N_8216,N_8186);
and U8781 (N_8781,N_8473,N_8050);
or U8782 (N_8782,N_8453,N_8263);
nor U8783 (N_8783,N_8114,N_8416);
nor U8784 (N_8784,N_8000,N_8479);
xnor U8785 (N_8785,N_8223,N_8417);
and U8786 (N_8786,N_8309,N_8317);
nand U8787 (N_8787,N_8417,N_8032);
xnor U8788 (N_8788,N_8181,N_8469);
and U8789 (N_8789,N_8037,N_8283);
or U8790 (N_8790,N_8154,N_8300);
and U8791 (N_8791,N_8184,N_8216);
and U8792 (N_8792,N_8077,N_8036);
nand U8793 (N_8793,N_8493,N_8188);
and U8794 (N_8794,N_8210,N_8211);
or U8795 (N_8795,N_8489,N_8129);
or U8796 (N_8796,N_8459,N_8073);
xor U8797 (N_8797,N_8327,N_8242);
xnor U8798 (N_8798,N_8426,N_8359);
or U8799 (N_8799,N_8247,N_8135);
nor U8800 (N_8800,N_8095,N_8421);
nand U8801 (N_8801,N_8142,N_8151);
and U8802 (N_8802,N_8116,N_8375);
or U8803 (N_8803,N_8488,N_8061);
nor U8804 (N_8804,N_8480,N_8447);
xnor U8805 (N_8805,N_8096,N_8404);
nand U8806 (N_8806,N_8020,N_8309);
and U8807 (N_8807,N_8455,N_8405);
xor U8808 (N_8808,N_8487,N_8347);
and U8809 (N_8809,N_8408,N_8315);
xnor U8810 (N_8810,N_8049,N_8285);
nor U8811 (N_8811,N_8265,N_8156);
or U8812 (N_8812,N_8071,N_8137);
nand U8813 (N_8813,N_8374,N_8325);
or U8814 (N_8814,N_8194,N_8299);
or U8815 (N_8815,N_8422,N_8365);
and U8816 (N_8816,N_8215,N_8246);
nor U8817 (N_8817,N_8180,N_8228);
and U8818 (N_8818,N_8176,N_8090);
and U8819 (N_8819,N_8344,N_8066);
xnor U8820 (N_8820,N_8275,N_8238);
and U8821 (N_8821,N_8162,N_8481);
xnor U8822 (N_8822,N_8193,N_8452);
xor U8823 (N_8823,N_8358,N_8130);
nor U8824 (N_8824,N_8469,N_8130);
xor U8825 (N_8825,N_8331,N_8389);
and U8826 (N_8826,N_8408,N_8003);
nor U8827 (N_8827,N_8120,N_8414);
nand U8828 (N_8828,N_8369,N_8492);
nor U8829 (N_8829,N_8047,N_8348);
nor U8830 (N_8830,N_8279,N_8487);
xor U8831 (N_8831,N_8379,N_8275);
nand U8832 (N_8832,N_8477,N_8386);
nand U8833 (N_8833,N_8034,N_8201);
nand U8834 (N_8834,N_8315,N_8373);
nand U8835 (N_8835,N_8303,N_8014);
and U8836 (N_8836,N_8366,N_8146);
nand U8837 (N_8837,N_8237,N_8330);
xnor U8838 (N_8838,N_8470,N_8287);
and U8839 (N_8839,N_8426,N_8486);
nor U8840 (N_8840,N_8411,N_8219);
nand U8841 (N_8841,N_8176,N_8268);
or U8842 (N_8842,N_8261,N_8286);
xnor U8843 (N_8843,N_8398,N_8364);
nor U8844 (N_8844,N_8110,N_8333);
and U8845 (N_8845,N_8227,N_8416);
xnor U8846 (N_8846,N_8293,N_8171);
and U8847 (N_8847,N_8052,N_8220);
nor U8848 (N_8848,N_8011,N_8127);
nand U8849 (N_8849,N_8184,N_8339);
and U8850 (N_8850,N_8161,N_8331);
or U8851 (N_8851,N_8288,N_8366);
xnor U8852 (N_8852,N_8334,N_8366);
nor U8853 (N_8853,N_8128,N_8354);
xor U8854 (N_8854,N_8470,N_8375);
and U8855 (N_8855,N_8018,N_8297);
and U8856 (N_8856,N_8486,N_8264);
nor U8857 (N_8857,N_8207,N_8012);
xor U8858 (N_8858,N_8225,N_8153);
or U8859 (N_8859,N_8423,N_8408);
or U8860 (N_8860,N_8090,N_8386);
and U8861 (N_8861,N_8009,N_8454);
or U8862 (N_8862,N_8424,N_8280);
or U8863 (N_8863,N_8037,N_8175);
nand U8864 (N_8864,N_8347,N_8032);
and U8865 (N_8865,N_8170,N_8270);
and U8866 (N_8866,N_8335,N_8216);
nor U8867 (N_8867,N_8105,N_8342);
and U8868 (N_8868,N_8063,N_8002);
nand U8869 (N_8869,N_8213,N_8300);
nor U8870 (N_8870,N_8192,N_8015);
and U8871 (N_8871,N_8378,N_8011);
and U8872 (N_8872,N_8211,N_8412);
or U8873 (N_8873,N_8268,N_8414);
xor U8874 (N_8874,N_8404,N_8064);
nor U8875 (N_8875,N_8070,N_8201);
or U8876 (N_8876,N_8263,N_8027);
xnor U8877 (N_8877,N_8232,N_8236);
and U8878 (N_8878,N_8046,N_8234);
or U8879 (N_8879,N_8095,N_8382);
or U8880 (N_8880,N_8309,N_8242);
or U8881 (N_8881,N_8068,N_8118);
xnor U8882 (N_8882,N_8307,N_8081);
xor U8883 (N_8883,N_8234,N_8230);
and U8884 (N_8884,N_8184,N_8354);
nand U8885 (N_8885,N_8176,N_8487);
nand U8886 (N_8886,N_8154,N_8387);
nor U8887 (N_8887,N_8440,N_8136);
nand U8888 (N_8888,N_8069,N_8396);
xor U8889 (N_8889,N_8295,N_8333);
and U8890 (N_8890,N_8375,N_8165);
or U8891 (N_8891,N_8481,N_8360);
or U8892 (N_8892,N_8355,N_8447);
xor U8893 (N_8893,N_8397,N_8112);
nand U8894 (N_8894,N_8041,N_8394);
xnor U8895 (N_8895,N_8456,N_8220);
or U8896 (N_8896,N_8313,N_8088);
and U8897 (N_8897,N_8214,N_8451);
and U8898 (N_8898,N_8037,N_8483);
nor U8899 (N_8899,N_8214,N_8136);
or U8900 (N_8900,N_8193,N_8441);
and U8901 (N_8901,N_8363,N_8383);
nor U8902 (N_8902,N_8287,N_8255);
nor U8903 (N_8903,N_8373,N_8275);
and U8904 (N_8904,N_8188,N_8019);
or U8905 (N_8905,N_8018,N_8396);
nand U8906 (N_8906,N_8311,N_8070);
xnor U8907 (N_8907,N_8126,N_8420);
and U8908 (N_8908,N_8371,N_8115);
nand U8909 (N_8909,N_8217,N_8002);
nand U8910 (N_8910,N_8374,N_8353);
nor U8911 (N_8911,N_8182,N_8073);
or U8912 (N_8912,N_8244,N_8404);
nor U8913 (N_8913,N_8055,N_8432);
nand U8914 (N_8914,N_8103,N_8470);
or U8915 (N_8915,N_8193,N_8277);
and U8916 (N_8916,N_8119,N_8393);
and U8917 (N_8917,N_8416,N_8164);
or U8918 (N_8918,N_8461,N_8294);
xor U8919 (N_8919,N_8432,N_8167);
and U8920 (N_8920,N_8004,N_8106);
and U8921 (N_8921,N_8131,N_8075);
xnor U8922 (N_8922,N_8359,N_8476);
or U8923 (N_8923,N_8314,N_8264);
nand U8924 (N_8924,N_8153,N_8484);
nor U8925 (N_8925,N_8294,N_8373);
nor U8926 (N_8926,N_8350,N_8168);
and U8927 (N_8927,N_8212,N_8140);
xnor U8928 (N_8928,N_8080,N_8040);
nor U8929 (N_8929,N_8174,N_8037);
and U8930 (N_8930,N_8446,N_8205);
or U8931 (N_8931,N_8324,N_8101);
and U8932 (N_8932,N_8248,N_8072);
or U8933 (N_8933,N_8319,N_8231);
nand U8934 (N_8934,N_8322,N_8351);
or U8935 (N_8935,N_8421,N_8108);
or U8936 (N_8936,N_8462,N_8472);
or U8937 (N_8937,N_8146,N_8007);
xnor U8938 (N_8938,N_8304,N_8466);
xor U8939 (N_8939,N_8457,N_8195);
nand U8940 (N_8940,N_8290,N_8296);
xnor U8941 (N_8941,N_8488,N_8043);
nor U8942 (N_8942,N_8067,N_8453);
and U8943 (N_8943,N_8222,N_8001);
and U8944 (N_8944,N_8419,N_8351);
and U8945 (N_8945,N_8337,N_8494);
nor U8946 (N_8946,N_8206,N_8292);
xnor U8947 (N_8947,N_8286,N_8297);
and U8948 (N_8948,N_8490,N_8297);
or U8949 (N_8949,N_8491,N_8130);
xor U8950 (N_8950,N_8488,N_8354);
nor U8951 (N_8951,N_8272,N_8051);
nand U8952 (N_8952,N_8152,N_8420);
and U8953 (N_8953,N_8089,N_8141);
xor U8954 (N_8954,N_8117,N_8190);
or U8955 (N_8955,N_8391,N_8362);
or U8956 (N_8956,N_8269,N_8452);
xor U8957 (N_8957,N_8491,N_8062);
nor U8958 (N_8958,N_8198,N_8403);
or U8959 (N_8959,N_8469,N_8045);
nand U8960 (N_8960,N_8029,N_8419);
and U8961 (N_8961,N_8021,N_8058);
nor U8962 (N_8962,N_8187,N_8228);
or U8963 (N_8963,N_8184,N_8097);
or U8964 (N_8964,N_8464,N_8105);
or U8965 (N_8965,N_8494,N_8272);
nor U8966 (N_8966,N_8031,N_8444);
nor U8967 (N_8967,N_8193,N_8321);
xor U8968 (N_8968,N_8131,N_8142);
nor U8969 (N_8969,N_8273,N_8236);
nand U8970 (N_8970,N_8183,N_8382);
and U8971 (N_8971,N_8240,N_8142);
and U8972 (N_8972,N_8358,N_8333);
nand U8973 (N_8973,N_8154,N_8117);
nor U8974 (N_8974,N_8155,N_8457);
nor U8975 (N_8975,N_8101,N_8097);
and U8976 (N_8976,N_8465,N_8425);
xnor U8977 (N_8977,N_8350,N_8391);
or U8978 (N_8978,N_8093,N_8283);
nor U8979 (N_8979,N_8347,N_8034);
and U8980 (N_8980,N_8019,N_8208);
or U8981 (N_8981,N_8455,N_8339);
or U8982 (N_8982,N_8419,N_8128);
and U8983 (N_8983,N_8184,N_8361);
nand U8984 (N_8984,N_8042,N_8477);
nor U8985 (N_8985,N_8343,N_8416);
xor U8986 (N_8986,N_8351,N_8308);
nand U8987 (N_8987,N_8487,N_8458);
or U8988 (N_8988,N_8166,N_8118);
or U8989 (N_8989,N_8156,N_8235);
nor U8990 (N_8990,N_8496,N_8448);
or U8991 (N_8991,N_8419,N_8288);
nor U8992 (N_8992,N_8195,N_8102);
nor U8993 (N_8993,N_8340,N_8250);
or U8994 (N_8994,N_8473,N_8031);
nor U8995 (N_8995,N_8292,N_8129);
nor U8996 (N_8996,N_8141,N_8238);
nand U8997 (N_8997,N_8328,N_8169);
nand U8998 (N_8998,N_8190,N_8010);
or U8999 (N_8999,N_8226,N_8014);
or U9000 (N_9000,N_8669,N_8878);
nor U9001 (N_9001,N_8985,N_8573);
nor U9002 (N_9002,N_8677,N_8501);
nor U9003 (N_9003,N_8900,N_8974);
xnor U9004 (N_9004,N_8751,N_8515);
xnor U9005 (N_9005,N_8534,N_8951);
and U9006 (N_9006,N_8858,N_8828);
xnor U9007 (N_9007,N_8724,N_8948);
and U9008 (N_9008,N_8558,N_8904);
nand U9009 (N_9009,N_8770,N_8876);
nand U9010 (N_9010,N_8772,N_8520);
nand U9011 (N_9011,N_8693,N_8964);
and U9012 (N_9012,N_8714,N_8877);
or U9013 (N_9013,N_8711,N_8608);
nand U9014 (N_9014,N_8566,N_8620);
nor U9015 (N_9015,N_8622,N_8969);
nor U9016 (N_9016,N_8519,N_8953);
nor U9017 (N_9017,N_8894,N_8837);
and U9018 (N_9018,N_8710,N_8618);
xnor U9019 (N_9019,N_8797,N_8745);
nand U9020 (N_9020,N_8827,N_8753);
or U9021 (N_9021,N_8958,N_8848);
xor U9022 (N_9022,N_8962,N_8979);
nand U9023 (N_9023,N_8991,N_8800);
nor U9024 (N_9024,N_8606,N_8726);
or U9025 (N_9025,N_8988,N_8756);
nand U9026 (N_9026,N_8532,N_8516);
xor U9027 (N_9027,N_8981,N_8671);
xnor U9028 (N_9028,N_8766,N_8998);
nor U9029 (N_9029,N_8779,N_8597);
or U9030 (N_9030,N_8860,N_8587);
nor U9031 (N_9031,N_8773,N_8783);
or U9032 (N_9032,N_8917,N_8560);
xor U9033 (N_9033,N_8987,N_8862);
or U9034 (N_9034,N_8718,N_8530);
and U9035 (N_9035,N_8752,N_8994);
or U9036 (N_9036,N_8840,N_8518);
or U9037 (N_9037,N_8812,N_8505);
or U9038 (N_9038,N_8905,N_8972);
xor U9039 (N_9039,N_8805,N_8557);
nor U9040 (N_9040,N_8938,N_8742);
nand U9041 (N_9041,N_8562,N_8799);
nor U9042 (N_9042,N_8638,N_8689);
nand U9043 (N_9043,N_8619,N_8910);
and U9044 (N_9044,N_8932,N_8760);
or U9045 (N_9045,N_8621,N_8629);
xor U9046 (N_9046,N_8954,N_8583);
nand U9047 (N_9047,N_8645,N_8959);
nand U9048 (N_9048,N_8913,N_8536);
or U9049 (N_9049,N_8699,N_8685);
nand U9050 (N_9050,N_8814,N_8871);
or U9051 (N_9051,N_8657,N_8684);
xor U9052 (N_9052,N_8648,N_8561);
nor U9053 (N_9053,N_8914,N_8774);
or U9054 (N_9054,N_8603,N_8949);
or U9055 (N_9055,N_8879,N_8895);
nor U9056 (N_9056,N_8723,N_8780);
xor U9057 (N_9057,N_8855,N_8705);
and U9058 (N_9058,N_8983,N_8755);
and U9059 (N_9059,N_8836,N_8874);
or U9060 (N_9060,N_8602,N_8916);
xnor U9061 (N_9061,N_8784,N_8839);
and U9062 (N_9062,N_8738,N_8931);
xor U9063 (N_9063,N_8527,N_8634);
and U9064 (N_9064,N_8844,N_8811);
nand U9065 (N_9065,N_8970,N_8986);
and U9066 (N_9066,N_8864,N_8552);
nand U9067 (N_9067,N_8600,N_8748);
nand U9068 (N_9068,N_8887,N_8731);
and U9069 (N_9069,N_8643,N_8715);
nor U9070 (N_9070,N_8801,N_8502);
or U9071 (N_9071,N_8506,N_8884);
nand U9072 (N_9072,N_8851,N_8513);
or U9073 (N_9073,N_8686,N_8789);
nand U9074 (N_9074,N_8624,N_8984);
nand U9075 (N_9075,N_8806,N_8737);
and U9076 (N_9076,N_8803,N_8713);
nand U9077 (N_9077,N_8509,N_8944);
nand U9078 (N_9078,N_8888,N_8775);
xor U9079 (N_9079,N_8612,N_8907);
and U9080 (N_9080,N_8936,N_8517);
and U9081 (N_9081,N_8886,N_8798);
or U9082 (N_9082,N_8882,N_8842);
and U9083 (N_9083,N_8651,N_8531);
nor U9084 (N_9084,N_8546,N_8673);
or U9085 (N_9085,N_8598,N_8720);
xnor U9086 (N_9086,N_8976,N_8898);
or U9087 (N_9087,N_8540,N_8880);
nand U9088 (N_9088,N_8892,N_8535);
xnor U9089 (N_9089,N_8909,N_8754);
nand U9090 (N_9090,N_8952,N_8529);
nand U9091 (N_9091,N_8630,N_8666);
and U9092 (N_9092,N_8971,N_8746);
and U9093 (N_9093,N_8616,N_8642);
nor U9094 (N_9094,N_8586,N_8615);
or U9095 (N_9095,N_8694,N_8869);
nor U9096 (N_9096,N_8835,N_8596);
or U9097 (N_9097,N_8649,N_8639);
nor U9098 (N_9098,N_8605,N_8792);
or U9099 (N_9099,N_8687,N_8890);
and U9100 (N_9100,N_8730,N_8889);
or U9101 (N_9101,N_8763,N_8701);
and U9102 (N_9102,N_8523,N_8500);
or U9103 (N_9103,N_8940,N_8568);
nand U9104 (N_9104,N_8833,N_8908);
xor U9105 (N_9105,N_8853,N_8729);
nand U9106 (N_9106,N_8607,N_8691);
nand U9107 (N_9107,N_8628,N_8734);
and U9108 (N_9108,N_8967,N_8924);
nand U9109 (N_9109,N_8650,N_8778);
or U9110 (N_9110,N_8740,N_8942);
xnor U9111 (N_9111,N_8928,N_8526);
or U9112 (N_9112,N_8662,N_8989);
nand U9113 (N_9113,N_8982,N_8881);
and U9114 (N_9114,N_8999,N_8845);
or U9115 (N_9115,N_8681,N_8589);
and U9116 (N_9116,N_8926,N_8852);
and U9117 (N_9117,N_8747,N_8863);
nor U9118 (N_9118,N_8764,N_8576);
nor U9119 (N_9119,N_8849,N_8679);
or U9120 (N_9120,N_8721,N_8604);
and U9121 (N_9121,N_8966,N_8593);
nor U9122 (N_9122,N_8857,N_8582);
and U9123 (N_9123,N_8564,N_8594);
or U9124 (N_9124,N_8824,N_8930);
nand U9125 (N_9125,N_8978,N_8539);
nor U9126 (N_9126,N_8595,N_8725);
nand U9127 (N_9127,N_8659,N_8965);
xnor U9128 (N_9128,N_8788,N_8521);
nor U9129 (N_9129,N_8524,N_8556);
and U9130 (N_9130,N_8504,N_8533);
or U9131 (N_9131,N_8588,N_8676);
xnor U9132 (N_9132,N_8759,N_8787);
nand U9133 (N_9133,N_8633,N_8703);
nor U9134 (N_9134,N_8816,N_8941);
nor U9135 (N_9135,N_8765,N_8584);
nand U9136 (N_9136,N_8945,N_8617);
nor U9137 (N_9137,N_8591,N_8743);
nor U9138 (N_9138,N_8717,N_8739);
nand U9139 (N_9139,N_8868,N_8599);
nor U9140 (N_9140,N_8761,N_8777);
nand U9141 (N_9141,N_8667,N_8578);
or U9142 (N_9142,N_8702,N_8990);
or U9143 (N_9143,N_8866,N_8934);
nor U9144 (N_9144,N_8802,N_8522);
or U9145 (N_9145,N_8963,N_8525);
and U9146 (N_9146,N_8911,N_8654);
xor U9147 (N_9147,N_8925,N_8832);
xor U9148 (N_9148,N_8512,N_8867);
and U9149 (N_9149,N_8581,N_8744);
nand U9150 (N_9150,N_8885,N_8810);
xnor U9151 (N_9151,N_8611,N_8712);
xor U9152 (N_9152,N_8683,N_8767);
xor U9153 (N_9153,N_8899,N_8728);
nand U9154 (N_9154,N_8856,N_8897);
nor U9155 (N_9155,N_8793,N_8585);
nand U9156 (N_9156,N_8923,N_8825);
or U9157 (N_9157,N_8538,N_8569);
nor U9158 (N_9158,N_8861,N_8707);
and U9159 (N_9159,N_8809,N_8804);
nand U9160 (N_9160,N_8918,N_8592);
xnor U9161 (N_9161,N_8785,N_8846);
xnor U9162 (N_9162,N_8975,N_8507);
xor U9163 (N_9163,N_8826,N_8946);
nor U9164 (N_9164,N_8996,N_8635);
and U9165 (N_9165,N_8570,N_8510);
xnor U9166 (N_9166,N_8870,N_8841);
and U9167 (N_9167,N_8631,N_8813);
or U9168 (N_9168,N_8661,N_8933);
or U9169 (N_9169,N_8977,N_8609);
nor U9170 (N_9170,N_8716,N_8980);
nand U9171 (N_9171,N_8563,N_8750);
xnor U9172 (N_9172,N_8912,N_8791);
or U9173 (N_9173,N_8947,N_8769);
xor U9174 (N_9174,N_8610,N_8575);
xor U9175 (N_9175,N_8646,N_8697);
nor U9176 (N_9176,N_8819,N_8652);
or U9177 (N_9177,N_8614,N_8993);
nand U9178 (N_9178,N_8854,N_8922);
or U9179 (N_9179,N_8957,N_8950);
or U9180 (N_9180,N_8937,N_8902);
and U9181 (N_9181,N_8572,N_8735);
xnor U9182 (N_9182,N_8919,N_8579);
nor U9183 (N_9183,N_8555,N_8503);
xor U9184 (N_9184,N_8830,N_8786);
nand U9185 (N_9185,N_8927,N_8901);
nand U9186 (N_9186,N_8623,N_8537);
and U9187 (N_9187,N_8554,N_8719);
or U9188 (N_9188,N_8542,N_8665);
or U9189 (N_9189,N_8647,N_8722);
or U9190 (N_9190,N_8807,N_8818);
and U9191 (N_9191,N_8921,N_8843);
nor U9192 (N_9192,N_8995,N_8511);
xor U9193 (N_9193,N_8571,N_8636);
or U9194 (N_9194,N_8758,N_8749);
xor U9195 (N_9195,N_8675,N_8656);
or U9196 (N_9196,N_8961,N_8829);
or U9197 (N_9197,N_8664,N_8653);
or U9198 (N_9198,N_8821,N_8822);
and U9199 (N_9199,N_8762,N_8815);
nor U9200 (N_9200,N_8790,N_8794);
xnor U9201 (N_9201,N_8968,N_8574);
xnor U9202 (N_9202,N_8680,N_8929);
or U9203 (N_9203,N_8960,N_8688);
and U9204 (N_9204,N_8733,N_8590);
xor U9205 (N_9205,N_8709,N_8732);
nand U9206 (N_9206,N_8973,N_8640);
and U9207 (N_9207,N_8943,N_8613);
or U9208 (N_9208,N_8670,N_8674);
xor U9209 (N_9209,N_8655,N_8831);
nand U9210 (N_9210,N_8915,N_8920);
nor U9211 (N_9211,N_8820,N_8808);
and U9212 (N_9212,N_8997,N_8741);
xor U9213 (N_9213,N_8883,N_8906);
nand U9214 (N_9214,N_8865,N_8823);
or U9215 (N_9215,N_8956,N_8939);
and U9216 (N_9216,N_8872,N_8838);
nand U9217 (N_9217,N_8727,N_8796);
and U9218 (N_9218,N_8601,N_8644);
and U9219 (N_9219,N_8708,N_8577);
nor U9220 (N_9220,N_8850,N_8658);
xnor U9221 (N_9221,N_8893,N_8955);
and U9222 (N_9222,N_8781,N_8528);
and U9223 (N_9223,N_8875,N_8549);
nor U9224 (N_9224,N_8696,N_8627);
nand U9225 (N_9225,N_8678,N_8632);
or U9226 (N_9226,N_8847,N_8626);
xnor U9227 (N_9227,N_8668,N_8859);
nand U9228 (N_9228,N_8682,N_8776);
nand U9229 (N_9229,N_8565,N_8543);
nor U9230 (N_9230,N_8690,N_8771);
or U9231 (N_9231,N_8873,N_8551);
or U9232 (N_9232,N_8663,N_8641);
nor U9233 (N_9233,N_8550,N_8935);
nand U9234 (N_9234,N_8757,N_8704);
nand U9235 (N_9235,N_8545,N_8817);
nand U9236 (N_9236,N_8541,N_8514);
nand U9237 (N_9237,N_8567,N_8695);
xor U9238 (N_9238,N_8795,N_8782);
and U9239 (N_9239,N_8637,N_8625);
xnor U9240 (N_9240,N_8692,N_8834);
or U9241 (N_9241,N_8903,N_8706);
or U9242 (N_9242,N_8559,N_8553);
xor U9243 (N_9243,N_8768,N_8508);
and U9244 (N_9244,N_8660,N_8891);
or U9245 (N_9245,N_8992,N_8580);
nand U9246 (N_9246,N_8896,N_8698);
or U9247 (N_9247,N_8736,N_8672);
and U9248 (N_9248,N_8547,N_8700);
nor U9249 (N_9249,N_8544,N_8548);
nand U9250 (N_9250,N_8793,N_8744);
nor U9251 (N_9251,N_8733,N_8792);
nand U9252 (N_9252,N_8783,N_8545);
nand U9253 (N_9253,N_8659,N_8820);
nor U9254 (N_9254,N_8834,N_8518);
or U9255 (N_9255,N_8866,N_8585);
xnor U9256 (N_9256,N_8723,N_8819);
and U9257 (N_9257,N_8717,N_8892);
nand U9258 (N_9258,N_8902,N_8899);
and U9259 (N_9259,N_8576,N_8691);
nor U9260 (N_9260,N_8507,N_8832);
or U9261 (N_9261,N_8754,N_8518);
and U9262 (N_9262,N_8811,N_8940);
nor U9263 (N_9263,N_8989,N_8528);
xor U9264 (N_9264,N_8529,N_8669);
or U9265 (N_9265,N_8976,N_8841);
or U9266 (N_9266,N_8507,N_8697);
and U9267 (N_9267,N_8778,N_8654);
or U9268 (N_9268,N_8803,N_8596);
xnor U9269 (N_9269,N_8746,N_8857);
xor U9270 (N_9270,N_8816,N_8993);
and U9271 (N_9271,N_8744,N_8976);
and U9272 (N_9272,N_8699,N_8928);
and U9273 (N_9273,N_8947,N_8962);
and U9274 (N_9274,N_8684,N_8685);
or U9275 (N_9275,N_8780,N_8552);
xnor U9276 (N_9276,N_8536,N_8608);
or U9277 (N_9277,N_8933,N_8870);
nand U9278 (N_9278,N_8935,N_8608);
or U9279 (N_9279,N_8896,N_8954);
xor U9280 (N_9280,N_8936,N_8866);
nor U9281 (N_9281,N_8878,N_8968);
and U9282 (N_9282,N_8812,N_8829);
nor U9283 (N_9283,N_8615,N_8942);
xnor U9284 (N_9284,N_8666,N_8777);
or U9285 (N_9285,N_8699,N_8709);
xor U9286 (N_9286,N_8868,N_8555);
xnor U9287 (N_9287,N_8538,N_8571);
nand U9288 (N_9288,N_8603,N_8792);
xor U9289 (N_9289,N_8772,N_8677);
xor U9290 (N_9290,N_8507,N_8755);
nand U9291 (N_9291,N_8922,N_8818);
and U9292 (N_9292,N_8801,N_8869);
nor U9293 (N_9293,N_8865,N_8534);
nor U9294 (N_9294,N_8750,N_8759);
nand U9295 (N_9295,N_8934,N_8952);
nand U9296 (N_9296,N_8764,N_8900);
or U9297 (N_9297,N_8615,N_8706);
xnor U9298 (N_9298,N_8854,N_8780);
nand U9299 (N_9299,N_8817,N_8544);
or U9300 (N_9300,N_8978,N_8586);
or U9301 (N_9301,N_8769,N_8819);
or U9302 (N_9302,N_8624,N_8831);
xor U9303 (N_9303,N_8536,N_8609);
or U9304 (N_9304,N_8984,N_8651);
and U9305 (N_9305,N_8575,N_8642);
nor U9306 (N_9306,N_8957,N_8808);
and U9307 (N_9307,N_8809,N_8550);
or U9308 (N_9308,N_8561,N_8521);
nor U9309 (N_9309,N_8821,N_8791);
or U9310 (N_9310,N_8527,N_8641);
and U9311 (N_9311,N_8582,N_8577);
or U9312 (N_9312,N_8570,N_8895);
or U9313 (N_9313,N_8557,N_8710);
xnor U9314 (N_9314,N_8805,N_8700);
nand U9315 (N_9315,N_8556,N_8981);
nor U9316 (N_9316,N_8805,N_8511);
and U9317 (N_9317,N_8932,N_8532);
or U9318 (N_9318,N_8921,N_8956);
and U9319 (N_9319,N_8903,N_8692);
and U9320 (N_9320,N_8825,N_8521);
nand U9321 (N_9321,N_8677,N_8551);
nand U9322 (N_9322,N_8571,N_8808);
nand U9323 (N_9323,N_8574,N_8707);
xor U9324 (N_9324,N_8584,N_8641);
xnor U9325 (N_9325,N_8894,N_8705);
nand U9326 (N_9326,N_8890,N_8649);
xor U9327 (N_9327,N_8738,N_8831);
nor U9328 (N_9328,N_8791,N_8745);
nor U9329 (N_9329,N_8928,N_8744);
or U9330 (N_9330,N_8512,N_8593);
and U9331 (N_9331,N_8632,N_8753);
nand U9332 (N_9332,N_8980,N_8902);
and U9333 (N_9333,N_8777,N_8890);
nand U9334 (N_9334,N_8979,N_8605);
xnor U9335 (N_9335,N_8687,N_8898);
xor U9336 (N_9336,N_8995,N_8709);
or U9337 (N_9337,N_8598,N_8976);
or U9338 (N_9338,N_8987,N_8968);
xor U9339 (N_9339,N_8875,N_8625);
nand U9340 (N_9340,N_8911,N_8699);
xor U9341 (N_9341,N_8917,N_8982);
nand U9342 (N_9342,N_8735,N_8772);
or U9343 (N_9343,N_8841,N_8788);
or U9344 (N_9344,N_8938,N_8574);
xnor U9345 (N_9345,N_8590,N_8991);
and U9346 (N_9346,N_8744,N_8589);
nand U9347 (N_9347,N_8504,N_8912);
and U9348 (N_9348,N_8533,N_8906);
xor U9349 (N_9349,N_8703,N_8940);
nand U9350 (N_9350,N_8769,N_8567);
nor U9351 (N_9351,N_8946,N_8647);
nor U9352 (N_9352,N_8723,N_8921);
xor U9353 (N_9353,N_8600,N_8959);
and U9354 (N_9354,N_8900,N_8530);
nor U9355 (N_9355,N_8981,N_8706);
or U9356 (N_9356,N_8550,N_8768);
nand U9357 (N_9357,N_8974,N_8995);
nand U9358 (N_9358,N_8837,N_8849);
and U9359 (N_9359,N_8834,N_8989);
nor U9360 (N_9360,N_8527,N_8750);
nand U9361 (N_9361,N_8941,N_8887);
nor U9362 (N_9362,N_8676,N_8948);
and U9363 (N_9363,N_8957,N_8799);
nand U9364 (N_9364,N_8921,N_8893);
xnor U9365 (N_9365,N_8722,N_8531);
and U9366 (N_9366,N_8644,N_8822);
and U9367 (N_9367,N_8596,N_8920);
xor U9368 (N_9368,N_8929,N_8526);
nand U9369 (N_9369,N_8902,N_8642);
and U9370 (N_9370,N_8569,N_8658);
or U9371 (N_9371,N_8958,N_8584);
and U9372 (N_9372,N_8753,N_8696);
nor U9373 (N_9373,N_8682,N_8749);
nand U9374 (N_9374,N_8978,N_8691);
nand U9375 (N_9375,N_8978,N_8952);
xor U9376 (N_9376,N_8834,N_8745);
nand U9377 (N_9377,N_8500,N_8640);
and U9378 (N_9378,N_8616,N_8835);
nor U9379 (N_9379,N_8535,N_8814);
xnor U9380 (N_9380,N_8995,N_8923);
and U9381 (N_9381,N_8900,N_8759);
or U9382 (N_9382,N_8580,N_8834);
xnor U9383 (N_9383,N_8565,N_8662);
and U9384 (N_9384,N_8805,N_8766);
xor U9385 (N_9385,N_8850,N_8909);
or U9386 (N_9386,N_8625,N_8565);
and U9387 (N_9387,N_8732,N_8586);
nor U9388 (N_9388,N_8576,N_8607);
or U9389 (N_9389,N_8824,N_8704);
and U9390 (N_9390,N_8725,N_8905);
nor U9391 (N_9391,N_8548,N_8801);
xnor U9392 (N_9392,N_8909,N_8601);
nor U9393 (N_9393,N_8908,N_8642);
or U9394 (N_9394,N_8958,N_8673);
or U9395 (N_9395,N_8549,N_8544);
nor U9396 (N_9396,N_8640,N_8514);
and U9397 (N_9397,N_8549,N_8945);
nor U9398 (N_9398,N_8751,N_8902);
xor U9399 (N_9399,N_8813,N_8871);
xnor U9400 (N_9400,N_8800,N_8957);
xor U9401 (N_9401,N_8816,N_8902);
xor U9402 (N_9402,N_8569,N_8885);
nor U9403 (N_9403,N_8962,N_8839);
and U9404 (N_9404,N_8587,N_8740);
xor U9405 (N_9405,N_8906,N_8775);
nor U9406 (N_9406,N_8826,N_8515);
and U9407 (N_9407,N_8845,N_8589);
nand U9408 (N_9408,N_8975,N_8974);
xor U9409 (N_9409,N_8862,N_8648);
nand U9410 (N_9410,N_8726,N_8788);
xor U9411 (N_9411,N_8962,N_8801);
or U9412 (N_9412,N_8731,N_8939);
nor U9413 (N_9413,N_8968,N_8737);
nor U9414 (N_9414,N_8947,N_8508);
and U9415 (N_9415,N_8944,N_8850);
nor U9416 (N_9416,N_8985,N_8595);
nand U9417 (N_9417,N_8696,N_8607);
or U9418 (N_9418,N_8814,N_8751);
and U9419 (N_9419,N_8795,N_8915);
or U9420 (N_9420,N_8779,N_8950);
or U9421 (N_9421,N_8675,N_8653);
xnor U9422 (N_9422,N_8924,N_8949);
xnor U9423 (N_9423,N_8736,N_8890);
or U9424 (N_9424,N_8713,N_8800);
xnor U9425 (N_9425,N_8622,N_8577);
xor U9426 (N_9426,N_8726,N_8735);
or U9427 (N_9427,N_8633,N_8984);
and U9428 (N_9428,N_8838,N_8607);
or U9429 (N_9429,N_8775,N_8908);
nor U9430 (N_9430,N_8877,N_8957);
nand U9431 (N_9431,N_8601,N_8816);
and U9432 (N_9432,N_8531,N_8938);
xnor U9433 (N_9433,N_8839,N_8865);
nor U9434 (N_9434,N_8688,N_8530);
nor U9435 (N_9435,N_8525,N_8777);
and U9436 (N_9436,N_8692,N_8864);
and U9437 (N_9437,N_8710,N_8617);
or U9438 (N_9438,N_8835,N_8597);
nand U9439 (N_9439,N_8754,N_8883);
or U9440 (N_9440,N_8656,N_8730);
nor U9441 (N_9441,N_8848,N_8937);
and U9442 (N_9442,N_8998,N_8749);
and U9443 (N_9443,N_8862,N_8709);
and U9444 (N_9444,N_8886,N_8992);
nor U9445 (N_9445,N_8901,N_8689);
nand U9446 (N_9446,N_8848,N_8713);
nor U9447 (N_9447,N_8625,N_8911);
and U9448 (N_9448,N_8957,N_8820);
nor U9449 (N_9449,N_8567,N_8835);
xnor U9450 (N_9450,N_8718,N_8725);
xnor U9451 (N_9451,N_8851,N_8604);
and U9452 (N_9452,N_8600,N_8794);
nor U9453 (N_9453,N_8524,N_8952);
and U9454 (N_9454,N_8645,N_8870);
and U9455 (N_9455,N_8564,N_8661);
nor U9456 (N_9456,N_8931,N_8904);
or U9457 (N_9457,N_8747,N_8627);
and U9458 (N_9458,N_8919,N_8899);
nor U9459 (N_9459,N_8994,N_8713);
and U9460 (N_9460,N_8867,N_8712);
nand U9461 (N_9461,N_8940,N_8742);
nand U9462 (N_9462,N_8808,N_8921);
nand U9463 (N_9463,N_8944,N_8676);
nand U9464 (N_9464,N_8934,N_8911);
nand U9465 (N_9465,N_8803,N_8929);
nand U9466 (N_9466,N_8812,N_8988);
nand U9467 (N_9467,N_8584,N_8734);
nand U9468 (N_9468,N_8844,N_8568);
nor U9469 (N_9469,N_8973,N_8560);
nor U9470 (N_9470,N_8522,N_8687);
xor U9471 (N_9471,N_8744,N_8820);
or U9472 (N_9472,N_8805,N_8787);
xor U9473 (N_9473,N_8710,N_8742);
xor U9474 (N_9474,N_8765,N_8979);
nor U9475 (N_9475,N_8694,N_8582);
nor U9476 (N_9476,N_8794,N_8672);
and U9477 (N_9477,N_8647,N_8821);
nand U9478 (N_9478,N_8689,N_8968);
nor U9479 (N_9479,N_8534,N_8846);
and U9480 (N_9480,N_8718,N_8975);
or U9481 (N_9481,N_8641,N_8631);
xor U9482 (N_9482,N_8550,N_8770);
and U9483 (N_9483,N_8738,N_8851);
xor U9484 (N_9484,N_8742,N_8650);
xnor U9485 (N_9485,N_8899,N_8657);
nor U9486 (N_9486,N_8803,N_8760);
nand U9487 (N_9487,N_8823,N_8752);
and U9488 (N_9488,N_8672,N_8692);
or U9489 (N_9489,N_8886,N_8988);
xnor U9490 (N_9490,N_8949,N_8819);
or U9491 (N_9491,N_8861,N_8764);
nor U9492 (N_9492,N_8722,N_8811);
xnor U9493 (N_9493,N_8643,N_8778);
nand U9494 (N_9494,N_8986,N_8727);
or U9495 (N_9495,N_8990,N_8767);
nand U9496 (N_9496,N_8512,N_8533);
nand U9497 (N_9497,N_8583,N_8849);
nand U9498 (N_9498,N_8589,N_8915);
and U9499 (N_9499,N_8716,N_8657);
or U9500 (N_9500,N_9178,N_9438);
or U9501 (N_9501,N_9246,N_9453);
nor U9502 (N_9502,N_9160,N_9034);
nor U9503 (N_9503,N_9465,N_9389);
nand U9504 (N_9504,N_9352,N_9461);
nor U9505 (N_9505,N_9113,N_9027);
or U9506 (N_9506,N_9316,N_9054);
or U9507 (N_9507,N_9159,N_9230);
nand U9508 (N_9508,N_9399,N_9362);
nor U9509 (N_9509,N_9142,N_9222);
xnor U9510 (N_9510,N_9340,N_9294);
or U9511 (N_9511,N_9249,N_9244);
nor U9512 (N_9512,N_9322,N_9212);
or U9513 (N_9513,N_9351,N_9006);
xnor U9514 (N_9514,N_9470,N_9037);
nand U9515 (N_9515,N_9269,N_9187);
xnor U9516 (N_9516,N_9121,N_9384);
nand U9517 (N_9517,N_9432,N_9281);
or U9518 (N_9518,N_9098,N_9161);
and U9519 (N_9519,N_9140,N_9395);
or U9520 (N_9520,N_9185,N_9261);
and U9521 (N_9521,N_9000,N_9063);
and U9522 (N_9522,N_9367,N_9218);
xnor U9523 (N_9523,N_9475,N_9349);
xor U9524 (N_9524,N_9495,N_9048);
xor U9525 (N_9525,N_9297,N_9401);
xnor U9526 (N_9526,N_9118,N_9286);
xor U9527 (N_9527,N_9100,N_9266);
nor U9528 (N_9528,N_9107,N_9087);
nor U9529 (N_9529,N_9138,N_9109);
xor U9530 (N_9530,N_9035,N_9152);
and U9531 (N_9531,N_9471,N_9365);
nor U9532 (N_9532,N_9179,N_9278);
nand U9533 (N_9533,N_9148,N_9439);
or U9534 (N_9534,N_9386,N_9491);
nand U9535 (N_9535,N_9477,N_9426);
nand U9536 (N_9536,N_9213,N_9420);
nand U9537 (N_9537,N_9225,N_9162);
nor U9538 (N_9538,N_9361,N_9317);
nand U9539 (N_9539,N_9102,N_9117);
or U9540 (N_9540,N_9207,N_9364);
or U9541 (N_9541,N_9277,N_9283);
xnor U9542 (N_9542,N_9088,N_9354);
and U9543 (N_9543,N_9074,N_9265);
and U9544 (N_9544,N_9275,N_9315);
xnor U9545 (N_9545,N_9350,N_9338);
xnor U9546 (N_9546,N_9360,N_9196);
nand U9547 (N_9547,N_9312,N_9070);
and U9548 (N_9548,N_9156,N_9072);
nand U9549 (N_9549,N_9309,N_9190);
nor U9550 (N_9550,N_9032,N_9154);
or U9551 (N_9551,N_9067,N_9268);
nor U9552 (N_9552,N_9305,N_9062);
or U9553 (N_9553,N_9488,N_9262);
xor U9554 (N_9554,N_9056,N_9176);
or U9555 (N_9555,N_9443,N_9164);
nand U9556 (N_9556,N_9293,N_9104);
nand U9557 (N_9557,N_9031,N_9163);
xnor U9558 (N_9558,N_9348,N_9095);
or U9559 (N_9559,N_9137,N_9481);
and U9560 (N_9560,N_9436,N_9084);
nand U9561 (N_9561,N_9221,N_9479);
nor U9562 (N_9562,N_9450,N_9357);
nand U9563 (N_9563,N_9096,N_9325);
xor U9564 (N_9564,N_9380,N_9374);
and U9565 (N_9565,N_9373,N_9289);
nor U9566 (N_9566,N_9009,N_9235);
or U9567 (N_9567,N_9310,N_9066);
nand U9568 (N_9568,N_9369,N_9451);
xor U9569 (N_9569,N_9129,N_9279);
xor U9570 (N_9570,N_9051,N_9007);
nand U9571 (N_9571,N_9366,N_9347);
nand U9572 (N_9572,N_9460,N_9273);
nand U9573 (N_9573,N_9363,N_9149);
xor U9574 (N_9574,N_9346,N_9206);
nand U9575 (N_9575,N_9445,N_9321);
and U9576 (N_9576,N_9257,N_9301);
and U9577 (N_9577,N_9043,N_9039);
or U9578 (N_9578,N_9248,N_9433);
and U9579 (N_9579,N_9409,N_9318);
xor U9580 (N_9580,N_9157,N_9329);
xnor U9581 (N_9581,N_9038,N_9252);
nand U9582 (N_9582,N_9448,N_9308);
nor U9583 (N_9583,N_9036,N_9328);
nor U9584 (N_9584,N_9482,N_9444);
xor U9585 (N_9585,N_9476,N_9280);
nor U9586 (N_9586,N_9334,N_9175);
nand U9587 (N_9587,N_9441,N_9105);
or U9588 (N_9588,N_9402,N_9424);
or U9589 (N_9589,N_9320,N_9091);
and U9590 (N_9590,N_9492,N_9274);
nand U9591 (N_9591,N_9342,N_9040);
nor U9592 (N_9592,N_9458,N_9016);
or U9593 (N_9593,N_9023,N_9064);
nand U9594 (N_9594,N_9430,N_9180);
nor U9595 (N_9595,N_9473,N_9122);
nand U9596 (N_9596,N_9123,N_9454);
xor U9597 (N_9597,N_9172,N_9391);
and U9598 (N_9598,N_9189,N_9429);
nor U9599 (N_9599,N_9025,N_9397);
nand U9600 (N_9600,N_9018,N_9004);
nor U9601 (N_9601,N_9171,N_9082);
nor U9602 (N_9602,N_9131,N_9215);
nand U9603 (N_9603,N_9272,N_9422);
and U9604 (N_9604,N_9169,N_9073);
or U9605 (N_9605,N_9353,N_9344);
nor U9606 (N_9606,N_9290,N_9300);
and U9607 (N_9607,N_9400,N_9396);
nand U9608 (N_9608,N_9153,N_9241);
and U9609 (N_9609,N_9228,N_9442);
xnor U9610 (N_9610,N_9437,N_9217);
or U9611 (N_9611,N_9144,N_9472);
and U9612 (N_9612,N_9201,N_9114);
and U9613 (N_9613,N_9489,N_9327);
and U9614 (N_9614,N_9143,N_9381);
nor U9615 (N_9615,N_9242,N_9141);
and U9616 (N_9616,N_9498,N_9449);
and U9617 (N_9617,N_9227,N_9194);
or U9618 (N_9618,N_9343,N_9387);
nand U9619 (N_9619,N_9053,N_9403);
xor U9620 (N_9620,N_9182,N_9464);
xnor U9621 (N_9621,N_9166,N_9306);
nand U9622 (N_9622,N_9484,N_9077);
nor U9623 (N_9623,N_9052,N_9015);
and U9624 (N_9624,N_9013,N_9417);
and U9625 (N_9625,N_9174,N_9247);
and U9626 (N_9626,N_9223,N_9145);
xor U9627 (N_9627,N_9003,N_9239);
nand U9628 (N_9628,N_9057,N_9370);
and U9629 (N_9629,N_9427,N_9184);
xor U9630 (N_9630,N_9251,N_9295);
xnor U9631 (N_9631,N_9382,N_9001);
and U9632 (N_9632,N_9155,N_9012);
nor U9633 (N_9633,N_9292,N_9368);
nand U9634 (N_9634,N_9326,N_9355);
or U9635 (N_9635,N_9462,N_9250);
xnor U9636 (N_9636,N_9068,N_9376);
and U9637 (N_9637,N_9493,N_9177);
nor U9638 (N_9638,N_9419,N_9094);
nand U9639 (N_9639,N_9276,N_9005);
xnor U9640 (N_9640,N_9020,N_9455);
nand U9641 (N_9641,N_9393,N_9423);
nand U9642 (N_9642,N_9336,N_9385);
nand U9643 (N_9643,N_9256,N_9496);
xnor U9644 (N_9644,N_9047,N_9079);
and U9645 (N_9645,N_9049,N_9377);
nor U9646 (N_9646,N_9134,N_9126);
and U9647 (N_9647,N_9214,N_9099);
nand U9648 (N_9648,N_9410,N_9209);
or U9649 (N_9649,N_9490,N_9264);
xor U9650 (N_9650,N_9447,N_9407);
or U9651 (N_9651,N_9093,N_9135);
xnor U9652 (N_9652,N_9486,N_9375);
nand U9653 (N_9653,N_9383,N_9390);
nor U9654 (N_9654,N_9237,N_9452);
and U9655 (N_9655,N_9243,N_9487);
and U9656 (N_9656,N_9434,N_9319);
nand U9657 (N_9657,N_9245,N_9284);
or U9658 (N_9658,N_9128,N_9089);
xor U9659 (N_9659,N_9372,N_9081);
xor U9660 (N_9660,N_9071,N_9080);
xor U9661 (N_9661,N_9440,N_9119);
nor U9662 (N_9662,N_9229,N_9467);
nand U9663 (N_9663,N_9226,N_9075);
or U9664 (N_9664,N_9263,N_9002);
xor U9665 (N_9665,N_9466,N_9193);
nand U9666 (N_9666,N_9483,N_9045);
and U9667 (N_9667,N_9050,N_9158);
nand U9668 (N_9668,N_9415,N_9323);
or U9669 (N_9669,N_9147,N_9435);
nand U9670 (N_9670,N_9398,N_9203);
xor U9671 (N_9671,N_9008,N_9202);
or U9672 (N_9672,N_9431,N_9033);
xor U9673 (N_9673,N_9414,N_9287);
or U9674 (N_9674,N_9041,N_9494);
or U9675 (N_9675,N_9210,N_9186);
and U9676 (N_9676,N_9115,N_9028);
and U9677 (N_9677,N_9026,N_9059);
xor U9678 (N_9678,N_9061,N_9331);
xnor U9679 (N_9679,N_9330,N_9236);
xnor U9680 (N_9680,N_9224,N_9371);
nand U9681 (N_9681,N_9234,N_9307);
and U9682 (N_9682,N_9112,N_9181);
or U9683 (N_9683,N_9388,N_9055);
and U9684 (N_9684,N_9200,N_9103);
nand U9685 (N_9685,N_9233,N_9024);
xor U9686 (N_9686,N_9042,N_9133);
or U9687 (N_9687,N_9416,N_9165);
nand U9688 (N_9688,N_9232,N_9267);
xnor U9689 (N_9689,N_9299,N_9069);
xnor U9690 (N_9690,N_9463,N_9421);
and U9691 (N_9691,N_9204,N_9345);
xnor U9692 (N_9692,N_9120,N_9205);
and U9693 (N_9693,N_9271,N_9044);
nor U9694 (N_9694,N_9311,N_9046);
or U9695 (N_9695,N_9335,N_9425);
and U9696 (N_9696,N_9499,N_9379);
xor U9697 (N_9697,N_9468,N_9092);
nor U9698 (N_9698,N_9394,N_9240);
nand U9699 (N_9699,N_9168,N_9456);
xnor U9700 (N_9700,N_9459,N_9405);
nand U9701 (N_9701,N_9085,N_9378);
nand U9702 (N_9702,N_9136,N_9296);
and U9703 (N_9703,N_9220,N_9192);
nor U9704 (N_9704,N_9197,N_9198);
and U9705 (N_9705,N_9358,N_9413);
nor U9706 (N_9706,N_9078,N_9339);
xnor U9707 (N_9707,N_9259,N_9058);
xnor U9708 (N_9708,N_9288,N_9108);
nand U9709 (N_9709,N_9076,N_9332);
or U9710 (N_9710,N_9337,N_9208);
nand U9711 (N_9711,N_9116,N_9151);
or U9712 (N_9712,N_9457,N_9480);
and U9713 (N_9713,N_9086,N_9406);
nand U9714 (N_9714,N_9132,N_9412);
or U9715 (N_9715,N_9183,N_9010);
nand U9716 (N_9716,N_9188,N_9497);
and U9717 (N_9717,N_9392,N_9474);
xor U9718 (N_9718,N_9060,N_9173);
nand U9719 (N_9719,N_9341,N_9285);
xor U9720 (N_9720,N_9021,N_9324);
or U9721 (N_9721,N_9097,N_9022);
nor U9722 (N_9722,N_9408,N_9170);
nand U9723 (N_9723,N_9030,N_9313);
nor U9724 (N_9724,N_9139,N_9258);
xor U9725 (N_9725,N_9110,N_9211);
or U9726 (N_9726,N_9333,N_9199);
nand U9727 (N_9727,N_9359,N_9304);
nand U9728 (N_9728,N_9146,N_9418);
xor U9729 (N_9729,N_9260,N_9191);
nand U9730 (N_9730,N_9101,N_9124);
nand U9731 (N_9731,N_9019,N_9111);
nand U9732 (N_9732,N_9195,N_9253);
nor U9733 (N_9733,N_9127,N_9090);
and U9734 (N_9734,N_9029,N_9106);
nor U9735 (N_9735,N_9282,N_9254);
xnor U9736 (N_9736,N_9404,N_9298);
xor U9737 (N_9737,N_9469,N_9303);
nor U9738 (N_9738,N_9130,N_9017);
nor U9739 (N_9739,N_9216,N_9314);
and U9740 (N_9740,N_9255,N_9428);
nor U9741 (N_9741,N_9270,N_9238);
xor U9742 (N_9742,N_9011,N_9083);
xnor U9743 (N_9743,N_9446,N_9014);
and U9744 (N_9744,N_9411,N_9167);
xor U9745 (N_9745,N_9291,N_9219);
nor U9746 (N_9746,N_9065,N_9485);
or U9747 (N_9747,N_9478,N_9125);
or U9748 (N_9748,N_9231,N_9302);
nor U9749 (N_9749,N_9356,N_9150);
xor U9750 (N_9750,N_9215,N_9400);
xor U9751 (N_9751,N_9062,N_9227);
nor U9752 (N_9752,N_9383,N_9375);
and U9753 (N_9753,N_9486,N_9148);
and U9754 (N_9754,N_9097,N_9039);
nand U9755 (N_9755,N_9347,N_9255);
nand U9756 (N_9756,N_9006,N_9238);
nor U9757 (N_9757,N_9109,N_9014);
and U9758 (N_9758,N_9010,N_9127);
or U9759 (N_9759,N_9052,N_9014);
nand U9760 (N_9760,N_9122,N_9467);
nor U9761 (N_9761,N_9081,N_9498);
and U9762 (N_9762,N_9227,N_9403);
or U9763 (N_9763,N_9146,N_9316);
xor U9764 (N_9764,N_9148,N_9275);
xor U9765 (N_9765,N_9184,N_9014);
nand U9766 (N_9766,N_9101,N_9218);
or U9767 (N_9767,N_9437,N_9481);
and U9768 (N_9768,N_9310,N_9451);
or U9769 (N_9769,N_9373,N_9321);
nor U9770 (N_9770,N_9214,N_9008);
xor U9771 (N_9771,N_9297,N_9290);
nand U9772 (N_9772,N_9015,N_9023);
nand U9773 (N_9773,N_9094,N_9498);
xor U9774 (N_9774,N_9249,N_9377);
nor U9775 (N_9775,N_9268,N_9091);
or U9776 (N_9776,N_9042,N_9101);
and U9777 (N_9777,N_9057,N_9115);
nor U9778 (N_9778,N_9015,N_9255);
nor U9779 (N_9779,N_9284,N_9431);
and U9780 (N_9780,N_9026,N_9003);
or U9781 (N_9781,N_9446,N_9284);
nor U9782 (N_9782,N_9261,N_9465);
xor U9783 (N_9783,N_9191,N_9352);
or U9784 (N_9784,N_9460,N_9471);
xnor U9785 (N_9785,N_9479,N_9447);
xor U9786 (N_9786,N_9308,N_9286);
nor U9787 (N_9787,N_9044,N_9395);
and U9788 (N_9788,N_9230,N_9170);
nand U9789 (N_9789,N_9176,N_9093);
xor U9790 (N_9790,N_9387,N_9370);
nor U9791 (N_9791,N_9080,N_9338);
or U9792 (N_9792,N_9312,N_9380);
nor U9793 (N_9793,N_9332,N_9194);
xnor U9794 (N_9794,N_9353,N_9131);
xnor U9795 (N_9795,N_9162,N_9087);
and U9796 (N_9796,N_9092,N_9109);
and U9797 (N_9797,N_9156,N_9452);
and U9798 (N_9798,N_9255,N_9397);
xor U9799 (N_9799,N_9288,N_9201);
nand U9800 (N_9800,N_9051,N_9383);
nor U9801 (N_9801,N_9228,N_9230);
or U9802 (N_9802,N_9401,N_9114);
or U9803 (N_9803,N_9286,N_9377);
nor U9804 (N_9804,N_9252,N_9260);
nand U9805 (N_9805,N_9027,N_9452);
nor U9806 (N_9806,N_9498,N_9132);
xnor U9807 (N_9807,N_9311,N_9004);
or U9808 (N_9808,N_9123,N_9464);
and U9809 (N_9809,N_9277,N_9275);
xor U9810 (N_9810,N_9182,N_9162);
nand U9811 (N_9811,N_9414,N_9439);
and U9812 (N_9812,N_9197,N_9176);
nand U9813 (N_9813,N_9223,N_9026);
nand U9814 (N_9814,N_9424,N_9080);
xnor U9815 (N_9815,N_9243,N_9348);
or U9816 (N_9816,N_9253,N_9017);
nand U9817 (N_9817,N_9019,N_9051);
xor U9818 (N_9818,N_9026,N_9216);
and U9819 (N_9819,N_9328,N_9084);
nand U9820 (N_9820,N_9368,N_9229);
nor U9821 (N_9821,N_9473,N_9389);
xor U9822 (N_9822,N_9202,N_9183);
nand U9823 (N_9823,N_9410,N_9491);
xnor U9824 (N_9824,N_9044,N_9468);
nor U9825 (N_9825,N_9205,N_9024);
nand U9826 (N_9826,N_9479,N_9457);
xor U9827 (N_9827,N_9318,N_9274);
nand U9828 (N_9828,N_9442,N_9390);
xor U9829 (N_9829,N_9113,N_9323);
or U9830 (N_9830,N_9368,N_9012);
xnor U9831 (N_9831,N_9110,N_9270);
xor U9832 (N_9832,N_9078,N_9208);
nand U9833 (N_9833,N_9014,N_9471);
nor U9834 (N_9834,N_9021,N_9373);
nand U9835 (N_9835,N_9005,N_9418);
xor U9836 (N_9836,N_9031,N_9458);
xor U9837 (N_9837,N_9368,N_9456);
xor U9838 (N_9838,N_9333,N_9100);
or U9839 (N_9839,N_9169,N_9493);
or U9840 (N_9840,N_9023,N_9269);
or U9841 (N_9841,N_9366,N_9119);
nor U9842 (N_9842,N_9490,N_9347);
nor U9843 (N_9843,N_9337,N_9014);
and U9844 (N_9844,N_9122,N_9033);
xor U9845 (N_9845,N_9001,N_9246);
or U9846 (N_9846,N_9261,N_9444);
nor U9847 (N_9847,N_9171,N_9454);
and U9848 (N_9848,N_9138,N_9419);
or U9849 (N_9849,N_9205,N_9207);
nand U9850 (N_9850,N_9420,N_9317);
or U9851 (N_9851,N_9124,N_9272);
nand U9852 (N_9852,N_9004,N_9050);
nand U9853 (N_9853,N_9485,N_9272);
nand U9854 (N_9854,N_9182,N_9314);
nand U9855 (N_9855,N_9472,N_9017);
or U9856 (N_9856,N_9053,N_9257);
and U9857 (N_9857,N_9069,N_9013);
nor U9858 (N_9858,N_9027,N_9129);
nand U9859 (N_9859,N_9078,N_9298);
and U9860 (N_9860,N_9070,N_9155);
and U9861 (N_9861,N_9138,N_9184);
nor U9862 (N_9862,N_9343,N_9084);
nand U9863 (N_9863,N_9295,N_9080);
xor U9864 (N_9864,N_9335,N_9337);
and U9865 (N_9865,N_9481,N_9403);
nand U9866 (N_9866,N_9145,N_9217);
and U9867 (N_9867,N_9477,N_9154);
nand U9868 (N_9868,N_9169,N_9154);
xnor U9869 (N_9869,N_9498,N_9044);
nor U9870 (N_9870,N_9368,N_9133);
nand U9871 (N_9871,N_9345,N_9198);
nor U9872 (N_9872,N_9304,N_9435);
nor U9873 (N_9873,N_9105,N_9421);
xnor U9874 (N_9874,N_9000,N_9331);
nand U9875 (N_9875,N_9341,N_9475);
and U9876 (N_9876,N_9020,N_9442);
and U9877 (N_9877,N_9259,N_9459);
nand U9878 (N_9878,N_9479,N_9491);
nor U9879 (N_9879,N_9322,N_9378);
or U9880 (N_9880,N_9146,N_9244);
nand U9881 (N_9881,N_9111,N_9132);
or U9882 (N_9882,N_9067,N_9402);
or U9883 (N_9883,N_9497,N_9430);
or U9884 (N_9884,N_9276,N_9012);
or U9885 (N_9885,N_9070,N_9463);
xnor U9886 (N_9886,N_9370,N_9105);
or U9887 (N_9887,N_9312,N_9319);
xnor U9888 (N_9888,N_9202,N_9316);
and U9889 (N_9889,N_9484,N_9141);
nand U9890 (N_9890,N_9278,N_9144);
and U9891 (N_9891,N_9211,N_9287);
nand U9892 (N_9892,N_9147,N_9334);
nand U9893 (N_9893,N_9354,N_9489);
or U9894 (N_9894,N_9105,N_9195);
nor U9895 (N_9895,N_9478,N_9466);
xor U9896 (N_9896,N_9302,N_9327);
xor U9897 (N_9897,N_9042,N_9360);
and U9898 (N_9898,N_9108,N_9116);
nor U9899 (N_9899,N_9458,N_9250);
or U9900 (N_9900,N_9216,N_9485);
and U9901 (N_9901,N_9115,N_9487);
and U9902 (N_9902,N_9211,N_9436);
or U9903 (N_9903,N_9400,N_9333);
xor U9904 (N_9904,N_9026,N_9491);
nand U9905 (N_9905,N_9287,N_9283);
and U9906 (N_9906,N_9020,N_9411);
nand U9907 (N_9907,N_9153,N_9148);
xor U9908 (N_9908,N_9142,N_9180);
nand U9909 (N_9909,N_9446,N_9199);
and U9910 (N_9910,N_9177,N_9038);
nor U9911 (N_9911,N_9426,N_9205);
xnor U9912 (N_9912,N_9008,N_9225);
xnor U9913 (N_9913,N_9234,N_9483);
or U9914 (N_9914,N_9273,N_9016);
nand U9915 (N_9915,N_9108,N_9259);
nand U9916 (N_9916,N_9047,N_9089);
nor U9917 (N_9917,N_9225,N_9073);
nor U9918 (N_9918,N_9132,N_9321);
xor U9919 (N_9919,N_9458,N_9290);
and U9920 (N_9920,N_9483,N_9343);
xnor U9921 (N_9921,N_9360,N_9037);
nand U9922 (N_9922,N_9089,N_9434);
xnor U9923 (N_9923,N_9186,N_9302);
nand U9924 (N_9924,N_9452,N_9064);
or U9925 (N_9925,N_9009,N_9268);
nor U9926 (N_9926,N_9286,N_9125);
xor U9927 (N_9927,N_9439,N_9271);
or U9928 (N_9928,N_9485,N_9089);
nor U9929 (N_9929,N_9329,N_9001);
or U9930 (N_9930,N_9409,N_9193);
nand U9931 (N_9931,N_9007,N_9264);
nand U9932 (N_9932,N_9169,N_9415);
xor U9933 (N_9933,N_9482,N_9364);
or U9934 (N_9934,N_9468,N_9396);
xnor U9935 (N_9935,N_9073,N_9474);
nor U9936 (N_9936,N_9148,N_9304);
or U9937 (N_9937,N_9149,N_9071);
and U9938 (N_9938,N_9330,N_9484);
xnor U9939 (N_9939,N_9403,N_9262);
or U9940 (N_9940,N_9468,N_9470);
or U9941 (N_9941,N_9151,N_9257);
xnor U9942 (N_9942,N_9188,N_9272);
nand U9943 (N_9943,N_9317,N_9233);
and U9944 (N_9944,N_9024,N_9011);
nand U9945 (N_9945,N_9102,N_9052);
or U9946 (N_9946,N_9329,N_9238);
and U9947 (N_9947,N_9118,N_9141);
or U9948 (N_9948,N_9307,N_9109);
xor U9949 (N_9949,N_9287,N_9251);
nor U9950 (N_9950,N_9063,N_9240);
or U9951 (N_9951,N_9169,N_9189);
nor U9952 (N_9952,N_9165,N_9239);
or U9953 (N_9953,N_9165,N_9245);
nor U9954 (N_9954,N_9058,N_9017);
nor U9955 (N_9955,N_9489,N_9471);
nor U9956 (N_9956,N_9210,N_9037);
nor U9957 (N_9957,N_9086,N_9043);
nand U9958 (N_9958,N_9100,N_9345);
and U9959 (N_9959,N_9252,N_9346);
xor U9960 (N_9960,N_9178,N_9234);
or U9961 (N_9961,N_9438,N_9050);
nor U9962 (N_9962,N_9442,N_9100);
xnor U9963 (N_9963,N_9121,N_9391);
xor U9964 (N_9964,N_9045,N_9046);
nor U9965 (N_9965,N_9000,N_9458);
xnor U9966 (N_9966,N_9240,N_9445);
nand U9967 (N_9967,N_9337,N_9226);
or U9968 (N_9968,N_9417,N_9159);
or U9969 (N_9969,N_9334,N_9183);
and U9970 (N_9970,N_9125,N_9179);
nand U9971 (N_9971,N_9440,N_9181);
xnor U9972 (N_9972,N_9192,N_9058);
nor U9973 (N_9973,N_9262,N_9309);
xnor U9974 (N_9974,N_9014,N_9130);
and U9975 (N_9975,N_9466,N_9277);
xor U9976 (N_9976,N_9171,N_9263);
nand U9977 (N_9977,N_9460,N_9370);
and U9978 (N_9978,N_9201,N_9165);
nand U9979 (N_9979,N_9433,N_9027);
xor U9980 (N_9980,N_9294,N_9339);
and U9981 (N_9981,N_9273,N_9066);
nand U9982 (N_9982,N_9329,N_9278);
nor U9983 (N_9983,N_9344,N_9243);
and U9984 (N_9984,N_9301,N_9148);
nor U9985 (N_9985,N_9380,N_9175);
nor U9986 (N_9986,N_9113,N_9481);
or U9987 (N_9987,N_9391,N_9151);
xor U9988 (N_9988,N_9141,N_9100);
xor U9989 (N_9989,N_9012,N_9334);
or U9990 (N_9990,N_9351,N_9302);
xnor U9991 (N_9991,N_9310,N_9265);
xnor U9992 (N_9992,N_9234,N_9264);
xor U9993 (N_9993,N_9334,N_9173);
xnor U9994 (N_9994,N_9371,N_9112);
nor U9995 (N_9995,N_9435,N_9270);
nand U9996 (N_9996,N_9029,N_9475);
nor U9997 (N_9997,N_9057,N_9465);
nor U9998 (N_9998,N_9114,N_9317);
nor U9999 (N_9999,N_9218,N_9425);
nand U10000 (N_10000,N_9964,N_9752);
or U10001 (N_10001,N_9785,N_9853);
xor U10002 (N_10002,N_9616,N_9695);
or U10003 (N_10003,N_9520,N_9645);
and U10004 (N_10004,N_9801,N_9915);
or U10005 (N_10005,N_9704,N_9787);
nand U10006 (N_10006,N_9910,N_9939);
and U10007 (N_10007,N_9795,N_9943);
nor U10008 (N_10008,N_9686,N_9771);
or U10009 (N_10009,N_9602,N_9879);
and U10010 (N_10010,N_9619,N_9625);
and U10011 (N_10011,N_9657,N_9623);
or U10012 (N_10012,N_9767,N_9663);
xor U10013 (N_10013,N_9539,N_9710);
and U10014 (N_10014,N_9703,N_9847);
and U10015 (N_10015,N_9630,N_9569);
xor U10016 (N_10016,N_9983,N_9803);
and U10017 (N_10017,N_9747,N_9749);
or U10018 (N_10018,N_9639,N_9541);
nor U10019 (N_10019,N_9917,N_9502);
xnor U10020 (N_10020,N_9932,N_9624);
xnor U10021 (N_10021,N_9978,N_9885);
or U10022 (N_10022,N_9789,N_9620);
and U10023 (N_10023,N_9726,N_9953);
nor U10024 (N_10024,N_9537,N_9603);
xor U10025 (N_10025,N_9936,N_9841);
and U10026 (N_10026,N_9924,N_9600);
and U10027 (N_10027,N_9890,N_9865);
nand U10028 (N_10028,N_9552,N_9986);
nor U10029 (N_10029,N_9941,N_9974);
nand U10030 (N_10030,N_9618,N_9842);
or U10031 (N_10031,N_9768,N_9857);
xnor U10032 (N_10032,N_9884,N_9582);
xnor U10033 (N_10033,N_9678,N_9891);
xor U10034 (N_10034,N_9558,N_9652);
nor U10035 (N_10035,N_9594,N_9866);
nand U10036 (N_10036,N_9700,N_9685);
nand U10037 (N_10037,N_9731,N_9806);
or U10038 (N_10038,N_9674,N_9680);
nand U10039 (N_10039,N_9590,N_9863);
or U10040 (N_10040,N_9732,N_9957);
nor U10041 (N_10041,N_9778,N_9599);
nor U10042 (N_10042,N_9506,N_9770);
or U10043 (N_10043,N_9959,N_9548);
xnor U10044 (N_10044,N_9893,N_9969);
or U10045 (N_10045,N_9561,N_9693);
nand U10046 (N_10046,N_9780,N_9500);
or U10047 (N_10047,N_9887,N_9870);
nor U10048 (N_10048,N_9567,N_9533);
xor U10049 (N_10049,N_9738,N_9777);
xnor U10050 (N_10050,N_9553,N_9912);
nand U10051 (N_10051,N_9702,N_9937);
nor U10052 (N_10052,N_9748,N_9916);
or U10053 (N_10053,N_9889,N_9819);
or U10054 (N_10054,N_9952,N_9570);
or U10055 (N_10055,N_9595,N_9968);
and U10056 (N_10056,N_9990,N_9642);
and U10057 (N_10057,N_9508,N_9888);
xor U10058 (N_10058,N_9689,N_9880);
nor U10059 (N_10059,N_9825,N_9766);
xnor U10060 (N_10060,N_9810,N_9804);
nand U10061 (N_10061,N_9566,N_9858);
or U10062 (N_10062,N_9903,N_9907);
or U10063 (N_10063,N_9719,N_9756);
and U10064 (N_10064,N_9737,N_9579);
nand U10065 (N_10065,N_9995,N_9942);
nor U10066 (N_10066,N_9871,N_9572);
nor U10067 (N_10067,N_9892,N_9975);
or U10068 (N_10068,N_9784,N_9683);
or U10069 (N_10069,N_9805,N_9744);
nor U10070 (N_10070,N_9633,N_9587);
nor U10071 (N_10071,N_9922,N_9631);
or U10072 (N_10072,N_9928,N_9746);
xnor U10073 (N_10073,N_9614,N_9517);
or U10074 (N_10074,N_9989,N_9850);
xnor U10075 (N_10075,N_9714,N_9741);
and U10076 (N_10076,N_9809,N_9628);
nand U10077 (N_10077,N_9965,N_9906);
and U10078 (N_10078,N_9963,N_9796);
or U10079 (N_10079,N_9905,N_9988);
xnor U10080 (N_10080,N_9755,N_9724);
or U10081 (N_10081,N_9585,N_9708);
nand U10082 (N_10082,N_9834,N_9949);
and U10083 (N_10083,N_9504,N_9881);
nor U10084 (N_10084,N_9882,N_9859);
and U10085 (N_10085,N_9711,N_9627);
nor U10086 (N_10086,N_9532,N_9934);
nor U10087 (N_10087,N_9929,N_9687);
xor U10088 (N_10088,N_9876,N_9641);
nand U10089 (N_10089,N_9926,N_9800);
nor U10090 (N_10090,N_9586,N_9705);
and U10091 (N_10091,N_9947,N_9516);
or U10092 (N_10092,N_9560,N_9985);
nor U10093 (N_10093,N_9846,N_9608);
nor U10094 (N_10094,N_9546,N_9886);
nand U10095 (N_10095,N_9933,N_9513);
and U10096 (N_10096,N_9675,N_9528);
and U10097 (N_10097,N_9763,N_9643);
or U10098 (N_10098,N_9644,N_9543);
and U10099 (N_10099,N_9946,N_9831);
or U10100 (N_10100,N_9820,N_9909);
nand U10101 (N_10101,N_9691,N_9571);
nand U10102 (N_10102,N_9525,N_9613);
nor U10103 (N_10103,N_9725,N_9505);
nand U10104 (N_10104,N_9733,N_9824);
nand U10105 (N_10105,N_9984,N_9815);
or U10106 (N_10106,N_9832,N_9813);
and U10107 (N_10107,N_9735,N_9765);
or U10108 (N_10108,N_9655,N_9617);
nor U10109 (N_10109,N_9651,N_9901);
or U10110 (N_10110,N_9722,N_9837);
xor U10111 (N_10111,N_9707,N_9666);
nor U10112 (N_10112,N_9826,N_9745);
nand U10113 (N_10113,N_9510,N_9697);
or U10114 (N_10114,N_9874,N_9734);
xor U10115 (N_10115,N_9632,N_9716);
and U10116 (N_10116,N_9640,N_9764);
xnor U10117 (N_10117,N_9998,N_9592);
or U10118 (N_10118,N_9896,N_9883);
xnor U10119 (N_10119,N_9701,N_9754);
xnor U10120 (N_10120,N_9951,N_9781);
or U10121 (N_10121,N_9682,N_9667);
xnor U10122 (N_10122,N_9769,N_9607);
nand U10123 (N_10123,N_9650,N_9718);
nand U10124 (N_10124,N_9565,N_9563);
and U10125 (N_10125,N_9753,N_9501);
and U10126 (N_10126,N_9669,N_9549);
and U10127 (N_10127,N_9576,N_9958);
nor U10128 (N_10128,N_9811,N_9739);
nand U10129 (N_10129,N_9862,N_9908);
or U10130 (N_10130,N_9783,N_9659);
nand U10131 (N_10131,N_9527,N_9554);
nand U10132 (N_10132,N_9730,N_9798);
and U10133 (N_10133,N_9830,N_9559);
and U10134 (N_10134,N_9994,N_9698);
or U10135 (N_10135,N_9791,N_9914);
xnor U10136 (N_10136,N_9930,N_9720);
or U10137 (N_10137,N_9817,N_9868);
nor U10138 (N_10138,N_9997,N_9772);
nor U10139 (N_10139,N_9851,N_9526);
and U10140 (N_10140,N_9668,N_9977);
and U10141 (N_10141,N_9751,N_9971);
xnor U10142 (N_10142,N_9966,N_9931);
or U10143 (N_10143,N_9814,N_9944);
or U10144 (N_10144,N_9935,N_9979);
and U10145 (N_10145,N_9962,N_9911);
and U10146 (N_10146,N_9653,N_9564);
or U10147 (N_10147,N_9597,N_9544);
nand U10148 (N_10148,N_9635,N_9514);
xor U10149 (N_10149,N_9521,N_9773);
or U10150 (N_10150,N_9845,N_9855);
nand U10151 (N_10151,N_9503,N_9799);
or U10152 (N_10152,N_9774,N_9793);
and U10153 (N_10153,N_9878,N_9981);
xnor U10154 (N_10154,N_9950,N_9583);
and U10155 (N_10155,N_9728,N_9670);
xor U10156 (N_10156,N_9869,N_9665);
xnor U10157 (N_10157,N_9828,N_9588);
or U10158 (N_10158,N_9736,N_9536);
nand U10159 (N_10159,N_9991,N_9818);
or U10160 (N_10160,N_9976,N_9925);
xor U10161 (N_10161,N_9993,N_9894);
xor U10162 (N_10162,N_9601,N_9822);
xnor U10163 (N_10163,N_9530,N_9581);
or U10164 (N_10164,N_9522,N_9696);
xor U10165 (N_10165,N_9664,N_9758);
or U10166 (N_10166,N_9584,N_9551);
and U10167 (N_10167,N_9895,N_9821);
nor U10168 (N_10168,N_9872,N_9775);
or U10169 (N_10169,N_9550,N_9762);
and U10170 (N_10170,N_9512,N_9534);
or U10171 (N_10171,N_9694,N_9577);
and U10172 (N_10172,N_9555,N_9538);
xnor U10173 (N_10173,N_9761,N_9699);
xor U10174 (N_10174,N_9591,N_9898);
and U10175 (N_10175,N_9759,N_9626);
or U10176 (N_10176,N_9829,N_9750);
nor U10177 (N_10177,N_9604,N_9634);
and U10178 (N_10178,N_9786,N_9838);
and U10179 (N_10179,N_9709,N_9684);
xor U10180 (N_10180,N_9545,N_9511);
xnor U10181 (N_10181,N_9899,N_9518);
and U10182 (N_10182,N_9960,N_9970);
and U10183 (N_10183,N_9556,N_9854);
or U10184 (N_10184,N_9575,N_9927);
nor U10185 (N_10185,N_9992,N_9676);
xor U10186 (N_10186,N_9794,N_9861);
and U10187 (N_10187,N_9557,N_9921);
nand U10188 (N_10188,N_9788,N_9948);
nand U10189 (N_10189,N_9835,N_9562);
nor U10190 (N_10190,N_9515,N_9679);
nand U10191 (N_10191,N_9833,N_9982);
nand U10192 (N_10192,N_9742,N_9816);
or U10193 (N_10193,N_9622,N_9776);
and U10194 (N_10194,N_9823,N_9972);
and U10195 (N_10195,N_9647,N_9523);
nor U10196 (N_10196,N_9540,N_9802);
nor U10197 (N_10197,N_9839,N_9904);
nor U10198 (N_10198,N_9743,N_9568);
nor U10199 (N_10199,N_9656,N_9938);
xor U10200 (N_10200,N_9797,N_9973);
xor U10201 (N_10201,N_9860,N_9790);
or U10202 (N_10202,N_9596,N_9638);
and U10203 (N_10203,N_9649,N_9864);
xor U10204 (N_10204,N_9715,N_9808);
nand U10205 (N_10205,N_9648,N_9849);
nor U10206 (N_10206,N_9509,N_9856);
nor U10207 (N_10207,N_9945,N_9706);
or U10208 (N_10208,N_9612,N_9661);
nor U10209 (N_10209,N_9573,N_9672);
nor U10210 (N_10210,N_9782,N_9923);
xor U10211 (N_10211,N_9918,N_9987);
nor U10212 (N_10212,N_9692,N_9877);
nand U10213 (N_10213,N_9920,N_9843);
or U10214 (N_10214,N_9615,N_9673);
and U10215 (N_10215,N_9717,N_9507);
nor U10216 (N_10216,N_9723,N_9690);
nand U10217 (N_10217,N_9519,N_9848);
and U10218 (N_10218,N_9812,N_9713);
or U10219 (N_10219,N_9955,N_9897);
and U10220 (N_10220,N_9902,N_9807);
and U10221 (N_10221,N_9688,N_9636);
and U10222 (N_10222,N_9792,N_9681);
and U10223 (N_10223,N_9873,N_9721);
xor U10224 (N_10224,N_9660,N_9956);
xor U10225 (N_10225,N_9840,N_9760);
xor U10226 (N_10226,N_9605,N_9578);
and U10227 (N_10227,N_9646,N_9740);
nor U10228 (N_10228,N_9867,N_9658);
xnor U10229 (N_10229,N_9712,N_9727);
nor U10230 (N_10230,N_9779,N_9629);
nand U10231 (N_10231,N_9580,N_9827);
and U10232 (N_10232,N_9940,N_9729);
and U10233 (N_10233,N_9980,N_9852);
and U10234 (N_10234,N_9875,N_9542);
nor U10235 (N_10235,N_9913,N_9637);
xnor U10236 (N_10236,N_9606,N_9677);
xor U10237 (N_10237,N_9593,N_9999);
xor U10238 (N_10238,N_9535,N_9919);
or U10239 (N_10239,N_9757,N_9967);
or U10240 (N_10240,N_9671,N_9961);
and U10241 (N_10241,N_9996,N_9621);
nand U10242 (N_10242,N_9547,N_9610);
nor U10243 (N_10243,N_9589,N_9529);
and U10244 (N_10244,N_9654,N_9836);
and U10245 (N_10245,N_9609,N_9844);
or U10246 (N_10246,N_9954,N_9598);
and U10247 (N_10247,N_9574,N_9524);
and U10248 (N_10248,N_9662,N_9611);
and U10249 (N_10249,N_9531,N_9900);
xnor U10250 (N_10250,N_9954,N_9742);
or U10251 (N_10251,N_9583,N_9903);
nor U10252 (N_10252,N_9734,N_9650);
nand U10253 (N_10253,N_9525,N_9524);
nand U10254 (N_10254,N_9503,N_9918);
xor U10255 (N_10255,N_9537,N_9885);
and U10256 (N_10256,N_9856,N_9569);
xor U10257 (N_10257,N_9859,N_9653);
and U10258 (N_10258,N_9832,N_9984);
nand U10259 (N_10259,N_9601,N_9977);
nand U10260 (N_10260,N_9952,N_9547);
nor U10261 (N_10261,N_9765,N_9798);
xnor U10262 (N_10262,N_9861,N_9601);
nor U10263 (N_10263,N_9550,N_9617);
xor U10264 (N_10264,N_9850,N_9660);
nand U10265 (N_10265,N_9587,N_9825);
and U10266 (N_10266,N_9866,N_9742);
xnor U10267 (N_10267,N_9879,N_9562);
nand U10268 (N_10268,N_9861,N_9910);
or U10269 (N_10269,N_9566,N_9876);
and U10270 (N_10270,N_9845,N_9545);
and U10271 (N_10271,N_9991,N_9591);
nor U10272 (N_10272,N_9974,N_9641);
nand U10273 (N_10273,N_9853,N_9721);
nand U10274 (N_10274,N_9550,N_9952);
nand U10275 (N_10275,N_9626,N_9550);
nand U10276 (N_10276,N_9740,N_9803);
nor U10277 (N_10277,N_9706,N_9652);
xnor U10278 (N_10278,N_9783,N_9832);
xor U10279 (N_10279,N_9955,N_9928);
nand U10280 (N_10280,N_9651,N_9520);
xor U10281 (N_10281,N_9603,N_9809);
nand U10282 (N_10282,N_9739,N_9664);
nand U10283 (N_10283,N_9735,N_9734);
and U10284 (N_10284,N_9702,N_9841);
and U10285 (N_10285,N_9953,N_9903);
xnor U10286 (N_10286,N_9507,N_9723);
or U10287 (N_10287,N_9525,N_9586);
or U10288 (N_10288,N_9612,N_9937);
xor U10289 (N_10289,N_9802,N_9662);
and U10290 (N_10290,N_9948,N_9763);
nor U10291 (N_10291,N_9745,N_9564);
xnor U10292 (N_10292,N_9541,N_9957);
or U10293 (N_10293,N_9892,N_9748);
nand U10294 (N_10294,N_9634,N_9515);
nand U10295 (N_10295,N_9986,N_9663);
and U10296 (N_10296,N_9587,N_9907);
xnor U10297 (N_10297,N_9861,N_9597);
or U10298 (N_10298,N_9691,N_9923);
and U10299 (N_10299,N_9759,N_9737);
xor U10300 (N_10300,N_9664,N_9977);
nand U10301 (N_10301,N_9559,N_9892);
nand U10302 (N_10302,N_9676,N_9701);
nor U10303 (N_10303,N_9825,N_9943);
nand U10304 (N_10304,N_9555,N_9780);
and U10305 (N_10305,N_9568,N_9590);
and U10306 (N_10306,N_9815,N_9657);
and U10307 (N_10307,N_9843,N_9817);
xnor U10308 (N_10308,N_9638,N_9517);
nand U10309 (N_10309,N_9660,N_9634);
and U10310 (N_10310,N_9911,N_9959);
and U10311 (N_10311,N_9825,N_9707);
and U10312 (N_10312,N_9863,N_9793);
nand U10313 (N_10313,N_9565,N_9512);
xnor U10314 (N_10314,N_9589,N_9944);
and U10315 (N_10315,N_9731,N_9598);
nand U10316 (N_10316,N_9638,N_9717);
nor U10317 (N_10317,N_9659,N_9883);
and U10318 (N_10318,N_9575,N_9710);
xnor U10319 (N_10319,N_9884,N_9896);
and U10320 (N_10320,N_9946,N_9641);
xnor U10321 (N_10321,N_9563,N_9808);
nand U10322 (N_10322,N_9562,N_9857);
nand U10323 (N_10323,N_9777,N_9617);
nor U10324 (N_10324,N_9560,N_9895);
and U10325 (N_10325,N_9821,N_9777);
xnor U10326 (N_10326,N_9550,N_9669);
nor U10327 (N_10327,N_9911,N_9884);
and U10328 (N_10328,N_9565,N_9935);
nand U10329 (N_10329,N_9710,N_9754);
xor U10330 (N_10330,N_9576,N_9660);
nand U10331 (N_10331,N_9517,N_9502);
xnor U10332 (N_10332,N_9936,N_9805);
or U10333 (N_10333,N_9594,N_9724);
nor U10334 (N_10334,N_9549,N_9667);
or U10335 (N_10335,N_9936,N_9788);
nor U10336 (N_10336,N_9863,N_9677);
nand U10337 (N_10337,N_9696,N_9999);
or U10338 (N_10338,N_9753,N_9648);
xor U10339 (N_10339,N_9664,N_9874);
nor U10340 (N_10340,N_9906,N_9753);
nor U10341 (N_10341,N_9988,N_9907);
nand U10342 (N_10342,N_9934,N_9770);
nor U10343 (N_10343,N_9974,N_9797);
nor U10344 (N_10344,N_9566,N_9739);
xor U10345 (N_10345,N_9875,N_9609);
nor U10346 (N_10346,N_9736,N_9624);
nor U10347 (N_10347,N_9776,N_9568);
nand U10348 (N_10348,N_9857,N_9629);
and U10349 (N_10349,N_9920,N_9611);
and U10350 (N_10350,N_9591,N_9685);
nor U10351 (N_10351,N_9726,N_9617);
nand U10352 (N_10352,N_9687,N_9954);
nand U10353 (N_10353,N_9906,N_9548);
or U10354 (N_10354,N_9708,N_9863);
nand U10355 (N_10355,N_9903,N_9566);
nor U10356 (N_10356,N_9821,N_9633);
or U10357 (N_10357,N_9993,N_9576);
nand U10358 (N_10358,N_9709,N_9918);
or U10359 (N_10359,N_9935,N_9593);
nor U10360 (N_10360,N_9897,N_9608);
or U10361 (N_10361,N_9744,N_9860);
nor U10362 (N_10362,N_9962,N_9720);
nand U10363 (N_10363,N_9759,N_9971);
and U10364 (N_10364,N_9752,N_9597);
or U10365 (N_10365,N_9722,N_9815);
nand U10366 (N_10366,N_9634,N_9629);
nor U10367 (N_10367,N_9872,N_9871);
nand U10368 (N_10368,N_9618,N_9926);
nor U10369 (N_10369,N_9949,N_9734);
or U10370 (N_10370,N_9751,N_9543);
and U10371 (N_10371,N_9605,N_9833);
or U10372 (N_10372,N_9870,N_9512);
nand U10373 (N_10373,N_9673,N_9665);
and U10374 (N_10374,N_9902,N_9756);
or U10375 (N_10375,N_9724,N_9870);
and U10376 (N_10376,N_9923,N_9767);
xor U10377 (N_10377,N_9778,N_9817);
nor U10378 (N_10378,N_9988,N_9948);
nor U10379 (N_10379,N_9945,N_9715);
nor U10380 (N_10380,N_9891,N_9974);
xor U10381 (N_10381,N_9693,N_9868);
and U10382 (N_10382,N_9979,N_9896);
xor U10383 (N_10383,N_9558,N_9560);
xnor U10384 (N_10384,N_9897,N_9547);
and U10385 (N_10385,N_9817,N_9892);
xor U10386 (N_10386,N_9616,N_9870);
nor U10387 (N_10387,N_9916,N_9654);
nand U10388 (N_10388,N_9561,N_9980);
nor U10389 (N_10389,N_9791,N_9906);
nor U10390 (N_10390,N_9613,N_9787);
nor U10391 (N_10391,N_9792,N_9888);
and U10392 (N_10392,N_9751,N_9705);
and U10393 (N_10393,N_9517,N_9578);
or U10394 (N_10394,N_9623,N_9603);
nor U10395 (N_10395,N_9742,N_9695);
nor U10396 (N_10396,N_9704,N_9717);
nand U10397 (N_10397,N_9826,N_9649);
nor U10398 (N_10398,N_9935,N_9913);
or U10399 (N_10399,N_9840,N_9775);
or U10400 (N_10400,N_9728,N_9845);
nor U10401 (N_10401,N_9959,N_9963);
nand U10402 (N_10402,N_9980,N_9986);
nand U10403 (N_10403,N_9625,N_9924);
nand U10404 (N_10404,N_9845,N_9839);
xnor U10405 (N_10405,N_9719,N_9517);
nor U10406 (N_10406,N_9787,N_9660);
nor U10407 (N_10407,N_9966,N_9929);
xor U10408 (N_10408,N_9939,N_9842);
and U10409 (N_10409,N_9806,N_9923);
xor U10410 (N_10410,N_9867,N_9936);
xor U10411 (N_10411,N_9610,N_9539);
nor U10412 (N_10412,N_9552,N_9575);
xnor U10413 (N_10413,N_9564,N_9884);
and U10414 (N_10414,N_9625,N_9862);
nand U10415 (N_10415,N_9564,N_9587);
nand U10416 (N_10416,N_9862,N_9851);
xnor U10417 (N_10417,N_9725,N_9747);
nor U10418 (N_10418,N_9593,N_9756);
nand U10419 (N_10419,N_9636,N_9694);
nor U10420 (N_10420,N_9919,N_9733);
and U10421 (N_10421,N_9554,N_9862);
and U10422 (N_10422,N_9736,N_9854);
nor U10423 (N_10423,N_9926,N_9685);
xor U10424 (N_10424,N_9665,N_9625);
or U10425 (N_10425,N_9945,N_9828);
nor U10426 (N_10426,N_9929,N_9570);
and U10427 (N_10427,N_9960,N_9907);
nand U10428 (N_10428,N_9976,N_9952);
nand U10429 (N_10429,N_9546,N_9872);
and U10430 (N_10430,N_9833,N_9500);
xnor U10431 (N_10431,N_9783,N_9566);
and U10432 (N_10432,N_9618,N_9651);
or U10433 (N_10433,N_9850,N_9778);
nor U10434 (N_10434,N_9741,N_9529);
or U10435 (N_10435,N_9991,N_9689);
or U10436 (N_10436,N_9658,N_9546);
and U10437 (N_10437,N_9553,N_9775);
and U10438 (N_10438,N_9565,N_9662);
or U10439 (N_10439,N_9667,N_9848);
nand U10440 (N_10440,N_9632,N_9807);
nand U10441 (N_10441,N_9936,N_9861);
nor U10442 (N_10442,N_9631,N_9714);
and U10443 (N_10443,N_9780,N_9898);
nand U10444 (N_10444,N_9891,N_9551);
xor U10445 (N_10445,N_9983,N_9511);
and U10446 (N_10446,N_9520,N_9825);
nand U10447 (N_10447,N_9570,N_9648);
and U10448 (N_10448,N_9928,N_9553);
nand U10449 (N_10449,N_9912,N_9649);
nor U10450 (N_10450,N_9815,N_9616);
or U10451 (N_10451,N_9945,N_9760);
and U10452 (N_10452,N_9652,N_9768);
or U10453 (N_10453,N_9659,N_9542);
nand U10454 (N_10454,N_9597,N_9872);
xor U10455 (N_10455,N_9740,N_9548);
nand U10456 (N_10456,N_9827,N_9600);
or U10457 (N_10457,N_9876,N_9801);
and U10458 (N_10458,N_9885,N_9681);
or U10459 (N_10459,N_9672,N_9635);
or U10460 (N_10460,N_9639,N_9928);
and U10461 (N_10461,N_9700,N_9869);
xor U10462 (N_10462,N_9784,N_9633);
xor U10463 (N_10463,N_9783,N_9945);
xnor U10464 (N_10464,N_9916,N_9709);
xnor U10465 (N_10465,N_9714,N_9547);
or U10466 (N_10466,N_9722,N_9655);
and U10467 (N_10467,N_9555,N_9659);
xnor U10468 (N_10468,N_9834,N_9587);
xnor U10469 (N_10469,N_9934,N_9812);
nand U10470 (N_10470,N_9932,N_9621);
nand U10471 (N_10471,N_9878,N_9859);
xor U10472 (N_10472,N_9821,N_9929);
or U10473 (N_10473,N_9661,N_9943);
xnor U10474 (N_10474,N_9810,N_9991);
or U10475 (N_10475,N_9596,N_9606);
or U10476 (N_10476,N_9750,N_9634);
or U10477 (N_10477,N_9800,N_9832);
nor U10478 (N_10478,N_9601,N_9913);
nor U10479 (N_10479,N_9998,N_9553);
nand U10480 (N_10480,N_9607,N_9647);
nor U10481 (N_10481,N_9691,N_9837);
nand U10482 (N_10482,N_9974,N_9630);
nand U10483 (N_10483,N_9523,N_9760);
nand U10484 (N_10484,N_9759,N_9830);
nand U10485 (N_10485,N_9637,N_9964);
nor U10486 (N_10486,N_9520,N_9562);
nor U10487 (N_10487,N_9611,N_9656);
and U10488 (N_10488,N_9652,N_9783);
and U10489 (N_10489,N_9513,N_9664);
xnor U10490 (N_10490,N_9718,N_9706);
nor U10491 (N_10491,N_9916,N_9754);
and U10492 (N_10492,N_9505,N_9826);
nor U10493 (N_10493,N_9926,N_9601);
xor U10494 (N_10494,N_9794,N_9937);
or U10495 (N_10495,N_9900,N_9983);
or U10496 (N_10496,N_9896,N_9504);
and U10497 (N_10497,N_9990,N_9783);
or U10498 (N_10498,N_9576,N_9520);
xor U10499 (N_10499,N_9885,N_9584);
nand U10500 (N_10500,N_10416,N_10111);
nand U10501 (N_10501,N_10085,N_10353);
or U10502 (N_10502,N_10094,N_10272);
nand U10503 (N_10503,N_10122,N_10341);
xor U10504 (N_10504,N_10171,N_10036);
xor U10505 (N_10505,N_10069,N_10449);
or U10506 (N_10506,N_10189,N_10246);
nor U10507 (N_10507,N_10237,N_10390);
nor U10508 (N_10508,N_10498,N_10467);
nand U10509 (N_10509,N_10109,N_10385);
xor U10510 (N_10510,N_10399,N_10215);
nor U10511 (N_10511,N_10082,N_10490);
nor U10512 (N_10512,N_10361,N_10130);
or U10513 (N_10513,N_10305,N_10414);
nor U10514 (N_10514,N_10410,N_10205);
nor U10515 (N_10515,N_10167,N_10168);
nand U10516 (N_10516,N_10123,N_10116);
xor U10517 (N_10517,N_10285,N_10125);
and U10518 (N_10518,N_10183,N_10201);
nand U10519 (N_10519,N_10006,N_10476);
xor U10520 (N_10520,N_10232,N_10281);
or U10521 (N_10521,N_10436,N_10386);
nand U10522 (N_10522,N_10198,N_10277);
or U10523 (N_10523,N_10179,N_10045);
and U10524 (N_10524,N_10087,N_10202);
xor U10525 (N_10525,N_10051,N_10014);
xor U10526 (N_10526,N_10273,N_10304);
xor U10527 (N_10527,N_10342,N_10288);
nand U10528 (N_10528,N_10029,N_10250);
nor U10529 (N_10529,N_10450,N_10474);
and U10530 (N_10530,N_10265,N_10119);
or U10531 (N_10531,N_10354,N_10058);
nor U10532 (N_10532,N_10487,N_10221);
nor U10533 (N_10533,N_10294,N_10121);
xnor U10534 (N_10534,N_10317,N_10157);
or U10535 (N_10535,N_10211,N_10040);
xor U10536 (N_10536,N_10351,N_10411);
nor U10537 (N_10537,N_10268,N_10015);
xnor U10538 (N_10538,N_10401,N_10113);
and U10539 (N_10539,N_10453,N_10327);
and U10540 (N_10540,N_10472,N_10076);
nor U10541 (N_10541,N_10177,N_10251);
or U10542 (N_10542,N_10149,N_10310);
nand U10543 (N_10543,N_10061,N_10465);
nor U10544 (N_10544,N_10016,N_10028);
or U10545 (N_10545,N_10117,N_10331);
nor U10546 (N_10546,N_10428,N_10235);
nor U10547 (N_10547,N_10050,N_10153);
or U10548 (N_10548,N_10306,N_10233);
nand U10549 (N_10549,N_10260,N_10154);
nor U10550 (N_10550,N_10378,N_10388);
and U10551 (N_10551,N_10146,N_10442);
or U10552 (N_10552,N_10494,N_10278);
or U10553 (N_10553,N_10430,N_10187);
nor U10554 (N_10554,N_10274,N_10344);
and U10555 (N_10555,N_10375,N_10067);
nor U10556 (N_10556,N_10266,N_10387);
nor U10557 (N_10557,N_10170,N_10226);
nor U10558 (N_10558,N_10196,N_10079);
nand U10559 (N_10559,N_10486,N_10321);
xor U10560 (N_10560,N_10263,N_10114);
or U10561 (N_10561,N_10276,N_10106);
and U10562 (N_10562,N_10395,N_10185);
nand U10563 (N_10563,N_10102,N_10407);
or U10564 (N_10564,N_10290,N_10270);
or U10565 (N_10565,N_10257,N_10133);
nor U10566 (N_10566,N_10418,N_10218);
xnor U10567 (N_10567,N_10220,N_10362);
nor U10568 (N_10568,N_10330,N_10223);
and U10569 (N_10569,N_10297,N_10289);
nand U10570 (N_10570,N_10077,N_10066);
or U10571 (N_10571,N_10481,N_10021);
nand U10572 (N_10572,N_10359,N_10318);
xnor U10573 (N_10573,N_10404,N_10248);
nand U10574 (N_10574,N_10495,N_10315);
xor U10575 (N_10575,N_10325,N_10460);
nand U10576 (N_10576,N_10323,N_10026);
xnor U10577 (N_10577,N_10483,N_10010);
xor U10578 (N_10578,N_10160,N_10355);
and U10579 (N_10579,N_10097,N_10155);
xor U10580 (N_10580,N_10178,N_10497);
or U10581 (N_10581,N_10195,N_10340);
and U10582 (N_10582,N_10346,N_10143);
nand U10583 (N_10583,N_10070,N_10212);
nand U10584 (N_10584,N_10057,N_10134);
nand U10585 (N_10585,N_10271,N_10064);
and U10586 (N_10586,N_10227,N_10164);
xnor U10587 (N_10587,N_10374,N_10009);
or U10588 (N_10588,N_10056,N_10239);
or U10589 (N_10589,N_10142,N_10255);
and U10590 (N_10590,N_10286,N_10384);
and U10591 (N_10591,N_10048,N_10482);
nor U10592 (N_10592,N_10124,N_10437);
xor U10593 (N_10593,N_10150,N_10194);
nand U10594 (N_10594,N_10243,N_10105);
nor U10595 (N_10595,N_10034,N_10457);
xnor U10596 (N_10596,N_10471,N_10192);
nor U10597 (N_10597,N_10332,N_10366);
nand U10598 (N_10598,N_10242,N_10103);
nor U10599 (N_10599,N_10267,N_10209);
xnor U10600 (N_10600,N_10072,N_10406);
xor U10601 (N_10601,N_10367,N_10368);
or U10602 (N_10602,N_10408,N_10145);
and U10603 (N_10603,N_10120,N_10249);
nor U10604 (N_10604,N_10204,N_10333);
or U10605 (N_10605,N_10207,N_10458);
or U10606 (N_10606,N_10080,N_10400);
nor U10607 (N_10607,N_10132,N_10347);
xnor U10608 (N_10608,N_10025,N_10397);
nor U10609 (N_10609,N_10261,N_10313);
or U10610 (N_10610,N_10151,N_10165);
and U10611 (N_10611,N_10162,N_10055);
xor U10612 (N_10612,N_10104,N_10329);
xor U10613 (N_10613,N_10431,N_10035);
xor U10614 (N_10614,N_10307,N_10033);
xor U10615 (N_10615,N_10489,N_10083);
and U10616 (N_10616,N_10463,N_10295);
nor U10617 (N_10617,N_10454,N_10370);
xor U10618 (N_10618,N_10314,N_10225);
xor U10619 (N_10619,N_10075,N_10047);
and U10620 (N_10620,N_10475,N_10396);
or U10621 (N_10621,N_10380,N_10413);
or U10622 (N_10622,N_10383,N_10175);
nor U10623 (N_10623,N_10065,N_10063);
and U10624 (N_10624,N_10335,N_10345);
nor U10625 (N_10625,N_10247,N_10293);
nor U10626 (N_10626,N_10138,N_10446);
or U10627 (N_10627,N_10349,N_10089);
or U10628 (N_10628,N_10485,N_10451);
and U10629 (N_10629,N_10308,N_10296);
nor U10630 (N_10630,N_10445,N_10254);
or U10631 (N_10631,N_10012,N_10090);
nor U10632 (N_10632,N_10181,N_10348);
or U10633 (N_10633,N_10377,N_10180);
or U10634 (N_10634,N_10427,N_10499);
and U10635 (N_10635,N_10280,N_10043);
and U10636 (N_10636,N_10099,N_10173);
and U10637 (N_10637,N_10203,N_10379);
and U10638 (N_10638,N_10128,N_10493);
nand U10639 (N_10639,N_10405,N_10208);
xor U10640 (N_10640,N_10419,N_10206);
and U10641 (N_10641,N_10219,N_10302);
or U10642 (N_10642,N_10275,N_10484);
or U10643 (N_10643,N_10328,N_10197);
or U10644 (N_10644,N_10269,N_10262);
or U10645 (N_10645,N_10452,N_10007);
nor U10646 (N_10646,N_10129,N_10320);
nand U10647 (N_10647,N_10391,N_10244);
and U10648 (N_10648,N_10073,N_10455);
xnor U10649 (N_10649,N_10496,N_10024);
or U10650 (N_10650,N_10358,N_10127);
nor U10651 (N_10651,N_10199,N_10364);
and U10652 (N_10652,N_10415,N_10312);
or U10653 (N_10653,N_10441,N_10322);
nor U10654 (N_10654,N_10300,N_10110);
or U10655 (N_10655,N_10352,N_10213);
and U10656 (N_10656,N_10283,N_10190);
nor U10657 (N_10657,N_10477,N_10214);
nor U10658 (N_10658,N_10301,N_10422);
xor U10659 (N_10659,N_10373,N_10139);
or U10660 (N_10660,N_10447,N_10444);
or U10661 (N_10661,N_10032,N_10393);
and U10662 (N_10662,N_10005,N_10041);
and U10663 (N_10663,N_10381,N_10469);
xnor U10664 (N_10664,N_10107,N_10238);
nand U10665 (N_10665,N_10424,N_10023);
or U10666 (N_10666,N_10147,N_10030);
nor U10667 (N_10667,N_10144,N_10081);
nand U10668 (N_10668,N_10264,N_10360);
nand U10669 (N_10669,N_10479,N_10159);
nor U10670 (N_10670,N_10062,N_10287);
or U10671 (N_10671,N_10284,N_10152);
xnor U10672 (N_10672,N_10088,N_10037);
or U10673 (N_10673,N_10052,N_10042);
and U10674 (N_10674,N_10324,N_10319);
nor U10675 (N_10675,N_10417,N_10074);
nor U10676 (N_10676,N_10291,N_10326);
or U10677 (N_10677,N_10311,N_10093);
nand U10678 (N_10678,N_10018,N_10001);
nand U10679 (N_10679,N_10402,N_10459);
or U10680 (N_10680,N_10389,N_10112);
or U10681 (N_10681,N_10245,N_10118);
xnor U10682 (N_10682,N_10158,N_10435);
or U10683 (N_10683,N_10100,N_10019);
nor U10684 (N_10684,N_10163,N_10365);
and U10685 (N_10685,N_10443,N_10473);
or U10686 (N_10686,N_10426,N_10240);
nor U10687 (N_10687,N_10464,N_10131);
nor U10688 (N_10688,N_10176,N_10337);
and U10689 (N_10689,N_10008,N_10282);
xnor U10690 (N_10690,N_10086,N_10234);
nor U10691 (N_10691,N_10013,N_10421);
and U10692 (N_10692,N_10470,N_10191);
xnor U10693 (N_10693,N_10098,N_10182);
xor U10694 (N_10694,N_10394,N_10038);
or U10695 (N_10695,N_10096,N_10303);
or U10696 (N_10696,N_10438,N_10403);
xor U10697 (N_10697,N_10292,N_10039);
or U10698 (N_10698,N_10140,N_10309);
xnor U10699 (N_10699,N_10174,N_10161);
or U10700 (N_10700,N_10188,N_10084);
xnor U10701 (N_10701,N_10434,N_10135);
and U10702 (N_10702,N_10224,N_10166);
and U10703 (N_10703,N_10002,N_10236);
xnor U10704 (N_10704,N_10363,N_10108);
nor U10705 (N_10705,N_10372,N_10049);
nor U10706 (N_10706,N_10253,N_10156);
nand U10707 (N_10707,N_10299,N_10371);
nand U10708 (N_10708,N_10092,N_10461);
or U10709 (N_10709,N_10141,N_10027);
xnor U10710 (N_10710,N_10020,N_10115);
and U10711 (N_10711,N_10091,N_10022);
or U10712 (N_10712,N_10184,N_10193);
or U10713 (N_10713,N_10456,N_10488);
xnor U10714 (N_10714,N_10433,N_10044);
nand U10715 (N_10715,N_10210,N_10231);
nand U10716 (N_10716,N_10356,N_10429);
xor U10717 (N_10717,N_10228,N_10252);
and U10718 (N_10718,N_10382,N_10298);
or U10719 (N_10719,N_10003,N_10229);
and U10720 (N_10720,N_10186,N_10054);
nand U10721 (N_10721,N_10423,N_10412);
xor U10722 (N_10722,N_10492,N_10480);
and U10723 (N_10723,N_10439,N_10136);
xor U10724 (N_10724,N_10060,N_10126);
and U10725 (N_10725,N_10491,N_10334);
and U10726 (N_10726,N_10068,N_10222);
and U10727 (N_10727,N_10316,N_10409);
nand U10728 (N_10728,N_10357,N_10350);
nor U10729 (N_10729,N_10095,N_10420);
and U10730 (N_10730,N_10425,N_10376);
nor U10731 (N_10731,N_10241,N_10216);
nor U10732 (N_10732,N_10059,N_10462);
nand U10733 (N_10733,N_10392,N_10101);
and U10734 (N_10734,N_10468,N_10398);
nand U10735 (N_10735,N_10478,N_10230);
nor U10736 (N_10736,N_10338,N_10046);
xnor U10737 (N_10737,N_10011,N_10259);
nor U10738 (N_10738,N_10053,N_10172);
or U10739 (N_10739,N_10336,N_10432);
nand U10740 (N_10740,N_10448,N_10137);
or U10741 (N_10741,N_10017,N_10466);
or U10742 (N_10742,N_10217,N_10169);
and U10743 (N_10743,N_10343,N_10004);
nand U10744 (N_10744,N_10148,N_10000);
and U10745 (N_10745,N_10279,N_10440);
nor U10746 (N_10746,N_10258,N_10256);
xnor U10747 (N_10747,N_10339,N_10071);
or U10748 (N_10748,N_10200,N_10031);
nand U10749 (N_10749,N_10369,N_10078);
or U10750 (N_10750,N_10250,N_10108);
or U10751 (N_10751,N_10289,N_10248);
nor U10752 (N_10752,N_10489,N_10354);
nor U10753 (N_10753,N_10285,N_10141);
and U10754 (N_10754,N_10038,N_10148);
xor U10755 (N_10755,N_10152,N_10415);
and U10756 (N_10756,N_10070,N_10284);
nand U10757 (N_10757,N_10223,N_10440);
nor U10758 (N_10758,N_10042,N_10341);
nor U10759 (N_10759,N_10261,N_10141);
xnor U10760 (N_10760,N_10464,N_10200);
or U10761 (N_10761,N_10405,N_10325);
or U10762 (N_10762,N_10091,N_10237);
and U10763 (N_10763,N_10236,N_10491);
nor U10764 (N_10764,N_10269,N_10418);
xnor U10765 (N_10765,N_10399,N_10360);
or U10766 (N_10766,N_10485,N_10350);
nor U10767 (N_10767,N_10091,N_10355);
nand U10768 (N_10768,N_10480,N_10406);
nor U10769 (N_10769,N_10260,N_10385);
nor U10770 (N_10770,N_10282,N_10118);
and U10771 (N_10771,N_10189,N_10203);
nor U10772 (N_10772,N_10254,N_10036);
nor U10773 (N_10773,N_10240,N_10283);
and U10774 (N_10774,N_10222,N_10004);
and U10775 (N_10775,N_10312,N_10368);
and U10776 (N_10776,N_10404,N_10423);
xnor U10777 (N_10777,N_10110,N_10229);
nand U10778 (N_10778,N_10296,N_10092);
or U10779 (N_10779,N_10095,N_10418);
or U10780 (N_10780,N_10424,N_10074);
nand U10781 (N_10781,N_10343,N_10295);
xor U10782 (N_10782,N_10204,N_10005);
and U10783 (N_10783,N_10460,N_10429);
and U10784 (N_10784,N_10039,N_10115);
and U10785 (N_10785,N_10079,N_10418);
nand U10786 (N_10786,N_10496,N_10064);
nand U10787 (N_10787,N_10193,N_10037);
or U10788 (N_10788,N_10247,N_10133);
and U10789 (N_10789,N_10092,N_10185);
nand U10790 (N_10790,N_10360,N_10152);
xnor U10791 (N_10791,N_10486,N_10298);
nand U10792 (N_10792,N_10381,N_10137);
nor U10793 (N_10793,N_10485,N_10093);
and U10794 (N_10794,N_10416,N_10443);
and U10795 (N_10795,N_10068,N_10232);
and U10796 (N_10796,N_10181,N_10124);
nor U10797 (N_10797,N_10189,N_10151);
nand U10798 (N_10798,N_10118,N_10399);
nor U10799 (N_10799,N_10005,N_10074);
nand U10800 (N_10800,N_10233,N_10005);
and U10801 (N_10801,N_10152,N_10320);
and U10802 (N_10802,N_10108,N_10362);
or U10803 (N_10803,N_10435,N_10037);
nand U10804 (N_10804,N_10349,N_10374);
or U10805 (N_10805,N_10170,N_10199);
xnor U10806 (N_10806,N_10281,N_10033);
or U10807 (N_10807,N_10499,N_10168);
nand U10808 (N_10808,N_10099,N_10113);
xnor U10809 (N_10809,N_10286,N_10073);
nand U10810 (N_10810,N_10117,N_10238);
or U10811 (N_10811,N_10289,N_10338);
xor U10812 (N_10812,N_10360,N_10176);
nand U10813 (N_10813,N_10015,N_10276);
xnor U10814 (N_10814,N_10114,N_10477);
or U10815 (N_10815,N_10083,N_10164);
xnor U10816 (N_10816,N_10121,N_10088);
xnor U10817 (N_10817,N_10234,N_10160);
and U10818 (N_10818,N_10431,N_10053);
and U10819 (N_10819,N_10396,N_10305);
and U10820 (N_10820,N_10347,N_10349);
or U10821 (N_10821,N_10333,N_10248);
nand U10822 (N_10822,N_10434,N_10040);
nand U10823 (N_10823,N_10129,N_10391);
nor U10824 (N_10824,N_10406,N_10371);
xnor U10825 (N_10825,N_10427,N_10289);
or U10826 (N_10826,N_10082,N_10268);
xor U10827 (N_10827,N_10158,N_10153);
xor U10828 (N_10828,N_10107,N_10293);
and U10829 (N_10829,N_10157,N_10194);
or U10830 (N_10830,N_10065,N_10175);
nand U10831 (N_10831,N_10157,N_10400);
nor U10832 (N_10832,N_10331,N_10327);
or U10833 (N_10833,N_10093,N_10103);
nor U10834 (N_10834,N_10013,N_10370);
or U10835 (N_10835,N_10026,N_10442);
or U10836 (N_10836,N_10361,N_10150);
and U10837 (N_10837,N_10069,N_10084);
nand U10838 (N_10838,N_10422,N_10054);
xor U10839 (N_10839,N_10137,N_10210);
and U10840 (N_10840,N_10177,N_10181);
xnor U10841 (N_10841,N_10317,N_10366);
nor U10842 (N_10842,N_10293,N_10121);
xnor U10843 (N_10843,N_10061,N_10161);
and U10844 (N_10844,N_10324,N_10265);
nand U10845 (N_10845,N_10401,N_10381);
nand U10846 (N_10846,N_10304,N_10462);
nand U10847 (N_10847,N_10367,N_10030);
nand U10848 (N_10848,N_10393,N_10471);
or U10849 (N_10849,N_10266,N_10144);
or U10850 (N_10850,N_10414,N_10300);
nand U10851 (N_10851,N_10350,N_10471);
nand U10852 (N_10852,N_10207,N_10470);
and U10853 (N_10853,N_10324,N_10202);
or U10854 (N_10854,N_10266,N_10157);
or U10855 (N_10855,N_10385,N_10463);
and U10856 (N_10856,N_10499,N_10398);
and U10857 (N_10857,N_10161,N_10436);
and U10858 (N_10858,N_10181,N_10029);
xor U10859 (N_10859,N_10186,N_10194);
nor U10860 (N_10860,N_10228,N_10453);
nand U10861 (N_10861,N_10111,N_10234);
nand U10862 (N_10862,N_10045,N_10419);
nor U10863 (N_10863,N_10111,N_10239);
or U10864 (N_10864,N_10176,N_10046);
or U10865 (N_10865,N_10374,N_10227);
or U10866 (N_10866,N_10245,N_10433);
or U10867 (N_10867,N_10010,N_10150);
nand U10868 (N_10868,N_10012,N_10163);
nor U10869 (N_10869,N_10304,N_10415);
xnor U10870 (N_10870,N_10237,N_10207);
and U10871 (N_10871,N_10106,N_10498);
nand U10872 (N_10872,N_10299,N_10055);
and U10873 (N_10873,N_10457,N_10031);
nand U10874 (N_10874,N_10096,N_10497);
nor U10875 (N_10875,N_10383,N_10381);
or U10876 (N_10876,N_10459,N_10091);
or U10877 (N_10877,N_10345,N_10209);
and U10878 (N_10878,N_10186,N_10386);
xor U10879 (N_10879,N_10126,N_10077);
nand U10880 (N_10880,N_10293,N_10452);
nand U10881 (N_10881,N_10205,N_10499);
xor U10882 (N_10882,N_10429,N_10087);
xnor U10883 (N_10883,N_10352,N_10481);
xnor U10884 (N_10884,N_10332,N_10081);
and U10885 (N_10885,N_10246,N_10201);
and U10886 (N_10886,N_10450,N_10473);
nand U10887 (N_10887,N_10339,N_10185);
nand U10888 (N_10888,N_10147,N_10427);
and U10889 (N_10889,N_10206,N_10285);
and U10890 (N_10890,N_10174,N_10108);
xnor U10891 (N_10891,N_10064,N_10155);
or U10892 (N_10892,N_10069,N_10214);
and U10893 (N_10893,N_10162,N_10062);
xnor U10894 (N_10894,N_10099,N_10186);
and U10895 (N_10895,N_10255,N_10371);
nor U10896 (N_10896,N_10207,N_10203);
and U10897 (N_10897,N_10212,N_10176);
xor U10898 (N_10898,N_10401,N_10158);
or U10899 (N_10899,N_10217,N_10188);
and U10900 (N_10900,N_10081,N_10208);
and U10901 (N_10901,N_10324,N_10067);
xor U10902 (N_10902,N_10405,N_10365);
and U10903 (N_10903,N_10426,N_10036);
or U10904 (N_10904,N_10113,N_10173);
or U10905 (N_10905,N_10405,N_10299);
xor U10906 (N_10906,N_10252,N_10355);
and U10907 (N_10907,N_10187,N_10147);
or U10908 (N_10908,N_10360,N_10151);
and U10909 (N_10909,N_10312,N_10262);
xnor U10910 (N_10910,N_10470,N_10351);
or U10911 (N_10911,N_10128,N_10421);
and U10912 (N_10912,N_10241,N_10487);
nand U10913 (N_10913,N_10058,N_10303);
xnor U10914 (N_10914,N_10429,N_10449);
or U10915 (N_10915,N_10490,N_10260);
and U10916 (N_10916,N_10243,N_10340);
nand U10917 (N_10917,N_10041,N_10296);
xnor U10918 (N_10918,N_10350,N_10484);
nand U10919 (N_10919,N_10209,N_10188);
or U10920 (N_10920,N_10255,N_10471);
nand U10921 (N_10921,N_10262,N_10031);
nand U10922 (N_10922,N_10377,N_10302);
or U10923 (N_10923,N_10352,N_10404);
and U10924 (N_10924,N_10344,N_10069);
xnor U10925 (N_10925,N_10369,N_10353);
or U10926 (N_10926,N_10482,N_10151);
nand U10927 (N_10927,N_10091,N_10239);
nor U10928 (N_10928,N_10332,N_10466);
or U10929 (N_10929,N_10371,N_10481);
and U10930 (N_10930,N_10120,N_10356);
and U10931 (N_10931,N_10387,N_10172);
xor U10932 (N_10932,N_10096,N_10473);
nand U10933 (N_10933,N_10028,N_10348);
xnor U10934 (N_10934,N_10480,N_10125);
and U10935 (N_10935,N_10242,N_10288);
nand U10936 (N_10936,N_10410,N_10152);
and U10937 (N_10937,N_10000,N_10277);
or U10938 (N_10938,N_10237,N_10415);
nand U10939 (N_10939,N_10140,N_10125);
nor U10940 (N_10940,N_10466,N_10181);
xnor U10941 (N_10941,N_10253,N_10098);
and U10942 (N_10942,N_10020,N_10151);
xnor U10943 (N_10943,N_10465,N_10407);
and U10944 (N_10944,N_10201,N_10304);
nand U10945 (N_10945,N_10249,N_10462);
nor U10946 (N_10946,N_10486,N_10279);
or U10947 (N_10947,N_10435,N_10341);
xor U10948 (N_10948,N_10364,N_10041);
nand U10949 (N_10949,N_10256,N_10050);
or U10950 (N_10950,N_10284,N_10458);
nor U10951 (N_10951,N_10369,N_10230);
nor U10952 (N_10952,N_10217,N_10183);
or U10953 (N_10953,N_10380,N_10430);
nand U10954 (N_10954,N_10204,N_10188);
nand U10955 (N_10955,N_10270,N_10288);
and U10956 (N_10956,N_10106,N_10442);
nand U10957 (N_10957,N_10172,N_10382);
or U10958 (N_10958,N_10190,N_10173);
nand U10959 (N_10959,N_10242,N_10035);
and U10960 (N_10960,N_10314,N_10001);
nand U10961 (N_10961,N_10255,N_10467);
and U10962 (N_10962,N_10458,N_10371);
and U10963 (N_10963,N_10179,N_10005);
xnor U10964 (N_10964,N_10323,N_10437);
xnor U10965 (N_10965,N_10047,N_10207);
and U10966 (N_10966,N_10368,N_10035);
nor U10967 (N_10967,N_10133,N_10220);
or U10968 (N_10968,N_10489,N_10313);
nor U10969 (N_10969,N_10054,N_10479);
or U10970 (N_10970,N_10137,N_10073);
and U10971 (N_10971,N_10256,N_10113);
nand U10972 (N_10972,N_10338,N_10366);
nor U10973 (N_10973,N_10099,N_10331);
nor U10974 (N_10974,N_10104,N_10485);
xor U10975 (N_10975,N_10348,N_10304);
and U10976 (N_10976,N_10240,N_10059);
and U10977 (N_10977,N_10049,N_10099);
nand U10978 (N_10978,N_10221,N_10455);
and U10979 (N_10979,N_10386,N_10168);
nand U10980 (N_10980,N_10407,N_10038);
nand U10981 (N_10981,N_10192,N_10459);
xor U10982 (N_10982,N_10027,N_10257);
and U10983 (N_10983,N_10495,N_10382);
nand U10984 (N_10984,N_10319,N_10126);
or U10985 (N_10985,N_10314,N_10326);
and U10986 (N_10986,N_10110,N_10461);
xnor U10987 (N_10987,N_10423,N_10469);
xnor U10988 (N_10988,N_10292,N_10029);
nor U10989 (N_10989,N_10318,N_10369);
xor U10990 (N_10990,N_10360,N_10443);
nand U10991 (N_10991,N_10317,N_10064);
nand U10992 (N_10992,N_10276,N_10090);
nor U10993 (N_10993,N_10046,N_10416);
xor U10994 (N_10994,N_10094,N_10414);
or U10995 (N_10995,N_10163,N_10090);
nand U10996 (N_10996,N_10128,N_10263);
and U10997 (N_10997,N_10195,N_10410);
and U10998 (N_10998,N_10196,N_10091);
and U10999 (N_10999,N_10209,N_10223);
or U11000 (N_11000,N_10692,N_10672);
xnor U11001 (N_11001,N_10988,N_10690);
nand U11002 (N_11002,N_10733,N_10643);
nor U11003 (N_11003,N_10644,N_10572);
nor U11004 (N_11004,N_10822,N_10786);
and U11005 (N_11005,N_10696,N_10561);
or U11006 (N_11006,N_10542,N_10548);
or U11007 (N_11007,N_10916,N_10889);
nor U11008 (N_11008,N_10607,N_10848);
nand U11009 (N_11009,N_10769,N_10566);
nor U11010 (N_11010,N_10519,N_10784);
nor U11011 (N_11011,N_10789,N_10703);
or U11012 (N_11012,N_10544,N_10509);
and U11013 (N_11013,N_10899,N_10759);
and U11014 (N_11014,N_10637,N_10511);
nand U11015 (N_11015,N_10730,N_10755);
or U11016 (N_11016,N_10907,N_10807);
nor U11017 (N_11017,N_10657,N_10795);
and U11018 (N_11018,N_10876,N_10568);
xor U11019 (N_11019,N_10628,N_10772);
nor U11020 (N_11020,N_10977,N_10638);
and U11021 (N_11021,N_10560,N_10714);
and U11022 (N_11022,N_10586,N_10629);
or U11023 (N_11023,N_10526,N_10716);
or U11024 (N_11024,N_10990,N_10964);
and U11025 (N_11025,N_10861,N_10559);
xor U11026 (N_11026,N_10891,N_10982);
and U11027 (N_11027,N_10513,N_10894);
and U11028 (N_11028,N_10871,N_10865);
xor U11029 (N_11029,N_10870,N_10507);
nor U11030 (N_11030,N_10588,N_10743);
nand U11031 (N_11031,N_10806,N_10677);
or U11032 (N_11032,N_10660,N_10585);
or U11033 (N_11033,N_10664,N_10661);
and U11034 (N_11034,N_10869,N_10771);
nand U11035 (N_11035,N_10847,N_10997);
xnor U11036 (N_11036,N_10911,N_10785);
xor U11037 (N_11037,N_10597,N_10550);
xnor U11038 (N_11038,N_10831,N_10909);
nand U11039 (N_11039,N_10739,N_10875);
or U11040 (N_11040,N_10545,N_10591);
xor U11041 (N_11041,N_10781,N_10906);
or U11042 (N_11042,N_10797,N_10926);
and U11043 (N_11043,N_10808,N_10898);
and U11044 (N_11044,N_10540,N_10543);
or U11045 (N_11045,N_10860,N_10726);
xor U11046 (N_11046,N_10980,N_10592);
and U11047 (N_11047,N_10652,N_10611);
nor U11048 (N_11048,N_10882,N_10681);
nand U11049 (N_11049,N_10727,N_10745);
or U11050 (N_11050,N_10910,N_10972);
and U11051 (N_11051,N_10843,N_10636);
nor U11052 (N_11052,N_10842,N_10541);
nor U11053 (N_11053,N_10828,N_10646);
nand U11054 (N_11054,N_10760,N_10697);
or U11055 (N_11055,N_10930,N_10707);
nor U11056 (N_11056,N_10883,N_10874);
nor U11057 (N_11057,N_10959,N_10546);
xor U11058 (N_11058,N_10558,N_10617);
or U11059 (N_11059,N_10709,N_10500);
xor U11060 (N_11060,N_10694,N_10944);
and U11061 (N_11061,N_10937,N_10956);
or U11062 (N_11062,N_10762,N_10927);
nand U11063 (N_11063,N_10804,N_10616);
and U11064 (N_11064,N_10567,N_10678);
or U11065 (N_11065,N_10684,N_10634);
and U11066 (N_11066,N_10656,N_10994);
nor U11067 (N_11067,N_10897,N_10817);
or U11068 (N_11068,N_10605,N_10724);
and U11069 (N_11069,N_10867,N_10763);
nand U11070 (N_11070,N_10734,N_10987);
xor U11071 (N_11071,N_10649,N_10823);
or U11072 (N_11072,N_10630,N_10565);
nor U11073 (N_11073,N_10878,N_10764);
nor U11074 (N_11074,N_10779,N_10814);
nand U11075 (N_11075,N_10737,N_10534);
nor U11076 (N_11076,N_10527,N_10928);
xnor U11077 (N_11077,N_10603,N_10816);
and U11078 (N_11078,N_10662,N_10648);
or U11079 (N_11079,N_10529,N_10711);
xnor U11080 (N_11080,N_10936,N_10757);
nor U11081 (N_11081,N_10720,N_10675);
or U11082 (N_11082,N_10986,N_10820);
and U11083 (N_11083,N_10575,N_10756);
xor U11084 (N_11084,N_10556,N_10587);
xor U11085 (N_11085,N_10901,N_10788);
nand U11086 (N_11086,N_10794,N_10787);
xnor U11087 (N_11087,N_10551,N_10969);
and U11088 (N_11088,N_10706,N_10562);
nor U11089 (N_11089,N_10674,N_10908);
nand U11090 (N_11090,N_10925,N_10792);
or U11091 (N_11091,N_10800,N_10844);
xnor U11092 (N_11092,N_10516,N_10905);
and U11093 (N_11093,N_10531,N_10502);
and U11094 (N_11094,N_10705,N_10836);
nand U11095 (N_11095,N_10922,N_10945);
and U11096 (N_11096,N_10748,N_10967);
nand U11097 (N_11097,N_10879,N_10719);
xnor U11098 (N_11098,N_10921,N_10647);
or U11099 (N_11099,N_10829,N_10695);
or U11100 (N_11100,N_10934,N_10608);
xnor U11101 (N_11101,N_10975,N_10515);
xor U11102 (N_11102,N_10949,N_10991);
nand U11103 (N_11103,N_10614,N_10747);
or U11104 (N_11104,N_10583,N_10783);
xor U11105 (N_11105,N_10824,N_10951);
and U11106 (N_11106,N_10581,N_10753);
and U11107 (N_11107,N_10538,N_10810);
and U11108 (N_11108,N_10974,N_10573);
nand U11109 (N_11109,N_10752,N_10732);
nor U11110 (N_11110,N_10669,N_10963);
or U11111 (N_11111,N_10853,N_10774);
nand U11112 (N_11112,N_10852,N_10738);
or U11113 (N_11113,N_10746,N_10893);
or U11114 (N_11114,N_10813,N_10731);
nor U11115 (N_11115,N_10532,N_10593);
and U11116 (N_11116,N_10621,N_10523);
xor U11117 (N_11117,N_10995,N_10520);
nand U11118 (N_11118,N_10576,N_10710);
nand U11119 (N_11119,N_10873,N_10768);
or U11120 (N_11120,N_10650,N_10954);
or U11121 (N_11121,N_10903,N_10506);
or U11122 (N_11122,N_10832,N_10815);
or U11123 (N_11123,N_10924,N_10658);
and U11124 (N_11124,N_10863,N_10984);
nor U11125 (N_11125,N_10704,N_10553);
xor U11126 (N_11126,N_10659,N_10501);
nand U11127 (N_11127,N_10943,N_10862);
and U11128 (N_11128,N_10686,N_10931);
nor U11129 (N_11129,N_10596,N_10981);
and U11130 (N_11130,N_10849,N_10979);
or U11131 (N_11131,N_10670,N_10840);
and U11132 (N_11132,N_10618,N_10761);
or U11133 (N_11133,N_10868,N_10537);
nand U11134 (N_11134,N_10758,N_10654);
and U11135 (N_11135,N_10968,N_10741);
nor U11136 (N_11136,N_10530,N_10725);
nand U11137 (N_11137,N_10947,N_10610);
xor U11138 (N_11138,N_10613,N_10850);
xor U11139 (N_11139,N_10595,N_10778);
and U11140 (N_11140,N_10996,N_10971);
or U11141 (N_11141,N_10521,N_10885);
xnor U11142 (N_11142,N_10715,N_10655);
and U11143 (N_11143,N_10735,N_10938);
nor U11144 (N_11144,N_10549,N_10582);
xor U11145 (N_11145,N_10528,N_10533);
xor U11146 (N_11146,N_10872,N_10625);
nand U11147 (N_11147,N_10750,N_10590);
or U11148 (N_11148,N_10612,N_10830);
and U11149 (N_11149,N_10913,N_10886);
and U11150 (N_11150,N_10970,N_10615);
or U11151 (N_11151,N_10881,N_10525);
xor U11152 (N_11152,N_10798,N_10594);
and U11153 (N_11153,N_10702,N_10554);
and U11154 (N_11154,N_10536,N_10819);
nand U11155 (N_11155,N_10856,N_10888);
and U11156 (N_11156,N_10973,N_10833);
nor U11157 (N_11157,N_10604,N_10791);
nor U11158 (N_11158,N_10939,N_10834);
or U11159 (N_11159,N_10854,N_10818);
or U11160 (N_11160,N_10632,N_10866);
and U11161 (N_11161,N_10622,N_10505);
nand U11162 (N_11162,N_10915,N_10689);
nor U11163 (N_11163,N_10929,N_10917);
nand U11164 (N_11164,N_10811,N_10701);
xor U11165 (N_11165,N_10522,N_10920);
or U11166 (N_11166,N_10902,N_10639);
and U11167 (N_11167,N_10932,N_10952);
nand U11168 (N_11168,N_10742,N_10671);
nor U11169 (N_11169,N_10827,N_10773);
and U11170 (N_11170,N_10645,N_10524);
xnor U11171 (N_11171,N_10775,N_10978);
or U11172 (N_11172,N_10599,N_10635);
or U11173 (N_11173,N_10691,N_10896);
nor U11174 (N_11174,N_10626,N_10600);
nand U11175 (N_11175,N_10744,N_10623);
nor U11176 (N_11176,N_10557,N_10825);
xnor U11177 (N_11177,N_10942,N_10729);
nor U11178 (N_11178,N_10989,N_10601);
nor U11179 (N_11179,N_10589,N_10858);
and U11180 (N_11180,N_10957,N_10780);
nand U11181 (N_11181,N_10579,N_10803);
xnor U11182 (N_11182,N_10877,N_10514);
or U11183 (N_11183,N_10777,N_10776);
xnor U11184 (N_11184,N_10712,N_10754);
nand U11185 (N_11185,N_10721,N_10552);
xor U11186 (N_11186,N_10838,N_10682);
or U11187 (N_11187,N_10539,N_10884);
nand U11188 (N_11188,N_10687,N_10580);
and U11189 (N_11189,N_10976,N_10736);
or U11190 (N_11190,N_10676,N_10950);
xnor U11191 (N_11191,N_10578,N_10518);
and U11192 (N_11192,N_10504,N_10574);
nor U11193 (N_11193,N_10890,N_10793);
nor U11194 (N_11194,N_10673,N_10683);
xnor U11195 (N_11195,N_10722,N_10801);
nand U11196 (N_11196,N_10700,N_10598);
or U11197 (N_11197,N_10919,N_10923);
or U11198 (N_11198,N_10713,N_10627);
or U11199 (N_11199,N_10826,N_10508);
or U11200 (N_11200,N_10992,N_10859);
or U11201 (N_11201,N_10892,N_10855);
nand U11202 (N_11202,N_10966,N_10584);
and U11203 (N_11203,N_10728,N_10510);
and U11204 (N_11204,N_10953,N_10851);
xor U11205 (N_11205,N_10933,N_10985);
or U11206 (N_11206,N_10837,N_10993);
nor U11207 (N_11207,N_10631,N_10941);
nand U11208 (N_11208,N_10503,N_10961);
nand U11209 (N_11209,N_10609,N_10846);
xnor U11210 (N_11210,N_10965,N_10679);
and U11211 (N_11211,N_10708,N_10606);
nand U11212 (N_11212,N_10718,N_10940);
nor U11213 (N_11213,N_10960,N_10958);
nand U11214 (N_11214,N_10749,N_10571);
nor U11215 (N_11215,N_10802,N_10962);
nand U11216 (N_11216,N_10914,N_10563);
nor U11217 (N_11217,N_10577,N_10880);
xor U11218 (N_11218,N_10895,N_10935);
nor U11219 (N_11219,N_10887,N_10766);
nor U11220 (N_11220,N_10983,N_10782);
and U11221 (N_11221,N_10619,N_10620);
or U11222 (N_11222,N_10821,N_10946);
nor U11223 (N_11223,N_10717,N_10767);
nand U11224 (N_11224,N_10805,N_10665);
and U11225 (N_11225,N_10955,N_10640);
and U11226 (N_11226,N_10948,N_10998);
nand U11227 (N_11227,N_10688,N_10845);
nand U11228 (N_11228,N_10564,N_10624);
nor U11229 (N_11229,N_10751,N_10642);
nor U11230 (N_11230,N_10680,N_10740);
nand U11231 (N_11231,N_10685,N_10693);
or U11232 (N_11232,N_10839,N_10602);
nor U11233 (N_11233,N_10723,N_10770);
nor U11234 (N_11234,N_10812,N_10912);
nand U11235 (N_11235,N_10651,N_10790);
xor U11236 (N_11236,N_10918,N_10512);
nor U11237 (N_11237,N_10799,N_10765);
or U11238 (N_11238,N_10663,N_10547);
and U11239 (N_11239,N_10698,N_10666);
nor U11240 (N_11240,N_10517,N_10570);
xnor U11241 (N_11241,N_10904,N_10900);
and U11242 (N_11242,N_10653,N_10535);
or U11243 (N_11243,N_10667,N_10857);
nand U11244 (N_11244,N_10796,N_10555);
xnor U11245 (N_11245,N_10835,N_10569);
nand U11246 (N_11246,N_10641,N_10809);
or U11247 (N_11247,N_10864,N_10699);
nor U11248 (N_11248,N_10668,N_10633);
and U11249 (N_11249,N_10841,N_10999);
nand U11250 (N_11250,N_10940,N_10563);
and U11251 (N_11251,N_10560,N_10850);
xor U11252 (N_11252,N_10780,N_10804);
nor U11253 (N_11253,N_10927,N_10889);
nor U11254 (N_11254,N_10941,N_10865);
nand U11255 (N_11255,N_10707,N_10830);
and U11256 (N_11256,N_10586,N_10542);
and U11257 (N_11257,N_10532,N_10917);
xnor U11258 (N_11258,N_10566,N_10928);
nand U11259 (N_11259,N_10882,N_10877);
nand U11260 (N_11260,N_10628,N_10950);
and U11261 (N_11261,N_10506,N_10746);
and U11262 (N_11262,N_10808,N_10592);
and U11263 (N_11263,N_10577,N_10908);
and U11264 (N_11264,N_10902,N_10804);
nor U11265 (N_11265,N_10892,N_10789);
nand U11266 (N_11266,N_10863,N_10734);
and U11267 (N_11267,N_10641,N_10672);
nand U11268 (N_11268,N_10785,N_10875);
xnor U11269 (N_11269,N_10886,N_10517);
nand U11270 (N_11270,N_10874,N_10535);
xnor U11271 (N_11271,N_10956,N_10933);
nor U11272 (N_11272,N_10946,N_10650);
and U11273 (N_11273,N_10568,N_10789);
xnor U11274 (N_11274,N_10528,N_10621);
xnor U11275 (N_11275,N_10919,N_10737);
nand U11276 (N_11276,N_10505,N_10659);
xor U11277 (N_11277,N_10685,N_10779);
and U11278 (N_11278,N_10756,N_10937);
or U11279 (N_11279,N_10529,N_10779);
or U11280 (N_11280,N_10821,N_10559);
or U11281 (N_11281,N_10613,N_10912);
xnor U11282 (N_11282,N_10837,N_10603);
nand U11283 (N_11283,N_10781,N_10757);
xnor U11284 (N_11284,N_10744,N_10811);
xnor U11285 (N_11285,N_10732,N_10560);
nor U11286 (N_11286,N_10511,N_10709);
and U11287 (N_11287,N_10720,N_10528);
and U11288 (N_11288,N_10535,N_10652);
xor U11289 (N_11289,N_10793,N_10764);
nand U11290 (N_11290,N_10619,N_10559);
or U11291 (N_11291,N_10953,N_10982);
xor U11292 (N_11292,N_10956,N_10543);
nor U11293 (N_11293,N_10724,N_10751);
nor U11294 (N_11294,N_10610,N_10847);
xnor U11295 (N_11295,N_10736,N_10754);
nand U11296 (N_11296,N_10545,N_10922);
or U11297 (N_11297,N_10980,N_10567);
xor U11298 (N_11298,N_10669,N_10657);
nor U11299 (N_11299,N_10854,N_10639);
and U11300 (N_11300,N_10628,N_10773);
and U11301 (N_11301,N_10948,N_10558);
and U11302 (N_11302,N_10589,N_10622);
nand U11303 (N_11303,N_10948,N_10679);
nand U11304 (N_11304,N_10992,N_10578);
nand U11305 (N_11305,N_10983,N_10649);
nor U11306 (N_11306,N_10850,N_10579);
and U11307 (N_11307,N_10699,N_10737);
xor U11308 (N_11308,N_10821,N_10572);
nor U11309 (N_11309,N_10974,N_10729);
and U11310 (N_11310,N_10794,N_10600);
nand U11311 (N_11311,N_10640,N_10861);
xnor U11312 (N_11312,N_10824,N_10559);
and U11313 (N_11313,N_10585,N_10941);
and U11314 (N_11314,N_10840,N_10690);
nor U11315 (N_11315,N_10659,N_10920);
nand U11316 (N_11316,N_10639,N_10920);
xor U11317 (N_11317,N_10566,N_10975);
or U11318 (N_11318,N_10841,N_10829);
and U11319 (N_11319,N_10603,N_10735);
nand U11320 (N_11320,N_10742,N_10790);
xnor U11321 (N_11321,N_10947,N_10873);
and U11322 (N_11322,N_10792,N_10963);
nor U11323 (N_11323,N_10848,N_10915);
nor U11324 (N_11324,N_10900,N_10768);
nand U11325 (N_11325,N_10590,N_10600);
nor U11326 (N_11326,N_10571,N_10712);
nand U11327 (N_11327,N_10847,N_10871);
and U11328 (N_11328,N_10676,N_10530);
xnor U11329 (N_11329,N_10570,N_10936);
nor U11330 (N_11330,N_10875,N_10673);
and U11331 (N_11331,N_10777,N_10821);
nor U11332 (N_11332,N_10994,N_10883);
nor U11333 (N_11333,N_10877,N_10804);
nand U11334 (N_11334,N_10692,N_10635);
xor U11335 (N_11335,N_10794,N_10762);
nor U11336 (N_11336,N_10593,N_10621);
or U11337 (N_11337,N_10869,N_10728);
or U11338 (N_11338,N_10550,N_10760);
nor U11339 (N_11339,N_10715,N_10992);
nand U11340 (N_11340,N_10941,N_10743);
nand U11341 (N_11341,N_10900,N_10824);
nand U11342 (N_11342,N_10674,N_10850);
nand U11343 (N_11343,N_10621,N_10574);
nor U11344 (N_11344,N_10859,N_10729);
and U11345 (N_11345,N_10930,N_10654);
and U11346 (N_11346,N_10702,N_10572);
and U11347 (N_11347,N_10888,N_10712);
or U11348 (N_11348,N_10897,N_10900);
or U11349 (N_11349,N_10864,N_10745);
xnor U11350 (N_11350,N_10891,N_10723);
nor U11351 (N_11351,N_10546,N_10822);
or U11352 (N_11352,N_10546,N_10536);
and U11353 (N_11353,N_10508,N_10581);
and U11354 (N_11354,N_10992,N_10846);
nand U11355 (N_11355,N_10840,N_10760);
and U11356 (N_11356,N_10672,N_10732);
nand U11357 (N_11357,N_10859,N_10539);
nand U11358 (N_11358,N_10682,N_10839);
nand U11359 (N_11359,N_10622,N_10950);
and U11360 (N_11360,N_10902,N_10832);
and U11361 (N_11361,N_10884,N_10646);
or U11362 (N_11362,N_10723,N_10669);
xnor U11363 (N_11363,N_10900,N_10689);
xnor U11364 (N_11364,N_10534,N_10566);
xor U11365 (N_11365,N_10572,N_10720);
and U11366 (N_11366,N_10815,N_10772);
or U11367 (N_11367,N_10580,N_10574);
and U11368 (N_11368,N_10505,N_10734);
and U11369 (N_11369,N_10972,N_10627);
or U11370 (N_11370,N_10692,N_10997);
nand U11371 (N_11371,N_10587,N_10989);
nand U11372 (N_11372,N_10514,N_10983);
or U11373 (N_11373,N_10751,N_10812);
nand U11374 (N_11374,N_10748,N_10825);
or U11375 (N_11375,N_10626,N_10875);
nand U11376 (N_11376,N_10997,N_10631);
nor U11377 (N_11377,N_10685,N_10856);
xor U11378 (N_11378,N_10971,N_10912);
nand U11379 (N_11379,N_10621,N_10575);
nand U11380 (N_11380,N_10880,N_10772);
nor U11381 (N_11381,N_10539,N_10822);
and U11382 (N_11382,N_10935,N_10522);
nand U11383 (N_11383,N_10714,N_10512);
xor U11384 (N_11384,N_10612,N_10868);
xnor U11385 (N_11385,N_10666,N_10911);
and U11386 (N_11386,N_10916,N_10614);
or U11387 (N_11387,N_10852,N_10581);
and U11388 (N_11388,N_10919,N_10633);
nor U11389 (N_11389,N_10925,N_10576);
nor U11390 (N_11390,N_10633,N_10682);
nor U11391 (N_11391,N_10623,N_10821);
and U11392 (N_11392,N_10732,N_10523);
xnor U11393 (N_11393,N_10814,N_10888);
xor U11394 (N_11394,N_10774,N_10735);
or U11395 (N_11395,N_10715,N_10793);
nor U11396 (N_11396,N_10638,N_10631);
nor U11397 (N_11397,N_10675,N_10823);
nor U11398 (N_11398,N_10773,N_10741);
xnor U11399 (N_11399,N_10934,N_10833);
nor U11400 (N_11400,N_10737,N_10513);
nor U11401 (N_11401,N_10867,N_10992);
nand U11402 (N_11402,N_10645,N_10705);
nand U11403 (N_11403,N_10787,N_10995);
xor U11404 (N_11404,N_10922,N_10780);
and U11405 (N_11405,N_10520,N_10999);
and U11406 (N_11406,N_10864,N_10618);
and U11407 (N_11407,N_10595,N_10535);
and U11408 (N_11408,N_10559,N_10926);
and U11409 (N_11409,N_10839,N_10555);
and U11410 (N_11410,N_10626,N_10677);
xor U11411 (N_11411,N_10906,N_10716);
and U11412 (N_11412,N_10596,N_10736);
or U11413 (N_11413,N_10557,N_10827);
and U11414 (N_11414,N_10612,N_10757);
nor U11415 (N_11415,N_10587,N_10729);
nor U11416 (N_11416,N_10986,N_10753);
xor U11417 (N_11417,N_10767,N_10704);
or U11418 (N_11418,N_10696,N_10570);
or U11419 (N_11419,N_10947,N_10875);
nor U11420 (N_11420,N_10934,N_10685);
and U11421 (N_11421,N_10942,N_10825);
xor U11422 (N_11422,N_10896,N_10731);
and U11423 (N_11423,N_10950,N_10679);
xnor U11424 (N_11424,N_10658,N_10879);
or U11425 (N_11425,N_10703,N_10981);
or U11426 (N_11426,N_10870,N_10616);
nor U11427 (N_11427,N_10523,N_10718);
and U11428 (N_11428,N_10813,N_10938);
nor U11429 (N_11429,N_10587,N_10535);
nand U11430 (N_11430,N_10664,N_10884);
or U11431 (N_11431,N_10864,N_10844);
or U11432 (N_11432,N_10669,N_10796);
nor U11433 (N_11433,N_10840,N_10789);
nand U11434 (N_11434,N_10716,N_10943);
and U11435 (N_11435,N_10580,N_10749);
or U11436 (N_11436,N_10724,N_10967);
or U11437 (N_11437,N_10831,N_10562);
or U11438 (N_11438,N_10735,N_10845);
and U11439 (N_11439,N_10761,N_10957);
and U11440 (N_11440,N_10862,N_10551);
or U11441 (N_11441,N_10783,N_10777);
nand U11442 (N_11442,N_10654,N_10904);
or U11443 (N_11443,N_10533,N_10896);
or U11444 (N_11444,N_10578,N_10559);
nor U11445 (N_11445,N_10996,N_10853);
nand U11446 (N_11446,N_10578,N_10678);
nor U11447 (N_11447,N_10652,N_10621);
xnor U11448 (N_11448,N_10836,N_10738);
nor U11449 (N_11449,N_10684,N_10548);
nand U11450 (N_11450,N_10966,N_10707);
xnor U11451 (N_11451,N_10668,N_10636);
nor U11452 (N_11452,N_10730,N_10524);
nor U11453 (N_11453,N_10506,N_10564);
nor U11454 (N_11454,N_10555,N_10634);
nand U11455 (N_11455,N_10784,N_10988);
and U11456 (N_11456,N_10682,N_10910);
nand U11457 (N_11457,N_10757,N_10503);
or U11458 (N_11458,N_10622,N_10900);
or U11459 (N_11459,N_10574,N_10883);
nor U11460 (N_11460,N_10671,N_10623);
nand U11461 (N_11461,N_10644,N_10781);
or U11462 (N_11462,N_10595,N_10729);
nor U11463 (N_11463,N_10802,N_10873);
or U11464 (N_11464,N_10618,N_10678);
nor U11465 (N_11465,N_10933,N_10731);
nand U11466 (N_11466,N_10902,N_10630);
xnor U11467 (N_11467,N_10947,N_10775);
and U11468 (N_11468,N_10839,N_10897);
nand U11469 (N_11469,N_10981,N_10777);
or U11470 (N_11470,N_10881,N_10503);
and U11471 (N_11471,N_10725,N_10524);
and U11472 (N_11472,N_10657,N_10774);
xnor U11473 (N_11473,N_10948,N_10673);
nor U11474 (N_11474,N_10658,N_10682);
nand U11475 (N_11475,N_10844,N_10874);
nand U11476 (N_11476,N_10551,N_10631);
nor U11477 (N_11477,N_10558,N_10574);
nand U11478 (N_11478,N_10584,N_10634);
nor U11479 (N_11479,N_10631,N_10711);
and U11480 (N_11480,N_10548,N_10960);
and U11481 (N_11481,N_10625,N_10526);
or U11482 (N_11482,N_10900,N_10975);
nand U11483 (N_11483,N_10814,N_10957);
nor U11484 (N_11484,N_10550,N_10775);
xor U11485 (N_11485,N_10925,N_10961);
and U11486 (N_11486,N_10620,N_10608);
and U11487 (N_11487,N_10588,N_10826);
xnor U11488 (N_11488,N_10827,N_10623);
or U11489 (N_11489,N_10981,N_10694);
xnor U11490 (N_11490,N_10600,N_10645);
or U11491 (N_11491,N_10554,N_10526);
and U11492 (N_11492,N_10704,N_10841);
nand U11493 (N_11493,N_10740,N_10986);
and U11494 (N_11494,N_10643,N_10846);
nor U11495 (N_11495,N_10606,N_10787);
xnor U11496 (N_11496,N_10878,N_10766);
or U11497 (N_11497,N_10865,N_10717);
nor U11498 (N_11498,N_10870,N_10642);
or U11499 (N_11499,N_10801,N_10952);
and U11500 (N_11500,N_11393,N_11263);
or U11501 (N_11501,N_11243,N_11394);
xnor U11502 (N_11502,N_11097,N_11045);
xnor U11503 (N_11503,N_11140,N_11298);
or U11504 (N_11504,N_11012,N_11061);
xnor U11505 (N_11505,N_11201,N_11025);
or U11506 (N_11506,N_11489,N_11161);
nor U11507 (N_11507,N_11316,N_11146);
or U11508 (N_11508,N_11129,N_11408);
nor U11509 (N_11509,N_11446,N_11141);
xor U11510 (N_11510,N_11155,N_11160);
nand U11511 (N_11511,N_11142,N_11016);
nor U11512 (N_11512,N_11057,N_11418);
or U11513 (N_11513,N_11184,N_11080);
or U11514 (N_11514,N_11403,N_11302);
xor U11515 (N_11515,N_11048,N_11163);
nor U11516 (N_11516,N_11203,N_11284);
and U11517 (N_11517,N_11391,N_11037);
or U11518 (N_11518,N_11247,N_11328);
nand U11519 (N_11519,N_11484,N_11369);
nand U11520 (N_11520,N_11255,N_11389);
xor U11521 (N_11521,N_11426,N_11058);
or U11522 (N_11522,N_11390,N_11370);
or U11523 (N_11523,N_11183,N_11003);
or U11524 (N_11524,N_11182,N_11299);
or U11525 (N_11525,N_11329,N_11013);
nor U11526 (N_11526,N_11018,N_11111);
nand U11527 (N_11527,N_11441,N_11306);
and U11528 (N_11528,N_11417,N_11377);
and U11529 (N_11529,N_11262,N_11259);
nand U11530 (N_11530,N_11082,N_11421);
nand U11531 (N_11531,N_11143,N_11271);
or U11532 (N_11532,N_11482,N_11404);
nand U11533 (N_11533,N_11215,N_11004);
or U11534 (N_11534,N_11176,N_11413);
or U11535 (N_11535,N_11312,N_11093);
nand U11536 (N_11536,N_11480,N_11091);
nand U11537 (N_11537,N_11440,N_11110);
or U11538 (N_11538,N_11116,N_11118);
or U11539 (N_11539,N_11322,N_11314);
nor U11540 (N_11540,N_11467,N_11291);
and U11541 (N_11541,N_11127,N_11121);
nand U11542 (N_11542,N_11252,N_11178);
and U11543 (N_11543,N_11226,N_11049);
xor U11544 (N_11544,N_11383,N_11065);
and U11545 (N_11545,N_11425,N_11149);
and U11546 (N_11546,N_11485,N_11472);
and U11547 (N_11547,N_11199,N_11217);
or U11548 (N_11548,N_11433,N_11214);
nand U11549 (N_11549,N_11092,N_11332);
and U11550 (N_11550,N_11128,N_11056);
xor U11551 (N_11551,N_11313,N_11274);
or U11552 (N_11552,N_11248,N_11185);
xor U11553 (N_11553,N_11242,N_11103);
xnor U11554 (N_11554,N_11188,N_11179);
or U11555 (N_11555,N_11060,N_11340);
xor U11556 (N_11556,N_11281,N_11364);
and U11557 (N_11557,N_11437,N_11304);
or U11558 (N_11558,N_11114,N_11339);
nand U11559 (N_11559,N_11374,N_11290);
xor U11560 (N_11560,N_11210,N_11360);
nor U11561 (N_11561,N_11450,N_11158);
or U11562 (N_11562,N_11466,N_11355);
and U11563 (N_11563,N_11131,N_11153);
xor U11564 (N_11564,N_11094,N_11227);
or U11565 (N_11565,N_11442,N_11495);
or U11566 (N_11566,N_11475,N_11363);
nor U11567 (N_11567,N_11001,N_11388);
and U11568 (N_11568,N_11245,N_11028);
or U11569 (N_11569,N_11194,N_11017);
and U11570 (N_11570,N_11026,N_11499);
and U11571 (N_11571,N_11392,N_11137);
nor U11572 (N_11572,N_11070,N_11007);
and U11573 (N_11573,N_11401,N_11445);
xnor U11574 (N_11574,N_11098,N_11488);
xor U11575 (N_11575,N_11198,N_11019);
nor U11576 (N_11576,N_11323,N_11106);
nand U11577 (N_11577,N_11120,N_11409);
xnor U11578 (N_11578,N_11071,N_11341);
and U11579 (N_11579,N_11486,N_11324);
nand U11580 (N_11580,N_11261,N_11231);
xor U11581 (N_11581,N_11285,N_11186);
and U11582 (N_11582,N_11411,N_11320);
nand U11583 (N_11583,N_11085,N_11397);
xnor U11584 (N_11584,N_11073,N_11213);
and U11585 (N_11585,N_11372,N_11102);
xnor U11586 (N_11586,N_11030,N_11211);
nand U11587 (N_11587,N_11354,N_11478);
or U11588 (N_11588,N_11277,N_11135);
nand U11589 (N_11589,N_11218,N_11496);
or U11590 (N_11590,N_11064,N_11474);
and U11591 (N_11591,N_11069,N_11385);
nand U11592 (N_11592,N_11416,N_11113);
or U11593 (N_11593,N_11258,N_11487);
nand U11594 (N_11594,N_11310,N_11047);
or U11595 (N_11595,N_11221,N_11344);
xnor U11596 (N_11596,N_11222,N_11463);
nor U11597 (N_11597,N_11471,N_11470);
nand U11598 (N_11598,N_11379,N_11134);
or U11599 (N_11599,N_11387,N_11288);
and U11600 (N_11600,N_11432,N_11011);
nor U11601 (N_11601,N_11196,N_11024);
or U11602 (N_11602,N_11335,N_11154);
and U11603 (N_11603,N_11138,N_11205);
nand U11604 (N_11604,N_11462,N_11272);
xnor U11605 (N_11605,N_11415,N_11447);
nor U11606 (N_11606,N_11077,N_11398);
or U11607 (N_11607,N_11336,N_11190);
xnor U11608 (N_11608,N_11165,N_11189);
nand U11609 (N_11609,N_11431,N_11105);
or U11610 (N_11610,N_11150,N_11086);
and U11611 (N_11611,N_11349,N_11075);
or U11612 (N_11612,N_11167,N_11197);
xnor U11613 (N_11613,N_11237,N_11358);
xor U11614 (N_11614,N_11251,N_11300);
xor U11615 (N_11615,N_11101,N_11187);
xor U11616 (N_11616,N_11400,N_11125);
xnor U11617 (N_11617,N_11351,N_11407);
and U11618 (N_11618,N_11207,N_11052);
and U11619 (N_11619,N_11395,N_11157);
and U11620 (N_11620,N_11457,N_11266);
xnor U11621 (N_11621,N_11162,N_11228);
nand U11622 (N_11622,N_11321,N_11130);
nand U11623 (N_11623,N_11273,N_11356);
xor U11624 (N_11624,N_11095,N_11151);
and U11625 (N_11625,N_11023,N_11250);
or U11626 (N_11626,N_11216,N_11419);
nor U11627 (N_11627,N_11380,N_11027);
or U11628 (N_11628,N_11294,N_11424);
and U11629 (N_11629,N_11144,N_11133);
xnor U11630 (N_11630,N_11076,N_11078);
nand U11631 (N_11631,N_11260,N_11494);
xnor U11632 (N_11632,N_11410,N_11206);
xor U11633 (N_11633,N_11059,N_11399);
nor U11634 (N_11634,N_11034,N_11000);
nand U11635 (N_11635,N_11469,N_11422);
or U11636 (N_11636,N_11072,N_11122);
and U11637 (N_11637,N_11054,N_11292);
xor U11638 (N_11638,N_11365,N_11204);
or U11639 (N_11639,N_11223,N_11362);
nor U11640 (N_11640,N_11287,N_11046);
and U11641 (N_11641,N_11337,N_11386);
and U11642 (N_11642,N_11347,N_11089);
nand U11643 (N_11643,N_11453,N_11366);
nand U11644 (N_11644,N_11283,N_11238);
xor U11645 (N_11645,N_11212,N_11346);
xor U11646 (N_11646,N_11333,N_11170);
nand U11647 (N_11647,N_11191,N_11074);
or U11648 (N_11648,N_11353,N_11278);
or U11649 (N_11649,N_11303,N_11456);
nor U11650 (N_11650,N_11270,N_11343);
nor U11651 (N_11651,N_11008,N_11051);
nand U11652 (N_11652,N_11483,N_11021);
xnor U11653 (N_11653,N_11208,N_11438);
or U11654 (N_11654,N_11234,N_11326);
xnor U11655 (N_11655,N_11402,N_11139);
nand U11656 (N_11656,N_11036,N_11233);
or U11657 (N_11657,N_11434,N_11330);
nor U11658 (N_11658,N_11493,N_11220);
or U11659 (N_11659,N_11430,N_11327);
and U11660 (N_11660,N_11331,N_11068);
and U11661 (N_11661,N_11342,N_11219);
nand U11662 (N_11662,N_11200,N_11014);
nand U11663 (N_11663,N_11156,N_11334);
xnor U11664 (N_11664,N_11297,N_11177);
nor U11665 (N_11665,N_11429,N_11002);
xor U11666 (N_11666,N_11038,N_11053);
and U11667 (N_11667,N_11293,N_11180);
xor U11668 (N_11668,N_11239,N_11264);
and U11669 (N_11669,N_11465,N_11175);
nor U11670 (N_11670,N_11032,N_11378);
xnor U11671 (N_11671,N_11477,N_11296);
and U11672 (N_11672,N_11083,N_11371);
nand U11673 (N_11673,N_11193,N_11498);
xnor U11674 (N_11674,N_11009,N_11381);
xor U11675 (N_11675,N_11172,N_11230);
nor U11676 (N_11676,N_11375,N_11241);
xnor U11677 (N_11677,N_11100,N_11455);
and U11678 (N_11678,N_11136,N_11240);
nand U11679 (N_11679,N_11229,N_11338);
nor U11680 (N_11680,N_11420,N_11435);
and U11681 (N_11681,N_11029,N_11084);
and U11682 (N_11682,N_11359,N_11159);
or U11683 (N_11683,N_11490,N_11225);
nor U11684 (N_11684,N_11254,N_11152);
xor U11685 (N_11685,N_11145,N_11050);
and U11686 (N_11686,N_11020,N_11168);
and U11687 (N_11687,N_11081,N_11265);
nor U11688 (N_11688,N_11439,N_11479);
and U11689 (N_11689,N_11148,N_11040);
xor U11690 (N_11690,N_11124,N_11473);
and U11691 (N_11691,N_11373,N_11309);
nand U11692 (N_11692,N_11041,N_11348);
xnor U11693 (N_11693,N_11224,N_11126);
nand U11694 (N_11694,N_11115,N_11209);
and U11695 (N_11695,N_11382,N_11452);
nand U11696 (N_11696,N_11436,N_11491);
xnor U11697 (N_11697,N_11311,N_11448);
nor U11698 (N_11698,N_11361,N_11276);
nor U11699 (N_11699,N_11010,N_11042);
or U11700 (N_11700,N_11181,N_11067);
xor U11701 (N_11701,N_11192,N_11171);
and U11702 (N_11702,N_11414,N_11268);
nand U11703 (N_11703,N_11232,N_11253);
and U11704 (N_11704,N_11350,N_11256);
and U11705 (N_11705,N_11236,N_11280);
or U11706 (N_11706,N_11345,N_11269);
nor U11707 (N_11707,N_11460,N_11427);
or U11708 (N_11708,N_11289,N_11461);
and U11709 (N_11709,N_11096,N_11301);
and U11710 (N_11710,N_11164,N_11035);
and U11711 (N_11711,N_11295,N_11428);
and U11712 (N_11712,N_11099,N_11315);
xor U11713 (N_11713,N_11444,N_11132);
nor U11714 (N_11714,N_11235,N_11044);
nand U11715 (N_11715,N_11033,N_11282);
nand U11716 (N_11716,N_11055,N_11492);
nand U11717 (N_11717,N_11062,N_11279);
nand U11718 (N_11718,N_11318,N_11481);
nor U11719 (N_11719,N_11244,N_11119);
xnor U11720 (N_11720,N_11468,N_11079);
nor U11721 (N_11721,N_11376,N_11423);
xor U11722 (N_11722,N_11497,N_11015);
xor U11723 (N_11723,N_11405,N_11246);
nor U11724 (N_11724,N_11325,N_11451);
nor U11725 (N_11725,N_11464,N_11384);
nor U11726 (N_11726,N_11104,N_11202);
xnor U11727 (N_11727,N_11123,N_11173);
and U11728 (N_11728,N_11147,N_11367);
nand U11729 (N_11729,N_11443,N_11368);
nor U11730 (N_11730,N_11112,N_11396);
nand U11731 (N_11731,N_11412,N_11039);
nand U11732 (N_11732,N_11169,N_11087);
nor U11733 (N_11733,N_11454,N_11249);
and U11734 (N_11734,N_11195,N_11305);
nand U11735 (N_11735,N_11117,N_11066);
and U11736 (N_11736,N_11458,N_11174);
and U11737 (N_11737,N_11107,N_11006);
or U11738 (N_11738,N_11275,N_11286);
or U11739 (N_11739,N_11005,N_11109);
or U11740 (N_11740,N_11317,N_11267);
xnor U11741 (N_11741,N_11449,N_11043);
nor U11742 (N_11742,N_11031,N_11063);
and U11743 (N_11743,N_11406,N_11022);
xnor U11744 (N_11744,N_11357,N_11108);
nand U11745 (N_11745,N_11308,N_11088);
xnor U11746 (N_11746,N_11257,N_11319);
nand U11747 (N_11747,N_11476,N_11459);
nor U11748 (N_11748,N_11352,N_11166);
nor U11749 (N_11749,N_11307,N_11090);
xnor U11750 (N_11750,N_11258,N_11136);
and U11751 (N_11751,N_11110,N_11215);
nor U11752 (N_11752,N_11336,N_11039);
nand U11753 (N_11753,N_11258,N_11481);
or U11754 (N_11754,N_11166,N_11389);
xor U11755 (N_11755,N_11462,N_11103);
nor U11756 (N_11756,N_11283,N_11467);
xor U11757 (N_11757,N_11422,N_11262);
nor U11758 (N_11758,N_11077,N_11209);
xnor U11759 (N_11759,N_11124,N_11385);
or U11760 (N_11760,N_11247,N_11397);
and U11761 (N_11761,N_11374,N_11352);
xnor U11762 (N_11762,N_11286,N_11190);
and U11763 (N_11763,N_11289,N_11476);
xor U11764 (N_11764,N_11250,N_11173);
nor U11765 (N_11765,N_11184,N_11491);
nand U11766 (N_11766,N_11326,N_11351);
nand U11767 (N_11767,N_11278,N_11382);
nor U11768 (N_11768,N_11171,N_11228);
xor U11769 (N_11769,N_11007,N_11163);
and U11770 (N_11770,N_11179,N_11119);
xnor U11771 (N_11771,N_11234,N_11361);
xnor U11772 (N_11772,N_11149,N_11497);
or U11773 (N_11773,N_11412,N_11389);
xnor U11774 (N_11774,N_11013,N_11102);
nand U11775 (N_11775,N_11111,N_11161);
nor U11776 (N_11776,N_11379,N_11328);
and U11777 (N_11777,N_11067,N_11194);
and U11778 (N_11778,N_11246,N_11274);
xnor U11779 (N_11779,N_11106,N_11282);
nor U11780 (N_11780,N_11117,N_11049);
nor U11781 (N_11781,N_11272,N_11006);
and U11782 (N_11782,N_11424,N_11402);
xor U11783 (N_11783,N_11357,N_11403);
and U11784 (N_11784,N_11382,N_11342);
nand U11785 (N_11785,N_11119,N_11213);
or U11786 (N_11786,N_11042,N_11344);
nand U11787 (N_11787,N_11355,N_11484);
xor U11788 (N_11788,N_11024,N_11456);
nand U11789 (N_11789,N_11082,N_11177);
nand U11790 (N_11790,N_11122,N_11211);
nand U11791 (N_11791,N_11070,N_11028);
xnor U11792 (N_11792,N_11050,N_11475);
nor U11793 (N_11793,N_11215,N_11088);
or U11794 (N_11794,N_11181,N_11271);
or U11795 (N_11795,N_11204,N_11063);
xnor U11796 (N_11796,N_11009,N_11208);
nor U11797 (N_11797,N_11231,N_11331);
xor U11798 (N_11798,N_11002,N_11295);
or U11799 (N_11799,N_11497,N_11068);
or U11800 (N_11800,N_11401,N_11399);
and U11801 (N_11801,N_11119,N_11040);
nand U11802 (N_11802,N_11368,N_11238);
and U11803 (N_11803,N_11256,N_11145);
nand U11804 (N_11804,N_11034,N_11425);
nor U11805 (N_11805,N_11167,N_11481);
or U11806 (N_11806,N_11309,N_11124);
nor U11807 (N_11807,N_11244,N_11409);
nor U11808 (N_11808,N_11276,N_11286);
nand U11809 (N_11809,N_11047,N_11328);
or U11810 (N_11810,N_11029,N_11404);
nand U11811 (N_11811,N_11371,N_11491);
or U11812 (N_11812,N_11397,N_11478);
xor U11813 (N_11813,N_11342,N_11124);
or U11814 (N_11814,N_11078,N_11497);
and U11815 (N_11815,N_11087,N_11399);
and U11816 (N_11816,N_11189,N_11090);
nand U11817 (N_11817,N_11319,N_11079);
xor U11818 (N_11818,N_11380,N_11001);
nand U11819 (N_11819,N_11291,N_11410);
xnor U11820 (N_11820,N_11471,N_11293);
xor U11821 (N_11821,N_11017,N_11330);
nand U11822 (N_11822,N_11362,N_11439);
and U11823 (N_11823,N_11272,N_11050);
nand U11824 (N_11824,N_11106,N_11261);
nand U11825 (N_11825,N_11257,N_11265);
or U11826 (N_11826,N_11220,N_11321);
xnor U11827 (N_11827,N_11264,N_11262);
nor U11828 (N_11828,N_11292,N_11420);
and U11829 (N_11829,N_11021,N_11124);
and U11830 (N_11830,N_11366,N_11246);
nor U11831 (N_11831,N_11085,N_11079);
nor U11832 (N_11832,N_11224,N_11261);
and U11833 (N_11833,N_11306,N_11165);
or U11834 (N_11834,N_11332,N_11359);
nor U11835 (N_11835,N_11111,N_11397);
and U11836 (N_11836,N_11243,N_11409);
or U11837 (N_11837,N_11410,N_11368);
nand U11838 (N_11838,N_11146,N_11247);
nand U11839 (N_11839,N_11161,N_11176);
nor U11840 (N_11840,N_11421,N_11346);
nor U11841 (N_11841,N_11244,N_11495);
and U11842 (N_11842,N_11108,N_11074);
and U11843 (N_11843,N_11408,N_11146);
xor U11844 (N_11844,N_11323,N_11376);
or U11845 (N_11845,N_11046,N_11094);
xnor U11846 (N_11846,N_11067,N_11175);
nand U11847 (N_11847,N_11199,N_11226);
and U11848 (N_11848,N_11123,N_11071);
xor U11849 (N_11849,N_11403,N_11217);
xnor U11850 (N_11850,N_11462,N_11410);
nand U11851 (N_11851,N_11115,N_11402);
nor U11852 (N_11852,N_11100,N_11428);
nand U11853 (N_11853,N_11208,N_11112);
and U11854 (N_11854,N_11485,N_11057);
or U11855 (N_11855,N_11119,N_11450);
xnor U11856 (N_11856,N_11265,N_11102);
and U11857 (N_11857,N_11316,N_11321);
nand U11858 (N_11858,N_11141,N_11283);
nor U11859 (N_11859,N_11031,N_11025);
or U11860 (N_11860,N_11344,N_11441);
and U11861 (N_11861,N_11239,N_11284);
nor U11862 (N_11862,N_11482,N_11215);
nand U11863 (N_11863,N_11190,N_11264);
or U11864 (N_11864,N_11445,N_11369);
or U11865 (N_11865,N_11277,N_11249);
xor U11866 (N_11866,N_11262,N_11367);
or U11867 (N_11867,N_11363,N_11230);
xor U11868 (N_11868,N_11018,N_11168);
and U11869 (N_11869,N_11289,N_11470);
xor U11870 (N_11870,N_11223,N_11179);
nor U11871 (N_11871,N_11387,N_11035);
and U11872 (N_11872,N_11007,N_11039);
or U11873 (N_11873,N_11004,N_11448);
nand U11874 (N_11874,N_11065,N_11062);
or U11875 (N_11875,N_11167,N_11196);
xnor U11876 (N_11876,N_11369,N_11116);
xor U11877 (N_11877,N_11465,N_11498);
or U11878 (N_11878,N_11199,N_11329);
or U11879 (N_11879,N_11095,N_11060);
nor U11880 (N_11880,N_11211,N_11032);
or U11881 (N_11881,N_11454,N_11004);
nand U11882 (N_11882,N_11150,N_11201);
nand U11883 (N_11883,N_11191,N_11416);
or U11884 (N_11884,N_11411,N_11212);
or U11885 (N_11885,N_11436,N_11112);
nor U11886 (N_11886,N_11028,N_11195);
nor U11887 (N_11887,N_11037,N_11231);
xnor U11888 (N_11888,N_11075,N_11182);
nand U11889 (N_11889,N_11368,N_11096);
nor U11890 (N_11890,N_11345,N_11148);
nand U11891 (N_11891,N_11270,N_11085);
and U11892 (N_11892,N_11435,N_11106);
nand U11893 (N_11893,N_11358,N_11372);
nor U11894 (N_11894,N_11188,N_11021);
xnor U11895 (N_11895,N_11364,N_11012);
xor U11896 (N_11896,N_11234,N_11446);
nor U11897 (N_11897,N_11365,N_11352);
xor U11898 (N_11898,N_11356,N_11396);
or U11899 (N_11899,N_11400,N_11017);
and U11900 (N_11900,N_11074,N_11411);
xnor U11901 (N_11901,N_11233,N_11348);
and U11902 (N_11902,N_11151,N_11174);
xor U11903 (N_11903,N_11392,N_11243);
nand U11904 (N_11904,N_11156,N_11070);
xnor U11905 (N_11905,N_11212,N_11431);
nor U11906 (N_11906,N_11165,N_11382);
xnor U11907 (N_11907,N_11405,N_11268);
and U11908 (N_11908,N_11331,N_11304);
xor U11909 (N_11909,N_11455,N_11434);
and U11910 (N_11910,N_11158,N_11202);
nand U11911 (N_11911,N_11075,N_11137);
nand U11912 (N_11912,N_11022,N_11145);
and U11913 (N_11913,N_11051,N_11404);
nor U11914 (N_11914,N_11085,N_11281);
and U11915 (N_11915,N_11060,N_11075);
nand U11916 (N_11916,N_11472,N_11333);
or U11917 (N_11917,N_11264,N_11165);
and U11918 (N_11918,N_11445,N_11101);
and U11919 (N_11919,N_11074,N_11166);
nand U11920 (N_11920,N_11134,N_11492);
nand U11921 (N_11921,N_11473,N_11237);
nor U11922 (N_11922,N_11452,N_11003);
or U11923 (N_11923,N_11136,N_11135);
and U11924 (N_11924,N_11416,N_11132);
or U11925 (N_11925,N_11387,N_11080);
or U11926 (N_11926,N_11005,N_11063);
and U11927 (N_11927,N_11115,N_11316);
xnor U11928 (N_11928,N_11263,N_11138);
and U11929 (N_11929,N_11112,N_11100);
nor U11930 (N_11930,N_11194,N_11426);
nor U11931 (N_11931,N_11340,N_11140);
xor U11932 (N_11932,N_11271,N_11458);
and U11933 (N_11933,N_11241,N_11408);
nand U11934 (N_11934,N_11317,N_11025);
or U11935 (N_11935,N_11004,N_11254);
nor U11936 (N_11936,N_11246,N_11463);
or U11937 (N_11937,N_11291,N_11364);
nand U11938 (N_11938,N_11007,N_11457);
xnor U11939 (N_11939,N_11060,N_11143);
and U11940 (N_11940,N_11353,N_11101);
xor U11941 (N_11941,N_11429,N_11361);
and U11942 (N_11942,N_11332,N_11448);
xnor U11943 (N_11943,N_11452,N_11320);
or U11944 (N_11944,N_11084,N_11039);
nand U11945 (N_11945,N_11133,N_11022);
and U11946 (N_11946,N_11006,N_11062);
or U11947 (N_11947,N_11003,N_11393);
nand U11948 (N_11948,N_11116,N_11496);
nor U11949 (N_11949,N_11208,N_11161);
xor U11950 (N_11950,N_11246,N_11191);
or U11951 (N_11951,N_11446,N_11066);
and U11952 (N_11952,N_11070,N_11423);
nor U11953 (N_11953,N_11305,N_11264);
and U11954 (N_11954,N_11134,N_11062);
nand U11955 (N_11955,N_11447,N_11358);
xor U11956 (N_11956,N_11098,N_11282);
xor U11957 (N_11957,N_11376,N_11146);
xnor U11958 (N_11958,N_11333,N_11283);
and U11959 (N_11959,N_11018,N_11333);
or U11960 (N_11960,N_11176,N_11069);
xor U11961 (N_11961,N_11110,N_11489);
or U11962 (N_11962,N_11496,N_11282);
nor U11963 (N_11963,N_11206,N_11207);
nand U11964 (N_11964,N_11062,N_11219);
nor U11965 (N_11965,N_11333,N_11084);
and U11966 (N_11966,N_11045,N_11340);
nor U11967 (N_11967,N_11008,N_11077);
nor U11968 (N_11968,N_11275,N_11405);
and U11969 (N_11969,N_11178,N_11086);
nand U11970 (N_11970,N_11435,N_11281);
nor U11971 (N_11971,N_11195,N_11351);
xor U11972 (N_11972,N_11335,N_11165);
or U11973 (N_11973,N_11123,N_11024);
and U11974 (N_11974,N_11072,N_11110);
nor U11975 (N_11975,N_11130,N_11404);
and U11976 (N_11976,N_11319,N_11228);
nor U11977 (N_11977,N_11209,N_11375);
nand U11978 (N_11978,N_11099,N_11305);
or U11979 (N_11979,N_11424,N_11327);
xnor U11980 (N_11980,N_11380,N_11127);
nand U11981 (N_11981,N_11395,N_11269);
and U11982 (N_11982,N_11010,N_11369);
or U11983 (N_11983,N_11141,N_11388);
nand U11984 (N_11984,N_11105,N_11133);
xnor U11985 (N_11985,N_11468,N_11298);
nor U11986 (N_11986,N_11224,N_11039);
or U11987 (N_11987,N_11138,N_11492);
xnor U11988 (N_11988,N_11418,N_11205);
or U11989 (N_11989,N_11238,N_11159);
xnor U11990 (N_11990,N_11451,N_11415);
nand U11991 (N_11991,N_11248,N_11414);
nor U11992 (N_11992,N_11297,N_11154);
or U11993 (N_11993,N_11004,N_11346);
or U11994 (N_11994,N_11414,N_11004);
or U11995 (N_11995,N_11139,N_11047);
nor U11996 (N_11996,N_11083,N_11476);
or U11997 (N_11997,N_11033,N_11247);
nand U11998 (N_11998,N_11012,N_11330);
or U11999 (N_11999,N_11443,N_11230);
nand U12000 (N_12000,N_11754,N_11991);
xnor U12001 (N_12001,N_11997,N_11785);
nor U12002 (N_12002,N_11981,N_11564);
nor U12003 (N_12003,N_11512,N_11670);
xnor U12004 (N_12004,N_11976,N_11777);
or U12005 (N_12005,N_11745,N_11518);
and U12006 (N_12006,N_11787,N_11811);
and U12007 (N_12007,N_11943,N_11590);
nand U12008 (N_12008,N_11611,N_11626);
nor U12009 (N_12009,N_11729,N_11678);
nor U12010 (N_12010,N_11555,N_11772);
nor U12011 (N_12011,N_11990,N_11524);
nor U12012 (N_12012,N_11685,N_11683);
and U12013 (N_12013,N_11520,N_11834);
nor U12014 (N_12014,N_11816,N_11868);
or U12015 (N_12015,N_11610,N_11743);
nand U12016 (N_12016,N_11882,N_11750);
or U12017 (N_12017,N_11582,N_11917);
nor U12018 (N_12018,N_11533,N_11881);
nand U12019 (N_12019,N_11936,N_11778);
xor U12020 (N_12020,N_11986,N_11843);
nand U12021 (N_12021,N_11988,N_11738);
or U12022 (N_12022,N_11856,N_11660);
nor U12023 (N_12023,N_11783,N_11607);
nor U12024 (N_12024,N_11562,N_11871);
or U12025 (N_12025,N_11643,N_11874);
or U12026 (N_12026,N_11515,N_11539);
xor U12027 (N_12027,N_11961,N_11715);
xor U12028 (N_12028,N_11673,N_11503);
nor U12029 (N_12029,N_11691,N_11613);
nand U12030 (N_12030,N_11795,N_11711);
nand U12031 (N_12031,N_11937,N_11975);
and U12032 (N_12032,N_11773,N_11846);
and U12033 (N_12033,N_11940,N_11526);
and U12034 (N_12034,N_11665,N_11629);
nand U12035 (N_12035,N_11823,N_11575);
and U12036 (N_12036,N_11807,N_11726);
nand U12037 (N_12037,N_11813,N_11977);
nor U12038 (N_12038,N_11779,N_11775);
or U12039 (N_12039,N_11657,N_11585);
nand U12040 (N_12040,N_11935,N_11630);
xor U12041 (N_12041,N_11609,N_11593);
and U12042 (N_12042,N_11719,N_11722);
or U12043 (N_12043,N_11752,N_11573);
nand U12044 (N_12044,N_11956,N_11648);
nand U12045 (N_12045,N_11644,N_11909);
nand U12046 (N_12046,N_11634,N_11727);
nand U12047 (N_12047,N_11734,N_11764);
and U12048 (N_12048,N_11746,N_11616);
xor U12049 (N_12049,N_11747,N_11650);
xor U12050 (N_12050,N_11840,N_11911);
and U12051 (N_12051,N_11788,N_11791);
nand U12052 (N_12052,N_11805,N_11511);
or U12053 (N_12053,N_11501,N_11681);
xnor U12054 (N_12054,N_11700,N_11675);
nand U12055 (N_12055,N_11867,N_11989);
or U12056 (N_12056,N_11951,N_11896);
xnor U12057 (N_12057,N_11725,N_11632);
and U12058 (N_12058,N_11680,N_11712);
xnor U12059 (N_12059,N_11748,N_11706);
xor U12060 (N_12060,N_11869,N_11589);
and U12061 (N_12061,N_11994,N_11864);
xnor U12062 (N_12062,N_11568,N_11821);
and U12063 (N_12063,N_11849,N_11510);
or U12064 (N_12064,N_11853,N_11567);
xnor U12065 (N_12065,N_11649,N_11766);
or U12066 (N_12066,N_11705,N_11699);
or U12067 (N_12067,N_11931,N_11693);
or U12068 (N_12068,N_11504,N_11969);
and U12069 (N_12069,N_11857,N_11525);
xnor U12070 (N_12070,N_11659,N_11891);
nor U12071 (N_12071,N_11591,N_11944);
and U12072 (N_12072,N_11808,N_11702);
nand U12073 (N_12073,N_11756,N_11838);
nor U12074 (N_12074,N_11854,N_11605);
or U12075 (N_12075,N_11963,N_11519);
nand U12076 (N_12076,N_11862,N_11652);
or U12077 (N_12077,N_11641,N_11737);
and U12078 (N_12078,N_11790,N_11530);
or U12079 (N_12079,N_11875,N_11627);
nand U12080 (N_12080,N_11762,N_11887);
nand U12081 (N_12081,N_11651,N_11910);
nor U12082 (N_12082,N_11758,N_11946);
nand U12083 (N_12083,N_11529,N_11916);
nand U12084 (N_12084,N_11588,N_11701);
xnor U12085 (N_12085,N_11947,N_11730);
or U12086 (N_12086,N_11508,N_11930);
xor U12087 (N_12087,N_11604,N_11755);
xnor U12088 (N_12088,N_11522,N_11866);
or U12089 (N_12089,N_11802,N_11962);
xnor U12090 (N_12090,N_11682,N_11577);
nand U12091 (N_12091,N_11537,N_11674);
and U12092 (N_12092,N_11985,N_11970);
nand U12093 (N_12093,N_11538,N_11662);
xnor U12094 (N_12094,N_11572,N_11560);
and U12095 (N_12095,N_11804,N_11833);
xor U12096 (N_12096,N_11559,N_11635);
nand U12097 (N_12097,N_11602,N_11718);
or U12098 (N_12098,N_11561,N_11847);
xor U12099 (N_12099,N_11516,N_11580);
nor U12100 (N_12100,N_11806,N_11809);
and U12101 (N_12101,N_11797,N_11586);
or U12102 (N_12102,N_11993,N_11850);
or U12103 (N_12103,N_11599,N_11959);
and U12104 (N_12104,N_11724,N_11579);
or U12105 (N_12105,N_11631,N_11713);
xor U12106 (N_12106,N_11556,N_11995);
nor U12107 (N_12107,N_11566,N_11897);
nor U12108 (N_12108,N_11733,N_11922);
nor U12109 (N_12109,N_11848,N_11984);
or U12110 (N_12110,N_11927,N_11603);
nor U12111 (N_12111,N_11886,N_11957);
nor U12112 (N_12112,N_11625,N_11780);
and U12113 (N_12113,N_11983,N_11655);
and U12114 (N_12114,N_11782,N_11873);
nor U12115 (N_12115,N_11633,N_11967);
or U12116 (N_12116,N_11606,N_11776);
and U12117 (N_12117,N_11812,N_11664);
nor U12118 (N_12118,N_11831,N_11953);
and U12119 (N_12119,N_11569,N_11661);
nor U12120 (N_12120,N_11803,N_11528);
xor U12121 (N_12121,N_11717,N_11624);
nand U12122 (N_12122,N_11842,N_11669);
and U12123 (N_12123,N_11926,N_11689);
or U12124 (N_12124,N_11679,N_11945);
nor U12125 (N_12125,N_11958,N_11587);
nand U12126 (N_12126,N_11794,N_11837);
nor U12127 (N_12127,N_11571,N_11768);
and U12128 (N_12128,N_11878,N_11894);
nand U12129 (N_12129,N_11551,N_11974);
and U12130 (N_12130,N_11570,N_11690);
xor U12131 (N_12131,N_11732,N_11647);
and U12132 (N_12132,N_11547,N_11941);
and U12133 (N_12133,N_11924,N_11858);
xnor U12134 (N_12134,N_11541,N_11980);
and U12135 (N_12135,N_11565,N_11949);
and U12136 (N_12136,N_11720,N_11545);
or U12137 (N_12137,N_11999,N_11709);
xor U12138 (N_12138,N_11832,N_11968);
and U12139 (N_12139,N_11902,N_11623);
and U12140 (N_12140,N_11898,N_11751);
and U12141 (N_12141,N_11932,N_11596);
or U12142 (N_12142,N_11656,N_11513);
and U12143 (N_12143,N_11905,N_11904);
or U12144 (N_12144,N_11908,N_11550);
and U12145 (N_12145,N_11663,N_11505);
or U12146 (N_12146,N_11695,N_11535);
and U12147 (N_12147,N_11915,N_11948);
and U12148 (N_12148,N_11861,N_11880);
nand U12149 (N_12149,N_11827,N_11507);
nand U12150 (N_12150,N_11741,N_11899);
nand U12151 (N_12151,N_11865,N_11761);
and U12152 (N_12152,N_11536,N_11696);
and U12153 (N_12153,N_11594,N_11760);
nand U12154 (N_12154,N_11870,N_11893);
and U12155 (N_12155,N_11584,N_11933);
xnor U12156 (N_12156,N_11578,N_11598);
nand U12157 (N_12157,N_11548,N_11820);
and U12158 (N_12158,N_11697,N_11676);
xor U12159 (N_12159,N_11771,N_11500);
and U12160 (N_12160,N_11987,N_11892);
nand U12161 (N_12161,N_11703,N_11671);
nor U12162 (N_12162,N_11714,N_11636);
and U12163 (N_12163,N_11825,N_11534);
and U12164 (N_12164,N_11774,N_11694);
nor U12165 (N_12165,N_11792,N_11549);
nand U12166 (N_12166,N_11757,N_11934);
xor U12167 (N_12167,N_11913,N_11998);
xnor U12168 (N_12168,N_11814,N_11759);
xor U12169 (N_12169,N_11723,N_11799);
nor U12170 (N_12170,N_11620,N_11742);
nand U12171 (N_12171,N_11521,N_11971);
xor U12172 (N_12172,N_11841,N_11639);
or U12173 (N_12173,N_11844,N_11769);
xnor U12174 (N_12174,N_11828,N_11531);
nand U12175 (N_12175,N_11698,N_11923);
and U12176 (N_12176,N_11736,N_11770);
and U12177 (N_12177,N_11688,N_11686);
and U12178 (N_12178,N_11744,N_11890);
nor U12179 (N_12179,N_11879,N_11996);
xor U12180 (N_12180,N_11637,N_11982);
or U12181 (N_12181,N_11563,N_11860);
xor U12182 (N_12182,N_11900,N_11684);
or U12183 (N_12183,N_11514,N_11667);
xnor U12184 (N_12184,N_11830,N_11654);
nand U12185 (N_12185,N_11824,N_11796);
or U12186 (N_12186,N_11835,N_11704);
xnor U12187 (N_12187,N_11979,N_11658);
nor U12188 (N_12188,N_11731,N_11852);
and U12189 (N_12189,N_11966,N_11544);
nor U12190 (N_12190,N_11557,N_11542);
xor U12191 (N_12191,N_11653,N_11716);
nand U12192 (N_12192,N_11540,N_11888);
and U12193 (N_12193,N_11640,N_11954);
nor U12194 (N_12194,N_11558,N_11789);
xor U12195 (N_12195,N_11928,N_11919);
nand U12196 (N_12196,N_11884,N_11749);
and U12197 (N_12197,N_11920,N_11527);
nand U12198 (N_12198,N_11576,N_11964);
nor U12199 (N_12199,N_11883,N_11543);
xor U12200 (N_12200,N_11517,N_11885);
and U12201 (N_12201,N_11597,N_11960);
or U12202 (N_12202,N_11642,N_11581);
nand U12203 (N_12203,N_11595,N_11786);
nor U12204 (N_12204,N_11767,N_11784);
xor U12205 (N_12205,N_11687,N_11906);
xor U12206 (N_12206,N_11622,N_11921);
or U12207 (N_12207,N_11739,N_11826);
and U12208 (N_12208,N_11592,N_11895);
nand U12209 (N_12209,N_11618,N_11829);
or U12210 (N_12210,N_11818,N_11950);
and U12211 (N_12211,N_11646,N_11800);
xnor U12212 (N_12212,N_11668,N_11583);
nand U12213 (N_12213,N_11973,N_11863);
nor U12214 (N_12214,N_11612,N_11692);
xnor U12215 (N_12215,N_11672,N_11628);
nand U12216 (N_12216,N_11872,N_11608);
xnor U12217 (N_12217,N_11901,N_11877);
nand U12218 (N_12218,N_11876,N_11810);
xnor U12219 (N_12219,N_11819,N_11532);
and U12220 (N_12220,N_11710,N_11666);
nand U12221 (N_12221,N_11942,N_11506);
xnor U12222 (N_12222,N_11855,N_11793);
or U12223 (N_12223,N_11822,N_11753);
nor U12224 (N_12224,N_11600,N_11801);
and U12225 (N_12225,N_11638,N_11546);
nor U12226 (N_12226,N_11938,N_11972);
or U12227 (N_12227,N_11836,N_11845);
nand U12228 (N_12228,N_11552,N_11817);
and U12229 (N_12229,N_11907,N_11955);
xnor U12230 (N_12230,N_11708,N_11992);
nand U12231 (N_12231,N_11574,N_11735);
nand U12232 (N_12232,N_11965,N_11617);
or U12233 (N_12233,N_11601,N_11614);
nor U12234 (N_12234,N_11925,N_11952);
and U12235 (N_12235,N_11765,N_11815);
or U12236 (N_12236,N_11645,N_11621);
nand U12237 (N_12237,N_11914,N_11859);
or U12238 (N_12238,N_11839,N_11523);
nor U12239 (N_12239,N_11918,N_11554);
nand U12240 (N_12240,N_11502,N_11677);
and U12241 (N_12241,N_11798,N_11939);
xor U12242 (N_12242,N_11615,N_11553);
or U12243 (N_12243,N_11912,N_11721);
and U12244 (N_12244,N_11728,N_11781);
or U12245 (N_12245,N_11978,N_11707);
nand U12246 (N_12246,N_11929,N_11851);
or U12247 (N_12247,N_11619,N_11740);
nor U12248 (N_12248,N_11889,N_11903);
or U12249 (N_12249,N_11509,N_11763);
nand U12250 (N_12250,N_11608,N_11972);
nor U12251 (N_12251,N_11523,N_11617);
or U12252 (N_12252,N_11664,N_11546);
and U12253 (N_12253,N_11622,N_11646);
and U12254 (N_12254,N_11975,N_11888);
xor U12255 (N_12255,N_11733,N_11939);
nor U12256 (N_12256,N_11905,N_11992);
nor U12257 (N_12257,N_11578,N_11601);
or U12258 (N_12258,N_11541,N_11644);
xnor U12259 (N_12259,N_11951,N_11644);
or U12260 (N_12260,N_11650,N_11903);
and U12261 (N_12261,N_11877,N_11501);
or U12262 (N_12262,N_11696,N_11855);
xor U12263 (N_12263,N_11509,N_11539);
and U12264 (N_12264,N_11637,N_11962);
and U12265 (N_12265,N_11647,N_11625);
nand U12266 (N_12266,N_11825,N_11971);
xnor U12267 (N_12267,N_11670,N_11600);
nand U12268 (N_12268,N_11818,N_11965);
nand U12269 (N_12269,N_11855,N_11618);
nand U12270 (N_12270,N_11514,N_11518);
and U12271 (N_12271,N_11961,N_11775);
nand U12272 (N_12272,N_11635,N_11861);
or U12273 (N_12273,N_11979,N_11681);
nand U12274 (N_12274,N_11858,N_11770);
nand U12275 (N_12275,N_11714,N_11912);
nand U12276 (N_12276,N_11654,N_11694);
nand U12277 (N_12277,N_11915,N_11634);
and U12278 (N_12278,N_11970,N_11672);
or U12279 (N_12279,N_11980,N_11601);
and U12280 (N_12280,N_11513,N_11603);
nand U12281 (N_12281,N_11658,N_11626);
xor U12282 (N_12282,N_11857,N_11664);
and U12283 (N_12283,N_11726,N_11868);
or U12284 (N_12284,N_11558,N_11799);
xor U12285 (N_12285,N_11986,N_11619);
xnor U12286 (N_12286,N_11876,N_11940);
xor U12287 (N_12287,N_11875,N_11748);
nand U12288 (N_12288,N_11982,N_11839);
xnor U12289 (N_12289,N_11921,N_11801);
xor U12290 (N_12290,N_11702,N_11872);
and U12291 (N_12291,N_11600,N_11697);
or U12292 (N_12292,N_11591,N_11850);
xor U12293 (N_12293,N_11901,N_11957);
nand U12294 (N_12294,N_11666,N_11651);
nand U12295 (N_12295,N_11859,N_11641);
nor U12296 (N_12296,N_11857,N_11757);
xnor U12297 (N_12297,N_11630,N_11544);
nand U12298 (N_12298,N_11919,N_11792);
nand U12299 (N_12299,N_11664,N_11609);
nor U12300 (N_12300,N_11914,N_11582);
nand U12301 (N_12301,N_11753,N_11772);
nor U12302 (N_12302,N_11622,N_11579);
nor U12303 (N_12303,N_11692,N_11735);
and U12304 (N_12304,N_11998,N_11787);
nor U12305 (N_12305,N_11913,N_11719);
nor U12306 (N_12306,N_11680,N_11951);
and U12307 (N_12307,N_11987,N_11675);
and U12308 (N_12308,N_11873,N_11999);
or U12309 (N_12309,N_11523,N_11805);
xor U12310 (N_12310,N_11706,N_11583);
nand U12311 (N_12311,N_11718,N_11613);
and U12312 (N_12312,N_11561,N_11740);
and U12313 (N_12313,N_11551,N_11824);
nor U12314 (N_12314,N_11964,N_11867);
or U12315 (N_12315,N_11524,N_11639);
or U12316 (N_12316,N_11800,N_11911);
nand U12317 (N_12317,N_11585,N_11862);
or U12318 (N_12318,N_11836,N_11799);
nand U12319 (N_12319,N_11648,N_11713);
nand U12320 (N_12320,N_11531,N_11971);
nand U12321 (N_12321,N_11981,N_11548);
xor U12322 (N_12322,N_11793,N_11871);
or U12323 (N_12323,N_11635,N_11774);
or U12324 (N_12324,N_11770,N_11781);
nand U12325 (N_12325,N_11941,N_11720);
xnor U12326 (N_12326,N_11840,N_11522);
xor U12327 (N_12327,N_11657,N_11714);
and U12328 (N_12328,N_11799,N_11707);
or U12329 (N_12329,N_11974,N_11858);
nor U12330 (N_12330,N_11586,N_11847);
nand U12331 (N_12331,N_11922,N_11616);
and U12332 (N_12332,N_11689,N_11632);
xnor U12333 (N_12333,N_11656,N_11614);
nor U12334 (N_12334,N_11769,N_11523);
nand U12335 (N_12335,N_11568,N_11576);
nor U12336 (N_12336,N_11743,N_11949);
nand U12337 (N_12337,N_11535,N_11807);
xor U12338 (N_12338,N_11544,N_11987);
or U12339 (N_12339,N_11970,N_11976);
nand U12340 (N_12340,N_11550,N_11515);
nor U12341 (N_12341,N_11508,N_11699);
nor U12342 (N_12342,N_11556,N_11885);
nand U12343 (N_12343,N_11883,N_11845);
and U12344 (N_12344,N_11886,N_11652);
or U12345 (N_12345,N_11833,N_11818);
or U12346 (N_12346,N_11678,N_11782);
and U12347 (N_12347,N_11982,N_11866);
nor U12348 (N_12348,N_11571,N_11828);
xor U12349 (N_12349,N_11534,N_11562);
or U12350 (N_12350,N_11777,N_11667);
xor U12351 (N_12351,N_11503,N_11856);
xor U12352 (N_12352,N_11911,N_11885);
nor U12353 (N_12353,N_11687,N_11994);
and U12354 (N_12354,N_11690,N_11935);
nand U12355 (N_12355,N_11604,N_11739);
xor U12356 (N_12356,N_11658,N_11716);
or U12357 (N_12357,N_11641,N_11693);
and U12358 (N_12358,N_11625,N_11622);
or U12359 (N_12359,N_11786,N_11765);
nand U12360 (N_12360,N_11729,N_11565);
or U12361 (N_12361,N_11637,N_11665);
nand U12362 (N_12362,N_11943,N_11910);
nand U12363 (N_12363,N_11724,N_11742);
and U12364 (N_12364,N_11537,N_11784);
xor U12365 (N_12365,N_11773,N_11512);
xor U12366 (N_12366,N_11939,N_11620);
xnor U12367 (N_12367,N_11529,N_11545);
nand U12368 (N_12368,N_11672,N_11539);
nand U12369 (N_12369,N_11628,N_11890);
xnor U12370 (N_12370,N_11886,N_11646);
or U12371 (N_12371,N_11628,N_11924);
or U12372 (N_12372,N_11710,N_11739);
nand U12373 (N_12373,N_11890,N_11769);
nand U12374 (N_12374,N_11876,N_11928);
nand U12375 (N_12375,N_11686,N_11826);
xor U12376 (N_12376,N_11644,N_11764);
nor U12377 (N_12377,N_11604,N_11717);
xnor U12378 (N_12378,N_11784,N_11936);
nor U12379 (N_12379,N_11973,N_11587);
nand U12380 (N_12380,N_11963,N_11822);
and U12381 (N_12381,N_11744,N_11824);
or U12382 (N_12382,N_11536,N_11581);
nor U12383 (N_12383,N_11635,N_11965);
xor U12384 (N_12384,N_11816,N_11657);
nor U12385 (N_12385,N_11849,N_11993);
and U12386 (N_12386,N_11500,N_11840);
nand U12387 (N_12387,N_11917,N_11795);
nand U12388 (N_12388,N_11646,N_11802);
and U12389 (N_12389,N_11600,N_11703);
and U12390 (N_12390,N_11891,N_11953);
nand U12391 (N_12391,N_11550,N_11507);
nand U12392 (N_12392,N_11658,N_11613);
xnor U12393 (N_12393,N_11816,N_11846);
nand U12394 (N_12394,N_11566,N_11812);
and U12395 (N_12395,N_11697,N_11558);
and U12396 (N_12396,N_11605,N_11533);
and U12397 (N_12397,N_11641,N_11789);
nand U12398 (N_12398,N_11925,N_11885);
or U12399 (N_12399,N_11782,N_11975);
and U12400 (N_12400,N_11600,N_11756);
xnor U12401 (N_12401,N_11830,N_11761);
and U12402 (N_12402,N_11884,N_11830);
nor U12403 (N_12403,N_11789,N_11918);
or U12404 (N_12404,N_11923,N_11808);
nor U12405 (N_12405,N_11736,N_11633);
nand U12406 (N_12406,N_11566,N_11608);
xor U12407 (N_12407,N_11524,N_11607);
xnor U12408 (N_12408,N_11570,N_11695);
nand U12409 (N_12409,N_11644,N_11700);
nor U12410 (N_12410,N_11897,N_11899);
xor U12411 (N_12411,N_11869,N_11805);
or U12412 (N_12412,N_11505,N_11728);
xnor U12413 (N_12413,N_11513,N_11700);
nand U12414 (N_12414,N_11941,N_11571);
or U12415 (N_12415,N_11535,N_11522);
or U12416 (N_12416,N_11796,N_11615);
nor U12417 (N_12417,N_11981,N_11688);
nand U12418 (N_12418,N_11581,N_11631);
nor U12419 (N_12419,N_11759,N_11780);
and U12420 (N_12420,N_11631,N_11628);
nand U12421 (N_12421,N_11717,N_11817);
xor U12422 (N_12422,N_11639,N_11902);
xor U12423 (N_12423,N_11579,N_11810);
or U12424 (N_12424,N_11638,N_11587);
nor U12425 (N_12425,N_11807,N_11840);
or U12426 (N_12426,N_11834,N_11642);
xor U12427 (N_12427,N_11821,N_11998);
nor U12428 (N_12428,N_11703,N_11824);
and U12429 (N_12429,N_11973,N_11935);
xnor U12430 (N_12430,N_11966,N_11748);
and U12431 (N_12431,N_11871,N_11600);
or U12432 (N_12432,N_11635,N_11517);
nor U12433 (N_12433,N_11956,N_11754);
nand U12434 (N_12434,N_11713,N_11634);
nor U12435 (N_12435,N_11865,N_11601);
and U12436 (N_12436,N_11864,N_11783);
nand U12437 (N_12437,N_11732,N_11556);
or U12438 (N_12438,N_11881,N_11678);
nand U12439 (N_12439,N_11966,N_11514);
or U12440 (N_12440,N_11551,N_11687);
xnor U12441 (N_12441,N_11934,N_11587);
and U12442 (N_12442,N_11575,N_11664);
nor U12443 (N_12443,N_11611,N_11628);
xnor U12444 (N_12444,N_11884,N_11997);
xnor U12445 (N_12445,N_11797,N_11789);
or U12446 (N_12446,N_11605,N_11630);
and U12447 (N_12447,N_11545,N_11657);
and U12448 (N_12448,N_11953,N_11707);
xor U12449 (N_12449,N_11936,N_11630);
or U12450 (N_12450,N_11725,N_11654);
nand U12451 (N_12451,N_11599,N_11915);
and U12452 (N_12452,N_11935,N_11701);
xnor U12453 (N_12453,N_11514,N_11564);
and U12454 (N_12454,N_11997,N_11515);
nor U12455 (N_12455,N_11646,N_11694);
or U12456 (N_12456,N_11796,N_11806);
or U12457 (N_12457,N_11808,N_11701);
nand U12458 (N_12458,N_11961,N_11601);
nand U12459 (N_12459,N_11838,N_11996);
or U12460 (N_12460,N_11824,N_11889);
or U12461 (N_12461,N_11821,N_11806);
nor U12462 (N_12462,N_11796,N_11803);
nand U12463 (N_12463,N_11704,N_11607);
nor U12464 (N_12464,N_11624,N_11544);
and U12465 (N_12465,N_11760,N_11596);
and U12466 (N_12466,N_11998,N_11878);
xor U12467 (N_12467,N_11956,N_11895);
and U12468 (N_12468,N_11526,N_11948);
or U12469 (N_12469,N_11692,N_11508);
nor U12470 (N_12470,N_11666,N_11703);
or U12471 (N_12471,N_11996,N_11610);
nand U12472 (N_12472,N_11651,N_11526);
nor U12473 (N_12473,N_11993,N_11605);
or U12474 (N_12474,N_11775,N_11803);
nand U12475 (N_12475,N_11802,N_11677);
xnor U12476 (N_12476,N_11735,N_11914);
nand U12477 (N_12477,N_11836,N_11760);
nand U12478 (N_12478,N_11882,N_11851);
xnor U12479 (N_12479,N_11960,N_11992);
xnor U12480 (N_12480,N_11976,N_11841);
nor U12481 (N_12481,N_11870,N_11988);
xnor U12482 (N_12482,N_11761,N_11740);
or U12483 (N_12483,N_11615,N_11704);
nor U12484 (N_12484,N_11791,N_11853);
and U12485 (N_12485,N_11684,N_11775);
nand U12486 (N_12486,N_11862,N_11852);
or U12487 (N_12487,N_11524,N_11901);
and U12488 (N_12488,N_11942,N_11586);
nand U12489 (N_12489,N_11591,N_11537);
nand U12490 (N_12490,N_11744,N_11796);
xor U12491 (N_12491,N_11902,N_11565);
nand U12492 (N_12492,N_11978,N_11688);
or U12493 (N_12493,N_11837,N_11867);
or U12494 (N_12494,N_11758,N_11568);
nand U12495 (N_12495,N_11566,N_11816);
xnor U12496 (N_12496,N_11797,N_11792);
or U12497 (N_12497,N_11581,N_11724);
or U12498 (N_12498,N_11738,N_11755);
xor U12499 (N_12499,N_11750,N_11795);
or U12500 (N_12500,N_12072,N_12481);
and U12501 (N_12501,N_12265,N_12381);
xor U12502 (N_12502,N_12200,N_12147);
nor U12503 (N_12503,N_12492,N_12003);
and U12504 (N_12504,N_12386,N_12294);
nor U12505 (N_12505,N_12301,N_12292);
xor U12506 (N_12506,N_12393,N_12367);
nor U12507 (N_12507,N_12279,N_12220);
nor U12508 (N_12508,N_12010,N_12176);
nor U12509 (N_12509,N_12373,N_12196);
xnor U12510 (N_12510,N_12051,N_12026);
xor U12511 (N_12511,N_12322,N_12224);
or U12512 (N_12512,N_12420,N_12160);
or U12513 (N_12513,N_12483,N_12319);
or U12514 (N_12514,N_12317,N_12298);
and U12515 (N_12515,N_12474,N_12087);
nand U12516 (N_12516,N_12172,N_12201);
or U12517 (N_12517,N_12495,N_12288);
nor U12518 (N_12518,N_12098,N_12199);
nand U12519 (N_12519,N_12375,N_12485);
nor U12520 (N_12520,N_12077,N_12327);
nor U12521 (N_12521,N_12192,N_12361);
nor U12522 (N_12522,N_12364,N_12324);
xnor U12523 (N_12523,N_12249,N_12073);
nor U12524 (N_12524,N_12437,N_12053);
xor U12525 (N_12525,N_12491,N_12180);
or U12526 (N_12526,N_12457,N_12012);
xnor U12527 (N_12527,N_12312,N_12031);
or U12528 (N_12528,N_12422,N_12114);
nor U12529 (N_12529,N_12260,N_12038);
nand U12530 (N_12530,N_12445,N_12307);
nor U12531 (N_12531,N_12146,N_12133);
and U12532 (N_12532,N_12349,N_12497);
nor U12533 (N_12533,N_12309,N_12158);
xor U12534 (N_12534,N_12238,N_12430);
and U12535 (N_12535,N_12377,N_12149);
and U12536 (N_12536,N_12332,N_12231);
xnor U12537 (N_12537,N_12496,N_12423);
nand U12538 (N_12538,N_12454,N_12449);
xor U12539 (N_12539,N_12218,N_12226);
and U12540 (N_12540,N_12023,N_12058);
xnor U12541 (N_12541,N_12335,N_12447);
and U12542 (N_12542,N_12069,N_12066);
nand U12543 (N_12543,N_12246,N_12126);
nor U12544 (N_12544,N_12369,N_12243);
or U12545 (N_12545,N_12384,N_12156);
xor U12546 (N_12546,N_12438,N_12020);
and U12547 (N_12547,N_12019,N_12101);
xor U12548 (N_12548,N_12297,N_12376);
xnor U12549 (N_12549,N_12305,N_12444);
xor U12550 (N_12550,N_12223,N_12253);
nand U12551 (N_12551,N_12263,N_12217);
xor U12552 (N_12552,N_12308,N_12366);
nand U12553 (N_12553,N_12435,N_12125);
xnor U12554 (N_12554,N_12235,N_12267);
nand U12555 (N_12555,N_12167,N_12175);
nand U12556 (N_12556,N_12410,N_12144);
xnor U12557 (N_12557,N_12042,N_12278);
or U12558 (N_12558,N_12266,N_12314);
and U12559 (N_12559,N_12034,N_12321);
or U12560 (N_12560,N_12443,N_12106);
or U12561 (N_12561,N_12416,N_12448);
xnor U12562 (N_12562,N_12441,N_12390);
xor U12563 (N_12563,N_12436,N_12465);
nor U12564 (N_12564,N_12385,N_12303);
nand U12565 (N_12565,N_12245,N_12221);
nor U12566 (N_12566,N_12184,N_12493);
nand U12567 (N_12567,N_12228,N_12459);
and U12568 (N_12568,N_12000,N_12434);
nand U12569 (N_12569,N_12343,N_12396);
or U12570 (N_12570,N_12124,N_12388);
xor U12571 (N_12571,N_12372,N_12382);
and U12572 (N_12572,N_12313,N_12426);
nand U12573 (N_12573,N_12100,N_12183);
nor U12574 (N_12574,N_12212,N_12011);
nand U12575 (N_12575,N_12214,N_12287);
and U12576 (N_12576,N_12189,N_12090);
xnor U12577 (N_12577,N_12295,N_12320);
and U12578 (N_12578,N_12452,N_12211);
or U12579 (N_12579,N_12048,N_12387);
xor U12580 (N_12580,N_12479,N_12113);
xor U12581 (N_12581,N_12052,N_12431);
and U12582 (N_12582,N_12118,N_12174);
and U12583 (N_12583,N_12137,N_12346);
or U12584 (N_12584,N_12272,N_12208);
nand U12585 (N_12585,N_12419,N_12132);
xor U12586 (N_12586,N_12151,N_12049);
nand U12587 (N_12587,N_12425,N_12362);
nand U12588 (N_12588,N_12164,N_12232);
or U12589 (N_12589,N_12254,N_12115);
and U12590 (N_12590,N_12275,N_12001);
nor U12591 (N_12591,N_12472,N_12236);
nand U12592 (N_12592,N_12143,N_12155);
nor U12593 (N_12593,N_12475,N_12400);
or U12594 (N_12594,N_12405,N_12401);
xor U12595 (N_12595,N_12008,N_12379);
xor U12596 (N_12596,N_12055,N_12188);
and U12597 (N_12597,N_12458,N_12061);
xnor U12598 (N_12598,N_12467,N_12096);
nor U12599 (N_12599,N_12354,N_12383);
or U12600 (N_12600,N_12194,N_12138);
xnor U12601 (N_12601,N_12103,N_12112);
nand U12602 (N_12602,N_12097,N_12075);
and U12603 (N_12603,N_12281,N_12002);
or U12604 (N_12604,N_12229,N_12271);
nand U12605 (N_12605,N_12136,N_12094);
nand U12606 (N_12606,N_12262,N_12099);
and U12607 (N_12607,N_12351,N_12499);
nor U12608 (N_12608,N_12230,N_12463);
and U12609 (N_12609,N_12412,N_12006);
nor U12610 (N_12610,N_12045,N_12325);
nor U12611 (N_12611,N_12358,N_12213);
and U12612 (N_12612,N_12484,N_12380);
xor U12613 (N_12613,N_12290,N_12065);
nand U12614 (N_12614,N_12148,N_12153);
nor U12615 (N_12615,N_12378,N_12190);
and U12616 (N_12616,N_12178,N_12169);
or U12617 (N_12617,N_12399,N_12209);
nand U12618 (N_12618,N_12070,N_12326);
and U12619 (N_12619,N_12395,N_12127);
nand U12620 (N_12620,N_12198,N_12004);
and U12621 (N_12621,N_12269,N_12140);
xor U12622 (N_12622,N_12170,N_12131);
xnor U12623 (N_12623,N_12086,N_12119);
and U12624 (N_12624,N_12123,N_12007);
xnor U12625 (N_12625,N_12284,N_12202);
and U12626 (N_12626,N_12080,N_12216);
xnor U12627 (N_12627,N_12227,N_12330);
and U12628 (N_12628,N_12110,N_12043);
or U12629 (N_12629,N_12345,N_12067);
or U12630 (N_12630,N_12340,N_12024);
and U12631 (N_12631,N_12233,N_12046);
xnor U12632 (N_12632,N_12259,N_12062);
or U12633 (N_12633,N_12421,N_12344);
xnor U12634 (N_12634,N_12471,N_12413);
nor U12635 (N_12635,N_12427,N_12187);
or U12636 (N_12636,N_12025,N_12432);
nand U12637 (N_12637,N_12063,N_12109);
nor U12638 (N_12638,N_12050,N_12121);
or U12639 (N_12639,N_12215,N_12311);
nand U12640 (N_12640,N_12182,N_12244);
nor U12641 (N_12641,N_12280,N_12270);
nand U12642 (N_12642,N_12370,N_12365);
and U12643 (N_12643,N_12108,N_12145);
nand U12644 (N_12644,N_12092,N_12173);
nor U12645 (N_12645,N_12300,N_12139);
xnor U12646 (N_12646,N_12161,N_12059);
and U12647 (N_12647,N_12261,N_12195);
and U12648 (N_12648,N_12022,N_12154);
nor U12649 (N_12649,N_12391,N_12021);
nand U12650 (N_12650,N_12466,N_12071);
and U12651 (N_12651,N_12282,N_12250);
nand U12652 (N_12652,N_12339,N_12453);
nand U12653 (N_12653,N_12179,N_12342);
and U12654 (N_12654,N_12206,N_12473);
or U12655 (N_12655,N_12018,N_12219);
nor U12656 (N_12656,N_12424,N_12442);
and U12657 (N_12657,N_12181,N_12408);
nand U12658 (N_12658,N_12350,N_12464);
xor U12659 (N_12659,N_12363,N_12450);
and U12660 (N_12660,N_12009,N_12237);
and U12661 (N_12661,N_12197,N_12392);
xnor U12662 (N_12662,N_12456,N_12296);
nand U12663 (N_12663,N_12141,N_12035);
and U12664 (N_12664,N_12163,N_12005);
or U12665 (N_12665,N_12418,N_12286);
xnor U12666 (N_12666,N_12397,N_12368);
nand U12667 (N_12667,N_12304,N_12283);
and U12668 (N_12668,N_12177,N_12039);
or U12669 (N_12669,N_12347,N_12478);
and U12670 (N_12670,N_12036,N_12468);
nand U12671 (N_12671,N_12374,N_12060);
and U12672 (N_12672,N_12451,N_12079);
and U12673 (N_12673,N_12205,N_12470);
xnor U12674 (N_12674,N_12085,N_12460);
nand U12675 (N_12675,N_12204,N_12057);
nor U12676 (N_12676,N_12247,N_12498);
or U12677 (N_12677,N_12264,N_12054);
xor U12678 (N_12678,N_12040,N_12355);
and U12679 (N_12679,N_12166,N_12122);
nand U12680 (N_12680,N_12248,N_12476);
xnor U12681 (N_12681,N_12028,N_12360);
nand U12682 (N_12682,N_12047,N_12255);
and U12683 (N_12683,N_12352,N_12406);
or U12684 (N_12684,N_12277,N_12095);
and U12685 (N_12685,N_12013,N_12193);
nor U12686 (N_12686,N_12241,N_12257);
or U12687 (N_12687,N_12191,N_12135);
and U12688 (N_12688,N_12064,N_12486);
or U12689 (N_12689,N_12403,N_12029);
xor U12690 (N_12690,N_12433,N_12168);
xor U12691 (N_12691,N_12044,N_12033);
and U12692 (N_12692,N_12323,N_12015);
nor U12693 (N_12693,N_12328,N_12076);
and U12694 (N_12694,N_12494,N_12078);
and U12695 (N_12695,N_12134,N_12276);
xnor U12696 (N_12696,N_12081,N_12310);
and U12697 (N_12697,N_12348,N_12251);
xnor U12698 (N_12698,N_12185,N_12318);
nor U12699 (N_12699,N_12203,N_12084);
xor U12700 (N_12700,N_12274,N_12299);
and U12701 (N_12701,N_12171,N_12315);
or U12702 (N_12702,N_12091,N_12159);
nand U12703 (N_12703,N_12482,N_12428);
nand U12704 (N_12704,N_12489,N_12240);
nor U12705 (N_12705,N_12252,N_12041);
nor U12706 (N_12706,N_12293,N_12337);
nand U12707 (N_12707,N_12116,N_12117);
nand U12708 (N_12708,N_12338,N_12027);
or U12709 (N_12709,N_12341,N_12477);
nand U12710 (N_12710,N_12017,N_12402);
nand U12711 (N_12711,N_12331,N_12032);
and U12712 (N_12712,N_12074,N_12407);
or U12713 (N_12713,N_12152,N_12030);
or U12714 (N_12714,N_12334,N_12336);
or U12715 (N_12715,N_12356,N_12234);
or U12716 (N_12716,N_12120,N_12102);
nand U12717 (N_12717,N_12439,N_12239);
nand U12718 (N_12718,N_12371,N_12107);
and U12719 (N_12719,N_12487,N_12105);
nand U12720 (N_12720,N_12088,N_12165);
or U12721 (N_12721,N_12273,N_12333);
and U12722 (N_12722,N_12225,N_12289);
xor U12723 (N_12723,N_12291,N_12480);
or U12724 (N_12724,N_12414,N_12268);
or U12725 (N_12725,N_12316,N_12186);
and U12726 (N_12726,N_12207,N_12083);
or U12727 (N_12727,N_12222,N_12285);
xor U12728 (N_12728,N_12469,N_12461);
and U12729 (N_12729,N_12429,N_12082);
or U12730 (N_12730,N_12142,N_12446);
or U12731 (N_12731,N_12306,N_12389);
nor U12732 (N_12732,N_12357,N_12014);
and U12733 (N_12733,N_12398,N_12488);
nand U12734 (N_12734,N_12415,N_12068);
nand U12735 (N_12735,N_12089,N_12462);
nor U12736 (N_12736,N_12104,N_12157);
or U12737 (N_12737,N_12353,N_12111);
nor U12738 (N_12738,N_12130,N_12329);
nor U12739 (N_12739,N_12150,N_12359);
and U12740 (N_12740,N_12411,N_12394);
or U12741 (N_12741,N_12417,N_12440);
xor U12742 (N_12742,N_12256,N_12404);
nor U12743 (N_12743,N_12016,N_12258);
or U12744 (N_12744,N_12037,N_12093);
xnor U12745 (N_12745,N_12409,N_12302);
nand U12746 (N_12746,N_12162,N_12056);
nand U12747 (N_12747,N_12128,N_12455);
and U12748 (N_12748,N_12129,N_12210);
nor U12749 (N_12749,N_12242,N_12490);
or U12750 (N_12750,N_12249,N_12378);
or U12751 (N_12751,N_12065,N_12013);
xor U12752 (N_12752,N_12183,N_12493);
nor U12753 (N_12753,N_12170,N_12071);
xor U12754 (N_12754,N_12428,N_12157);
and U12755 (N_12755,N_12258,N_12252);
nor U12756 (N_12756,N_12256,N_12317);
and U12757 (N_12757,N_12034,N_12254);
xor U12758 (N_12758,N_12027,N_12030);
or U12759 (N_12759,N_12380,N_12129);
nand U12760 (N_12760,N_12216,N_12073);
xnor U12761 (N_12761,N_12210,N_12009);
or U12762 (N_12762,N_12125,N_12086);
xor U12763 (N_12763,N_12486,N_12471);
xor U12764 (N_12764,N_12218,N_12320);
xor U12765 (N_12765,N_12389,N_12371);
nor U12766 (N_12766,N_12093,N_12254);
and U12767 (N_12767,N_12014,N_12133);
nand U12768 (N_12768,N_12187,N_12268);
nor U12769 (N_12769,N_12304,N_12045);
xor U12770 (N_12770,N_12174,N_12004);
or U12771 (N_12771,N_12444,N_12325);
nor U12772 (N_12772,N_12451,N_12261);
nand U12773 (N_12773,N_12349,N_12131);
or U12774 (N_12774,N_12256,N_12030);
or U12775 (N_12775,N_12063,N_12098);
or U12776 (N_12776,N_12107,N_12047);
and U12777 (N_12777,N_12412,N_12066);
nand U12778 (N_12778,N_12034,N_12187);
nor U12779 (N_12779,N_12102,N_12150);
or U12780 (N_12780,N_12020,N_12024);
nor U12781 (N_12781,N_12055,N_12119);
and U12782 (N_12782,N_12174,N_12395);
or U12783 (N_12783,N_12087,N_12191);
nor U12784 (N_12784,N_12008,N_12132);
nor U12785 (N_12785,N_12422,N_12407);
or U12786 (N_12786,N_12471,N_12129);
or U12787 (N_12787,N_12248,N_12037);
nand U12788 (N_12788,N_12064,N_12422);
and U12789 (N_12789,N_12305,N_12021);
xor U12790 (N_12790,N_12016,N_12105);
or U12791 (N_12791,N_12442,N_12433);
nand U12792 (N_12792,N_12011,N_12311);
nand U12793 (N_12793,N_12240,N_12244);
or U12794 (N_12794,N_12221,N_12195);
or U12795 (N_12795,N_12459,N_12178);
nand U12796 (N_12796,N_12348,N_12490);
nor U12797 (N_12797,N_12074,N_12451);
xnor U12798 (N_12798,N_12237,N_12496);
or U12799 (N_12799,N_12175,N_12147);
nor U12800 (N_12800,N_12311,N_12308);
or U12801 (N_12801,N_12006,N_12304);
or U12802 (N_12802,N_12302,N_12173);
nor U12803 (N_12803,N_12270,N_12129);
nand U12804 (N_12804,N_12476,N_12404);
xnor U12805 (N_12805,N_12344,N_12114);
nor U12806 (N_12806,N_12155,N_12160);
nand U12807 (N_12807,N_12322,N_12332);
xor U12808 (N_12808,N_12261,N_12061);
or U12809 (N_12809,N_12463,N_12086);
or U12810 (N_12810,N_12201,N_12459);
and U12811 (N_12811,N_12141,N_12407);
nor U12812 (N_12812,N_12344,N_12225);
xnor U12813 (N_12813,N_12182,N_12386);
nand U12814 (N_12814,N_12303,N_12309);
xor U12815 (N_12815,N_12251,N_12241);
or U12816 (N_12816,N_12357,N_12171);
or U12817 (N_12817,N_12034,N_12437);
or U12818 (N_12818,N_12068,N_12352);
xor U12819 (N_12819,N_12243,N_12079);
and U12820 (N_12820,N_12140,N_12151);
nand U12821 (N_12821,N_12477,N_12457);
and U12822 (N_12822,N_12227,N_12381);
xor U12823 (N_12823,N_12030,N_12127);
nor U12824 (N_12824,N_12128,N_12239);
nor U12825 (N_12825,N_12415,N_12250);
nand U12826 (N_12826,N_12466,N_12134);
xnor U12827 (N_12827,N_12267,N_12215);
or U12828 (N_12828,N_12086,N_12095);
and U12829 (N_12829,N_12138,N_12483);
nand U12830 (N_12830,N_12233,N_12121);
or U12831 (N_12831,N_12308,N_12483);
nand U12832 (N_12832,N_12170,N_12166);
nand U12833 (N_12833,N_12131,N_12001);
or U12834 (N_12834,N_12008,N_12080);
or U12835 (N_12835,N_12281,N_12453);
xnor U12836 (N_12836,N_12341,N_12161);
xor U12837 (N_12837,N_12256,N_12373);
and U12838 (N_12838,N_12286,N_12282);
nor U12839 (N_12839,N_12375,N_12092);
nor U12840 (N_12840,N_12290,N_12069);
xnor U12841 (N_12841,N_12003,N_12441);
or U12842 (N_12842,N_12308,N_12175);
nand U12843 (N_12843,N_12464,N_12032);
or U12844 (N_12844,N_12227,N_12106);
nor U12845 (N_12845,N_12469,N_12196);
or U12846 (N_12846,N_12284,N_12081);
xnor U12847 (N_12847,N_12406,N_12271);
nand U12848 (N_12848,N_12198,N_12318);
nor U12849 (N_12849,N_12284,N_12432);
xnor U12850 (N_12850,N_12204,N_12326);
or U12851 (N_12851,N_12072,N_12160);
and U12852 (N_12852,N_12273,N_12038);
xor U12853 (N_12853,N_12147,N_12241);
nor U12854 (N_12854,N_12307,N_12117);
or U12855 (N_12855,N_12346,N_12144);
and U12856 (N_12856,N_12447,N_12237);
and U12857 (N_12857,N_12294,N_12167);
and U12858 (N_12858,N_12466,N_12215);
xor U12859 (N_12859,N_12096,N_12047);
and U12860 (N_12860,N_12128,N_12318);
or U12861 (N_12861,N_12204,N_12049);
or U12862 (N_12862,N_12414,N_12467);
or U12863 (N_12863,N_12294,N_12300);
and U12864 (N_12864,N_12124,N_12334);
nand U12865 (N_12865,N_12460,N_12020);
nand U12866 (N_12866,N_12319,N_12070);
nor U12867 (N_12867,N_12465,N_12220);
or U12868 (N_12868,N_12395,N_12006);
xnor U12869 (N_12869,N_12003,N_12317);
and U12870 (N_12870,N_12357,N_12315);
or U12871 (N_12871,N_12353,N_12079);
nand U12872 (N_12872,N_12345,N_12415);
xnor U12873 (N_12873,N_12350,N_12361);
nand U12874 (N_12874,N_12367,N_12397);
xnor U12875 (N_12875,N_12173,N_12156);
nor U12876 (N_12876,N_12417,N_12369);
nand U12877 (N_12877,N_12054,N_12232);
or U12878 (N_12878,N_12230,N_12112);
nor U12879 (N_12879,N_12006,N_12383);
nand U12880 (N_12880,N_12482,N_12011);
and U12881 (N_12881,N_12098,N_12289);
or U12882 (N_12882,N_12334,N_12428);
and U12883 (N_12883,N_12117,N_12246);
or U12884 (N_12884,N_12137,N_12244);
nand U12885 (N_12885,N_12322,N_12074);
nor U12886 (N_12886,N_12068,N_12142);
and U12887 (N_12887,N_12033,N_12300);
or U12888 (N_12888,N_12415,N_12243);
nor U12889 (N_12889,N_12353,N_12004);
nor U12890 (N_12890,N_12374,N_12258);
and U12891 (N_12891,N_12170,N_12463);
and U12892 (N_12892,N_12141,N_12038);
xor U12893 (N_12893,N_12479,N_12412);
nor U12894 (N_12894,N_12348,N_12144);
xor U12895 (N_12895,N_12122,N_12393);
or U12896 (N_12896,N_12015,N_12437);
and U12897 (N_12897,N_12219,N_12033);
nor U12898 (N_12898,N_12278,N_12424);
or U12899 (N_12899,N_12036,N_12212);
or U12900 (N_12900,N_12064,N_12175);
nand U12901 (N_12901,N_12329,N_12152);
or U12902 (N_12902,N_12169,N_12321);
nand U12903 (N_12903,N_12260,N_12026);
xnor U12904 (N_12904,N_12377,N_12471);
or U12905 (N_12905,N_12391,N_12333);
nand U12906 (N_12906,N_12426,N_12016);
nand U12907 (N_12907,N_12427,N_12300);
nand U12908 (N_12908,N_12302,N_12330);
xnor U12909 (N_12909,N_12490,N_12154);
nor U12910 (N_12910,N_12161,N_12320);
or U12911 (N_12911,N_12082,N_12416);
or U12912 (N_12912,N_12423,N_12441);
and U12913 (N_12913,N_12225,N_12195);
xor U12914 (N_12914,N_12058,N_12448);
nand U12915 (N_12915,N_12058,N_12033);
nand U12916 (N_12916,N_12132,N_12118);
xor U12917 (N_12917,N_12291,N_12497);
and U12918 (N_12918,N_12161,N_12379);
xnor U12919 (N_12919,N_12284,N_12323);
nor U12920 (N_12920,N_12390,N_12179);
nand U12921 (N_12921,N_12025,N_12043);
nand U12922 (N_12922,N_12344,N_12196);
and U12923 (N_12923,N_12351,N_12105);
nor U12924 (N_12924,N_12323,N_12467);
and U12925 (N_12925,N_12013,N_12435);
or U12926 (N_12926,N_12057,N_12026);
and U12927 (N_12927,N_12399,N_12133);
nor U12928 (N_12928,N_12395,N_12428);
xnor U12929 (N_12929,N_12200,N_12326);
and U12930 (N_12930,N_12294,N_12168);
nand U12931 (N_12931,N_12138,N_12001);
nand U12932 (N_12932,N_12170,N_12122);
and U12933 (N_12933,N_12269,N_12105);
nor U12934 (N_12934,N_12223,N_12466);
xor U12935 (N_12935,N_12104,N_12105);
nand U12936 (N_12936,N_12163,N_12467);
and U12937 (N_12937,N_12009,N_12068);
nand U12938 (N_12938,N_12177,N_12414);
nand U12939 (N_12939,N_12138,N_12492);
and U12940 (N_12940,N_12186,N_12420);
nor U12941 (N_12941,N_12447,N_12443);
nand U12942 (N_12942,N_12008,N_12460);
or U12943 (N_12943,N_12403,N_12499);
and U12944 (N_12944,N_12012,N_12455);
nand U12945 (N_12945,N_12300,N_12353);
or U12946 (N_12946,N_12291,N_12477);
nand U12947 (N_12947,N_12162,N_12294);
or U12948 (N_12948,N_12269,N_12406);
and U12949 (N_12949,N_12428,N_12327);
and U12950 (N_12950,N_12326,N_12269);
nor U12951 (N_12951,N_12184,N_12386);
nor U12952 (N_12952,N_12288,N_12205);
nor U12953 (N_12953,N_12144,N_12293);
nor U12954 (N_12954,N_12406,N_12347);
and U12955 (N_12955,N_12384,N_12130);
nor U12956 (N_12956,N_12096,N_12466);
nor U12957 (N_12957,N_12086,N_12248);
xnor U12958 (N_12958,N_12442,N_12362);
or U12959 (N_12959,N_12476,N_12268);
nand U12960 (N_12960,N_12217,N_12381);
nor U12961 (N_12961,N_12202,N_12159);
nand U12962 (N_12962,N_12226,N_12320);
nor U12963 (N_12963,N_12279,N_12084);
or U12964 (N_12964,N_12389,N_12227);
and U12965 (N_12965,N_12311,N_12118);
or U12966 (N_12966,N_12420,N_12155);
nor U12967 (N_12967,N_12296,N_12458);
or U12968 (N_12968,N_12199,N_12301);
and U12969 (N_12969,N_12004,N_12357);
xor U12970 (N_12970,N_12314,N_12339);
or U12971 (N_12971,N_12215,N_12290);
xor U12972 (N_12972,N_12463,N_12471);
nor U12973 (N_12973,N_12175,N_12003);
xor U12974 (N_12974,N_12092,N_12238);
or U12975 (N_12975,N_12391,N_12222);
nor U12976 (N_12976,N_12178,N_12061);
and U12977 (N_12977,N_12320,N_12212);
nor U12978 (N_12978,N_12391,N_12353);
or U12979 (N_12979,N_12231,N_12001);
nand U12980 (N_12980,N_12356,N_12014);
and U12981 (N_12981,N_12441,N_12333);
nand U12982 (N_12982,N_12429,N_12487);
nand U12983 (N_12983,N_12115,N_12475);
nand U12984 (N_12984,N_12411,N_12049);
xnor U12985 (N_12985,N_12305,N_12225);
and U12986 (N_12986,N_12136,N_12113);
xnor U12987 (N_12987,N_12190,N_12280);
nand U12988 (N_12988,N_12035,N_12423);
xnor U12989 (N_12989,N_12228,N_12355);
nand U12990 (N_12990,N_12249,N_12209);
and U12991 (N_12991,N_12282,N_12251);
nand U12992 (N_12992,N_12307,N_12035);
xnor U12993 (N_12993,N_12096,N_12057);
nand U12994 (N_12994,N_12049,N_12312);
nor U12995 (N_12995,N_12394,N_12091);
nand U12996 (N_12996,N_12337,N_12454);
and U12997 (N_12997,N_12061,N_12149);
or U12998 (N_12998,N_12377,N_12388);
nand U12999 (N_12999,N_12168,N_12245);
or U13000 (N_13000,N_12938,N_12691);
xnor U13001 (N_13001,N_12931,N_12895);
or U13002 (N_13002,N_12943,N_12884);
or U13003 (N_13003,N_12799,N_12589);
xor U13004 (N_13004,N_12784,N_12665);
and U13005 (N_13005,N_12526,N_12578);
xnor U13006 (N_13006,N_12743,N_12758);
and U13007 (N_13007,N_12571,N_12876);
xor U13008 (N_13008,N_12704,N_12961);
xor U13009 (N_13009,N_12654,N_12970);
nor U13010 (N_13010,N_12637,N_12983);
xnor U13011 (N_13011,N_12671,N_12683);
nand U13012 (N_13012,N_12832,N_12998);
xnor U13013 (N_13013,N_12669,N_12639);
or U13014 (N_13014,N_12753,N_12993);
or U13015 (N_13015,N_12772,N_12502);
xnor U13016 (N_13016,N_12768,N_12607);
or U13017 (N_13017,N_12825,N_12694);
nor U13018 (N_13018,N_12572,N_12558);
or U13019 (N_13019,N_12527,N_12985);
and U13020 (N_13020,N_12932,N_12664);
xnor U13021 (N_13021,N_12569,N_12650);
xor U13022 (N_13022,N_12816,N_12532);
xor U13023 (N_13023,N_12919,N_12969);
nor U13024 (N_13024,N_12543,N_12765);
nand U13025 (N_13025,N_12864,N_12666);
xor U13026 (N_13026,N_12732,N_12830);
xnor U13027 (N_13027,N_12869,N_12673);
xor U13028 (N_13028,N_12723,N_12838);
nor U13029 (N_13029,N_12531,N_12847);
nand U13030 (N_13030,N_12951,N_12802);
and U13031 (N_13031,N_12924,N_12793);
or U13032 (N_13032,N_12903,N_12948);
nor U13033 (N_13033,N_12600,N_12894);
nor U13034 (N_13034,N_12892,N_12852);
nor U13035 (N_13035,N_12696,N_12806);
nand U13036 (N_13036,N_12862,N_12634);
xnor U13037 (N_13037,N_12672,N_12522);
xnor U13038 (N_13038,N_12503,N_12795);
nand U13039 (N_13039,N_12556,N_12833);
and U13040 (N_13040,N_12831,N_12785);
and U13041 (N_13041,N_12926,N_12810);
xor U13042 (N_13042,N_12557,N_12929);
xor U13043 (N_13043,N_12540,N_12706);
or U13044 (N_13044,N_12984,N_12877);
nor U13045 (N_13045,N_12939,N_12563);
nor U13046 (N_13046,N_12697,N_12724);
nor U13047 (N_13047,N_12937,N_12656);
or U13048 (N_13048,N_12515,N_12859);
nand U13049 (N_13049,N_12609,N_12834);
nand U13050 (N_13050,N_12570,N_12875);
or U13051 (N_13051,N_12586,N_12850);
xnor U13052 (N_13052,N_12788,N_12813);
nand U13053 (N_13053,N_12516,N_12963);
and U13054 (N_13054,N_12628,N_12837);
xor U13055 (N_13055,N_12674,N_12818);
and U13056 (N_13056,N_12787,N_12521);
xnor U13057 (N_13057,N_12510,N_12551);
nor U13058 (N_13058,N_12716,N_12766);
and U13059 (N_13059,N_12685,N_12509);
nand U13060 (N_13060,N_12635,N_12855);
nor U13061 (N_13061,N_12541,N_12804);
xor U13062 (N_13062,N_12646,N_12579);
nand U13063 (N_13063,N_12536,N_12524);
xnor U13064 (N_13064,N_12715,N_12982);
nand U13065 (N_13065,N_12575,N_12971);
or U13066 (N_13066,N_12559,N_12775);
nand U13067 (N_13067,N_12588,N_12949);
and U13068 (N_13068,N_12667,N_12501);
or U13069 (N_13069,N_12591,N_12690);
nor U13070 (N_13070,N_12812,N_12796);
nand U13071 (N_13071,N_12987,N_12921);
and U13072 (N_13072,N_12678,N_12631);
nand U13073 (N_13073,N_12920,N_12616);
and U13074 (N_13074,N_12925,N_12670);
and U13075 (N_13075,N_12566,N_12722);
nor U13076 (N_13076,N_12955,N_12528);
and U13077 (N_13077,N_12822,N_12729);
or U13078 (N_13078,N_12801,N_12781);
or U13079 (N_13079,N_12930,N_12885);
or U13080 (N_13080,N_12956,N_12596);
nand U13081 (N_13081,N_12618,N_12874);
or U13082 (N_13082,N_12611,N_12771);
or U13083 (N_13083,N_12786,N_12720);
or U13084 (N_13084,N_12908,N_12861);
and U13085 (N_13085,N_12725,N_12649);
and U13086 (N_13086,N_12907,N_12583);
or U13087 (N_13087,N_12811,N_12975);
and U13088 (N_13088,N_12703,N_12546);
nor U13089 (N_13089,N_12817,N_12750);
xnor U13090 (N_13090,N_12657,N_12549);
and U13091 (N_13091,N_12644,N_12742);
nor U13092 (N_13092,N_12538,N_12680);
nor U13093 (N_13093,N_12594,N_12564);
nand U13094 (N_13094,N_12782,N_12809);
or U13095 (N_13095,N_12581,N_12870);
nor U13096 (N_13096,N_12805,N_12980);
nor U13097 (N_13097,N_12945,N_12610);
nor U13098 (N_13098,N_12574,N_12829);
xnor U13099 (N_13099,N_12681,N_12573);
nand U13100 (N_13100,N_12641,N_12994);
xor U13101 (N_13101,N_12916,N_12887);
and U13102 (N_13102,N_12754,N_12560);
and U13103 (N_13103,N_12647,N_12880);
or U13104 (N_13104,N_12783,N_12867);
or U13105 (N_13105,N_12648,N_12555);
nand U13106 (N_13106,N_12617,N_12719);
and U13107 (N_13107,N_12651,N_12709);
and U13108 (N_13108,N_12584,N_12565);
nor U13109 (N_13109,N_12845,N_12606);
nor U13110 (N_13110,N_12652,N_12827);
nor U13111 (N_13111,N_12953,N_12632);
nand U13112 (N_13112,N_12890,N_12590);
or U13113 (N_13113,N_12899,N_12917);
xor U13114 (N_13114,N_12821,N_12530);
and U13115 (N_13115,N_12624,N_12506);
nor U13116 (N_13116,N_12577,N_12967);
xnor U13117 (N_13117,N_12554,N_12730);
nand U13118 (N_13118,N_12776,N_12941);
and U13119 (N_13119,N_12707,N_12755);
xor U13120 (N_13120,N_12645,N_12759);
or U13121 (N_13121,N_12595,N_12815);
nor U13122 (N_13122,N_12737,N_12636);
or U13123 (N_13123,N_12947,N_12547);
nor U13124 (N_13124,N_12981,N_12886);
nor U13125 (N_13125,N_12711,N_12901);
xnor U13126 (N_13126,N_12918,N_12507);
nand U13127 (N_13127,N_12604,N_12905);
nor U13128 (N_13128,N_12620,N_12902);
and U13129 (N_13129,N_12798,N_12760);
or U13130 (N_13130,N_12705,N_12548);
nand U13131 (N_13131,N_12807,N_12841);
or U13132 (N_13132,N_12512,N_12800);
or U13133 (N_13133,N_12585,N_12687);
and U13134 (N_13134,N_12655,N_12602);
nor U13135 (N_13135,N_12839,N_12593);
nand U13136 (N_13136,N_12851,N_12950);
nor U13137 (N_13137,N_12819,N_12519);
nor U13138 (N_13138,N_12973,N_12601);
or U13139 (N_13139,N_12679,N_12576);
xnor U13140 (N_13140,N_12525,N_12808);
and U13141 (N_13141,N_12695,N_12935);
xor U13142 (N_13142,N_12702,N_12746);
xor U13143 (N_13143,N_12848,N_12965);
nor U13144 (N_13144,N_12944,N_12523);
xnor U13145 (N_13145,N_12625,N_12996);
nand U13146 (N_13146,N_12844,N_12520);
xor U13147 (N_13147,N_12535,N_12853);
and U13148 (N_13148,N_12627,N_12739);
and U13149 (N_13149,N_12708,N_12741);
nor U13150 (N_13150,N_12764,N_12779);
and U13151 (N_13151,N_12643,N_12675);
or U13152 (N_13152,N_12663,N_12888);
or U13153 (N_13153,N_12964,N_12789);
nor U13154 (N_13154,N_12505,N_12717);
nor U13155 (N_13155,N_12668,N_12659);
nor U13156 (N_13156,N_12909,N_12605);
and U13157 (N_13157,N_12952,N_12774);
and U13158 (N_13158,N_12626,N_12726);
or U13159 (N_13159,N_12959,N_12979);
or U13160 (N_13160,N_12871,N_12721);
or U13161 (N_13161,N_12684,N_12824);
xnor U13162 (N_13162,N_12597,N_12769);
and U13163 (N_13163,N_12913,N_12912);
nand U13164 (N_13164,N_12962,N_12533);
nor U13165 (N_13165,N_12738,N_12748);
and U13166 (N_13166,N_12968,N_12797);
nor U13167 (N_13167,N_12803,N_12761);
nand U13168 (N_13168,N_12992,N_12794);
and U13169 (N_13169,N_12836,N_12910);
and U13170 (N_13170,N_12988,N_12991);
xnor U13171 (N_13171,N_12661,N_12642);
and U13172 (N_13172,N_12791,N_12835);
nor U13173 (N_13173,N_12872,N_12744);
nor U13174 (N_13174,N_12727,N_12599);
and U13175 (N_13175,N_12915,N_12603);
nand U13176 (N_13176,N_12904,N_12517);
and U13177 (N_13177,N_12922,N_12828);
nand U13178 (N_13178,N_12677,N_12692);
and U13179 (N_13179,N_12820,N_12640);
and U13180 (N_13180,N_12733,N_12728);
xnor U13181 (N_13181,N_12686,N_12700);
nor U13182 (N_13182,N_12508,N_12749);
xor U13183 (N_13183,N_12747,N_12972);
and U13184 (N_13184,N_12553,N_12658);
and U13185 (N_13185,N_12545,N_12843);
nand U13186 (N_13186,N_12978,N_12736);
nand U13187 (N_13187,N_12986,N_12745);
nand U13188 (N_13188,N_12762,N_12757);
and U13189 (N_13189,N_12500,N_12714);
xnor U13190 (N_13190,N_12633,N_12814);
nor U13191 (N_13191,N_12638,N_12630);
nor U13192 (N_13192,N_12731,N_12756);
and U13193 (N_13193,N_12740,N_12712);
and U13194 (N_13194,N_12866,N_12999);
nand U13195 (N_13195,N_12580,N_12790);
and U13196 (N_13196,N_12752,N_12763);
nor U13197 (N_13197,N_12878,N_12954);
xnor U13198 (N_13198,N_12623,N_12881);
xor U13199 (N_13199,N_12621,N_12896);
and U13200 (N_13200,N_12868,N_12863);
or U13201 (N_13201,N_12842,N_12928);
nor U13202 (N_13202,N_12568,N_12898);
xor U13203 (N_13203,N_12865,N_12858);
xnor U13204 (N_13204,N_12770,N_12662);
nand U13205 (N_13205,N_12966,N_12989);
or U13206 (N_13206,N_12936,N_12561);
and U13207 (N_13207,N_12735,N_12792);
or U13208 (N_13208,N_12823,N_12734);
xnor U13209 (N_13209,N_12552,N_12882);
nor U13210 (N_13210,N_12544,N_12897);
nor U13211 (N_13211,N_12710,N_12906);
xor U13212 (N_13212,N_12854,N_12511);
nand U13213 (N_13213,N_12539,N_12562);
or U13214 (N_13214,N_12856,N_12653);
xnor U13215 (N_13215,N_12958,N_12693);
nor U13216 (N_13216,N_12614,N_12718);
xor U13217 (N_13217,N_12587,N_12960);
and U13218 (N_13218,N_12629,N_12891);
and U13219 (N_13219,N_12780,N_12701);
and U13220 (N_13220,N_12934,N_12777);
nor U13221 (N_13221,N_12826,N_12598);
nand U13222 (N_13222,N_12612,N_12608);
and U13223 (N_13223,N_12840,N_12615);
and U13224 (N_13224,N_12582,N_12900);
and U13225 (N_13225,N_12550,N_12860);
or U13226 (N_13226,N_12518,N_12622);
nand U13227 (N_13227,N_12514,N_12914);
xnor U13228 (N_13228,N_12873,N_12889);
nor U13229 (N_13229,N_12676,N_12688);
nand U13230 (N_13230,N_12773,N_12857);
and U13231 (N_13231,N_12592,N_12534);
nor U13232 (N_13232,N_12542,N_12751);
or U13233 (N_13233,N_12923,N_12849);
and U13234 (N_13234,N_12974,N_12619);
nand U13235 (N_13235,N_12879,N_12976);
nand U13236 (N_13236,N_12911,N_12957);
and U13237 (N_13237,N_12990,N_12940);
nand U13238 (N_13238,N_12942,N_12537);
or U13239 (N_13239,N_12504,N_12946);
or U13240 (N_13240,N_12660,N_12699);
and U13241 (N_13241,N_12689,N_12682);
nor U13242 (N_13242,N_12933,N_12997);
or U13243 (N_13243,N_12977,N_12767);
xor U13244 (N_13244,N_12613,N_12698);
xor U13245 (N_13245,N_12883,N_12713);
or U13246 (N_13246,N_12778,N_12995);
xor U13247 (N_13247,N_12846,N_12893);
nor U13248 (N_13248,N_12567,N_12513);
xor U13249 (N_13249,N_12529,N_12927);
xor U13250 (N_13250,N_12608,N_12782);
nor U13251 (N_13251,N_12633,N_12701);
xnor U13252 (N_13252,N_12852,N_12591);
xnor U13253 (N_13253,N_12639,N_12589);
or U13254 (N_13254,N_12793,N_12576);
and U13255 (N_13255,N_12535,N_12716);
and U13256 (N_13256,N_12656,N_12839);
nor U13257 (N_13257,N_12705,N_12935);
nand U13258 (N_13258,N_12727,N_12820);
nand U13259 (N_13259,N_12555,N_12691);
xnor U13260 (N_13260,N_12643,N_12823);
or U13261 (N_13261,N_12758,N_12692);
xor U13262 (N_13262,N_12515,N_12616);
xor U13263 (N_13263,N_12922,N_12505);
nand U13264 (N_13264,N_12525,N_12773);
or U13265 (N_13265,N_12679,N_12634);
nor U13266 (N_13266,N_12995,N_12944);
xor U13267 (N_13267,N_12583,N_12561);
xor U13268 (N_13268,N_12520,N_12944);
nand U13269 (N_13269,N_12999,N_12535);
nand U13270 (N_13270,N_12740,N_12868);
nand U13271 (N_13271,N_12884,N_12730);
nor U13272 (N_13272,N_12897,N_12972);
nor U13273 (N_13273,N_12978,N_12861);
xnor U13274 (N_13274,N_12613,N_12972);
or U13275 (N_13275,N_12600,N_12897);
nor U13276 (N_13276,N_12841,N_12731);
nor U13277 (N_13277,N_12627,N_12770);
or U13278 (N_13278,N_12580,N_12621);
nor U13279 (N_13279,N_12541,N_12730);
nand U13280 (N_13280,N_12568,N_12883);
and U13281 (N_13281,N_12500,N_12509);
and U13282 (N_13282,N_12601,N_12980);
xnor U13283 (N_13283,N_12554,N_12941);
nand U13284 (N_13284,N_12554,N_12991);
and U13285 (N_13285,N_12717,N_12763);
nor U13286 (N_13286,N_12888,N_12792);
and U13287 (N_13287,N_12914,N_12670);
nand U13288 (N_13288,N_12734,N_12707);
nand U13289 (N_13289,N_12522,N_12912);
nor U13290 (N_13290,N_12710,N_12636);
or U13291 (N_13291,N_12710,N_12786);
or U13292 (N_13292,N_12951,N_12558);
nor U13293 (N_13293,N_12824,N_12530);
or U13294 (N_13294,N_12590,N_12653);
xor U13295 (N_13295,N_12709,N_12500);
or U13296 (N_13296,N_12961,N_12510);
xor U13297 (N_13297,N_12950,N_12986);
and U13298 (N_13298,N_12704,N_12536);
nand U13299 (N_13299,N_12552,N_12801);
nor U13300 (N_13300,N_12683,N_12829);
xor U13301 (N_13301,N_12778,N_12595);
nand U13302 (N_13302,N_12701,N_12536);
and U13303 (N_13303,N_12879,N_12956);
xor U13304 (N_13304,N_12677,N_12985);
or U13305 (N_13305,N_12701,N_12951);
xor U13306 (N_13306,N_12917,N_12722);
nor U13307 (N_13307,N_12508,N_12506);
nand U13308 (N_13308,N_12982,N_12808);
and U13309 (N_13309,N_12753,N_12942);
and U13310 (N_13310,N_12642,N_12610);
and U13311 (N_13311,N_12525,N_12915);
nand U13312 (N_13312,N_12925,N_12705);
nand U13313 (N_13313,N_12964,N_12835);
or U13314 (N_13314,N_12578,N_12644);
nor U13315 (N_13315,N_12997,N_12881);
nor U13316 (N_13316,N_12523,N_12510);
nand U13317 (N_13317,N_12959,N_12778);
nor U13318 (N_13318,N_12610,N_12648);
nand U13319 (N_13319,N_12507,N_12641);
nand U13320 (N_13320,N_12836,N_12596);
or U13321 (N_13321,N_12514,N_12959);
and U13322 (N_13322,N_12928,N_12536);
xnor U13323 (N_13323,N_12692,N_12948);
xor U13324 (N_13324,N_12861,N_12977);
nor U13325 (N_13325,N_12649,N_12922);
nor U13326 (N_13326,N_12925,N_12654);
and U13327 (N_13327,N_12974,N_12582);
nand U13328 (N_13328,N_12722,N_12907);
nand U13329 (N_13329,N_12702,N_12846);
nand U13330 (N_13330,N_12527,N_12763);
or U13331 (N_13331,N_12680,N_12803);
and U13332 (N_13332,N_12747,N_12578);
nor U13333 (N_13333,N_12610,N_12715);
and U13334 (N_13334,N_12724,N_12888);
nand U13335 (N_13335,N_12517,N_12509);
xor U13336 (N_13336,N_12774,N_12708);
nand U13337 (N_13337,N_12972,N_12925);
and U13338 (N_13338,N_12546,N_12828);
nor U13339 (N_13339,N_12671,N_12551);
or U13340 (N_13340,N_12543,N_12678);
nand U13341 (N_13341,N_12642,N_12905);
nor U13342 (N_13342,N_12618,N_12915);
nand U13343 (N_13343,N_12945,N_12988);
nor U13344 (N_13344,N_12954,N_12676);
nor U13345 (N_13345,N_12990,N_12974);
nor U13346 (N_13346,N_12735,N_12956);
and U13347 (N_13347,N_12713,N_12962);
and U13348 (N_13348,N_12872,N_12538);
nor U13349 (N_13349,N_12964,N_12688);
and U13350 (N_13350,N_12635,N_12719);
and U13351 (N_13351,N_12845,N_12536);
nor U13352 (N_13352,N_12801,N_12661);
and U13353 (N_13353,N_12735,N_12592);
nand U13354 (N_13354,N_12827,N_12935);
or U13355 (N_13355,N_12866,N_12569);
nand U13356 (N_13356,N_12802,N_12584);
or U13357 (N_13357,N_12762,N_12821);
and U13358 (N_13358,N_12797,N_12757);
nor U13359 (N_13359,N_12669,N_12749);
or U13360 (N_13360,N_12823,N_12944);
nor U13361 (N_13361,N_12542,N_12899);
xor U13362 (N_13362,N_12997,N_12943);
and U13363 (N_13363,N_12661,N_12843);
nor U13364 (N_13364,N_12534,N_12917);
xnor U13365 (N_13365,N_12851,N_12747);
and U13366 (N_13366,N_12634,N_12945);
xor U13367 (N_13367,N_12891,N_12507);
xnor U13368 (N_13368,N_12728,N_12865);
and U13369 (N_13369,N_12865,N_12765);
nor U13370 (N_13370,N_12541,N_12855);
or U13371 (N_13371,N_12773,N_12677);
nand U13372 (N_13372,N_12792,N_12896);
nand U13373 (N_13373,N_12750,N_12531);
or U13374 (N_13374,N_12914,N_12805);
xnor U13375 (N_13375,N_12878,N_12609);
nor U13376 (N_13376,N_12621,N_12574);
xnor U13377 (N_13377,N_12502,N_12848);
xor U13378 (N_13378,N_12954,N_12898);
and U13379 (N_13379,N_12667,N_12943);
nor U13380 (N_13380,N_12770,N_12610);
and U13381 (N_13381,N_12886,N_12973);
nor U13382 (N_13382,N_12657,N_12868);
nor U13383 (N_13383,N_12602,N_12548);
nand U13384 (N_13384,N_12962,N_12851);
nor U13385 (N_13385,N_12827,N_12922);
xor U13386 (N_13386,N_12897,N_12743);
xnor U13387 (N_13387,N_12860,N_12948);
nand U13388 (N_13388,N_12624,N_12857);
nand U13389 (N_13389,N_12888,N_12849);
nor U13390 (N_13390,N_12886,N_12681);
xor U13391 (N_13391,N_12562,N_12502);
xor U13392 (N_13392,N_12971,N_12792);
or U13393 (N_13393,N_12867,N_12670);
nand U13394 (N_13394,N_12882,N_12820);
or U13395 (N_13395,N_12575,N_12641);
xor U13396 (N_13396,N_12993,N_12693);
nor U13397 (N_13397,N_12989,N_12611);
nor U13398 (N_13398,N_12512,N_12852);
and U13399 (N_13399,N_12692,N_12845);
and U13400 (N_13400,N_12817,N_12555);
and U13401 (N_13401,N_12974,N_12696);
and U13402 (N_13402,N_12955,N_12735);
nor U13403 (N_13403,N_12681,N_12652);
and U13404 (N_13404,N_12886,N_12953);
and U13405 (N_13405,N_12924,N_12873);
xor U13406 (N_13406,N_12647,N_12651);
nor U13407 (N_13407,N_12901,N_12778);
and U13408 (N_13408,N_12730,N_12656);
nand U13409 (N_13409,N_12635,N_12544);
nand U13410 (N_13410,N_12929,N_12514);
xor U13411 (N_13411,N_12540,N_12841);
nor U13412 (N_13412,N_12921,N_12789);
nand U13413 (N_13413,N_12721,N_12913);
or U13414 (N_13414,N_12939,N_12606);
or U13415 (N_13415,N_12604,N_12960);
nor U13416 (N_13416,N_12828,N_12932);
xnor U13417 (N_13417,N_12713,N_12721);
xor U13418 (N_13418,N_12813,N_12785);
nor U13419 (N_13419,N_12704,N_12843);
xnor U13420 (N_13420,N_12617,N_12961);
and U13421 (N_13421,N_12739,N_12552);
nand U13422 (N_13422,N_12845,N_12669);
or U13423 (N_13423,N_12884,N_12521);
xor U13424 (N_13424,N_12712,N_12666);
nor U13425 (N_13425,N_12626,N_12693);
nand U13426 (N_13426,N_12761,N_12608);
or U13427 (N_13427,N_12572,N_12960);
nand U13428 (N_13428,N_12725,N_12557);
or U13429 (N_13429,N_12775,N_12629);
nor U13430 (N_13430,N_12975,N_12574);
or U13431 (N_13431,N_12840,N_12566);
xor U13432 (N_13432,N_12769,N_12680);
nor U13433 (N_13433,N_12710,N_12886);
or U13434 (N_13434,N_12763,N_12973);
nor U13435 (N_13435,N_12558,N_12542);
xor U13436 (N_13436,N_12700,N_12941);
or U13437 (N_13437,N_12836,N_12824);
and U13438 (N_13438,N_12788,N_12632);
and U13439 (N_13439,N_12769,N_12929);
nand U13440 (N_13440,N_12654,N_12560);
and U13441 (N_13441,N_12830,N_12502);
or U13442 (N_13442,N_12884,N_12899);
nand U13443 (N_13443,N_12833,N_12682);
and U13444 (N_13444,N_12701,N_12588);
nor U13445 (N_13445,N_12526,N_12678);
xnor U13446 (N_13446,N_12964,N_12862);
and U13447 (N_13447,N_12891,N_12889);
nor U13448 (N_13448,N_12943,N_12729);
nand U13449 (N_13449,N_12795,N_12782);
nor U13450 (N_13450,N_12772,N_12784);
and U13451 (N_13451,N_12632,N_12663);
nor U13452 (N_13452,N_12610,N_12534);
and U13453 (N_13453,N_12632,N_12998);
xor U13454 (N_13454,N_12725,N_12882);
or U13455 (N_13455,N_12951,N_12735);
xnor U13456 (N_13456,N_12856,N_12767);
nand U13457 (N_13457,N_12986,N_12584);
nor U13458 (N_13458,N_12789,N_12832);
and U13459 (N_13459,N_12917,N_12683);
xor U13460 (N_13460,N_12650,N_12636);
nand U13461 (N_13461,N_12940,N_12861);
nor U13462 (N_13462,N_12772,N_12647);
xor U13463 (N_13463,N_12959,N_12720);
nand U13464 (N_13464,N_12784,N_12716);
xnor U13465 (N_13465,N_12630,N_12686);
or U13466 (N_13466,N_12939,N_12514);
nor U13467 (N_13467,N_12941,N_12785);
xor U13468 (N_13468,N_12540,N_12578);
and U13469 (N_13469,N_12507,N_12931);
nand U13470 (N_13470,N_12828,N_12838);
or U13471 (N_13471,N_12742,N_12761);
nand U13472 (N_13472,N_12592,N_12952);
xor U13473 (N_13473,N_12756,N_12893);
and U13474 (N_13474,N_12849,N_12668);
or U13475 (N_13475,N_12850,N_12821);
nor U13476 (N_13476,N_12953,N_12959);
and U13477 (N_13477,N_12811,N_12567);
nand U13478 (N_13478,N_12616,N_12505);
and U13479 (N_13479,N_12576,N_12874);
nand U13480 (N_13480,N_12654,N_12667);
nand U13481 (N_13481,N_12588,N_12674);
nor U13482 (N_13482,N_12975,N_12639);
nand U13483 (N_13483,N_12963,N_12964);
xor U13484 (N_13484,N_12827,N_12982);
xor U13485 (N_13485,N_12635,N_12785);
and U13486 (N_13486,N_12820,N_12691);
and U13487 (N_13487,N_12884,N_12584);
or U13488 (N_13488,N_12593,N_12792);
or U13489 (N_13489,N_12843,N_12654);
xnor U13490 (N_13490,N_12961,N_12873);
and U13491 (N_13491,N_12526,N_12906);
xor U13492 (N_13492,N_12673,N_12901);
or U13493 (N_13493,N_12663,N_12837);
or U13494 (N_13494,N_12985,N_12714);
or U13495 (N_13495,N_12879,N_12970);
nand U13496 (N_13496,N_12709,N_12818);
nor U13497 (N_13497,N_12632,N_12640);
and U13498 (N_13498,N_12998,N_12909);
xor U13499 (N_13499,N_12749,N_12989);
nand U13500 (N_13500,N_13287,N_13108);
and U13501 (N_13501,N_13116,N_13064);
nor U13502 (N_13502,N_13051,N_13142);
or U13503 (N_13503,N_13313,N_13053);
and U13504 (N_13504,N_13424,N_13425);
xor U13505 (N_13505,N_13411,N_13414);
and U13506 (N_13506,N_13401,N_13333);
nand U13507 (N_13507,N_13429,N_13056);
nor U13508 (N_13508,N_13303,N_13216);
xnor U13509 (N_13509,N_13473,N_13240);
xnor U13510 (N_13510,N_13081,N_13392);
xor U13511 (N_13511,N_13140,N_13006);
xnor U13512 (N_13512,N_13161,N_13422);
xnor U13513 (N_13513,N_13295,N_13267);
nand U13514 (N_13514,N_13219,N_13471);
xnor U13515 (N_13515,N_13011,N_13222);
nor U13516 (N_13516,N_13404,N_13003);
nor U13517 (N_13517,N_13171,N_13032);
xor U13518 (N_13518,N_13420,N_13399);
xnor U13519 (N_13519,N_13445,N_13463);
or U13520 (N_13520,N_13251,N_13130);
nand U13521 (N_13521,N_13403,N_13169);
xor U13522 (N_13522,N_13435,N_13364);
nor U13523 (N_13523,N_13484,N_13259);
and U13524 (N_13524,N_13211,N_13210);
and U13525 (N_13525,N_13063,N_13482);
nor U13526 (N_13526,N_13234,N_13119);
or U13527 (N_13527,N_13460,N_13481);
nand U13528 (N_13528,N_13025,N_13122);
nand U13529 (N_13529,N_13451,N_13163);
and U13530 (N_13530,N_13256,N_13237);
xnor U13531 (N_13531,N_13474,N_13136);
nand U13532 (N_13532,N_13241,N_13078);
xor U13533 (N_13533,N_13383,N_13491);
xor U13534 (N_13534,N_13490,N_13173);
and U13535 (N_13535,N_13479,N_13397);
or U13536 (N_13536,N_13348,N_13407);
xnor U13537 (N_13537,N_13191,N_13047);
nand U13538 (N_13538,N_13109,N_13209);
xnor U13539 (N_13539,N_13076,N_13027);
or U13540 (N_13540,N_13286,N_13376);
nand U13541 (N_13541,N_13325,N_13465);
nor U13542 (N_13542,N_13203,N_13280);
xor U13543 (N_13543,N_13035,N_13070);
nor U13544 (N_13544,N_13091,N_13117);
nand U13545 (N_13545,N_13049,N_13158);
and U13546 (N_13546,N_13493,N_13029);
nand U13547 (N_13547,N_13396,N_13264);
xnor U13548 (N_13548,N_13293,N_13466);
nand U13549 (N_13549,N_13436,N_13176);
nor U13550 (N_13550,N_13023,N_13265);
or U13551 (N_13551,N_13455,N_13099);
nor U13552 (N_13552,N_13012,N_13005);
nor U13553 (N_13553,N_13120,N_13339);
nand U13554 (N_13554,N_13440,N_13377);
nor U13555 (N_13555,N_13329,N_13462);
nor U13556 (N_13556,N_13446,N_13379);
nand U13557 (N_13557,N_13357,N_13456);
nand U13558 (N_13558,N_13292,N_13269);
xnor U13559 (N_13559,N_13250,N_13262);
xnor U13560 (N_13560,N_13074,N_13384);
xnor U13561 (N_13561,N_13041,N_13478);
and U13562 (N_13562,N_13139,N_13487);
nand U13563 (N_13563,N_13118,N_13268);
xnor U13564 (N_13564,N_13337,N_13288);
or U13565 (N_13565,N_13338,N_13432);
nor U13566 (N_13566,N_13363,N_13060);
or U13567 (N_13567,N_13381,N_13415);
xor U13568 (N_13568,N_13194,N_13385);
and U13569 (N_13569,N_13188,N_13245);
and U13570 (N_13570,N_13492,N_13167);
and U13571 (N_13571,N_13180,N_13152);
and U13572 (N_13572,N_13184,N_13413);
and U13573 (N_13573,N_13165,N_13495);
or U13574 (N_13574,N_13110,N_13395);
or U13575 (N_13575,N_13423,N_13405);
nor U13576 (N_13576,N_13249,N_13106);
nand U13577 (N_13577,N_13497,N_13257);
nand U13578 (N_13578,N_13092,N_13443);
or U13579 (N_13579,N_13030,N_13202);
or U13580 (N_13580,N_13274,N_13312);
nand U13581 (N_13581,N_13278,N_13208);
nand U13582 (N_13582,N_13344,N_13052);
nand U13583 (N_13583,N_13190,N_13086);
xnor U13584 (N_13584,N_13387,N_13104);
xnor U13585 (N_13585,N_13496,N_13146);
xor U13586 (N_13586,N_13282,N_13254);
or U13587 (N_13587,N_13195,N_13416);
and U13588 (N_13588,N_13024,N_13013);
nor U13589 (N_13589,N_13389,N_13393);
nor U13590 (N_13590,N_13192,N_13149);
xor U13591 (N_13591,N_13227,N_13266);
nand U13592 (N_13592,N_13458,N_13285);
xor U13593 (N_13593,N_13230,N_13138);
nand U13594 (N_13594,N_13038,N_13084);
xnor U13595 (N_13595,N_13309,N_13224);
nor U13596 (N_13596,N_13472,N_13341);
nand U13597 (N_13597,N_13353,N_13271);
xor U13598 (N_13598,N_13150,N_13143);
and U13599 (N_13599,N_13059,N_13077);
or U13600 (N_13600,N_13105,N_13225);
nand U13601 (N_13601,N_13043,N_13372);
nand U13602 (N_13602,N_13151,N_13369);
and U13603 (N_13603,N_13131,N_13419);
nand U13604 (N_13604,N_13009,N_13248);
or U13605 (N_13605,N_13002,N_13328);
and U13606 (N_13606,N_13181,N_13326);
xor U13607 (N_13607,N_13068,N_13028);
nor U13608 (N_13608,N_13065,N_13441);
or U13609 (N_13609,N_13016,N_13010);
nand U13610 (N_13610,N_13375,N_13175);
or U13611 (N_13611,N_13261,N_13449);
nand U13612 (N_13612,N_13229,N_13067);
or U13613 (N_13613,N_13489,N_13058);
and U13614 (N_13614,N_13289,N_13126);
nand U13615 (N_13615,N_13367,N_13098);
or U13616 (N_13616,N_13483,N_13217);
nand U13617 (N_13617,N_13072,N_13159);
and U13618 (N_13618,N_13121,N_13147);
nand U13619 (N_13619,N_13356,N_13400);
nor U13620 (N_13620,N_13374,N_13470);
nand U13621 (N_13621,N_13236,N_13018);
nor U13622 (N_13622,N_13370,N_13014);
xor U13623 (N_13623,N_13444,N_13362);
nand U13624 (N_13624,N_13039,N_13112);
nor U13625 (N_13625,N_13431,N_13461);
and U13626 (N_13626,N_13101,N_13457);
or U13627 (N_13627,N_13323,N_13186);
and U13628 (N_13628,N_13168,N_13214);
xor U13629 (N_13629,N_13200,N_13365);
or U13630 (N_13630,N_13132,N_13480);
nand U13631 (N_13631,N_13322,N_13307);
xnor U13632 (N_13632,N_13319,N_13223);
nand U13633 (N_13633,N_13177,N_13090);
xor U13634 (N_13634,N_13258,N_13380);
nand U13635 (N_13635,N_13426,N_13315);
and U13636 (N_13636,N_13239,N_13089);
or U13637 (N_13637,N_13127,N_13166);
xor U13638 (N_13638,N_13004,N_13113);
xnor U13639 (N_13639,N_13226,N_13438);
xor U13640 (N_13640,N_13349,N_13141);
nand U13641 (N_13641,N_13135,N_13020);
or U13642 (N_13642,N_13061,N_13097);
or U13643 (N_13643,N_13170,N_13398);
and U13644 (N_13644,N_13042,N_13125);
and U13645 (N_13645,N_13207,N_13082);
or U13646 (N_13646,N_13096,N_13442);
xor U13647 (N_13647,N_13270,N_13178);
or U13648 (N_13648,N_13001,N_13279);
xor U13649 (N_13649,N_13083,N_13342);
nor U13650 (N_13650,N_13347,N_13088);
and U13651 (N_13651,N_13154,N_13368);
xnor U13652 (N_13652,N_13201,N_13244);
and U13653 (N_13653,N_13182,N_13300);
and U13654 (N_13654,N_13459,N_13133);
xnor U13655 (N_13655,N_13253,N_13093);
or U13656 (N_13656,N_13033,N_13144);
or U13657 (N_13657,N_13187,N_13448);
nand U13658 (N_13658,N_13281,N_13304);
xnor U13659 (N_13659,N_13085,N_13447);
nand U13660 (N_13660,N_13410,N_13045);
xor U13661 (N_13661,N_13145,N_13071);
nand U13662 (N_13662,N_13475,N_13346);
xnor U13663 (N_13663,N_13046,N_13235);
or U13664 (N_13664,N_13197,N_13213);
and U13665 (N_13665,N_13102,N_13358);
or U13666 (N_13666,N_13311,N_13366);
xor U13667 (N_13667,N_13305,N_13069);
or U13668 (N_13668,N_13232,N_13382);
nand U13669 (N_13669,N_13402,N_13137);
xor U13670 (N_13670,N_13469,N_13233);
nor U13671 (N_13671,N_13094,N_13238);
and U13672 (N_13672,N_13297,N_13452);
nand U13673 (N_13673,N_13160,N_13134);
nand U13674 (N_13674,N_13324,N_13164);
nor U13675 (N_13675,N_13412,N_13277);
or U13676 (N_13676,N_13022,N_13153);
nand U13677 (N_13677,N_13428,N_13351);
nand U13678 (N_13678,N_13031,N_13345);
or U13679 (N_13679,N_13468,N_13048);
xor U13680 (N_13680,N_13100,N_13485);
and U13681 (N_13681,N_13080,N_13156);
xnor U13682 (N_13682,N_13486,N_13418);
nor U13683 (N_13683,N_13331,N_13019);
xnor U13684 (N_13684,N_13050,N_13284);
nor U13685 (N_13685,N_13212,N_13062);
or U13686 (N_13686,N_13294,N_13095);
and U13687 (N_13687,N_13488,N_13206);
xor U13688 (N_13688,N_13111,N_13057);
xnor U13689 (N_13689,N_13332,N_13196);
nand U13690 (N_13690,N_13296,N_13408);
xnor U13691 (N_13691,N_13394,N_13406);
and U13692 (N_13692,N_13198,N_13390);
nand U13693 (N_13693,N_13179,N_13476);
nand U13694 (N_13694,N_13359,N_13290);
nand U13695 (N_13695,N_13075,N_13129);
and U13696 (N_13696,N_13228,N_13157);
xnor U13697 (N_13697,N_13242,N_13283);
xor U13698 (N_13698,N_13427,N_13247);
xor U13699 (N_13699,N_13291,N_13123);
and U13700 (N_13700,N_13220,N_13308);
nand U13701 (N_13701,N_13433,N_13330);
nor U13702 (N_13702,N_13352,N_13361);
nor U13703 (N_13703,N_13318,N_13391);
nor U13704 (N_13704,N_13148,N_13464);
xor U13705 (N_13705,N_13044,N_13343);
xnor U13706 (N_13706,N_13272,N_13174);
nand U13707 (N_13707,N_13371,N_13055);
and U13708 (N_13708,N_13115,N_13040);
xor U13709 (N_13709,N_13000,N_13316);
nand U13710 (N_13710,N_13302,N_13409);
and U13711 (N_13711,N_13155,N_13355);
nor U13712 (N_13712,N_13494,N_13350);
nor U13713 (N_13713,N_13306,N_13360);
xnor U13714 (N_13714,N_13114,N_13298);
xnor U13715 (N_13715,N_13015,N_13317);
xnor U13716 (N_13716,N_13499,N_13373);
nor U13717 (N_13717,N_13036,N_13378);
nor U13718 (N_13718,N_13079,N_13189);
or U13719 (N_13719,N_13453,N_13299);
xor U13720 (N_13720,N_13386,N_13467);
nor U13721 (N_13721,N_13007,N_13434);
nand U13722 (N_13722,N_13477,N_13107);
nand U13723 (N_13723,N_13021,N_13231);
and U13724 (N_13724,N_13066,N_13437);
and U13725 (N_13725,N_13263,N_13199);
nor U13726 (N_13726,N_13275,N_13205);
and U13727 (N_13727,N_13439,N_13215);
xor U13728 (N_13728,N_13320,N_13172);
or U13729 (N_13729,N_13037,N_13301);
and U13730 (N_13730,N_13260,N_13221);
nand U13731 (N_13731,N_13314,N_13321);
nand U13732 (N_13732,N_13388,N_13310);
nand U13733 (N_13733,N_13336,N_13124);
nand U13734 (N_13734,N_13421,N_13498);
or U13735 (N_13735,N_13273,N_13162);
xor U13736 (N_13736,N_13430,N_13454);
or U13737 (N_13737,N_13026,N_13246);
xor U13738 (N_13738,N_13034,N_13008);
nor U13739 (N_13739,N_13204,N_13193);
xor U13740 (N_13740,N_13103,N_13218);
or U13741 (N_13741,N_13335,N_13276);
nand U13742 (N_13742,N_13255,N_13017);
and U13743 (N_13743,N_13327,N_13334);
xnor U13744 (N_13744,N_13252,N_13185);
nor U13745 (N_13745,N_13128,N_13183);
nor U13746 (N_13746,N_13054,N_13340);
nand U13747 (N_13747,N_13354,N_13243);
xnor U13748 (N_13748,N_13417,N_13073);
nand U13749 (N_13749,N_13450,N_13087);
and U13750 (N_13750,N_13170,N_13226);
nor U13751 (N_13751,N_13489,N_13094);
nand U13752 (N_13752,N_13345,N_13007);
nor U13753 (N_13753,N_13095,N_13262);
xor U13754 (N_13754,N_13485,N_13185);
or U13755 (N_13755,N_13059,N_13491);
and U13756 (N_13756,N_13159,N_13423);
or U13757 (N_13757,N_13138,N_13266);
or U13758 (N_13758,N_13254,N_13310);
or U13759 (N_13759,N_13230,N_13206);
and U13760 (N_13760,N_13021,N_13203);
nor U13761 (N_13761,N_13211,N_13365);
and U13762 (N_13762,N_13098,N_13059);
or U13763 (N_13763,N_13117,N_13074);
nor U13764 (N_13764,N_13380,N_13017);
or U13765 (N_13765,N_13267,N_13085);
or U13766 (N_13766,N_13482,N_13340);
nor U13767 (N_13767,N_13334,N_13405);
nand U13768 (N_13768,N_13154,N_13354);
and U13769 (N_13769,N_13188,N_13132);
nor U13770 (N_13770,N_13130,N_13391);
nand U13771 (N_13771,N_13001,N_13389);
xnor U13772 (N_13772,N_13369,N_13165);
nor U13773 (N_13773,N_13203,N_13455);
nor U13774 (N_13774,N_13492,N_13124);
or U13775 (N_13775,N_13414,N_13044);
and U13776 (N_13776,N_13460,N_13496);
nand U13777 (N_13777,N_13159,N_13249);
xor U13778 (N_13778,N_13106,N_13163);
nor U13779 (N_13779,N_13353,N_13166);
or U13780 (N_13780,N_13437,N_13112);
xor U13781 (N_13781,N_13171,N_13276);
and U13782 (N_13782,N_13473,N_13138);
nand U13783 (N_13783,N_13350,N_13377);
nor U13784 (N_13784,N_13231,N_13290);
nor U13785 (N_13785,N_13192,N_13074);
xnor U13786 (N_13786,N_13425,N_13387);
or U13787 (N_13787,N_13022,N_13200);
nand U13788 (N_13788,N_13178,N_13400);
nand U13789 (N_13789,N_13299,N_13406);
nand U13790 (N_13790,N_13002,N_13051);
and U13791 (N_13791,N_13145,N_13458);
and U13792 (N_13792,N_13369,N_13187);
or U13793 (N_13793,N_13350,N_13352);
nand U13794 (N_13794,N_13392,N_13151);
or U13795 (N_13795,N_13311,N_13017);
nand U13796 (N_13796,N_13235,N_13393);
nand U13797 (N_13797,N_13202,N_13031);
and U13798 (N_13798,N_13007,N_13300);
and U13799 (N_13799,N_13334,N_13144);
xnor U13800 (N_13800,N_13184,N_13438);
nor U13801 (N_13801,N_13465,N_13399);
nand U13802 (N_13802,N_13068,N_13111);
and U13803 (N_13803,N_13044,N_13473);
and U13804 (N_13804,N_13347,N_13111);
and U13805 (N_13805,N_13051,N_13295);
and U13806 (N_13806,N_13319,N_13455);
or U13807 (N_13807,N_13291,N_13250);
or U13808 (N_13808,N_13095,N_13057);
nand U13809 (N_13809,N_13129,N_13056);
and U13810 (N_13810,N_13287,N_13111);
and U13811 (N_13811,N_13480,N_13301);
and U13812 (N_13812,N_13323,N_13283);
or U13813 (N_13813,N_13407,N_13388);
nor U13814 (N_13814,N_13422,N_13460);
or U13815 (N_13815,N_13391,N_13472);
nand U13816 (N_13816,N_13067,N_13480);
or U13817 (N_13817,N_13353,N_13445);
nand U13818 (N_13818,N_13372,N_13079);
xnor U13819 (N_13819,N_13075,N_13438);
xnor U13820 (N_13820,N_13341,N_13226);
nor U13821 (N_13821,N_13145,N_13188);
and U13822 (N_13822,N_13197,N_13063);
nor U13823 (N_13823,N_13135,N_13105);
or U13824 (N_13824,N_13341,N_13234);
and U13825 (N_13825,N_13419,N_13183);
and U13826 (N_13826,N_13325,N_13346);
nand U13827 (N_13827,N_13122,N_13241);
or U13828 (N_13828,N_13460,N_13426);
or U13829 (N_13829,N_13110,N_13161);
nor U13830 (N_13830,N_13058,N_13322);
nor U13831 (N_13831,N_13411,N_13438);
nor U13832 (N_13832,N_13106,N_13010);
xor U13833 (N_13833,N_13472,N_13081);
or U13834 (N_13834,N_13249,N_13134);
xor U13835 (N_13835,N_13386,N_13130);
xnor U13836 (N_13836,N_13208,N_13462);
and U13837 (N_13837,N_13399,N_13491);
xnor U13838 (N_13838,N_13192,N_13326);
or U13839 (N_13839,N_13024,N_13057);
nor U13840 (N_13840,N_13304,N_13453);
nor U13841 (N_13841,N_13441,N_13395);
and U13842 (N_13842,N_13478,N_13499);
xor U13843 (N_13843,N_13223,N_13328);
nor U13844 (N_13844,N_13307,N_13328);
and U13845 (N_13845,N_13493,N_13239);
xnor U13846 (N_13846,N_13034,N_13121);
nand U13847 (N_13847,N_13232,N_13240);
and U13848 (N_13848,N_13268,N_13487);
or U13849 (N_13849,N_13011,N_13151);
nand U13850 (N_13850,N_13305,N_13254);
nand U13851 (N_13851,N_13419,N_13433);
nor U13852 (N_13852,N_13222,N_13412);
nor U13853 (N_13853,N_13430,N_13205);
xor U13854 (N_13854,N_13143,N_13220);
or U13855 (N_13855,N_13098,N_13470);
xnor U13856 (N_13856,N_13164,N_13109);
or U13857 (N_13857,N_13186,N_13071);
nor U13858 (N_13858,N_13103,N_13031);
nor U13859 (N_13859,N_13420,N_13197);
xor U13860 (N_13860,N_13340,N_13436);
and U13861 (N_13861,N_13423,N_13356);
or U13862 (N_13862,N_13232,N_13370);
and U13863 (N_13863,N_13293,N_13315);
or U13864 (N_13864,N_13466,N_13024);
nand U13865 (N_13865,N_13470,N_13299);
nor U13866 (N_13866,N_13346,N_13103);
nor U13867 (N_13867,N_13477,N_13072);
xor U13868 (N_13868,N_13364,N_13267);
nand U13869 (N_13869,N_13284,N_13037);
or U13870 (N_13870,N_13137,N_13260);
nor U13871 (N_13871,N_13132,N_13150);
or U13872 (N_13872,N_13459,N_13023);
or U13873 (N_13873,N_13108,N_13185);
nand U13874 (N_13874,N_13246,N_13012);
nor U13875 (N_13875,N_13038,N_13444);
and U13876 (N_13876,N_13065,N_13484);
nor U13877 (N_13877,N_13208,N_13331);
nor U13878 (N_13878,N_13020,N_13162);
and U13879 (N_13879,N_13055,N_13291);
nor U13880 (N_13880,N_13012,N_13015);
nand U13881 (N_13881,N_13403,N_13327);
nor U13882 (N_13882,N_13465,N_13301);
and U13883 (N_13883,N_13251,N_13047);
nand U13884 (N_13884,N_13409,N_13338);
and U13885 (N_13885,N_13143,N_13241);
nand U13886 (N_13886,N_13199,N_13160);
nand U13887 (N_13887,N_13137,N_13361);
or U13888 (N_13888,N_13433,N_13448);
xor U13889 (N_13889,N_13337,N_13107);
nor U13890 (N_13890,N_13232,N_13135);
or U13891 (N_13891,N_13256,N_13045);
or U13892 (N_13892,N_13153,N_13284);
xnor U13893 (N_13893,N_13447,N_13443);
nand U13894 (N_13894,N_13026,N_13492);
nand U13895 (N_13895,N_13039,N_13253);
nor U13896 (N_13896,N_13147,N_13170);
nor U13897 (N_13897,N_13030,N_13121);
and U13898 (N_13898,N_13034,N_13358);
or U13899 (N_13899,N_13176,N_13029);
nand U13900 (N_13900,N_13064,N_13468);
and U13901 (N_13901,N_13227,N_13192);
and U13902 (N_13902,N_13309,N_13162);
xnor U13903 (N_13903,N_13260,N_13279);
and U13904 (N_13904,N_13057,N_13468);
nand U13905 (N_13905,N_13377,N_13470);
xnor U13906 (N_13906,N_13277,N_13495);
nor U13907 (N_13907,N_13239,N_13375);
nor U13908 (N_13908,N_13452,N_13199);
xor U13909 (N_13909,N_13479,N_13136);
and U13910 (N_13910,N_13063,N_13152);
nand U13911 (N_13911,N_13138,N_13145);
and U13912 (N_13912,N_13276,N_13036);
nand U13913 (N_13913,N_13358,N_13372);
xor U13914 (N_13914,N_13176,N_13171);
and U13915 (N_13915,N_13139,N_13269);
nand U13916 (N_13916,N_13192,N_13381);
or U13917 (N_13917,N_13114,N_13006);
nand U13918 (N_13918,N_13271,N_13061);
nand U13919 (N_13919,N_13200,N_13171);
nand U13920 (N_13920,N_13249,N_13382);
nor U13921 (N_13921,N_13291,N_13256);
nor U13922 (N_13922,N_13020,N_13015);
nand U13923 (N_13923,N_13294,N_13115);
nor U13924 (N_13924,N_13336,N_13090);
nand U13925 (N_13925,N_13082,N_13168);
nor U13926 (N_13926,N_13174,N_13346);
xor U13927 (N_13927,N_13232,N_13075);
and U13928 (N_13928,N_13330,N_13408);
nand U13929 (N_13929,N_13126,N_13311);
or U13930 (N_13930,N_13253,N_13110);
nor U13931 (N_13931,N_13381,N_13244);
nor U13932 (N_13932,N_13023,N_13125);
xnor U13933 (N_13933,N_13372,N_13472);
nand U13934 (N_13934,N_13239,N_13212);
nor U13935 (N_13935,N_13062,N_13330);
and U13936 (N_13936,N_13471,N_13042);
nor U13937 (N_13937,N_13434,N_13322);
nand U13938 (N_13938,N_13038,N_13249);
and U13939 (N_13939,N_13046,N_13171);
nor U13940 (N_13940,N_13061,N_13427);
xor U13941 (N_13941,N_13196,N_13002);
xnor U13942 (N_13942,N_13143,N_13289);
and U13943 (N_13943,N_13437,N_13279);
xnor U13944 (N_13944,N_13229,N_13274);
nor U13945 (N_13945,N_13282,N_13168);
nor U13946 (N_13946,N_13301,N_13114);
xnor U13947 (N_13947,N_13435,N_13160);
nand U13948 (N_13948,N_13450,N_13014);
or U13949 (N_13949,N_13495,N_13263);
or U13950 (N_13950,N_13455,N_13467);
or U13951 (N_13951,N_13405,N_13417);
and U13952 (N_13952,N_13105,N_13282);
nand U13953 (N_13953,N_13204,N_13001);
nand U13954 (N_13954,N_13186,N_13345);
and U13955 (N_13955,N_13293,N_13342);
nand U13956 (N_13956,N_13093,N_13277);
or U13957 (N_13957,N_13457,N_13092);
xnor U13958 (N_13958,N_13218,N_13371);
xor U13959 (N_13959,N_13081,N_13062);
nand U13960 (N_13960,N_13167,N_13334);
or U13961 (N_13961,N_13049,N_13397);
nor U13962 (N_13962,N_13361,N_13243);
xnor U13963 (N_13963,N_13336,N_13346);
or U13964 (N_13964,N_13092,N_13338);
xnor U13965 (N_13965,N_13334,N_13148);
nor U13966 (N_13966,N_13036,N_13405);
nor U13967 (N_13967,N_13128,N_13394);
nand U13968 (N_13968,N_13055,N_13461);
nand U13969 (N_13969,N_13014,N_13375);
nor U13970 (N_13970,N_13140,N_13296);
nand U13971 (N_13971,N_13029,N_13318);
or U13972 (N_13972,N_13453,N_13326);
nand U13973 (N_13973,N_13462,N_13483);
and U13974 (N_13974,N_13491,N_13070);
xnor U13975 (N_13975,N_13119,N_13446);
or U13976 (N_13976,N_13073,N_13273);
or U13977 (N_13977,N_13186,N_13138);
xor U13978 (N_13978,N_13352,N_13487);
nor U13979 (N_13979,N_13360,N_13036);
nor U13980 (N_13980,N_13300,N_13447);
nand U13981 (N_13981,N_13306,N_13129);
or U13982 (N_13982,N_13123,N_13465);
nor U13983 (N_13983,N_13455,N_13206);
nor U13984 (N_13984,N_13103,N_13027);
xnor U13985 (N_13985,N_13492,N_13474);
or U13986 (N_13986,N_13260,N_13321);
and U13987 (N_13987,N_13208,N_13118);
or U13988 (N_13988,N_13265,N_13048);
and U13989 (N_13989,N_13025,N_13024);
or U13990 (N_13990,N_13151,N_13176);
nand U13991 (N_13991,N_13350,N_13356);
and U13992 (N_13992,N_13411,N_13356);
nor U13993 (N_13993,N_13206,N_13462);
xor U13994 (N_13994,N_13085,N_13130);
nand U13995 (N_13995,N_13146,N_13350);
xnor U13996 (N_13996,N_13292,N_13497);
nand U13997 (N_13997,N_13220,N_13102);
nor U13998 (N_13998,N_13356,N_13080);
xnor U13999 (N_13999,N_13420,N_13475);
or U14000 (N_14000,N_13849,N_13914);
xnor U14001 (N_14001,N_13564,N_13814);
and U14002 (N_14002,N_13944,N_13553);
or U14003 (N_14003,N_13671,N_13662);
and U14004 (N_14004,N_13781,N_13867);
xnor U14005 (N_14005,N_13659,N_13767);
or U14006 (N_14006,N_13750,N_13856);
nand U14007 (N_14007,N_13802,N_13545);
nand U14008 (N_14008,N_13576,N_13886);
nor U14009 (N_14009,N_13560,N_13890);
or U14010 (N_14010,N_13834,N_13863);
or U14011 (N_14011,N_13820,N_13971);
nand U14012 (N_14012,N_13656,N_13809);
nor U14013 (N_14013,N_13556,N_13652);
or U14014 (N_14014,N_13725,N_13512);
or U14015 (N_14015,N_13788,N_13684);
or U14016 (N_14016,N_13990,N_13633);
nor U14017 (N_14017,N_13661,N_13989);
nand U14018 (N_14018,N_13765,N_13581);
or U14019 (N_14019,N_13784,N_13951);
xnor U14020 (N_14020,N_13693,N_13689);
nand U14021 (N_14021,N_13594,N_13575);
and U14022 (N_14022,N_13598,N_13509);
nor U14023 (N_14023,N_13783,N_13739);
xnor U14024 (N_14024,N_13579,N_13715);
nand U14025 (N_14025,N_13775,N_13969);
xor U14026 (N_14026,N_13612,N_13995);
and U14027 (N_14027,N_13591,N_13694);
nor U14028 (N_14028,N_13701,N_13713);
or U14029 (N_14029,N_13621,N_13908);
nor U14030 (N_14030,N_13630,N_13976);
nand U14031 (N_14031,N_13573,N_13862);
and U14032 (N_14032,N_13720,N_13826);
or U14033 (N_14033,N_13919,N_13929);
nand U14034 (N_14034,N_13870,N_13940);
xnor U14035 (N_14035,N_13806,N_13947);
nor U14036 (N_14036,N_13972,N_13646);
and U14037 (N_14037,N_13709,N_13836);
or U14038 (N_14038,N_13687,N_13742);
and U14039 (N_14039,N_13546,N_13510);
nor U14040 (N_14040,N_13879,N_13761);
xnor U14041 (N_14041,N_13670,N_13620);
and U14042 (N_14042,N_13970,N_13839);
nand U14043 (N_14043,N_13614,N_13845);
xor U14044 (N_14044,N_13780,N_13640);
nor U14045 (N_14045,N_13736,N_13956);
nand U14046 (N_14046,N_13803,N_13801);
nand U14047 (N_14047,N_13592,N_13584);
xor U14048 (N_14048,N_13930,N_13558);
nand U14049 (N_14049,N_13619,N_13732);
nor U14050 (N_14050,N_13945,N_13854);
or U14051 (N_14051,N_13999,N_13747);
or U14052 (N_14052,N_13651,N_13571);
or U14053 (N_14053,N_13859,N_13681);
nand U14054 (N_14054,N_13757,N_13825);
xor U14055 (N_14055,N_13596,N_13899);
or U14056 (N_14056,N_13514,N_13601);
or U14057 (N_14057,N_13866,N_13695);
nand U14058 (N_14058,N_13878,N_13853);
xnor U14059 (N_14059,N_13603,N_13717);
or U14060 (N_14060,N_13962,N_13881);
nor U14061 (N_14061,N_13634,N_13738);
and U14062 (N_14062,N_13719,N_13915);
nor U14063 (N_14063,N_13602,N_13615);
and U14064 (N_14064,N_13638,N_13618);
xor U14065 (N_14065,N_13655,N_13751);
nand U14066 (N_14066,N_13843,N_13505);
nor U14067 (N_14067,N_13888,N_13683);
nor U14068 (N_14068,N_13986,N_13799);
nor U14069 (N_14069,N_13599,N_13666);
nand U14070 (N_14070,N_13743,N_13653);
or U14071 (N_14071,N_13696,N_13798);
xor U14072 (N_14072,N_13937,N_13504);
xor U14073 (N_14073,N_13844,N_13896);
nor U14074 (N_14074,N_13790,N_13658);
nand U14075 (N_14075,N_13741,N_13794);
xnor U14076 (N_14076,N_13552,N_13680);
or U14077 (N_14077,N_13549,N_13669);
nor U14078 (N_14078,N_13534,N_13570);
nand U14079 (N_14079,N_13542,N_13708);
or U14080 (N_14080,N_13964,N_13833);
nor U14081 (N_14081,N_13500,N_13622);
or U14082 (N_14082,N_13647,N_13793);
nand U14083 (N_14083,N_13916,N_13942);
xnor U14084 (N_14084,N_13627,N_13818);
and U14085 (N_14085,N_13926,N_13745);
or U14086 (N_14086,N_13918,N_13894);
xnor U14087 (N_14087,N_13768,N_13774);
and U14088 (N_14088,N_13557,N_13502);
nand U14089 (N_14089,N_13957,N_13616);
nand U14090 (N_14090,N_13513,N_13804);
nor U14091 (N_14091,N_13797,N_13786);
or U14092 (N_14092,N_13812,N_13568);
and U14093 (N_14093,N_13532,N_13731);
nor U14094 (N_14094,N_13777,N_13846);
and U14095 (N_14095,N_13993,N_13643);
nand U14096 (N_14096,N_13562,N_13764);
and U14097 (N_14097,N_13977,N_13726);
or U14098 (N_14098,N_13714,N_13855);
nand U14099 (N_14099,N_13984,N_13737);
and U14100 (N_14100,N_13850,N_13852);
nor U14101 (N_14101,N_13980,N_13882);
and U14102 (N_14102,N_13950,N_13588);
or U14103 (N_14103,N_13722,N_13838);
xnor U14104 (N_14104,N_13537,N_13858);
or U14105 (N_14105,N_13981,N_13756);
xnor U14106 (N_14106,N_13815,N_13796);
or U14107 (N_14107,N_13679,N_13928);
or U14108 (N_14108,N_13936,N_13954);
and U14109 (N_14109,N_13665,N_13938);
or U14110 (N_14110,N_13823,N_13516);
xor U14111 (N_14111,N_13831,N_13994);
xnor U14112 (N_14112,N_13718,N_13868);
and U14113 (N_14113,N_13566,N_13948);
nand U14114 (N_14114,N_13730,N_13550);
nor U14115 (N_14115,N_13567,N_13608);
or U14116 (N_14116,N_13906,N_13586);
xor U14117 (N_14117,N_13952,N_13922);
xor U14118 (N_14118,N_13527,N_13735);
and U14119 (N_14119,N_13729,N_13960);
nor U14120 (N_14120,N_13706,N_13885);
nor U14121 (N_14121,N_13985,N_13835);
xnor U14122 (N_14122,N_13606,N_13965);
xnor U14123 (N_14123,N_13744,N_13685);
xor U14124 (N_14124,N_13590,N_13934);
or U14125 (N_14125,N_13779,N_13975);
nand U14126 (N_14126,N_13626,N_13880);
and U14127 (N_14127,N_13789,N_13595);
nand U14128 (N_14128,N_13829,N_13958);
and U14129 (N_14129,N_13808,N_13526);
nand U14130 (N_14130,N_13507,N_13773);
or U14131 (N_14131,N_13587,N_13724);
or U14132 (N_14132,N_13766,N_13759);
xor U14133 (N_14133,N_13518,N_13521);
xor U14134 (N_14134,N_13536,N_13538);
nor U14135 (N_14135,N_13522,N_13541);
and U14136 (N_14136,N_13664,N_13700);
nand U14137 (N_14137,N_13607,N_13668);
nand U14138 (N_14138,N_13821,N_13749);
nand U14139 (N_14139,N_13963,N_13923);
nand U14140 (N_14140,N_13710,N_13876);
and U14141 (N_14141,N_13520,N_13811);
and U14142 (N_14142,N_13941,N_13682);
or U14143 (N_14143,N_13924,N_13686);
and U14144 (N_14144,N_13597,N_13887);
xor U14145 (N_14145,N_13611,N_13905);
and U14146 (N_14146,N_13840,N_13582);
nand U14147 (N_14147,N_13525,N_13645);
and U14148 (N_14148,N_13654,N_13589);
nand U14149 (N_14149,N_13988,N_13569);
nor U14150 (N_14150,N_13540,N_13657);
and U14151 (N_14151,N_13943,N_13555);
and U14152 (N_14152,N_13996,N_13883);
xor U14153 (N_14153,N_13872,N_13810);
nor U14154 (N_14154,N_13754,N_13974);
and U14155 (N_14155,N_13782,N_13968);
and U14156 (N_14156,N_13580,N_13966);
nor U14157 (N_14157,N_13642,N_13605);
xnor U14158 (N_14158,N_13979,N_13644);
or U14159 (N_14159,N_13959,N_13753);
and U14160 (N_14160,N_13508,N_13830);
nand U14161 (N_14161,N_13932,N_13763);
nor U14162 (N_14162,N_13698,N_13703);
or U14163 (N_14163,N_13551,N_13842);
nor U14164 (N_14164,N_13559,N_13901);
and U14165 (N_14165,N_13561,N_13690);
nor U14166 (N_14166,N_13746,N_13639);
and U14167 (N_14167,N_13857,N_13841);
xor U14168 (N_14168,N_13921,N_13824);
nand U14169 (N_14169,N_13624,N_13702);
or U14170 (N_14170,N_13998,N_13748);
and U14171 (N_14171,N_13813,N_13641);
nand U14172 (N_14172,N_13903,N_13667);
xor U14173 (N_14173,N_13544,N_13931);
and U14174 (N_14174,N_13727,N_13913);
xor U14175 (N_14175,N_13832,N_13828);
or U14176 (N_14176,N_13851,N_13819);
nand U14177 (N_14177,N_13517,N_13623);
nand U14178 (N_14178,N_13891,N_13762);
nor U14179 (N_14179,N_13752,N_13902);
or U14180 (N_14180,N_13791,N_13983);
or U14181 (N_14181,N_13503,N_13673);
nor U14182 (N_14182,N_13528,N_13600);
or U14183 (N_14183,N_13860,N_13704);
nor U14184 (N_14184,N_13933,N_13678);
xnor U14185 (N_14185,N_13795,N_13917);
xor U14186 (N_14186,N_13547,N_13707);
xor U14187 (N_14187,N_13873,N_13712);
xnor U14188 (N_14188,N_13519,N_13939);
xor U14189 (N_14189,N_13617,N_13716);
or U14190 (N_14190,N_13897,N_13613);
nand U14191 (N_14191,N_13884,N_13877);
xnor U14192 (N_14192,N_13721,N_13827);
nand U14193 (N_14193,N_13817,N_13609);
nand U14194 (N_14194,N_13530,N_13875);
and U14195 (N_14195,N_13900,N_13847);
or U14196 (N_14196,N_13637,N_13848);
nand U14197 (N_14197,N_13593,N_13676);
nand U14198 (N_14198,N_13524,N_13535);
nor U14199 (N_14199,N_13604,N_13663);
nand U14200 (N_14200,N_13805,N_13991);
and U14201 (N_14201,N_13515,N_13692);
nand U14202 (N_14202,N_13792,N_13501);
nand U14203 (N_14203,N_13800,N_13740);
nor U14204 (N_14204,N_13649,N_13769);
xor U14205 (N_14205,N_13911,N_13961);
nand U14206 (N_14206,N_13978,N_13892);
nand U14207 (N_14207,N_13785,N_13955);
nor U14208 (N_14208,N_13699,N_13688);
or U14209 (N_14209,N_13889,N_13864);
nor U14210 (N_14210,N_13771,N_13992);
xnor U14211 (N_14211,N_13760,N_13997);
and U14212 (N_14212,N_13973,N_13631);
nor U14213 (N_14213,N_13565,N_13787);
nor U14214 (N_14214,N_13660,N_13728);
nor U14215 (N_14215,N_13946,N_13907);
xor U14216 (N_14216,N_13904,N_13577);
nand U14217 (N_14217,N_13629,N_13861);
nor U14218 (N_14218,N_13628,N_13987);
nor U14219 (N_14219,N_13935,N_13648);
nor U14220 (N_14220,N_13982,N_13672);
nor U14221 (N_14221,N_13554,N_13927);
nand U14222 (N_14222,N_13563,N_13636);
and U14223 (N_14223,N_13572,N_13920);
xnor U14224 (N_14224,N_13531,N_13755);
or U14225 (N_14225,N_13677,N_13691);
nand U14226 (N_14226,N_13865,N_13871);
xnor U14227 (N_14227,N_13837,N_13778);
nand U14228 (N_14228,N_13893,N_13583);
nand U14229 (N_14229,N_13529,N_13711);
or U14230 (N_14230,N_13625,N_13539);
or U14231 (N_14231,N_13953,N_13898);
or U14232 (N_14232,N_13675,N_13807);
xor U14233 (N_14233,N_13967,N_13734);
nand U14234 (N_14234,N_13650,N_13610);
nand U14235 (N_14235,N_13733,N_13697);
nor U14236 (N_14236,N_13772,N_13705);
and U14237 (N_14237,N_13895,N_13822);
or U14238 (N_14238,N_13506,N_13869);
and U14239 (N_14239,N_13543,N_13635);
nand U14240 (N_14240,N_13533,N_13770);
nand U14241 (N_14241,N_13925,N_13912);
nor U14242 (N_14242,N_13776,N_13758);
xnor U14243 (N_14243,N_13548,N_13909);
nand U14244 (N_14244,N_13723,N_13523);
nand U14245 (N_14245,N_13585,N_13674);
or U14246 (N_14246,N_13949,N_13511);
xnor U14247 (N_14247,N_13874,N_13632);
nor U14248 (N_14248,N_13578,N_13910);
nand U14249 (N_14249,N_13816,N_13574);
nand U14250 (N_14250,N_13605,N_13844);
and U14251 (N_14251,N_13771,N_13856);
or U14252 (N_14252,N_13725,N_13959);
nor U14253 (N_14253,N_13658,N_13679);
nor U14254 (N_14254,N_13592,N_13990);
xnor U14255 (N_14255,N_13818,N_13728);
nor U14256 (N_14256,N_13775,N_13829);
nor U14257 (N_14257,N_13793,N_13973);
xor U14258 (N_14258,N_13809,N_13939);
xnor U14259 (N_14259,N_13564,N_13687);
or U14260 (N_14260,N_13935,N_13612);
nand U14261 (N_14261,N_13968,N_13681);
and U14262 (N_14262,N_13593,N_13534);
nand U14263 (N_14263,N_13918,N_13904);
and U14264 (N_14264,N_13879,N_13707);
nor U14265 (N_14265,N_13915,N_13931);
nand U14266 (N_14266,N_13686,N_13884);
xor U14267 (N_14267,N_13553,N_13801);
or U14268 (N_14268,N_13717,N_13530);
xor U14269 (N_14269,N_13636,N_13854);
or U14270 (N_14270,N_13531,N_13561);
and U14271 (N_14271,N_13861,N_13854);
nor U14272 (N_14272,N_13672,N_13881);
nand U14273 (N_14273,N_13781,N_13537);
nor U14274 (N_14274,N_13741,N_13960);
nand U14275 (N_14275,N_13992,N_13717);
and U14276 (N_14276,N_13683,N_13839);
and U14277 (N_14277,N_13979,N_13759);
nor U14278 (N_14278,N_13735,N_13650);
xnor U14279 (N_14279,N_13892,N_13767);
and U14280 (N_14280,N_13864,N_13854);
nand U14281 (N_14281,N_13580,N_13726);
nand U14282 (N_14282,N_13944,N_13873);
xnor U14283 (N_14283,N_13809,N_13678);
nand U14284 (N_14284,N_13789,N_13629);
and U14285 (N_14285,N_13849,N_13923);
nand U14286 (N_14286,N_13771,N_13999);
nand U14287 (N_14287,N_13581,N_13959);
xnor U14288 (N_14288,N_13834,N_13518);
xor U14289 (N_14289,N_13601,N_13518);
or U14290 (N_14290,N_13995,N_13883);
xor U14291 (N_14291,N_13597,N_13743);
and U14292 (N_14292,N_13555,N_13773);
nand U14293 (N_14293,N_13704,N_13911);
xnor U14294 (N_14294,N_13804,N_13566);
nand U14295 (N_14295,N_13901,N_13932);
nor U14296 (N_14296,N_13818,N_13770);
nand U14297 (N_14297,N_13559,N_13797);
or U14298 (N_14298,N_13575,N_13858);
nand U14299 (N_14299,N_13665,N_13955);
nor U14300 (N_14300,N_13973,N_13502);
nand U14301 (N_14301,N_13855,N_13946);
xnor U14302 (N_14302,N_13823,N_13762);
xnor U14303 (N_14303,N_13912,N_13755);
and U14304 (N_14304,N_13569,N_13961);
and U14305 (N_14305,N_13667,N_13545);
xor U14306 (N_14306,N_13781,N_13914);
nand U14307 (N_14307,N_13812,N_13729);
nand U14308 (N_14308,N_13793,N_13577);
nor U14309 (N_14309,N_13560,N_13668);
and U14310 (N_14310,N_13525,N_13914);
or U14311 (N_14311,N_13730,N_13879);
nor U14312 (N_14312,N_13835,N_13913);
xor U14313 (N_14313,N_13718,N_13500);
xnor U14314 (N_14314,N_13892,N_13504);
nor U14315 (N_14315,N_13923,N_13723);
nand U14316 (N_14316,N_13544,N_13915);
and U14317 (N_14317,N_13645,N_13817);
xnor U14318 (N_14318,N_13874,N_13627);
nor U14319 (N_14319,N_13541,N_13908);
and U14320 (N_14320,N_13958,N_13825);
and U14321 (N_14321,N_13594,N_13545);
or U14322 (N_14322,N_13881,N_13870);
xnor U14323 (N_14323,N_13551,N_13671);
nand U14324 (N_14324,N_13651,N_13863);
and U14325 (N_14325,N_13536,N_13966);
xor U14326 (N_14326,N_13874,N_13757);
xor U14327 (N_14327,N_13961,N_13694);
xor U14328 (N_14328,N_13695,N_13706);
xnor U14329 (N_14329,N_13762,N_13720);
nor U14330 (N_14330,N_13718,N_13698);
nand U14331 (N_14331,N_13741,N_13909);
or U14332 (N_14332,N_13793,N_13983);
or U14333 (N_14333,N_13853,N_13905);
xnor U14334 (N_14334,N_13773,N_13512);
nand U14335 (N_14335,N_13726,N_13708);
or U14336 (N_14336,N_13632,N_13841);
xnor U14337 (N_14337,N_13607,N_13920);
xor U14338 (N_14338,N_13589,N_13754);
xnor U14339 (N_14339,N_13579,N_13588);
or U14340 (N_14340,N_13607,N_13667);
nor U14341 (N_14341,N_13595,N_13630);
nor U14342 (N_14342,N_13912,N_13548);
xor U14343 (N_14343,N_13845,N_13920);
or U14344 (N_14344,N_13539,N_13810);
and U14345 (N_14345,N_13605,N_13606);
or U14346 (N_14346,N_13575,N_13943);
and U14347 (N_14347,N_13986,N_13704);
nor U14348 (N_14348,N_13748,N_13944);
nor U14349 (N_14349,N_13816,N_13993);
or U14350 (N_14350,N_13680,N_13800);
xnor U14351 (N_14351,N_13581,N_13580);
or U14352 (N_14352,N_13822,N_13761);
nor U14353 (N_14353,N_13660,N_13628);
nand U14354 (N_14354,N_13885,N_13675);
nand U14355 (N_14355,N_13875,N_13746);
xnor U14356 (N_14356,N_13702,N_13594);
or U14357 (N_14357,N_13841,N_13548);
nor U14358 (N_14358,N_13581,N_13713);
nor U14359 (N_14359,N_13971,N_13829);
nand U14360 (N_14360,N_13834,N_13917);
nand U14361 (N_14361,N_13960,N_13914);
nand U14362 (N_14362,N_13571,N_13815);
nand U14363 (N_14363,N_13981,N_13613);
nor U14364 (N_14364,N_13877,N_13904);
and U14365 (N_14365,N_13816,N_13850);
nor U14366 (N_14366,N_13716,N_13918);
and U14367 (N_14367,N_13954,N_13698);
or U14368 (N_14368,N_13976,N_13911);
nor U14369 (N_14369,N_13869,N_13925);
and U14370 (N_14370,N_13973,N_13503);
xor U14371 (N_14371,N_13512,N_13821);
nand U14372 (N_14372,N_13790,N_13635);
xor U14373 (N_14373,N_13990,N_13676);
xnor U14374 (N_14374,N_13664,N_13612);
nor U14375 (N_14375,N_13706,N_13815);
nor U14376 (N_14376,N_13693,N_13646);
or U14377 (N_14377,N_13571,N_13864);
or U14378 (N_14378,N_13859,N_13663);
nand U14379 (N_14379,N_13668,N_13784);
nor U14380 (N_14380,N_13727,N_13776);
or U14381 (N_14381,N_13665,N_13608);
or U14382 (N_14382,N_13765,N_13678);
xnor U14383 (N_14383,N_13655,N_13558);
or U14384 (N_14384,N_13949,N_13602);
nor U14385 (N_14385,N_13550,N_13583);
and U14386 (N_14386,N_13817,N_13691);
or U14387 (N_14387,N_13750,N_13960);
and U14388 (N_14388,N_13607,N_13996);
nor U14389 (N_14389,N_13627,N_13966);
and U14390 (N_14390,N_13873,N_13872);
and U14391 (N_14391,N_13554,N_13793);
or U14392 (N_14392,N_13883,N_13882);
and U14393 (N_14393,N_13882,N_13634);
xnor U14394 (N_14394,N_13981,N_13537);
and U14395 (N_14395,N_13527,N_13985);
nor U14396 (N_14396,N_13963,N_13897);
xnor U14397 (N_14397,N_13780,N_13631);
and U14398 (N_14398,N_13645,N_13832);
and U14399 (N_14399,N_13774,N_13784);
and U14400 (N_14400,N_13680,N_13666);
and U14401 (N_14401,N_13951,N_13530);
or U14402 (N_14402,N_13508,N_13775);
and U14403 (N_14403,N_13905,N_13966);
or U14404 (N_14404,N_13997,N_13919);
nor U14405 (N_14405,N_13777,N_13764);
nor U14406 (N_14406,N_13647,N_13537);
nand U14407 (N_14407,N_13609,N_13893);
and U14408 (N_14408,N_13609,N_13542);
or U14409 (N_14409,N_13613,N_13710);
nor U14410 (N_14410,N_13923,N_13953);
nor U14411 (N_14411,N_13521,N_13795);
nor U14412 (N_14412,N_13931,N_13516);
xnor U14413 (N_14413,N_13722,N_13517);
nand U14414 (N_14414,N_13851,N_13922);
nor U14415 (N_14415,N_13784,N_13681);
nor U14416 (N_14416,N_13766,N_13633);
xnor U14417 (N_14417,N_13864,N_13893);
and U14418 (N_14418,N_13820,N_13645);
or U14419 (N_14419,N_13530,N_13802);
or U14420 (N_14420,N_13925,N_13934);
nor U14421 (N_14421,N_13515,N_13928);
and U14422 (N_14422,N_13524,N_13816);
xnor U14423 (N_14423,N_13718,N_13934);
xor U14424 (N_14424,N_13868,N_13958);
nand U14425 (N_14425,N_13772,N_13760);
or U14426 (N_14426,N_13721,N_13708);
nand U14427 (N_14427,N_13591,N_13663);
or U14428 (N_14428,N_13732,N_13839);
and U14429 (N_14429,N_13694,N_13681);
and U14430 (N_14430,N_13793,N_13537);
xor U14431 (N_14431,N_13797,N_13831);
nand U14432 (N_14432,N_13976,N_13562);
and U14433 (N_14433,N_13892,N_13712);
nand U14434 (N_14434,N_13879,N_13556);
nand U14435 (N_14435,N_13860,N_13515);
nand U14436 (N_14436,N_13935,N_13944);
xnor U14437 (N_14437,N_13605,N_13835);
or U14438 (N_14438,N_13718,N_13666);
or U14439 (N_14439,N_13992,N_13723);
nand U14440 (N_14440,N_13528,N_13898);
and U14441 (N_14441,N_13512,N_13573);
xor U14442 (N_14442,N_13932,N_13773);
or U14443 (N_14443,N_13746,N_13939);
and U14444 (N_14444,N_13597,N_13547);
xor U14445 (N_14445,N_13625,N_13940);
xor U14446 (N_14446,N_13870,N_13926);
and U14447 (N_14447,N_13777,N_13932);
nor U14448 (N_14448,N_13957,N_13798);
and U14449 (N_14449,N_13595,N_13544);
or U14450 (N_14450,N_13660,N_13897);
nor U14451 (N_14451,N_13904,N_13856);
or U14452 (N_14452,N_13748,N_13740);
xnor U14453 (N_14453,N_13691,N_13883);
nor U14454 (N_14454,N_13796,N_13874);
xnor U14455 (N_14455,N_13906,N_13560);
nand U14456 (N_14456,N_13898,N_13601);
or U14457 (N_14457,N_13580,N_13546);
nand U14458 (N_14458,N_13795,N_13865);
xnor U14459 (N_14459,N_13580,N_13919);
or U14460 (N_14460,N_13909,N_13631);
and U14461 (N_14461,N_13605,N_13688);
and U14462 (N_14462,N_13950,N_13511);
and U14463 (N_14463,N_13966,N_13780);
xnor U14464 (N_14464,N_13602,N_13945);
and U14465 (N_14465,N_13926,N_13619);
and U14466 (N_14466,N_13696,N_13603);
or U14467 (N_14467,N_13957,N_13964);
nand U14468 (N_14468,N_13626,N_13658);
and U14469 (N_14469,N_13874,N_13962);
or U14470 (N_14470,N_13544,N_13503);
or U14471 (N_14471,N_13604,N_13565);
nand U14472 (N_14472,N_13670,N_13827);
xnor U14473 (N_14473,N_13997,N_13900);
nand U14474 (N_14474,N_13611,N_13622);
or U14475 (N_14475,N_13543,N_13697);
nor U14476 (N_14476,N_13507,N_13541);
nor U14477 (N_14477,N_13715,N_13697);
or U14478 (N_14478,N_13746,N_13895);
xnor U14479 (N_14479,N_13592,N_13942);
and U14480 (N_14480,N_13893,N_13871);
nand U14481 (N_14481,N_13942,N_13660);
xor U14482 (N_14482,N_13549,N_13589);
or U14483 (N_14483,N_13858,N_13748);
nor U14484 (N_14484,N_13686,N_13776);
nor U14485 (N_14485,N_13863,N_13749);
nand U14486 (N_14486,N_13785,N_13681);
nand U14487 (N_14487,N_13775,N_13618);
nor U14488 (N_14488,N_13902,N_13849);
xor U14489 (N_14489,N_13752,N_13686);
nand U14490 (N_14490,N_13853,N_13931);
nor U14491 (N_14491,N_13559,N_13535);
and U14492 (N_14492,N_13748,N_13592);
and U14493 (N_14493,N_13909,N_13673);
and U14494 (N_14494,N_13906,N_13942);
nand U14495 (N_14495,N_13615,N_13817);
nor U14496 (N_14496,N_13665,N_13767);
nand U14497 (N_14497,N_13997,N_13842);
nor U14498 (N_14498,N_13842,N_13726);
and U14499 (N_14499,N_13778,N_13576);
nand U14500 (N_14500,N_14498,N_14380);
and U14501 (N_14501,N_14054,N_14001);
xnor U14502 (N_14502,N_14475,N_14157);
and U14503 (N_14503,N_14269,N_14360);
or U14504 (N_14504,N_14108,N_14385);
and U14505 (N_14505,N_14388,N_14201);
and U14506 (N_14506,N_14392,N_14373);
nand U14507 (N_14507,N_14186,N_14184);
nor U14508 (N_14508,N_14488,N_14248);
xnor U14509 (N_14509,N_14456,N_14403);
or U14510 (N_14510,N_14176,N_14436);
nand U14511 (N_14511,N_14073,N_14194);
nor U14512 (N_14512,N_14361,N_14134);
and U14513 (N_14513,N_14152,N_14441);
nand U14514 (N_14514,N_14449,N_14314);
or U14515 (N_14515,N_14442,N_14323);
nor U14516 (N_14516,N_14247,N_14092);
nor U14517 (N_14517,N_14187,N_14325);
xnor U14518 (N_14518,N_14082,N_14408);
and U14519 (N_14519,N_14457,N_14034);
nor U14520 (N_14520,N_14133,N_14103);
and U14521 (N_14521,N_14478,N_14274);
nor U14522 (N_14522,N_14149,N_14026);
and U14523 (N_14523,N_14094,N_14292);
and U14524 (N_14524,N_14017,N_14287);
and U14525 (N_14525,N_14452,N_14422);
nor U14526 (N_14526,N_14341,N_14443);
xnor U14527 (N_14527,N_14455,N_14322);
nand U14528 (N_14528,N_14178,N_14407);
and U14529 (N_14529,N_14379,N_14420);
and U14530 (N_14530,N_14047,N_14042);
and U14531 (N_14531,N_14020,N_14437);
nand U14532 (N_14532,N_14291,N_14007);
or U14533 (N_14533,N_14353,N_14041);
xor U14534 (N_14534,N_14162,N_14175);
and U14535 (N_14535,N_14354,N_14044);
xor U14536 (N_14536,N_14210,N_14172);
nor U14537 (N_14537,N_14473,N_14096);
xor U14538 (N_14538,N_14124,N_14273);
nor U14539 (N_14539,N_14004,N_14363);
or U14540 (N_14540,N_14435,N_14290);
nor U14541 (N_14541,N_14352,N_14233);
or U14542 (N_14542,N_14153,N_14382);
and U14543 (N_14543,N_14261,N_14396);
or U14544 (N_14544,N_14340,N_14107);
xor U14545 (N_14545,N_14119,N_14177);
nor U14546 (N_14546,N_14234,N_14327);
nand U14547 (N_14547,N_14220,N_14052);
and U14548 (N_14548,N_14029,N_14083);
or U14549 (N_14549,N_14114,N_14245);
xnor U14550 (N_14550,N_14458,N_14196);
nor U14551 (N_14551,N_14242,N_14057);
xnor U14552 (N_14552,N_14275,N_14333);
and U14553 (N_14553,N_14204,N_14117);
and U14554 (N_14554,N_14021,N_14019);
nor U14555 (N_14555,N_14069,N_14470);
xor U14556 (N_14556,N_14421,N_14135);
and U14557 (N_14557,N_14123,N_14072);
nand U14558 (N_14558,N_14148,N_14387);
and U14559 (N_14559,N_14100,N_14008);
nor U14560 (N_14560,N_14237,N_14180);
and U14561 (N_14561,N_14058,N_14466);
nor U14562 (N_14562,N_14376,N_14075);
and U14563 (N_14563,N_14329,N_14131);
and U14564 (N_14564,N_14336,N_14143);
and U14565 (N_14565,N_14005,N_14055);
xor U14566 (N_14566,N_14032,N_14413);
nor U14567 (N_14567,N_14426,N_14334);
and U14568 (N_14568,N_14061,N_14332);
or U14569 (N_14569,N_14289,N_14159);
xor U14570 (N_14570,N_14451,N_14218);
xnor U14571 (N_14571,N_14091,N_14030);
nand U14572 (N_14572,N_14056,N_14105);
nand U14573 (N_14573,N_14424,N_14390);
nor U14574 (N_14574,N_14499,N_14307);
xnor U14575 (N_14575,N_14039,N_14038);
and U14576 (N_14576,N_14465,N_14067);
xor U14577 (N_14577,N_14080,N_14397);
or U14578 (N_14578,N_14348,N_14406);
or U14579 (N_14579,N_14139,N_14484);
nand U14580 (N_14580,N_14110,N_14367);
or U14581 (N_14581,N_14163,N_14267);
and U14582 (N_14582,N_14433,N_14182);
nor U14583 (N_14583,N_14491,N_14192);
xnor U14584 (N_14584,N_14012,N_14104);
xnor U14585 (N_14585,N_14324,N_14285);
or U14586 (N_14586,N_14035,N_14338);
nor U14587 (N_14587,N_14320,N_14399);
nand U14588 (N_14588,N_14253,N_14010);
nor U14589 (N_14589,N_14350,N_14339);
or U14590 (N_14590,N_14479,N_14276);
or U14591 (N_14591,N_14393,N_14126);
or U14592 (N_14592,N_14115,N_14223);
and U14593 (N_14593,N_14137,N_14239);
xor U14594 (N_14594,N_14489,N_14212);
xnor U14595 (N_14595,N_14427,N_14065);
nor U14596 (N_14596,N_14068,N_14154);
and U14597 (N_14597,N_14369,N_14402);
or U14598 (N_14598,N_14036,N_14444);
and U14599 (N_14599,N_14174,N_14481);
and U14600 (N_14600,N_14270,N_14089);
nand U14601 (N_14601,N_14351,N_14303);
and U14602 (N_14602,N_14404,N_14425);
nor U14603 (N_14603,N_14265,N_14193);
and U14604 (N_14604,N_14011,N_14249);
nand U14605 (N_14605,N_14130,N_14118);
xor U14606 (N_14606,N_14372,N_14308);
nor U14607 (N_14607,N_14293,N_14202);
or U14608 (N_14608,N_14485,N_14281);
nand U14609 (N_14609,N_14326,N_14099);
nor U14610 (N_14610,N_14195,N_14469);
and U14611 (N_14611,N_14347,N_14410);
xnor U14612 (N_14612,N_14145,N_14496);
and U14613 (N_14613,N_14302,N_14160);
xor U14614 (N_14614,N_14200,N_14025);
nor U14615 (N_14615,N_14411,N_14389);
nand U14616 (N_14616,N_14279,N_14310);
nor U14617 (N_14617,N_14282,N_14171);
nor U14618 (N_14618,N_14400,N_14227);
xnor U14619 (N_14619,N_14024,N_14098);
and U14620 (N_14620,N_14037,N_14450);
nor U14621 (N_14621,N_14417,N_14432);
or U14622 (N_14622,N_14043,N_14431);
xor U14623 (N_14623,N_14088,N_14474);
or U14624 (N_14624,N_14283,N_14191);
or U14625 (N_14625,N_14295,N_14365);
and U14626 (N_14626,N_14045,N_14482);
or U14627 (N_14627,N_14070,N_14125);
or U14628 (N_14628,N_14492,N_14483);
or U14629 (N_14629,N_14121,N_14093);
xor U14630 (N_14630,N_14066,N_14102);
and U14631 (N_14631,N_14120,N_14357);
and U14632 (N_14632,N_14003,N_14216);
or U14633 (N_14633,N_14079,N_14053);
and U14634 (N_14634,N_14028,N_14151);
nand U14635 (N_14635,N_14240,N_14301);
nand U14636 (N_14636,N_14471,N_14343);
or U14637 (N_14637,N_14198,N_14230);
nand U14638 (N_14638,N_14048,N_14147);
xnor U14639 (N_14639,N_14023,N_14467);
or U14640 (N_14640,N_14002,N_14183);
xnor U14641 (N_14641,N_14490,N_14359);
nor U14642 (N_14642,N_14246,N_14062);
xnor U14643 (N_14643,N_14236,N_14296);
nor U14644 (N_14644,N_14084,N_14430);
nor U14645 (N_14645,N_14087,N_14375);
nor U14646 (N_14646,N_14181,N_14000);
or U14647 (N_14647,N_14486,N_14132);
nor U14648 (N_14648,N_14169,N_14342);
and U14649 (N_14649,N_14112,N_14311);
nor U14650 (N_14650,N_14356,N_14166);
or U14651 (N_14651,N_14221,N_14262);
xnor U14652 (N_14652,N_14304,N_14146);
or U14653 (N_14653,N_14378,N_14286);
and U14654 (N_14654,N_14497,N_14277);
nand U14655 (N_14655,N_14167,N_14271);
or U14656 (N_14656,N_14031,N_14016);
nor U14657 (N_14657,N_14266,N_14232);
and U14658 (N_14658,N_14377,N_14063);
and U14659 (N_14659,N_14416,N_14165);
nor U14660 (N_14660,N_14051,N_14368);
xor U14661 (N_14661,N_14476,N_14086);
or U14662 (N_14662,N_14257,N_14203);
nor U14663 (N_14663,N_14013,N_14009);
and U14664 (N_14664,N_14472,N_14229);
xor U14665 (N_14665,N_14337,N_14164);
nand U14666 (N_14666,N_14040,N_14190);
nand U14667 (N_14667,N_14254,N_14280);
nor U14668 (N_14668,N_14453,N_14033);
and U14669 (N_14669,N_14116,N_14170);
nor U14670 (N_14670,N_14459,N_14468);
and U14671 (N_14671,N_14440,N_14462);
and U14672 (N_14672,N_14208,N_14409);
and U14673 (N_14673,N_14022,N_14129);
nand U14674 (N_14674,N_14331,N_14217);
xnor U14675 (N_14675,N_14150,N_14315);
or U14676 (N_14676,N_14423,N_14255);
nor U14677 (N_14677,N_14398,N_14386);
nor U14678 (N_14678,N_14142,N_14414);
xor U14679 (N_14679,N_14077,N_14394);
xnor U14680 (N_14680,N_14074,N_14081);
xor U14681 (N_14681,N_14412,N_14213);
and U14682 (N_14682,N_14140,N_14345);
nand U14683 (N_14683,N_14370,N_14321);
and U14684 (N_14684,N_14439,N_14278);
nor U14685 (N_14685,N_14260,N_14224);
nor U14686 (N_14686,N_14298,N_14109);
nand U14687 (N_14687,N_14155,N_14346);
nor U14688 (N_14688,N_14374,N_14349);
nor U14689 (N_14689,N_14128,N_14014);
and U14690 (N_14690,N_14328,N_14294);
nand U14691 (N_14691,N_14018,N_14306);
nand U14692 (N_14692,N_14252,N_14446);
nand U14693 (N_14693,N_14335,N_14391);
or U14694 (N_14694,N_14447,N_14251);
nor U14695 (N_14695,N_14330,N_14144);
or U14696 (N_14696,N_14111,N_14222);
and U14697 (N_14697,N_14384,N_14078);
and U14698 (N_14698,N_14318,N_14197);
xnor U14699 (N_14699,N_14460,N_14226);
nor U14700 (N_14700,N_14272,N_14006);
nor U14701 (N_14701,N_14136,N_14173);
nor U14702 (N_14702,N_14015,N_14059);
nand U14703 (N_14703,N_14415,N_14071);
and U14704 (N_14704,N_14429,N_14156);
nand U14705 (N_14705,N_14316,N_14214);
xnor U14706 (N_14706,N_14185,N_14258);
xnor U14707 (N_14707,N_14264,N_14445);
or U14708 (N_14708,N_14487,N_14313);
nand U14709 (N_14709,N_14209,N_14463);
nor U14710 (N_14710,N_14179,N_14494);
xnor U14711 (N_14711,N_14064,N_14161);
nor U14712 (N_14712,N_14493,N_14219);
nor U14713 (N_14713,N_14418,N_14480);
and U14714 (N_14714,N_14122,N_14231);
or U14715 (N_14715,N_14309,N_14250);
nand U14716 (N_14716,N_14027,N_14188);
and U14717 (N_14717,N_14215,N_14383);
and U14718 (N_14718,N_14419,N_14095);
nor U14719 (N_14719,N_14395,N_14464);
nor U14720 (N_14720,N_14060,N_14050);
and U14721 (N_14721,N_14243,N_14381);
and U14722 (N_14722,N_14362,N_14299);
or U14723 (N_14723,N_14244,N_14205);
nand U14724 (N_14724,N_14312,N_14238);
nand U14725 (N_14725,N_14113,N_14358);
or U14726 (N_14726,N_14235,N_14206);
nor U14727 (N_14727,N_14461,N_14207);
or U14728 (N_14728,N_14259,N_14495);
or U14729 (N_14729,N_14371,N_14090);
nor U14730 (N_14730,N_14284,N_14438);
xor U14731 (N_14731,N_14097,N_14241);
xor U14732 (N_14732,N_14288,N_14199);
and U14733 (N_14733,N_14355,N_14138);
and U14734 (N_14734,N_14300,N_14085);
or U14735 (N_14735,N_14305,N_14106);
nor U14736 (N_14736,N_14401,N_14428);
nand U14737 (N_14737,N_14263,N_14344);
nor U14738 (N_14738,N_14319,N_14448);
and U14739 (N_14739,N_14101,N_14256);
or U14740 (N_14740,N_14366,N_14434);
and U14741 (N_14741,N_14076,N_14127);
nor U14742 (N_14742,N_14317,N_14225);
nand U14743 (N_14743,N_14189,N_14158);
or U14744 (N_14744,N_14364,N_14228);
and U14745 (N_14745,N_14046,N_14454);
or U14746 (N_14746,N_14477,N_14297);
nand U14747 (N_14747,N_14049,N_14268);
nand U14748 (N_14748,N_14211,N_14405);
and U14749 (N_14749,N_14141,N_14168);
and U14750 (N_14750,N_14422,N_14220);
nor U14751 (N_14751,N_14199,N_14347);
nand U14752 (N_14752,N_14416,N_14375);
or U14753 (N_14753,N_14362,N_14497);
nor U14754 (N_14754,N_14458,N_14469);
or U14755 (N_14755,N_14096,N_14150);
xnor U14756 (N_14756,N_14270,N_14425);
nor U14757 (N_14757,N_14395,N_14055);
nand U14758 (N_14758,N_14108,N_14357);
and U14759 (N_14759,N_14035,N_14065);
and U14760 (N_14760,N_14130,N_14202);
or U14761 (N_14761,N_14081,N_14192);
xor U14762 (N_14762,N_14398,N_14066);
or U14763 (N_14763,N_14429,N_14063);
xor U14764 (N_14764,N_14213,N_14492);
and U14765 (N_14765,N_14355,N_14035);
or U14766 (N_14766,N_14034,N_14154);
and U14767 (N_14767,N_14483,N_14370);
nand U14768 (N_14768,N_14032,N_14035);
nand U14769 (N_14769,N_14462,N_14079);
nand U14770 (N_14770,N_14380,N_14080);
nand U14771 (N_14771,N_14416,N_14415);
nand U14772 (N_14772,N_14044,N_14279);
and U14773 (N_14773,N_14016,N_14375);
nor U14774 (N_14774,N_14011,N_14398);
nand U14775 (N_14775,N_14481,N_14437);
or U14776 (N_14776,N_14051,N_14463);
and U14777 (N_14777,N_14397,N_14179);
nand U14778 (N_14778,N_14161,N_14042);
nand U14779 (N_14779,N_14056,N_14018);
xor U14780 (N_14780,N_14215,N_14389);
nor U14781 (N_14781,N_14127,N_14430);
or U14782 (N_14782,N_14119,N_14427);
nand U14783 (N_14783,N_14375,N_14301);
nor U14784 (N_14784,N_14380,N_14442);
nand U14785 (N_14785,N_14304,N_14255);
and U14786 (N_14786,N_14016,N_14138);
nor U14787 (N_14787,N_14248,N_14122);
xor U14788 (N_14788,N_14249,N_14402);
xnor U14789 (N_14789,N_14422,N_14302);
nor U14790 (N_14790,N_14391,N_14403);
nor U14791 (N_14791,N_14411,N_14316);
xor U14792 (N_14792,N_14455,N_14425);
nand U14793 (N_14793,N_14331,N_14279);
nor U14794 (N_14794,N_14283,N_14293);
and U14795 (N_14795,N_14244,N_14307);
or U14796 (N_14796,N_14114,N_14074);
xnor U14797 (N_14797,N_14348,N_14128);
xor U14798 (N_14798,N_14184,N_14153);
nor U14799 (N_14799,N_14414,N_14007);
nand U14800 (N_14800,N_14288,N_14106);
xnor U14801 (N_14801,N_14082,N_14110);
or U14802 (N_14802,N_14351,N_14141);
or U14803 (N_14803,N_14222,N_14458);
xnor U14804 (N_14804,N_14249,N_14471);
and U14805 (N_14805,N_14033,N_14422);
nor U14806 (N_14806,N_14114,N_14004);
nor U14807 (N_14807,N_14430,N_14449);
xor U14808 (N_14808,N_14373,N_14065);
and U14809 (N_14809,N_14425,N_14414);
and U14810 (N_14810,N_14118,N_14111);
xnor U14811 (N_14811,N_14452,N_14226);
xor U14812 (N_14812,N_14059,N_14355);
nor U14813 (N_14813,N_14348,N_14365);
and U14814 (N_14814,N_14493,N_14492);
nand U14815 (N_14815,N_14262,N_14325);
xor U14816 (N_14816,N_14082,N_14080);
nor U14817 (N_14817,N_14054,N_14158);
or U14818 (N_14818,N_14487,N_14445);
or U14819 (N_14819,N_14415,N_14424);
nor U14820 (N_14820,N_14357,N_14467);
and U14821 (N_14821,N_14122,N_14280);
and U14822 (N_14822,N_14388,N_14033);
nand U14823 (N_14823,N_14084,N_14126);
or U14824 (N_14824,N_14255,N_14078);
nand U14825 (N_14825,N_14277,N_14014);
nor U14826 (N_14826,N_14483,N_14268);
and U14827 (N_14827,N_14295,N_14063);
and U14828 (N_14828,N_14225,N_14440);
nand U14829 (N_14829,N_14390,N_14092);
and U14830 (N_14830,N_14274,N_14300);
nor U14831 (N_14831,N_14118,N_14354);
nor U14832 (N_14832,N_14453,N_14393);
and U14833 (N_14833,N_14387,N_14097);
nor U14834 (N_14834,N_14386,N_14223);
and U14835 (N_14835,N_14455,N_14134);
and U14836 (N_14836,N_14165,N_14365);
and U14837 (N_14837,N_14073,N_14422);
or U14838 (N_14838,N_14353,N_14107);
nand U14839 (N_14839,N_14121,N_14496);
nand U14840 (N_14840,N_14100,N_14455);
nand U14841 (N_14841,N_14018,N_14376);
nor U14842 (N_14842,N_14283,N_14196);
xnor U14843 (N_14843,N_14265,N_14238);
or U14844 (N_14844,N_14410,N_14308);
nand U14845 (N_14845,N_14245,N_14134);
and U14846 (N_14846,N_14050,N_14137);
nand U14847 (N_14847,N_14356,N_14086);
or U14848 (N_14848,N_14330,N_14351);
or U14849 (N_14849,N_14164,N_14383);
and U14850 (N_14850,N_14441,N_14173);
and U14851 (N_14851,N_14099,N_14087);
nor U14852 (N_14852,N_14245,N_14159);
xnor U14853 (N_14853,N_14114,N_14035);
and U14854 (N_14854,N_14313,N_14157);
nor U14855 (N_14855,N_14407,N_14245);
xnor U14856 (N_14856,N_14276,N_14456);
nor U14857 (N_14857,N_14349,N_14339);
nand U14858 (N_14858,N_14487,N_14196);
nor U14859 (N_14859,N_14258,N_14171);
nor U14860 (N_14860,N_14046,N_14465);
nand U14861 (N_14861,N_14167,N_14059);
and U14862 (N_14862,N_14145,N_14459);
nor U14863 (N_14863,N_14406,N_14267);
or U14864 (N_14864,N_14354,N_14476);
and U14865 (N_14865,N_14279,N_14459);
nand U14866 (N_14866,N_14168,N_14440);
or U14867 (N_14867,N_14308,N_14359);
nor U14868 (N_14868,N_14364,N_14464);
nor U14869 (N_14869,N_14367,N_14182);
or U14870 (N_14870,N_14197,N_14056);
nand U14871 (N_14871,N_14060,N_14124);
and U14872 (N_14872,N_14404,N_14233);
and U14873 (N_14873,N_14371,N_14004);
nor U14874 (N_14874,N_14121,N_14092);
xnor U14875 (N_14875,N_14125,N_14492);
nor U14876 (N_14876,N_14433,N_14356);
nor U14877 (N_14877,N_14263,N_14364);
or U14878 (N_14878,N_14384,N_14281);
and U14879 (N_14879,N_14140,N_14235);
xor U14880 (N_14880,N_14437,N_14043);
or U14881 (N_14881,N_14332,N_14463);
or U14882 (N_14882,N_14400,N_14155);
xor U14883 (N_14883,N_14236,N_14416);
nor U14884 (N_14884,N_14450,N_14123);
xor U14885 (N_14885,N_14282,N_14310);
xnor U14886 (N_14886,N_14484,N_14001);
and U14887 (N_14887,N_14075,N_14013);
nand U14888 (N_14888,N_14471,N_14485);
nor U14889 (N_14889,N_14259,N_14463);
or U14890 (N_14890,N_14198,N_14335);
nand U14891 (N_14891,N_14315,N_14454);
xor U14892 (N_14892,N_14286,N_14444);
nand U14893 (N_14893,N_14290,N_14246);
nor U14894 (N_14894,N_14292,N_14127);
or U14895 (N_14895,N_14263,N_14123);
xnor U14896 (N_14896,N_14145,N_14301);
nand U14897 (N_14897,N_14100,N_14298);
nor U14898 (N_14898,N_14159,N_14489);
or U14899 (N_14899,N_14243,N_14235);
or U14900 (N_14900,N_14382,N_14267);
and U14901 (N_14901,N_14194,N_14071);
nand U14902 (N_14902,N_14326,N_14086);
or U14903 (N_14903,N_14072,N_14142);
nor U14904 (N_14904,N_14244,N_14287);
nand U14905 (N_14905,N_14291,N_14204);
xor U14906 (N_14906,N_14365,N_14120);
and U14907 (N_14907,N_14401,N_14209);
and U14908 (N_14908,N_14173,N_14256);
xor U14909 (N_14909,N_14296,N_14026);
nor U14910 (N_14910,N_14218,N_14478);
nor U14911 (N_14911,N_14324,N_14277);
xor U14912 (N_14912,N_14135,N_14081);
and U14913 (N_14913,N_14359,N_14090);
nor U14914 (N_14914,N_14166,N_14202);
and U14915 (N_14915,N_14488,N_14261);
and U14916 (N_14916,N_14382,N_14433);
xor U14917 (N_14917,N_14421,N_14001);
nand U14918 (N_14918,N_14115,N_14148);
nand U14919 (N_14919,N_14135,N_14365);
xnor U14920 (N_14920,N_14252,N_14009);
and U14921 (N_14921,N_14034,N_14499);
and U14922 (N_14922,N_14021,N_14179);
or U14923 (N_14923,N_14314,N_14464);
or U14924 (N_14924,N_14001,N_14383);
or U14925 (N_14925,N_14216,N_14389);
or U14926 (N_14926,N_14032,N_14467);
xor U14927 (N_14927,N_14359,N_14124);
or U14928 (N_14928,N_14301,N_14329);
nor U14929 (N_14929,N_14349,N_14106);
and U14930 (N_14930,N_14498,N_14003);
nor U14931 (N_14931,N_14243,N_14434);
nand U14932 (N_14932,N_14462,N_14415);
nand U14933 (N_14933,N_14130,N_14229);
or U14934 (N_14934,N_14092,N_14471);
nor U14935 (N_14935,N_14471,N_14040);
nand U14936 (N_14936,N_14106,N_14187);
nor U14937 (N_14937,N_14350,N_14019);
xnor U14938 (N_14938,N_14006,N_14193);
or U14939 (N_14939,N_14402,N_14112);
or U14940 (N_14940,N_14276,N_14352);
nand U14941 (N_14941,N_14409,N_14337);
or U14942 (N_14942,N_14464,N_14206);
and U14943 (N_14943,N_14340,N_14493);
or U14944 (N_14944,N_14399,N_14256);
nand U14945 (N_14945,N_14242,N_14220);
nor U14946 (N_14946,N_14268,N_14082);
nor U14947 (N_14947,N_14375,N_14025);
and U14948 (N_14948,N_14473,N_14040);
or U14949 (N_14949,N_14327,N_14407);
nor U14950 (N_14950,N_14457,N_14449);
nor U14951 (N_14951,N_14286,N_14021);
xnor U14952 (N_14952,N_14053,N_14481);
or U14953 (N_14953,N_14364,N_14146);
nor U14954 (N_14954,N_14456,N_14342);
and U14955 (N_14955,N_14274,N_14159);
nor U14956 (N_14956,N_14122,N_14062);
or U14957 (N_14957,N_14191,N_14460);
xnor U14958 (N_14958,N_14368,N_14028);
or U14959 (N_14959,N_14318,N_14440);
xnor U14960 (N_14960,N_14352,N_14157);
or U14961 (N_14961,N_14127,N_14097);
and U14962 (N_14962,N_14313,N_14190);
or U14963 (N_14963,N_14351,N_14457);
nand U14964 (N_14964,N_14460,N_14348);
xnor U14965 (N_14965,N_14254,N_14185);
nor U14966 (N_14966,N_14208,N_14473);
nand U14967 (N_14967,N_14150,N_14276);
nor U14968 (N_14968,N_14312,N_14117);
or U14969 (N_14969,N_14309,N_14459);
or U14970 (N_14970,N_14175,N_14454);
and U14971 (N_14971,N_14183,N_14335);
nand U14972 (N_14972,N_14456,N_14347);
and U14973 (N_14973,N_14132,N_14217);
and U14974 (N_14974,N_14487,N_14367);
nand U14975 (N_14975,N_14372,N_14001);
nor U14976 (N_14976,N_14188,N_14377);
and U14977 (N_14977,N_14220,N_14137);
nor U14978 (N_14978,N_14373,N_14317);
and U14979 (N_14979,N_14010,N_14401);
xnor U14980 (N_14980,N_14062,N_14326);
nand U14981 (N_14981,N_14326,N_14341);
nand U14982 (N_14982,N_14491,N_14451);
or U14983 (N_14983,N_14464,N_14016);
xnor U14984 (N_14984,N_14459,N_14303);
nand U14985 (N_14985,N_14398,N_14290);
and U14986 (N_14986,N_14356,N_14041);
or U14987 (N_14987,N_14308,N_14337);
or U14988 (N_14988,N_14094,N_14344);
xor U14989 (N_14989,N_14044,N_14375);
or U14990 (N_14990,N_14034,N_14317);
xnor U14991 (N_14991,N_14187,N_14049);
or U14992 (N_14992,N_14142,N_14290);
and U14993 (N_14993,N_14164,N_14084);
nor U14994 (N_14994,N_14294,N_14351);
or U14995 (N_14995,N_14326,N_14048);
nand U14996 (N_14996,N_14345,N_14370);
and U14997 (N_14997,N_14216,N_14083);
and U14998 (N_14998,N_14237,N_14276);
xor U14999 (N_14999,N_14117,N_14120);
xnor U15000 (N_15000,N_14781,N_14520);
and U15001 (N_15001,N_14915,N_14775);
nand U15002 (N_15002,N_14827,N_14691);
or U15003 (N_15003,N_14560,N_14729);
nor U15004 (N_15004,N_14661,N_14649);
xor U15005 (N_15005,N_14888,N_14767);
nor U15006 (N_15006,N_14702,N_14993);
nor U15007 (N_15007,N_14917,N_14923);
xor U15008 (N_15008,N_14864,N_14608);
and U15009 (N_15009,N_14554,N_14654);
and U15010 (N_15010,N_14591,N_14938);
or U15011 (N_15011,N_14823,N_14668);
xor U15012 (N_15012,N_14958,N_14934);
and U15013 (N_15013,N_14518,N_14943);
nand U15014 (N_15014,N_14969,N_14904);
and U15015 (N_15015,N_14564,N_14863);
or U15016 (N_15016,N_14881,N_14513);
and U15017 (N_15017,N_14652,N_14737);
or U15018 (N_15018,N_14879,N_14524);
nand U15019 (N_15019,N_14736,N_14964);
nand U15020 (N_15020,N_14629,N_14862);
and U15021 (N_15021,N_14821,N_14714);
and U15022 (N_15022,N_14562,N_14657);
or U15023 (N_15023,N_14713,N_14880);
nand U15024 (N_15024,N_14538,N_14916);
or U15025 (N_15025,N_14968,N_14859);
nand U15026 (N_15026,N_14996,N_14906);
or U15027 (N_15027,N_14532,N_14505);
nand U15028 (N_15028,N_14644,N_14635);
or U15029 (N_15029,N_14517,N_14632);
and U15030 (N_15030,N_14876,N_14975);
and U15031 (N_15031,N_14620,N_14832);
and U15032 (N_15032,N_14616,N_14986);
and U15033 (N_15033,N_14609,N_14959);
and U15034 (N_15034,N_14667,N_14642);
nor U15035 (N_15035,N_14614,N_14724);
or U15036 (N_15036,N_14739,N_14779);
xnor U15037 (N_15037,N_14857,N_14741);
xnor U15038 (N_15038,N_14646,N_14553);
xor U15039 (N_15039,N_14810,N_14860);
xor U15040 (N_15040,N_14761,N_14809);
and U15041 (N_15041,N_14953,N_14950);
xor U15042 (N_15042,N_14613,N_14659);
nor U15043 (N_15043,N_14547,N_14673);
nand U15044 (N_15044,N_14971,N_14634);
nand U15045 (N_15045,N_14542,N_14941);
and U15046 (N_15046,N_14872,N_14748);
nor U15047 (N_15047,N_14587,N_14569);
or U15048 (N_15048,N_14704,N_14588);
and U15049 (N_15049,N_14678,N_14636);
and U15050 (N_15050,N_14597,N_14840);
xnor U15051 (N_15051,N_14565,N_14617);
and U15052 (N_15052,N_14626,N_14793);
nor U15053 (N_15053,N_14638,N_14526);
nand U15054 (N_15054,N_14987,N_14798);
and U15055 (N_15055,N_14786,N_14817);
and U15056 (N_15056,N_14794,N_14692);
nor U15057 (N_15057,N_14769,N_14552);
xnor U15058 (N_15058,N_14948,N_14776);
xnor U15059 (N_15059,N_14967,N_14728);
nor U15060 (N_15060,N_14624,N_14603);
nor U15061 (N_15061,N_14960,N_14537);
nand U15062 (N_15062,N_14585,N_14628);
or U15063 (N_15063,N_14965,N_14666);
nand U15064 (N_15064,N_14839,N_14842);
nor U15065 (N_15065,N_14921,N_14605);
xor U15066 (N_15066,N_14725,N_14858);
nor U15067 (N_15067,N_14818,N_14508);
nand U15068 (N_15068,N_14995,N_14695);
or U15069 (N_15069,N_14892,N_14674);
nand U15070 (N_15070,N_14604,N_14662);
xor U15071 (N_15071,N_14716,N_14787);
or U15072 (N_15072,N_14530,N_14581);
and U15073 (N_15073,N_14961,N_14510);
and U15074 (N_15074,N_14730,N_14789);
or U15075 (N_15075,N_14825,N_14722);
xor U15076 (N_15076,N_14621,N_14648);
or U15077 (N_15077,N_14602,N_14875);
xor U15078 (N_15078,N_14877,N_14759);
and U15079 (N_15079,N_14852,N_14544);
xnor U15080 (N_15080,N_14801,N_14531);
nor U15081 (N_15081,N_14846,N_14751);
and U15082 (N_15082,N_14523,N_14966);
nor U15083 (N_15083,N_14803,N_14850);
xor U15084 (N_15084,N_14952,N_14516);
nand U15085 (N_15085,N_14791,N_14972);
nand U15086 (N_15086,N_14985,N_14782);
xnor U15087 (N_15087,N_14910,N_14549);
nor U15088 (N_15088,N_14559,N_14945);
or U15089 (N_15089,N_14844,N_14509);
xnor U15090 (N_15090,N_14732,N_14521);
and U15091 (N_15091,N_14738,N_14784);
and U15092 (N_15092,N_14999,N_14593);
nor U15093 (N_15093,N_14816,N_14762);
or U15094 (N_15094,N_14944,N_14541);
nand U15095 (N_15095,N_14785,N_14643);
nand U15096 (N_15096,N_14705,N_14687);
or U15097 (N_15097,N_14677,N_14914);
and U15098 (N_15098,N_14765,N_14719);
or U15099 (N_15099,N_14824,N_14992);
nor U15100 (N_15100,N_14778,N_14500);
nand U15101 (N_15101,N_14755,N_14685);
xnor U15102 (N_15102,N_14694,N_14957);
xor U15103 (N_15103,N_14693,N_14932);
xnor U15104 (N_15104,N_14973,N_14780);
nor U15105 (N_15105,N_14925,N_14893);
nor U15106 (N_15106,N_14865,N_14894);
xor U15107 (N_15107,N_14718,N_14856);
nor U15108 (N_15108,N_14774,N_14631);
xnor U15109 (N_15109,N_14672,N_14820);
xnor U15110 (N_15110,N_14637,N_14918);
and U15111 (N_15111,N_14535,N_14670);
nor U15112 (N_15112,N_14773,N_14903);
nor U15113 (N_15113,N_14507,N_14754);
or U15114 (N_15114,N_14777,N_14954);
xor U15115 (N_15115,N_14895,N_14701);
nor U15116 (N_15116,N_14655,N_14570);
xor U15117 (N_15117,N_14706,N_14586);
nor U15118 (N_15118,N_14897,N_14578);
xnor U15119 (N_15119,N_14989,N_14805);
nand U15120 (N_15120,N_14703,N_14909);
xnor U15121 (N_15121,N_14527,N_14561);
or U15122 (N_15122,N_14911,N_14633);
nor U15123 (N_15123,N_14502,N_14887);
and U15124 (N_15124,N_14851,N_14822);
and U15125 (N_15125,N_14800,N_14788);
xor U15126 (N_15126,N_14760,N_14815);
or U15127 (N_15127,N_14883,N_14749);
nand U15128 (N_15128,N_14556,N_14885);
and U15129 (N_15129,N_14772,N_14830);
nand U15130 (N_15130,N_14550,N_14981);
xor U15131 (N_15131,N_14905,N_14841);
or U15132 (N_15132,N_14506,N_14861);
and U15133 (N_15133,N_14874,N_14574);
nand U15134 (N_15134,N_14884,N_14924);
nor U15135 (N_15135,N_14976,N_14997);
and U15136 (N_15136,N_14849,N_14807);
and U15137 (N_15137,N_14831,N_14834);
xor U15138 (N_15138,N_14653,N_14675);
xnor U15139 (N_15139,N_14843,N_14828);
nor U15140 (N_15140,N_14869,N_14912);
nand U15141 (N_15141,N_14625,N_14600);
xnor U15142 (N_15142,N_14650,N_14567);
nor U15143 (N_15143,N_14770,N_14866);
nand U15144 (N_15144,N_14717,N_14684);
and U15145 (N_15145,N_14899,N_14937);
xnor U15146 (N_15146,N_14835,N_14814);
or U15147 (N_15147,N_14630,N_14745);
xor U15148 (N_15148,N_14512,N_14826);
xnor U15149 (N_15149,N_14598,N_14720);
or U15150 (N_15150,N_14991,N_14853);
nand U15151 (N_15151,N_14536,N_14726);
nand U15152 (N_15152,N_14868,N_14927);
nand U15153 (N_15153,N_14902,N_14599);
xnor U15154 (N_15154,N_14699,N_14886);
or U15155 (N_15155,N_14721,N_14922);
nand U15156 (N_15156,N_14504,N_14688);
and U15157 (N_15157,N_14572,N_14664);
xor U15158 (N_15158,N_14882,N_14896);
nand U15159 (N_15159,N_14682,N_14790);
nor U15160 (N_15160,N_14974,N_14514);
and U15161 (N_15161,N_14533,N_14583);
nor U15162 (N_15162,N_14764,N_14756);
nor U15163 (N_15163,N_14982,N_14689);
or U15164 (N_15164,N_14566,N_14946);
nand U15165 (N_15165,N_14811,N_14796);
nand U15166 (N_15166,N_14848,N_14949);
nor U15167 (N_15167,N_14658,N_14519);
nor U15168 (N_15168,N_14998,N_14898);
nand U15169 (N_15169,N_14891,N_14802);
nor U15170 (N_15170,N_14928,N_14819);
or U15171 (N_15171,N_14837,N_14931);
nand U15172 (N_15172,N_14576,N_14980);
xnor U15173 (N_15173,N_14766,N_14539);
nand U15174 (N_15174,N_14935,N_14596);
and U15175 (N_15175,N_14607,N_14690);
or U15176 (N_15176,N_14577,N_14540);
or U15177 (N_15177,N_14994,N_14669);
or U15178 (N_15178,N_14771,N_14686);
xnor U15179 (N_15179,N_14584,N_14829);
nand U15180 (N_15180,N_14988,N_14715);
or U15181 (N_15181,N_14511,N_14676);
and U15182 (N_15182,N_14697,N_14663);
xor U15183 (N_15183,N_14836,N_14733);
nand U15184 (N_15184,N_14696,N_14873);
nor U15185 (N_15185,N_14813,N_14501);
and U15186 (N_15186,N_14907,N_14568);
or U15187 (N_15187,N_14618,N_14855);
and U15188 (N_15188,N_14528,N_14610);
nor U15189 (N_15189,N_14947,N_14571);
and U15190 (N_15190,N_14752,N_14707);
or U15191 (N_15191,N_14792,N_14795);
nand U15192 (N_15192,N_14601,N_14930);
and U15193 (N_15193,N_14743,N_14742);
or U15194 (N_15194,N_14747,N_14783);
nand U15195 (N_15195,N_14639,N_14623);
nor U15196 (N_15196,N_14919,N_14845);
or U15197 (N_15197,N_14750,N_14606);
xor U15198 (N_15198,N_14970,N_14983);
nand U15199 (N_15199,N_14595,N_14627);
or U15200 (N_15200,N_14525,N_14589);
or U15201 (N_15201,N_14665,N_14529);
nor U15202 (N_15202,N_14956,N_14977);
or U15203 (N_15203,N_14647,N_14580);
nor U15204 (N_15204,N_14763,N_14575);
and U15205 (N_15205,N_14579,N_14723);
xnor U15206 (N_15206,N_14812,N_14515);
nand U15207 (N_15207,N_14592,N_14731);
xor U15208 (N_15208,N_14753,N_14735);
nor U15209 (N_15209,N_14838,N_14979);
xor U15210 (N_15210,N_14545,N_14942);
and U15211 (N_15211,N_14590,N_14870);
and U15212 (N_15212,N_14808,N_14867);
xor U15213 (N_15213,N_14619,N_14622);
nor U15214 (N_15214,N_14711,N_14727);
nor U15215 (N_15215,N_14854,N_14551);
or U15216 (N_15216,N_14656,N_14913);
and U15217 (N_15217,N_14920,N_14744);
nand U15218 (N_15218,N_14871,N_14546);
or U15219 (N_15219,N_14615,N_14757);
xnor U15220 (N_15220,N_14984,N_14963);
nor U15221 (N_15221,N_14878,N_14683);
and U15222 (N_15222,N_14962,N_14522);
nand U15223 (N_15223,N_14908,N_14712);
nand U15224 (N_15224,N_14594,N_14833);
and U15225 (N_15225,N_14804,N_14698);
or U15226 (N_15226,N_14955,N_14563);
or U15227 (N_15227,N_14951,N_14641);
and U15228 (N_15228,N_14543,N_14645);
xor U15229 (N_15229,N_14573,N_14890);
xor U15230 (N_15230,N_14582,N_14901);
xor U15231 (N_15231,N_14799,N_14660);
nor U15232 (N_15232,N_14768,N_14681);
nor U15233 (N_15233,N_14651,N_14940);
nor U15234 (N_15234,N_14555,N_14534);
or U15235 (N_15235,N_14700,N_14936);
xnor U15236 (N_15236,N_14709,N_14640);
nor U15237 (N_15237,N_14612,N_14900);
or U15238 (N_15238,N_14933,N_14680);
or U15239 (N_15239,N_14558,N_14990);
xor U15240 (N_15240,N_14926,N_14746);
nand U15241 (N_15241,N_14557,N_14797);
xor U15242 (N_15242,N_14889,N_14847);
or U15243 (N_15243,N_14758,N_14671);
nor U15244 (N_15244,N_14806,N_14740);
or U15245 (N_15245,N_14611,N_14503);
or U15246 (N_15246,N_14978,N_14679);
and U15247 (N_15247,N_14734,N_14548);
nor U15248 (N_15248,N_14708,N_14710);
nor U15249 (N_15249,N_14929,N_14939);
nand U15250 (N_15250,N_14550,N_14608);
and U15251 (N_15251,N_14555,N_14993);
xor U15252 (N_15252,N_14775,N_14723);
or U15253 (N_15253,N_14941,N_14652);
nor U15254 (N_15254,N_14795,N_14978);
and U15255 (N_15255,N_14554,N_14826);
nor U15256 (N_15256,N_14838,N_14650);
and U15257 (N_15257,N_14509,N_14997);
or U15258 (N_15258,N_14955,N_14523);
and U15259 (N_15259,N_14603,N_14664);
xor U15260 (N_15260,N_14541,N_14609);
or U15261 (N_15261,N_14769,N_14965);
and U15262 (N_15262,N_14541,N_14510);
or U15263 (N_15263,N_14885,N_14935);
or U15264 (N_15264,N_14669,N_14561);
nand U15265 (N_15265,N_14672,N_14720);
xnor U15266 (N_15266,N_14965,N_14991);
nand U15267 (N_15267,N_14731,N_14765);
nand U15268 (N_15268,N_14908,N_14806);
nor U15269 (N_15269,N_14642,N_14790);
nor U15270 (N_15270,N_14717,N_14705);
nand U15271 (N_15271,N_14911,N_14803);
or U15272 (N_15272,N_14991,N_14960);
nor U15273 (N_15273,N_14863,N_14709);
xor U15274 (N_15274,N_14732,N_14630);
or U15275 (N_15275,N_14875,N_14933);
nand U15276 (N_15276,N_14533,N_14962);
or U15277 (N_15277,N_14834,N_14610);
nand U15278 (N_15278,N_14503,N_14889);
or U15279 (N_15279,N_14617,N_14819);
or U15280 (N_15280,N_14562,N_14532);
and U15281 (N_15281,N_14704,N_14587);
and U15282 (N_15282,N_14868,N_14600);
xnor U15283 (N_15283,N_14797,N_14568);
nor U15284 (N_15284,N_14941,N_14705);
or U15285 (N_15285,N_14995,N_14711);
nor U15286 (N_15286,N_14883,N_14988);
nor U15287 (N_15287,N_14506,N_14661);
and U15288 (N_15288,N_14660,N_14997);
nor U15289 (N_15289,N_14712,N_14847);
xnor U15290 (N_15290,N_14543,N_14521);
and U15291 (N_15291,N_14541,N_14922);
xnor U15292 (N_15292,N_14900,N_14715);
or U15293 (N_15293,N_14891,N_14725);
and U15294 (N_15294,N_14501,N_14525);
nand U15295 (N_15295,N_14643,N_14852);
or U15296 (N_15296,N_14617,N_14584);
and U15297 (N_15297,N_14548,N_14820);
and U15298 (N_15298,N_14724,N_14569);
nand U15299 (N_15299,N_14883,N_14666);
nand U15300 (N_15300,N_14500,N_14710);
and U15301 (N_15301,N_14696,N_14677);
nand U15302 (N_15302,N_14747,N_14764);
nand U15303 (N_15303,N_14811,N_14923);
xnor U15304 (N_15304,N_14896,N_14506);
and U15305 (N_15305,N_14532,N_14958);
or U15306 (N_15306,N_14517,N_14933);
and U15307 (N_15307,N_14652,N_14636);
nor U15308 (N_15308,N_14691,N_14709);
nor U15309 (N_15309,N_14727,N_14995);
nand U15310 (N_15310,N_14949,N_14665);
nand U15311 (N_15311,N_14789,N_14808);
and U15312 (N_15312,N_14522,N_14820);
xnor U15313 (N_15313,N_14916,N_14541);
and U15314 (N_15314,N_14576,N_14835);
xnor U15315 (N_15315,N_14742,N_14754);
nand U15316 (N_15316,N_14696,N_14588);
nor U15317 (N_15317,N_14582,N_14921);
or U15318 (N_15318,N_14898,N_14666);
xor U15319 (N_15319,N_14955,N_14660);
xor U15320 (N_15320,N_14727,N_14856);
xor U15321 (N_15321,N_14563,N_14908);
and U15322 (N_15322,N_14502,N_14899);
nand U15323 (N_15323,N_14872,N_14854);
nand U15324 (N_15324,N_14772,N_14889);
xnor U15325 (N_15325,N_14863,N_14901);
or U15326 (N_15326,N_14695,N_14789);
and U15327 (N_15327,N_14969,N_14939);
or U15328 (N_15328,N_14822,N_14803);
and U15329 (N_15329,N_14935,N_14517);
and U15330 (N_15330,N_14570,N_14690);
nor U15331 (N_15331,N_14544,N_14792);
nand U15332 (N_15332,N_14713,N_14929);
xor U15333 (N_15333,N_14692,N_14906);
or U15334 (N_15334,N_14652,N_14841);
nor U15335 (N_15335,N_14845,N_14761);
and U15336 (N_15336,N_14688,N_14816);
nand U15337 (N_15337,N_14827,N_14607);
nor U15338 (N_15338,N_14763,N_14697);
nand U15339 (N_15339,N_14889,N_14654);
nor U15340 (N_15340,N_14917,N_14693);
and U15341 (N_15341,N_14604,N_14848);
and U15342 (N_15342,N_14656,N_14953);
nor U15343 (N_15343,N_14638,N_14819);
xnor U15344 (N_15344,N_14501,N_14506);
xnor U15345 (N_15345,N_14703,N_14983);
or U15346 (N_15346,N_14715,N_14998);
xor U15347 (N_15347,N_14934,N_14770);
nand U15348 (N_15348,N_14606,N_14664);
and U15349 (N_15349,N_14839,N_14682);
nor U15350 (N_15350,N_14934,N_14624);
nor U15351 (N_15351,N_14698,N_14846);
xnor U15352 (N_15352,N_14593,N_14889);
nand U15353 (N_15353,N_14711,N_14870);
nor U15354 (N_15354,N_14830,N_14788);
nor U15355 (N_15355,N_14621,N_14900);
nand U15356 (N_15356,N_14601,N_14631);
nand U15357 (N_15357,N_14757,N_14721);
and U15358 (N_15358,N_14592,N_14857);
and U15359 (N_15359,N_14633,N_14573);
nor U15360 (N_15360,N_14726,N_14830);
nand U15361 (N_15361,N_14505,N_14931);
and U15362 (N_15362,N_14784,N_14890);
or U15363 (N_15363,N_14884,N_14957);
xnor U15364 (N_15364,N_14644,N_14620);
xor U15365 (N_15365,N_14877,N_14920);
xnor U15366 (N_15366,N_14939,N_14591);
nor U15367 (N_15367,N_14960,N_14838);
xnor U15368 (N_15368,N_14503,N_14586);
nand U15369 (N_15369,N_14827,N_14829);
nand U15370 (N_15370,N_14666,N_14845);
or U15371 (N_15371,N_14774,N_14876);
nand U15372 (N_15372,N_14785,N_14793);
xor U15373 (N_15373,N_14794,N_14805);
and U15374 (N_15374,N_14862,N_14967);
nor U15375 (N_15375,N_14991,N_14813);
or U15376 (N_15376,N_14734,N_14880);
or U15377 (N_15377,N_14605,N_14854);
or U15378 (N_15378,N_14980,N_14626);
xor U15379 (N_15379,N_14621,N_14691);
and U15380 (N_15380,N_14552,N_14966);
nand U15381 (N_15381,N_14717,N_14844);
nand U15382 (N_15382,N_14535,N_14875);
xnor U15383 (N_15383,N_14552,N_14637);
or U15384 (N_15384,N_14589,N_14885);
xor U15385 (N_15385,N_14853,N_14510);
or U15386 (N_15386,N_14535,N_14509);
xor U15387 (N_15387,N_14970,N_14974);
xor U15388 (N_15388,N_14511,N_14744);
nor U15389 (N_15389,N_14596,N_14567);
and U15390 (N_15390,N_14794,N_14851);
nand U15391 (N_15391,N_14863,N_14612);
nand U15392 (N_15392,N_14925,N_14963);
nand U15393 (N_15393,N_14675,N_14925);
and U15394 (N_15394,N_14547,N_14761);
nor U15395 (N_15395,N_14522,N_14650);
and U15396 (N_15396,N_14590,N_14831);
xor U15397 (N_15397,N_14747,N_14689);
nor U15398 (N_15398,N_14686,N_14976);
and U15399 (N_15399,N_14689,N_14646);
nand U15400 (N_15400,N_14554,N_14969);
nor U15401 (N_15401,N_14508,N_14580);
and U15402 (N_15402,N_14856,N_14662);
nor U15403 (N_15403,N_14965,N_14959);
or U15404 (N_15404,N_14722,N_14691);
nand U15405 (N_15405,N_14559,N_14745);
or U15406 (N_15406,N_14867,N_14655);
or U15407 (N_15407,N_14831,N_14916);
and U15408 (N_15408,N_14724,N_14811);
nor U15409 (N_15409,N_14554,N_14559);
and U15410 (N_15410,N_14741,N_14558);
and U15411 (N_15411,N_14913,N_14774);
nor U15412 (N_15412,N_14738,N_14657);
or U15413 (N_15413,N_14821,N_14633);
or U15414 (N_15414,N_14603,N_14763);
nor U15415 (N_15415,N_14748,N_14565);
or U15416 (N_15416,N_14560,N_14770);
or U15417 (N_15417,N_14888,N_14737);
or U15418 (N_15418,N_14565,N_14782);
or U15419 (N_15419,N_14553,N_14771);
nor U15420 (N_15420,N_14702,N_14915);
nand U15421 (N_15421,N_14812,N_14934);
nor U15422 (N_15422,N_14525,N_14987);
and U15423 (N_15423,N_14644,N_14762);
nor U15424 (N_15424,N_14884,N_14863);
and U15425 (N_15425,N_14553,N_14558);
or U15426 (N_15426,N_14624,N_14579);
and U15427 (N_15427,N_14601,N_14958);
nor U15428 (N_15428,N_14501,N_14934);
and U15429 (N_15429,N_14917,N_14734);
and U15430 (N_15430,N_14888,N_14677);
and U15431 (N_15431,N_14779,N_14671);
xor U15432 (N_15432,N_14697,N_14861);
xnor U15433 (N_15433,N_14849,N_14508);
nor U15434 (N_15434,N_14717,N_14834);
xnor U15435 (N_15435,N_14691,N_14546);
or U15436 (N_15436,N_14606,N_14861);
or U15437 (N_15437,N_14848,N_14861);
and U15438 (N_15438,N_14672,N_14892);
or U15439 (N_15439,N_14671,N_14991);
or U15440 (N_15440,N_14621,N_14802);
nor U15441 (N_15441,N_14608,N_14553);
nand U15442 (N_15442,N_14602,N_14516);
xor U15443 (N_15443,N_14624,N_14538);
nand U15444 (N_15444,N_14951,N_14841);
or U15445 (N_15445,N_14781,N_14880);
nand U15446 (N_15446,N_14552,N_14554);
or U15447 (N_15447,N_14546,N_14745);
nor U15448 (N_15448,N_14914,N_14754);
nand U15449 (N_15449,N_14642,N_14823);
nand U15450 (N_15450,N_14936,N_14986);
xor U15451 (N_15451,N_14693,N_14620);
nand U15452 (N_15452,N_14938,N_14542);
and U15453 (N_15453,N_14680,N_14840);
xor U15454 (N_15454,N_14825,N_14609);
xnor U15455 (N_15455,N_14605,N_14975);
xnor U15456 (N_15456,N_14892,N_14887);
nor U15457 (N_15457,N_14774,N_14586);
or U15458 (N_15458,N_14651,N_14739);
nor U15459 (N_15459,N_14611,N_14606);
and U15460 (N_15460,N_14763,N_14988);
nand U15461 (N_15461,N_14906,N_14697);
xnor U15462 (N_15462,N_14838,N_14651);
nor U15463 (N_15463,N_14743,N_14860);
and U15464 (N_15464,N_14822,N_14663);
and U15465 (N_15465,N_14982,N_14935);
nand U15466 (N_15466,N_14716,N_14702);
xnor U15467 (N_15467,N_14777,N_14879);
or U15468 (N_15468,N_14525,N_14885);
and U15469 (N_15469,N_14544,N_14618);
nor U15470 (N_15470,N_14608,N_14520);
and U15471 (N_15471,N_14956,N_14650);
nor U15472 (N_15472,N_14778,N_14986);
or U15473 (N_15473,N_14509,N_14661);
and U15474 (N_15474,N_14602,N_14821);
nand U15475 (N_15475,N_14545,N_14909);
nor U15476 (N_15476,N_14997,N_14891);
nor U15477 (N_15477,N_14710,N_14835);
or U15478 (N_15478,N_14698,N_14713);
and U15479 (N_15479,N_14703,N_14614);
nor U15480 (N_15480,N_14578,N_14522);
xnor U15481 (N_15481,N_14797,N_14837);
xnor U15482 (N_15482,N_14728,N_14589);
or U15483 (N_15483,N_14837,N_14921);
and U15484 (N_15484,N_14550,N_14797);
nor U15485 (N_15485,N_14650,N_14700);
nor U15486 (N_15486,N_14972,N_14826);
or U15487 (N_15487,N_14858,N_14964);
and U15488 (N_15488,N_14943,N_14513);
and U15489 (N_15489,N_14608,N_14676);
and U15490 (N_15490,N_14973,N_14798);
nand U15491 (N_15491,N_14923,N_14655);
nor U15492 (N_15492,N_14759,N_14767);
and U15493 (N_15493,N_14704,N_14646);
xnor U15494 (N_15494,N_14667,N_14707);
and U15495 (N_15495,N_14667,N_14724);
or U15496 (N_15496,N_14574,N_14952);
nand U15497 (N_15497,N_14742,N_14780);
nor U15498 (N_15498,N_14745,N_14721);
nand U15499 (N_15499,N_14904,N_14766);
nand U15500 (N_15500,N_15190,N_15438);
nand U15501 (N_15501,N_15077,N_15089);
xor U15502 (N_15502,N_15234,N_15224);
or U15503 (N_15503,N_15161,N_15499);
or U15504 (N_15504,N_15176,N_15251);
and U15505 (N_15505,N_15377,N_15189);
xnor U15506 (N_15506,N_15146,N_15264);
nor U15507 (N_15507,N_15180,N_15462);
nor U15508 (N_15508,N_15047,N_15247);
xnor U15509 (N_15509,N_15380,N_15030);
nor U15510 (N_15510,N_15246,N_15254);
xnor U15511 (N_15511,N_15059,N_15043);
and U15512 (N_15512,N_15450,N_15464);
or U15513 (N_15513,N_15303,N_15442);
or U15514 (N_15514,N_15471,N_15472);
nand U15515 (N_15515,N_15400,N_15424);
xnor U15516 (N_15516,N_15166,N_15045);
nor U15517 (N_15517,N_15277,N_15355);
and U15518 (N_15518,N_15091,N_15087);
or U15519 (N_15519,N_15330,N_15009);
nand U15520 (N_15520,N_15186,N_15396);
and U15521 (N_15521,N_15323,N_15114);
nand U15522 (N_15522,N_15178,N_15308);
xnor U15523 (N_15523,N_15065,N_15299);
or U15524 (N_15524,N_15199,N_15405);
and U15525 (N_15525,N_15390,N_15134);
xor U15526 (N_15526,N_15426,N_15011);
or U15527 (N_15527,N_15031,N_15122);
xor U15528 (N_15528,N_15155,N_15286);
or U15529 (N_15529,N_15078,N_15226);
xor U15530 (N_15530,N_15468,N_15337);
nor U15531 (N_15531,N_15446,N_15113);
and U15532 (N_15532,N_15002,N_15076);
nand U15533 (N_15533,N_15205,N_15035);
nand U15534 (N_15534,N_15276,N_15084);
xnor U15535 (N_15535,N_15149,N_15202);
nand U15536 (N_15536,N_15128,N_15184);
nand U15537 (N_15537,N_15130,N_15174);
and U15538 (N_15538,N_15051,N_15253);
xor U15539 (N_15539,N_15217,N_15369);
xnor U15540 (N_15540,N_15452,N_15448);
and U15541 (N_15541,N_15340,N_15402);
and U15542 (N_15542,N_15016,N_15278);
or U15543 (N_15543,N_15231,N_15039);
and U15544 (N_15544,N_15328,N_15111);
nor U15545 (N_15545,N_15025,N_15046);
nor U15546 (N_15546,N_15107,N_15275);
and U15547 (N_15547,N_15159,N_15463);
nand U15548 (N_15548,N_15201,N_15342);
xnor U15549 (N_15549,N_15054,N_15353);
and U15550 (N_15550,N_15133,N_15191);
or U15551 (N_15551,N_15026,N_15170);
or U15552 (N_15552,N_15080,N_15418);
or U15553 (N_15553,N_15071,N_15129);
nand U15554 (N_15554,N_15187,N_15235);
or U15555 (N_15555,N_15348,N_15358);
nor U15556 (N_15556,N_15478,N_15289);
or U15557 (N_15557,N_15346,N_15257);
or U15558 (N_15558,N_15237,N_15371);
nand U15559 (N_15559,N_15086,N_15142);
xor U15560 (N_15560,N_15344,N_15301);
and U15561 (N_15561,N_15496,N_15072);
xnor U15562 (N_15562,N_15236,N_15392);
or U15563 (N_15563,N_15391,N_15458);
nand U15564 (N_15564,N_15415,N_15104);
nand U15565 (N_15565,N_15175,N_15284);
nand U15566 (N_15566,N_15304,N_15221);
or U15567 (N_15567,N_15449,N_15145);
xnor U15568 (N_15568,N_15085,N_15465);
or U15569 (N_15569,N_15197,N_15341);
or U15570 (N_15570,N_15292,N_15296);
nand U15571 (N_15571,N_15003,N_15117);
and U15572 (N_15572,N_15439,N_15131);
xnor U15573 (N_15573,N_15230,N_15469);
or U15574 (N_15574,N_15153,N_15193);
or U15575 (N_15575,N_15282,N_15399);
xnor U15576 (N_15576,N_15293,N_15165);
nand U15577 (N_15577,N_15056,N_15135);
xnor U15578 (N_15578,N_15171,N_15300);
and U15579 (N_15579,N_15315,N_15313);
and U15580 (N_15580,N_15032,N_15225);
xor U15581 (N_15581,N_15349,N_15382);
or U15582 (N_15582,N_15352,N_15356);
nand U15583 (N_15583,N_15447,N_15028);
or U15584 (N_15584,N_15453,N_15021);
nor U15585 (N_15585,N_15433,N_15474);
xnor U15586 (N_15586,N_15379,N_15115);
nor U15587 (N_15587,N_15416,N_15376);
nor U15588 (N_15588,N_15411,N_15419);
nor U15589 (N_15589,N_15069,N_15198);
nand U15590 (N_15590,N_15229,N_15258);
xor U15591 (N_15591,N_15177,N_15432);
or U15592 (N_15592,N_15015,N_15261);
xnor U15593 (N_15593,N_15157,N_15037);
or U15594 (N_15594,N_15470,N_15409);
and U15595 (N_15595,N_15154,N_15211);
or U15596 (N_15596,N_15126,N_15112);
nand U15597 (N_15597,N_15314,N_15033);
xnor U15598 (N_15598,N_15027,N_15057);
and U15599 (N_15599,N_15457,N_15403);
or U15600 (N_15600,N_15359,N_15298);
nand U15601 (N_15601,N_15218,N_15102);
or U15602 (N_15602,N_15367,N_15454);
nand U15603 (N_15603,N_15479,N_15081);
nand U15604 (N_15604,N_15417,N_15119);
and U15605 (N_15605,N_15412,N_15173);
and U15606 (N_15606,N_15188,N_15147);
nand U15607 (N_15607,N_15004,N_15013);
or U15608 (N_15608,N_15140,N_15326);
xor U15609 (N_15609,N_15196,N_15106);
or U15610 (N_15610,N_15260,N_15006);
and U15611 (N_15611,N_15481,N_15475);
and U15612 (N_15612,N_15339,N_15074);
xor U15613 (N_15613,N_15374,N_15351);
nor U15614 (N_15614,N_15386,N_15158);
xor U15615 (N_15615,N_15487,N_15216);
nand U15616 (N_15616,N_15305,N_15480);
nand U15617 (N_15617,N_15017,N_15441);
and U15618 (N_15618,N_15413,N_15431);
and U15619 (N_15619,N_15492,N_15148);
nor U15620 (N_15620,N_15241,N_15034);
and U15621 (N_15621,N_15014,N_15389);
xnor U15622 (N_15622,N_15443,N_15421);
xor U15623 (N_15623,N_15120,N_15408);
nor U15624 (N_15624,N_15336,N_15451);
xor U15625 (N_15625,N_15212,N_15317);
nand U15626 (N_15626,N_15223,N_15169);
nor U15627 (N_15627,N_15101,N_15363);
and U15628 (N_15628,N_15295,N_15040);
nand U15629 (N_15629,N_15401,N_15271);
nor U15630 (N_15630,N_15200,N_15082);
or U15631 (N_15631,N_15250,N_15309);
nand U15632 (N_15632,N_15052,N_15209);
nand U15633 (N_15633,N_15381,N_15100);
or U15634 (N_15634,N_15268,N_15321);
nand U15635 (N_15635,N_15375,N_15486);
nand U15636 (N_15636,N_15207,N_15497);
nor U15637 (N_15637,N_15372,N_15370);
xnor U15638 (N_15638,N_15123,N_15378);
xor U15639 (N_15639,N_15324,N_15310);
xor U15640 (N_15640,N_15092,N_15108);
or U15641 (N_15641,N_15345,N_15262);
nor U15642 (N_15642,N_15322,N_15210);
or U15643 (N_15643,N_15428,N_15194);
and U15644 (N_15644,N_15050,N_15498);
nand U15645 (N_15645,N_15285,N_15023);
nor U15646 (N_15646,N_15204,N_15150);
xnor U15647 (N_15647,N_15407,N_15182);
nand U15648 (N_15648,N_15110,N_15429);
nand U15649 (N_15649,N_15430,N_15063);
or U15650 (N_15650,N_15279,N_15167);
or U15651 (N_15651,N_15088,N_15215);
and U15652 (N_15652,N_15136,N_15090);
nor U15653 (N_15653,N_15272,N_15287);
or U15654 (N_15654,N_15311,N_15185);
nand U15655 (N_15655,N_15240,N_15493);
nand U15656 (N_15656,N_15312,N_15095);
xnor U15657 (N_15657,N_15327,N_15192);
xnor U15658 (N_15658,N_15066,N_15332);
nand U15659 (N_15659,N_15044,N_15083);
nand U15660 (N_15660,N_15476,N_15228);
nand U15661 (N_15661,N_15270,N_15297);
and U15662 (N_15662,N_15163,N_15488);
or U15663 (N_15663,N_15125,N_15001);
nor U15664 (N_15664,N_15164,N_15319);
and U15665 (N_15665,N_15259,N_15103);
and U15666 (N_15666,N_15096,N_15022);
nor U15667 (N_15667,N_15291,N_15109);
nor U15668 (N_15668,N_15427,N_15160);
xnor U15669 (N_15669,N_15099,N_15280);
and U15670 (N_15670,N_15141,N_15362);
nand U15671 (N_15671,N_15067,N_15219);
and U15672 (N_15672,N_15144,N_15124);
and U15673 (N_15673,N_15172,N_15121);
xor U15674 (N_15674,N_15306,N_15455);
xor U15675 (N_15675,N_15334,N_15220);
xnor U15676 (N_15676,N_15012,N_15393);
nand U15677 (N_15677,N_15325,N_15206);
and U15678 (N_15678,N_15238,N_15132);
xor U15679 (N_15679,N_15203,N_15385);
or U15680 (N_15680,N_15010,N_15440);
and U15681 (N_15681,N_15294,N_15435);
and U15682 (N_15682,N_15423,N_15459);
or U15683 (N_15683,N_15302,N_15307);
nand U15684 (N_15684,N_15288,N_15118);
and U15685 (N_15685,N_15064,N_15425);
and U15686 (N_15686,N_15460,N_15036);
and U15687 (N_15687,N_15456,N_15331);
and U15688 (N_15688,N_15473,N_15232);
and U15689 (N_15689,N_15137,N_15434);
or U15690 (N_15690,N_15490,N_15151);
nor U15691 (N_15691,N_15227,N_15061);
nor U15692 (N_15692,N_15213,N_15406);
nand U15693 (N_15693,N_15365,N_15055);
or U15694 (N_15694,N_15482,N_15138);
nor U15695 (N_15695,N_15179,N_15414);
nor U15696 (N_15696,N_15422,N_15263);
nand U15697 (N_15697,N_15152,N_15181);
and U15698 (N_15698,N_15373,N_15483);
and U15699 (N_15699,N_15444,N_15420);
xnor U15700 (N_15700,N_15366,N_15094);
nor U15701 (N_15701,N_15394,N_15368);
and U15702 (N_15702,N_15195,N_15244);
nand U15703 (N_15703,N_15222,N_15269);
nor U15704 (N_15704,N_15489,N_15343);
nand U15705 (N_15705,N_15384,N_15183);
or U15706 (N_15706,N_15333,N_15273);
xor U15707 (N_15707,N_15398,N_15461);
xor U15708 (N_15708,N_15255,N_15239);
nor U15709 (N_15709,N_15041,N_15274);
xnor U15710 (N_15710,N_15156,N_15397);
nand U15711 (N_15711,N_15008,N_15020);
nor U15712 (N_15712,N_15208,N_15053);
xnor U15713 (N_15713,N_15243,N_15005);
nor U15714 (N_15714,N_15338,N_15049);
nand U15715 (N_15715,N_15466,N_15316);
or U15716 (N_15716,N_15350,N_15073);
nand U15717 (N_15717,N_15256,N_15048);
and U15718 (N_15718,N_15242,N_15168);
or U15719 (N_15719,N_15248,N_15098);
xor U15720 (N_15720,N_15245,N_15029);
and U15721 (N_15721,N_15019,N_15105);
or U15722 (N_15722,N_15266,N_15068);
and U15723 (N_15723,N_15364,N_15070);
nor U15724 (N_15724,N_15007,N_15038);
nor U15725 (N_15725,N_15410,N_15062);
xor U15726 (N_15726,N_15281,N_15116);
or U15727 (N_15727,N_15097,N_15075);
and U15728 (N_15728,N_15143,N_15024);
nand U15729 (N_15729,N_15360,N_15437);
or U15730 (N_15730,N_15467,N_15162);
nand U15731 (N_15731,N_15495,N_15093);
nor U15732 (N_15732,N_15127,N_15357);
nand U15733 (N_15733,N_15491,N_15318);
or U15734 (N_15734,N_15042,N_15484);
or U15735 (N_15735,N_15436,N_15320);
nor U15736 (N_15736,N_15265,N_15139);
nor U15737 (N_15737,N_15477,N_15290);
or U15738 (N_15738,N_15335,N_15267);
xnor U15739 (N_15739,N_15347,N_15445);
nand U15740 (N_15740,N_15000,N_15214);
nand U15741 (N_15741,N_15494,N_15404);
nand U15742 (N_15742,N_15233,N_15387);
nor U15743 (N_15743,N_15485,N_15383);
and U15744 (N_15744,N_15249,N_15079);
xor U15745 (N_15745,N_15388,N_15354);
and U15746 (N_15746,N_15361,N_15060);
or U15747 (N_15747,N_15018,N_15252);
nor U15748 (N_15748,N_15329,N_15283);
nand U15749 (N_15749,N_15058,N_15395);
xor U15750 (N_15750,N_15200,N_15479);
and U15751 (N_15751,N_15338,N_15365);
or U15752 (N_15752,N_15196,N_15333);
nand U15753 (N_15753,N_15481,N_15494);
xor U15754 (N_15754,N_15268,N_15276);
and U15755 (N_15755,N_15462,N_15146);
and U15756 (N_15756,N_15229,N_15414);
and U15757 (N_15757,N_15239,N_15283);
or U15758 (N_15758,N_15087,N_15387);
and U15759 (N_15759,N_15322,N_15331);
nor U15760 (N_15760,N_15100,N_15234);
nand U15761 (N_15761,N_15191,N_15431);
xor U15762 (N_15762,N_15066,N_15427);
nand U15763 (N_15763,N_15492,N_15386);
nand U15764 (N_15764,N_15022,N_15217);
nor U15765 (N_15765,N_15015,N_15339);
and U15766 (N_15766,N_15388,N_15475);
or U15767 (N_15767,N_15124,N_15482);
or U15768 (N_15768,N_15361,N_15058);
and U15769 (N_15769,N_15173,N_15458);
xnor U15770 (N_15770,N_15071,N_15332);
or U15771 (N_15771,N_15084,N_15078);
nand U15772 (N_15772,N_15453,N_15304);
xor U15773 (N_15773,N_15152,N_15429);
nor U15774 (N_15774,N_15068,N_15483);
and U15775 (N_15775,N_15046,N_15192);
and U15776 (N_15776,N_15314,N_15389);
nand U15777 (N_15777,N_15144,N_15026);
and U15778 (N_15778,N_15297,N_15211);
nor U15779 (N_15779,N_15040,N_15245);
or U15780 (N_15780,N_15155,N_15369);
nand U15781 (N_15781,N_15111,N_15317);
and U15782 (N_15782,N_15450,N_15468);
or U15783 (N_15783,N_15133,N_15302);
and U15784 (N_15784,N_15115,N_15327);
xnor U15785 (N_15785,N_15447,N_15106);
and U15786 (N_15786,N_15487,N_15049);
or U15787 (N_15787,N_15317,N_15149);
xor U15788 (N_15788,N_15445,N_15066);
xnor U15789 (N_15789,N_15351,N_15104);
and U15790 (N_15790,N_15268,N_15493);
nor U15791 (N_15791,N_15351,N_15455);
xnor U15792 (N_15792,N_15211,N_15345);
and U15793 (N_15793,N_15282,N_15244);
and U15794 (N_15794,N_15332,N_15230);
nor U15795 (N_15795,N_15453,N_15005);
xor U15796 (N_15796,N_15113,N_15123);
nor U15797 (N_15797,N_15407,N_15475);
or U15798 (N_15798,N_15066,N_15226);
and U15799 (N_15799,N_15294,N_15317);
xnor U15800 (N_15800,N_15097,N_15463);
nor U15801 (N_15801,N_15378,N_15067);
xnor U15802 (N_15802,N_15444,N_15264);
nand U15803 (N_15803,N_15034,N_15289);
and U15804 (N_15804,N_15200,N_15277);
nor U15805 (N_15805,N_15491,N_15179);
and U15806 (N_15806,N_15342,N_15336);
or U15807 (N_15807,N_15397,N_15394);
nor U15808 (N_15808,N_15453,N_15287);
and U15809 (N_15809,N_15026,N_15194);
and U15810 (N_15810,N_15079,N_15386);
or U15811 (N_15811,N_15156,N_15197);
or U15812 (N_15812,N_15211,N_15145);
nand U15813 (N_15813,N_15037,N_15161);
and U15814 (N_15814,N_15337,N_15132);
xor U15815 (N_15815,N_15137,N_15287);
nand U15816 (N_15816,N_15219,N_15129);
and U15817 (N_15817,N_15345,N_15401);
and U15818 (N_15818,N_15057,N_15420);
or U15819 (N_15819,N_15298,N_15029);
or U15820 (N_15820,N_15230,N_15006);
or U15821 (N_15821,N_15429,N_15136);
nand U15822 (N_15822,N_15410,N_15334);
xor U15823 (N_15823,N_15363,N_15015);
xor U15824 (N_15824,N_15252,N_15152);
xnor U15825 (N_15825,N_15441,N_15257);
and U15826 (N_15826,N_15438,N_15033);
nand U15827 (N_15827,N_15395,N_15150);
nand U15828 (N_15828,N_15144,N_15482);
nand U15829 (N_15829,N_15146,N_15253);
nor U15830 (N_15830,N_15272,N_15249);
and U15831 (N_15831,N_15071,N_15205);
or U15832 (N_15832,N_15162,N_15088);
nand U15833 (N_15833,N_15176,N_15364);
and U15834 (N_15834,N_15179,N_15412);
xnor U15835 (N_15835,N_15345,N_15326);
xnor U15836 (N_15836,N_15190,N_15197);
and U15837 (N_15837,N_15183,N_15276);
nor U15838 (N_15838,N_15225,N_15399);
nor U15839 (N_15839,N_15219,N_15405);
xor U15840 (N_15840,N_15443,N_15066);
nand U15841 (N_15841,N_15438,N_15195);
xnor U15842 (N_15842,N_15243,N_15057);
nand U15843 (N_15843,N_15384,N_15015);
nor U15844 (N_15844,N_15160,N_15340);
or U15845 (N_15845,N_15008,N_15079);
nor U15846 (N_15846,N_15376,N_15469);
nor U15847 (N_15847,N_15134,N_15495);
nand U15848 (N_15848,N_15329,N_15066);
nor U15849 (N_15849,N_15407,N_15379);
and U15850 (N_15850,N_15348,N_15078);
and U15851 (N_15851,N_15150,N_15041);
xnor U15852 (N_15852,N_15085,N_15370);
xor U15853 (N_15853,N_15252,N_15176);
or U15854 (N_15854,N_15464,N_15091);
xor U15855 (N_15855,N_15478,N_15496);
and U15856 (N_15856,N_15298,N_15135);
or U15857 (N_15857,N_15103,N_15372);
nor U15858 (N_15858,N_15263,N_15121);
nand U15859 (N_15859,N_15376,N_15194);
and U15860 (N_15860,N_15485,N_15155);
or U15861 (N_15861,N_15072,N_15497);
xnor U15862 (N_15862,N_15248,N_15244);
and U15863 (N_15863,N_15274,N_15426);
nand U15864 (N_15864,N_15086,N_15012);
or U15865 (N_15865,N_15173,N_15292);
and U15866 (N_15866,N_15486,N_15073);
nor U15867 (N_15867,N_15379,N_15381);
nand U15868 (N_15868,N_15206,N_15005);
and U15869 (N_15869,N_15343,N_15342);
and U15870 (N_15870,N_15002,N_15239);
nor U15871 (N_15871,N_15442,N_15415);
or U15872 (N_15872,N_15351,N_15353);
xnor U15873 (N_15873,N_15228,N_15173);
nor U15874 (N_15874,N_15206,N_15026);
and U15875 (N_15875,N_15000,N_15375);
nor U15876 (N_15876,N_15244,N_15102);
nor U15877 (N_15877,N_15003,N_15255);
or U15878 (N_15878,N_15330,N_15070);
xor U15879 (N_15879,N_15228,N_15482);
and U15880 (N_15880,N_15059,N_15091);
and U15881 (N_15881,N_15478,N_15308);
nand U15882 (N_15882,N_15175,N_15338);
nand U15883 (N_15883,N_15355,N_15214);
nand U15884 (N_15884,N_15033,N_15196);
nand U15885 (N_15885,N_15388,N_15409);
or U15886 (N_15886,N_15193,N_15283);
nand U15887 (N_15887,N_15193,N_15391);
nor U15888 (N_15888,N_15155,N_15184);
and U15889 (N_15889,N_15376,N_15280);
nand U15890 (N_15890,N_15153,N_15175);
and U15891 (N_15891,N_15194,N_15390);
xor U15892 (N_15892,N_15188,N_15016);
nor U15893 (N_15893,N_15325,N_15472);
xnor U15894 (N_15894,N_15280,N_15423);
nor U15895 (N_15895,N_15072,N_15152);
nand U15896 (N_15896,N_15345,N_15410);
nand U15897 (N_15897,N_15343,N_15425);
and U15898 (N_15898,N_15285,N_15137);
xnor U15899 (N_15899,N_15096,N_15023);
and U15900 (N_15900,N_15129,N_15200);
nand U15901 (N_15901,N_15384,N_15302);
nor U15902 (N_15902,N_15236,N_15267);
and U15903 (N_15903,N_15201,N_15376);
or U15904 (N_15904,N_15314,N_15448);
and U15905 (N_15905,N_15151,N_15011);
or U15906 (N_15906,N_15228,N_15126);
nor U15907 (N_15907,N_15155,N_15041);
and U15908 (N_15908,N_15375,N_15407);
nand U15909 (N_15909,N_15003,N_15412);
or U15910 (N_15910,N_15493,N_15450);
nor U15911 (N_15911,N_15227,N_15195);
nor U15912 (N_15912,N_15290,N_15141);
nor U15913 (N_15913,N_15205,N_15037);
or U15914 (N_15914,N_15267,N_15132);
nand U15915 (N_15915,N_15094,N_15003);
nor U15916 (N_15916,N_15113,N_15427);
nand U15917 (N_15917,N_15181,N_15432);
xor U15918 (N_15918,N_15143,N_15470);
and U15919 (N_15919,N_15168,N_15424);
and U15920 (N_15920,N_15464,N_15361);
nand U15921 (N_15921,N_15255,N_15109);
nand U15922 (N_15922,N_15213,N_15447);
nor U15923 (N_15923,N_15371,N_15315);
nand U15924 (N_15924,N_15182,N_15158);
xor U15925 (N_15925,N_15007,N_15175);
or U15926 (N_15926,N_15021,N_15197);
nand U15927 (N_15927,N_15384,N_15258);
or U15928 (N_15928,N_15321,N_15247);
nand U15929 (N_15929,N_15048,N_15274);
and U15930 (N_15930,N_15063,N_15171);
nor U15931 (N_15931,N_15258,N_15048);
nor U15932 (N_15932,N_15353,N_15309);
nor U15933 (N_15933,N_15112,N_15006);
xnor U15934 (N_15934,N_15042,N_15057);
or U15935 (N_15935,N_15202,N_15053);
nor U15936 (N_15936,N_15091,N_15446);
and U15937 (N_15937,N_15030,N_15142);
nor U15938 (N_15938,N_15373,N_15242);
and U15939 (N_15939,N_15434,N_15145);
nand U15940 (N_15940,N_15177,N_15197);
and U15941 (N_15941,N_15215,N_15059);
nand U15942 (N_15942,N_15225,N_15181);
or U15943 (N_15943,N_15493,N_15030);
or U15944 (N_15944,N_15187,N_15473);
xnor U15945 (N_15945,N_15249,N_15299);
nand U15946 (N_15946,N_15351,N_15103);
nand U15947 (N_15947,N_15411,N_15041);
and U15948 (N_15948,N_15209,N_15468);
or U15949 (N_15949,N_15127,N_15470);
nand U15950 (N_15950,N_15303,N_15076);
xnor U15951 (N_15951,N_15300,N_15080);
nor U15952 (N_15952,N_15006,N_15313);
or U15953 (N_15953,N_15185,N_15313);
nor U15954 (N_15954,N_15110,N_15210);
and U15955 (N_15955,N_15318,N_15019);
or U15956 (N_15956,N_15232,N_15239);
or U15957 (N_15957,N_15084,N_15289);
nor U15958 (N_15958,N_15344,N_15455);
and U15959 (N_15959,N_15117,N_15332);
nor U15960 (N_15960,N_15273,N_15174);
or U15961 (N_15961,N_15146,N_15003);
or U15962 (N_15962,N_15443,N_15135);
xnor U15963 (N_15963,N_15104,N_15119);
and U15964 (N_15964,N_15160,N_15376);
xnor U15965 (N_15965,N_15033,N_15036);
nor U15966 (N_15966,N_15146,N_15080);
xnor U15967 (N_15967,N_15285,N_15205);
and U15968 (N_15968,N_15357,N_15364);
nor U15969 (N_15969,N_15082,N_15048);
nand U15970 (N_15970,N_15067,N_15472);
xor U15971 (N_15971,N_15274,N_15208);
or U15972 (N_15972,N_15352,N_15082);
nand U15973 (N_15973,N_15248,N_15045);
and U15974 (N_15974,N_15081,N_15480);
xnor U15975 (N_15975,N_15323,N_15087);
or U15976 (N_15976,N_15220,N_15389);
nand U15977 (N_15977,N_15496,N_15139);
or U15978 (N_15978,N_15461,N_15005);
nor U15979 (N_15979,N_15009,N_15434);
nand U15980 (N_15980,N_15484,N_15105);
nand U15981 (N_15981,N_15396,N_15187);
nand U15982 (N_15982,N_15187,N_15414);
nand U15983 (N_15983,N_15493,N_15235);
nand U15984 (N_15984,N_15408,N_15135);
nand U15985 (N_15985,N_15416,N_15142);
or U15986 (N_15986,N_15156,N_15324);
or U15987 (N_15987,N_15392,N_15172);
or U15988 (N_15988,N_15410,N_15395);
xor U15989 (N_15989,N_15184,N_15347);
nor U15990 (N_15990,N_15210,N_15089);
nor U15991 (N_15991,N_15104,N_15196);
and U15992 (N_15992,N_15335,N_15493);
and U15993 (N_15993,N_15039,N_15438);
nor U15994 (N_15994,N_15286,N_15147);
and U15995 (N_15995,N_15194,N_15475);
and U15996 (N_15996,N_15268,N_15416);
or U15997 (N_15997,N_15363,N_15197);
nor U15998 (N_15998,N_15235,N_15157);
and U15999 (N_15999,N_15392,N_15441);
nor U16000 (N_16000,N_15979,N_15702);
nand U16001 (N_16001,N_15845,N_15866);
xor U16002 (N_16002,N_15950,N_15563);
or U16003 (N_16003,N_15697,N_15712);
or U16004 (N_16004,N_15896,N_15568);
nor U16005 (N_16005,N_15564,N_15974);
or U16006 (N_16006,N_15973,N_15927);
nor U16007 (N_16007,N_15801,N_15941);
nor U16008 (N_16008,N_15537,N_15769);
or U16009 (N_16009,N_15682,N_15604);
nand U16010 (N_16010,N_15643,N_15555);
or U16011 (N_16011,N_15890,N_15882);
nor U16012 (N_16012,N_15990,N_15899);
nor U16013 (N_16013,N_15730,N_15918);
or U16014 (N_16014,N_15736,N_15581);
and U16015 (N_16015,N_15930,N_15764);
nand U16016 (N_16016,N_15820,N_15806);
or U16017 (N_16017,N_15638,N_15887);
nor U16018 (N_16018,N_15759,N_15575);
xor U16019 (N_16019,N_15931,N_15800);
xnor U16020 (N_16020,N_15876,N_15893);
nand U16021 (N_16021,N_15636,N_15963);
and U16022 (N_16022,N_15955,N_15543);
nand U16023 (N_16023,N_15623,N_15840);
nand U16024 (N_16024,N_15592,N_15583);
and U16025 (N_16025,N_15945,N_15711);
and U16026 (N_16026,N_15891,N_15559);
xnor U16027 (N_16027,N_15874,N_15617);
nor U16028 (N_16028,N_15809,N_15722);
and U16029 (N_16029,N_15902,N_15889);
xnor U16030 (N_16030,N_15777,N_15539);
xor U16031 (N_16031,N_15818,N_15762);
or U16032 (N_16032,N_15724,N_15506);
and U16033 (N_16033,N_15938,N_15821);
xor U16034 (N_16034,N_15673,N_15726);
and U16035 (N_16035,N_15576,N_15970);
or U16036 (N_16036,N_15886,N_15956);
and U16037 (N_16037,N_15854,N_15629);
or U16038 (N_16038,N_15785,N_15980);
xnor U16039 (N_16039,N_15901,N_15842);
xnor U16040 (N_16040,N_15758,N_15699);
nand U16041 (N_16041,N_15837,N_15528);
nand U16042 (N_16042,N_15529,N_15879);
nor U16043 (N_16043,N_15547,N_15860);
or U16044 (N_16044,N_15598,N_15792);
nand U16045 (N_16045,N_15844,N_15793);
nand U16046 (N_16046,N_15656,N_15784);
xnor U16047 (N_16047,N_15994,N_15753);
xor U16048 (N_16048,N_15632,N_15709);
nor U16049 (N_16049,N_15939,N_15805);
nor U16050 (N_16050,N_15765,N_15767);
nand U16051 (N_16051,N_15520,N_15650);
and U16052 (N_16052,N_15992,N_15962);
and U16053 (N_16053,N_15834,N_15881);
xor U16054 (N_16054,N_15525,N_15967);
or U16055 (N_16055,N_15982,N_15752);
xnor U16056 (N_16056,N_15734,N_15846);
nor U16057 (N_16057,N_15501,N_15557);
nor U16058 (N_16058,N_15908,N_15947);
or U16059 (N_16059,N_15684,N_15851);
and U16060 (N_16060,N_15880,N_15906);
or U16061 (N_16061,N_15668,N_15605);
or U16062 (N_16062,N_15634,N_15517);
nand U16063 (N_16063,N_15695,N_15553);
xor U16064 (N_16064,N_15716,N_15934);
xor U16065 (N_16065,N_15863,N_15612);
or U16066 (N_16066,N_15704,N_15572);
nand U16067 (N_16067,N_15571,N_15781);
nand U16068 (N_16068,N_15959,N_15871);
nor U16069 (N_16069,N_15855,N_15952);
and U16070 (N_16070,N_15674,N_15802);
or U16071 (N_16071,N_15878,N_15903);
and U16072 (N_16072,N_15868,N_15507);
nor U16073 (N_16073,N_15649,N_15922);
or U16074 (N_16074,N_15685,N_15535);
or U16075 (N_16075,N_15524,N_15664);
xor U16076 (N_16076,N_15676,N_15989);
xnor U16077 (N_16077,N_15620,N_15745);
nor U16078 (N_16078,N_15940,N_15628);
and U16079 (N_16079,N_15833,N_15751);
and U16080 (N_16080,N_15900,N_15771);
xor U16081 (N_16081,N_15857,N_15663);
and U16082 (N_16082,N_15971,N_15949);
nor U16083 (N_16083,N_15723,N_15627);
nand U16084 (N_16084,N_15741,N_15786);
nor U16085 (N_16085,N_15558,N_15953);
nand U16086 (N_16086,N_15826,N_15912);
nand U16087 (N_16087,N_15678,N_15590);
nand U16088 (N_16088,N_15740,N_15746);
nand U16089 (N_16089,N_15782,N_15582);
nand U16090 (N_16090,N_15509,N_15819);
nand U16091 (N_16091,N_15630,N_15679);
xnor U16092 (N_16092,N_15835,N_15502);
xnor U16093 (N_16093,N_15748,N_15708);
xor U16094 (N_16094,N_15850,N_15925);
nand U16095 (N_16095,N_15579,N_15607);
xnor U16096 (N_16096,N_15895,N_15768);
nand U16097 (N_16097,N_15964,N_15983);
or U16098 (N_16098,N_15984,N_15968);
xor U16099 (N_16099,N_15856,N_15905);
nor U16100 (N_16100,N_15957,N_15538);
and U16101 (N_16101,N_15926,N_15648);
xnor U16102 (N_16102,N_15587,N_15616);
nand U16103 (N_16103,N_15586,N_15591);
and U16104 (N_16104,N_15534,N_15776);
xor U16105 (N_16105,N_15613,N_15614);
xor U16106 (N_16106,N_15681,N_15827);
and U16107 (N_16107,N_15817,N_15594);
nor U16108 (N_16108,N_15694,N_15904);
or U16109 (N_16109,N_15545,N_15810);
xnor U16110 (N_16110,N_15830,N_15611);
and U16111 (N_16111,N_15670,N_15864);
xnor U16112 (N_16112,N_15935,N_15892);
or U16113 (N_16113,N_15633,N_15812);
nor U16114 (N_16114,N_15943,N_15798);
and U16115 (N_16115,N_15873,N_15606);
nand U16116 (N_16116,N_15503,N_15774);
xor U16117 (N_16117,N_15839,N_15631);
or U16118 (N_16118,N_15909,N_15573);
or U16119 (N_16119,N_15719,N_15862);
or U16120 (N_16120,N_15500,N_15677);
nor U16121 (N_16121,N_15518,N_15701);
and U16122 (N_16122,N_15640,N_15703);
and U16123 (N_16123,N_15595,N_15825);
and U16124 (N_16124,N_15698,N_15732);
xnor U16125 (N_16125,N_15706,N_15933);
nand U16126 (N_16126,N_15823,N_15907);
or U16127 (N_16127,N_15683,N_15513);
or U16128 (N_16128,N_15660,N_15512);
nand U16129 (N_16129,N_15742,N_15618);
xor U16130 (N_16130,N_15843,N_15960);
or U16131 (N_16131,N_15756,N_15584);
nand U16132 (N_16132,N_15877,N_15526);
nor U16133 (N_16133,N_15665,N_15853);
xor U16134 (N_16134,N_15675,N_15519);
nor U16135 (N_16135,N_15965,N_15936);
nand U16136 (N_16136,N_15621,N_15847);
xor U16137 (N_16137,N_15779,N_15996);
xnor U16138 (N_16138,N_15937,N_15511);
xor U16139 (N_16139,N_15822,N_15692);
xor U16140 (N_16140,N_15888,N_15666);
nor U16141 (N_16141,N_15549,N_15527);
and U16142 (N_16142,N_15915,N_15811);
and U16143 (N_16143,N_15735,N_15977);
xor U16144 (N_16144,N_15754,N_15689);
and U16145 (N_16145,N_15574,N_15929);
nor U16146 (N_16146,N_15521,N_15978);
xnor U16147 (N_16147,N_15848,N_15763);
xor U16148 (N_16148,N_15790,N_15505);
xnor U16149 (N_16149,N_15911,N_15794);
or U16150 (N_16150,N_15787,N_15551);
xor U16151 (N_16151,N_15804,N_15687);
xnor U16152 (N_16152,N_15803,N_15609);
xnor U16153 (N_16153,N_15789,N_15791);
nor U16154 (N_16154,N_15816,N_15870);
nand U16155 (N_16155,N_15797,N_15757);
and U16156 (N_16156,N_15731,N_15775);
or U16157 (N_16157,N_15898,N_15642);
nand U16158 (N_16158,N_15924,N_15836);
xnor U16159 (N_16159,N_15690,N_15639);
xor U16160 (N_16160,N_15829,N_15920);
and U16161 (N_16161,N_15700,N_15867);
xnor U16162 (N_16162,N_15608,N_15921);
and U16163 (N_16163,N_15885,N_15986);
and U16164 (N_16164,N_15662,N_15913);
and U16165 (N_16165,N_15747,N_15593);
nor U16166 (N_16166,N_15966,N_15696);
nand U16167 (N_16167,N_15749,N_15991);
or U16168 (N_16168,N_15667,N_15714);
and U16169 (N_16169,N_15766,N_15672);
nor U16170 (N_16170,N_15654,N_15588);
or U16171 (N_16171,N_15733,N_15715);
nor U16172 (N_16172,N_15619,N_15807);
xor U16173 (N_16173,N_15824,N_15993);
xnor U16174 (N_16174,N_15884,N_15958);
xnor U16175 (N_16175,N_15651,N_15669);
and U16176 (N_16176,N_15596,N_15849);
nor U16177 (N_16177,N_15705,N_15969);
nor U16178 (N_16178,N_15727,N_15540);
xor U16179 (N_16179,N_15644,N_15721);
or U16180 (N_16180,N_15624,N_15508);
and U16181 (N_16181,N_15577,N_15815);
and U16182 (N_16182,N_15671,N_15772);
nand U16183 (N_16183,N_15795,N_15999);
xor U16184 (N_16184,N_15661,N_15869);
xor U16185 (N_16185,N_15658,N_15522);
nand U16186 (N_16186,N_15897,N_15917);
nand U16187 (N_16187,N_15602,N_15626);
nor U16188 (N_16188,N_15972,N_15928);
nor U16189 (N_16189,N_15883,N_15760);
nor U16190 (N_16190,N_15635,N_15585);
nand U16191 (N_16191,N_15916,N_15813);
nand U16192 (N_16192,N_15961,N_15561);
xor U16193 (N_16193,N_15570,N_15985);
nand U16194 (N_16194,N_15707,N_15975);
nor U16195 (N_16195,N_15770,N_15637);
and U16196 (N_16196,N_15910,N_15875);
or U16197 (N_16197,N_15566,N_15743);
and U16198 (N_16198,N_15828,N_15814);
nor U16199 (N_16199,N_15569,N_15976);
nor U16200 (N_16200,N_15546,N_15542);
and U16201 (N_16201,N_15646,N_15544);
nand U16202 (N_16202,N_15783,N_15514);
or U16203 (N_16203,N_15995,N_15615);
xnor U16204 (N_16204,N_15680,N_15567);
nand U16205 (N_16205,N_15718,N_15531);
or U16206 (N_16206,N_15686,N_15773);
and U16207 (N_16207,N_15720,N_15923);
or U16208 (N_16208,N_15641,N_15516);
and U16209 (N_16209,N_15778,N_15796);
nor U16210 (N_16210,N_15652,N_15536);
or U16211 (N_16211,N_15647,N_15914);
or U16212 (N_16212,N_15831,N_15523);
and U16213 (N_16213,N_15548,N_15859);
and U16214 (N_16214,N_15562,N_15659);
nor U16215 (N_16215,N_15894,N_15738);
xor U16216 (N_16216,N_15541,N_15530);
or U16217 (N_16217,N_15865,N_15515);
xor U16218 (N_16218,N_15988,N_15578);
nor U16219 (N_16219,N_15554,N_15932);
or U16220 (N_16220,N_15841,N_15597);
and U16221 (N_16221,N_15954,N_15981);
or U16222 (N_16222,N_15655,N_15852);
and U16223 (N_16223,N_15589,N_15750);
or U16224 (N_16224,N_15838,N_15737);
nor U16225 (N_16225,N_15951,N_15691);
and U16226 (N_16226,N_15601,N_15550);
and U16227 (N_16227,N_15808,N_15560);
xor U16228 (N_16228,N_15713,N_15603);
xor U16229 (N_16229,N_15556,N_15645);
and U16230 (N_16230,N_15739,N_15600);
xor U16231 (N_16231,N_15944,N_15533);
xnor U16232 (N_16232,N_15693,N_15610);
and U16233 (N_16233,N_15755,N_15780);
or U16234 (N_16234,N_15653,N_15919);
xnor U16235 (N_16235,N_15622,N_15717);
and U16236 (N_16236,N_15504,N_15657);
or U16237 (N_16237,N_15728,N_15725);
and U16238 (N_16238,N_15832,N_15625);
or U16239 (N_16239,N_15710,N_15788);
or U16240 (N_16240,N_15942,N_15872);
and U16241 (N_16241,N_15946,N_15729);
nand U16242 (N_16242,N_15858,N_15688);
and U16243 (N_16243,N_15861,N_15998);
xnor U16244 (N_16244,N_15948,N_15532);
nor U16245 (N_16245,N_15799,N_15997);
or U16246 (N_16246,N_15580,N_15552);
or U16247 (N_16247,N_15565,N_15510);
or U16248 (N_16248,N_15761,N_15987);
xor U16249 (N_16249,N_15599,N_15744);
xor U16250 (N_16250,N_15963,N_15745);
xnor U16251 (N_16251,N_15541,N_15729);
xnor U16252 (N_16252,N_15581,N_15548);
nor U16253 (N_16253,N_15831,N_15666);
nor U16254 (N_16254,N_15965,N_15911);
or U16255 (N_16255,N_15887,N_15503);
nor U16256 (N_16256,N_15891,N_15924);
and U16257 (N_16257,N_15817,N_15603);
nand U16258 (N_16258,N_15760,N_15920);
xnor U16259 (N_16259,N_15654,N_15919);
nor U16260 (N_16260,N_15842,N_15781);
and U16261 (N_16261,N_15672,N_15554);
nand U16262 (N_16262,N_15557,N_15774);
and U16263 (N_16263,N_15984,N_15996);
nand U16264 (N_16264,N_15789,N_15799);
or U16265 (N_16265,N_15923,N_15984);
or U16266 (N_16266,N_15713,N_15884);
and U16267 (N_16267,N_15760,N_15533);
nor U16268 (N_16268,N_15619,N_15806);
or U16269 (N_16269,N_15942,N_15710);
nor U16270 (N_16270,N_15776,N_15566);
nand U16271 (N_16271,N_15869,N_15567);
and U16272 (N_16272,N_15769,N_15717);
or U16273 (N_16273,N_15870,N_15874);
or U16274 (N_16274,N_15720,N_15897);
xnor U16275 (N_16275,N_15631,N_15686);
xnor U16276 (N_16276,N_15882,N_15585);
and U16277 (N_16277,N_15738,N_15646);
xor U16278 (N_16278,N_15959,N_15812);
nor U16279 (N_16279,N_15887,N_15803);
or U16280 (N_16280,N_15505,N_15863);
or U16281 (N_16281,N_15740,N_15620);
nor U16282 (N_16282,N_15850,N_15684);
xnor U16283 (N_16283,N_15907,N_15788);
and U16284 (N_16284,N_15621,N_15669);
nor U16285 (N_16285,N_15723,N_15630);
xor U16286 (N_16286,N_15980,N_15752);
xor U16287 (N_16287,N_15802,N_15633);
or U16288 (N_16288,N_15938,N_15607);
and U16289 (N_16289,N_15898,N_15992);
nor U16290 (N_16290,N_15514,N_15525);
xor U16291 (N_16291,N_15564,N_15589);
or U16292 (N_16292,N_15680,N_15989);
and U16293 (N_16293,N_15551,N_15643);
nand U16294 (N_16294,N_15841,N_15655);
nor U16295 (N_16295,N_15845,N_15605);
or U16296 (N_16296,N_15527,N_15692);
nor U16297 (N_16297,N_15824,N_15808);
nor U16298 (N_16298,N_15604,N_15908);
xor U16299 (N_16299,N_15568,N_15540);
and U16300 (N_16300,N_15969,N_15564);
xnor U16301 (N_16301,N_15539,N_15679);
xnor U16302 (N_16302,N_15883,N_15712);
and U16303 (N_16303,N_15978,N_15764);
or U16304 (N_16304,N_15624,N_15602);
nand U16305 (N_16305,N_15695,N_15509);
xor U16306 (N_16306,N_15986,N_15899);
xor U16307 (N_16307,N_15881,N_15792);
or U16308 (N_16308,N_15890,N_15889);
xor U16309 (N_16309,N_15531,N_15638);
nand U16310 (N_16310,N_15998,N_15603);
and U16311 (N_16311,N_15825,N_15817);
and U16312 (N_16312,N_15919,N_15834);
nand U16313 (N_16313,N_15713,N_15734);
nor U16314 (N_16314,N_15877,N_15556);
and U16315 (N_16315,N_15628,N_15769);
and U16316 (N_16316,N_15977,N_15985);
nor U16317 (N_16317,N_15572,N_15763);
nor U16318 (N_16318,N_15999,N_15981);
nand U16319 (N_16319,N_15771,N_15741);
nor U16320 (N_16320,N_15926,N_15832);
nor U16321 (N_16321,N_15859,N_15755);
nor U16322 (N_16322,N_15576,N_15912);
and U16323 (N_16323,N_15640,N_15565);
or U16324 (N_16324,N_15819,N_15706);
nand U16325 (N_16325,N_15837,N_15518);
or U16326 (N_16326,N_15523,N_15516);
xnor U16327 (N_16327,N_15679,N_15577);
nor U16328 (N_16328,N_15647,N_15943);
or U16329 (N_16329,N_15711,N_15869);
or U16330 (N_16330,N_15653,N_15793);
and U16331 (N_16331,N_15898,N_15966);
and U16332 (N_16332,N_15811,N_15515);
xnor U16333 (N_16333,N_15841,N_15651);
or U16334 (N_16334,N_15625,N_15866);
and U16335 (N_16335,N_15989,N_15594);
or U16336 (N_16336,N_15684,N_15656);
nor U16337 (N_16337,N_15635,N_15807);
and U16338 (N_16338,N_15727,N_15681);
and U16339 (N_16339,N_15595,N_15837);
nand U16340 (N_16340,N_15689,N_15816);
nand U16341 (N_16341,N_15502,N_15656);
nand U16342 (N_16342,N_15951,N_15614);
nor U16343 (N_16343,N_15895,N_15604);
nor U16344 (N_16344,N_15919,N_15683);
and U16345 (N_16345,N_15783,N_15564);
nand U16346 (N_16346,N_15907,N_15876);
xor U16347 (N_16347,N_15553,N_15555);
nand U16348 (N_16348,N_15969,N_15852);
and U16349 (N_16349,N_15608,N_15581);
nor U16350 (N_16350,N_15652,N_15703);
and U16351 (N_16351,N_15625,N_15589);
xor U16352 (N_16352,N_15756,N_15838);
xnor U16353 (N_16353,N_15755,N_15533);
nor U16354 (N_16354,N_15682,N_15613);
nor U16355 (N_16355,N_15885,N_15519);
nand U16356 (N_16356,N_15598,N_15678);
or U16357 (N_16357,N_15950,N_15922);
nor U16358 (N_16358,N_15942,N_15650);
nor U16359 (N_16359,N_15841,N_15590);
xnor U16360 (N_16360,N_15793,N_15748);
or U16361 (N_16361,N_15844,N_15799);
nand U16362 (N_16362,N_15908,N_15911);
and U16363 (N_16363,N_15567,N_15508);
xor U16364 (N_16364,N_15552,N_15729);
or U16365 (N_16365,N_15841,N_15770);
nor U16366 (N_16366,N_15838,N_15689);
xnor U16367 (N_16367,N_15545,N_15526);
nand U16368 (N_16368,N_15514,N_15966);
xor U16369 (N_16369,N_15927,N_15715);
or U16370 (N_16370,N_15916,N_15963);
nor U16371 (N_16371,N_15983,N_15579);
and U16372 (N_16372,N_15795,N_15857);
and U16373 (N_16373,N_15761,N_15615);
or U16374 (N_16374,N_15655,N_15648);
and U16375 (N_16375,N_15837,N_15630);
or U16376 (N_16376,N_15810,N_15768);
nor U16377 (N_16377,N_15660,N_15889);
nand U16378 (N_16378,N_15690,N_15799);
and U16379 (N_16379,N_15735,N_15877);
xor U16380 (N_16380,N_15877,N_15936);
and U16381 (N_16381,N_15828,N_15929);
or U16382 (N_16382,N_15702,N_15593);
or U16383 (N_16383,N_15885,N_15831);
nor U16384 (N_16384,N_15764,N_15883);
or U16385 (N_16385,N_15507,N_15596);
nand U16386 (N_16386,N_15801,N_15656);
nor U16387 (N_16387,N_15812,N_15960);
xor U16388 (N_16388,N_15571,N_15834);
xnor U16389 (N_16389,N_15647,N_15986);
nor U16390 (N_16390,N_15919,N_15569);
or U16391 (N_16391,N_15801,N_15760);
or U16392 (N_16392,N_15525,N_15641);
nor U16393 (N_16393,N_15593,N_15974);
nand U16394 (N_16394,N_15977,N_15780);
xnor U16395 (N_16395,N_15576,N_15502);
nor U16396 (N_16396,N_15970,N_15674);
nor U16397 (N_16397,N_15785,N_15511);
xnor U16398 (N_16398,N_15859,N_15903);
nand U16399 (N_16399,N_15942,N_15589);
xor U16400 (N_16400,N_15895,N_15516);
nor U16401 (N_16401,N_15719,N_15595);
nor U16402 (N_16402,N_15965,N_15880);
or U16403 (N_16403,N_15899,N_15588);
nand U16404 (N_16404,N_15873,N_15897);
nand U16405 (N_16405,N_15685,N_15526);
or U16406 (N_16406,N_15592,N_15822);
or U16407 (N_16407,N_15781,N_15587);
nor U16408 (N_16408,N_15502,N_15725);
and U16409 (N_16409,N_15789,N_15790);
xnor U16410 (N_16410,N_15769,N_15889);
or U16411 (N_16411,N_15700,N_15559);
nand U16412 (N_16412,N_15657,N_15780);
nor U16413 (N_16413,N_15629,N_15950);
nor U16414 (N_16414,N_15719,N_15645);
nand U16415 (N_16415,N_15882,N_15773);
xnor U16416 (N_16416,N_15510,N_15646);
xnor U16417 (N_16417,N_15683,N_15503);
xnor U16418 (N_16418,N_15734,N_15858);
nor U16419 (N_16419,N_15681,N_15931);
and U16420 (N_16420,N_15937,N_15549);
nor U16421 (N_16421,N_15659,N_15727);
nand U16422 (N_16422,N_15614,N_15875);
nor U16423 (N_16423,N_15652,N_15533);
nor U16424 (N_16424,N_15913,N_15830);
nor U16425 (N_16425,N_15560,N_15513);
and U16426 (N_16426,N_15606,N_15920);
nor U16427 (N_16427,N_15851,N_15580);
xor U16428 (N_16428,N_15980,N_15669);
nand U16429 (N_16429,N_15570,N_15919);
nor U16430 (N_16430,N_15812,N_15740);
nor U16431 (N_16431,N_15748,N_15904);
or U16432 (N_16432,N_15653,N_15744);
or U16433 (N_16433,N_15566,N_15645);
nand U16434 (N_16434,N_15509,N_15580);
and U16435 (N_16435,N_15676,N_15966);
nor U16436 (N_16436,N_15575,N_15711);
and U16437 (N_16437,N_15741,N_15543);
or U16438 (N_16438,N_15792,N_15687);
xnor U16439 (N_16439,N_15733,N_15816);
nor U16440 (N_16440,N_15797,N_15940);
or U16441 (N_16441,N_15535,N_15968);
xnor U16442 (N_16442,N_15614,N_15631);
xnor U16443 (N_16443,N_15983,N_15620);
or U16444 (N_16444,N_15866,N_15962);
or U16445 (N_16445,N_15901,N_15703);
or U16446 (N_16446,N_15678,N_15829);
nand U16447 (N_16447,N_15687,N_15673);
nor U16448 (N_16448,N_15853,N_15828);
and U16449 (N_16449,N_15616,N_15639);
xor U16450 (N_16450,N_15705,N_15895);
nand U16451 (N_16451,N_15626,N_15802);
nand U16452 (N_16452,N_15913,N_15502);
and U16453 (N_16453,N_15595,N_15912);
and U16454 (N_16454,N_15823,N_15732);
nand U16455 (N_16455,N_15588,N_15806);
and U16456 (N_16456,N_15674,N_15638);
nand U16457 (N_16457,N_15887,N_15515);
xnor U16458 (N_16458,N_15541,N_15581);
or U16459 (N_16459,N_15713,N_15958);
nor U16460 (N_16460,N_15901,N_15877);
and U16461 (N_16461,N_15795,N_15781);
xor U16462 (N_16462,N_15996,N_15968);
nand U16463 (N_16463,N_15600,N_15867);
and U16464 (N_16464,N_15607,N_15897);
nand U16465 (N_16465,N_15752,N_15538);
and U16466 (N_16466,N_15541,N_15852);
nand U16467 (N_16467,N_15837,N_15869);
or U16468 (N_16468,N_15795,N_15750);
nand U16469 (N_16469,N_15796,N_15828);
xnor U16470 (N_16470,N_15595,N_15832);
nand U16471 (N_16471,N_15737,N_15632);
and U16472 (N_16472,N_15638,N_15792);
and U16473 (N_16473,N_15791,N_15608);
or U16474 (N_16474,N_15661,N_15837);
nor U16475 (N_16475,N_15748,N_15631);
and U16476 (N_16476,N_15805,N_15974);
xor U16477 (N_16477,N_15534,N_15778);
xor U16478 (N_16478,N_15906,N_15659);
nor U16479 (N_16479,N_15506,N_15707);
and U16480 (N_16480,N_15504,N_15678);
and U16481 (N_16481,N_15544,N_15564);
nor U16482 (N_16482,N_15956,N_15912);
xnor U16483 (N_16483,N_15660,N_15764);
nand U16484 (N_16484,N_15889,N_15993);
xor U16485 (N_16485,N_15633,N_15721);
nand U16486 (N_16486,N_15994,N_15534);
or U16487 (N_16487,N_15680,N_15597);
nand U16488 (N_16488,N_15666,N_15781);
nand U16489 (N_16489,N_15903,N_15728);
and U16490 (N_16490,N_15856,N_15611);
nand U16491 (N_16491,N_15502,N_15807);
nor U16492 (N_16492,N_15506,N_15528);
or U16493 (N_16493,N_15946,N_15627);
nor U16494 (N_16494,N_15701,N_15525);
xor U16495 (N_16495,N_15796,N_15543);
nor U16496 (N_16496,N_15859,N_15632);
nand U16497 (N_16497,N_15966,N_15886);
nand U16498 (N_16498,N_15987,N_15621);
or U16499 (N_16499,N_15994,N_15872);
nand U16500 (N_16500,N_16297,N_16069);
nand U16501 (N_16501,N_16389,N_16077);
or U16502 (N_16502,N_16393,N_16133);
and U16503 (N_16503,N_16129,N_16383);
nand U16504 (N_16504,N_16411,N_16064);
or U16505 (N_16505,N_16198,N_16169);
nor U16506 (N_16506,N_16179,N_16422);
nand U16507 (N_16507,N_16127,N_16194);
or U16508 (N_16508,N_16040,N_16280);
nand U16509 (N_16509,N_16227,N_16363);
and U16510 (N_16510,N_16080,N_16405);
nor U16511 (N_16511,N_16017,N_16081);
nand U16512 (N_16512,N_16023,N_16355);
nor U16513 (N_16513,N_16448,N_16335);
nor U16514 (N_16514,N_16395,N_16387);
nand U16515 (N_16515,N_16111,N_16073);
and U16516 (N_16516,N_16254,N_16273);
nor U16517 (N_16517,N_16088,N_16174);
xor U16518 (N_16518,N_16191,N_16244);
or U16519 (N_16519,N_16486,N_16249);
or U16520 (N_16520,N_16430,N_16454);
nand U16521 (N_16521,N_16431,N_16105);
or U16522 (N_16522,N_16022,N_16413);
nor U16523 (N_16523,N_16160,N_16250);
nand U16524 (N_16524,N_16106,N_16235);
and U16525 (N_16525,N_16154,N_16305);
and U16526 (N_16526,N_16240,N_16404);
xnor U16527 (N_16527,N_16139,N_16007);
nand U16528 (N_16528,N_16427,N_16217);
or U16529 (N_16529,N_16408,N_16074);
or U16530 (N_16530,N_16200,N_16177);
and U16531 (N_16531,N_16165,N_16376);
nand U16532 (N_16532,N_16110,N_16167);
and U16533 (N_16533,N_16156,N_16053);
nand U16534 (N_16534,N_16168,N_16175);
or U16535 (N_16535,N_16450,N_16409);
nor U16536 (N_16536,N_16406,N_16205);
nand U16537 (N_16537,N_16079,N_16418);
or U16538 (N_16538,N_16400,N_16157);
nor U16539 (N_16539,N_16076,N_16224);
and U16540 (N_16540,N_16123,N_16455);
and U16541 (N_16541,N_16050,N_16340);
xnor U16542 (N_16542,N_16365,N_16233);
or U16543 (N_16543,N_16102,N_16043);
and U16544 (N_16544,N_16483,N_16229);
nand U16545 (N_16545,N_16270,N_16095);
nor U16546 (N_16546,N_16407,N_16225);
or U16547 (N_16547,N_16461,N_16371);
xor U16548 (N_16548,N_16444,N_16159);
xor U16549 (N_16549,N_16412,N_16442);
nand U16550 (N_16550,N_16460,N_16281);
xor U16551 (N_16551,N_16319,N_16143);
or U16552 (N_16552,N_16014,N_16184);
nor U16553 (N_16553,N_16354,N_16417);
nor U16554 (N_16554,N_16187,N_16420);
or U16555 (N_16555,N_16377,N_16247);
nor U16556 (N_16556,N_16149,N_16024);
xor U16557 (N_16557,N_16309,N_16341);
or U16558 (N_16558,N_16364,N_16279);
xnor U16559 (N_16559,N_16001,N_16013);
nor U16560 (N_16560,N_16057,N_16269);
or U16561 (N_16561,N_16338,N_16379);
nor U16562 (N_16562,N_16031,N_16367);
and U16563 (N_16563,N_16181,N_16164);
nor U16564 (N_16564,N_16099,N_16325);
xor U16565 (N_16565,N_16401,N_16180);
xnor U16566 (N_16566,N_16055,N_16429);
xnor U16567 (N_16567,N_16182,N_16278);
and U16568 (N_16568,N_16234,N_16189);
or U16569 (N_16569,N_16343,N_16092);
nor U16570 (N_16570,N_16294,N_16476);
nor U16571 (N_16571,N_16265,N_16403);
nor U16572 (N_16572,N_16054,N_16000);
xor U16573 (N_16573,N_16202,N_16005);
and U16574 (N_16574,N_16494,N_16262);
or U16575 (N_16575,N_16375,N_16342);
or U16576 (N_16576,N_16004,N_16210);
nand U16577 (N_16577,N_16251,N_16370);
and U16578 (N_16578,N_16495,N_16231);
and U16579 (N_16579,N_16292,N_16109);
xor U16580 (N_16580,N_16246,N_16472);
nand U16581 (N_16581,N_16360,N_16300);
or U16582 (N_16582,N_16378,N_16333);
and U16583 (N_16583,N_16303,N_16438);
or U16584 (N_16584,N_16385,N_16314);
xnor U16585 (N_16585,N_16021,N_16259);
nand U16586 (N_16586,N_16298,N_16185);
and U16587 (N_16587,N_16415,N_16103);
nand U16588 (N_16588,N_16299,N_16451);
xor U16589 (N_16589,N_16214,N_16452);
or U16590 (N_16590,N_16318,N_16242);
xor U16591 (N_16591,N_16356,N_16489);
and U16592 (N_16592,N_16170,N_16045);
and U16593 (N_16593,N_16256,N_16381);
nand U16594 (N_16594,N_16394,N_16302);
nor U16595 (N_16595,N_16382,N_16222);
and U16596 (N_16596,N_16039,N_16380);
or U16597 (N_16597,N_16082,N_16130);
nor U16598 (N_16598,N_16087,N_16153);
xor U16599 (N_16599,N_16487,N_16331);
or U16600 (N_16600,N_16261,N_16386);
nor U16601 (N_16601,N_16197,N_16276);
nand U16602 (N_16602,N_16480,N_16195);
or U16603 (N_16603,N_16492,N_16332);
or U16604 (N_16604,N_16316,N_16308);
and U16605 (N_16605,N_16052,N_16232);
nor U16606 (N_16606,N_16439,N_16124);
or U16607 (N_16607,N_16078,N_16172);
or U16608 (N_16608,N_16146,N_16100);
nand U16609 (N_16609,N_16101,N_16090);
and U16610 (N_16610,N_16469,N_16238);
nand U16611 (N_16611,N_16361,N_16060);
nor U16612 (N_16612,N_16446,N_16042);
nand U16613 (N_16613,N_16277,N_16148);
xor U16614 (N_16614,N_16490,N_16009);
nor U16615 (N_16615,N_16061,N_16436);
and U16616 (N_16616,N_16034,N_16038);
nor U16617 (N_16617,N_16058,N_16288);
nand U16618 (N_16618,N_16132,N_16067);
nand U16619 (N_16619,N_16098,N_16253);
or U16620 (N_16620,N_16443,N_16398);
xor U16621 (N_16621,N_16134,N_16020);
or U16622 (N_16622,N_16230,N_16019);
or U16623 (N_16623,N_16243,N_16131);
xor U16624 (N_16624,N_16350,N_16018);
nand U16625 (N_16625,N_16028,N_16334);
nor U16626 (N_16626,N_16437,N_16056);
xor U16627 (N_16627,N_16268,N_16362);
nand U16628 (N_16628,N_16128,N_16328);
nor U16629 (N_16629,N_16388,N_16321);
nor U16630 (N_16630,N_16173,N_16093);
xnor U16631 (N_16631,N_16327,N_16208);
nor U16632 (N_16632,N_16215,N_16317);
nand U16633 (N_16633,N_16147,N_16207);
nand U16634 (N_16634,N_16104,N_16463);
xnor U16635 (N_16635,N_16245,N_16337);
nor U16636 (N_16636,N_16322,N_16445);
xor U16637 (N_16637,N_16065,N_16122);
and U16638 (N_16638,N_16479,N_16071);
xnor U16639 (N_16639,N_16390,N_16112);
or U16640 (N_16640,N_16324,N_16059);
nand U16641 (N_16641,N_16323,N_16135);
and U16642 (N_16642,N_16310,N_16041);
or U16643 (N_16643,N_16125,N_16313);
nand U16644 (N_16644,N_16199,N_16206);
xor U16645 (N_16645,N_16228,N_16115);
nor U16646 (N_16646,N_16025,N_16477);
nand U16647 (N_16647,N_16141,N_16188);
or U16648 (N_16648,N_16237,N_16347);
nand U16649 (N_16649,N_16307,N_16084);
xnor U16650 (N_16650,N_16008,N_16145);
nor U16651 (N_16651,N_16201,N_16274);
nor U16652 (N_16652,N_16044,N_16171);
and U16653 (N_16653,N_16330,N_16462);
nand U16654 (N_16654,N_16236,N_16116);
xnor U16655 (N_16655,N_16425,N_16449);
and U16656 (N_16656,N_16392,N_16326);
nor U16657 (N_16657,N_16290,N_16283);
nor U16658 (N_16658,N_16161,N_16289);
and U16659 (N_16659,N_16424,N_16275);
or U16660 (N_16660,N_16068,N_16284);
or U16661 (N_16661,N_16083,N_16315);
or U16662 (N_16662,N_16306,N_16359);
nor U16663 (N_16663,N_16351,N_16271);
nand U16664 (N_16664,N_16475,N_16121);
and U16665 (N_16665,N_16026,N_16296);
xor U16666 (N_16666,N_16155,N_16140);
nand U16667 (N_16667,N_16352,N_16484);
or U16668 (N_16668,N_16459,N_16282);
or U16669 (N_16669,N_16119,N_16311);
and U16670 (N_16670,N_16027,N_16464);
or U16671 (N_16671,N_16190,N_16163);
or U16672 (N_16672,N_16030,N_16485);
xor U16673 (N_16673,N_16440,N_16075);
and U16674 (N_16674,N_16183,N_16468);
or U16675 (N_16675,N_16416,N_16166);
or U16676 (N_16676,N_16258,N_16470);
nand U16677 (N_16677,N_16066,N_16032);
xnor U16678 (N_16678,N_16113,N_16441);
or U16679 (N_16679,N_16178,N_16349);
nor U16680 (N_16680,N_16272,N_16266);
or U16681 (N_16681,N_16397,N_16414);
or U16682 (N_16682,N_16482,N_16046);
and U16683 (N_16683,N_16036,N_16108);
nor U16684 (N_16684,N_16051,N_16366);
or U16685 (N_16685,N_16150,N_16072);
and U16686 (N_16686,N_16434,N_16496);
xnor U16687 (N_16687,N_16094,N_16357);
nor U16688 (N_16688,N_16037,N_16426);
or U16689 (N_16689,N_16118,N_16428);
nor U16690 (N_16690,N_16257,N_16493);
nor U16691 (N_16691,N_16295,N_16176);
and U16692 (N_16692,N_16291,N_16384);
nand U16693 (N_16693,N_16456,N_16186);
xnor U16694 (N_16694,N_16117,N_16089);
and U16695 (N_16695,N_16248,N_16474);
xor U16696 (N_16696,N_16301,N_16263);
and U16697 (N_16697,N_16458,N_16126);
nor U16698 (N_16698,N_16223,N_16120);
or U16699 (N_16699,N_16216,N_16062);
or U16700 (N_16700,N_16287,N_16264);
or U16701 (N_16701,N_16433,N_16252);
or U16702 (N_16702,N_16497,N_16304);
or U16703 (N_16703,N_16226,N_16086);
nand U16704 (N_16704,N_16312,N_16158);
or U16705 (N_16705,N_16465,N_16070);
and U16706 (N_16706,N_16035,N_16396);
xnor U16707 (N_16707,N_16419,N_16137);
nand U16708 (N_16708,N_16447,N_16011);
xnor U16709 (N_16709,N_16491,N_16348);
nor U16710 (N_16710,N_16218,N_16221);
nand U16711 (N_16711,N_16260,N_16471);
nand U16712 (N_16712,N_16285,N_16432);
and U16713 (N_16713,N_16402,N_16410);
or U16714 (N_16714,N_16091,N_16049);
and U16715 (N_16715,N_16466,N_16097);
nor U16716 (N_16716,N_16029,N_16033);
xor U16717 (N_16717,N_16346,N_16286);
and U16718 (N_16718,N_16255,N_16399);
nand U16719 (N_16719,N_16107,N_16015);
or U16720 (N_16720,N_16473,N_16293);
nand U16721 (N_16721,N_16423,N_16391);
xnor U16722 (N_16722,N_16003,N_16372);
nor U16723 (N_16723,N_16162,N_16138);
and U16724 (N_16724,N_16192,N_16012);
nand U16725 (N_16725,N_16114,N_16353);
or U16726 (N_16726,N_16336,N_16344);
xor U16727 (N_16727,N_16435,N_16329);
or U16728 (N_16728,N_16213,N_16239);
xnor U16729 (N_16729,N_16320,N_16453);
nand U16730 (N_16730,N_16142,N_16063);
xor U16731 (N_16731,N_16048,N_16203);
nor U16732 (N_16732,N_16096,N_16481);
nand U16733 (N_16733,N_16345,N_16369);
nor U16734 (N_16734,N_16211,N_16002);
or U16735 (N_16735,N_16219,N_16136);
nor U16736 (N_16736,N_16498,N_16499);
or U16737 (N_16737,N_16144,N_16010);
and U16738 (N_16738,N_16339,N_16358);
xor U16739 (N_16739,N_16421,N_16016);
or U16740 (N_16740,N_16006,N_16374);
nor U16741 (N_16741,N_16220,N_16368);
and U16742 (N_16742,N_16193,N_16488);
nand U16743 (N_16743,N_16085,N_16209);
nand U16744 (N_16744,N_16478,N_16047);
nor U16745 (N_16745,N_16151,N_16373);
nand U16746 (N_16746,N_16204,N_16196);
or U16747 (N_16747,N_16457,N_16212);
xnor U16748 (N_16748,N_16152,N_16467);
and U16749 (N_16749,N_16241,N_16267);
nand U16750 (N_16750,N_16043,N_16332);
nor U16751 (N_16751,N_16278,N_16458);
nand U16752 (N_16752,N_16332,N_16053);
nand U16753 (N_16753,N_16281,N_16105);
nor U16754 (N_16754,N_16316,N_16182);
nand U16755 (N_16755,N_16199,N_16009);
xor U16756 (N_16756,N_16473,N_16325);
nor U16757 (N_16757,N_16485,N_16062);
nand U16758 (N_16758,N_16345,N_16307);
nand U16759 (N_16759,N_16121,N_16099);
or U16760 (N_16760,N_16325,N_16242);
xnor U16761 (N_16761,N_16237,N_16161);
or U16762 (N_16762,N_16437,N_16121);
nand U16763 (N_16763,N_16258,N_16255);
nand U16764 (N_16764,N_16457,N_16287);
xor U16765 (N_16765,N_16174,N_16143);
xor U16766 (N_16766,N_16225,N_16357);
and U16767 (N_16767,N_16391,N_16463);
or U16768 (N_16768,N_16065,N_16134);
and U16769 (N_16769,N_16180,N_16434);
nor U16770 (N_16770,N_16460,N_16015);
or U16771 (N_16771,N_16027,N_16396);
nand U16772 (N_16772,N_16295,N_16443);
and U16773 (N_16773,N_16363,N_16171);
nor U16774 (N_16774,N_16281,N_16308);
nand U16775 (N_16775,N_16029,N_16117);
or U16776 (N_16776,N_16342,N_16048);
or U16777 (N_16777,N_16400,N_16189);
nand U16778 (N_16778,N_16256,N_16046);
xor U16779 (N_16779,N_16385,N_16401);
and U16780 (N_16780,N_16239,N_16023);
nand U16781 (N_16781,N_16341,N_16395);
and U16782 (N_16782,N_16062,N_16374);
xor U16783 (N_16783,N_16466,N_16427);
nand U16784 (N_16784,N_16212,N_16305);
nand U16785 (N_16785,N_16383,N_16429);
nor U16786 (N_16786,N_16457,N_16153);
or U16787 (N_16787,N_16426,N_16035);
xor U16788 (N_16788,N_16143,N_16047);
or U16789 (N_16789,N_16219,N_16438);
and U16790 (N_16790,N_16488,N_16334);
or U16791 (N_16791,N_16239,N_16416);
and U16792 (N_16792,N_16489,N_16472);
and U16793 (N_16793,N_16173,N_16335);
and U16794 (N_16794,N_16280,N_16174);
xor U16795 (N_16795,N_16318,N_16400);
and U16796 (N_16796,N_16378,N_16361);
or U16797 (N_16797,N_16272,N_16062);
nand U16798 (N_16798,N_16185,N_16136);
nor U16799 (N_16799,N_16390,N_16420);
and U16800 (N_16800,N_16015,N_16037);
or U16801 (N_16801,N_16280,N_16199);
or U16802 (N_16802,N_16377,N_16267);
nand U16803 (N_16803,N_16328,N_16335);
xor U16804 (N_16804,N_16447,N_16456);
nor U16805 (N_16805,N_16459,N_16018);
nor U16806 (N_16806,N_16007,N_16499);
nor U16807 (N_16807,N_16074,N_16041);
xnor U16808 (N_16808,N_16436,N_16499);
and U16809 (N_16809,N_16385,N_16410);
xnor U16810 (N_16810,N_16068,N_16099);
and U16811 (N_16811,N_16079,N_16399);
and U16812 (N_16812,N_16278,N_16408);
nand U16813 (N_16813,N_16448,N_16356);
nand U16814 (N_16814,N_16420,N_16309);
and U16815 (N_16815,N_16060,N_16177);
and U16816 (N_16816,N_16291,N_16272);
xor U16817 (N_16817,N_16422,N_16154);
and U16818 (N_16818,N_16068,N_16280);
and U16819 (N_16819,N_16368,N_16496);
nor U16820 (N_16820,N_16005,N_16354);
and U16821 (N_16821,N_16279,N_16190);
nor U16822 (N_16822,N_16027,N_16290);
or U16823 (N_16823,N_16330,N_16286);
and U16824 (N_16824,N_16171,N_16294);
xnor U16825 (N_16825,N_16440,N_16181);
and U16826 (N_16826,N_16328,N_16098);
xnor U16827 (N_16827,N_16117,N_16420);
nand U16828 (N_16828,N_16352,N_16369);
or U16829 (N_16829,N_16094,N_16103);
xnor U16830 (N_16830,N_16419,N_16135);
nor U16831 (N_16831,N_16475,N_16024);
nor U16832 (N_16832,N_16303,N_16356);
xor U16833 (N_16833,N_16313,N_16406);
and U16834 (N_16834,N_16232,N_16171);
nor U16835 (N_16835,N_16132,N_16247);
nand U16836 (N_16836,N_16328,N_16235);
xor U16837 (N_16837,N_16130,N_16405);
and U16838 (N_16838,N_16120,N_16297);
nor U16839 (N_16839,N_16158,N_16258);
nand U16840 (N_16840,N_16274,N_16064);
nor U16841 (N_16841,N_16255,N_16499);
and U16842 (N_16842,N_16054,N_16202);
nor U16843 (N_16843,N_16224,N_16025);
or U16844 (N_16844,N_16131,N_16309);
nand U16845 (N_16845,N_16475,N_16132);
and U16846 (N_16846,N_16006,N_16249);
or U16847 (N_16847,N_16300,N_16194);
xor U16848 (N_16848,N_16253,N_16033);
or U16849 (N_16849,N_16012,N_16264);
or U16850 (N_16850,N_16493,N_16105);
xnor U16851 (N_16851,N_16033,N_16165);
xor U16852 (N_16852,N_16348,N_16115);
xor U16853 (N_16853,N_16090,N_16079);
nand U16854 (N_16854,N_16236,N_16285);
and U16855 (N_16855,N_16492,N_16273);
or U16856 (N_16856,N_16254,N_16438);
nor U16857 (N_16857,N_16062,N_16249);
nand U16858 (N_16858,N_16179,N_16433);
nor U16859 (N_16859,N_16350,N_16283);
nand U16860 (N_16860,N_16401,N_16265);
xor U16861 (N_16861,N_16266,N_16021);
and U16862 (N_16862,N_16070,N_16430);
xnor U16863 (N_16863,N_16180,N_16076);
and U16864 (N_16864,N_16431,N_16320);
nor U16865 (N_16865,N_16157,N_16046);
nand U16866 (N_16866,N_16181,N_16106);
nor U16867 (N_16867,N_16203,N_16310);
and U16868 (N_16868,N_16443,N_16139);
xor U16869 (N_16869,N_16482,N_16247);
nand U16870 (N_16870,N_16098,N_16263);
and U16871 (N_16871,N_16001,N_16331);
xnor U16872 (N_16872,N_16191,N_16087);
and U16873 (N_16873,N_16394,N_16416);
nand U16874 (N_16874,N_16267,N_16000);
or U16875 (N_16875,N_16214,N_16001);
and U16876 (N_16876,N_16432,N_16001);
nor U16877 (N_16877,N_16062,N_16205);
xor U16878 (N_16878,N_16333,N_16476);
nor U16879 (N_16879,N_16298,N_16221);
or U16880 (N_16880,N_16448,N_16426);
nor U16881 (N_16881,N_16185,N_16043);
nand U16882 (N_16882,N_16459,N_16234);
nor U16883 (N_16883,N_16403,N_16397);
nand U16884 (N_16884,N_16039,N_16278);
nor U16885 (N_16885,N_16335,N_16439);
xor U16886 (N_16886,N_16298,N_16256);
or U16887 (N_16887,N_16358,N_16199);
nor U16888 (N_16888,N_16032,N_16014);
xnor U16889 (N_16889,N_16488,N_16474);
nor U16890 (N_16890,N_16195,N_16211);
and U16891 (N_16891,N_16358,N_16007);
xnor U16892 (N_16892,N_16237,N_16198);
xnor U16893 (N_16893,N_16026,N_16338);
xor U16894 (N_16894,N_16449,N_16360);
nand U16895 (N_16895,N_16044,N_16047);
nor U16896 (N_16896,N_16468,N_16347);
and U16897 (N_16897,N_16071,N_16455);
nand U16898 (N_16898,N_16328,N_16392);
nand U16899 (N_16899,N_16463,N_16103);
xnor U16900 (N_16900,N_16143,N_16069);
and U16901 (N_16901,N_16042,N_16312);
nor U16902 (N_16902,N_16249,N_16087);
nand U16903 (N_16903,N_16303,N_16182);
xnor U16904 (N_16904,N_16245,N_16192);
or U16905 (N_16905,N_16492,N_16490);
nand U16906 (N_16906,N_16063,N_16420);
nor U16907 (N_16907,N_16032,N_16381);
or U16908 (N_16908,N_16086,N_16422);
nor U16909 (N_16909,N_16427,N_16373);
or U16910 (N_16910,N_16092,N_16328);
nand U16911 (N_16911,N_16196,N_16149);
nand U16912 (N_16912,N_16213,N_16432);
and U16913 (N_16913,N_16283,N_16420);
nor U16914 (N_16914,N_16058,N_16394);
xnor U16915 (N_16915,N_16188,N_16155);
nor U16916 (N_16916,N_16438,N_16026);
or U16917 (N_16917,N_16090,N_16371);
or U16918 (N_16918,N_16423,N_16082);
xnor U16919 (N_16919,N_16222,N_16215);
and U16920 (N_16920,N_16296,N_16338);
xor U16921 (N_16921,N_16459,N_16213);
and U16922 (N_16922,N_16205,N_16417);
and U16923 (N_16923,N_16145,N_16330);
and U16924 (N_16924,N_16301,N_16279);
or U16925 (N_16925,N_16479,N_16383);
and U16926 (N_16926,N_16428,N_16270);
nor U16927 (N_16927,N_16370,N_16044);
nor U16928 (N_16928,N_16258,N_16489);
nand U16929 (N_16929,N_16230,N_16499);
and U16930 (N_16930,N_16432,N_16375);
xor U16931 (N_16931,N_16371,N_16166);
and U16932 (N_16932,N_16318,N_16388);
xor U16933 (N_16933,N_16171,N_16126);
xnor U16934 (N_16934,N_16169,N_16230);
or U16935 (N_16935,N_16010,N_16366);
nor U16936 (N_16936,N_16302,N_16483);
nor U16937 (N_16937,N_16422,N_16296);
xnor U16938 (N_16938,N_16126,N_16034);
nand U16939 (N_16939,N_16324,N_16182);
nor U16940 (N_16940,N_16234,N_16021);
nor U16941 (N_16941,N_16111,N_16358);
xnor U16942 (N_16942,N_16006,N_16048);
nor U16943 (N_16943,N_16374,N_16116);
nand U16944 (N_16944,N_16271,N_16476);
or U16945 (N_16945,N_16365,N_16269);
nand U16946 (N_16946,N_16477,N_16222);
nor U16947 (N_16947,N_16492,N_16304);
nand U16948 (N_16948,N_16097,N_16321);
nor U16949 (N_16949,N_16480,N_16076);
xnor U16950 (N_16950,N_16157,N_16176);
nand U16951 (N_16951,N_16299,N_16026);
nand U16952 (N_16952,N_16150,N_16262);
or U16953 (N_16953,N_16299,N_16379);
and U16954 (N_16954,N_16072,N_16436);
nand U16955 (N_16955,N_16026,N_16407);
or U16956 (N_16956,N_16484,N_16016);
or U16957 (N_16957,N_16382,N_16205);
nand U16958 (N_16958,N_16109,N_16130);
xor U16959 (N_16959,N_16347,N_16048);
xnor U16960 (N_16960,N_16295,N_16182);
or U16961 (N_16961,N_16128,N_16212);
and U16962 (N_16962,N_16189,N_16040);
or U16963 (N_16963,N_16097,N_16256);
nand U16964 (N_16964,N_16006,N_16252);
or U16965 (N_16965,N_16356,N_16462);
xnor U16966 (N_16966,N_16364,N_16281);
or U16967 (N_16967,N_16004,N_16335);
and U16968 (N_16968,N_16122,N_16263);
or U16969 (N_16969,N_16354,N_16071);
nor U16970 (N_16970,N_16171,N_16434);
nand U16971 (N_16971,N_16049,N_16288);
xor U16972 (N_16972,N_16081,N_16341);
and U16973 (N_16973,N_16038,N_16448);
nand U16974 (N_16974,N_16164,N_16060);
xor U16975 (N_16975,N_16171,N_16464);
nand U16976 (N_16976,N_16110,N_16313);
and U16977 (N_16977,N_16210,N_16368);
xnor U16978 (N_16978,N_16297,N_16347);
xor U16979 (N_16979,N_16152,N_16388);
nand U16980 (N_16980,N_16399,N_16267);
or U16981 (N_16981,N_16492,N_16434);
and U16982 (N_16982,N_16190,N_16100);
nor U16983 (N_16983,N_16249,N_16309);
or U16984 (N_16984,N_16400,N_16047);
and U16985 (N_16985,N_16271,N_16474);
and U16986 (N_16986,N_16337,N_16094);
or U16987 (N_16987,N_16022,N_16386);
or U16988 (N_16988,N_16415,N_16271);
and U16989 (N_16989,N_16105,N_16465);
and U16990 (N_16990,N_16384,N_16396);
nand U16991 (N_16991,N_16374,N_16011);
or U16992 (N_16992,N_16489,N_16481);
xnor U16993 (N_16993,N_16482,N_16227);
nor U16994 (N_16994,N_16414,N_16458);
xor U16995 (N_16995,N_16168,N_16132);
nand U16996 (N_16996,N_16252,N_16397);
and U16997 (N_16997,N_16175,N_16348);
xor U16998 (N_16998,N_16402,N_16441);
nor U16999 (N_16999,N_16395,N_16018);
nor U17000 (N_17000,N_16896,N_16800);
nor U17001 (N_17001,N_16940,N_16534);
nor U17002 (N_17002,N_16808,N_16691);
nand U17003 (N_17003,N_16576,N_16763);
nand U17004 (N_17004,N_16533,N_16816);
xnor U17005 (N_17005,N_16560,N_16875);
and U17006 (N_17006,N_16585,N_16858);
or U17007 (N_17007,N_16575,N_16636);
nor U17008 (N_17008,N_16837,N_16857);
or U17009 (N_17009,N_16684,N_16545);
nor U17010 (N_17010,N_16685,N_16941);
and U17011 (N_17011,N_16934,N_16726);
and U17012 (N_17012,N_16955,N_16775);
nand U17013 (N_17013,N_16944,N_16511);
xnor U17014 (N_17014,N_16503,N_16661);
and U17015 (N_17015,N_16989,N_16504);
nand U17016 (N_17016,N_16584,N_16796);
nand U17017 (N_17017,N_16531,N_16739);
and U17018 (N_17018,N_16566,N_16959);
xor U17019 (N_17019,N_16977,N_16785);
or U17020 (N_17020,N_16734,N_16624);
and U17021 (N_17021,N_16614,N_16530);
nor U17022 (N_17022,N_16819,N_16906);
xnor U17023 (N_17023,N_16957,N_16563);
and U17024 (N_17024,N_16604,N_16922);
nor U17025 (N_17025,N_16931,N_16956);
and U17026 (N_17026,N_16842,N_16998);
xnor U17027 (N_17027,N_16610,N_16778);
nand U17028 (N_17028,N_16539,N_16645);
nand U17029 (N_17029,N_16618,N_16973);
nor U17030 (N_17030,N_16911,N_16701);
or U17031 (N_17031,N_16501,N_16730);
and U17032 (N_17032,N_16917,N_16830);
or U17033 (N_17033,N_16523,N_16946);
nor U17034 (N_17034,N_16892,N_16916);
xor U17035 (N_17035,N_16707,N_16932);
and U17036 (N_17036,N_16861,N_16535);
xnor U17037 (N_17037,N_16804,N_16786);
or U17038 (N_17038,N_16652,N_16718);
xnor U17039 (N_17039,N_16666,N_16589);
nor U17040 (N_17040,N_16949,N_16655);
or U17041 (N_17041,N_16706,N_16822);
or U17042 (N_17042,N_16647,N_16769);
or U17043 (N_17043,N_16543,N_16554);
or U17044 (N_17044,N_16512,N_16960);
nand U17045 (N_17045,N_16635,N_16884);
and U17046 (N_17046,N_16650,N_16752);
or U17047 (N_17047,N_16926,N_16653);
xor U17048 (N_17048,N_16628,N_16735);
nand U17049 (N_17049,N_16901,N_16724);
or U17050 (N_17050,N_16755,N_16754);
or U17051 (N_17051,N_16799,N_16947);
xnor U17052 (N_17052,N_16626,N_16813);
xnor U17053 (N_17053,N_16620,N_16717);
nand U17054 (N_17054,N_16565,N_16849);
nor U17055 (N_17055,N_16728,N_16606);
nor U17056 (N_17056,N_16893,N_16880);
xnor U17057 (N_17057,N_16981,N_16985);
nand U17058 (N_17058,N_16818,N_16721);
nor U17059 (N_17059,N_16826,N_16725);
nor U17060 (N_17060,N_16526,N_16600);
nor U17061 (N_17061,N_16633,N_16648);
nand U17062 (N_17062,N_16747,N_16742);
and U17063 (N_17063,N_16748,N_16736);
xor U17064 (N_17064,N_16710,N_16513);
xnor U17065 (N_17065,N_16845,N_16757);
nor U17066 (N_17066,N_16783,N_16683);
nor U17067 (N_17067,N_16870,N_16608);
xnor U17068 (N_17068,N_16829,N_16966);
nand U17069 (N_17069,N_16988,N_16673);
or U17070 (N_17070,N_16638,N_16867);
nand U17071 (N_17071,N_16918,N_16743);
xnor U17072 (N_17072,N_16741,N_16928);
nand U17073 (N_17073,N_16525,N_16640);
or U17074 (N_17074,N_16553,N_16823);
nand U17075 (N_17075,N_16854,N_16510);
xor U17076 (N_17076,N_16781,N_16855);
xor U17077 (N_17077,N_16852,N_16711);
nor U17078 (N_17078,N_16883,N_16617);
and U17079 (N_17079,N_16549,N_16603);
nand U17080 (N_17080,N_16756,N_16943);
or U17081 (N_17081,N_16637,N_16997);
nor U17082 (N_17082,N_16679,N_16681);
nand U17083 (N_17083,N_16887,N_16676);
and U17084 (N_17084,N_16599,N_16987);
or U17085 (N_17085,N_16773,N_16851);
nand U17086 (N_17086,N_16557,N_16664);
and U17087 (N_17087,N_16570,N_16621);
or U17088 (N_17088,N_16662,N_16846);
or U17089 (N_17089,N_16992,N_16713);
and U17090 (N_17090,N_16882,N_16954);
or U17091 (N_17091,N_16625,N_16948);
nand U17092 (N_17092,N_16794,N_16874);
nand U17093 (N_17093,N_16871,N_16579);
or U17094 (N_17094,N_16587,N_16719);
and U17095 (N_17095,N_16853,N_16564);
or U17096 (N_17096,N_16933,N_16979);
xor U17097 (N_17097,N_16529,N_16657);
and U17098 (N_17098,N_16623,N_16792);
xnor U17099 (N_17099,N_16964,N_16695);
xnor U17100 (N_17100,N_16723,N_16542);
nor U17101 (N_17101,N_16612,N_16521);
or U17102 (N_17102,N_16990,N_16898);
nand U17103 (N_17103,N_16850,N_16528);
or U17104 (N_17104,N_16974,N_16862);
xor U17105 (N_17105,N_16962,N_16712);
and U17106 (N_17106,N_16975,N_16894);
and U17107 (N_17107,N_16651,N_16772);
nor U17108 (N_17108,N_16817,N_16594);
nor U17109 (N_17109,N_16924,N_16699);
xor U17110 (N_17110,N_16765,N_16895);
nor U17111 (N_17111,N_16642,N_16694);
or U17112 (N_17112,N_16868,N_16812);
nand U17113 (N_17113,N_16700,N_16688);
nor U17114 (N_17114,N_16629,N_16833);
nand U17115 (N_17115,N_16986,N_16703);
nor U17116 (N_17116,N_16680,N_16889);
nand U17117 (N_17117,N_16595,N_16537);
nand U17118 (N_17118,N_16961,N_16929);
xnor U17119 (N_17119,N_16945,N_16506);
or U17120 (N_17120,N_16507,N_16815);
or U17121 (N_17121,N_16574,N_16672);
xor U17122 (N_17122,N_16905,N_16939);
or U17123 (N_17123,N_16968,N_16878);
xor U17124 (N_17124,N_16784,N_16925);
xor U17125 (N_17125,N_16514,N_16908);
and U17126 (N_17126,N_16869,N_16779);
nor U17127 (N_17127,N_16978,N_16583);
and U17128 (N_17128,N_16890,N_16518);
xor U17129 (N_17129,N_16580,N_16984);
and U17130 (N_17130,N_16991,N_16588);
nor U17131 (N_17131,N_16809,N_16698);
nor U17132 (N_17132,N_16787,N_16971);
nand U17133 (N_17133,N_16750,N_16524);
xnor U17134 (N_17134,N_16611,N_16522);
or U17135 (N_17135,N_16722,N_16914);
nand U17136 (N_17136,N_16689,N_16505);
xnor U17137 (N_17137,N_16821,N_16631);
or U17138 (N_17138,N_16582,N_16668);
and U17139 (N_17139,N_16913,N_16716);
nor U17140 (N_17140,N_16831,N_16863);
nand U17141 (N_17141,N_16641,N_16798);
or U17142 (N_17142,N_16733,N_16644);
nand U17143 (N_17143,N_16619,N_16864);
or U17144 (N_17144,N_16745,N_16578);
and U17145 (N_17145,N_16630,N_16972);
or U17146 (N_17146,N_16865,N_16807);
and U17147 (N_17147,N_16659,N_16993);
xnor U17148 (N_17148,N_16788,N_16760);
nand U17149 (N_17149,N_16970,N_16705);
xnor U17150 (N_17150,N_16885,N_16935);
or U17151 (N_17151,N_16834,N_16544);
nor U17152 (N_17152,N_16586,N_16758);
or U17153 (N_17153,N_16793,N_16909);
or U17154 (N_17154,N_16923,N_16795);
and U17155 (N_17155,N_16872,N_16936);
nand U17156 (N_17156,N_16873,N_16824);
and U17157 (N_17157,N_16771,N_16670);
or U17158 (N_17158,N_16910,N_16886);
or U17159 (N_17159,N_16682,N_16904);
nand U17160 (N_17160,N_16519,N_16843);
xor U17161 (N_17161,N_16877,N_16556);
nand U17162 (N_17162,N_16841,N_16573);
or U17163 (N_17163,N_16654,N_16753);
and U17164 (N_17164,N_16592,N_16567);
nand U17165 (N_17165,N_16900,N_16561);
nand U17166 (N_17166,N_16791,N_16920);
nor U17167 (N_17167,N_16558,N_16622);
and U17168 (N_17168,N_16678,N_16801);
nand U17169 (N_17169,N_16782,N_16532);
nand U17170 (N_17170,N_16836,N_16616);
nand U17171 (N_17171,N_16761,N_16921);
or U17172 (N_17172,N_16562,N_16536);
nand U17173 (N_17173,N_16596,N_16520);
and U17174 (N_17174,N_16738,N_16996);
xor U17175 (N_17175,N_16967,N_16602);
and U17176 (N_17176,N_16593,N_16774);
nand U17177 (N_17177,N_16571,N_16903);
or U17178 (N_17178,N_16942,N_16615);
or U17179 (N_17179,N_16696,N_16559);
xnor U17180 (N_17180,N_16790,N_16983);
nand U17181 (N_17181,N_16714,N_16919);
and U17182 (N_17182,N_16601,N_16547);
and U17183 (N_17183,N_16540,N_16762);
and U17184 (N_17184,N_16999,N_16671);
xnor U17185 (N_17185,N_16667,N_16690);
nor U17186 (N_17186,N_16897,N_16749);
and U17187 (N_17187,N_16969,N_16768);
nand U17188 (N_17188,N_16777,N_16902);
or U17189 (N_17189,N_16881,N_16572);
or U17190 (N_17190,N_16839,N_16632);
nand U17191 (N_17191,N_16709,N_16744);
or U17192 (N_17192,N_16899,N_16825);
or U17193 (N_17193,N_16591,N_16789);
xor U17194 (N_17194,N_16767,N_16810);
xor U17195 (N_17195,N_16500,N_16692);
nor U17196 (N_17196,N_16720,N_16731);
nor U17197 (N_17197,N_16550,N_16879);
nor U17198 (N_17198,N_16976,N_16704);
and U17199 (N_17199,N_16737,N_16646);
nor U17200 (N_17200,N_16994,N_16891);
nor U17201 (N_17201,N_16953,N_16876);
nand U17202 (N_17202,N_16938,N_16627);
nand U17203 (N_17203,N_16590,N_16598);
nor U17204 (N_17204,N_16803,N_16927);
xor U17205 (N_17205,N_16832,N_16609);
and U17206 (N_17206,N_16546,N_16605);
and U17207 (N_17207,N_16766,N_16820);
xor U17208 (N_17208,N_16995,N_16963);
xnor U17209 (N_17209,N_16538,N_16828);
and U17210 (N_17210,N_16838,N_16780);
nand U17211 (N_17211,N_16727,N_16860);
nand U17212 (N_17212,N_16802,N_16859);
nor U17213 (N_17213,N_16658,N_16930);
xnor U17214 (N_17214,N_16607,N_16751);
nand U17215 (N_17215,N_16634,N_16674);
or U17216 (N_17216,N_16665,N_16915);
and U17217 (N_17217,N_16677,N_16643);
or U17218 (N_17218,N_16663,N_16950);
or U17219 (N_17219,N_16764,N_16888);
and U17220 (N_17220,N_16597,N_16555);
nor U17221 (N_17221,N_16848,N_16515);
nor U17222 (N_17222,N_16965,N_16568);
or U17223 (N_17223,N_16746,N_16982);
and U17224 (N_17224,N_16806,N_16776);
xnor U17225 (N_17225,N_16840,N_16814);
nand U17226 (N_17226,N_16856,N_16729);
and U17227 (N_17227,N_16639,N_16516);
xnor U17228 (N_17228,N_16805,N_16660);
nand U17229 (N_17229,N_16702,N_16669);
and U17230 (N_17230,N_16958,N_16656);
and U17231 (N_17231,N_16686,N_16759);
nor U17232 (N_17232,N_16509,N_16912);
and U17233 (N_17233,N_16827,N_16835);
nor U17234 (N_17234,N_16844,N_16866);
nand U17235 (N_17235,N_16697,N_16907);
xnor U17236 (N_17236,N_16937,N_16649);
nor U17237 (N_17237,N_16502,N_16951);
and U17238 (N_17238,N_16715,N_16693);
nand U17239 (N_17239,N_16508,N_16770);
nor U17240 (N_17240,N_16797,N_16517);
xnor U17241 (N_17241,N_16569,N_16708);
and U17242 (N_17242,N_16980,N_16581);
nor U17243 (N_17243,N_16527,N_16811);
nand U17244 (N_17244,N_16847,N_16551);
or U17245 (N_17245,N_16577,N_16687);
nand U17246 (N_17246,N_16952,N_16740);
nor U17247 (N_17247,N_16732,N_16541);
or U17248 (N_17248,N_16552,N_16675);
and U17249 (N_17249,N_16548,N_16613);
and U17250 (N_17250,N_16574,N_16677);
xnor U17251 (N_17251,N_16847,N_16959);
or U17252 (N_17252,N_16965,N_16651);
xnor U17253 (N_17253,N_16600,N_16905);
or U17254 (N_17254,N_16672,N_16950);
or U17255 (N_17255,N_16507,N_16973);
nand U17256 (N_17256,N_16578,N_16992);
or U17257 (N_17257,N_16744,N_16838);
nor U17258 (N_17258,N_16502,N_16679);
nor U17259 (N_17259,N_16514,N_16569);
nand U17260 (N_17260,N_16618,N_16546);
and U17261 (N_17261,N_16824,N_16775);
xor U17262 (N_17262,N_16913,N_16880);
nor U17263 (N_17263,N_16781,N_16633);
nor U17264 (N_17264,N_16678,N_16581);
or U17265 (N_17265,N_16660,N_16520);
or U17266 (N_17266,N_16695,N_16648);
nand U17267 (N_17267,N_16703,N_16602);
or U17268 (N_17268,N_16659,N_16935);
nor U17269 (N_17269,N_16650,N_16757);
or U17270 (N_17270,N_16875,N_16692);
and U17271 (N_17271,N_16542,N_16925);
nand U17272 (N_17272,N_16663,N_16754);
or U17273 (N_17273,N_16807,N_16720);
or U17274 (N_17274,N_16574,N_16586);
nor U17275 (N_17275,N_16928,N_16619);
or U17276 (N_17276,N_16959,N_16713);
or U17277 (N_17277,N_16980,N_16783);
nor U17278 (N_17278,N_16742,N_16829);
xnor U17279 (N_17279,N_16632,N_16837);
or U17280 (N_17280,N_16734,N_16627);
and U17281 (N_17281,N_16638,N_16913);
xor U17282 (N_17282,N_16653,N_16724);
and U17283 (N_17283,N_16892,N_16527);
nand U17284 (N_17284,N_16912,N_16712);
xnor U17285 (N_17285,N_16742,N_16688);
and U17286 (N_17286,N_16995,N_16834);
or U17287 (N_17287,N_16560,N_16949);
nand U17288 (N_17288,N_16977,N_16969);
xor U17289 (N_17289,N_16631,N_16679);
nor U17290 (N_17290,N_16714,N_16636);
or U17291 (N_17291,N_16942,N_16603);
nor U17292 (N_17292,N_16574,N_16957);
xnor U17293 (N_17293,N_16812,N_16726);
nand U17294 (N_17294,N_16568,N_16578);
nand U17295 (N_17295,N_16796,N_16865);
and U17296 (N_17296,N_16830,N_16860);
nand U17297 (N_17297,N_16887,N_16741);
or U17298 (N_17298,N_16703,N_16823);
or U17299 (N_17299,N_16820,N_16602);
xnor U17300 (N_17300,N_16994,N_16500);
and U17301 (N_17301,N_16631,N_16915);
xor U17302 (N_17302,N_16849,N_16803);
xnor U17303 (N_17303,N_16880,N_16983);
and U17304 (N_17304,N_16507,N_16918);
or U17305 (N_17305,N_16899,N_16530);
or U17306 (N_17306,N_16577,N_16604);
nand U17307 (N_17307,N_16937,N_16897);
or U17308 (N_17308,N_16872,N_16905);
and U17309 (N_17309,N_16975,N_16707);
xor U17310 (N_17310,N_16846,N_16586);
nor U17311 (N_17311,N_16624,N_16823);
nor U17312 (N_17312,N_16719,N_16586);
nor U17313 (N_17313,N_16924,N_16898);
xor U17314 (N_17314,N_16828,N_16508);
nor U17315 (N_17315,N_16875,N_16667);
nand U17316 (N_17316,N_16648,N_16552);
or U17317 (N_17317,N_16549,N_16701);
xor U17318 (N_17318,N_16826,N_16685);
or U17319 (N_17319,N_16561,N_16811);
nor U17320 (N_17320,N_16661,N_16658);
and U17321 (N_17321,N_16785,N_16914);
or U17322 (N_17322,N_16915,N_16667);
or U17323 (N_17323,N_16834,N_16588);
or U17324 (N_17324,N_16970,N_16574);
and U17325 (N_17325,N_16505,N_16922);
nand U17326 (N_17326,N_16814,N_16722);
nand U17327 (N_17327,N_16594,N_16761);
nand U17328 (N_17328,N_16544,N_16637);
xnor U17329 (N_17329,N_16582,N_16868);
nor U17330 (N_17330,N_16802,N_16922);
nand U17331 (N_17331,N_16891,N_16598);
or U17332 (N_17332,N_16564,N_16611);
xor U17333 (N_17333,N_16647,N_16934);
nand U17334 (N_17334,N_16702,N_16792);
nor U17335 (N_17335,N_16563,N_16898);
xor U17336 (N_17336,N_16588,N_16814);
nor U17337 (N_17337,N_16746,N_16912);
and U17338 (N_17338,N_16614,N_16608);
nand U17339 (N_17339,N_16907,N_16708);
or U17340 (N_17340,N_16806,N_16861);
nand U17341 (N_17341,N_16763,N_16682);
xor U17342 (N_17342,N_16697,N_16813);
xnor U17343 (N_17343,N_16786,N_16517);
xnor U17344 (N_17344,N_16710,N_16905);
nand U17345 (N_17345,N_16534,N_16887);
nand U17346 (N_17346,N_16990,N_16923);
nand U17347 (N_17347,N_16713,N_16771);
nor U17348 (N_17348,N_16767,N_16567);
or U17349 (N_17349,N_16598,N_16605);
and U17350 (N_17350,N_16905,N_16975);
xnor U17351 (N_17351,N_16614,N_16657);
and U17352 (N_17352,N_16991,N_16646);
and U17353 (N_17353,N_16501,N_16633);
or U17354 (N_17354,N_16554,N_16508);
and U17355 (N_17355,N_16913,N_16550);
nand U17356 (N_17356,N_16587,N_16513);
or U17357 (N_17357,N_16760,N_16882);
and U17358 (N_17358,N_16963,N_16588);
or U17359 (N_17359,N_16537,N_16992);
or U17360 (N_17360,N_16930,N_16976);
xor U17361 (N_17361,N_16657,N_16915);
xor U17362 (N_17362,N_16819,N_16940);
or U17363 (N_17363,N_16696,N_16747);
and U17364 (N_17364,N_16751,N_16866);
xnor U17365 (N_17365,N_16586,N_16633);
nor U17366 (N_17366,N_16601,N_16624);
xnor U17367 (N_17367,N_16707,N_16781);
nor U17368 (N_17368,N_16761,N_16978);
and U17369 (N_17369,N_16759,N_16834);
or U17370 (N_17370,N_16951,N_16866);
or U17371 (N_17371,N_16635,N_16811);
and U17372 (N_17372,N_16792,N_16574);
or U17373 (N_17373,N_16814,N_16584);
nand U17374 (N_17374,N_16841,N_16616);
xnor U17375 (N_17375,N_16843,N_16985);
nand U17376 (N_17376,N_16674,N_16730);
nand U17377 (N_17377,N_16800,N_16819);
xor U17378 (N_17378,N_16841,N_16529);
xor U17379 (N_17379,N_16862,N_16782);
xnor U17380 (N_17380,N_16792,N_16504);
nor U17381 (N_17381,N_16921,N_16986);
or U17382 (N_17382,N_16972,N_16774);
or U17383 (N_17383,N_16536,N_16638);
and U17384 (N_17384,N_16765,N_16596);
xnor U17385 (N_17385,N_16808,N_16972);
nand U17386 (N_17386,N_16526,N_16718);
or U17387 (N_17387,N_16831,N_16694);
or U17388 (N_17388,N_16698,N_16631);
nor U17389 (N_17389,N_16608,N_16628);
or U17390 (N_17390,N_16923,N_16942);
nor U17391 (N_17391,N_16994,N_16711);
and U17392 (N_17392,N_16582,N_16556);
or U17393 (N_17393,N_16576,N_16553);
and U17394 (N_17394,N_16748,N_16699);
nand U17395 (N_17395,N_16502,N_16980);
nor U17396 (N_17396,N_16872,N_16660);
nand U17397 (N_17397,N_16825,N_16978);
or U17398 (N_17398,N_16672,N_16706);
nor U17399 (N_17399,N_16821,N_16800);
or U17400 (N_17400,N_16909,N_16955);
nor U17401 (N_17401,N_16920,N_16647);
nor U17402 (N_17402,N_16701,N_16965);
nor U17403 (N_17403,N_16703,N_16800);
xor U17404 (N_17404,N_16981,N_16601);
nand U17405 (N_17405,N_16569,N_16541);
and U17406 (N_17406,N_16709,N_16783);
nor U17407 (N_17407,N_16818,N_16535);
and U17408 (N_17408,N_16507,N_16907);
nor U17409 (N_17409,N_16664,N_16544);
nor U17410 (N_17410,N_16837,N_16906);
and U17411 (N_17411,N_16518,N_16742);
or U17412 (N_17412,N_16810,N_16935);
xor U17413 (N_17413,N_16656,N_16645);
nor U17414 (N_17414,N_16815,N_16545);
or U17415 (N_17415,N_16935,N_16506);
xnor U17416 (N_17416,N_16689,N_16961);
nand U17417 (N_17417,N_16961,N_16507);
or U17418 (N_17418,N_16734,N_16945);
nor U17419 (N_17419,N_16818,N_16863);
or U17420 (N_17420,N_16932,N_16983);
xor U17421 (N_17421,N_16983,N_16612);
and U17422 (N_17422,N_16591,N_16839);
xor U17423 (N_17423,N_16922,N_16812);
or U17424 (N_17424,N_16837,N_16656);
and U17425 (N_17425,N_16870,N_16510);
nor U17426 (N_17426,N_16531,N_16606);
or U17427 (N_17427,N_16844,N_16620);
nand U17428 (N_17428,N_16595,N_16886);
and U17429 (N_17429,N_16967,N_16560);
nor U17430 (N_17430,N_16910,N_16515);
xor U17431 (N_17431,N_16638,N_16909);
nor U17432 (N_17432,N_16596,N_16560);
or U17433 (N_17433,N_16837,N_16858);
and U17434 (N_17434,N_16683,N_16967);
and U17435 (N_17435,N_16955,N_16521);
or U17436 (N_17436,N_16571,N_16935);
xor U17437 (N_17437,N_16592,N_16766);
and U17438 (N_17438,N_16674,N_16670);
nor U17439 (N_17439,N_16758,N_16920);
and U17440 (N_17440,N_16693,N_16560);
xnor U17441 (N_17441,N_16813,N_16750);
nor U17442 (N_17442,N_16651,N_16845);
nor U17443 (N_17443,N_16780,N_16947);
nor U17444 (N_17444,N_16799,N_16967);
xnor U17445 (N_17445,N_16631,N_16883);
xnor U17446 (N_17446,N_16741,N_16715);
nand U17447 (N_17447,N_16935,N_16918);
nor U17448 (N_17448,N_16748,N_16717);
or U17449 (N_17449,N_16680,N_16507);
nor U17450 (N_17450,N_16577,N_16677);
xor U17451 (N_17451,N_16852,N_16622);
nor U17452 (N_17452,N_16952,N_16713);
nor U17453 (N_17453,N_16998,N_16934);
or U17454 (N_17454,N_16545,N_16906);
xnor U17455 (N_17455,N_16735,N_16711);
xor U17456 (N_17456,N_16981,N_16834);
and U17457 (N_17457,N_16517,N_16710);
xor U17458 (N_17458,N_16660,N_16921);
nand U17459 (N_17459,N_16653,N_16535);
xor U17460 (N_17460,N_16520,N_16988);
nand U17461 (N_17461,N_16990,N_16622);
nand U17462 (N_17462,N_16658,N_16598);
nand U17463 (N_17463,N_16856,N_16617);
and U17464 (N_17464,N_16758,N_16714);
nor U17465 (N_17465,N_16662,N_16574);
xor U17466 (N_17466,N_16507,N_16594);
nor U17467 (N_17467,N_16588,N_16674);
nand U17468 (N_17468,N_16974,N_16665);
and U17469 (N_17469,N_16764,N_16563);
xor U17470 (N_17470,N_16561,N_16839);
xnor U17471 (N_17471,N_16966,N_16590);
xnor U17472 (N_17472,N_16878,N_16632);
or U17473 (N_17473,N_16681,N_16795);
nand U17474 (N_17474,N_16666,N_16562);
and U17475 (N_17475,N_16861,N_16757);
xor U17476 (N_17476,N_16603,N_16655);
xnor U17477 (N_17477,N_16645,N_16788);
nor U17478 (N_17478,N_16808,N_16864);
nor U17479 (N_17479,N_16952,N_16805);
or U17480 (N_17480,N_16743,N_16665);
xnor U17481 (N_17481,N_16536,N_16864);
and U17482 (N_17482,N_16766,N_16705);
nor U17483 (N_17483,N_16770,N_16517);
nor U17484 (N_17484,N_16556,N_16974);
xnor U17485 (N_17485,N_16729,N_16527);
and U17486 (N_17486,N_16521,N_16925);
nor U17487 (N_17487,N_16601,N_16521);
xor U17488 (N_17488,N_16976,N_16895);
nor U17489 (N_17489,N_16515,N_16924);
and U17490 (N_17490,N_16882,N_16896);
nand U17491 (N_17491,N_16850,N_16789);
xnor U17492 (N_17492,N_16519,N_16735);
and U17493 (N_17493,N_16501,N_16555);
nor U17494 (N_17494,N_16511,N_16708);
nand U17495 (N_17495,N_16569,N_16822);
nor U17496 (N_17496,N_16620,N_16688);
nand U17497 (N_17497,N_16801,N_16743);
or U17498 (N_17498,N_16618,N_16945);
or U17499 (N_17499,N_16571,N_16714);
and U17500 (N_17500,N_17282,N_17105);
and U17501 (N_17501,N_17413,N_17198);
and U17502 (N_17502,N_17455,N_17378);
xnor U17503 (N_17503,N_17442,N_17172);
nor U17504 (N_17504,N_17489,N_17152);
xnor U17505 (N_17505,N_17066,N_17011);
and U17506 (N_17506,N_17322,N_17113);
and U17507 (N_17507,N_17313,N_17386);
or U17508 (N_17508,N_17159,N_17070);
or U17509 (N_17509,N_17437,N_17047);
xnor U17510 (N_17510,N_17209,N_17171);
xor U17511 (N_17511,N_17382,N_17167);
and U17512 (N_17512,N_17057,N_17216);
nor U17513 (N_17513,N_17075,N_17220);
or U17514 (N_17514,N_17032,N_17132);
nand U17515 (N_17515,N_17016,N_17466);
nand U17516 (N_17516,N_17059,N_17324);
xor U17517 (N_17517,N_17223,N_17284);
or U17518 (N_17518,N_17402,N_17488);
nor U17519 (N_17519,N_17243,N_17131);
and U17520 (N_17520,N_17036,N_17088);
and U17521 (N_17521,N_17205,N_17069);
xnor U17522 (N_17522,N_17161,N_17136);
nor U17523 (N_17523,N_17250,N_17174);
nand U17524 (N_17524,N_17229,N_17221);
nand U17525 (N_17525,N_17078,N_17026);
and U17526 (N_17526,N_17380,N_17496);
xnor U17527 (N_17527,N_17118,N_17404);
nand U17528 (N_17528,N_17037,N_17043);
xor U17529 (N_17529,N_17003,N_17332);
or U17530 (N_17530,N_17438,N_17308);
nor U17531 (N_17531,N_17231,N_17014);
nand U17532 (N_17532,N_17232,N_17317);
and U17533 (N_17533,N_17129,N_17352);
xor U17534 (N_17534,N_17117,N_17477);
or U17535 (N_17535,N_17010,N_17389);
nand U17536 (N_17536,N_17293,N_17370);
nand U17537 (N_17537,N_17120,N_17044);
and U17538 (N_17538,N_17429,N_17381);
xnor U17539 (N_17539,N_17416,N_17082);
and U17540 (N_17540,N_17056,N_17168);
nor U17541 (N_17541,N_17298,N_17089);
and U17542 (N_17542,N_17201,N_17025);
and U17543 (N_17543,N_17028,N_17270);
or U17544 (N_17544,N_17369,N_17435);
or U17545 (N_17545,N_17158,N_17235);
nand U17546 (N_17546,N_17187,N_17185);
nand U17547 (N_17547,N_17417,N_17111);
nor U17548 (N_17548,N_17050,N_17004);
xor U17549 (N_17549,N_17049,N_17234);
nand U17550 (N_17550,N_17134,N_17375);
xnor U17551 (N_17551,N_17412,N_17206);
and U17552 (N_17552,N_17268,N_17385);
nand U17553 (N_17553,N_17343,N_17067);
or U17554 (N_17554,N_17263,N_17482);
and U17555 (N_17555,N_17051,N_17331);
nand U17556 (N_17556,N_17106,N_17207);
nor U17557 (N_17557,N_17012,N_17362);
nor U17558 (N_17558,N_17068,N_17304);
xnor U17559 (N_17559,N_17169,N_17017);
nor U17560 (N_17560,N_17176,N_17361);
and U17561 (N_17561,N_17251,N_17238);
nor U17562 (N_17562,N_17009,N_17367);
nand U17563 (N_17563,N_17421,N_17296);
xnor U17564 (N_17564,N_17023,N_17247);
nand U17565 (N_17565,N_17290,N_17264);
xnor U17566 (N_17566,N_17170,N_17276);
xnor U17567 (N_17567,N_17253,N_17432);
and U17568 (N_17568,N_17143,N_17471);
and U17569 (N_17569,N_17408,N_17191);
nor U17570 (N_17570,N_17237,N_17186);
and U17571 (N_17571,N_17301,N_17395);
nor U17572 (N_17572,N_17262,N_17195);
or U17573 (N_17573,N_17436,N_17485);
nand U17574 (N_17574,N_17156,N_17230);
or U17575 (N_17575,N_17193,N_17355);
or U17576 (N_17576,N_17394,N_17165);
and U17577 (N_17577,N_17203,N_17085);
or U17578 (N_17578,N_17020,N_17063);
or U17579 (N_17579,N_17181,N_17288);
nand U17580 (N_17580,N_17312,N_17080);
xnor U17581 (N_17581,N_17034,N_17336);
xor U17582 (N_17582,N_17439,N_17388);
and U17583 (N_17583,N_17039,N_17052);
nor U17584 (N_17584,N_17227,N_17151);
nor U17585 (N_17585,N_17015,N_17103);
nor U17586 (N_17586,N_17473,N_17374);
nand U17587 (N_17587,N_17122,N_17107);
xor U17588 (N_17588,N_17101,N_17495);
or U17589 (N_17589,N_17024,N_17498);
and U17590 (N_17590,N_17194,N_17147);
nand U17591 (N_17591,N_17445,N_17218);
xnor U17592 (N_17592,N_17456,N_17222);
or U17593 (N_17593,N_17319,N_17157);
xor U17594 (N_17594,N_17487,N_17449);
nand U17595 (N_17595,N_17210,N_17054);
nand U17596 (N_17596,N_17470,N_17360);
nor U17597 (N_17597,N_17182,N_17283);
or U17598 (N_17598,N_17465,N_17040);
xor U17599 (N_17599,N_17329,N_17358);
nand U17600 (N_17600,N_17000,N_17245);
nor U17601 (N_17601,N_17259,N_17104);
nand U17602 (N_17602,N_17046,N_17398);
or U17603 (N_17603,N_17476,N_17430);
or U17604 (N_17604,N_17166,N_17249);
nand U17605 (N_17605,N_17379,N_17490);
or U17606 (N_17606,N_17341,N_17196);
nor U17607 (N_17607,N_17347,N_17001);
and U17608 (N_17608,N_17178,N_17190);
and U17609 (N_17609,N_17225,N_17390);
nand U17610 (N_17610,N_17224,N_17325);
and U17611 (N_17611,N_17373,N_17002);
nand U17612 (N_17612,N_17365,N_17140);
xnor U17613 (N_17613,N_17095,N_17256);
nor U17614 (N_17614,N_17060,N_17180);
nor U17615 (N_17615,N_17109,N_17200);
nand U17616 (N_17616,N_17215,N_17440);
nor U17617 (N_17617,N_17266,N_17255);
xor U17618 (N_17618,N_17345,N_17213);
nor U17619 (N_17619,N_17314,N_17204);
xor U17620 (N_17620,N_17330,N_17302);
nand U17621 (N_17621,N_17226,N_17139);
and U17622 (N_17622,N_17123,N_17099);
or U17623 (N_17623,N_17072,N_17300);
and U17624 (N_17624,N_17141,N_17108);
or U17625 (N_17625,N_17474,N_17353);
xnor U17626 (N_17626,N_17354,N_17124);
or U17627 (N_17627,N_17297,N_17497);
or U17628 (N_17628,N_17045,N_17184);
nor U17629 (N_17629,N_17457,N_17348);
nor U17630 (N_17630,N_17071,N_17499);
xor U17631 (N_17631,N_17125,N_17393);
nand U17632 (N_17632,N_17338,N_17400);
nor U17633 (N_17633,N_17464,N_17252);
nand U17634 (N_17634,N_17019,N_17031);
nor U17635 (N_17635,N_17008,N_17278);
or U17636 (N_17636,N_17469,N_17146);
and U17637 (N_17637,N_17177,N_17115);
xor U17638 (N_17638,N_17423,N_17428);
or U17639 (N_17639,N_17461,N_17397);
nand U17640 (N_17640,N_17081,N_17384);
nand U17641 (N_17641,N_17275,N_17486);
xor U17642 (N_17642,N_17160,N_17260);
or U17643 (N_17643,N_17053,N_17042);
nand U17644 (N_17644,N_17173,N_17350);
nor U17645 (N_17645,N_17292,N_17406);
nor U17646 (N_17646,N_17006,N_17383);
xor U17647 (N_17647,N_17309,N_17175);
nor U17648 (N_17648,N_17133,N_17018);
and U17649 (N_17649,N_17097,N_17422);
nand U17650 (N_17650,N_17463,N_17116);
or U17651 (N_17651,N_17007,N_17217);
or U17652 (N_17652,N_17299,N_17119);
nor U17653 (N_17653,N_17038,N_17077);
and U17654 (N_17654,N_17327,N_17443);
and U17655 (N_17655,N_17092,N_17492);
or U17656 (N_17656,N_17448,N_17022);
nand U17657 (N_17657,N_17419,N_17315);
xor U17658 (N_17658,N_17079,N_17441);
nor U17659 (N_17659,N_17005,N_17310);
xnor U17660 (N_17660,N_17162,N_17407);
xnor U17661 (N_17661,N_17340,N_17246);
and U17662 (N_17662,N_17468,N_17326);
nand U17663 (N_17663,N_17418,N_17472);
xor U17664 (N_17664,N_17065,N_17493);
nand U17665 (N_17665,N_17294,N_17074);
xor U17666 (N_17666,N_17228,N_17055);
nor U17667 (N_17667,N_17346,N_17392);
nor U17668 (N_17668,N_17265,N_17414);
and U17669 (N_17669,N_17121,N_17269);
xor U17670 (N_17670,N_17100,N_17149);
or U17671 (N_17671,N_17183,N_17127);
or U17672 (N_17672,N_17316,N_17277);
nor U17673 (N_17673,N_17164,N_17454);
and U17674 (N_17674,N_17258,N_17144);
nor U17675 (N_17675,N_17145,N_17459);
and U17676 (N_17676,N_17285,N_17013);
and U17677 (N_17677,N_17202,N_17344);
nand U17678 (N_17678,N_17377,N_17188);
xor U17679 (N_17679,N_17321,N_17475);
nor U17680 (N_17680,N_17391,N_17096);
xor U17681 (N_17681,N_17356,N_17371);
xor U17682 (N_17682,N_17110,N_17199);
or U17683 (N_17683,N_17357,N_17084);
xor U17684 (N_17684,N_17318,N_17211);
nand U17685 (N_17685,N_17098,N_17112);
nor U17686 (N_17686,N_17163,N_17363);
nor U17687 (N_17687,N_17433,N_17453);
nor U17688 (N_17688,N_17281,N_17076);
nand U17689 (N_17689,N_17090,N_17148);
nand U17690 (N_17690,N_17086,N_17431);
nor U17691 (N_17691,N_17307,N_17359);
nor U17692 (N_17692,N_17286,N_17287);
nor U17693 (N_17693,N_17420,N_17102);
and U17694 (N_17694,N_17279,N_17335);
nor U17695 (N_17695,N_17236,N_17244);
and U17696 (N_17696,N_17219,N_17150);
and U17697 (N_17697,N_17444,N_17267);
nand U17698 (N_17698,N_17271,N_17342);
nand U17699 (N_17699,N_17087,N_17242);
nor U17700 (N_17700,N_17323,N_17058);
xnor U17701 (N_17701,N_17272,N_17403);
nor U17702 (N_17702,N_17368,N_17334);
nor U17703 (N_17703,N_17254,N_17376);
xnor U17704 (N_17704,N_17452,N_17467);
xor U17705 (N_17705,N_17434,N_17339);
nand U17706 (N_17706,N_17303,N_17179);
or U17707 (N_17707,N_17426,N_17241);
or U17708 (N_17708,N_17154,N_17083);
or U17709 (N_17709,N_17349,N_17479);
and U17710 (N_17710,N_17130,N_17447);
nand U17711 (N_17711,N_17295,N_17411);
nand U17712 (N_17712,N_17484,N_17399);
and U17713 (N_17713,N_17239,N_17305);
nor U17714 (N_17714,N_17481,N_17483);
nand U17715 (N_17715,N_17189,N_17333);
xnor U17716 (N_17716,N_17409,N_17289);
nor U17717 (N_17717,N_17048,N_17212);
xor U17718 (N_17718,N_17451,N_17274);
and U17719 (N_17719,N_17280,N_17030);
or U17720 (N_17720,N_17491,N_17257);
nand U17721 (N_17721,N_17311,N_17041);
nand U17722 (N_17722,N_17091,N_17138);
nand U17723 (N_17723,N_17460,N_17273);
xnor U17724 (N_17724,N_17197,N_17450);
nand U17725 (N_17725,N_17320,N_17458);
xor U17726 (N_17726,N_17446,N_17061);
and U17727 (N_17727,N_17233,N_17064);
or U17728 (N_17728,N_17291,N_17073);
and U17729 (N_17729,N_17029,N_17478);
and U17730 (N_17730,N_17135,N_17427);
nand U17731 (N_17731,N_17337,N_17480);
nand U17732 (N_17732,N_17396,N_17062);
nand U17733 (N_17733,N_17208,N_17410);
or U17734 (N_17734,N_17387,N_17366);
and U17735 (N_17735,N_17137,N_17021);
xnor U17736 (N_17736,N_17261,N_17128);
and U17737 (N_17737,N_17153,N_17462);
nand U17738 (N_17738,N_17328,N_17425);
xor U17739 (N_17739,N_17415,N_17306);
or U17740 (N_17740,N_17192,N_17494);
and U17741 (N_17741,N_17240,N_17126);
xor U17742 (N_17742,N_17093,N_17094);
or U17743 (N_17743,N_17027,N_17033);
nand U17744 (N_17744,N_17248,N_17035);
nand U17745 (N_17745,N_17401,N_17142);
nand U17746 (N_17746,N_17155,N_17114);
xor U17747 (N_17747,N_17405,N_17372);
nor U17748 (N_17748,N_17424,N_17364);
nor U17749 (N_17749,N_17351,N_17214);
xor U17750 (N_17750,N_17473,N_17076);
or U17751 (N_17751,N_17473,N_17134);
nor U17752 (N_17752,N_17381,N_17202);
xor U17753 (N_17753,N_17175,N_17332);
nor U17754 (N_17754,N_17411,N_17242);
or U17755 (N_17755,N_17123,N_17428);
xor U17756 (N_17756,N_17296,N_17418);
nor U17757 (N_17757,N_17097,N_17421);
and U17758 (N_17758,N_17499,N_17126);
and U17759 (N_17759,N_17174,N_17364);
and U17760 (N_17760,N_17156,N_17277);
and U17761 (N_17761,N_17155,N_17460);
or U17762 (N_17762,N_17440,N_17250);
xor U17763 (N_17763,N_17417,N_17178);
nand U17764 (N_17764,N_17027,N_17103);
and U17765 (N_17765,N_17336,N_17314);
and U17766 (N_17766,N_17194,N_17065);
nor U17767 (N_17767,N_17387,N_17381);
and U17768 (N_17768,N_17031,N_17217);
nand U17769 (N_17769,N_17418,N_17318);
and U17770 (N_17770,N_17175,N_17344);
nor U17771 (N_17771,N_17280,N_17441);
nor U17772 (N_17772,N_17210,N_17169);
or U17773 (N_17773,N_17397,N_17254);
nor U17774 (N_17774,N_17306,N_17302);
nand U17775 (N_17775,N_17462,N_17286);
or U17776 (N_17776,N_17319,N_17488);
and U17777 (N_17777,N_17191,N_17143);
xnor U17778 (N_17778,N_17131,N_17253);
nand U17779 (N_17779,N_17085,N_17429);
or U17780 (N_17780,N_17113,N_17387);
nand U17781 (N_17781,N_17428,N_17178);
and U17782 (N_17782,N_17036,N_17134);
nand U17783 (N_17783,N_17172,N_17221);
or U17784 (N_17784,N_17383,N_17014);
nor U17785 (N_17785,N_17488,N_17137);
nor U17786 (N_17786,N_17338,N_17109);
nor U17787 (N_17787,N_17431,N_17441);
or U17788 (N_17788,N_17482,N_17334);
nor U17789 (N_17789,N_17233,N_17037);
nor U17790 (N_17790,N_17297,N_17021);
and U17791 (N_17791,N_17156,N_17256);
xnor U17792 (N_17792,N_17444,N_17410);
or U17793 (N_17793,N_17229,N_17466);
and U17794 (N_17794,N_17469,N_17227);
or U17795 (N_17795,N_17475,N_17128);
or U17796 (N_17796,N_17206,N_17346);
and U17797 (N_17797,N_17043,N_17067);
and U17798 (N_17798,N_17385,N_17426);
nand U17799 (N_17799,N_17469,N_17377);
and U17800 (N_17800,N_17318,N_17120);
and U17801 (N_17801,N_17081,N_17074);
or U17802 (N_17802,N_17366,N_17439);
nor U17803 (N_17803,N_17061,N_17303);
nor U17804 (N_17804,N_17118,N_17110);
nand U17805 (N_17805,N_17190,N_17244);
or U17806 (N_17806,N_17449,N_17457);
nor U17807 (N_17807,N_17328,N_17061);
xor U17808 (N_17808,N_17239,N_17039);
or U17809 (N_17809,N_17066,N_17381);
and U17810 (N_17810,N_17322,N_17108);
or U17811 (N_17811,N_17222,N_17013);
nand U17812 (N_17812,N_17409,N_17199);
nand U17813 (N_17813,N_17311,N_17265);
and U17814 (N_17814,N_17474,N_17182);
or U17815 (N_17815,N_17435,N_17139);
nor U17816 (N_17816,N_17090,N_17230);
or U17817 (N_17817,N_17266,N_17203);
xnor U17818 (N_17818,N_17403,N_17287);
xor U17819 (N_17819,N_17378,N_17191);
and U17820 (N_17820,N_17125,N_17230);
nor U17821 (N_17821,N_17245,N_17247);
nor U17822 (N_17822,N_17266,N_17084);
nand U17823 (N_17823,N_17162,N_17368);
nor U17824 (N_17824,N_17005,N_17291);
nor U17825 (N_17825,N_17224,N_17196);
xnor U17826 (N_17826,N_17135,N_17265);
xor U17827 (N_17827,N_17314,N_17420);
or U17828 (N_17828,N_17260,N_17138);
xor U17829 (N_17829,N_17412,N_17281);
xnor U17830 (N_17830,N_17122,N_17217);
and U17831 (N_17831,N_17148,N_17138);
nor U17832 (N_17832,N_17069,N_17233);
or U17833 (N_17833,N_17064,N_17379);
nand U17834 (N_17834,N_17271,N_17038);
nand U17835 (N_17835,N_17161,N_17455);
and U17836 (N_17836,N_17292,N_17242);
or U17837 (N_17837,N_17259,N_17070);
nor U17838 (N_17838,N_17055,N_17133);
and U17839 (N_17839,N_17252,N_17359);
or U17840 (N_17840,N_17183,N_17314);
nor U17841 (N_17841,N_17496,N_17422);
nor U17842 (N_17842,N_17084,N_17216);
nand U17843 (N_17843,N_17478,N_17428);
nor U17844 (N_17844,N_17241,N_17133);
nand U17845 (N_17845,N_17220,N_17179);
or U17846 (N_17846,N_17345,N_17491);
nand U17847 (N_17847,N_17344,N_17354);
or U17848 (N_17848,N_17258,N_17416);
xnor U17849 (N_17849,N_17365,N_17327);
or U17850 (N_17850,N_17441,N_17124);
xnor U17851 (N_17851,N_17427,N_17302);
nor U17852 (N_17852,N_17412,N_17329);
nor U17853 (N_17853,N_17140,N_17405);
nor U17854 (N_17854,N_17142,N_17042);
nor U17855 (N_17855,N_17075,N_17358);
xnor U17856 (N_17856,N_17389,N_17330);
nand U17857 (N_17857,N_17240,N_17170);
or U17858 (N_17858,N_17349,N_17340);
nor U17859 (N_17859,N_17271,N_17492);
xor U17860 (N_17860,N_17316,N_17106);
or U17861 (N_17861,N_17241,N_17002);
and U17862 (N_17862,N_17424,N_17436);
nand U17863 (N_17863,N_17147,N_17351);
and U17864 (N_17864,N_17389,N_17220);
xor U17865 (N_17865,N_17064,N_17451);
or U17866 (N_17866,N_17129,N_17341);
or U17867 (N_17867,N_17190,N_17431);
xnor U17868 (N_17868,N_17257,N_17028);
and U17869 (N_17869,N_17204,N_17236);
nand U17870 (N_17870,N_17186,N_17119);
nor U17871 (N_17871,N_17153,N_17410);
nand U17872 (N_17872,N_17040,N_17219);
or U17873 (N_17873,N_17047,N_17252);
nand U17874 (N_17874,N_17245,N_17243);
xnor U17875 (N_17875,N_17305,N_17071);
or U17876 (N_17876,N_17333,N_17464);
nand U17877 (N_17877,N_17023,N_17178);
nand U17878 (N_17878,N_17244,N_17385);
or U17879 (N_17879,N_17004,N_17496);
and U17880 (N_17880,N_17169,N_17424);
or U17881 (N_17881,N_17064,N_17230);
or U17882 (N_17882,N_17084,N_17445);
xor U17883 (N_17883,N_17273,N_17194);
and U17884 (N_17884,N_17226,N_17270);
or U17885 (N_17885,N_17492,N_17489);
or U17886 (N_17886,N_17426,N_17200);
nand U17887 (N_17887,N_17498,N_17138);
xor U17888 (N_17888,N_17097,N_17177);
nor U17889 (N_17889,N_17417,N_17472);
or U17890 (N_17890,N_17338,N_17125);
nor U17891 (N_17891,N_17010,N_17175);
and U17892 (N_17892,N_17038,N_17425);
xnor U17893 (N_17893,N_17329,N_17325);
nor U17894 (N_17894,N_17387,N_17497);
or U17895 (N_17895,N_17292,N_17300);
nor U17896 (N_17896,N_17242,N_17037);
nand U17897 (N_17897,N_17421,N_17488);
nor U17898 (N_17898,N_17382,N_17082);
and U17899 (N_17899,N_17333,N_17121);
nand U17900 (N_17900,N_17312,N_17200);
nor U17901 (N_17901,N_17287,N_17358);
nor U17902 (N_17902,N_17491,N_17267);
or U17903 (N_17903,N_17025,N_17030);
or U17904 (N_17904,N_17072,N_17145);
xor U17905 (N_17905,N_17089,N_17328);
nor U17906 (N_17906,N_17486,N_17086);
nor U17907 (N_17907,N_17176,N_17199);
and U17908 (N_17908,N_17433,N_17286);
and U17909 (N_17909,N_17323,N_17086);
nor U17910 (N_17910,N_17388,N_17340);
xor U17911 (N_17911,N_17378,N_17399);
nor U17912 (N_17912,N_17125,N_17414);
xor U17913 (N_17913,N_17183,N_17442);
or U17914 (N_17914,N_17117,N_17359);
xnor U17915 (N_17915,N_17389,N_17031);
or U17916 (N_17916,N_17007,N_17041);
nor U17917 (N_17917,N_17304,N_17153);
nor U17918 (N_17918,N_17477,N_17128);
nand U17919 (N_17919,N_17279,N_17083);
xnor U17920 (N_17920,N_17312,N_17461);
nor U17921 (N_17921,N_17336,N_17352);
xnor U17922 (N_17922,N_17254,N_17196);
xor U17923 (N_17923,N_17031,N_17162);
nand U17924 (N_17924,N_17433,N_17036);
nor U17925 (N_17925,N_17341,N_17228);
nand U17926 (N_17926,N_17453,N_17214);
xnor U17927 (N_17927,N_17306,N_17173);
nand U17928 (N_17928,N_17287,N_17240);
xor U17929 (N_17929,N_17019,N_17022);
and U17930 (N_17930,N_17038,N_17410);
nor U17931 (N_17931,N_17499,N_17022);
and U17932 (N_17932,N_17230,N_17084);
and U17933 (N_17933,N_17138,N_17196);
nand U17934 (N_17934,N_17353,N_17019);
nor U17935 (N_17935,N_17251,N_17039);
nor U17936 (N_17936,N_17227,N_17287);
and U17937 (N_17937,N_17342,N_17404);
or U17938 (N_17938,N_17458,N_17466);
and U17939 (N_17939,N_17369,N_17077);
nand U17940 (N_17940,N_17017,N_17281);
nand U17941 (N_17941,N_17057,N_17347);
or U17942 (N_17942,N_17163,N_17258);
nand U17943 (N_17943,N_17026,N_17481);
xnor U17944 (N_17944,N_17398,N_17456);
nand U17945 (N_17945,N_17173,N_17091);
nor U17946 (N_17946,N_17420,N_17106);
nor U17947 (N_17947,N_17123,N_17125);
or U17948 (N_17948,N_17420,N_17327);
nor U17949 (N_17949,N_17427,N_17394);
or U17950 (N_17950,N_17476,N_17047);
xnor U17951 (N_17951,N_17351,N_17121);
xor U17952 (N_17952,N_17405,N_17301);
nand U17953 (N_17953,N_17313,N_17303);
or U17954 (N_17954,N_17231,N_17329);
nand U17955 (N_17955,N_17005,N_17320);
or U17956 (N_17956,N_17389,N_17290);
and U17957 (N_17957,N_17045,N_17434);
or U17958 (N_17958,N_17322,N_17144);
nor U17959 (N_17959,N_17357,N_17439);
and U17960 (N_17960,N_17041,N_17048);
nor U17961 (N_17961,N_17451,N_17037);
and U17962 (N_17962,N_17339,N_17079);
xor U17963 (N_17963,N_17001,N_17123);
nand U17964 (N_17964,N_17175,N_17485);
xor U17965 (N_17965,N_17222,N_17453);
nand U17966 (N_17966,N_17056,N_17162);
or U17967 (N_17967,N_17157,N_17101);
nand U17968 (N_17968,N_17341,N_17472);
nand U17969 (N_17969,N_17031,N_17264);
nand U17970 (N_17970,N_17438,N_17414);
xnor U17971 (N_17971,N_17319,N_17362);
xnor U17972 (N_17972,N_17327,N_17272);
nor U17973 (N_17973,N_17181,N_17310);
nor U17974 (N_17974,N_17285,N_17041);
xnor U17975 (N_17975,N_17034,N_17377);
nor U17976 (N_17976,N_17385,N_17260);
nor U17977 (N_17977,N_17397,N_17257);
xor U17978 (N_17978,N_17143,N_17054);
nor U17979 (N_17979,N_17415,N_17260);
xor U17980 (N_17980,N_17395,N_17210);
xnor U17981 (N_17981,N_17391,N_17077);
nor U17982 (N_17982,N_17290,N_17228);
xor U17983 (N_17983,N_17446,N_17241);
xnor U17984 (N_17984,N_17127,N_17162);
and U17985 (N_17985,N_17074,N_17275);
nor U17986 (N_17986,N_17494,N_17408);
or U17987 (N_17987,N_17093,N_17024);
or U17988 (N_17988,N_17188,N_17337);
or U17989 (N_17989,N_17402,N_17098);
xor U17990 (N_17990,N_17466,N_17036);
nand U17991 (N_17991,N_17016,N_17138);
and U17992 (N_17992,N_17334,N_17356);
xnor U17993 (N_17993,N_17406,N_17295);
nand U17994 (N_17994,N_17036,N_17013);
nor U17995 (N_17995,N_17291,N_17165);
nor U17996 (N_17996,N_17332,N_17407);
and U17997 (N_17997,N_17304,N_17381);
xor U17998 (N_17998,N_17280,N_17477);
or U17999 (N_17999,N_17141,N_17260);
nand U18000 (N_18000,N_17664,N_17651);
or U18001 (N_18001,N_17976,N_17569);
and U18002 (N_18002,N_17905,N_17719);
or U18003 (N_18003,N_17791,N_17622);
xnor U18004 (N_18004,N_17812,N_17689);
nor U18005 (N_18005,N_17534,N_17598);
xnor U18006 (N_18006,N_17885,N_17959);
or U18007 (N_18007,N_17659,N_17724);
or U18008 (N_18008,N_17743,N_17736);
and U18009 (N_18009,N_17560,N_17803);
or U18010 (N_18010,N_17815,N_17605);
and U18011 (N_18011,N_17876,N_17553);
nand U18012 (N_18012,N_17541,N_17741);
and U18013 (N_18013,N_17878,N_17817);
or U18014 (N_18014,N_17846,N_17708);
xnor U18015 (N_18015,N_17980,N_17747);
nand U18016 (N_18016,N_17582,N_17643);
and U18017 (N_18017,N_17686,N_17562);
and U18018 (N_18018,N_17587,N_17754);
or U18019 (N_18019,N_17536,N_17678);
nor U18020 (N_18020,N_17910,N_17839);
nor U18021 (N_18021,N_17793,N_17662);
or U18022 (N_18022,N_17833,N_17915);
and U18023 (N_18023,N_17813,N_17775);
nand U18024 (N_18024,N_17852,N_17781);
xor U18025 (N_18025,N_17575,N_17933);
and U18026 (N_18026,N_17973,N_17772);
nor U18027 (N_18027,N_17840,N_17897);
xnor U18028 (N_18028,N_17591,N_17932);
and U18029 (N_18029,N_17695,N_17668);
and U18030 (N_18030,N_17784,N_17554);
or U18031 (N_18031,N_17821,N_17956);
nand U18032 (N_18032,N_17913,N_17880);
and U18033 (N_18033,N_17751,N_17700);
and U18034 (N_18034,N_17967,N_17794);
nand U18035 (N_18035,N_17893,N_17685);
and U18036 (N_18036,N_17525,N_17938);
and U18037 (N_18037,N_17584,N_17916);
nand U18038 (N_18038,N_17944,N_17675);
or U18039 (N_18039,N_17998,N_17638);
xor U18040 (N_18040,N_17861,N_17513);
and U18041 (N_18041,N_17504,N_17807);
nor U18042 (N_18042,N_17767,N_17986);
xor U18043 (N_18043,N_17646,N_17609);
and U18044 (N_18044,N_17515,N_17978);
nor U18045 (N_18045,N_17538,N_17723);
xor U18046 (N_18046,N_17969,N_17863);
nor U18047 (N_18047,N_17540,N_17750);
and U18048 (N_18048,N_17629,N_17691);
or U18049 (N_18049,N_17838,N_17583);
nor U18050 (N_18050,N_17697,N_17542);
nor U18051 (N_18051,N_17982,N_17581);
or U18052 (N_18052,N_17883,N_17529);
nor U18053 (N_18053,N_17955,N_17585);
nand U18054 (N_18054,N_17626,N_17783);
nor U18055 (N_18055,N_17602,N_17924);
or U18056 (N_18056,N_17901,N_17687);
nor U18057 (N_18057,N_17755,N_17623);
xnor U18058 (N_18058,N_17782,N_17669);
or U18059 (N_18059,N_17828,N_17665);
xnor U18060 (N_18060,N_17844,N_17672);
xnor U18061 (N_18061,N_17725,N_17818);
nor U18062 (N_18062,N_17884,N_17537);
xor U18063 (N_18063,N_17929,N_17552);
nand U18064 (N_18064,N_17713,N_17709);
or U18065 (N_18065,N_17765,N_17548);
nor U18066 (N_18066,N_17522,N_17683);
or U18067 (N_18067,N_17710,N_17787);
nand U18068 (N_18068,N_17640,N_17653);
nand U18069 (N_18069,N_17612,N_17912);
nand U18070 (N_18070,N_17991,N_17699);
xor U18071 (N_18071,N_17706,N_17798);
or U18072 (N_18072,N_17825,N_17737);
xnor U18073 (N_18073,N_17777,N_17788);
xor U18074 (N_18074,N_17879,N_17805);
nor U18075 (N_18075,N_17610,N_17845);
and U18076 (N_18076,N_17799,N_17501);
and U18077 (N_18077,N_17759,N_17822);
nand U18078 (N_18078,N_17981,N_17512);
xor U18079 (N_18079,N_17667,N_17567);
xnor U18080 (N_18080,N_17946,N_17826);
nor U18081 (N_18081,N_17832,N_17628);
nand U18082 (N_18082,N_17677,N_17875);
or U18083 (N_18083,N_17680,N_17649);
and U18084 (N_18084,N_17892,N_17977);
and U18085 (N_18085,N_17881,N_17722);
nand U18086 (N_18086,N_17681,N_17958);
or U18087 (N_18087,N_17570,N_17682);
nor U18088 (N_18088,N_17596,N_17556);
or U18089 (N_18089,N_17975,N_17843);
nor U18090 (N_18090,N_17898,N_17589);
xnor U18091 (N_18091,N_17972,N_17608);
or U18092 (N_18092,N_17731,N_17939);
or U18093 (N_18093,N_17831,N_17714);
xor U18094 (N_18094,N_17907,N_17797);
nand U18095 (N_18095,N_17851,N_17717);
and U18096 (N_18096,N_17827,N_17999);
xor U18097 (N_18097,N_17874,N_17864);
and U18098 (N_18098,N_17847,N_17850);
nor U18099 (N_18099,N_17568,N_17524);
nand U18100 (N_18100,N_17992,N_17745);
and U18101 (N_18101,N_17547,N_17670);
and U18102 (N_18102,N_17948,N_17510);
or U18103 (N_18103,N_17776,N_17964);
nand U18104 (N_18104,N_17518,N_17962);
xnor U18105 (N_18105,N_17987,N_17579);
or U18106 (N_18106,N_17871,N_17648);
and U18107 (N_18107,N_17970,N_17774);
nor U18108 (N_18108,N_17533,N_17882);
nand U18109 (N_18109,N_17592,N_17974);
nand U18110 (N_18110,N_17597,N_17923);
or U18111 (N_18111,N_17746,N_17740);
nand U18112 (N_18112,N_17661,N_17641);
or U18113 (N_18113,N_17961,N_17925);
nand U18114 (N_18114,N_17823,N_17773);
or U18115 (N_18115,N_17989,N_17849);
or U18116 (N_18116,N_17914,N_17645);
xor U18117 (N_18117,N_17888,N_17919);
nor U18118 (N_18118,N_17634,N_17853);
nor U18119 (N_18119,N_17792,N_17808);
nand U18120 (N_18120,N_17877,N_17588);
nand U18121 (N_18121,N_17637,N_17804);
nor U18122 (N_18122,N_17993,N_17559);
or U18123 (N_18123,N_17715,N_17656);
xnor U18124 (N_18124,N_17756,N_17997);
nor U18125 (N_18125,N_17809,N_17968);
nand U18126 (N_18126,N_17894,N_17701);
xor U18127 (N_18127,N_17618,N_17632);
nor U18128 (N_18128,N_17721,N_17927);
and U18129 (N_18129,N_17786,N_17523);
or U18130 (N_18130,N_17862,N_17505);
nand U18131 (N_18131,N_17620,N_17551);
nor U18132 (N_18132,N_17996,N_17684);
or U18133 (N_18133,N_17720,N_17899);
nand U18134 (N_18134,N_17762,N_17744);
nor U18135 (N_18135,N_17950,N_17814);
nand U18136 (N_18136,N_17800,N_17544);
or U18137 (N_18137,N_17930,N_17995);
nor U18138 (N_18138,N_17866,N_17696);
nor U18139 (N_18139,N_17577,N_17702);
nand U18140 (N_18140,N_17984,N_17621);
or U18141 (N_18141,N_17752,N_17937);
nand U18142 (N_18142,N_17819,N_17748);
nand U18143 (N_18143,N_17574,N_17966);
and U18144 (N_18144,N_17855,N_17566);
xor U18145 (N_18145,N_17558,N_17789);
nand U18146 (N_18146,N_17539,N_17726);
and U18147 (N_18147,N_17769,N_17858);
and U18148 (N_18148,N_17636,N_17945);
and U18149 (N_18149,N_17698,N_17619);
and U18150 (N_18150,N_17896,N_17988);
nand U18151 (N_18151,N_17902,N_17834);
and U18152 (N_18152,N_17796,N_17642);
or U18153 (N_18153,N_17688,N_17630);
xor U18154 (N_18154,N_17546,N_17514);
nand U18155 (N_18155,N_17705,N_17650);
or U18156 (N_18156,N_17860,N_17761);
and U18157 (N_18157,N_17857,N_17604);
nor U18158 (N_18158,N_17942,N_17595);
nor U18159 (N_18159,N_17795,N_17811);
and U18160 (N_18160,N_17571,N_17671);
nand U18161 (N_18161,N_17749,N_17531);
nand U18162 (N_18162,N_17704,N_17507);
nand U18163 (N_18163,N_17509,N_17586);
or U18164 (N_18164,N_17594,N_17564);
nand U18165 (N_18165,N_17886,N_17763);
nand U18166 (N_18166,N_17841,N_17528);
nand U18167 (N_18167,N_17949,N_17517);
nand U18168 (N_18168,N_17526,N_17947);
nor U18169 (N_18169,N_17868,N_17790);
nand U18170 (N_18170,N_17895,N_17545);
nor U18171 (N_18171,N_17519,N_17960);
nor U18172 (N_18172,N_17644,N_17936);
nand U18173 (N_18173,N_17918,N_17718);
and U18174 (N_18174,N_17733,N_17611);
xor U18175 (N_18175,N_17829,N_17830);
or U18176 (N_18176,N_17511,N_17957);
or U18177 (N_18177,N_17920,N_17965);
nor U18178 (N_18178,N_17909,N_17854);
xor U18179 (N_18179,N_17785,N_17867);
and U18180 (N_18180,N_17806,N_17676);
and U18181 (N_18181,N_17703,N_17666);
xor U18182 (N_18182,N_17951,N_17768);
nor U18183 (N_18183,N_17613,N_17801);
nand U18184 (N_18184,N_17931,N_17917);
xor U18185 (N_18185,N_17766,N_17658);
nor U18186 (N_18186,N_17565,N_17660);
and U18187 (N_18187,N_17624,N_17625);
nand U18188 (N_18188,N_17607,N_17563);
and U18189 (N_18189,N_17707,N_17810);
and U18190 (N_18190,N_17940,N_17837);
or U18191 (N_18191,N_17663,N_17963);
or U18192 (N_18192,N_17983,N_17764);
nand U18193 (N_18193,N_17779,N_17780);
and U18194 (N_18194,N_17657,N_17599);
nor U18195 (N_18195,N_17728,N_17820);
or U18196 (N_18196,N_17652,N_17500);
and U18197 (N_18197,N_17716,N_17502);
nor U18198 (N_18198,N_17971,N_17994);
nor U18199 (N_18199,N_17758,N_17617);
xnor U18200 (N_18200,N_17616,N_17603);
and U18201 (N_18201,N_17906,N_17601);
nand U18202 (N_18202,N_17941,N_17836);
and U18203 (N_18203,N_17614,N_17848);
or U18204 (N_18204,N_17631,N_17859);
nor U18205 (N_18205,N_17615,N_17921);
nor U18206 (N_18206,N_17727,N_17690);
and U18207 (N_18207,N_17979,N_17580);
nand U18208 (N_18208,N_17856,N_17865);
and U18209 (N_18209,N_17954,N_17985);
and U18210 (N_18210,N_17816,N_17550);
nand U18211 (N_18211,N_17757,N_17889);
and U18212 (N_18212,N_17633,N_17742);
xor U18213 (N_18213,N_17576,N_17647);
or U18214 (N_18214,N_17770,N_17760);
and U18215 (N_18215,N_17928,N_17900);
nor U18216 (N_18216,N_17869,N_17872);
nor U18217 (N_18217,N_17887,N_17935);
and U18218 (N_18218,N_17903,N_17655);
nor U18219 (N_18219,N_17926,N_17654);
or U18220 (N_18220,N_17911,N_17890);
and U18221 (N_18221,N_17934,N_17835);
and U18222 (N_18222,N_17572,N_17952);
xnor U18223 (N_18223,N_17557,N_17503);
nor U18224 (N_18224,N_17870,N_17549);
and U18225 (N_18225,N_17692,N_17543);
nor U18226 (N_18226,N_17730,N_17590);
or U18227 (N_18227,N_17527,N_17508);
or U18228 (N_18228,N_17694,N_17530);
nor U18229 (N_18229,N_17735,N_17639);
or U18230 (N_18230,N_17738,N_17674);
xnor U18231 (N_18231,N_17516,N_17842);
xor U18232 (N_18232,N_17600,N_17943);
or U18233 (N_18233,N_17673,N_17778);
xnor U18234 (N_18234,N_17753,N_17739);
nand U18235 (N_18235,N_17904,N_17990);
and U18236 (N_18236,N_17578,N_17593);
nor U18237 (N_18237,N_17711,N_17635);
and U18238 (N_18238,N_17824,N_17535);
xor U18239 (N_18239,N_17532,N_17732);
nor U18240 (N_18240,N_17873,N_17953);
or U18241 (N_18241,N_17734,N_17606);
nor U18242 (N_18242,N_17922,N_17771);
or U18243 (N_18243,N_17555,N_17908);
nor U18244 (N_18244,N_17891,N_17520);
nor U18245 (N_18245,N_17802,N_17693);
and U18246 (N_18246,N_17561,N_17521);
xor U18247 (N_18247,N_17573,N_17506);
and U18248 (N_18248,N_17679,N_17729);
nor U18249 (N_18249,N_17712,N_17627);
and U18250 (N_18250,N_17863,N_17886);
or U18251 (N_18251,N_17964,N_17939);
xor U18252 (N_18252,N_17579,N_17696);
nand U18253 (N_18253,N_17530,N_17679);
nor U18254 (N_18254,N_17589,N_17601);
xor U18255 (N_18255,N_17780,N_17748);
xor U18256 (N_18256,N_17564,N_17639);
nand U18257 (N_18257,N_17776,N_17933);
or U18258 (N_18258,N_17760,N_17651);
nor U18259 (N_18259,N_17938,N_17638);
and U18260 (N_18260,N_17761,N_17898);
and U18261 (N_18261,N_17509,N_17773);
nor U18262 (N_18262,N_17691,N_17964);
or U18263 (N_18263,N_17958,N_17980);
and U18264 (N_18264,N_17939,N_17747);
nor U18265 (N_18265,N_17526,N_17634);
and U18266 (N_18266,N_17774,N_17570);
xor U18267 (N_18267,N_17927,N_17539);
nand U18268 (N_18268,N_17598,N_17562);
xor U18269 (N_18269,N_17984,N_17898);
nand U18270 (N_18270,N_17932,N_17784);
xnor U18271 (N_18271,N_17856,N_17697);
nand U18272 (N_18272,N_17873,N_17847);
nand U18273 (N_18273,N_17513,N_17630);
or U18274 (N_18274,N_17548,N_17734);
xnor U18275 (N_18275,N_17541,N_17771);
and U18276 (N_18276,N_17744,N_17966);
or U18277 (N_18277,N_17630,N_17762);
or U18278 (N_18278,N_17653,N_17857);
and U18279 (N_18279,N_17693,N_17505);
xor U18280 (N_18280,N_17902,N_17616);
xor U18281 (N_18281,N_17975,N_17649);
or U18282 (N_18282,N_17554,N_17997);
nand U18283 (N_18283,N_17558,N_17954);
or U18284 (N_18284,N_17519,N_17722);
or U18285 (N_18285,N_17643,N_17684);
nor U18286 (N_18286,N_17603,N_17739);
nor U18287 (N_18287,N_17793,N_17735);
and U18288 (N_18288,N_17970,N_17546);
and U18289 (N_18289,N_17800,N_17797);
and U18290 (N_18290,N_17730,N_17791);
or U18291 (N_18291,N_17711,N_17559);
or U18292 (N_18292,N_17533,N_17649);
nor U18293 (N_18293,N_17898,N_17771);
and U18294 (N_18294,N_17966,N_17585);
or U18295 (N_18295,N_17647,N_17809);
nor U18296 (N_18296,N_17542,N_17887);
nor U18297 (N_18297,N_17877,N_17556);
nor U18298 (N_18298,N_17849,N_17662);
nand U18299 (N_18299,N_17981,N_17842);
or U18300 (N_18300,N_17710,N_17928);
nor U18301 (N_18301,N_17834,N_17982);
nand U18302 (N_18302,N_17537,N_17980);
nand U18303 (N_18303,N_17926,N_17800);
nand U18304 (N_18304,N_17584,N_17825);
or U18305 (N_18305,N_17763,N_17742);
and U18306 (N_18306,N_17772,N_17639);
or U18307 (N_18307,N_17628,N_17913);
or U18308 (N_18308,N_17747,N_17630);
xnor U18309 (N_18309,N_17668,N_17993);
nand U18310 (N_18310,N_17607,N_17929);
nor U18311 (N_18311,N_17541,N_17540);
and U18312 (N_18312,N_17593,N_17814);
nand U18313 (N_18313,N_17920,N_17615);
nor U18314 (N_18314,N_17536,N_17655);
nand U18315 (N_18315,N_17640,N_17749);
or U18316 (N_18316,N_17944,N_17780);
nor U18317 (N_18317,N_17676,N_17892);
nor U18318 (N_18318,N_17905,N_17861);
nor U18319 (N_18319,N_17721,N_17884);
nand U18320 (N_18320,N_17538,N_17531);
xnor U18321 (N_18321,N_17901,N_17995);
nor U18322 (N_18322,N_17520,N_17531);
or U18323 (N_18323,N_17639,N_17983);
nand U18324 (N_18324,N_17822,N_17938);
nand U18325 (N_18325,N_17550,N_17561);
nand U18326 (N_18326,N_17717,N_17895);
and U18327 (N_18327,N_17826,N_17817);
xor U18328 (N_18328,N_17628,N_17655);
nor U18329 (N_18329,N_17803,N_17873);
and U18330 (N_18330,N_17877,N_17943);
nor U18331 (N_18331,N_17811,N_17893);
xnor U18332 (N_18332,N_17579,N_17746);
xnor U18333 (N_18333,N_17805,N_17848);
xnor U18334 (N_18334,N_17776,N_17705);
xnor U18335 (N_18335,N_17889,N_17816);
or U18336 (N_18336,N_17512,N_17893);
nor U18337 (N_18337,N_17595,N_17807);
nand U18338 (N_18338,N_17565,N_17887);
nand U18339 (N_18339,N_17742,N_17687);
nand U18340 (N_18340,N_17664,N_17524);
nor U18341 (N_18341,N_17997,N_17936);
and U18342 (N_18342,N_17940,N_17724);
nor U18343 (N_18343,N_17990,N_17597);
nand U18344 (N_18344,N_17525,N_17642);
nand U18345 (N_18345,N_17534,N_17516);
xnor U18346 (N_18346,N_17751,N_17678);
nor U18347 (N_18347,N_17678,N_17740);
nor U18348 (N_18348,N_17739,N_17525);
and U18349 (N_18349,N_17880,N_17691);
nor U18350 (N_18350,N_17692,N_17841);
and U18351 (N_18351,N_17932,N_17909);
or U18352 (N_18352,N_17736,N_17888);
nor U18353 (N_18353,N_17642,N_17879);
nand U18354 (N_18354,N_17530,N_17993);
nand U18355 (N_18355,N_17816,N_17743);
xnor U18356 (N_18356,N_17912,N_17951);
xor U18357 (N_18357,N_17748,N_17707);
nor U18358 (N_18358,N_17700,N_17883);
xnor U18359 (N_18359,N_17862,N_17721);
and U18360 (N_18360,N_17858,N_17925);
nor U18361 (N_18361,N_17708,N_17795);
xnor U18362 (N_18362,N_17863,N_17564);
or U18363 (N_18363,N_17868,N_17762);
and U18364 (N_18364,N_17883,N_17859);
xor U18365 (N_18365,N_17752,N_17627);
or U18366 (N_18366,N_17574,N_17929);
or U18367 (N_18367,N_17888,N_17892);
and U18368 (N_18368,N_17754,N_17753);
xor U18369 (N_18369,N_17868,N_17797);
and U18370 (N_18370,N_17988,N_17612);
or U18371 (N_18371,N_17533,N_17879);
nor U18372 (N_18372,N_17589,N_17949);
or U18373 (N_18373,N_17779,N_17683);
and U18374 (N_18374,N_17996,N_17621);
nand U18375 (N_18375,N_17796,N_17747);
xnor U18376 (N_18376,N_17519,N_17620);
nor U18377 (N_18377,N_17993,N_17688);
nand U18378 (N_18378,N_17619,N_17548);
or U18379 (N_18379,N_17732,N_17513);
nor U18380 (N_18380,N_17644,N_17580);
xnor U18381 (N_18381,N_17852,N_17577);
xnor U18382 (N_18382,N_17866,N_17775);
or U18383 (N_18383,N_17583,N_17746);
or U18384 (N_18384,N_17580,N_17837);
nand U18385 (N_18385,N_17695,N_17507);
and U18386 (N_18386,N_17913,N_17649);
xnor U18387 (N_18387,N_17558,N_17526);
xor U18388 (N_18388,N_17982,N_17616);
xnor U18389 (N_18389,N_17505,N_17979);
nand U18390 (N_18390,N_17534,N_17527);
and U18391 (N_18391,N_17818,N_17667);
nor U18392 (N_18392,N_17698,N_17712);
and U18393 (N_18393,N_17959,N_17914);
or U18394 (N_18394,N_17561,N_17610);
nor U18395 (N_18395,N_17681,N_17776);
xnor U18396 (N_18396,N_17803,N_17791);
and U18397 (N_18397,N_17580,N_17801);
xor U18398 (N_18398,N_17643,N_17551);
or U18399 (N_18399,N_17858,N_17929);
nand U18400 (N_18400,N_17542,N_17879);
nand U18401 (N_18401,N_17536,N_17643);
xnor U18402 (N_18402,N_17587,N_17931);
or U18403 (N_18403,N_17732,N_17819);
and U18404 (N_18404,N_17667,N_17700);
nand U18405 (N_18405,N_17551,N_17882);
xnor U18406 (N_18406,N_17675,N_17921);
and U18407 (N_18407,N_17965,N_17919);
nand U18408 (N_18408,N_17558,N_17793);
and U18409 (N_18409,N_17649,N_17773);
and U18410 (N_18410,N_17692,N_17540);
nand U18411 (N_18411,N_17547,N_17728);
and U18412 (N_18412,N_17988,N_17775);
xnor U18413 (N_18413,N_17904,N_17891);
or U18414 (N_18414,N_17814,N_17808);
or U18415 (N_18415,N_17821,N_17886);
nor U18416 (N_18416,N_17782,N_17892);
xnor U18417 (N_18417,N_17752,N_17906);
nor U18418 (N_18418,N_17969,N_17930);
and U18419 (N_18419,N_17674,N_17954);
nor U18420 (N_18420,N_17596,N_17561);
nor U18421 (N_18421,N_17749,N_17527);
and U18422 (N_18422,N_17978,N_17798);
and U18423 (N_18423,N_17869,N_17940);
nand U18424 (N_18424,N_17701,N_17530);
and U18425 (N_18425,N_17648,N_17554);
nor U18426 (N_18426,N_17551,N_17860);
or U18427 (N_18427,N_17720,N_17997);
xor U18428 (N_18428,N_17623,N_17850);
and U18429 (N_18429,N_17521,N_17913);
xor U18430 (N_18430,N_17801,N_17852);
and U18431 (N_18431,N_17722,N_17983);
xor U18432 (N_18432,N_17856,N_17848);
or U18433 (N_18433,N_17934,N_17652);
and U18434 (N_18434,N_17789,N_17843);
nand U18435 (N_18435,N_17790,N_17848);
and U18436 (N_18436,N_17810,N_17979);
xor U18437 (N_18437,N_17581,N_17529);
and U18438 (N_18438,N_17827,N_17617);
or U18439 (N_18439,N_17951,N_17560);
or U18440 (N_18440,N_17804,N_17773);
or U18441 (N_18441,N_17713,N_17995);
nor U18442 (N_18442,N_17916,N_17976);
and U18443 (N_18443,N_17872,N_17934);
nor U18444 (N_18444,N_17888,N_17697);
or U18445 (N_18445,N_17595,N_17679);
or U18446 (N_18446,N_17782,N_17623);
or U18447 (N_18447,N_17639,N_17987);
xor U18448 (N_18448,N_17762,N_17808);
nor U18449 (N_18449,N_17970,N_17699);
nand U18450 (N_18450,N_17805,N_17649);
nor U18451 (N_18451,N_17593,N_17935);
or U18452 (N_18452,N_17579,N_17747);
or U18453 (N_18453,N_17662,N_17679);
nor U18454 (N_18454,N_17721,N_17612);
xnor U18455 (N_18455,N_17856,N_17835);
and U18456 (N_18456,N_17563,N_17851);
nor U18457 (N_18457,N_17618,N_17742);
and U18458 (N_18458,N_17967,N_17773);
or U18459 (N_18459,N_17853,N_17886);
or U18460 (N_18460,N_17672,N_17873);
nand U18461 (N_18461,N_17845,N_17980);
or U18462 (N_18462,N_17778,N_17576);
nor U18463 (N_18463,N_17865,N_17694);
nor U18464 (N_18464,N_17965,N_17656);
or U18465 (N_18465,N_17779,N_17893);
nor U18466 (N_18466,N_17641,N_17865);
nand U18467 (N_18467,N_17995,N_17906);
nor U18468 (N_18468,N_17964,N_17732);
nand U18469 (N_18469,N_17632,N_17969);
nor U18470 (N_18470,N_17970,N_17737);
nor U18471 (N_18471,N_17933,N_17615);
or U18472 (N_18472,N_17815,N_17754);
and U18473 (N_18473,N_17716,N_17507);
nor U18474 (N_18474,N_17971,N_17891);
xor U18475 (N_18475,N_17835,N_17766);
or U18476 (N_18476,N_17563,N_17737);
nand U18477 (N_18477,N_17596,N_17840);
and U18478 (N_18478,N_17823,N_17612);
or U18479 (N_18479,N_17694,N_17758);
nor U18480 (N_18480,N_17655,N_17695);
nand U18481 (N_18481,N_17623,N_17764);
nor U18482 (N_18482,N_17727,N_17852);
or U18483 (N_18483,N_17974,N_17927);
and U18484 (N_18484,N_17691,N_17593);
xor U18485 (N_18485,N_17633,N_17941);
and U18486 (N_18486,N_17500,N_17538);
nor U18487 (N_18487,N_17779,N_17877);
and U18488 (N_18488,N_17996,N_17955);
and U18489 (N_18489,N_17505,N_17617);
or U18490 (N_18490,N_17906,N_17938);
or U18491 (N_18491,N_17527,N_17883);
nand U18492 (N_18492,N_17768,N_17757);
and U18493 (N_18493,N_17727,N_17590);
nor U18494 (N_18494,N_17525,N_17544);
xnor U18495 (N_18495,N_17973,N_17809);
nor U18496 (N_18496,N_17843,N_17551);
nor U18497 (N_18497,N_17588,N_17558);
and U18498 (N_18498,N_17512,N_17859);
nand U18499 (N_18499,N_17580,N_17951);
or U18500 (N_18500,N_18346,N_18002);
and U18501 (N_18501,N_18100,N_18304);
and U18502 (N_18502,N_18081,N_18490);
xor U18503 (N_18503,N_18413,N_18156);
xor U18504 (N_18504,N_18141,N_18083);
or U18505 (N_18505,N_18395,N_18223);
nor U18506 (N_18506,N_18211,N_18308);
or U18507 (N_18507,N_18046,N_18466);
and U18508 (N_18508,N_18322,N_18228);
nor U18509 (N_18509,N_18377,N_18199);
or U18510 (N_18510,N_18414,N_18102);
and U18511 (N_18511,N_18142,N_18289);
or U18512 (N_18512,N_18122,N_18494);
nor U18513 (N_18513,N_18471,N_18441);
or U18514 (N_18514,N_18014,N_18135);
xnor U18515 (N_18515,N_18019,N_18138);
nor U18516 (N_18516,N_18434,N_18110);
xnor U18517 (N_18517,N_18012,N_18220);
nand U18518 (N_18518,N_18437,N_18341);
nor U18519 (N_18519,N_18253,N_18123);
nor U18520 (N_18520,N_18154,N_18003);
or U18521 (N_18521,N_18037,N_18005);
xnor U18522 (N_18522,N_18387,N_18070);
nand U18523 (N_18523,N_18239,N_18309);
and U18524 (N_18524,N_18167,N_18314);
nor U18525 (N_18525,N_18112,N_18354);
or U18526 (N_18526,N_18485,N_18139);
nand U18527 (N_18527,N_18349,N_18311);
xor U18528 (N_18528,N_18101,N_18085);
nor U18529 (N_18529,N_18491,N_18440);
and U18530 (N_18530,N_18399,N_18376);
and U18531 (N_18531,N_18040,N_18062);
xnor U18532 (N_18532,N_18416,N_18043);
and U18533 (N_18533,N_18408,N_18275);
xor U18534 (N_18534,N_18236,N_18451);
or U18535 (N_18535,N_18010,N_18045);
or U18536 (N_18536,N_18000,N_18237);
nand U18537 (N_18537,N_18233,N_18450);
nor U18538 (N_18538,N_18247,N_18128);
or U18539 (N_18539,N_18463,N_18018);
nor U18540 (N_18540,N_18210,N_18096);
and U18541 (N_18541,N_18386,N_18303);
nor U18542 (N_18542,N_18295,N_18205);
nand U18543 (N_18543,N_18367,N_18280);
nand U18544 (N_18544,N_18151,N_18079);
or U18545 (N_18545,N_18121,N_18360);
nand U18546 (N_18546,N_18125,N_18161);
and U18547 (N_18547,N_18366,N_18137);
and U18548 (N_18548,N_18011,N_18484);
nor U18549 (N_18549,N_18186,N_18301);
nand U18550 (N_18550,N_18152,N_18075);
nand U18551 (N_18551,N_18460,N_18179);
xor U18552 (N_18552,N_18472,N_18224);
nand U18553 (N_18553,N_18458,N_18444);
nor U18554 (N_18554,N_18283,N_18453);
nand U18555 (N_18555,N_18098,N_18315);
nor U18556 (N_18556,N_18063,N_18007);
xor U18557 (N_18557,N_18483,N_18392);
or U18558 (N_18558,N_18194,N_18113);
xnor U18559 (N_18559,N_18164,N_18323);
or U18560 (N_18560,N_18058,N_18118);
and U18561 (N_18561,N_18073,N_18061);
nor U18562 (N_18562,N_18254,N_18184);
nor U18563 (N_18563,N_18475,N_18391);
nand U18564 (N_18564,N_18221,N_18343);
or U18565 (N_18565,N_18262,N_18251);
and U18566 (N_18566,N_18325,N_18390);
nand U18567 (N_18567,N_18190,N_18207);
xnor U18568 (N_18568,N_18340,N_18243);
xor U18569 (N_18569,N_18449,N_18134);
and U18570 (N_18570,N_18189,N_18363);
and U18571 (N_18571,N_18024,N_18107);
xnor U18572 (N_18572,N_18424,N_18488);
or U18573 (N_18573,N_18278,N_18284);
and U18574 (N_18574,N_18307,N_18042);
and U18575 (N_18575,N_18027,N_18088);
and U18576 (N_18576,N_18418,N_18092);
xor U18577 (N_18577,N_18317,N_18039);
nor U18578 (N_18578,N_18192,N_18328);
nand U18579 (N_18579,N_18294,N_18389);
xnor U18580 (N_18580,N_18109,N_18162);
nor U18581 (N_18581,N_18230,N_18191);
or U18582 (N_18582,N_18312,N_18299);
xnor U18583 (N_18583,N_18267,N_18193);
xor U18584 (N_18584,N_18173,N_18182);
nand U18585 (N_18585,N_18359,N_18147);
nor U18586 (N_18586,N_18124,N_18271);
nor U18587 (N_18587,N_18131,N_18400);
nor U18588 (N_18588,N_18329,N_18248);
and U18589 (N_18589,N_18443,N_18175);
and U18590 (N_18590,N_18021,N_18293);
xor U18591 (N_18591,N_18302,N_18324);
nor U18592 (N_18592,N_18215,N_18263);
xnor U18593 (N_18593,N_18461,N_18266);
or U18594 (N_18594,N_18047,N_18404);
nand U18595 (N_18595,N_18127,N_18196);
and U18596 (N_18596,N_18214,N_18393);
or U18597 (N_18597,N_18222,N_18105);
nand U18598 (N_18598,N_18455,N_18212);
nand U18599 (N_18599,N_18203,N_18375);
nand U18600 (N_18600,N_18022,N_18041);
or U18601 (N_18601,N_18495,N_18468);
and U18602 (N_18602,N_18177,N_18069);
nand U18603 (N_18603,N_18218,N_18352);
nand U18604 (N_18604,N_18286,N_18067);
and U18605 (N_18605,N_18421,N_18195);
nor U18606 (N_18606,N_18038,N_18496);
or U18607 (N_18607,N_18094,N_18478);
or U18608 (N_18608,N_18025,N_18185);
and U18609 (N_18609,N_18180,N_18499);
or U18610 (N_18610,N_18227,N_18029);
and U18611 (N_18611,N_18355,N_18273);
xnor U18612 (N_18612,N_18330,N_18270);
xnor U18613 (N_18613,N_18454,N_18462);
or U18614 (N_18614,N_18445,N_18261);
and U18615 (N_18615,N_18398,N_18287);
nand U18616 (N_18616,N_18351,N_18467);
or U18617 (N_18617,N_18357,N_18257);
or U18618 (N_18618,N_18272,N_18411);
nand U18619 (N_18619,N_18310,N_18479);
nand U18620 (N_18620,N_18292,N_18417);
nand U18621 (N_18621,N_18091,N_18335);
and U18622 (N_18622,N_18422,N_18498);
or U18623 (N_18623,N_18300,N_18204);
nand U18624 (N_18624,N_18093,N_18115);
xnor U18625 (N_18625,N_18208,N_18406);
and U18626 (N_18626,N_18313,N_18249);
xor U18627 (N_18627,N_18350,N_18155);
xnor U18628 (N_18628,N_18241,N_18446);
xnor U18629 (N_18629,N_18049,N_18333);
nand U18630 (N_18630,N_18338,N_18051);
nand U18631 (N_18631,N_18053,N_18345);
and U18632 (N_18632,N_18415,N_18469);
or U18633 (N_18633,N_18183,N_18246);
or U18634 (N_18634,N_18370,N_18200);
or U18635 (N_18635,N_18332,N_18030);
nor U18636 (N_18636,N_18371,N_18419);
xor U18637 (N_18637,N_18126,N_18274);
xnor U18638 (N_18638,N_18265,N_18015);
nor U18639 (N_18639,N_18380,N_18202);
nand U18640 (N_18640,N_18448,N_18114);
nor U18641 (N_18641,N_18432,N_18068);
or U18642 (N_18642,N_18382,N_18379);
xor U18643 (N_18643,N_18285,N_18384);
or U18644 (N_18644,N_18482,N_18425);
nand U18645 (N_18645,N_18004,N_18321);
or U18646 (N_18646,N_18009,N_18396);
nand U18647 (N_18647,N_18433,N_18059);
nor U18648 (N_18648,N_18362,N_18470);
nand U18649 (N_18649,N_18402,N_18136);
or U18650 (N_18650,N_18072,N_18225);
nor U18651 (N_18651,N_18166,N_18158);
xnor U18652 (N_18652,N_18447,N_18279);
nand U18653 (N_18653,N_18157,N_18240);
nor U18654 (N_18654,N_18170,N_18439);
nand U18655 (N_18655,N_18242,N_18116);
xnor U18656 (N_18656,N_18486,N_18296);
or U18657 (N_18657,N_18008,N_18264);
nor U18658 (N_18658,N_18089,N_18487);
nor U18659 (N_18659,N_18132,N_18111);
nand U18660 (N_18660,N_18474,N_18036);
nor U18661 (N_18661,N_18130,N_18250);
nand U18662 (N_18662,N_18492,N_18368);
nand U18663 (N_18663,N_18056,N_18169);
nand U18664 (N_18664,N_18378,N_18097);
nor U18665 (N_18665,N_18168,N_18410);
nor U18666 (N_18666,N_18181,N_18099);
or U18667 (N_18667,N_18347,N_18342);
and U18668 (N_18668,N_18409,N_18106);
xnor U18669 (N_18669,N_18117,N_18327);
xnor U18670 (N_18670,N_18493,N_18054);
xor U18671 (N_18671,N_18305,N_18457);
nor U18672 (N_18672,N_18477,N_18397);
and U18673 (N_18673,N_18219,N_18129);
xnor U18674 (N_18674,N_18148,N_18133);
xor U18675 (N_18675,N_18201,N_18436);
nor U18676 (N_18676,N_18172,N_18381);
nor U18677 (N_18677,N_18035,N_18140);
or U18678 (N_18678,N_18481,N_18291);
nor U18679 (N_18679,N_18369,N_18331);
nand U18680 (N_18680,N_18497,N_18055);
or U18681 (N_18681,N_18276,N_18020);
or U18682 (N_18682,N_18339,N_18216);
xnor U18683 (N_18683,N_18071,N_18316);
nor U18684 (N_18684,N_18174,N_18160);
nor U18685 (N_18685,N_18420,N_18234);
nor U18686 (N_18686,N_18337,N_18050);
nand U18687 (N_18687,N_18412,N_18013);
xnor U18688 (N_18688,N_18277,N_18064);
nand U18689 (N_18689,N_18052,N_18429);
nor U18690 (N_18690,N_18016,N_18066);
and U18691 (N_18691,N_18076,N_18489);
nor U18692 (N_18692,N_18426,N_18260);
nand U18693 (N_18693,N_18394,N_18385);
nor U18694 (N_18694,N_18464,N_18153);
nor U18695 (N_18695,N_18281,N_18336);
nand U18696 (N_18696,N_18244,N_18374);
or U18697 (N_18697,N_18465,N_18229);
or U18698 (N_18698,N_18372,N_18306);
or U18699 (N_18699,N_18213,N_18407);
nor U18700 (N_18700,N_18187,N_18198);
and U18701 (N_18701,N_18034,N_18258);
nand U18702 (N_18702,N_18226,N_18048);
nand U18703 (N_18703,N_18057,N_18269);
nand U18704 (N_18704,N_18430,N_18320);
and U18705 (N_18705,N_18023,N_18209);
xnor U18706 (N_18706,N_18074,N_18356);
nand U18707 (N_18707,N_18149,N_18238);
xnor U18708 (N_18708,N_18435,N_18032);
and U18709 (N_18709,N_18087,N_18006);
nand U18710 (N_18710,N_18290,N_18119);
nor U18711 (N_18711,N_18476,N_18188);
nand U18712 (N_18712,N_18388,N_18104);
nand U18713 (N_18713,N_18255,N_18031);
nand U18714 (N_18714,N_18318,N_18145);
and U18715 (N_18715,N_18176,N_18288);
nor U18716 (N_18716,N_18017,N_18428);
nor U18717 (N_18717,N_18232,N_18403);
and U18718 (N_18718,N_18282,N_18326);
nand U18719 (N_18719,N_18268,N_18473);
and U18720 (N_18720,N_18373,N_18365);
xnor U18721 (N_18721,N_18060,N_18082);
nand U18722 (N_18722,N_18144,N_18065);
nor U18723 (N_18723,N_18361,N_18197);
xor U18724 (N_18724,N_18344,N_18103);
nor U18725 (N_18725,N_18028,N_18150);
nand U18726 (N_18726,N_18143,N_18078);
or U18727 (N_18727,N_18401,N_18334);
xnor U18728 (N_18728,N_18358,N_18252);
or U18729 (N_18729,N_18298,N_18456);
nor U18730 (N_18730,N_18427,N_18001);
nand U18731 (N_18731,N_18026,N_18178);
nand U18732 (N_18732,N_18077,N_18319);
nor U18733 (N_18733,N_18090,N_18146);
or U18734 (N_18734,N_18245,N_18423);
or U18735 (N_18735,N_18442,N_18431);
xnor U18736 (N_18736,N_18480,N_18165);
nand U18737 (N_18737,N_18095,N_18383);
nor U18738 (N_18738,N_18459,N_18256);
xor U18739 (N_18739,N_18159,N_18084);
nor U18740 (N_18740,N_18452,N_18364);
nor U18741 (N_18741,N_18080,N_18044);
and U18742 (N_18742,N_18217,N_18438);
nand U18743 (N_18743,N_18033,N_18120);
and U18744 (N_18744,N_18405,N_18297);
or U18745 (N_18745,N_18348,N_18108);
nor U18746 (N_18746,N_18163,N_18259);
xnor U18747 (N_18747,N_18235,N_18206);
nor U18748 (N_18748,N_18171,N_18231);
and U18749 (N_18749,N_18353,N_18086);
or U18750 (N_18750,N_18231,N_18295);
xor U18751 (N_18751,N_18208,N_18160);
or U18752 (N_18752,N_18423,N_18188);
or U18753 (N_18753,N_18456,N_18130);
nand U18754 (N_18754,N_18446,N_18123);
xor U18755 (N_18755,N_18080,N_18256);
nand U18756 (N_18756,N_18112,N_18477);
and U18757 (N_18757,N_18447,N_18375);
nor U18758 (N_18758,N_18176,N_18410);
and U18759 (N_18759,N_18218,N_18308);
or U18760 (N_18760,N_18196,N_18305);
and U18761 (N_18761,N_18178,N_18287);
and U18762 (N_18762,N_18433,N_18052);
or U18763 (N_18763,N_18203,N_18247);
nand U18764 (N_18764,N_18112,N_18445);
nor U18765 (N_18765,N_18007,N_18265);
xor U18766 (N_18766,N_18423,N_18401);
nand U18767 (N_18767,N_18200,N_18109);
or U18768 (N_18768,N_18434,N_18119);
xor U18769 (N_18769,N_18045,N_18180);
nor U18770 (N_18770,N_18263,N_18092);
xnor U18771 (N_18771,N_18156,N_18264);
nor U18772 (N_18772,N_18208,N_18148);
nor U18773 (N_18773,N_18059,N_18396);
or U18774 (N_18774,N_18125,N_18299);
and U18775 (N_18775,N_18103,N_18224);
xor U18776 (N_18776,N_18130,N_18379);
nand U18777 (N_18777,N_18213,N_18127);
xnor U18778 (N_18778,N_18071,N_18271);
xor U18779 (N_18779,N_18110,N_18263);
nor U18780 (N_18780,N_18030,N_18265);
and U18781 (N_18781,N_18299,N_18228);
xnor U18782 (N_18782,N_18116,N_18199);
and U18783 (N_18783,N_18383,N_18473);
or U18784 (N_18784,N_18236,N_18344);
or U18785 (N_18785,N_18227,N_18190);
or U18786 (N_18786,N_18470,N_18496);
and U18787 (N_18787,N_18433,N_18160);
nor U18788 (N_18788,N_18048,N_18213);
nor U18789 (N_18789,N_18312,N_18278);
nor U18790 (N_18790,N_18302,N_18223);
xor U18791 (N_18791,N_18173,N_18088);
nand U18792 (N_18792,N_18036,N_18019);
xor U18793 (N_18793,N_18067,N_18199);
nand U18794 (N_18794,N_18087,N_18194);
nor U18795 (N_18795,N_18468,N_18221);
and U18796 (N_18796,N_18257,N_18025);
or U18797 (N_18797,N_18198,N_18438);
nor U18798 (N_18798,N_18130,N_18118);
and U18799 (N_18799,N_18343,N_18099);
nand U18800 (N_18800,N_18015,N_18494);
and U18801 (N_18801,N_18482,N_18117);
and U18802 (N_18802,N_18379,N_18090);
nor U18803 (N_18803,N_18447,N_18402);
nand U18804 (N_18804,N_18051,N_18086);
nand U18805 (N_18805,N_18252,N_18189);
nand U18806 (N_18806,N_18023,N_18305);
xnor U18807 (N_18807,N_18307,N_18378);
xor U18808 (N_18808,N_18051,N_18251);
and U18809 (N_18809,N_18330,N_18360);
nor U18810 (N_18810,N_18239,N_18267);
nand U18811 (N_18811,N_18289,N_18296);
xor U18812 (N_18812,N_18411,N_18010);
nand U18813 (N_18813,N_18083,N_18243);
xor U18814 (N_18814,N_18342,N_18220);
and U18815 (N_18815,N_18280,N_18490);
and U18816 (N_18816,N_18023,N_18152);
and U18817 (N_18817,N_18289,N_18169);
nand U18818 (N_18818,N_18133,N_18481);
nor U18819 (N_18819,N_18040,N_18243);
nor U18820 (N_18820,N_18051,N_18096);
or U18821 (N_18821,N_18141,N_18454);
or U18822 (N_18822,N_18202,N_18011);
xnor U18823 (N_18823,N_18109,N_18327);
nand U18824 (N_18824,N_18123,N_18318);
nand U18825 (N_18825,N_18219,N_18326);
or U18826 (N_18826,N_18415,N_18130);
nand U18827 (N_18827,N_18126,N_18110);
or U18828 (N_18828,N_18056,N_18097);
xnor U18829 (N_18829,N_18388,N_18048);
and U18830 (N_18830,N_18362,N_18093);
and U18831 (N_18831,N_18360,N_18489);
nor U18832 (N_18832,N_18089,N_18458);
or U18833 (N_18833,N_18112,N_18141);
and U18834 (N_18834,N_18129,N_18302);
or U18835 (N_18835,N_18062,N_18199);
nor U18836 (N_18836,N_18052,N_18274);
nor U18837 (N_18837,N_18167,N_18032);
nand U18838 (N_18838,N_18489,N_18354);
nor U18839 (N_18839,N_18132,N_18428);
nor U18840 (N_18840,N_18398,N_18006);
nand U18841 (N_18841,N_18041,N_18285);
nand U18842 (N_18842,N_18380,N_18027);
nor U18843 (N_18843,N_18241,N_18432);
nor U18844 (N_18844,N_18135,N_18000);
and U18845 (N_18845,N_18052,N_18303);
nand U18846 (N_18846,N_18099,N_18471);
and U18847 (N_18847,N_18489,N_18383);
xnor U18848 (N_18848,N_18370,N_18256);
and U18849 (N_18849,N_18044,N_18348);
nor U18850 (N_18850,N_18347,N_18286);
and U18851 (N_18851,N_18279,N_18093);
or U18852 (N_18852,N_18201,N_18194);
nand U18853 (N_18853,N_18204,N_18063);
and U18854 (N_18854,N_18250,N_18040);
and U18855 (N_18855,N_18423,N_18139);
xor U18856 (N_18856,N_18217,N_18397);
and U18857 (N_18857,N_18261,N_18399);
or U18858 (N_18858,N_18479,N_18408);
xor U18859 (N_18859,N_18298,N_18280);
nand U18860 (N_18860,N_18275,N_18477);
and U18861 (N_18861,N_18263,N_18184);
nand U18862 (N_18862,N_18329,N_18018);
or U18863 (N_18863,N_18488,N_18164);
or U18864 (N_18864,N_18123,N_18457);
xnor U18865 (N_18865,N_18078,N_18233);
or U18866 (N_18866,N_18359,N_18407);
nand U18867 (N_18867,N_18398,N_18230);
xnor U18868 (N_18868,N_18046,N_18407);
and U18869 (N_18869,N_18395,N_18405);
or U18870 (N_18870,N_18250,N_18377);
nor U18871 (N_18871,N_18355,N_18196);
xnor U18872 (N_18872,N_18109,N_18271);
and U18873 (N_18873,N_18289,N_18476);
or U18874 (N_18874,N_18079,N_18417);
nand U18875 (N_18875,N_18004,N_18136);
nor U18876 (N_18876,N_18022,N_18138);
xnor U18877 (N_18877,N_18155,N_18395);
and U18878 (N_18878,N_18232,N_18171);
nor U18879 (N_18879,N_18138,N_18277);
xnor U18880 (N_18880,N_18077,N_18262);
nor U18881 (N_18881,N_18146,N_18460);
and U18882 (N_18882,N_18349,N_18060);
xnor U18883 (N_18883,N_18090,N_18383);
nand U18884 (N_18884,N_18471,N_18092);
nand U18885 (N_18885,N_18493,N_18006);
xor U18886 (N_18886,N_18113,N_18310);
or U18887 (N_18887,N_18306,N_18039);
nand U18888 (N_18888,N_18443,N_18049);
xor U18889 (N_18889,N_18327,N_18447);
xnor U18890 (N_18890,N_18298,N_18442);
nor U18891 (N_18891,N_18461,N_18301);
or U18892 (N_18892,N_18138,N_18468);
or U18893 (N_18893,N_18095,N_18069);
and U18894 (N_18894,N_18028,N_18421);
or U18895 (N_18895,N_18085,N_18204);
nand U18896 (N_18896,N_18451,N_18040);
nor U18897 (N_18897,N_18287,N_18461);
and U18898 (N_18898,N_18288,N_18106);
xor U18899 (N_18899,N_18453,N_18480);
or U18900 (N_18900,N_18285,N_18261);
and U18901 (N_18901,N_18232,N_18043);
and U18902 (N_18902,N_18319,N_18472);
nor U18903 (N_18903,N_18137,N_18271);
xnor U18904 (N_18904,N_18337,N_18307);
or U18905 (N_18905,N_18019,N_18107);
xor U18906 (N_18906,N_18072,N_18098);
and U18907 (N_18907,N_18001,N_18012);
nor U18908 (N_18908,N_18253,N_18024);
nand U18909 (N_18909,N_18120,N_18434);
xnor U18910 (N_18910,N_18199,N_18444);
nand U18911 (N_18911,N_18165,N_18393);
xnor U18912 (N_18912,N_18427,N_18264);
nand U18913 (N_18913,N_18367,N_18380);
nor U18914 (N_18914,N_18229,N_18475);
and U18915 (N_18915,N_18068,N_18462);
and U18916 (N_18916,N_18075,N_18037);
xor U18917 (N_18917,N_18356,N_18143);
and U18918 (N_18918,N_18421,N_18003);
and U18919 (N_18919,N_18221,N_18238);
xor U18920 (N_18920,N_18357,N_18416);
nand U18921 (N_18921,N_18105,N_18390);
and U18922 (N_18922,N_18482,N_18484);
xor U18923 (N_18923,N_18431,N_18358);
and U18924 (N_18924,N_18415,N_18461);
nand U18925 (N_18925,N_18422,N_18400);
or U18926 (N_18926,N_18481,N_18175);
nand U18927 (N_18927,N_18301,N_18419);
nand U18928 (N_18928,N_18130,N_18255);
xnor U18929 (N_18929,N_18352,N_18390);
xnor U18930 (N_18930,N_18044,N_18160);
or U18931 (N_18931,N_18348,N_18041);
or U18932 (N_18932,N_18116,N_18405);
and U18933 (N_18933,N_18274,N_18488);
nand U18934 (N_18934,N_18390,N_18379);
xor U18935 (N_18935,N_18495,N_18029);
xor U18936 (N_18936,N_18355,N_18311);
nor U18937 (N_18937,N_18064,N_18271);
and U18938 (N_18938,N_18284,N_18334);
nor U18939 (N_18939,N_18310,N_18251);
nor U18940 (N_18940,N_18272,N_18300);
xor U18941 (N_18941,N_18019,N_18055);
xnor U18942 (N_18942,N_18256,N_18212);
xnor U18943 (N_18943,N_18370,N_18248);
and U18944 (N_18944,N_18179,N_18008);
and U18945 (N_18945,N_18212,N_18017);
and U18946 (N_18946,N_18475,N_18128);
or U18947 (N_18947,N_18247,N_18166);
or U18948 (N_18948,N_18351,N_18083);
and U18949 (N_18949,N_18349,N_18459);
or U18950 (N_18950,N_18059,N_18000);
nor U18951 (N_18951,N_18429,N_18131);
nor U18952 (N_18952,N_18497,N_18256);
and U18953 (N_18953,N_18313,N_18180);
and U18954 (N_18954,N_18413,N_18112);
xor U18955 (N_18955,N_18342,N_18423);
xnor U18956 (N_18956,N_18470,N_18042);
xnor U18957 (N_18957,N_18463,N_18192);
nand U18958 (N_18958,N_18196,N_18403);
nor U18959 (N_18959,N_18247,N_18021);
xnor U18960 (N_18960,N_18427,N_18215);
nor U18961 (N_18961,N_18015,N_18114);
nor U18962 (N_18962,N_18396,N_18474);
and U18963 (N_18963,N_18282,N_18352);
nand U18964 (N_18964,N_18075,N_18196);
xnor U18965 (N_18965,N_18420,N_18276);
nor U18966 (N_18966,N_18216,N_18002);
nor U18967 (N_18967,N_18264,N_18472);
and U18968 (N_18968,N_18040,N_18293);
nand U18969 (N_18969,N_18148,N_18248);
nor U18970 (N_18970,N_18497,N_18271);
nor U18971 (N_18971,N_18272,N_18401);
xor U18972 (N_18972,N_18083,N_18457);
nand U18973 (N_18973,N_18248,N_18084);
or U18974 (N_18974,N_18395,N_18118);
and U18975 (N_18975,N_18470,N_18045);
and U18976 (N_18976,N_18456,N_18372);
and U18977 (N_18977,N_18217,N_18203);
nor U18978 (N_18978,N_18270,N_18391);
or U18979 (N_18979,N_18180,N_18009);
or U18980 (N_18980,N_18482,N_18219);
xor U18981 (N_18981,N_18091,N_18470);
nor U18982 (N_18982,N_18356,N_18366);
or U18983 (N_18983,N_18407,N_18189);
and U18984 (N_18984,N_18493,N_18178);
and U18985 (N_18985,N_18117,N_18020);
nor U18986 (N_18986,N_18390,N_18269);
nand U18987 (N_18987,N_18489,N_18338);
xor U18988 (N_18988,N_18417,N_18247);
or U18989 (N_18989,N_18331,N_18257);
and U18990 (N_18990,N_18004,N_18043);
xnor U18991 (N_18991,N_18148,N_18221);
and U18992 (N_18992,N_18290,N_18053);
nand U18993 (N_18993,N_18255,N_18452);
xor U18994 (N_18994,N_18262,N_18379);
and U18995 (N_18995,N_18097,N_18295);
xor U18996 (N_18996,N_18298,N_18231);
nand U18997 (N_18997,N_18124,N_18012);
or U18998 (N_18998,N_18138,N_18107);
nor U18999 (N_18999,N_18261,N_18463);
nor U19000 (N_19000,N_18903,N_18756);
xnor U19001 (N_19001,N_18672,N_18849);
or U19002 (N_19002,N_18997,N_18717);
nand U19003 (N_19003,N_18932,N_18562);
or U19004 (N_19004,N_18658,N_18784);
and U19005 (N_19005,N_18924,N_18986);
and U19006 (N_19006,N_18919,N_18881);
or U19007 (N_19007,N_18801,N_18628);
xnor U19008 (N_19008,N_18750,N_18871);
nand U19009 (N_19009,N_18963,N_18645);
or U19010 (N_19010,N_18720,N_18923);
xnor U19011 (N_19011,N_18882,N_18981);
xor U19012 (N_19012,N_18696,N_18677);
or U19013 (N_19013,N_18839,N_18859);
nand U19014 (N_19014,N_18836,N_18506);
and U19015 (N_19015,N_18889,N_18681);
xnor U19016 (N_19016,N_18691,N_18770);
nand U19017 (N_19017,N_18892,N_18771);
xor U19018 (N_19018,N_18548,N_18979);
nor U19019 (N_19019,N_18813,N_18917);
xor U19020 (N_19020,N_18608,N_18824);
nand U19021 (N_19021,N_18965,N_18577);
nor U19022 (N_19022,N_18583,N_18764);
nand U19023 (N_19023,N_18805,N_18897);
nor U19024 (N_19024,N_18906,N_18678);
or U19025 (N_19025,N_18729,N_18576);
or U19026 (N_19026,N_18854,N_18957);
xor U19027 (N_19027,N_18879,N_18954);
or U19028 (N_19028,N_18534,N_18961);
nor U19029 (N_19029,N_18683,N_18547);
nor U19030 (N_19030,N_18621,N_18984);
and U19031 (N_19031,N_18802,N_18690);
nor U19032 (N_19032,N_18996,N_18823);
and U19033 (N_19033,N_18557,N_18600);
xor U19034 (N_19034,N_18969,N_18694);
xnor U19035 (N_19035,N_18828,N_18816);
xnor U19036 (N_19036,N_18826,N_18657);
or U19037 (N_19037,N_18772,N_18795);
nor U19038 (N_19038,N_18604,N_18992);
and U19039 (N_19039,N_18833,N_18565);
nor U19040 (N_19040,N_18766,N_18762);
nand U19041 (N_19041,N_18514,N_18601);
nor U19042 (N_19042,N_18944,N_18737);
nand U19043 (N_19043,N_18618,N_18531);
xnor U19044 (N_19044,N_18679,N_18974);
or U19045 (N_19045,N_18735,N_18743);
nand U19046 (N_19046,N_18778,N_18680);
nand U19047 (N_19047,N_18977,N_18807);
or U19048 (N_19048,N_18960,N_18635);
nand U19049 (N_19049,N_18931,N_18788);
xor U19050 (N_19050,N_18858,N_18752);
nand U19051 (N_19051,N_18783,N_18905);
nand U19052 (N_19052,N_18662,N_18912);
and U19053 (N_19053,N_18508,N_18629);
nor U19054 (N_19054,N_18742,N_18939);
nand U19055 (N_19055,N_18509,N_18860);
or U19056 (N_19056,N_18806,N_18605);
nor U19057 (N_19057,N_18649,N_18718);
nor U19058 (N_19058,N_18582,N_18883);
and U19059 (N_19059,N_18949,N_18782);
nor U19060 (N_19060,N_18935,N_18799);
nand U19061 (N_19061,N_18885,N_18727);
or U19062 (N_19062,N_18513,N_18651);
or U19063 (N_19063,N_18950,N_18921);
nand U19064 (N_19064,N_18886,N_18511);
nor U19065 (N_19065,N_18934,N_18789);
or U19066 (N_19066,N_18744,N_18791);
xnor U19067 (N_19067,N_18962,N_18653);
and U19068 (N_19068,N_18559,N_18875);
xnor U19069 (N_19069,N_18704,N_18722);
nand U19070 (N_19070,N_18644,N_18627);
nand U19071 (N_19071,N_18941,N_18692);
xor U19072 (N_19072,N_18884,N_18516);
xor U19073 (N_19073,N_18529,N_18817);
or U19074 (N_19074,N_18993,N_18759);
xor U19075 (N_19075,N_18790,N_18555);
and U19076 (N_19076,N_18779,N_18517);
nor U19077 (N_19077,N_18834,N_18560);
xor U19078 (N_19078,N_18733,N_18995);
nor U19079 (N_19079,N_18872,N_18773);
and U19080 (N_19080,N_18646,N_18535);
nand U19081 (N_19081,N_18522,N_18573);
xnor U19082 (N_19082,N_18953,N_18641);
nor U19083 (N_19083,N_18930,N_18556);
nand U19084 (N_19084,N_18982,N_18874);
and U19085 (N_19085,N_18545,N_18687);
xor U19086 (N_19086,N_18580,N_18741);
nand U19087 (N_19087,N_18774,N_18617);
nor U19088 (N_19088,N_18537,N_18865);
nor U19089 (N_19089,N_18880,N_18708);
and U19090 (N_19090,N_18699,N_18916);
xor U19091 (N_19091,N_18714,N_18623);
or U19092 (N_19092,N_18948,N_18911);
nor U19093 (N_19093,N_18698,N_18847);
or U19094 (N_19094,N_18526,N_18561);
nand U19095 (N_19095,N_18611,N_18970);
or U19096 (N_19096,N_18734,N_18870);
xor U19097 (N_19097,N_18975,N_18814);
nor U19098 (N_19098,N_18850,N_18845);
nand U19099 (N_19099,N_18700,N_18838);
xor U19100 (N_19100,N_18887,N_18991);
or U19101 (N_19101,N_18607,N_18685);
nor U19102 (N_19102,N_18585,N_18819);
xnor U19103 (N_19103,N_18507,N_18825);
or U19104 (N_19104,N_18666,N_18612);
or U19105 (N_19105,N_18909,N_18890);
nand U19106 (N_19106,N_18758,N_18777);
nor U19107 (N_19107,N_18896,N_18837);
nand U19108 (N_19108,N_18978,N_18551);
or U19109 (N_19109,N_18829,N_18553);
xor U19110 (N_19110,N_18530,N_18877);
or U19111 (N_19111,N_18787,N_18863);
and U19112 (N_19112,N_18581,N_18810);
xnor U19113 (N_19113,N_18633,N_18940);
xor U19114 (N_19114,N_18913,N_18656);
nand U19115 (N_19115,N_18785,N_18546);
nand U19116 (N_19116,N_18637,N_18793);
xor U19117 (N_19117,N_18972,N_18908);
nand U19118 (N_19118,N_18732,N_18803);
or U19119 (N_19119,N_18579,N_18593);
nor U19120 (N_19120,N_18888,N_18663);
nand U19121 (N_19121,N_18693,N_18914);
nand U19122 (N_19122,N_18707,N_18634);
and U19123 (N_19123,N_18754,N_18808);
nand U19124 (N_19124,N_18609,N_18518);
nor U19125 (N_19125,N_18740,N_18625);
nor U19126 (N_19126,N_18552,N_18862);
nor U19127 (N_19127,N_18523,N_18521);
or U19128 (N_19128,N_18541,N_18985);
or U19129 (N_19129,N_18745,N_18739);
xnor U19130 (N_19130,N_18848,N_18959);
nand U19131 (N_19131,N_18857,N_18647);
nand U19132 (N_19132,N_18586,N_18851);
nor U19133 (N_19133,N_18780,N_18673);
and U19134 (N_19134,N_18809,N_18578);
or U19135 (N_19135,N_18763,N_18964);
nor U19136 (N_19136,N_18632,N_18724);
xnor U19137 (N_19137,N_18915,N_18792);
nor U19138 (N_19138,N_18544,N_18998);
nor U19139 (N_19139,N_18898,N_18500);
nand U19140 (N_19140,N_18602,N_18701);
xor U19141 (N_19141,N_18563,N_18542);
or U19142 (N_19142,N_18747,N_18527);
nor U19143 (N_19143,N_18661,N_18603);
nor U19144 (N_19144,N_18596,N_18775);
and U19145 (N_19145,N_18549,N_18706);
nand U19146 (N_19146,N_18515,N_18822);
and U19147 (N_19147,N_18512,N_18726);
nor U19148 (N_19148,N_18616,N_18613);
or U19149 (N_19149,N_18922,N_18861);
or U19150 (N_19150,N_18606,N_18564);
and U19151 (N_19151,N_18856,N_18648);
xnor U19152 (N_19152,N_18811,N_18804);
nand U19153 (N_19153,N_18505,N_18566);
or U19154 (N_19154,N_18827,N_18670);
xnor U19155 (N_19155,N_18768,N_18615);
and U19156 (N_19156,N_18894,N_18907);
nor U19157 (N_19157,N_18710,N_18660);
and U19158 (N_19158,N_18781,N_18504);
or U19159 (N_19159,N_18748,N_18840);
nand U19160 (N_19160,N_18574,N_18533);
nor U19161 (N_19161,N_18821,N_18757);
and U19162 (N_19162,N_18532,N_18818);
nand U19163 (N_19163,N_18925,N_18571);
and U19164 (N_19164,N_18835,N_18705);
nor U19165 (N_19165,N_18990,N_18971);
nand U19166 (N_19166,N_18667,N_18891);
nand U19167 (N_19167,N_18926,N_18719);
and U19168 (N_19168,N_18684,N_18502);
and U19169 (N_19169,N_18929,N_18587);
xor U19170 (N_19170,N_18820,N_18869);
xor U19171 (N_19171,N_18652,N_18753);
xnor U19172 (N_19172,N_18711,N_18540);
nor U19173 (N_19173,N_18844,N_18539);
and U19174 (N_19174,N_18760,N_18668);
nand U19175 (N_19175,N_18899,N_18968);
nor U19176 (N_19176,N_18832,N_18830);
nor U19177 (N_19177,N_18702,N_18873);
nor U19178 (N_19178,N_18584,N_18688);
nor U19179 (N_19179,N_18951,N_18731);
nand U19180 (N_19180,N_18642,N_18853);
and U19181 (N_19181,N_18864,N_18920);
or U19182 (N_19182,N_18786,N_18987);
and U19183 (N_19183,N_18958,N_18878);
xnor U19184 (N_19184,N_18855,N_18769);
or U19185 (N_19185,N_18842,N_18676);
or U19186 (N_19186,N_18592,N_18812);
nor U19187 (N_19187,N_18728,N_18746);
or U19188 (N_19188,N_18794,N_18945);
xnor U19189 (N_19189,N_18572,N_18619);
nand U19190 (N_19190,N_18638,N_18755);
nor U19191 (N_19191,N_18715,N_18665);
and U19192 (N_19192,N_18738,N_18598);
nor U19193 (N_19193,N_18868,N_18570);
or U19194 (N_19194,N_18943,N_18846);
or U19195 (N_19195,N_18620,N_18712);
nand U19196 (N_19196,N_18933,N_18866);
xnor U19197 (N_19197,N_18716,N_18674);
or U19198 (N_19198,N_18994,N_18636);
and U19199 (N_19199,N_18736,N_18988);
or U19200 (N_19200,N_18558,N_18852);
xnor U19201 (N_19201,N_18815,N_18761);
nand U19202 (N_19202,N_18893,N_18510);
or U19203 (N_19203,N_18589,N_18567);
nand U19204 (N_19204,N_18624,N_18900);
xor U19205 (N_19205,N_18622,N_18543);
or U19206 (N_19206,N_18639,N_18876);
and U19207 (N_19207,N_18765,N_18595);
nand U19208 (N_19208,N_18671,N_18501);
nand U19209 (N_19209,N_18675,N_18721);
or U19210 (N_19210,N_18631,N_18659);
nand U19211 (N_19211,N_18910,N_18682);
nor U19212 (N_19212,N_18928,N_18550);
and U19213 (N_19213,N_18640,N_18831);
xor U19214 (N_19214,N_18697,N_18655);
nor U19215 (N_19215,N_18695,N_18525);
nand U19216 (N_19216,N_18973,N_18536);
nand U19217 (N_19217,N_18937,N_18686);
nor U19218 (N_19218,N_18841,N_18524);
or U19219 (N_19219,N_18938,N_18796);
or U19220 (N_19220,N_18650,N_18843);
nand U19221 (N_19221,N_18703,N_18967);
xor U19222 (N_19222,N_18569,N_18751);
or U19223 (N_19223,N_18749,N_18901);
nand U19224 (N_19224,N_18904,N_18538);
xor U19225 (N_19225,N_18956,N_18946);
nor U19226 (N_19226,N_18800,N_18895);
xnor U19227 (N_19227,N_18723,N_18614);
or U19228 (N_19228,N_18713,N_18528);
or U19229 (N_19229,N_18730,N_18776);
nor U19230 (N_19230,N_18575,N_18626);
xor U19231 (N_19231,N_18709,N_18976);
xnor U19232 (N_19232,N_18610,N_18590);
or U19233 (N_19233,N_18725,N_18980);
and U19234 (N_19234,N_18902,N_18798);
or U19235 (N_19235,N_18983,N_18520);
nor U19236 (N_19236,N_18554,N_18599);
nand U19237 (N_19237,N_18568,N_18767);
nor U19238 (N_19238,N_18669,N_18630);
xnor U19239 (N_19239,N_18597,N_18643);
nor U19240 (N_19240,N_18918,N_18519);
and U19241 (N_19241,N_18594,N_18503);
nand U19242 (N_19242,N_18989,N_18867);
nand U19243 (N_19243,N_18952,N_18942);
and U19244 (N_19244,N_18936,N_18588);
or U19245 (N_19245,N_18797,N_18955);
or U19246 (N_19246,N_18966,N_18591);
or U19247 (N_19247,N_18654,N_18664);
xor U19248 (N_19248,N_18689,N_18947);
nand U19249 (N_19249,N_18999,N_18927);
and U19250 (N_19250,N_18873,N_18566);
nand U19251 (N_19251,N_18610,N_18669);
nand U19252 (N_19252,N_18637,N_18717);
and U19253 (N_19253,N_18599,N_18654);
nand U19254 (N_19254,N_18570,N_18648);
or U19255 (N_19255,N_18770,N_18612);
or U19256 (N_19256,N_18956,N_18858);
or U19257 (N_19257,N_18722,N_18849);
or U19258 (N_19258,N_18592,N_18751);
nand U19259 (N_19259,N_18723,N_18610);
or U19260 (N_19260,N_18589,N_18562);
or U19261 (N_19261,N_18754,N_18509);
or U19262 (N_19262,N_18845,N_18798);
nor U19263 (N_19263,N_18549,N_18613);
and U19264 (N_19264,N_18647,N_18601);
xor U19265 (N_19265,N_18784,N_18926);
nand U19266 (N_19266,N_18547,N_18749);
xor U19267 (N_19267,N_18765,N_18670);
nand U19268 (N_19268,N_18929,N_18950);
xnor U19269 (N_19269,N_18793,N_18853);
and U19270 (N_19270,N_18789,N_18990);
xnor U19271 (N_19271,N_18899,N_18984);
or U19272 (N_19272,N_18897,N_18750);
or U19273 (N_19273,N_18759,N_18959);
nand U19274 (N_19274,N_18949,N_18662);
nand U19275 (N_19275,N_18638,N_18725);
nand U19276 (N_19276,N_18736,N_18823);
nor U19277 (N_19277,N_18542,N_18527);
xnor U19278 (N_19278,N_18899,N_18831);
nor U19279 (N_19279,N_18698,N_18885);
or U19280 (N_19280,N_18862,N_18532);
nor U19281 (N_19281,N_18577,N_18532);
nand U19282 (N_19282,N_18977,N_18505);
and U19283 (N_19283,N_18789,N_18861);
nor U19284 (N_19284,N_18813,N_18831);
nand U19285 (N_19285,N_18881,N_18775);
and U19286 (N_19286,N_18523,N_18675);
nor U19287 (N_19287,N_18554,N_18729);
nor U19288 (N_19288,N_18976,N_18909);
or U19289 (N_19289,N_18506,N_18528);
nand U19290 (N_19290,N_18987,N_18608);
nor U19291 (N_19291,N_18906,N_18856);
xnor U19292 (N_19292,N_18553,N_18876);
xor U19293 (N_19293,N_18830,N_18553);
or U19294 (N_19294,N_18606,N_18586);
nor U19295 (N_19295,N_18930,N_18816);
nand U19296 (N_19296,N_18560,N_18931);
nor U19297 (N_19297,N_18928,N_18629);
xor U19298 (N_19298,N_18690,N_18667);
xor U19299 (N_19299,N_18948,N_18736);
xor U19300 (N_19300,N_18568,N_18617);
nor U19301 (N_19301,N_18529,N_18826);
and U19302 (N_19302,N_18745,N_18912);
xnor U19303 (N_19303,N_18643,N_18970);
nand U19304 (N_19304,N_18719,N_18559);
and U19305 (N_19305,N_18554,N_18818);
xor U19306 (N_19306,N_18854,N_18537);
nand U19307 (N_19307,N_18514,N_18736);
or U19308 (N_19308,N_18841,N_18987);
nor U19309 (N_19309,N_18899,N_18613);
nand U19310 (N_19310,N_18501,N_18532);
nand U19311 (N_19311,N_18561,N_18515);
xnor U19312 (N_19312,N_18913,N_18982);
nor U19313 (N_19313,N_18618,N_18979);
or U19314 (N_19314,N_18920,N_18544);
nand U19315 (N_19315,N_18560,N_18508);
xnor U19316 (N_19316,N_18724,N_18545);
or U19317 (N_19317,N_18627,N_18824);
and U19318 (N_19318,N_18666,N_18840);
xor U19319 (N_19319,N_18531,N_18711);
xor U19320 (N_19320,N_18822,N_18865);
and U19321 (N_19321,N_18657,N_18722);
nand U19322 (N_19322,N_18759,N_18659);
nor U19323 (N_19323,N_18947,N_18817);
or U19324 (N_19324,N_18956,N_18862);
xor U19325 (N_19325,N_18750,N_18779);
and U19326 (N_19326,N_18969,N_18659);
and U19327 (N_19327,N_18831,N_18865);
xnor U19328 (N_19328,N_18892,N_18989);
nand U19329 (N_19329,N_18958,N_18942);
xnor U19330 (N_19330,N_18654,N_18719);
nor U19331 (N_19331,N_18530,N_18776);
nor U19332 (N_19332,N_18900,N_18755);
or U19333 (N_19333,N_18732,N_18543);
xor U19334 (N_19334,N_18933,N_18808);
and U19335 (N_19335,N_18878,N_18537);
nand U19336 (N_19336,N_18854,N_18501);
nand U19337 (N_19337,N_18960,N_18934);
nand U19338 (N_19338,N_18819,N_18573);
nand U19339 (N_19339,N_18712,N_18846);
and U19340 (N_19340,N_18878,N_18894);
or U19341 (N_19341,N_18667,N_18651);
xor U19342 (N_19342,N_18837,N_18720);
and U19343 (N_19343,N_18737,N_18672);
or U19344 (N_19344,N_18504,N_18609);
nor U19345 (N_19345,N_18945,N_18849);
xor U19346 (N_19346,N_18523,N_18582);
nor U19347 (N_19347,N_18950,N_18941);
or U19348 (N_19348,N_18909,N_18510);
or U19349 (N_19349,N_18598,N_18939);
nor U19350 (N_19350,N_18783,N_18944);
nor U19351 (N_19351,N_18524,N_18902);
nor U19352 (N_19352,N_18506,N_18661);
xnor U19353 (N_19353,N_18731,N_18559);
and U19354 (N_19354,N_18595,N_18750);
nor U19355 (N_19355,N_18560,N_18782);
nand U19356 (N_19356,N_18505,N_18749);
or U19357 (N_19357,N_18816,N_18687);
and U19358 (N_19358,N_18984,N_18737);
nand U19359 (N_19359,N_18741,N_18507);
nor U19360 (N_19360,N_18923,N_18639);
xnor U19361 (N_19361,N_18580,N_18800);
and U19362 (N_19362,N_18610,N_18894);
xor U19363 (N_19363,N_18608,N_18661);
or U19364 (N_19364,N_18986,N_18693);
nand U19365 (N_19365,N_18834,N_18792);
nor U19366 (N_19366,N_18829,N_18655);
nand U19367 (N_19367,N_18739,N_18803);
nor U19368 (N_19368,N_18947,N_18858);
nor U19369 (N_19369,N_18763,N_18748);
nor U19370 (N_19370,N_18546,N_18991);
or U19371 (N_19371,N_18606,N_18536);
nor U19372 (N_19372,N_18647,N_18635);
and U19373 (N_19373,N_18820,N_18607);
nand U19374 (N_19374,N_18733,N_18503);
and U19375 (N_19375,N_18639,N_18711);
or U19376 (N_19376,N_18645,N_18678);
xnor U19377 (N_19377,N_18688,N_18939);
or U19378 (N_19378,N_18946,N_18978);
or U19379 (N_19379,N_18941,N_18843);
nor U19380 (N_19380,N_18692,N_18613);
nand U19381 (N_19381,N_18691,N_18765);
xnor U19382 (N_19382,N_18741,N_18555);
nand U19383 (N_19383,N_18929,N_18691);
and U19384 (N_19384,N_18974,N_18769);
nand U19385 (N_19385,N_18750,N_18845);
nand U19386 (N_19386,N_18703,N_18755);
nand U19387 (N_19387,N_18942,N_18726);
nand U19388 (N_19388,N_18688,N_18638);
xnor U19389 (N_19389,N_18558,N_18570);
xnor U19390 (N_19390,N_18830,N_18847);
nand U19391 (N_19391,N_18561,N_18951);
nor U19392 (N_19392,N_18763,N_18757);
or U19393 (N_19393,N_18576,N_18733);
xor U19394 (N_19394,N_18891,N_18720);
xor U19395 (N_19395,N_18879,N_18755);
or U19396 (N_19396,N_18810,N_18699);
nand U19397 (N_19397,N_18851,N_18615);
xor U19398 (N_19398,N_18688,N_18789);
nor U19399 (N_19399,N_18977,N_18840);
xnor U19400 (N_19400,N_18761,N_18993);
nor U19401 (N_19401,N_18805,N_18995);
nor U19402 (N_19402,N_18868,N_18964);
nand U19403 (N_19403,N_18913,N_18655);
nand U19404 (N_19404,N_18582,N_18658);
and U19405 (N_19405,N_18758,N_18865);
or U19406 (N_19406,N_18620,N_18901);
and U19407 (N_19407,N_18569,N_18945);
nand U19408 (N_19408,N_18604,N_18692);
nand U19409 (N_19409,N_18518,N_18867);
nor U19410 (N_19410,N_18638,N_18903);
nand U19411 (N_19411,N_18604,N_18960);
nor U19412 (N_19412,N_18927,N_18747);
nand U19413 (N_19413,N_18901,N_18688);
or U19414 (N_19414,N_18594,N_18892);
and U19415 (N_19415,N_18701,N_18910);
nor U19416 (N_19416,N_18570,N_18505);
nand U19417 (N_19417,N_18711,N_18984);
nand U19418 (N_19418,N_18717,N_18574);
or U19419 (N_19419,N_18547,N_18989);
nor U19420 (N_19420,N_18711,N_18701);
and U19421 (N_19421,N_18559,N_18870);
xor U19422 (N_19422,N_18645,N_18553);
or U19423 (N_19423,N_18742,N_18530);
nand U19424 (N_19424,N_18961,N_18781);
or U19425 (N_19425,N_18873,N_18712);
or U19426 (N_19426,N_18573,N_18991);
or U19427 (N_19427,N_18929,N_18582);
xnor U19428 (N_19428,N_18817,N_18876);
xnor U19429 (N_19429,N_18896,N_18817);
xor U19430 (N_19430,N_18766,N_18945);
nand U19431 (N_19431,N_18889,N_18791);
or U19432 (N_19432,N_18793,N_18586);
xor U19433 (N_19433,N_18691,N_18728);
nor U19434 (N_19434,N_18962,N_18807);
or U19435 (N_19435,N_18874,N_18772);
nand U19436 (N_19436,N_18940,N_18901);
xnor U19437 (N_19437,N_18665,N_18953);
xnor U19438 (N_19438,N_18644,N_18502);
or U19439 (N_19439,N_18521,N_18629);
xor U19440 (N_19440,N_18614,N_18865);
nor U19441 (N_19441,N_18660,N_18800);
or U19442 (N_19442,N_18661,N_18989);
xnor U19443 (N_19443,N_18829,N_18654);
xor U19444 (N_19444,N_18923,N_18700);
xnor U19445 (N_19445,N_18701,N_18584);
xor U19446 (N_19446,N_18757,N_18779);
nand U19447 (N_19447,N_18816,N_18635);
or U19448 (N_19448,N_18864,N_18790);
nand U19449 (N_19449,N_18792,N_18694);
nand U19450 (N_19450,N_18649,N_18783);
nor U19451 (N_19451,N_18943,N_18919);
xor U19452 (N_19452,N_18583,N_18696);
or U19453 (N_19453,N_18657,N_18534);
nand U19454 (N_19454,N_18772,N_18645);
and U19455 (N_19455,N_18771,N_18858);
nor U19456 (N_19456,N_18733,N_18747);
and U19457 (N_19457,N_18592,N_18913);
nor U19458 (N_19458,N_18882,N_18856);
or U19459 (N_19459,N_18589,N_18842);
or U19460 (N_19460,N_18551,N_18596);
xor U19461 (N_19461,N_18742,N_18830);
and U19462 (N_19462,N_18911,N_18629);
nand U19463 (N_19463,N_18711,N_18526);
nand U19464 (N_19464,N_18849,N_18836);
and U19465 (N_19465,N_18967,N_18597);
nor U19466 (N_19466,N_18893,N_18662);
nand U19467 (N_19467,N_18508,N_18970);
and U19468 (N_19468,N_18754,N_18612);
and U19469 (N_19469,N_18926,N_18806);
or U19470 (N_19470,N_18791,N_18866);
nand U19471 (N_19471,N_18843,N_18914);
and U19472 (N_19472,N_18902,N_18679);
or U19473 (N_19473,N_18987,N_18858);
or U19474 (N_19474,N_18698,N_18607);
and U19475 (N_19475,N_18967,N_18578);
nand U19476 (N_19476,N_18824,N_18700);
nor U19477 (N_19477,N_18610,N_18950);
nand U19478 (N_19478,N_18891,N_18582);
or U19479 (N_19479,N_18699,N_18633);
nand U19480 (N_19480,N_18911,N_18616);
and U19481 (N_19481,N_18531,N_18724);
nand U19482 (N_19482,N_18655,N_18798);
xor U19483 (N_19483,N_18637,N_18907);
xnor U19484 (N_19484,N_18739,N_18988);
nor U19485 (N_19485,N_18726,N_18532);
and U19486 (N_19486,N_18610,N_18903);
nor U19487 (N_19487,N_18631,N_18644);
or U19488 (N_19488,N_18574,N_18648);
and U19489 (N_19489,N_18753,N_18811);
and U19490 (N_19490,N_18674,N_18845);
nor U19491 (N_19491,N_18933,N_18709);
or U19492 (N_19492,N_18822,N_18715);
or U19493 (N_19493,N_18536,N_18965);
and U19494 (N_19494,N_18760,N_18523);
and U19495 (N_19495,N_18854,N_18736);
xnor U19496 (N_19496,N_18547,N_18528);
nand U19497 (N_19497,N_18994,N_18594);
xnor U19498 (N_19498,N_18629,N_18658);
nand U19499 (N_19499,N_18809,N_18624);
nand U19500 (N_19500,N_19039,N_19156);
nand U19501 (N_19501,N_19471,N_19406);
and U19502 (N_19502,N_19239,N_19004);
nand U19503 (N_19503,N_19070,N_19198);
and U19504 (N_19504,N_19058,N_19488);
nor U19505 (N_19505,N_19468,N_19451);
and U19506 (N_19506,N_19344,N_19258);
nand U19507 (N_19507,N_19150,N_19281);
nor U19508 (N_19508,N_19171,N_19262);
nor U19509 (N_19509,N_19118,N_19394);
and U19510 (N_19510,N_19135,N_19244);
xor U19511 (N_19511,N_19484,N_19028);
xnor U19512 (N_19512,N_19470,N_19287);
or U19513 (N_19513,N_19276,N_19243);
nor U19514 (N_19514,N_19013,N_19452);
nor U19515 (N_19515,N_19286,N_19222);
nor U19516 (N_19516,N_19352,N_19341);
nor U19517 (N_19517,N_19494,N_19428);
or U19518 (N_19518,N_19224,N_19020);
nand U19519 (N_19519,N_19082,N_19242);
and U19520 (N_19520,N_19404,N_19146);
nor U19521 (N_19521,N_19435,N_19040);
nand U19522 (N_19522,N_19154,N_19308);
nand U19523 (N_19523,N_19457,N_19097);
xnor U19524 (N_19524,N_19087,N_19057);
and U19525 (N_19525,N_19351,N_19195);
nor U19526 (N_19526,N_19003,N_19054);
and U19527 (N_19527,N_19279,N_19012);
xor U19528 (N_19528,N_19310,N_19173);
or U19529 (N_19529,N_19085,N_19424);
xor U19530 (N_19530,N_19208,N_19437);
nor U19531 (N_19531,N_19228,N_19438);
and U19532 (N_19532,N_19165,N_19177);
nand U19533 (N_19533,N_19260,N_19147);
nand U19534 (N_19534,N_19001,N_19014);
or U19535 (N_19535,N_19072,N_19292);
or U19536 (N_19536,N_19024,N_19130);
and U19537 (N_19537,N_19353,N_19053);
and U19538 (N_19538,N_19075,N_19196);
xor U19539 (N_19539,N_19304,N_19373);
or U19540 (N_19540,N_19176,N_19194);
nand U19541 (N_19541,N_19269,N_19267);
and U19542 (N_19542,N_19095,N_19375);
nand U19543 (N_19543,N_19343,N_19068);
or U19544 (N_19544,N_19491,N_19407);
nor U19545 (N_19545,N_19385,N_19137);
and U19546 (N_19546,N_19164,N_19285);
or U19547 (N_19547,N_19257,N_19300);
nand U19548 (N_19548,N_19172,N_19100);
nor U19549 (N_19549,N_19074,N_19030);
nor U19550 (N_19550,N_19056,N_19007);
and U19551 (N_19551,N_19124,N_19323);
nor U19552 (N_19552,N_19157,N_19337);
nand U19553 (N_19553,N_19212,N_19312);
nor U19554 (N_19554,N_19047,N_19240);
xor U19555 (N_19555,N_19380,N_19487);
and U19556 (N_19556,N_19210,N_19241);
nor U19557 (N_19557,N_19180,N_19005);
xor U19558 (N_19558,N_19339,N_19103);
nor U19559 (N_19559,N_19037,N_19334);
nand U19560 (N_19560,N_19393,N_19062);
xnor U19561 (N_19561,N_19220,N_19492);
xnor U19562 (N_19562,N_19099,N_19088);
xor U19563 (N_19563,N_19204,N_19255);
xnor U19564 (N_19564,N_19418,N_19076);
or U19565 (N_19565,N_19219,N_19271);
nor U19566 (N_19566,N_19283,N_19248);
or U19567 (N_19567,N_19402,N_19266);
xor U19568 (N_19568,N_19144,N_19361);
and U19569 (N_19569,N_19282,N_19356);
nand U19570 (N_19570,N_19307,N_19441);
or U19571 (N_19571,N_19066,N_19202);
nor U19572 (N_19572,N_19469,N_19446);
or U19573 (N_19573,N_19377,N_19387);
or U19574 (N_19574,N_19365,N_19277);
or U19575 (N_19575,N_19122,N_19139);
nand U19576 (N_19576,N_19134,N_19408);
or U19577 (N_19577,N_19372,N_19223);
xnor U19578 (N_19578,N_19415,N_19362);
nor U19579 (N_19579,N_19252,N_19495);
or U19580 (N_19580,N_19152,N_19386);
nor U19581 (N_19581,N_19143,N_19006);
xnor U19582 (N_19582,N_19273,N_19429);
or U19583 (N_19583,N_19297,N_19008);
nand U19584 (N_19584,N_19493,N_19083);
nand U19585 (N_19585,N_19367,N_19453);
nor U19586 (N_19586,N_19140,N_19280);
nor U19587 (N_19587,N_19116,N_19476);
or U19588 (N_19588,N_19059,N_19160);
nor U19589 (N_19589,N_19063,N_19060);
nor U19590 (N_19590,N_19187,N_19462);
nand U19591 (N_19591,N_19032,N_19482);
or U19592 (N_19592,N_19093,N_19168);
or U19593 (N_19593,N_19481,N_19268);
and U19594 (N_19594,N_19275,N_19483);
or U19595 (N_19595,N_19142,N_19159);
or U19596 (N_19596,N_19018,N_19138);
and U19597 (N_19597,N_19296,N_19309);
and U19598 (N_19598,N_19071,N_19126);
xor U19599 (N_19599,N_19169,N_19336);
and U19600 (N_19600,N_19274,N_19369);
or U19601 (N_19601,N_19213,N_19111);
xnor U19602 (N_19602,N_19426,N_19414);
xor U19603 (N_19603,N_19330,N_19403);
nor U19604 (N_19604,N_19236,N_19302);
xnor U19605 (N_19605,N_19325,N_19232);
or U19606 (N_19606,N_19349,N_19026);
xor U19607 (N_19607,N_19025,N_19329);
xor U19608 (N_19608,N_19303,N_19161);
xnor U19609 (N_19609,N_19129,N_19316);
nor U19610 (N_19610,N_19151,N_19199);
nand U19611 (N_19611,N_19288,N_19185);
and U19612 (N_19612,N_19413,N_19235);
or U19613 (N_19613,N_19259,N_19023);
and U19614 (N_19614,N_19479,N_19017);
xnor U19615 (N_19615,N_19324,N_19295);
nor U19616 (N_19616,N_19031,N_19158);
xor U19617 (N_19617,N_19460,N_19178);
and U19618 (N_19618,N_19465,N_19092);
xor U19619 (N_19619,N_19216,N_19132);
nand U19620 (N_19620,N_19427,N_19366);
or U19621 (N_19621,N_19350,N_19378);
xor U19622 (N_19622,N_19009,N_19278);
or U19623 (N_19623,N_19294,N_19077);
xnor U19624 (N_19624,N_19192,N_19474);
and U19625 (N_19625,N_19221,N_19417);
xnor U19626 (N_19626,N_19360,N_19049);
and U19627 (N_19627,N_19119,N_19061);
or U19628 (N_19628,N_19206,N_19027);
or U19629 (N_19629,N_19217,N_19141);
and U19630 (N_19630,N_19454,N_19321);
or U19631 (N_19631,N_19284,N_19133);
and U19632 (N_19632,N_19079,N_19496);
nand U19633 (N_19633,N_19015,N_19376);
or U19634 (N_19634,N_19473,N_19042);
nor U19635 (N_19635,N_19166,N_19382);
or U19636 (N_19636,N_19332,N_19211);
and U19637 (N_19637,N_19046,N_19113);
nor U19638 (N_19638,N_19225,N_19395);
and U19639 (N_19639,N_19123,N_19251);
nor U19640 (N_19640,N_19117,N_19357);
nor U19641 (N_19641,N_19253,N_19162);
or U19642 (N_19642,N_19209,N_19186);
nand U19643 (N_19643,N_19264,N_19010);
nand U19644 (N_19644,N_19080,N_19333);
and U19645 (N_19645,N_19226,N_19036);
and U19646 (N_19646,N_19381,N_19214);
nor U19647 (N_19647,N_19089,N_19348);
or U19648 (N_19648,N_19354,N_19145);
or U19649 (N_19649,N_19136,N_19421);
or U19650 (N_19650,N_19247,N_19254);
xor U19651 (N_19651,N_19110,N_19319);
nor U19652 (N_19652,N_19455,N_19043);
and U19653 (N_19653,N_19094,N_19197);
xor U19654 (N_19654,N_19355,N_19498);
xnor U19655 (N_19655,N_19101,N_19148);
nand U19656 (N_19656,N_19184,N_19272);
or U19657 (N_19657,N_19363,N_19250);
nor U19658 (N_19658,N_19411,N_19078);
and U19659 (N_19659,N_19112,N_19121);
nor U19660 (N_19660,N_19230,N_19106);
and U19661 (N_19661,N_19486,N_19301);
and U19662 (N_19662,N_19000,N_19489);
nand U19663 (N_19663,N_19359,N_19478);
or U19664 (N_19664,N_19218,N_19298);
nor U19665 (N_19665,N_19405,N_19327);
nand U19666 (N_19666,N_19463,N_19398);
and U19667 (N_19667,N_19442,N_19425);
nor U19668 (N_19668,N_19466,N_19290);
and U19669 (N_19669,N_19374,N_19090);
or U19670 (N_19670,N_19035,N_19423);
or U19671 (N_19671,N_19399,N_19033);
or U19672 (N_19672,N_19444,N_19081);
or U19673 (N_19673,N_19456,N_19238);
nand U19674 (N_19674,N_19389,N_19318);
nand U19675 (N_19675,N_19191,N_19055);
xor U19676 (N_19676,N_19167,N_19490);
nand U19677 (N_19677,N_19115,N_19193);
xnor U19678 (N_19678,N_19422,N_19419);
xor U19679 (N_19679,N_19261,N_19458);
nor U19680 (N_19680,N_19439,N_19201);
xnor U19681 (N_19681,N_19231,N_19342);
xnor U19682 (N_19682,N_19459,N_19155);
xor U19683 (N_19683,N_19170,N_19450);
or U19684 (N_19684,N_19189,N_19249);
and U19685 (N_19685,N_19091,N_19289);
and U19686 (N_19686,N_19125,N_19190);
nand U19687 (N_19687,N_19497,N_19434);
nor U19688 (N_19688,N_19461,N_19328);
or U19689 (N_19689,N_19396,N_19397);
and U19690 (N_19690,N_19364,N_19480);
or U19691 (N_19691,N_19345,N_19021);
nand U19692 (N_19692,N_19065,N_19163);
nand U19693 (N_19693,N_19041,N_19368);
xnor U19694 (N_19694,N_19207,N_19326);
or U19695 (N_19695,N_19270,N_19215);
and U19696 (N_19696,N_19313,N_19044);
nand U19697 (N_19697,N_19098,N_19420);
xnor U19698 (N_19698,N_19064,N_19051);
xnor U19699 (N_19699,N_19400,N_19379);
nor U19700 (N_19700,N_19346,N_19317);
or U19701 (N_19701,N_19069,N_19067);
and U19702 (N_19702,N_19485,N_19449);
nor U19703 (N_19703,N_19200,N_19002);
nand U19704 (N_19704,N_19314,N_19320);
or U19705 (N_19705,N_19096,N_19108);
nor U19706 (N_19706,N_19412,N_19305);
nand U19707 (N_19707,N_19315,N_19430);
nor U19708 (N_19708,N_19034,N_19467);
nand U19709 (N_19709,N_19011,N_19388);
nand U19710 (N_19710,N_19038,N_19390);
and U19711 (N_19711,N_19203,N_19183);
xnor U19712 (N_19712,N_19182,N_19464);
nor U19713 (N_19713,N_19401,N_19416);
and U19714 (N_19714,N_19358,N_19181);
nor U19715 (N_19715,N_19127,N_19149);
nand U19716 (N_19716,N_19477,N_19256);
nor U19717 (N_19717,N_19188,N_19107);
and U19718 (N_19718,N_19432,N_19246);
or U19719 (N_19719,N_19335,N_19436);
nor U19720 (N_19720,N_19306,N_19331);
and U19721 (N_19721,N_19174,N_19019);
or U19722 (N_19722,N_19073,N_19050);
xnor U19723 (N_19723,N_19131,N_19029);
xnor U19724 (N_19724,N_19371,N_19384);
and U19725 (N_19725,N_19120,N_19445);
nor U19726 (N_19726,N_19447,N_19052);
or U19727 (N_19727,N_19114,N_19048);
nor U19728 (N_19728,N_19499,N_19263);
nand U19729 (N_19729,N_19179,N_19392);
xnor U19730 (N_19730,N_19409,N_19265);
xor U19731 (N_19731,N_19299,N_19084);
or U19732 (N_19732,N_19233,N_19448);
and U19733 (N_19733,N_19022,N_19237);
xnor U19734 (N_19734,N_19234,N_19433);
or U19735 (N_19735,N_19370,N_19205);
or U19736 (N_19736,N_19475,N_19153);
and U19737 (N_19737,N_19322,N_19431);
xor U19738 (N_19738,N_19086,N_19383);
nand U19739 (N_19739,N_19391,N_19293);
nor U19740 (N_19740,N_19128,N_19045);
nor U19741 (N_19741,N_19229,N_19105);
nor U19742 (N_19742,N_19347,N_19104);
nor U19743 (N_19743,N_19443,N_19410);
xnor U19744 (N_19744,N_19291,N_19227);
nand U19745 (N_19745,N_19175,N_19472);
or U19746 (N_19746,N_19338,N_19340);
nor U19747 (N_19747,N_19245,N_19440);
nor U19748 (N_19748,N_19102,N_19311);
xnor U19749 (N_19749,N_19109,N_19016);
nand U19750 (N_19750,N_19434,N_19225);
and U19751 (N_19751,N_19056,N_19423);
xnor U19752 (N_19752,N_19344,N_19469);
or U19753 (N_19753,N_19159,N_19015);
nand U19754 (N_19754,N_19334,N_19171);
and U19755 (N_19755,N_19262,N_19257);
or U19756 (N_19756,N_19156,N_19103);
xor U19757 (N_19757,N_19222,N_19125);
xnor U19758 (N_19758,N_19082,N_19079);
nand U19759 (N_19759,N_19402,N_19142);
or U19760 (N_19760,N_19300,N_19379);
nor U19761 (N_19761,N_19092,N_19157);
or U19762 (N_19762,N_19441,N_19103);
or U19763 (N_19763,N_19250,N_19221);
nor U19764 (N_19764,N_19013,N_19017);
nor U19765 (N_19765,N_19180,N_19296);
and U19766 (N_19766,N_19191,N_19334);
xor U19767 (N_19767,N_19389,N_19464);
xor U19768 (N_19768,N_19147,N_19223);
nor U19769 (N_19769,N_19447,N_19013);
nor U19770 (N_19770,N_19174,N_19363);
or U19771 (N_19771,N_19314,N_19203);
or U19772 (N_19772,N_19282,N_19152);
xor U19773 (N_19773,N_19319,N_19279);
nand U19774 (N_19774,N_19308,N_19058);
nor U19775 (N_19775,N_19049,N_19064);
and U19776 (N_19776,N_19361,N_19213);
nand U19777 (N_19777,N_19214,N_19316);
nor U19778 (N_19778,N_19468,N_19218);
nor U19779 (N_19779,N_19289,N_19184);
or U19780 (N_19780,N_19358,N_19162);
or U19781 (N_19781,N_19311,N_19206);
nor U19782 (N_19782,N_19125,N_19421);
nand U19783 (N_19783,N_19130,N_19414);
nand U19784 (N_19784,N_19051,N_19067);
nand U19785 (N_19785,N_19243,N_19407);
nor U19786 (N_19786,N_19342,N_19381);
or U19787 (N_19787,N_19041,N_19460);
xor U19788 (N_19788,N_19088,N_19156);
nand U19789 (N_19789,N_19015,N_19311);
nand U19790 (N_19790,N_19311,N_19184);
xnor U19791 (N_19791,N_19250,N_19142);
xor U19792 (N_19792,N_19126,N_19477);
xnor U19793 (N_19793,N_19382,N_19491);
or U19794 (N_19794,N_19474,N_19180);
and U19795 (N_19795,N_19093,N_19247);
nor U19796 (N_19796,N_19301,N_19107);
or U19797 (N_19797,N_19091,N_19329);
nor U19798 (N_19798,N_19232,N_19282);
xor U19799 (N_19799,N_19301,N_19370);
xor U19800 (N_19800,N_19317,N_19343);
xnor U19801 (N_19801,N_19038,N_19401);
nand U19802 (N_19802,N_19111,N_19405);
nand U19803 (N_19803,N_19330,N_19198);
nand U19804 (N_19804,N_19154,N_19101);
and U19805 (N_19805,N_19303,N_19498);
and U19806 (N_19806,N_19040,N_19149);
or U19807 (N_19807,N_19257,N_19408);
or U19808 (N_19808,N_19452,N_19314);
and U19809 (N_19809,N_19135,N_19078);
or U19810 (N_19810,N_19152,N_19078);
and U19811 (N_19811,N_19431,N_19448);
nor U19812 (N_19812,N_19022,N_19081);
nor U19813 (N_19813,N_19403,N_19159);
and U19814 (N_19814,N_19214,N_19494);
nor U19815 (N_19815,N_19231,N_19242);
and U19816 (N_19816,N_19024,N_19058);
nor U19817 (N_19817,N_19248,N_19360);
nand U19818 (N_19818,N_19443,N_19368);
xor U19819 (N_19819,N_19049,N_19200);
nand U19820 (N_19820,N_19468,N_19353);
nand U19821 (N_19821,N_19131,N_19108);
and U19822 (N_19822,N_19158,N_19236);
nand U19823 (N_19823,N_19356,N_19131);
and U19824 (N_19824,N_19454,N_19331);
nand U19825 (N_19825,N_19349,N_19076);
and U19826 (N_19826,N_19243,N_19063);
nand U19827 (N_19827,N_19131,N_19217);
nor U19828 (N_19828,N_19449,N_19167);
xor U19829 (N_19829,N_19401,N_19325);
xnor U19830 (N_19830,N_19205,N_19387);
and U19831 (N_19831,N_19341,N_19253);
xnor U19832 (N_19832,N_19426,N_19320);
or U19833 (N_19833,N_19017,N_19160);
nor U19834 (N_19834,N_19062,N_19037);
or U19835 (N_19835,N_19437,N_19023);
nand U19836 (N_19836,N_19027,N_19467);
xnor U19837 (N_19837,N_19167,N_19351);
nor U19838 (N_19838,N_19362,N_19493);
nand U19839 (N_19839,N_19426,N_19397);
xnor U19840 (N_19840,N_19141,N_19199);
xnor U19841 (N_19841,N_19035,N_19030);
nand U19842 (N_19842,N_19102,N_19145);
xnor U19843 (N_19843,N_19112,N_19067);
nand U19844 (N_19844,N_19218,N_19082);
nand U19845 (N_19845,N_19462,N_19073);
nor U19846 (N_19846,N_19437,N_19317);
or U19847 (N_19847,N_19058,N_19125);
nand U19848 (N_19848,N_19441,N_19332);
nand U19849 (N_19849,N_19340,N_19482);
nor U19850 (N_19850,N_19108,N_19414);
nor U19851 (N_19851,N_19285,N_19427);
nor U19852 (N_19852,N_19426,N_19035);
nand U19853 (N_19853,N_19206,N_19354);
or U19854 (N_19854,N_19493,N_19343);
nor U19855 (N_19855,N_19063,N_19202);
and U19856 (N_19856,N_19246,N_19054);
and U19857 (N_19857,N_19280,N_19027);
nor U19858 (N_19858,N_19337,N_19320);
nor U19859 (N_19859,N_19446,N_19292);
nand U19860 (N_19860,N_19470,N_19358);
or U19861 (N_19861,N_19304,N_19191);
and U19862 (N_19862,N_19361,N_19461);
or U19863 (N_19863,N_19074,N_19426);
and U19864 (N_19864,N_19135,N_19347);
and U19865 (N_19865,N_19247,N_19200);
xnor U19866 (N_19866,N_19411,N_19352);
and U19867 (N_19867,N_19434,N_19243);
nor U19868 (N_19868,N_19409,N_19093);
and U19869 (N_19869,N_19177,N_19075);
nor U19870 (N_19870,N_19317,N_19246);
or U19871 (N_19871,N_19495,N_19496);
nor U19872 (N_19872,N_19285,N_19474);
xnor U19873 (N_19873,N_19394,N_19459);
xor U19874 (N_19874,N_19400,N_19468);
or U19875 (N_19875,N_19322,N_19302);
nand U19876 (N_19876,N_19301,N_19343);
and U19877 (N_19877,N_19276,N_19119);
and U19878 (N_19878,N_19227,N_19266);
xor U19879 (N_19879,N_19463,N_19355);
and U19880 (N_19880,N_19448,N_19488);
nor U19881 (N_19881,N_19033,N_19209);
nor U19882 (N_19882,N_19405,N_19029);
nor U19883 (N_19883,N_19231,N_19114);
and U19884 (N_19884,N_19226,N_19387);
or U19885 (N_19885,N_19187,N_19117);
and U19886 (N_19886,N_19333,N_19120);
or U19887 (N_19887,N_19066,N_19136);
nand U19888 (N_19888,N_19306,N_19075);
xor U19889 (N_19889,N_19360,N_19092);
or U19890 (N_19890,N_19423,N_19481);
or U19891 (N_19891,N_19266,N_19084);
nor U19892 (N_19892,N_19114,N_19422);
nor U19893 (N_19893,N_19257,N_19296);
and U19894 (N_19894,N_19010,N_19165);
xor U19895 (N_19895,N_19307,N_19429);
and U19896 (N_19896,N_19156,N_19157);
or U19897 (N_19897,N_19323,N_19401);
xnor U19898 (N_19898,N_19218,N_19401);
xnor U19899 (N_19899,N_19464,N_19345);
nor U19900 (N_19900,N_19487,N_19470);
nand U19901 (N_19901,N_19217,N_19340);
nand U19902 (N_19902,N_19047,N_19039);
nor U19903 (N_19903,N_19405,N_19488);
nor U19904 (N_19904,N_19447,N_19046);
nor U19905 (N_19905,N_19129,N_19452);
and U19906 (N_19906,N_19090,N_19115);
and U19907 (N_19907,N_19040,N_19371);
or U19908 (N_19908,N_19120,N_19385);
nand U19909 (N_19909,N_19458,N_19499);
or U19910 (N_19910,N_19351,N_19489);
nand U19911 (N_19911,N_19348,N_19016);
nand U19912 (N_19912,N_19186,N_19353);
nand U19913 (N_19913,N_19145,N_19269);
xnor U19914 (N_19914,N_19182,N_19384);
nor U19915 (N_19915,N_19492,N_19127);
xor U19916 (N_19916,N_19247,N_19447);
nor U19917 (N_19917,N_19041,N_19300);
nor U19918 (N_19918,N_19182,N_19111);
xor U19919 (N_19919,N_19442,N_19320);
nor U19920 (N_19920,N_19117,N_19317);
or U19921 (N_19921,N_19175,N_19149);
nor U19922 (N_19922,N_19479,N_19099);
nor U19923 (N_19923,N_19374,N_19423);
xor U19924 (N_19924,N_19014,N_19268);
xor U19925 (N_19925,N_19450,N_19405);
nor U19926 (N_19926,N_19107,N_19275);
nand U19927 (N_19927,N_19227,N_19332);
nor U19928 (N_19928,N_19458,N_19098);
nor U19929 (N_19929,N_19084,N_19306);
nand U19930 (N_19930,N_19127,N_19442);
or U19931 (N_19931,N_19196,N_19083);
nand U19932 (N_19932,N_19263,N_19168);
nand U19933 (N_19933,N_19109,N_19457);
or U19934 (N_19934,N_19178,N_19273);
or U19935 (N_19935,N_19231,N_19188);
or U19936 (N_19936,N_19312,N_19445);
or U19937 (N_19937,N_19023,N_19179);
nand U19938 (N_19938,N_19498,N_19366);
nor U19939 (N_19939,N_19083,N_19434);
xor U19940 (N_19940,N_19313,N_19096);
xnor U19941 (N_19941,N_19058,N_19314);
nor U19942 (N_19942,N_19264,N_19173);
and U19943 (N_19943,N_19231,N_19466);
xnor U19944 (N_19944,N_19012,N_19451);
and U19945 (N_19945,N_19379,N_19457);
or U19946 (N_19946,N_19355,N_19110);
or U19947 (N_19947,N_19422,N_19190);
or U19948 (N_19948,N_19469,N_19237);
nor U19949 (N_19949,N_19058,N_19331);
or U19950 (N_19950,N_19489,N_19481);
and U19951 (N_19951,N_19088,N_19137);
or U19952 (N_19952,N_19332,N_19225);
or U19953 (N_19953,N_19127,N_19488);
and U19954 (N_19954,N_19302,N_19432);
xor U19955 (N_19955,N_19446,N_19384);
or U19956 (N_19956,N_19102,N_19001);
xor U19957 (N_19957,N_19195,N_19162);
or U19958 (N_19958,N_19031,N_19285);
or U19959 (N_19959,N_19355,N_19123);
nor U19960 (N_19960,N_19482,N_19428);
nand U19961 (N_19961,N_19018,N_19259);
nand U19962 (N_19962,N_19064,N_19489);
xnor U19963 (N_19963,N_19190,N_19102);
nand U19964 (N_19964,N_19383,N_19368);
or U19965 (N_19965,N_19077,N_19107);
and U19966 (N_19966,N_19461,N_19142);
or U19967 (N_19967,N_19027,N_19279);
nor U19968 (N_19968,N_19008,N_19141);
xor U19969 (N_19969,N_19316,N_19010);
xnor U19970 (N_19970,N_19333,N_19264);
and U19971 (N_19971,N_19317,N_19210);
nor U19972 (N_19972,N_19308,N_19080);
nor U19973 (N_19973,N_19173,N_19249);
nand U19974 (N_19974,N_19135,N_19110);
nand U19975 (N_19975,N_19332,N_19498);
or U19976 (N_19976,N_19035,N_19184);
xnor U19977 (N_19977,N_19303,N_19356);
and U19978 (N_19978,N_19333,N_19188);
nor U19979 (N_19979,N_19153,N_19122);
xor U19980 (N_19980,N_19315,N_19369);
nand U19981 (N_19981,N_19027,N_19225);
and U19982 (N_19982,N_19398,N_19404);
or U19983 (N_19983,N_19097,N_19157);
or U19984 (N_19984,N_19056,N_19091);
and U19985 (N_19985,N_19056,N_19236);
nand U19986 (N_19986,N_19302,N_19064);
or U19987 (N_19987,N_19058,N_19332);
or U19988 (N_19988,N_19292,N_19014);
nor U19989 (N_19989,N_19026,N_19045);
nor U19990 (N_19990,N_19299,N_19083);
or U19991 (N_19991,N_19204,N_19353);
nand U19992 (N_19992,N_19299,N_19480);
and U19993 (N_19993,N_19353,N_19298);
or U19994 (N_19994,N_19441,N_19403);
and U19995 (N_19995,N_19145,N_19329);
and U19996 (N_19996,N_19368,N_19386);
and U19997 (N_19997,N_19020,N_19473);
or U19998 (N_19998,N_19409,N_19347);
or U19999 (N_19999,N_19153,N_19024);
xnor UO_0 (O_0,N_19810,N_19962);
nor UO_1 (O_1,N_19626,N_19539);
nand UO_2 (O_2,N_19970,N_19611);
or UO_3 (O_3,N_19955,N_19540);
or UO_4 (O_4,N_19673,N_19663);
or UO_5 (O_5,N_19922,N_19820);
and UO_6 (O_6,N_19590,N_19722);
nor UO_7 (O_7,N_19711,N_19812);
xnor UO_8 (O_8,N_19500,N_19901);
nor UO_9 (O_9,N_19522,N_19573);
nor UO_10 (O_10,N_19797,N_19681);
and UO_11 (O_11,N_19815,N_19583);
xnor UO_12 (O_12,N_19974,N_19758);
and UO_13 (O_13,N_19562,N_19998);
or UO_14 (O_14,N_19732,N_19730);
xor UO_15 (O_15,N_19863,N_19642);
nand UO_16 (O_16,N_19789,N_19875);
and UO_17 (O_17,N_19623,N_19734);
nor UO_18 (O_18,N_19741,N_19588);
or UO_19 (O_19,N_19825,N_19617);
and UO_20 (O_20,N_19826,N_19871);
xor UO_21 (O_21,N_19659,N_19733);
nor UO_22 (O_22,N_19802,N_19639);
and UO_23 (O_23,N_19740,N_19839);
and UO_24 (O_24,N_19912,N_19677);
or UO_25 (O_25,N_19838,N_19918);
nor UO_26 (O_26,N_19965,N_19716);
or UO_27 (O_27,N_19557,N_19902);
nand UO_28 (O_28,N_19641,N_19811);
nor UO_29 (O_29,N_19542,N_19571);
nor UO_30 (O_30,N_19682,N_19903);
or UO_31 (O_31,N_19742,N_19849);
xor UO_32 (O_32,N_19801,N_19896);
xor UO_33 (O_33,N_19745,N_19746);
or UO_34 (O_34,N_19701,N_19926);
xor UO_35 (O_35,N_19973,N_19579);
and UO_36 (O_36,N_19771,N_19782);
xor UO_37 (O_37,N_19967,N_19774);
nand UO_38 (O_38,N_19747,N_19691);
or UO_39 (O_39,N_19828,N_19845);
nand UO_40 (O_40,N_19976,N_19997);
nor UO_41 (O_41,N_19987,N_19989);
or UO_42 (O_42,N_19553,N_19505);
xnor UO_43 (O_43,N_19556,N_19808);
and UO_44 (O_44,N_19610,N_19616);
and UO_45 (O_45,N_19506,N_19514);
or UO_46 (O_46,N_19813,N_19925);
or UO_47 (O_47,N_19675,N_19531);
or UO_48 (O_48,N_19900,N_19979);
or UO_49 (O_49,N_19957,N_19543);
nor UO_50 (O_50,N_19868,N_19818);
nand UO_51 (O_51,N_19630,N_19859);
and UO_52 (O_52,N_19708,N_19763);
nand UO_53 (O_53,N_19893,N_19779);
or UO_54 (O_54,N_19585,N_19744);
nor UO_55 (O_55,N_19950,N_19717);
and UO_56 (O_56,N_19516,N_19510);
or UO_57 (O_57,N_19715,N_19991);
and UO_58 (O_58,N_19830,N_19767);
nor UO_59 (O_59,N_19575,N_19586);
and UO_60 (O_60,N_19589,N_19928);
or UO_61 (O_61,N_19622,N_19865);
and UO_62 (O_62,N_19930,N_19574);
nand UO_63 (O_63,N_19555,N_19651);
xnor UO_64 (O_64,N_19644,N_19853);
nor UO_65 (O_65,N_19934,N_19944);
or UO_66 (O_66,N_19618,N_19857);
and UO_67 (O_67,N_19735,N_19657);
or UO_68 (O_68,N_19569,N_19705);
xnor UO_69 (O_69,N_19702,N_19911);
or UO_70 (O_70,N_19524,N_19655);
nand UO_71 (O_71,N_19798,N_19939);
nand UO_72 (O_72,N_19827,N_19821);
nand UO_73 (O_73,N_19731,N_19951);
and UO_74 (O_74,N_19707,N_19534);
nand UO_75 (O_75,N_19561,N_19796);
nor UO_76 (O_76,N_19560,N_19870);
xnor UO_77 (O_77,N_19958,N_19723);
nand UO_78 (O_78,N_19605,N_19597);
nor UO_79 (O_79,N_19846,N_19704);
xnor UO_80 (O_80,N_19832,N_19995);
or UO_81 (O_81,N_19791,N_19861);
nand UO_82 (O_82,N_19817,N_19598);
xor UO_83 (O_83,N_19592,N_19567);
and UO_84 (O_84,N_19593,N_19885);
or UO_85 (O_85,N_19608,N_19703);
nor UO_86 (O_86,N_19761,N_19897);
and UO_87 (O_87,N_19554,N_19959);
nand UO_88 (O_88,N_19546,N_19753);
nand UO_89 (O_89,N_19806,N_19916);
or UO_90 (O_90,N_19609,N_19517);
nand UO_91 (O_91,N_19835,N_19643);
xor UO_92 (O_92,N_19519,N_19872);
nor UO_93 (O_93,N_19824,N_19719);
and UO_94 (O_94,N_19752,N_19972);
xnor UO_95 (O_95,N_19736,N_19945);
nor UO_96 (O_96,N_19727,N_19721);
and UO_97 (O_97,N_19678,N_19980);
xor UO_98 (O_98,N_19653,N_19607);
nor UO_99 (O_99,N_19750,N_19679);
and UO_100 (O_100,N_19757,N_19851);
nand UO_101 (O_101,N_19513,N_19956);
or UO_102 (O_102,N_19619,N_19794);
or UO_103 (O_103,N_19776,N_19843);
nor UO_104 (O_104,N_19684,N_19578);
or UO_105 (O_105,N_19512,N_19847);
or UO_106 (O_106,N_19581,N_19614);
nor UO_107 (O_107,N_19823,N_19528);
nor UO_108 (O_108,N_19541,N_19961);
or UO_109 (O_109,N_19867,N_19940);
nor UO_110 (O_110,N_19726,N_19850);
nand UO_111 (O_111,N_19809,N_19603);
nor UO_112 (O_112,N_19756,N_19565);
nand UO_113 (O_113,N_19503,N_19892);
xnor UO_114 (O_114,N_19645,N_19671);
or UO_115 (O_115,N_19532,N_19613);
nand UO_116 (O_116,N_19631,N_19993);
nand UO_117 (O_117,N_19566,N_19587);
nor UO_118 (O_118,N_19739,N_19669);
nand UO_119 (O_119,N_19869,N_19982);
xor UO_120 (O_120,N_19908,N_19595);
or UO_121 (O_121,N_19814,N_19706);
and UO_122 (O_122,N_19840,N_19693);
or UO_123 (O_123,N_19737,N_19931);
nand UO_124 (O_124,N_19772,N_19879);
and UO_125 (O_125,N_19996,N_19977);
xnor UO_126 (O_126,N_19915,N_19952);
xnor UO_127 (O_127,N_19530,N_19615);
and UO_128 (O_128,N_19692,N_19690);
nor UO_129 (O_129,N_19844,N_19936);
nand UO_130 (O_130,N_19625,N_19547);
xnor UO_131 (O_131,N_19518,N_19921);
and UO_132 (O_132,N_19538,N_19968);
and UO_133 (O_133,N_19985,N_19971);
nor UO_134 (O_134,N_19783,N_19699);
nor UO_135 (O_135,N_19949,N_19960);
xor UO_136 (O_136,N_19759,N_19769);
nor UO_137 (O_137,N_19942,N_19933);
or UO_138 (O_138,N_19520,N_19672);
or UO_139 (O_139,N_19891,N_19685);
and UO_140 (O_140,N_19548,N_19729);
and UO_141 (O_141,N_19596,N_19656);
xnor UO_142 (O_142,N_19632,N_19620);
xnor UO_143 (O_143,N_19990,N_19768);
or UO_144 (O_144,N_19697,N_19895);
and UO_145 (O_145,N_19509,N_19627);
nand UO_146 (O_146,N_19986,N_19793);
or UO_147 (O_147,N_19963,N_19700);
nor UO_148 (O_148,N_19680,N_19787);
and UO_149 (O_149,N_19841,N_19856);
nor UO_150 (O_150,N_19646,N_19833);
and UO_151 (O_151,N_19580,N_19640);
nand UO_152 (O_152,N_19834,N_19764);
and UO_153 (O_153,N_19923,N_19687);
nor UO_154 (O_154,N_19909,N_19635);
and UO_155 (O_155,N_19748,N_19545);
nor UO_156 (O_156,N_19720,N_19866);
and UO_157 (O_157,N_19910,N_19889);
or UO_158 (O_158,N_19696,N_19662);
or UO_159 (O_159,N_19890,N_19978);
xor UO_160 (O_160,N_19508,N_19572);
or UO_161 (O_161,N_19943,N_19906);
and UO_162 (O_162,N_19983,N_19822);
and UO_163 (O_163,N_19914,N_19591);
nor UO_164 (O_164,N_19504,N_19738);
nor UO_165 (O_165,N_19754,N_19762);
and UO_166 (O_166,N_19981,N_19724);
nor UO_167 (O_167,N_19594,N_19852);
nor UO_168 (O_168,N_19648,N_19709);
xor UO_169 (O_169,N_19638,N_19984);
or UO_170 (O_170,N_19946,N_19948);
or UO_171 (O_171,N_19999,N_19947);
nand UO_172 (O_172,N_19848,N_19803);
and UO_173 (O_173,N_19533,N_19913);
or UO_174 (O_174,N_19881,N_19837);
and UO_175 (O_175,N_19988,N_19507);
and UO_176 (O_176,N_19676,N_19935);
and UO_177 (O_177,N_19695,N_19552);
nand UO_178 (O_178,N_19932,N_19694);
xor UO_179 (O_179,N_19523,N_19670);
nor UO_180 (O_180,N_19831,N_19873);
nor UO_181 (O_181,N_19501,N_19650);
nor UO_182 (O_182,N_19599,N_19886);
and UO_183 (O_183,N_19966,N_19621);
xor UO_184 (O_184,N_19689,N_19884);
or UO_185 (O_185,N_19874,N_19601);
nand UO_186 (O_186,N_19629,N_19877);
or UO_187 (O_187,N_19536,N_19725);
nor UO_188 (O_188,N_19521,N_19698);
nor UO_189 (O_189,N_19927,N_19511);
nor UO_190 (O_190,N_19778,N_19860);
nor UO_191 (O_191,N_19864,N_19660);
nor UO_192 (O_192,N_19712,N_19953);
nor UO_193 (O_193,N_19862,N_19559);
or UO_194 (O_194,N_19855,N_19907);
nor UO_195 (O_195,N_19920,N_19937);
or UO_196 (O_196,N_19785,N_19600);
and UO_197 (O_197,N_19558,N_19876);
xnor UO_198 (O_198,N_19602,N_19502);
or UO_199 (O_199,N_19674,N_19842);
and UO_200 (O_200,N_19624,N_19647);
nand UO_201 (O_201,N_19938,N_19535);
nor UO_202 (O_202,N_19544,N_19688);
or UO_203 (O_203,N_19604,N_19924);
xor UO_204 (O_204,N_19654,N_19929);
xnor UO_205 (O_205,N_19975,N_19665);
and UO_206 (O_206,N_19816,N_19775);
nand UO_207 (O_207,N_19898,N_19661);
xnor UO_208 (O_208,N_19683,N_19612);
nor UO_209 (O_209,N_19883,N_19686);
and UO_210 (O_210,N_19905,N_19766);
or UO_211 (O_211,N_19550,N_19664);
or UO_212 (O_212,N_19634,N_19628);
or UO_213 (O_213,N_19551,N_19765);
and UO_214 (O_214,N_19515,N_19577);
or UO_215 (O_215,N_19658,N_19807);
xnor UO_216 (O_216,N_19713,N_19829);
nand UO_217 (O_217,N_19854,N_19668);
nand UO_218 (O_218,N_19882,N_19564);
nand UO_219 (O_219,N_19633,N_19964);
xor UO_220 (O_220,N_19743,N_19666);
nand UO_221 (O_221,N_19941,N_19888);
nand UO_222 (O_222,N_19549,N_19527);
and UO_223 (O_223,N_19529,N_19718);
xnor UO_224 (O_224,N_19584,N_19994);
xnor UO_225 (O_225,N_19919,N_19710);
nor UO_226 (O_226,N_19804,N_19637);
nand UO_227 (O_227,N_19790,N_19805);
nand UO_228 (O_228,N_19954,N_19786);
nand UO_229 (O_229,N_19749,N_19568);
or UO_230 (O_230,N_19780,N_19760);
or UO_231 (O_231,N_19969,N_19714);
xor UO_232 (O_232,N_19878,N_19652);
and UO_233 (O_233,N_19992,N_19799);
nor UO_234 (O_234,N_19755,N_19537);
and UO_235 (O_235,N_19795,N_19649);
nor UO_236 (O_236,N_19917,N_19836);
nor UO_237 (O_237,N_19525,N_19570);
nand UO_238 (O_238,N_19606,N_19751);
or UO_239 (O_239,N_19899,N_19819);
xor UO_240 (O_240,N_19563,N_19728);
nand UO_241 (O_241,N_19894,N_19904);
xor UO_242 (O_242,N_19858,N_19667);
nor UO_243 (O_243,N_19777,N_19788);
nand UO_244 (O_244,N_19880,N_19576);
and UO_245 (O_245,N_19526,N_19887);
and UO_246 (O_246,N_19770,N_19800);
and UO_247 (O_247,N_19792,N_19781);
and UO_248 (O_248,N_19636,N_19784);
nor UO_249 (O_249,N_19582,N_19773);
nand UO_250 (O_250,N_19593,N_19729);
or UO_251 (O_251,N_19852,N_19898);
or UO_252 (O_252,N_19764,N_19614);
nor UO_253 (O_253,N_19582,N_19604);
or UO_254 (O_254,N_19592,N_19808);
or UO_255 (O_255,N_19841,N_19604);
and UO_256 (O_256,N_19772,N_19666);
xor UO_257 (O_257,N_19599,N_19641);
or UO_258 (O_258,N_19909,N_19646);
or UO_259 (O_259,N_19718,N_19842);
xor UO_260 (O_260,N_19791,N_19592);
or UO_261 (O_261,N_19620,N_19878);
and UO_262 (O_262,N_19831,N_19794);
and UO_263 (O_263,N_19606,N_19640);
nor UO_264 (O_264,N_19747,N_19596);
and UO_265 (O_265,N_19796,N_19742);
xor UO_266 (O_266,N_19749,N_19848);
nand UO_267 (O_267,N_19806,N_19957);
nor UO_268 (O_268,N_19840,N_19758);
nor UO_269 (O_269,N_19901,N_19851);
nand UO_270 (O_270,N_19889,N_19623);
nand UO_271 (O_271,N_19741,N_19718);
nor UO_272 (O_272,N_19702,N_19934);
or UO_273 (O_273,N_19585,N_19953);
xor UO_274 (O_274,N_19648,N_19966);
and UO_275 (O_275,N_19643,N_19896);
nor UO_276 (O_276,N_19983,N_19574);
xor UO_277 (O_277,N_19706,N_19579);
nor UO_278 (O_278,N_19773,N_19514);
and UO_279 (O_279,N_19506,N_19845);
and UO_280 (O_280,N_19923,N_19560);
xor UO_281 (O_281,N_19626,N_19944);
and UO_282 (O_282,N_19697,N_19687);
nor UO_283 (O_283,N_19936,N_19627);
or UO_284 (O_284,N_19956,N_19509);
xnor UO_285 (O_285,N_19935,N_19829);
and UO_286 (O_286,N_19627,N_19632);
nor UO_287 (O_287,N_19548,N_19925);
nor UO_288 (O_288,N_19895,N_19718);
and UO_289 (O_289,N_19622,N_19647);
nand UO_290 (O_290,N_19943,N_19875);
or UO_291 (O_291,N_19663,N_19844);
or UO_292 (O_292,N_19882,N_19810);
or UO_293 (O_293,N_19630,N_19781);
or UO_294 (O_294,N_19519,N_19679);
nand UO_295 (O_295,N_19807,N_19811);
and UO_296 (O_296,N_19600,N_19992);
xnor UO_297 (O_297,N_19794,N_19647);
and UO_298 (O_298,N_19989,N_19714);
nor UO_299 (O_299,N_19709,N_19716);
xor UO_300 (O_300,N_19528,N_19852);
and UO_301 (O_301,N_19810,N_19824);
nand UO_302 (O_302,N_19743,N_19558);
or UO_303 (O_303,N_19606,N_19519);
nand UO_304 (O_304,N_19873,N_19987);
or UO_305 (O_305,N_19545,N_19719);
xor UO_306 (O_306,N_19759,N_19643);
and UO_307 (O_307,N_19511,N_19517);
xnor UO_308 (O_308,N_19953,N_19610);
or UO_309 (O_309,N_19521,N_19962);
nand UO_310 (O_310,N_19830,N_19727);
nor UO_311 (O_311,N_19655,N_19763);
or UO_312 (O_312,N_19939,N_19905);
xor UO_313 (O_313,N_19911,N_19882);
nor UO_314 (O_314,N_19753,N_19532);
nor UO_315 (O_315,N_19685,N_19926);
nand UO_316 (O_316,N_19835,N_19602);
nand UO_317 (O_317,N_19834,N_19707);
nand UO_318 (O_318,N_19749,N_19881);
xor UO_319 (O_319,N_19918,N_19933);
xor UO_320 (O_320,N_19674,N_19589);
nor UO_321 (O_321,N_19503,N_19827);
or UO_322 (O_322,N_19845,N_19851);
nor UO_323 (O_323,N_19597,N_19910);
and UO_324 (O_324,N_19775,N_19602);
and UO_325 (O_325,N_19832,N_19656);
xnor UO_326 (O_326,N_19862,N_19587);
nand UO_327 (O_327,N_19638,N_19603);
nand UO_328 (O_328,N_19651,N_19957);
xor UO_329 (O_329,N_19514,N_19754);
or UO_330 (O_330,N_19941,N_19768);
nand UO_331 (O_331,N_19777,N_19832);
nand UO_332 (O_332,N_19759,N_19794);
nor UO_333 (O_333,N_19836,N_19546);
nand UO_334 (O_334,N_19868,N_19912);
and UO_335 (O_335,N_19858,N_19949);
xor UO_336 (O_336,N_19774,N_19870);
nor UO_337 (O_337,N_19997,N_19570);
nor UO_338 (O_338,N_19880,N_19769);
xor UO_339 (O_339,N_19875,N_19880);
nor UO_340 (O_340,N_19508,N_19953);
and UO_341 (O_341,N_19644,N_19949);
and UO_342 (O_342,N_19598,N_19849);
nor UO_343 (O_343,N_19881,N_19769);
xnor UO_344 (O_344,N_19637,N_19776);
and UO_345 (O_345,N_19958,N_19844);
nand UO_346 (O_346,N_19766,N_19785);
nor UO_347 (O_347,N_19608,N_19768);
or UO_348 (O_348,N_19733,N_19563);
xnor UO_349 (O_349,N_19688,N_19807);
or UO_350 (O_350,N_19580,N_19864);
nor UO_351 (O_351,N_19956,N_19941);
nand UO_352 (O_352,N_19861,N_19561);
nand UO_353 (O_353,N_19505,N_19612);
and UO_354 (O_354,N_19622,N_19780);
nand UO_355 (O_355,N_19925,N_19852);
and UO_356 (O_356,N_19843,N_19747);
or UO_357 (O_357,N_19875,N_19516);
and UO_358 (O_358,N_19653,N_19956);
nand UO_359 (O_359,N_19795,N_19868);
and UO_360 (O_360,N_19526,N_19989);
or UO_361 (O_361,N_19688,N_19783);
and UO_362 (O_362,N_19604,N_19639);
or UO_363 (O_363,N_19780,N_19556);
and UO_364 (O_364,N_19900,N_19964);
or UO_365 (O_365,N_19898,N_19807);
xor UO_366 (O_366,N_19998,N_19935);
xor UO_367 (O_367,N_19571,N_19845);
or UO_368 (O_368,N_19689,N_19856);
and UO_369 (O_369,N_19592,N_19522);
nand UO_370 (O_370,N_19964,N_19844);
xnor UO_371 (O_371,N_19659,N_19985);
nand UO_372 (O_372,N_19977,N_19889);
nor UO_373 (O_373,N_19708,N_19788);
and UO_374 (O_374,N_19990,N_19603);
xnor UO_375 (O_375,N_19545,N_19661);
and UO_376 (O_376,N_19604,N_19693);
nor UO_377 (O_377,N_19667,N_19522);
nor UO_378 (O_378,N_19930,N_19685);
xor UO_379 (O_379,N_19905,N_19829);
xor UO_380 (O_380,N_19871,N_19719);
or UO_381 (O_381,N_19900,N_19715);
xnor UO_382 (O_382,N_19827,N_19750);
or UO_383 (O_383,N_19750,N_19735);
or UO_384 (O_384,N_19624,N_19986);
xnor UO_385 (O_385,N_19956,N_19763);
and UO_386 (O_386,N_19734,N_19768);
xnor UO_387 (O_387,N_19513,N_19739);
xnor UO_388 (O_388,N_19770,N_19818);
nor UO_389 (O_389,N_19596,N_19941);
nor UO_390 (O_390,N_19952,N_19948);
xor UO_391 (O_391,N_19969,N_19891);
xnor UO_392 (O_392,N_19594,N_19798);
xnor UO_393 (O_393,N_19541,N_19552);
nand UO_394 (O_394,N_19875,N_19503);
and UO_395 (O_395,N_19739,N_19544);
nor UO_396 (O_396,N_19847,N_19899);
and UO_397 (O_397,N_19909,N_19625);
nand UO_398 (O_398,N_19643,N_19703);
nor UO_399 (O_399,N_19763,N_19741);
nand UO_400 (O_400,N_19850,N_19682);
and UO_401 (O_401,N_19792,N_19558);
nor UO_402 (O_402,N_19700,N_19989);
nand UO_403 (O_403,N_19873,N_19637);
nor UO_404 (O_404,N_19900,N_19654);
xnor UO_405 (O_405,N_19927,N_19918);
nand UO_406 (O_406,N_19898,N_19703);
or UO_407 (O_407,N_19765,N_19743);
nand UO_408 (O_408,N_19650,N_19579);
and UO_409 (O_409,N_19568,N_19573);
and UO_410 (O_410,N_19668,N_19679);
and UO_411 (O_411,N_19667,N_19705);
nand UO_412 (O_412,N_19671,N_19514);
or UO_413 (O_413,N_19911,N_19997);
xnor UO_414 (O_414,N_19924,N_19801);
and UO_415 (O_415,N_19618,N_19521);
nor UO_416 (O_416,N_19879,N_19853);
and UO_417 (O_417,N_19581,N_19850);
nor UO_418 (O_418,N_19980,N_19577);
nor UO_419 (O_419,N_19564,N_19739);
nor UO_420 (O_420,N_19684,N_19863);
nor UO_421 (O_421,N_19512,N_19912);
nor UO_422 (O_422,N_19775,N_19646);
nor UO_423 (O_423,N_19657,N_19653);
or UO_424 (O_424,N_19849,N_19810);
or UO_425 (O_425,N_19993,N_19965);
nor UO_426 (O_426,N_19678,N_19700);
or UO_427 (O_427,N_19795,N_19879);
xnor UO_428 (O_428,N_19676,N_19956);
nand UO_429 (O_429,N_19549,N_19994);
nor UO_430 (O_430,N_19625,N_19711);
nand UO_431 (O_431,N_19997,N_19566);
xnor UO_432 (O_432,N_19685,N_19920);
and UO_433 (O_433,N_19600,N_19770);
xor UO_434 (O_434,N_19855,N_19658);
or UO_435 (O_435,N_19516,N_19850);
nand UO_436 (O_436,N_19557,N_19820);
or UO_437 (O_437,N_19570,N_19964);
xor UO_438 (O_438,N_19935,N_19582);
nor UO_439 (O_439,N_19843,N_19973);
or UO_440 (O_440,N_19963,N_19959);
nand UO_441 (O_441,N_19520,N_19915);
nand UO_442 (O_442,N_19591,N_19875);
nor UO_443 (O_443,N_19810,N_19534);
xor UO_444 (O_444,N_19799,N_19596);
nor UO_445 (O_445,N_19695,N_19799);
nand UO_446 (O_446,N_19789,N_19901);
nor UO_447 (O_447,N_19958,N_19699);
and UO_448 (O_448,N_19786,N_19779);
and UO_449 (O_449,N_19958,N_19540);
or UO_450 (O_450,N_19773,N_19882);
and UO_451 (O_451,N_19559,N_19712);
nor UO_452 (O_452,N_19895,N_19875);
nand UO_453 (O_453,N_19705,N_19998);
nor UO_454 (O_454,N_19973,N_19753);
nor UO_455 (O_455,N_19761,N_19986);
nand UO_456 (O_456,N_19836,N_19924);
or UO_457 (O_457,N_19690,N_19785);
xor UO_458 (O_458,N_19926,N_19851);
xor UO_459 (O_459,N_19531,N_19622);
nand UO_460 (O_460,N_19908,N_19812);
nand UO_461 (O_461,N_19835,N_19546);
or UO_462 (O_462,N_19690,N_19889);
and UO_463 (O_463,N_19602,N_19801);
xor UO_464 (O_464,N_19763,N_19886);
and UO_465 (O_465,N_19807,N_19818);
or UO_466 (O_466,N_19500,N_19665);
nand UO_467 (O_467,N_19839,N_19956);
xnor UO_468 (O_468,N_19893,N_19837);
and UO_469 (O_469,N_19539,N_19981);
or UO_470 (O_470,N_19697,N_19579);
and UO_471 (O_471,N_19971,N_19741);
or UO_472 (O_472,N_19818,N_19500);
nor UO_473 (O_473,N_19713,N_19995);
xor UO_474 (O_474,N_19930,N_19601);
nor UO_475 (O_475,N_19966,N_19558);
nor UO_476 (O_476,N_19644,N_19961);
xnor UO_477 (O_477,N_19805,N_19533);
xnor UO_478 (O_478,N_19519,N_19714);
nand UO_479 (O_479,N_19910,N_19776);
nand UO_480 (O_480,N_19672,N_19517);
xor UO_481 (O_481,N_19999,N_19585);
xor UO_482 (O_482,N_19847,N_19786);
and UO_483 (O_483,N_19929,N_19771);
xnor UO_484 (O_484,N_19688,N_19819);
and UO_485 (O_485,N_19809,N_19676);
xnor UO_486 (O_486,N_19782,N_19586);
or UO_487 (O_487,N_19620,N_19587);
nand UO_488 (O_488,N_19558,N_19957);
xnor UO_489 (O_489,N_19524,N_19875);
and UO_490 (O_490,N_19997,N_19757);
xnor UO_491 (O_491,N_19822,N_19988);
and UO_492 (O_492,N_19575,N_19951);
nor UO_493 (O_493,N_19835,N_19564);
or UO_494 (O_494,N_19964,N_19561);
and UO_495 (O_495,N_19585,N_19587);
nor UO_496 (O_496,N_19704,N_19514);
and UO_497 (O_497,N_19810,N_19689);
xor UO_498 (O_498,N_19616,N_19851);
nand UO_499 (O_499,N_19767,N_19731);
nand UO_500 (O_500,N_19954,N_19620);
nand UO_501 (O_501,N_19880,N_19650);
or UO_502 (O_502,N_19595,N_19584);
nand UO_503 (O_503,N_19985,N_19645);
or UO_504 (O_504,N_19785,N_19695);
nor UO_505 (O_505,N_19555,N_19809);
and UO_506 (O_506,N_19744,N_19755);
nand UO_507 (O_507,N_19621,N_19509);
nand UO_508 (O_508,N_19748,N_19805);
nand UO_509 (O_509,N_19745,N_19858);
xnor UO_510 (O_510,N_19751,N_19618);
nand UO_511 (O_511,N_19501,N_19815);
xnor UO_512 (O_512,N_19944,N_19509);
nand UO_513 (O_513,N_19710,N_19526);
xor UO_514 (O_514,N_19652,N_19623);
xnor UO_515 (O_515,N_19848,N_19832);
xor UO_516 (O_516,N_19811,N_19542);
or UO_517 (O_517,N_19780,N_19770);
nor UO_518 (O_518,N_19640,N_19768);
nand UO_519 (O_519,N_19667,N_19717);
or UO_520 (O_520,N_19984,N_19526);
nand UO_521 (O_521,N_19692,N_19551);
and UO_522 (O_522,N_19690,N_19630);
nor UO_523 (O_523,N_19950,N_19614);
and UO_524 (O_524,N_19700,N_19688);
or UO_525 (O_525,N_19511,N_19790);
nand UO_526 (O_526,N_19691,N_19586);
or UO_527 (O_527,N_19597,N_19966);
nor UO_528 (O_528,N_19602,N_19554);
nand UO_529 (O_529,N_19531,N_19873);
nand UO_530 (O_530,N_19667,N_19500);
xnor UO_531 (O_531,N_19817,N_19861);
and UO_532 (O_532,N_19925,N_19934);
and UO_533 (O_533,N_19918,N_19852);
nor UO_534 (O_534,N_19531,N_19980);
xnor UO_535 (O_535,N_19852,N_19509);
and UO_536 (O_536,N_19948,N_19813);
nor UO_537 (O_537,N_19934,N_19614);
nand UO_538 (O_538,N_19587,N_19627);
or UO_539 (O_539,N_19513,N_19776);
nand UO_540 (O_540,N_19656,N_19818);
or UO_541 (O_541,N_19806,N_19874);
nand UO_542 (O_542,N_19529,N_19566);
and UO_543 (O_543,N_19663,N_19618);
nor UO_544 (O_544,N_19574,N_19514);
nand UO_545 (O_545,N_19795,N_19954);
nand UO_546 (O_546,N_19860,N_19924);
nand UO_547 (O_547,N_19862,N_19909);
nor UO_548 (O_548,N_19822,N_19520);
nand UO_549 (O_549,N_19964,N_19574);
and UO_550 (O_550,N_19671,N_19653);
nor UO_551 (O_551,N_19530,N_19621);
and UO_552 (O_552,N_19852,N_19839);
and UO_553 (O_553,N_19633,N_19556);
xnor UO_554 (O_554,N_19760,N_19570);
nand UO_555 (O_555,N_19939,N_19734);
or UO_556 (O_556,N_19985,N_19905);
nor UO_557 (O_557,N_19678,N_19624);
or UO_558 (O_558,N_19954,N_19562);
nand UO_559 (O_559,N_19976,N_19737);
nor UO_560 (O_560,N_19940,N_19807);
nor UO_561 (O_561,N_19825,N_19653);
nand UO_562 (O_562,N_19651,N_19699);
or UO_563 (O_563,N_19523,N_19840);
nand UO_564 (O_564,N_19634,N_19725);
or UO_565 (O_565,N_19591,N_19781);
and UO_566 (O_566,N_19656,N_19648);
and UO_567 (O_567,N_19757,N_19634);
nand UO_568 (O_568,N_19655,N_19823);
or UO_569 (O_569,N_19612,N_19690);
nor UO_570 (O_570,N_19751,N_19910);
and UO_571 (O_571,N_19631,N_19678);
xor UO_572 (O_572,N_19517,N_19740);
nand UO_573 (O_573,N_19506,N_19538);
nor UO_574 (O_574,N_19904,N_19959);
nor UO_575 (O_575,N_19959,N_19708);
and UO_576 (O_576,N_19809,N_19794);
or UO_577 (O_577,N_19849,N_19557);
xor UO_578 (O_578,N_19598,N_19919);
nand UO_579 (O_579,N_19606,N_19578);
xnor UO_580 (O_580,N_19518,N_19899);
nor UO_581 (O_581,N_19662,N_19901);
and UO_582 (O_582,N_19729,N_19775);
nor UO_583 (O_583,N_19521,N_19895);
nor UO_584 (O_584,N_19828,N_19718);
xnor UO_585 (O_585,N_19666,N_19739);
nor UO_586 (O_586,N_19664,N_19973);
and UO_587 (O_587,N_19859,N_19854);
nor UO_588 (O_588,N_19640,N_19635);
xor UO_589 (O_589,N_19795,N_19669);
nand UO_590 (O_590,N_19763,N_19541);
nand UO_591 (O_591,N_19820,N_19998);
xor UO_592 (O_592,N_19886,N_19828);
or UO_593 (O_593,N_19836,N_19646);
or UO_594 (O_594,N_19899,N_19942);
nor UO_595 (O_595,N_19659,N_19888);
or UO_596 (O_596,N_19774,N_19645);
nand UO_597 (O_597,N_19936,N_19785);
or UO_598 (O_598,N_19819,N_19681);
or UO_599 (O_599,N_19867,N_19709);
and UO_600 (O_600,N_19746,N_19623);
nor UO_601 (O_601,N_19675,N_19706);
xor UO_602 (O_602,N_19739,N_19578);
xor UO_603 (O_603,N_19623,N_19856);
or UO_604 (O_604,N_19770,N_19671);
or UO_605 (O_605,N_19721,N_19582);
or UO_606 (O_606,N_19624,N_19562);
nand UO_607 (O_607,N_19661,N_19667);
xnor UO_608 (O_608,N_19747,N_19940);
nor UO_609 (O_609,N_19985,N_19624);
nand UO_610 (O_610,N_19565,N_19633);
nor UO_611 (O_611,N_19772,N_19596);
and UO_612 (O_612,N_19552,N_19543);
xnor UO_613 (O_613,N_19689,N_19694);
nor UO_614 (O_614,N_19883,N_19695);
nand UO_615 (O_615,N_19955,N_19749);
nor UO_616 (O_616,N_19594,N_19780);
nor UO_617 (O_617,N_19972,N_19860);
xnor UO_618 (O_618,N_19542,N_19971);
or UO_619 (O_619,N_19997,N_19557);
nand UO_620 (O_620,N_19845,N_19521);
nor UO_621 (O_621,N_19799,N_19626);
nor UO_622 (O_622,N_19528,N_19770);
nand UO_623 (O_623,N_19959,N_19912);
nor UO_624 (O_624,N_19797,N_19652);
nor UO_625 (O_625,N_19537,N_19738);
and UO_626 (O_626,N_19728,N_19886);
or UO_627 (O_627,N_19609,N_19906);
xnor UO_628 (O_628,N_19758,N_19697);
nand UO_629 (O_629,N_19708,N_19663);
nand UO_630 (O_630,N_19841,N_19758);
nor UO_631 (O_631,N_19544,N_19509);
nor UO_632 (O_632,N_19879,N_19992);
nand UO_633 (O_633,N_19662,N_19602);
or UO_634 (O_634,N_19942,N_19847);
and UO_635 (O_635,N_19731,N_19529);
nor UO_636 (O_636,N_19550,N_19893);
or UO_637 (O_637,N_19626,N_19914);
nand UO_638 (O_638,N_19892,N_19850);
or UO_639 (O_639,N_19618,N_19622);
or UO_640 (O_640,N_19627,N_19784);
nand UO_641 (O_641,N_19952,N_19737);
or UO_642 (O_642,N_19973,N_19531);
xor UO_643 (O_643,N_19797,N_19530);
xnor UO_644 (O_644,N_19964,N_19995);
or UO_645 (O_645,N_19700,N_19707);
or UO_646 (O_646,N_19625,N_19860);
and UO_647 (O_647,N_19558,N_19633);
nor UO_648 (O_648,N_19994,N_19755);
and UO_649 (O_649,N_19906,N_19827);
nand UO_650 (O_650,N_19999,N_19800);
and UO_651 (O_651,N_19643,N_19745);
nor UO_652 (O_652,N_19896,N_19914);
and UO_653 (O_653,N_19989,N_19511);
nand UO_654 (O_654,N_19773,N_19725);
nor UO_655 (O_655,N_19702,N_19756);
or UO_656 (O_656,N_19714,N_19612);
nand UO_657 (O_657,N_19538,N_19884);
nand UO_658 (O_658,N_19883,N_19873);
nand UO_659 (O_659,N_19611,N_19861);
nor UO_660 (O_660,N_19841,N_19775);
or UO_661 (O_661,N_19606,N_19692);
or UO_662 (O_662,N_19769,N_19758);
nand UO_663 (O_663,N_19557,N_19936);
and UO_664 (O_664,N_19649,N_19968);
or UO_665 (O_665,N_19795,N_19664);
xnor UO_666 (O_666,N_19584,N_19577);
nand UO_667 (O_667,N_19782,N_19626);
nand UO_668 (O_668,N_19883,N_19839);
nor UO_669 (O_669,N_19734,N_19751);
nor UO_670 (O_670,N_19783,N_19521);
nor UO_671 (O_671,N_19630,N_19760);
xor UO_672 (O_672,N_19582,N_19768);
and UO_673 (O_673,N_19666,N_19986);
and UO_674 (O_674,N_19846,N_19898);
xor UO_675 (O_675,N_19980,N_19773);
and UO_676 (O_676,N_19891,N_19833);
nand UO_677 (O_677,N_19862,N_19567);
nor UO_678 (O_678,N_19619,N_19863);
nor UO_679 (O_679,N_19700,N_19887);
or UO_680 (O_680,N_19873,N_19868);
or UO_681 (O_681,N_19802,N_19996);
nand UO_682 (O_682,N_19901,N_19603);
nor UO_683 (O_683,N_19611,N_19880);
xnor UO_684 (O_684,N_19897,N_19813);
and UO_685 (O_685,N_19572,N_19512);
nand UO_686 (O_686,N_19522,N_19869);
nand UO_687 (O_687,N_19731,N_19547);
nand UO_688 (O_688,N_19945,N_19609);
xnor UO_689 (O_689,N_19760,N_19858);
or UO_690 (O_690,N_19621,N_19805);
xnor UO_691 (O_691,N_19655,N_19826);
xor UO_692 (O_692,N_19908,N_19777);
xnor UO_693 (O_693,N_19905,N_19931);
nor UO_694 (O_694,N_19500,N_19942);
or UO_695 (O_695,N_19979,N_19560);
nor UO_696 (O_696,N_19756,N_19639);
and UO_697 (O_697,N_19572,N_19754);
xor UO_698 (O_698,N_19656,N_19536);
xor UO_699 (O_699,N_19665,N_19922);
xor UO_700 (O_700,N_19875,N_19637);
or UO_701 (O_701,N_19965,N_19997);
or UO_702 (O_702,N_19695,N_19644);
nor UO_703 (O_703,N_19582,N_19598);
nand UO_704 (O_704,N_19678,N_19909);
or UO_705 (O_705,N_19627,N_19798);
nand UO_706 (O_706,N_19690,N_19649);
or UO_707 (O_707,N_19595,N_19639);
xnor UO_708 (O_708,N_19790,N_19894);
and UO_709 (O_709,N_19912,N_19918);
and UO_710 (O_710,N_19956,N_19632);
xor UO_711 (O_711,N_19743,N_19961);
nor UO_712 (O_712,N_19636,N_19902);
nor UO_713 (O_713,N_19889,N_19700);
or UO_714 (O_714,N_19668,N_19716);
nand UO_715 (O_715,N_19809,N_19743);
and UO_716 (O_716,N_19874,N_19552);
or UO_717 (O_717,N_19677,N_19771);
and UO_718 (O_718,N_19724,N_19643);
xnor UO_719 (O_719,N_19912,N_19634);
or UO_720 (O_720,N_19883,N_19887);
or UO_721 (O_721,N_19992,N_19768);
xnor UO_722 (O_722,N_19543,N_19567);
xor UO_723 (O_723,N_19831,N_19879);
and UO_724 (O_724,N_19592,N_19829);
nor UO_725 (O_725,N_19941,N_19589);
xor UO_726 (O_726,N_19603,N_19617);
nor UO_727 (O_727,N_19933,N_19760);
nor UO_728 (O_728,N_19633,N_19853);
xnor UO_729 (O_729,N_19884,N_19516);
nor UO_730 (O_730,N_19834,N_19515);
nand UO_731 (O_731,N_19593,N_19822);
and UO_732 (O_732,N_19646,N_19579);
and UO_733 (O_733,N_19926,N_19975);
nor UO_734 (O_734,N_19690,N_19913);
or UO_735 (O_735,N_19835,N_19727);
xor UO_736 (O_736,N_19689,N_19893);
xor UO_737 (O_737,N_19732,N_19965);
xor UO_738 (O_738,N_19672,N_19954);
nor UO_739 (O_739,N_19946,N_19886);
nor UO_740 (O_740,N_19909,N_19614);
and UO_741 (O_741,N_19973,N_19819);
and UO_742 (O_742,N_19680,N_19844);
and UO_743 (O_743,N_19645,N_19847);
xnor UO_744 (O_744,N_19863,N_19994);
or UO_745 (O_745,N_19545,N_19759);
nor UO_746 (O_746,N_19965,N_19686);
and UO_747 (O_747,N_19908,N_19768);
nand UO_748 (O_748,N_19906,N_19588);
nor UO_749 (O_749,N_19800,N_19648);
and UO_750 (O_750,N_19667,N_19868);
nand UO_751 (O_751,N_19842,N_19540);
nor UO_752 (O_752,N_19611,N_19850);
and UO_753 (O_753,N_19570,N_19700);
xor UO_754 (O_754,N_19860,N_19671);
nand UO_755 (O_755,N_19700,N_19710);
nand UO_756 (O_756,N_19592,N_19573);
xnor UO_757 (O_757,N_19638,N_19525);
xnor UO_758 (O_758,N_19650,N_19783);
nand UO_759 (O_759,N_19814,N_19714);
or UO_760 (O_760,N_19915,N_19528);
xnor UO_761 (O_761,N_19852,N_19798);
and UO_762 (O_762,N_19552,N_19584);
or UO_763 (O_763,N_19959,N_19734);
xor UO_764 (O_764,N_19764,N_19577);
nand UO_765 (O_765,N_19941,N_19949);
or UO_766 (O_766,N_19734,N_19740);
xor UO_767 (O_767,N_19732,N_19889);
xnor UO_768 (O_768,N_19774,N_19925);
xor UO_769 (O_769,N_19635,N_19751);
nor UO_770 (O_770,N_19836,N_19644);
and UO_771 (O_771,N_19543,N_19661);
or UO_772 (O_772,N_19581,N_19706);
and UO_773 (O_773,N_19665,N_19824);
nor UO_774 (O_774,N_19714,N_19856);
xor UO_775 (O_775,N_19679,N_19579);
xnor UO_776 (O_776,N_19959,N_19916);
nand UO_777 (O_777,N_19832,N_19921);
xnor UO_778 (O_778,N_19980,N_19915);
nor UO_779 (O_779,N_19957,N_19838);
nand UO_780 (O_780,N_19760,N_19636);
xor UO_781 (O_781,N_19643,N_19942);
xor UO_782 (O_782,N_19927,N_19975);
nand UO_783 (O_783,N_19996,N_19853);
or UO_784 (O_784,N_19561,N_19944);
xor UO_785 (O_785,N_19651,N_19742);
nor UO_786 (O_786,N_19890,N_19878);
xnor UO_787 (O_787,N_19904,N_19578);
and UO_788 (O_788,N_19563,N_19579);
and UO_789 (O_789,N_19585,N_19562);
and UO_790 (O_790,N_19709,N_19972);
or UO_791 (O_791,N_19558,N_19963);
xor UO_792 (O_792,N_19965,N_19568);
nor UO_793 (O_793,N_19562,N_19630);
and UO_794 (O_794,N_19633,N_19531);
nor UO_795 (O_795,N_19511,N_19974);
nand UO_796 (O_796,N_19631,N_19518);
or UO_797 (O_797,N_19693,N_19741);
and UO_798 (O_798,N_19697,N_19597);
xnor UO_799 (O_799,N_19614,N_19894);
nand UO_800 (O_800,N_19621,N_19684);
and UO_801 (O_801,N_19864,N_19669);
nor UO_802 (O_802,N_19608,N_19865);
xor UO_803 (O_803,N_19738,N_19776);
nand UO_804 (O_804,N_19925,N_19821);
and UO_805 (O_805,N_19540,N_19657);
nor UO_806 (O_806,N_19567,N_19989);
nor UO_807 (O_807,N_19582,N_19938);
nand UO_808 (O_808,N_19768,N_19922);
nor UO_809 (O_809,N_19793,N_19731);
and UO_810 (O_810,N_19530,N_19829);
and UO_811 (O_811,N_19694,N_19793);
nand UO_812 (O_812,N_19636,N_19590);
and UO_813 (O_813,N_19537,N_19982);
or UO_814 (O_814,N_19846,N_19756);
nor UO_815 (O_815,N_19625,N_19820);
and UO_816 (O_816,N_19932,N_19891);
nand UO_817 (O_817,N_19969,N_19500);
nand UO_818 (O_818,N_19736,N_19818);
nor UO_819 (O_819,N_19661,N_19917);
nand UO_820 (O_820,N_19642,N_19623);
nand UO_821 (O_821,N_19913,N_19891);
nor UO_822 (O_822,N_19788,N_19660);
xor UO_823 (O_823,N_19980,N_19500);
and UO_824 (O_824,N_19892,N_19934);
xor UO_825 (O_825,N_19631,N_19929);
nand UO_826 (O_826,N_19676,N_19716);
nor UO_827 (O_827,N_19528,N_19843);
and UO_828 (O_828,N_19661,N_19698);
or UO_829 (O_829,N_19599,N_19676);
xnor UO_830 (O_830,N_19908,N_19973);
nand UO_831 (O_831,N_19934,N_19947);
or UO_832 (O_832,N_19805,N_19791);
xor UO_833 (O_833,N_19920,N_19900);
xor UO_834 (O_834,N_19627,N_19517);
and UO_835 (O_835,N_19743,N_19656);
xor UO_836 (O_836,N_19678,N_19823);
nand UO_837 (O_837,N_19998,N_19934);
nand UO_838 (O_838,N_19863,N_19705);
nor UO_839 (O_839,N_19817,N_19849);
and UO_840 (O_840,N_19657,N_19686);
xnor UO_841 (O_841,N_19730,N_19975);
nor UO_842 (O_842,N_19822,N_19901);
or UO_843 (O_843,N_19755,N_19958);
nand UO_844 (O_844,N_19578,N_19858);
and UO_845 (O_845,N_19849,N_19907);
or UO_846 (O_846,N_19600,N_19968);
xnor UO_847 (O_847,N_19836,N_19612);
nor UO_848 (O_848,N_19921,N_19513);
and UO_849 (O_849,N_19885,N_19701);
and UO_850 (O_850,N_19726,N_19907);
xnor UO_851 (O_851,N_19511,N_19679);
nand UO_852 (O_852,N_19718,N_19547);
nand UO_853 (O_853,N_19525,N_19718);
xnor UO_854 (O_854,N_19871,N_19815);
xnor UO_855 (O_855,N_19928,N_19757);
nand UO_856 (O_856,N_19925,N_19592);
or UO_857 (O_857,N_19932,N_19707);
nor UO_858 (O_858,N_19914,N_19650);
nand UO_859 (O_859,N_19665,N_19899);
and UO_860 (O_860,N_19887,N_19625);
nand UO_861 (O_861,N_19821,N_19695);
and UO_862 (O_862,N_19516,N_19741);
or UO_863 (O_863,N_19534,N_19645);
xnor UO_864 (O_864,N_19584,N_19926);
nor UO_865 (O_865,N_19960,N_19992);
or UO_866 (O_866,N_19971,N_19942);
xnor UO_867 (O_867,N_19812,N_19724);
xnor UO_868 (O_868,N_19581,N_19966);
or UO_869 (O_869,N_19957,N_19563);
and UO_870 (O_870,N_19547,N_19874);
or UO_871 (O_871,N_19556,N_19564);
and UO_872 (O_872,N_19801,N_19982);
and UO_873 (O_873,N_19933,N_19571);
nor UO_874 (O_874,N_19842,N_19735);
nand UO_875 (O_875,N_19781,N_19635);
xor UO_876 (O_876,N_19853,N_19614);
or UO_877 (O_877,N_19991,N_19899);
xnor UO_878 (O_878,N_19855,N_19606);
nor UO_879 (O_879,N_19804,N_19564);
or UO_880 (O_880,N_19780,N_19840);
or UO_881 (O_881,N_19900,N_19591);
or UO_882 (O_882,N_19832,N_19529);
nand UO_883 (O_883,N_19607,N_19892);
nor UO_884 (O_884,N_19508,N_19781);
and UO_885 (O_885,N_19707,N_19672);
nor UO_886 (O_886,N_19690,N_19936);
or UO_887 (O_887,N_19517,N_19945);
xor UO_888 (O_888,N_19514,N_19884);
xor UO_889 (O_889,N_19524,N_19724);
xnor UO_890 (O_890,N_19956,N_19796);
and UO_891 (O_891,N_19838,N_19700);
or UO_892 (O_892,N_19710,N_19567);
or UO_893 (O_893,N_19945,N_19715);
or UO_894 (O_894,N_19747,N_19699);
xor UO_895 (O_895,N_19954,N_19956);
and UO_896 (O_896,N_19515,N_19913);
nor UO_897 (O_897,N_19722,N_19812);
nand UO_898 (O_898,N_19644,N_19894);
and UO_899 (O_899,N_19862,N_19765);
and UO_900 (O_900,N_19952,N_19667);
and UO_901 (O_901,N_19698,N_19675);
or UO_902 (O_902,N_19890,N_19998);
xor UO_903 (O_903,N_19502,N_19825);
and UO_904 (O_904,N_19932,N_19808);
and UO_905 (O_905,N_19506,N_19522);
nor UO_906 (O_906,N_19513,N_19878);
or UO_907 (O_907,N_19649,N_19892);
xnor UO_908 (O_908,N_19554,N_19738);
nand UO_909 (O_909,N_19803,N_19885);
nor UO_910 (O_910,N_19666,N_19811);
nand UO_911 (O_911,N_19709,N_19901);
nor UO_912 (O_912,N_19893,N_19759);
nor UO_913 (O_913,N_19700,N_19522);
and UO_914 (O_914,N_19891,N_19592);
or UO_915 (O_915,N_19894,N_19870);
xor UO_916 (O_916,N_19631,N_19745);
xnor UO_917 (O_917,N_19750,N_19678);
nand UO_918 (O_918,N_19665,N_19759);
xnor UO_919 (O_919,N_19562,N_19516);
and UO_920 (O_920,N_19683,N_19644);
and UO_921 (O_921,N_19643,N_19731);
nor UO_922 (O_922,N_19937,N_19681);
nand UO_923 (O_923,N_19688,N_19984);
xor UO_924 (O_924,N_19707,N_19517);
nor UO_925 (O_925,N_19685,N_19854);
nand UO_926 (O_926,N_19758,N_19646);
nor UO_927 (O_927,N_19793,N_19633);
or UO_928 (O_928,N_19651,N_19503);
nor UO_929 (O_929,N_19723,N_19805);
nor UO_930 (O_930,N_19928,N_19561);
nand UO_931 (O_931,N_19942,N_19734);
and UO_932 (O_932,N_19814,N_19720);
and UO_933 (O_933,N_19679,N_19867);
nor UO_934 (O_934,N_19995,N_19871);
or UO_935 (O_935,N_19505,N_19537);
nand UO_936 (O_936,N_19558,N_19761);
and UO_937 (O_937,N_19985,N_19806);
nand UO_938 (O_938,N_19828,N_19772);
xnor UO_939 (O_939,N_19786,N_19546);
and UO_940 (O_940,N_19717,N_19896);
and UO_941 (O_941,N_19799,N_19970);
and UO_942 (O_942,N_19999,N_19602);
xor UO_943 (O_943,N_19847,N_19821);
nor UO_944 (O_944,N_19777,N_19819);
xor UO_945 (O_945,N_19535,N_19915);
and UO_946 (O_946,N_19579,N_19647);
or UO_947 (O_947,N_19722,N_19630);
xnor UO_948 (O_948,N_19770,N_19889);
and UO_949 (O_949,N_19518,N_19895);
and UO_950 (O_950,N_19631,N_19977);
nand UO_951 (O_951,N_19837,N_19834);
nand UO_952 (O_952,N_19842,N_19604);
nor UO_953 (O_953,N_19668,N_19811);
and UO_954 (O_954,N_19638,N_19505);
nand UO_955 (O_955,N_19547,N_19593);
nor UO_956 (O_956,N_19628,N_19536);
or UO_957 (O_957,N_19731,N_19947);
nand UO_958 (O_958,N_19944,N_19841);
and UO_959 (O_959,N_19570,N_19930);
nor UO_960 (O_960,N_19990,N_19543);
nor UO_961 (O_961,N_19625,N_19506);
nor UO_962 (O_962,N_19704,N_19646);
and UO_963 (O_963,N_19843,N_19778);
nor UO_964 (O_964,N_19666,N_19775);
xor UO_965 (O_965,N_19776,N_19658);
xnor UO_966 (O_966,N_19605,N_19878);
xnor UO_967 (O_967,N_19969,N_19917);
nand UO_968 (O_968,N_19812,N_19646);
nand UO_969 (O_969,N_19883,N_19809);
xnor UO_970 (O_970,N_19801,N_19963);
and UO_971 (O_971,N_19613,N_19794);
nor UO_972 (O_972,N_19545,N_19820);
or UO_973 (O_973,N_19596,N_19851);
and UO_974 (O_974,N_19882,N_19563);
nand UO_975 (O_975,N_19814,N_19961);
xor UO_976 (O_976,N_19980,N_19559);
nand UO_977 (O_977,N_19512,N_19942);
xnor UO_978 (O_978,N_19643,N_19646);
xnor UO_979 (O_979,N_19568,N_19799);
or UO_980 (O_980,N_19901,N_19521);
nand UO_981 (O_981,N_19809,N_19644);
nand UO_982 (O_982,N_19624,N_19737);
xnor UO_983 (O_983,N_19631,N_19876);
and UO_984 (O_984,N_19631,N_19969);
nand UO_985 (O_985,N_19776,N_19876);
nor UO_986 (O_986,N_19561,N_19708);
xor UO_987 (O_987,N_19502,N_19653);
or UO_988 (O_988,N_19976,N_19927);
nand UO_989 (O_989,N_19919,N_19975);
or UO_990 (O_990,N_19524,N_19692);
and UO_991 (O_991,N_19705,N_19971);
xnor UO_992 (O_992,N_19784,N_19993);
nand UO_993 (O_993,N_19917,N_19735);
and UO_994 (O_994,N_19955,N_19670);
xor UO_995 (O_995,N_19672,N_19690);
nor UO_996 (O_996,N_19718,N_19689);
xnor UO_997 (O_997,N_19918,N_19994);
or UO_998 (O_998,N_19861,N_19706);
nor UO_999 (O_999,N_19782,N_19628);
nand UO_1000 (O_1000,N_19588,N_19842);
nand UO_1001 (O_1001,N_19796,N_19989);
and UO_1002 (O_1002,N_19636,N_19873);
xnor UO_1003 (O_1003,N_19546,N_19872);
nor UO_1004 (O_1004,N_19683,N_19950);
nor UO_1005 (O_1005,N_19989,N_19620);
and UO_1006 (O_1006,N_19514,N_19655);
xnor UO_1007 (O_1007,N_19648,N_19704);
nand UO_1008 (O_1008,N_19655,N_19956);
or UO_1009 (O_1009,N_19700,N_19581);
and UO_1010 (O_1010,N_19706,N_19849);
nand UO_1011 (O_1011,N_19573,N_19806);
nor UO_1012 (O_1012,N_19737,N_19672);
nand UO_1013 (O_1013,N_19991,N_19826);
xnor UO_1014 (O_1014,N_19684,N_19789);
or UO_1015 (O_1015,N_19783,N_19861);
xnor UO_1016 (O_1016,N_19812,N_19994);
and UO_1017 (O_1017,N_19716,N_19504);
or UO_1018 (O_1018,N_19542,N_19713);
or UO_1019 (O_1019,N_19691,N_19500);
or UO_1020 (O_1020,N_19797,N_19897);
nor UO_1021 (O_1021,N_19695,N_19895);
xnor UO_1022 (O_1022,N_19565,N_19905);
nor UO_1023 (O_1023,N_19753,N_19996);
nor UO_1024 (O_1024,N_19642,N_19743);
nor UO_1025 (O_1025,N_19506,N_19950);
nand UO_1026 (O_1026,N_19735,N_19684);
nor UO_1027 (O_1027,N_19592,N_19886);
and UO_1028 (O_1028,N_19621,N_19824);
or UO_1029 (O_1029,N_19711,N_19660);
xnor UO_1030 (O_1030,N_19541,N_19906);
nor UO_1031 (O_1031,N_19761,N_19788);
or UO_1032 (O_1032,N_19926,N_19886);
nor UO_1033 (O_1033,N_19729,N_19936);
and UO_1034 (O_1034,N_19998,N_19520);
xnor UO_1035 (O_1035,N_19548,N_19631);
nand UO_1036 (O_1036,N_19652,N_19639);
and UO_1037 (O_1037,N_19682,N_19946);
or UO_1038 (O_1038,N_19891,N_19923);
nor UO_1039 (O_1039,N_19944,N_19758);
nor UO_1040 (O_1040,N_19781,N_19985);
nand UO_1041 (O_1041,N_19625,N_19524);
or UO_1042 (O_1042,N_19564,N_19969);
nor UO_1043 (O_1043,N_19825,N_19708);
and UO_1044 (O_1044,N_19808,N_19652);
xor UO_1045 (O_1045,N_19628,N_19729);
or UO_1046 (O_1046,N_19738,N_19712);
nand UO_1047 (O_1047,N_19877,N_19867);
or UO_1048 (O_1048,N_19553,N_19759);
xnor UO_1049 (O_1049,N_19619,N_19775);
xnor UO_1050 (O_1050,N_19955,N_19728);
and UO_1051 (O_1051,N_19750,N_19761);
nor UO_1052 (O_1052,N_19629,N_19671);
and UO_1053 (O_1053,N_19810,N_19608);
and UO_1054 (O_1054,N_19537,N_19555);
and UO_1055 (O_1055,N_19567,N_19969);
and UO_1056 (O_1056,N_19529,N_19503);
nor UO_1057 (O_1057,N_19700,N_19593);
nand UO_1058 (O_1058,N_19852,N_19776);
and UO_1059 (O_1059,N_19775,N_19996);
xor UO_1060 (O_1060,N_19526,N_19908);
and UO_1061 (O_1061,N_19839,N_19662);
nand UO_1062 (O_1062,N_19868,N_19645);
nand UO_1063 (O_1063,N_19946,N_19881);
nor UO_1064 (O_1064,N_19515,N_19541);
xnor UO_1065 (O_1065,N_19809,N_19698);
or UO_1066 (O_1066,N_19776,N_19859);
and UO_1067 (O_1067,N_19659,N_19764);
and UO_1068 (O_1068,N_19851,N_19636);
nand UO_1069 (O_1069,N_19599,N_19538);
nor UO_1070 (O_1070,N_19824,N_19746);
and UO_1071 (O_1071,N_19953,N_19754);
xnor UO_1072 (O_1072,N_19646,N_19792);
xor UO_1073 (O_1073,N_19660,N_19935);
and UO_1074 (O_1074,N_19704,N_19744);
and UO_1075 (O_1075,N_19666,N_19784);
xnor UO_1076 (O_1076,N_19786,N_19658);
nor UO_1077 (O_1077,N_19525,N_19600);
and UO_1078 (O_1078,N_19717,N_19577);
or UO_1079 (O_1079,N_19511,N_19746);
or UO_1080 (O_1080,N_19749,N_19827);
xnor UO_1081 (O_1081,N_19643,N_19962);
and UO_1082 (O_1082,N_19979,N_19882);
xor UO_1083 (O_1083,N_19610,N_19888);
or UO_1084 (O_1084,N_19547,N_19790);
xor UO_1085 (O_1085,N_19521,N_19941);
nor UO_1086 (O_1086,N_19573,N_19520);
and UO_1087 (O_1087,N_19672,N_19790);
or UO_1088 (O_1088,N_19518,N_19559);
and UO_1089 (O_1089,N_19811,N_19707);
xor UO_1090 (O_1090,N_19545,N_19535);
nor UO_1091 (O_1091,N_19933,N_19722);
nor UO_1092 (O_1092,N_19559,N_19514);
nor UO_1093 (O_1093,N_19960,N_19764);
and UO_1094 (O_1094,N_19807,N_19583);
and UO_1095 (O_1095,N_19933,N_19630);
and UO_1096 (O_1096,N_19879,N_19670);
and UO_1097 (O_1097,N_19838,N_19722);
nand UO_1098 (O_1098,N_19646,N_19930);
and UO_1099 (O_1099,N_19660,N_19916);
xnor UO_1100 (O_1100,N_19554,N_19859);
or UO_1101 (O_1101,N_19560,N_19819);
or UO_1102 (O_1102,N_19934,N_19783);
nand UO_1103 (O_1103,N_19617,N_19948);
nor UO_1104 (O_1104,N_19955,N_19938);
nand UO_1105 (O_1105,N_19774,N_19667);
or UO_1106 (O_1106,N_19799,N_19897);
xnor UO_1107 (O_1107,N_19678,N_19633);
nand UO_1108 (O_1108,N_19703,N_19528);
nand UO_1109 (O_1109,N_19689,N_19517);
xor UO_1110 (O_1110,N_19640,N_19505);
nor UO_1111 (O_1111,N_19811,N_19572);
and UO_1112 (O_1112,N_19940,N_19634);
and UO_1113 (O_1113,N_19960,N_19615);
and UO_1114 (O_1114,N_19718,N_19635);
xnor UO_1115 (O_1115,N_19591,N_19693);
and UO_1116 (O_1116,N_19566,N_19801);
nor UO_1117 (O_1117,N_19759,N_19592);
nor UO_1118 (O_1118,N_19658,N_19876);
nand UO_1119 (O_1119,N_19593,N_19763);
nor UO_1120 (O_1120,N_19769,N_19667);
and UO_1121 (O_1121,N_19972,N_19837);
nand UO_1122 (O_1122,N_19810,N_19650);
xnor UO_1123 (O_1123,N_19650,N_19702);
xnor UO_1124 (O_1124,N_19804,N_19877);
nand UO_1125 (O_1125,N_19631,N_19895);
nand UO_1126 (O_1126,N_19970,N_19694);
xnor UO_1127 (O_1127,N_19567,N_19943);
nand UO_1128 (O_1128,N_19597,N_19810);
nand UO_1129 (O_1129,N_19762,N_19845);
nor UO_1130 (O_1130,N_19904,N_19869);
or UO_1131 (O_1131,N_19880,N_19599);
and UO_1132 (O_1132,N_19655,N_19934);
or UO_1133 (O_1133,N_19596,N_19657);
or UO_1134 (O_1134,N_19855,N_19746);
and UO_1135 (O_1135,N_19603,N_19964);
xor UO_1136 (O_1136,N_19560,N_19568);
nand UO_1137 (O_1137,N_19696,N_19889);
or UO_1138 (O_1138,N_19759,N_19841);
or UO_1139 (O_1139,N_19758,N_19515);
or UO_1140 (O_1140,N_19855,N_19727);
nor UO_1141 (O_1141,N_19575,N_19986);
or UO_1142 (O_1142,N_19724,N_19749);
xnor UO_1143 (O_1143,N_19855,N_19642);
xor UO_1144 (O_1144,N_19857,N_19818);
nand UO_1145 (O_1145,N_19887,N_19628);
nand UO_1146 (O_1146,N_19575,N_19908);
and UO_1147 (O_1147,N_19954,N_19512);
or UO_1148 (O_1148,N_19949,N_19709);
nor UO_1149 (O_1149,N_19544,N_19696);
or UO_1150 (O_1150,N_19753,N_19560);
or UO_1151 (O_1151,N_19628,N_19502);
xnor UO_1152 (O_1152,N_19670,N_19995);
or UO_1153 (O_1153,N_19922,N_19829);
nand UO_1154 (O_1154,N_19540,N_19619);
xnor UO_1155 (O_1155,N_19963,N_19705);
nand UO_1156 (O_1156,N_19513,N_19907);
and UO_1157 (O_1157,N_19842,N_19786);
nand UO_1158 (O_1158,N_19689,N_19977);
or UO_1159 (O_1159,N_19736,N_19763);
nand UO_1160 (O_1160,N_19673,N_19651);
or UO_1161 (O_1161,N_19663,N_19701);
or UO_1162 (O_1162,N_19754,N_19926);
nand UO_1163 (O_1163,N_19791,N_19794);
and UO_1164 (O_1164,N_19965,N_19861);
xnor UO_1165 (O_1165,N_19898,N_19928);
and UO_1166 (O_1166,N_19661,N_19596);
and UO_1167 (O_1167,N_19729,N_19951);
nand UO_1168 (O_1168,N_19707,N_19941);
or UO_1169 (O_1169,N_19735,N_19816);
xnor UO_1170 (O_1170,N_19658,N_19696);
and UO_1171 (O_1171,N_19964,N_19793);
xnor UO_1172 (O_1172,N_19656,N_19541);
nand UO_1173 (O_1173,N_19645,N_19844);
nand UO_1174 (O_1174,N_19679,N_19861);
nand UO_1175 (O_1175,N_19826,N_19596);
nor UO_1176 (O_1176,N_19571,N_19912);
and UO_1177 (O_1177,N_19985,N_19958);
and UO_1178 (O_1178,N_19591,N_19750);
nand UO_1179 (O_1179,N_19905,N_19926);
and UO_1180 (O_1180,N_19742,N_19574);
xnor UO_1181 (O_1181,N_19906,N_19775);
xnor UO_1182 (O_1182,N_19930,N_19871);
xnor UO_1183 (O_1183,N_19867,N_19732);
and UO_1184 (O_1184,N_19944,N_19836);
or UO_1185 (O_1185,N_19860,N_19799);
and UO_1186 (O_1186,N_19618,N_19607);
nor UO_1187 (O_1187,N_19602,N_19731);
nor UO_1188 (O_1188,N_19598,N_19990);
or UO_1189 (O_1189,N_19728,N_19684);
xor UO_1190 (O_1190,N_19792,N_19639);
nand UO_1191 (O_1191,N_19631,N_19915);
nor UO_1192 (O_1192,N_19641,N_19716);
nand UO_1193 (O_1193,N_19891,N_19679);
xor UO_1194 (O_1194,N_19864,N_19842);
or UO_1195 (O_1195,N_19973,N_19631);
nand UO_1196 (O_1196,N_19854,N_19566);
and UO_1197 (O_1197,N_19583,N_19679);
nand UO_1198 (O_1198,N_19675,N_19511);
and UO_1199 (O_1199,N_19817,N_19546);
nor UO_1200 (O_1200,N_19611,N_19944);
and UO_1201 (O_1201,N_19508,N_19787);
or UO_1202 (O_1202,N_19667,N_19541);
xor UO_1203 (O_1203,N_19751,N_19888);
nand UO_1204 (O_1204,N_19608,N_19812);
or UO_1205 (O_1205,N_19843,N_19771);
nand UO_1206 (O_1206,N_19731,N_19672);
and UO_1207 (O_1207,N_19810,N_19637);
and UO_1208 (O_1208,N_19579,N_19975);
or UO_1209 (O_1209,N_19661,N_19892);
or UO_1210 (O_1210,N_19886,N_19552);
xnor UO_1211 (O_1211,N_19606,N_19776);
xor UO_1212 (O_1212,N_19689,N_19903);
xor UO_1213 (O_1213,N_19854,N_19699);
nand UO_1214 (O_1214,N_19612,N_19592);
and UO_1215 (O_1215,N_19556,N_19680);
or UO_1216 (O_1216,N_19528,N_19513);
nor UO_1217 (O_1217,N_19663,N_19653);
and UO_1218 (O_1218,N_19500,N_19603);
nor UO_1219 (O_1219,N_19921,N_19846);
nor UO_1220 (O_1220,N_19915,N_19519);
and UO_1221 (O_1221,N_19934,N_19569);
nor UO_1222 (O_1222,N_19704,N_19627);
xor UO_1223 (O_1223,N_19556,N_19565);
nor UO_1224 (O_1224,N_19781,N_19527);
nand UO_1225 (O_1225,N_19772,N_19839);
or UO_1226 (O_1226,N_19773,N_19651);
xor UO_1227 (O_1227,N_19583,N_19993);
nor UO_1228 (O_1228,N_19810,N_19683);
or UO_1229 (O_1229,N_19652,N_19536);
nand UO_1230 (O_1230,N_19833,N_19653);
and UO_1231 (O_1231,N_19994,N_19819);
nor UO_1232 (O_1232,N_19822,N_19553);
nand UO_1233 (O_1233,N_19873,N_19893);
and UO_1234 (O_1234,N_19944,N_19803);
and UO_1235 (O_1235,N_19974,N_19656);
nor UO_1236 (O_1236,N_19962,N_19528);
or UO_1237 (O_1237,N_19938,N_19542);
xor UO_1238 (O_1238,N_19526,N_19951);
and UO_1239 (O_1239,N_19603,N_19567);
nor UO_1240 (O_1240,N_19740,N_19795);
nor UO_1241 (O_1241,N_19856,N_19791);
or UO_1242 (O_1242,N_19763,N_19808);
xnor UO_1243 (O_1243,N_19527,N_19535);
and UO_1244 (O_1244,N_19591,N_19740);
or UO_1245 (O_1245,N_19745,N_19919);
and UO_1246 (O_1246,N_19676,N_19808);
and UO_1247 (O_1247,N_19667,N_19506);
xor UO_1248 (O_1248,N_19710,N_19642);
nor UO_1249 (O_1249,N_19938,N_19968);
or UO_1250 (O_1250,N_19570,N_19852);
nor UO_1251 (O_1251,N_19889,N_19653);
nand UO_1252 (O_1252,N_19981,N_19536);
xnor UO_1253 (O_1253,N_19623,N_19947);
nand UO_1254 (O_1254,N_19504,N_19879);
nand UO_1255 (O_1255,N_19622,N_19528);
xnor UO_1256 (O_1256,N_19985,N_19815);
and UO_1257 (O_1257,N_19686,N_19736);
or UO_1258 (O_1258,N_19920,N_19878);
xnor UO_1259 (O_1259,N_19841,N_19991);
and UO_1260 (O_1260,N_19693,N_19744);
xor UO_1261 (O_1261,N_19871,N_19808);
and UO_1262 (O_1262,N_19605,N_19980);
nor UO_1263 (O_1263,N_19670,N_19551);
nand UO_1264 (O_1264,N_19862,N_19965);
nand UO_1265 (O_1265,N_19660,N_19833);
or UO_1266 (O_1266,N_19623,N_19569);
nor UO_1267 (O_1267,N_19572,N_19792);
or UO_1268 (O_1268,N_19880,N_19915);
and UO_1269 (O_1269,N_19755,N_19751);
and UO_1270 (O_1270,N_19542,N_19894);
nand UO_1271 (O_1271,N_19605,N_19507);
nor UO_1272 (O_1272,N_19932,N_19580);
nand UO_1273 (O_1273,N_19831,N_19966);
nor UO_1274 (O_1274,N_19913,N_19753);
xor UO_1275 (O_1275,N_19597,N_19767);
nor UO_1276 (O_1276,N_19771,N_19879);
or UO_1277 (O_1277,N_19790,N_19621);
or UO_1278 (O_1278,N_19715,N_19784);
nor UO_1279 (O_1279,N_19902,N_19642);
or UO_1280 (O_1280,N_19969,N_19762);
nand UO_1281 (O_1281,N_19780,N_19567);
nor UO_1282 (O_1282,N_19832,N_19875);
or UO_1283 (O_1283,N_19577,N_19672);
xnor UO_1284 (O_1284,N_19542,N_19968);
xor UO_1285 (O_1285,N_19693,N_19768);
nand UO_1286 (O_1286,N_19988,N_19975);
and UO_1287 (O_1287,N_19604,N_19654);
or UO_1288 (O_1288,N_19626,N_19790);
or UO_1289 (O_1289,N_19689,N_19637);
and UO_1290 (O_1290,N_19894,N_19881);
nand UO_1291 (O_1291,N_19757,N_19854);
or UO_1292 (O_1292,N_19898,N_19593);
nand UO_1293 (O_1293,N_19591,N_19801);
nand UO_1294 (O_1294,N_19619,N_19552);
or UO_1295 (O_1295,N_19802,N_19553);
nand UO_1296 (O_1296,N_19866,N_19884);
or UO_1297 (O_1297,N_19948,N_19879);
or UO_1298 (O_1298,N_19514,N_19609);
xor UO_1299 (O_1299,N_19713,N_19777);
nand UO_1300 (O_1300,N_19773,N_19974);
xnor UO_1301 (O_1301,N_19775,N_19709);
nand UO_1302 (O_1302,N_19634,N_19746);
and UO_1303 (O_1303,N_19944,N_19871);
xor UO_1304 (O_1304,N_19697,N_19812);
or UO_1305 (O_1305,N_19517,N_19954);
xor UO_1306 (O_1306,N_19500,N_19971);
xor UO_1307 (O_1307,N_19521,N_19988);
nand UO_1308 (O_1308,N_19945,N_19737);
or UO_1309 (O_1309,N_19869,N_19960);
nor UO_1310 (O_1310,N_19855,N_19624);
or UO_1311 (O_1311,N_19879,N_19843);
nand UO_1312 (O_1312,N_19929,N_19765);
nor UO_1313 (O_1313,N_19939,N_19768);
xnor UO_1314 (O_1314,N_19913,N_19751);
or UO_1315 (O_1315,N_19750,N_19920);
xnor UO_1316 (O_1316,N_19961,N_19937);
xor UO_1317 (O_1317,N_19626,N_19735);
and UO_1318 (O_1318,N_19845,N_19704);
nand UO_1319 (O_1319,N_19544,N_19720);
nand UO_1320 (O_1320,N_19798,N_19876);
and UO_1321 (O_1321,N_19954,N_19555);
and UO_1322 (O_1322,N_19616,N_19624);
nor UO_1323 (O_1323,N_19782,N_19849);
and UO_1324 (O_1324,N_19706,N_19720);
xnor UO_1325 (O_1325,N_19684,N_19727);
or UO_1326 (O_1326,N_19662,N_19735);
xor UO_1327 (O_1327,N_19948,N_19599);
xor UO_1328 (O_1328,N_19612,N_19711);
or UO_1329 (O_1329,N_19520,N_19803);
nand UO_1330 (O_1330,N_19656,N_19575);
nor UO_1331 (O_1331,N_19690,N_19958);
or UO_1332 (O_1332,N_19654,N_19708);
or UO_1333 (O_1333,N_19574,N_19743);
nor UO_1334 (O_1334,N_19545,N_19979);
nor UO_1335 (O_1335,N_19773,N_19975);
xnor UO_1336 (O_1336,N_19980,N_19911);
or UO_1337 (O_1337,N_19623,N_19885);
nor UO_1338 (O_1338,N_19621,N_19629);
xor UO_1339 (O_1339,N_19552,N_19808);
nor UO_1340 (O_1340,N_19877,N_19579);
nor UO_1341 (O_1341,N_19528,N_19830);
xnor UO_1342 (O_1342,N_19701,N_19623);
and UO_1343 (O_1343,N_19935,N_19788);
and UO_1344 (O_1344,N_19851,N_19620);
and UO_1345 (O_1345,N_19846,N_19611);
nand UO_1346 (O_1346,N_19913,N_19669);
xor UO_1347 (O_1347,N_19974,N_19651);
or UO_1348 (O_1348,N_19960,N_19548);
xnor UO_1349 (O_1349,N_19663,N_19586);
and UO_1350 (O_1350,N_19612,N_19900);
nand UO_1351 (O_1351,N_19965,N_19598);
nor UO_1352 (O_1352,N_19818,N_19837);
or UO_1353 (O_1353,N_19743,N_19695);
xnor UO_1354 (O_1354,N_19799,N_19542);
and UO_1355 (O_1355,N_19667,N_19743);
xnor UO_1356 (O_1356,N_19719,N_19840);
or UO_1357 (O_1357,N_19987,N_19726);
nor UO_1358 (O_1358,N_19909,N_19939);
xor UO_1359 (O_1359,N_19974,N_19853);
nor UO_1360 (O_1360,N_19773,N_19890);
or UO_1361 (O_1361,N_19689,N_19899);
xor UO_1362 (O_1362,N_19948,N_19926);
xor UO_1363 (O_1363,N_19984,N_19683);
xor UO_1364 (O_1364,N_19710,N_19631);
nand UO_1365 (O_1365,N_19597,N_19512);
xor UO_1366 (O_1366,N_19661,N_19726);
and UO_1367 (O_1367,N_19801,N_19882);
nor UO_1368 (O_1368,N_19715,N_19978);
and UO_1369 (O_1369,N_19776,N_19517);
nor UO_1370 (O_1370,N_19989,N_19528);
nor UO_1371 (O_1371,N_19687,N_19896);
xor UO_1372 (O_1372,N_19835,N_19605);
or UO_1373 (O_1373,N_19739,N_19713);
or UO_1374 (O_1374,N_19832,N_19868);
nor UO_1375 (O_1375,N_19589,N_19526);
nor UO_1376 (O_1376,N_19549,N_19677);
xnor UO_1377 (O_1377,N_19911,N_19938);
nand UO_1378 (O_1378,N_19815,N_19887);
nand UO_1379 (O_1379,N_19716,N_19574);
and UO_1380 (O_1380,N_19620,N_19659);
and UO_1381 (O_1381,N_19728,N_19801);
or UO_1382 (O_1382,N_19501,N_19581);
nand UO_1383 (O_1383,N_19644,N_19587);
nand UO_1384 (O_1384,N_19956,N_19894);
and UO_1385 (O_1385,N_19679,N_19531);
and UO_1386 (O_1386,N_19883,N_19874);
xor UO_1387 (O_1387,N_19550,N_19585);
nand UO_1388 (O_1388,N_19547,N_19569);
nand UO_1389 (O_1389,N_19703,N_19924);
xor UO_1390 (O_1390,N_19648,N_19547);
nor UO_1391 (O_1391,N_19845,N_19659);
xnor UO_1392 (O_1392,N_19889,N_19804);
or UO_1393 (O_1393,N_19919,N_19925);
nand UO_1394 (O_1394,N_19583,N_19806);
or UO_1395 (O_1395,N_19805,N_19732);
or UO_1396 (O_1396,N_19665,N_19693);
nor UO_1397 (O_1397,N_19964,N_19889);
or UO_1398 (O_1398,N_19740,N_19777);
nor UO_1399 (O_1399,N_19703,N_19583);
nor UO_1400 (O_1400,N_19673,N_19632);
nor UO_1401 (O_1401,N_19858,N_19645);
and UO_1402 (O_1402,N_19624,N_19755);
nand UO_1403 (O_1403,N_19973,N_19995);
xor UO_1404 (O_1404,N_19921,N_19951);
xor UO_1405 (O_1405,N_19807,N_19837);
and UO_1406 (O_1406,N_19656,N_19665);
nand UO_1407 (O_1407,N_19591,N_19922);
nand UO_1408 (O_1408,N_19808,N_19847);
and UO_1409 (O_1409,N_19955,N_19722);
nor UO_1410 (O_1410,N_19826,N_19552);
nor UO_1411 (O_1411,N_19581,N_19830);
nor UO_1412 (O_1412,N_19872,N_19968);
or UO_1413 (O_1413,N_19537,N_19764);
nor UO_1414 (O_1414,N_19559,N_19624);
xnor UO_1415 (O_1415,N_19856,N_19766);
xor UO_1416 (O_1416,N_19709,N_19870);
xnor UO_1417 (O_1417,N_19856,N_19532);
nor UO_1418 (O_1418,N_19819,N_19792);
xnor UO_1419 (O_1419,N_19740,N_19810);
nand UO_1420 (O_1420,N_19526,N_19557);
nand UO_1421 (O_1421,N_19604,N_19695);
and UO_1422 (O_1422,N_19808,N_19880);
nand UO_1423 (O_1423,N_19821,N_19643);
xor UO_1424 (O_1424,N_19687,N_19615);
xor UO_1425 (O_1425,N_19798,N_19868);
and UO_1426 (O_1426,N_19521,N_19635);
nor UO_1427 (O_1427,N_19926,N_19982);
and UO_1428 (O_1428,N_19650,N_19831);
or UO_1429 (O_1429,N_19581,N_19510);
and UO_1430 (O_1430,N_19788,N_19937);
xor UO_1431 (O_1431,N_19626,N_19910);
and UO_1432 (O_1432,N_19943,N_19815);
nand UO_1433 (O_1433,N_19904,N_19957);
nor UO_1434 (O_1434,N_19534,N_19792);
nor UO_1435 (O_1435,N_19696,N_19602);
or UO_1436 (O_1436,N_19921,N_19714);
xnor UO_1437 (O_1437,N_19922,N_19819);
xor UO_1438 (O_1438,N_19791,N_19969);
nor UO_1439 (O_1439,N_19825,N_19999);
xnor UO_1440 (O_1440,N_19646,N_19651);
nand UO_1441 (O_1441,N_19919,N_19502);
nand UO_1442 (O_1442,N_19662,N_19516);
xnor UO_1443 (O_1443,N_19856,N_19968);
nand UO_1444 (O_1444,N_19767,N_19838);
nand UO_1445 (O_1445,N_19532,N_19976);
and UO_1446 (O_1446,N_19639,N_19844);
nand UO_1447 (O_1447,N_19971,N_19853);
and UO_1448 (O_1448,N_19606,N_19949);
and UO_1449 (O_1449,N_19545,N_19990);
nand UO_1450 (O_1450,N_19861,N_19887);
nor UO_1451 (O_1451,N_19988,N_19805);
xor UO_1452 (O_1452,N_19813,N_19554);
nand UO_1453 (O_1453,N_19821,N_19708);
nor UO_1454 (O_1454,N_19781,N_19679);
and UO_1455 (O_1455,N_19992,N_19506);
and UO_1456 (O_1456,N_19881,N_19756);
nor UO_1457 (O_1457,N_19851,N_19880);
and UO_1458 (O_1458,N_19615,N_19767);
nand UO_1459 (O_1459,N_19542,N_19501);
xor UO_1460 (O_1460,N_19913,N_19869);
nor UO_1461 (O_1461,N_19663,N_19889);
nand UO_1462 (O_1462,N_19919,N_19680);
xnor UO_1463 (O_1463,N_19926,N_19558);
xnor UO_1464 (O_1464,N_19881,N_19541);
nand UO_1465 (O_1465,N_19559,N_19871);
xor UO_1466 (O_1466,N_19647,N_19604);
and UO_1467 (O_1467,N_19856,N_19745);
and UO_1468 (O_1468,N_19718,N_19578);
nand UO_1469 (O_1469,N_19850,N_19658);
xor UO_1470 (O_1470,N_19515,N_19593);
nand UO_1471 (O_1471,N_19769,N_19624);
and UO_1472 (O_1472,N_19789,N_19769);
nor UO_1473 (O_1473,N_19509,N_19849);
or UO_1474 (O_1474,N_19781,N_19923);
nand UO_1475 (O_1475,N_19839,N_19586);
and UO_1476 (O_1476,N_19901,N_19994);
nor UO_1477 (O_1477,N_19830,N_19522);
nand UO_1478 (O_1478,N_19652,N_19912);
and UO_1479 (O_1479,N_19557,N_19856);
and UO_1480 (O_1480,N_19769,N_19706);
nand UO_1481 (O_1481,N_19601,N_19779);
xor UO_1482 (O_1482,N_19571,N_19779);
or UO_1483 (O_1483,N_19600,N_19500);
and UO_1484 (O_1484,N_19720,N_19822);
and UO_1485 (O_1485,N_19516,N_19755);
nor UO_1486 (O_1486,N_19632,N_19910);
nand UO_1487 (O_1487,N_19981,N_19625);
or UO_1488 (O_1488,N_19707,N_19750);
xnor UO_1489 (O_1489,N_19854,N_19803);
nand UO_1490 (O_1490,N_19790,N_19829);
nor UO_1491 (O_1491,N_19875,N_19888);
xnor UO_1492 (O_1492,N_19547,N_19539);
nor UO_1493 (O_1493,N_19836,N_19633);
nor UO_1494 (O_1494,N_19893,N_19673);
or UO_1495 (O_1495,N_19828,N_19636);
and UO_1496 (O_1496,N_19771,N_19628);
nand UO_1497 (O_1497,N_19992,N_19891);
nor UO_1498 (O_1498,N_19867,N_19752);
or UO_1499 (O_1499,N_19623,N_19543);
nor UO_1500 (O_1500,N_19645,N_19736);
and UO_1501 (O_1501,N_19745,N_19593);
nand UO_1502 (O_1502,N_19734,N_19660);
nor UO_1503 (O_1503,N_19724,N_19525);
nand UO_1504 (O_1504,N_19989,N_19934);
xnor UO_1505 (O_1505,N_19518,N_19778);
and UO_1506 (O_1506,N_19525,N_19779);
nand UO_1507 (O_1507,N_19873,N_19689);
and UO_1508 (O_1508,N_19911,N_19570);
xor UO_1509 (O_1509,N_19691,N_19686);
and UO_1510 (O_1510,N_19793,N_19527);
nand UO_1511 (O_1511,N_19973,N_19639);
nand UO_1512 (O_1512,N_19798,N_19925);
and UO_1513 (O_1513,N_19738,N_19624);
nand UO_1514 (O_1514,N_19968,N_19873);
nand UO_1515 (O_1515,N_19702,N_19651);
or UO_1516 (O_1516,N_19907,N_19936);
and UO_1517 (O_1517,N_19987,N_19592);
or UO_1518 (O_1518,N_19558,N_19793);
or UO_1519 (O_1519,N_19884,N_19634);
or UO_1520 (O_1520,N_19816,N_19799);
nand UO_1521 (O_1521,N_19676,N_19637);
and UO_1522 (O_1522,N_19513,N_19522);
nor UO_1523 (O_1523,N_19908,N_19969);
and UO_1524 (O_1524,N_19540,N_19560);
nand UO_1525 (O_1525,N_19533,N_19737);
xor UO_1526 (O_1526,N_19656,N_19994);
xnor UO_1527 (O_1527,N_19923,N_19693);
and UO_1528 (O_1528,N_19517,N_19654);
nor UO_1529 (O_1529,N_19715,N_19759);
and UO_1530 (O_1530,N_19873,N_19934);
and UO_1531 (O_1531,N_19768,N_19607);
nor UO_1532 (O_1532,N_19805,N_19675);
xor UO_1533 (O_1533,N_19746,N_19738);
nand UO_1534 (O_1534,N_19574,N_19749);
nand UO_1535 (O_1535,N_19991,N_19953);
nand UO_1536 (O_1536,N_19682,N_19863);
or UO_1537 (O_1537,N_19747,N_19918);
and UO_1538 (O_1538,N_19576,N_19892);
or UO_1539 (O_1539,N_19754,N_19956);
and UO_1540 (O_1540,N_19599,N_19998);
xor UO_1541 (O_1541,N_19692,N_19666);
and UO_1542 (O_1542,N_19551,N_19845);
nand UO_1543 (O_1543,N_19800,N_19757);
nor UO_1544 (O_1544,N_19722,N_19846);
nand UO_1545 (O_1545,N_19576,N_19847);
nor UO_1546 (O_1546,N_19644,N_19717);
or UO_1547 (O_1547,N_19718,N_19884);
and UO_1548 (O_1548,N_19611,N_19689);
nand UO_1549 (O_1549,N_19769,N_19599);
and UO_1550 (O_1550,N_19610,N_19738);
nand UO_1551 (O_1551,N_19654,N_19514);
nand UO_1552 (O_1552,N_19872,N_19504);
xnor UO_1553 (O_1553,N_19750,N_19720);
nand UO_1554 (O_1554,N_19730,N_19985);
xnor UO_1555 (O_1555,N_19533,N_19558);
or UO_1556 (O_1556,N_19863,N_19674);
or UO_1557 (O_1557,N_19624,N_19572);
nor UO_1558 (O_1558,N_19931,N_19812);
nor UO_1559 (O_1559,N_19963,N_19711);
xor UO_1560 (O_1560,N_19758,N_19880);
nor UO_1561 (O_1561,N_19737,N_19828);
xnor UO_1562 (O_1562,N_19529,N_19701);
or UO_1563 (O_1563,N_19675,N_19830);
xnor UO_1564 (O_1564,N_19574,N_19819);
xnor UO_1565 (O_1565,N_19751,N_19643);
or UO_1566 (O_1566,N_19829,N_19855);
xor UO_1567 (O_1567,N_19661,N_19718);
nand UO_1568 (O_1568,N_19779,N_19539);
nand UO_1569 (O_1569,N_19590,N_19671);
nor UO_1570 (O_1570,N_19614,N_19525);
and UO_1571 (O_1571,N_19918,N_19791);
and UO_1572 (O_1572,N_19705,N_19854);
nor UO_1573 (O_1573,N_19880,N_19517);
nand UO_1574 (O_1574,N_19686,N_19676);
xnor UO_1575 (O_1575,N_19694,N_19892);
nor UO_1576 (O_1576,N_19860,N_19636);
and UO_1577 (O_1577,N_19980,N_19843);
or UO_1578 (O_1578,N_19961,N_19778);
or UO_1579 (O_1579,N_19765,N_19982);
nand UO_1580 (O_1580,N_19693,N_19835);
nor UO_1581 (O_1581,N_19755,N_19908);
nand UO_1582 (O_1582,N_19832,N_19672);
nand UO_1583 (O_1583,N_19569,N_19840);
xor UO_1584 (O_1584,N_19862,N_19594);
nand UO_1585 (O_1585,N_19738,N_19626);
xnor UO_1586 (O_1586,N_19691,N_19779);
xor UO_1587 (O_1587,N_19606,N_19864);
nor UO_1588 (O_1588,N_19778,N_19525);
xor UO_1589 (O_1589,N_19550,N_19529);
and UO_1590 (O_1590,N_19984,N_19992);
or UO_1591 (O_1591,N_19843,N_19927);
nor UO_1592 (O_1592,N_19806,N_19588);
nand UO_1593 (O_1593,N_19644,N_19928);
or UO_1594 (O_1594,N_19518,N_19704);
nor UO_1595 (O_1595,N_19728,N_19589);
nor UO_1596 (O_1596,N_19774,N_19630);
and UO_1597 (O_1597,N_19755,N_19622);
xor UO_1598 (O_1598,N_19609,N_19606);
xnor UO_1599 (O_1599,N_19805,N_19840);
xor UO_1600 (O_1600,N_19589,N_19889);
or UO_1601 (O_1601,N_19602,N_19976);
nand UO_1602 (O_1602,N_19630,N_19538);
nand UO_1603 (O_1603,N_19780,N_19592);
nand UO_1604 (O_1604,N_19702,N_19774);
nand UO_1605 (O_1605,N_19529,N_19856);
nand UO_1606 (O_1606,N_19520,N_19766);
or UO_1607 (O_1607,N_19816,N_19878);
xnor UO_1608 (O_1608,N_19580,N_19791);
and UO_1609 (O_1609,N_19827,N_19508);
and UO_1610 (O_1610,N_19532,N_19947);
nand UO_1611 (O_1611,N_19776,N_19553);
nand UO_1612 (O_1612,N_19821,N_19948);
xnor UO_1613 (O_1613,N_19842,N_19885);
nand UO_1614 (O_1614,N_19741,N_19947);
nand UO_1615 (O_1615,N_19603,N_19518);
nor UO_1616 (O_1616,N_19783,N_19759);
nor UO_1617 (O_1617,N_19791,N_19910);
xnor UO_1618 (O_1618,N_19615,N_19901);
nor UO_1619 (O_1619,N_19717,N_19693);
nand UO_1620 (O_1620,N_19745,N_19501);
xnor UO_1621 (O_1621,N_19931,N_19773);
nand UO_1622 (O_1622,N_19689,N_19756);
or UO_1623 (O_1623,N_19561,N_19728);
xor UO_1624 (O_1624,N_19867,N_19771);
xnor UO_1625 (O_1625,N_19751,N_19664);
xor UO_1626 (O_1626,N_19668,N_19642);
nor UO_1627 (O_1627,N_19753,N_19692);
nand UO_1628 (O_1628,N_19616,N_19937);
nor UO_1629 (O_1629,N_19719,N_19820);
xor UO_1630 (O_1630,N_19921,N_19704);
nor UO_1631 (O_1631,N_19936,N_19504);
and UO_1632 (O_1632,N_19631,N_19916);
xnor UO_1633 (O_1633,N_19850,N_19758);
or UO_1634 (O_1634,N_19541,N_19804);
or UO_1635 (O_1635,N_19667,N_19936);
or UO_1636 (O_1636,N_19960,N_19558);
and UO_1637 (O_1637,N_19896,N_19635);
xnor UO_1638 (O_1638,N_19818,N_19549);
nand UO_1639 (O_1639,N_19933,N_19869);
xnor UO_1640 (O_1640,N_19862,N_19508);
xor UO_1641 (O_1641,N_19602,N_19691);
xor UO_1642 (O_1642,N_19739,N_19771);
xnor UO_1643 (O_1643,N_19665,N_19750);
or UO_1644 (O_1644,N_19985,N_19914);
nand UO_1645 (O_1645,N_19666,N_19567);
nor UO_1646 (O_1646,N_19579,N_19873);
nand UO_1647 (O_1647,N_19597,N_19912);
or UO_1648 (O_1648,N_19874,N_19915);
and UO_1649 (O_1649,N_19993,N_19651);
or UO_1650 (O_1650,N_19651,N_19843);
nand UO_1651 (O_1651,N_19771,N_19670);
and UO_1652 (O_1652,N_19896,N_19773);
and UO_1653 (O_1653,N_19666,N_19505);
and UO_1654 (O_1654,N_19928,N_19566);
nand UO_1655 (O_1655,N_19535,N_19595);
nor UO_1656 (O_1656,N_19748,N_19928);
and UO_1657 (O_1657,N_19505,N_19682);
nor UO_1658 (O_1658,N_19993,N_19972);
nand UO_1659 (O_1659,N_19881,N_19973);
or UO_1660 (O_1660,N_19963,N_19812);
xor UO_1661 (O_1661,N_19514,N_19674);
xnor UO_1662 (O_1662,N_19830,N_19989);
xor UO_1663 (O_1663,N_19711,N_19787);
and UO_1664 (O_1664,N_19872,N_19664);
and UO_1665 (O_1665,N_19561,N_19889);
xnor UO_1666 (O_1666,N_19895,N_19626);
or UO_1667 (O_1667,N_19677,N_19724);
nand UO_1668 (O_1668,N_19844,N_19910);
nor UO_1669 (O_1669,N_19554,N_19879);
and UO_1670 (O_1670,N_19724,N_19594);
or UO_1671 (O_1671,N_19600,N_19598);
or UO_1672 (O_1672,N_19780,N_19934);
nor UO_1673 (O_1673,N_19734,N_19748);
and UO_1674 (O_1674,N_19799,N_19767);
nor UO_1675 (O_1675,N_19669,N_19850);
nand UO_1676 (O_1676,N_19725,N_19857);
and UO_1677 (O_1677,N_19895,N_19975);
nand UO_1678 (O_1678,N_19785,N_19593);
and UO_1679 (O_1679,N_19878,N_19877);
nand UO_1680 (O_1680,N_19767,N_19904);
nor UO_1681 (O_1681,N_19746,N_19689);
or UO_1682 (O_1682,N_19545,N_19667);
or UO_1683 (O_1683,N_19823,N_19647);
nor UO_1684 (O_1684,N_19985,N_19904);
nand UO_1685 (O_1685,N_19745,N_19677);
or UO_1686 (O_1686,N_19632,N_19740);
and UO_1687 (O_1687,N_19985,N_19759);
or UO_1688 (O_1688,N_19712,N_19546);
and UO_1689 (O_1689,N_19587,N_19741);
nor UO_1690 (O_1690,N_19547,N_19635);
and UO_1691 (O_1691,N_19669,N_19910);
nand UO_1692 (O_1692,N_19736,N_19738);
xor UO_1693 (O_1693,N_19596,N_19736);
and UO_1694 (O_1694,N_19967,N_19702);
and UO_1695 (O_1695,N_19677,N_19593);
or UO_1696 (O_1696,N_19975,N_19610);
nor UO_1697 (O_1697,N_19566,N_19500);
and UO_1698 (O_1698,N_19560,N_19546);
and UO_1699 (O_1699,N_19980,N_19710);
nor UO_1700 (O_1700,N_19557,N_19687);
nor UO_1701 (O_1701,N_19965,N_19814);
or UO_1702 (O_1702,N_19985,N_19690);
nor UO_1703 (O_1703,N_19721,N_19539);
nand UO_1704 (O_1704,N_19920,N_19687);
nor UO_1705 (O_1705,N_19579,N_19558);
nor UO_1706 (O_1706,N_19787,N_19644);
nor UO_1707 (O_1707,N_19656,N_19674);
nand UO_1708 (O_1708,N_19944,N_19768);
or UO_1709 (O_1709,N_19809,N_19578);
and UO_1710 (O_1710,N_19767,N_19797);
nor UO_1711 (O_1711,N_19763,N_19702);
or UO_1712 (O_1712,N_19785,N_19934);
and UO_1713 (O_1713,N_19532,N_19950);
and UO_1714 (O_1714,N_19768,N_19526);
or UO_1715 (O_1715,N_19965,N_19800);
or UO_1716 (O_1716,N_19518,N_19836);
nand UO_1717 (O_1717,N_19739,N_19805);
xnor UO_1718 (O_1718,N_19852,N_19723);
nand UO_1719 (O_1719,N_19607,N_19745);
nand UO_1720 (O_1720,N_19752,N_19688);
nor UO_1721 (O_1721,N_19818,N_19957);
nand UO_1722 (O_1722,N_19779,N_19992);
or UO_1723 (O_1723,N_19815,N_19656);
nor UO_1724 (O_1724,N_19883,N_19521);
nor UO_1725 (O_1725,N_19953,N_19900);
xnor UO_1726 (O_1726,N_19568,N_19785);
or UO_1727 (O_1727,N_19742,N_19924);
or UO_1728 (O_1728,N_19871,N_19566);
and UO_1729 (O_1729,N_19900,N_19687);
nand UO_1730 (O_1730,N_19965,N_19681);
nand UO_1731 (O_1731,N_19531,N_19702);
xnor UO_1732 (O_1732,N_19801,N_19671);
and UO_1733 (O_1733,N_19717,N_19559);
and UO_1734 (O_1734,N_19598,N_19689);
and UO_1735 (O_1735,N_19998,N_19872);
xnor UO_1736 (O_1736,N_19902,N_19790);
xor UO_1737 (O_1737,N_19976,N_19911);
nand UO_1738 (O_1738,N_19680,N_19761);
xnor UO_1739 (O_1739,N_19666,N_19765);
and UO_1740 (O_1740,N_19910,N_19903);
or UO_1741 (O_1741,N_19560,N_19629);
xnor UO_1742 (O_1742,N_19770,N_19673);
nand UO_1743 (O_1743,N_19673,N_19740);
xor UO_1744 (O_1744,N_19541,N_19578);
nor UO_1745 (O_1745,N_19685,N_19668);
xor UO_1746 (O_1746,N_19696,N_19979);
and UO_1747 (O_1747,N_19692,N_19642);
nand UO_1748 (O_1748,N_19927,N_19896);
xor UO_1749 (O_1749,N_19905,N_19860);
xnor UO_1750 (O_1750,N_19914,N_19864);
and UO_1751 (O_1751,N_19901,N_19648);
nor UO_1752 (O_1752,N_19922,N_19844);
or UO_1753 (O_1753,N_19922,N_19750);
and UO_1754 (O_1754,N_19897,N_19907);
or UO_1755 (O_1755,N_19521,N_19693);
nand UO_1756 (O_1756,N_19739,N_19881);
nand UO_1757 (O_1757,N_19507,N_19504);
nand UO_1758 (O_1758,N_19759,N_19864);
or UO_1759 (O_1759,N_19531,N_19760);
and UO_1760 (O_1760,N_19756,N_19601);
nand UO_1761 (O_1761,N_19604,N_19708);
or UO_1762 (O_1762,N_19576,N_19725);
and UO_1763 (O_1763,N_19532,N_19604);
and UO_1764 (O_1764,N_19960,N_19981);
nand UO_1765 (O_1765,N_19847,N_19965);
nor UO_1766 (O_1766,N_19862,N_19627);
xor UO_1767 (O_1767,N_19934,N_19712);
or UO_1768 (O_1768,N_19834,N_19724);
nor UO_1769 (O_1769,N_19796,N_19500);
nand UO_1770 (O_1770,N_19536,N_19718);
and UO_1771 (O_1771,N_19713,N_19682);
or UO_1772 (O_1772,N_19788,N_19883);
xor UO_1773 (O_1773,N_19730,N_19939);
nor UO_1774 (O_1774,N_19717,N_19711);
or UO_1775 (O_1775,N_19661,N_19977);
xnor UO_1776 (O_1776,N_19701,N_19835);
and UO_1777 (O_1777,N_19807,N_19998);
nor UO_1778 (O_1778,N_19645,N_19503);
or UO_1779 (O_1779,N_19794,N_19843);
and UO_1780 (O_1780,N_19879,N_19960);
nor UO_1781 (O_1781,N_19868,N_19696);
nand UO_1782 (O_1782,N_19748,N_19802);
or UO_1783 (O_1783,N_19816,N_19543);
nand UO_1784 (O_1784,N_19608,N_19907);
and UO_1785 (O_1785,N_19937,N_19965);
nand UO_1786 (O_1786,N_19635,N_19623);
or UO_1787 (O_1787,N_19914,N_19801);
nor UO_1788 (O_1788,N_19797,N_19628);
and UO_1789 (O_1789,N_19588,N_19738);
and UO_1790 (O_1790,N_19714,N_19700);
xnor UO_1791 (O_1791,N_19708,N_19857);
nand UO_1792 (O_1792,N_19584,N_19769);
xnor UO_1793 (O_1793,N_19536,N_19813);
xnor UO_1794 (O_1794,N_19775,N_19662);
or UO_1795 (O_1795,N_19835,N_19676);
or UO_1796 (O_1796,N_19586,N_19733);
or UO_1797 (O_1797,N_19839,N_19761);
or UO_1798 (O_1798,N_19926,N_19601);
and UO_1799 (O_1799,N_19526,N_19745);
or UO_1800 (O_1800,N_19855,N_19819);
nor UO_1801 (O_1801,N_19991,N_19875);
and UO_1802 (O_1802,N_19991,N_19941);
or UO_1803 (O_1803,N_19908,N_19677);
or UO_1804 (O_1804,N_19854,N_19721);
nor UO_1805 (O_1805,N_19626,N_19562);
nand UO_1806 (O_1806,N_19901,N_19523);
or UO_1807 (O_1807,N_19797,N_19828);
xnor UO_1808 (O_1808,N_19867,N_19595);
nor UO_1809 (O_1809,N_19932,N_19611);
and UO_1810 (O_1810,N_19917,N_19626);
or UO_1811 (O_1811,N_19887,N_19551);
and UO_1812 (O_1812,N_19510,N_19904);
nand UO_1813 (O_1813,N_19695,N_19971);
nand UO_1814 (O_1814,N_19889,N_19810);
nand UO_1815 (O_1815,N_19574,N_19502);
and UO_1816 (O_1816,N_19849,N_19748);
xor UO_1817 (O_1817,N_19779,N_19987);
nor UO_1818 (O_1818,N_19873,N_19979);
and UO_1819 (O_1819,N_19729,N_19573);
xor UO_1820 (O_1820,N_19724,N_19701);
and UO_1821 (O_1821,N_19581,N_19975);
and UO_1822 (O_1822,N_19578,N_19632);
nand UO_1823 (O_1823,N_19678,N_19646);
xor UO_1824 (O_1824,N_19552,N_19977);
nor UO_1825 (O_1825,N_19776,N_19943);
or UO_1826 (O_1826,N_19856,N_19539);
xnor UO_1827 (O_1827,N_19848,N_19952);
nor UO_1828 (O_1828,N_19810,N_19798);
nor UO_1829 (O_1829,N_19942,N_19988);
nor UO_1830 (O_1830,N_19556,N_19900);
and UO_1831 (O_1831,N_19650,N_19547);
nor UO_1832 (O_1832,N_19595,N_19917);
xor UO_1833 (O_1833,N_19585,N_19991);
nor UO_1834 (O_1834,N_19909,N_19786);
nand UO_1835 (O_1835,N_19811,N_19695);
or UO_1836 (O_1836,N_19662,N_19715);
nand UO_1837 (O_1837,N_19742,N_19941);
nand UO_1838 (O_1838,N_19912,N_19610);
xor UO_1839 (O_1839,N_19649,N_19842);
nor UO_1840 (O_1840,N_19653,N_19856);
nor UO_1841 (O_1841,N_19958,N_19625);
or UO_1842 (O_1842,N_19594,N_19580);
and UO_1843 (O_1843,N_19619,N_19660);
and UO_1844 (O_1844,N_19854,N_19852);
and UO_1845 (O_1845,N_19846,N_19630);
xnor UO_1846 (O_1846,N_19721,N_19723);
and UO_1847 (O_1847,N_19562,N_19744);
and UO_1848 (O_1848,N_19500,N_19705);
nor UO_1849 (O_1849,N_19946,N_19523);
nor UO_1850 (O_1850,N_19558,N_19778);
or UO_1851 (O_1851,N_19631,N_19650);
and UO_1852 (O_1852,N_19909,N_19593);
xnor UO_1853 (O_1853,N_19703,N_19900);
nand UO_1854 (O_1854,N_19718,N_19827);
or UO_1855 (O_1855,N_19814,N_19667);
xnor UO_1856 (O_1856,N_19767,N_19785);
or UO_1857 (O_1857,N_19873,N_19965);
and UO_1858 (O_1858,N_19878,N_19533);
or UO_1859 (O_1859,N_19708,N_19697);
nand UO_1860 (O_1860,N_19832,N_19662);
or UO_1861 (O_1861,N_19993,N_19946);
and UO_1862 (O_1862,N_19903,N_19912);
and UO_1863 (O_1863,N_19563,N_19740);
and UO_1864 (O_1864,N_19730,N_19751);
nand UO_1865 (O_1865,N_19666,N_19664);
nor UO_1866 (O_1866,N_19960,N_19552);
nor UO_1867 (O_1867,N_19581,N_19604);
xor UO_1868 (O_1868,N_19890,N_19551);
nor UO_1869 (O_1869,N_19581,N_19982);
xnor UO_1870 (O_1870,N_19965,N_19725);
xor UO_1871 (O_1871,N_19638,N_19785);
or UO_1872 (O_1872,N_19553,N_19773);
xnor UO_1873 (O_1873,N_19777,N_19882);
and UO_1874 (O_1874,N_19681,N_19759);
xor UO_1875 (O_1875,N_19853,N_19517);
nor UO_1876 (O_1876,N_19962,N_19626);
or UO_1877 (O_1877,N_19919,N_19562);
nor UO_1878 (O_1878,N_19997,N_19823);
nor UO_1879 (O_1879,N_19757,N_19721);
or UO_1880 (O_1880,N_19921,N_19851);
xor UO_1881 (O_1881,N_19797,N_19880);
or UO_1882 (O_1882,N_19751,N_19839);
or UO_1883 (O_1883,N_19930,N_19740);
nand UO_1884 (O_1884,N_19834,N_19597);
and UO_1885 (O_1885,N_19875,N_19864);
xnor UO_1886 (O_1886,N_19808,N_19866);
and UO_1887 (O_1887,N_19960,N_19958);
xor UO_1888 (O_1888,N_19628,N_19614);
nor UO_1889 (O_1889,N_19701,N_19914);
and UO_1890 (O_1890,N_19752,N_19977);
xnor UO_1891 (O_1891,N_19890,N_19552);
nand UO_1892 (O_1892,N_19598,N_19753);
nand UO_1893 (O_1893,N_19704,N_19662);
nor UO_1894 (O_1894,N_19875,N_19707);
nand UO_1895 (O_1895,N_19853,N_19959);
nand UO_1896 (O_1896,N_19551,N_19769);
nor UO_1897 (O_1897,N_19597,N_19769);
nand UO_1898 (O_1898,N_19963,N_19623);
nand UO_1899 (O_1899,N_19904,N_19784);
xor UO_1900 (O_1900,N_19642,N_19812);
or UO_1901 (O_1901,N_19598,N_19940);
and UO_1902 (O_1902,N_19852,N_19834);
xnor UO_1903 (O_1903,N_19641,N_19775);
nand UO_1904 (O_1904,N_19778,N_19600);
nor UO_1905 (O_1905,N_19687,N_19640);
nor UO_1906 (O_1906,N_19699,N_19839);
nand UO_1907 (O_1907,N_19671,N_19859);
nor UO_1908 (O_1908,N_19851,N_19893);
nor UO_1909 (O_1909,N_19622,N_19790);
and UO_1910 (O_1910,N_19839,N_19820);
or UO_1911 (O_1911,N_19520,N_19831);
or UO_1912 (O_1912,N_19520,N_19625);
xnor UO_1913 (O_1913,N_19932,N_19961);
nand UO_1914 (O_1914,N_19792,N_19692);
nor UO_1915 (O_1915,N_19532,N_19530);
nor UO_1916 (O_1916,N_19770,N_19589);
and UO_1917 (O_1917,N_19741,N_19660);
nor UO_1918 (O_1918,N_19896,N_19971);
nand UO_1919 (O_1919,N_19547,N_19713);
nor UO_1920 (O_1920,N_19835,N_19717);
xnor UO_1921 (O_1921,N_19880,N_19985);
nor UO_1922 (O_1922,N_19885,N_19941);
nor UO_1923 (O_1923,N_19886,N_19579);
nand UO_1924 (O_1924,N_19853,N_19761);
and UO_1925 (O_1925,N_19985,N_19739);
xnor UO_1926 (O_1926,N_19674,N_19865);
nor UO_1927 (O_1927,N_19994,N_19996);
nand UO_1928 (O_1928,N_19706,N_19747);
or UO_1929 (O_1929,N_19970,N_19591);
nor UO_1930 (O_1930,N_19548,N_19870);
nand UO_1931 (O_1931,N_19647,N_19677);
or UO_1932 (O_1932,N_19803,N_19858);
nor UO_1933 (O_1933,N_19820,N_19624);
xnor UO_1934 (O_1934,N_19747,N_19671);
nor UO_1935 (O_1935,N_19552,N_19813);
nand UO_1936 (O_1936,N_19745,N_19559);
and UO_1937 (O_1937,N_19692,N_19860);
or UO_1938 (O_1938,N_19847,N_19602);
xor UO_1939 (O_1939,N_19571,N_19583);
and UO_1940 (O_1940,N_19764,N_19818);
nand UO_1941 (O_1941,N_19678,N_19958);
or UO_1942 (O_1942,N_19717,N_19530);
xnor UO_1943 (O_1943,N_19680,N_19585);
or UO_1944 (O_1944,N_19694,N_19723);
or UO_1945 (O_1945,N_19512,N_19809);
xnor UO_1946 (O_1946,N_19858,N_19670);
and UO_1947 (O_1947,N_19770,N_19621);
xor UO_1948 (O_1948,N_19845,N_19986);
and UO_1949 (O_1949,N_19597,N_19917);
nor UO_1950 (O_1950,N_19864,N_19927);
and UO_1951 (O_1951,N_19807,N_19780);
nor UO_1952 (O_1952,N_19631,N_19763);
xnor UO_1953 (O_1953,N_19822,N_19678);
or UO_1954 (O_1954,N_19824,N_19696);
or UO_1955 (O_1955,N_19730,N_19537);
or UO_1956 (O_1956,N_19770,N_19698);
nand UO_1957 (O_1957,N_19873,N_19668);
xnor UO_1958 (O_1958,N_19671,N_19524);
xnor UO_1959 (O_1959,N_19993,N_19963);
and UO_1960 (O_1960,N_19856,N_19850);
xnor UO_1961 (O_1961,N_19557,N_19581);
xor UO_1962 (O_1962,N_19963,N_19941);
nor UO_1963 (O_1963,N_19826,N_19642);
xor UO_1964 (O_1964,N_19847,N_19541);
and UO_1965 (O_1965,N_19829,N_19709);
nand UO_1966 (O_1966,N_19947,N_19799);
or UO_1967 (O_1967,N_19777,N_19623);
or UO_1968 (O_1968,N_19897,N_19711);
nor UO_1969 (O_1969,N_19736,N_19765);
and UO_1970 (O_1970,N_19763,N_19526);
or UO_1971 (O_1971,N_19500,N_19550);
and UO_1972 (O_1972,N_19779,N_19706);
xnor UO_1973 (O_1973,N_19823,N_19552);
xnor UO_1974 (O_1974,N_19862,N_19706);
or UO_1975 (O_1975,N_19646,N_19991);
nor UO_1976 (O_1976,N_19844,N_19646);
nand UO_1977 (O_1977,N_19688,N_19661);
xnor UO_1978 (O_1978,N_19919,N_19851);
nand UO_1979 (O_1979,N_19896,N_19669);
nand UO_1980 (O_1980,N_19823,N_19953);
nand UO_1981 (O_1981,N_19586,N_19673);
or UO_1982 (O_1982,N_19735,N_19924);
or UO_1983 (O_1983,N_19502,N_19645);
nand UO_1984 (O_1984,N_19665,N_19953);
nor UO_1985 (O_1985,N_19891,N_19647);
and UO_1986 (O_1986,N_19899,N_19934);
xnor UO_1987 (O_1987,N_19808,N_19662);
and UO_1988 (O_1988,N_19949,N_19922);
nor UO_1989 (O_1989,N_19980,N_19926);
xor UO_1990 (O_1990,N_19920,N_19872);
xor UO_1991 (O_1991,N_19787,N_19754);
or UO_1992 (O_1992,N_19863,N_19770);
nand UO_1993 (O_1993,N_19975,N_19626);
and UO_1994 (O_1994,N_19551,N_19917);
xor UO_1995 (O_1995,N_19506,N_19683);
nand UO_1996 (O_1996,N_19730,N_19694);
or UO_1997 (O_1997,N_19820,N_19739);
nand UO_1998 (O_1998,N_19670,N_19630);
or UO_1999 (O_1999,N_19700,N_19632);
and UO_2000 (O_2000,N_19912,N_19905);
xnor UO_2001 (O_2001,N_19860,N_19765);
nand UO_2002 (O_2002,N_19597,N_19890);
nor UO_2003 (O_2003,N_19900,N_19944);
and UO_2004 (O_2004,N_19614,N_19869);
and UO_2005 (O_2005,N_19571,N_19811);
xnor UO_2006 (O_2006,N_19674,N_19648);
nor UO_2007 (O_2007,N_19658,N_19941);
nand UO_2008 (O_2008,N_19946,N_19809);
xor UO_2009 (O_2009,N_19885,N_19859);
nand UO_2010 (O_2010,N_19569,N_19885);
and UO_2011 (O_2011,N_19788,N_19619);
and UO_2012 (O_2012,N_19866,N_19860);
nand UO_2013 (O_2013,N_19642,N_19835);
xnor UO_2014 (O_2014,N_19866,N_19700);
nand UO_2015 (O_2015,N_19812,N_19899);
nand UO_2016 (O_2016,N_19797,N_19551);
and UO_2017 (O_2017,N_19983,N_19601);
nor UO_2018 (O_2018,N_19907,N_19900);
nand UO_2019 (O_2019,N_19675,N_19728);
nand UO_2020 (O_2020,N_19578,N_19756);
or UO_2021 (O_2021,N_19976,N_19758);
or UO_2022 (O_2022,N_19812,N_19808);
nand UO_2023 (O_2023,N_19604,N_19537);
and UO_2024 (O_2024,N_19760,N_19919);
and UO_2025 (O_2025,N_19675,N_19801);
xnor UO_2026 (O_2026,N_19994,N_19512);
or UO_2027 (O_2027,N_19700,N_19811);
or UO_2028 (O_2028,N_19503,N_19869);
nand UO_2029 (O_2029,N_19633,N_19924);
xnor UO_2030 (O_2030,N_19814,N_19657);
nor UO_2031 (O_2031,N_19618,N_19950);
nand UO_2032 (O_2032,N_19766,N_19505);
and UO_2033 (O_2033,N_19800,N_19902);
nor UO_2034 (O_2034,N_19718,N_19816);
and UO_2035 (O_2035,N_19915,N_19956);
nor UO_2036 (O_2036,N_19845,N_19667);
and UO_2037 (O_2037,N_19715,N_19657);
nand UO_2038 (O_2038,N_19742,N_19575);
and UO_2039 (O_2039,N_19773,N_19744);
xnor UO_2040 (O_2040,N_19787,N_19766);
and UO_2041 (O_2041,N_19858,N_19867);
and UO_2042 (O_2042,N_19519,N_19529);
and UO_2043 (O_2043,N_19840,N_19606);
or UO_2044 (O_2044,N_19671,N_19565);
nand UO_2045 (O_2045,N_19655,N_19670);
and UO_2046 (O_2046,N_19620,N_19532);
and UO_2047 (O_2047,N_19679,N_19599);
nor UO_2048 (O_2048,N_19718,N_19988);
and UO_2049 (O_2049,N_19973,N_19757);
or UO_2050 (O_2050,N_19530,N_19618);
nand UO_2051 (O_2051,N_19901,N_19510);
and UO_2052 (O_2052,N_19694,N_19993);
or UO_2053 (O_2053,N_19625,N_19934);
nand UO_2054 (O_2054,N_19716,N_19687);
and UO_2055 (O_2055,N_19866,N_19942);
nand UO_2056 (O_2056,N_19529,N_19624);
xor UO_2057 (O_2057,N_19584,N_19816);
or UO_2058 (O_2058,N_19536,N_19675);
xnor UO_2059 (O_2059,N_19652,N_19833);
nand UO_2060 (O_2060,N_19948,N_19573);
xor UO_2061 (O_2061,N_19642,N_19718);
nor UO_2062 (O_2062,N_19624,N_19721);
and UO_2063 (O_2063,N_19586,N_19976);
or UO_2064 (O_2064,N_19589,N_19997);
and UO_2065 (O_2065,N_19831,N_19791);
and UO_2066 (O_2066,N_19594,N_19559);
nor UO_2067 (O_2067,N_19600,N_19510);
and UO_2068 (O_2068,N_19669,N_19847);
nor UO_2069 (O_2069,N_19907,N_19847);
or UO_2070 (O_2070,N_19662,N_19535);
xnor UO_2071 (O_2071,N_19734,N_19671);
nor UO_2072 (O_2072,N_19505,N_19966);
and UO_2073 (O_2073,N_19644,N_19808);
and UO_2074 (O_2074,N_19984,N_19820);
nand UO_2075 (O_2075,N_19562,N_19606);
nand UO_2076 (O_2076,N_19585,N_19950);
or UO_2077 (O_2077,N_19530,N_19898);
xor UO_2078 (O_2078,N_19794,N_19969);
or UO_2079 (O_2079,N_19813,N_19759);
or UO_2080 (O_2080,N_19673,N_19668);
and UO_2081 (O_2081,N_19687,N_19638);
nand UO_2082 (O_2082,N_19964,N_19656);
or UO_2083 (O_2083,N_19873,N_19583);
nand UO_2084 (O_2084,N_19965,N_19802);
xnor UO_2085 (O_2085,N_19859,N_19839);
nand UO_2086 (O_2086,N_19807,N_19757);
or UO_2087 (O_2087,N_19526,N_19964);
nand UO_2088 (O_2088,N_19878,N_19822);
nand UO_2089 (O_2089,N_19670,N_19563);
or UO_2090 (O_2090,N_19500,N_19681);
xnor UO_2091 (O_2091,N_19619,N_19562);
nand UO_2092 (O_2092,N_19607,N_19960);
nor UO_2093 (O_2093,N_19823,N_19842);
xor UO_2094 (O_2094,N_19963,N_19513);
nor UO_2095 (O_2095,N_19503,N_19996);
or UO_2096 (O_2096,N_19675,N_19542);
xor UO_2097 (O_2097,N_19533,N_19938);
nor UO_2098 (O_2098,N_19956,N_19799);
and UO_2099 (O_2099,N_19565,N_19822);
nor UO_2100 (O_2100,N_19989,N_19894);
nor UO_2101 (O_2101,N_19716,N_19644);
nor UO_2102 (O_2102,N_19699,N_19665);
nand UO_2103 (O_2103,N_19975,N_19753);
and UO_2104 (O_2104,N_19606,N_19518);
and UO_2105 (O_2105,N_19880,N_19607);
nand UO_2106 (O_2106,N_19958,N_19640);
xnor UO_2107 (O_2107,N_19621,N_19709);
and UO_2108 (O_2108,N_19611,N_19715);
nand UO_2109 (O_2109,N_19521,N_19911);
nand UO_2110 (O_2110,N_19548,N_19624);
and UO_2111 (O_2111,N_19815,N_19553);
and UO_2112 (O_2112,N_19581,N_19914);
and UO_2113 (O_2113,N_19879,N_19986);
xor UO_2114 (O_2114,N_19984,N_19715);
nor UO_2115 (O_2115,N_19977,N_19704);
xnor UO_2116 (O_2116,N_19723,N_19571);
or UO_2117 (O_2117,N_19678,N_19788);
or UO_2118 (O_2118,N_19577,N_19594);
nor UO_2119 (O_2119,N_19965,N_19593);
nor UO_2120 (O_2120,N_19921,N_19610);
xor UO_2121 (O_2121,N_19981,N_19901);
or UO_2122 (O_2122,N_19815,N_19904);
or UO_2123 (O_2123,N_19554,N_19906);
and UO_2124 (O_2124,N_19723,N_19798);
nand UO_2125 (O_2125,N_19645,N_19667);
and UO_2126 (O_2126,N_19621,N_19937);
nor UO_2127 (O_2127,N_19685,N_19951);
nand UO_2128 (O_2128,N_19553,N_19831);
nand UO_2129 (O_2129,N_19641,N_19899);
or UO_2130 (O_2130,N_19675,N_19546);
xnor UO_2131 (O_2131,N_19630,N_19988);
xor UO_2132 (O_2132,N_19710,N_19611);
nor UO_2133 (O_2133,N_19810,N_19875);
and UO_2134 (O_2134,N_19527,N_19513);
and UO_2135 (O_2135,N_19728,N_19610);
nand UO_2136 (O_2136,N_19952,N_19778);
xor UO_2137 (O_2137,N_19692,N_19589);
nor UO_2138 (O_2138,N_19688,N_19958);
nor UO_2139 (O_2139,N_19861,N_19821);
and UO_2140 (O_2140,N_19728,N_19922);
nor UO_2141 (O_2141,N_19623,N_19847);
xnor UO_2142 (O_2142,N_19988,N_19957);
xor UO_2143 (O_2143,N_19581,N_19880);
and UO_2144 (O_2144,N_19784,N_19521);
and UO_2145 (O_2145,N_19650,N_19536);
and UO_2146 (O_2146,N_19850,N_19863);
or UO_2147 (O_2147,N_19846,N_19619);
nor UO_2148 (O_2148,N_19695,N_19822);
nand UO_2149 (O_2149,N_19584,N_19570);
nand UO_2150 (O_2150,N_19774,N_19666);
xnor UO_2151 (O_2151,N_19754,N_19772);
and UO_2152 (O_2152,N_19631,N_19842);
or UO_2153 (O_2153,N_19707,N_19898);
xnor UO_2154 (O_2154,N_19698,N_19716);
nor UO_2155 (O_2155,N_19647,N_19894);
and UO_2156 (O_2156,N_19908,N_19627);
xor UO_2157 (O_2157,N_19509,N_19695);
nand UO_2158 (O_2158,N_19827,N_19594);
or UO_2159 (O_2159,N_19540,N_19581);
nand UO_2160 (O_2160,N_19840,N_19779);
xnor UO_2161 (O_2161,N_19939,N_19956);
or UO_2162 (O_2162,N_19908,N_19961);
xnor UO_2163 (O_2163,N_19615,N_19877);
or UO_2164 (O_2164,N_19853,N_19772);
nor UO_2165 (O_2165,N_19656,N_19796);
and UO_2166 (O_2166,N_19668,N_19500);
or UO_2167 (O_2167,N_19505,N_19671);
nor UO_2168 (O_2168,N_19522,N_19884);
nand UO_2169 (O_2169,N_19650,N_19540);
xor UO_2170 (O_2170,N_19966,N_19957);
or UO_2171 (O_2171,N_19841,N_19646);
and UO_2172 (O_2172,N_19811,N_19674);
or UO_2173 (O_2173,N_19514,N_19827);
nor UO_2174 (O_2174,N_19725,N_19612);
or UO_2175 (O_2175,N_19837,N_19591);
nand UO_2176 (O_2176,N_19977,N_19829);
xor UO_2177 (O_2177,N_19561,N_19778);
or UO_2178 (O_2178,N_19640,N_19642);
or UO_2179 (O_2179,N_19593,N_19568);
nor UO_2180 (O_2180,N_19833,N_19915);
nor UO_2181 (O_2181,N_19647,N_19642);
and UO_2182 (O_2182,N_19839,N_19750);
xor UO_2183 (O_2183,N_19742,N_19778);
xnor UO_2184 (O_2184,N_19750,N_19711);
nor UO_2185 (O_2185,N_19569,N_19555);
nor UO_2186 (O_2186,N_19563,N_19866);
and UO_2187 (O_2187,N_19650,N_19909);
xor UO_2188 (O_2188,N_19526,N_19523);
or UO_2189 (O_2189,N_19744,N_19903);
or UO_2190 (O_2190,N_19946,N_19507);
and UO_2191 (O_2191,N_19993,N_19962);
xnor UO_2192 (O_2192,N_19844,N_19874);
nor UO_2193 (O_2193,N_19860,N_19749);
or UO_2194 (O_2194,N_19754,N_19503);
nor UO_2195 (O_2195,N_19801,N_19752);
and UO_2196 (O_2196,N_19516,N_19920);
nand UO_2197 (O_2197,N_19573,N_19870);
or UO_2198 (O_2198,N_19916,N_19673);
and UO_2199 (O_2199,N_19509,N_19554);
nand UO_2200 (O_2200,N_19702,N_19916);
or UO_2201 (O_2201,N_19874,N_19633);
nor UO_2202 (O_2202,N_19595,N_19954);
nand UO_2203 (O_2203,N_19699,N_19964);
and UO_2204 (O_2204,N_19899,N_19693);
and UO_2205 (O_2205,N_19752,N_19587);
nand UO_2206 (O_2206,N_19849,N_19730);
nor UO_2207 (O_2207,N_19654,N_19827);
or UO_2208 (O_2208,N_19625,N_19858);
nor UO_2209 (O_2209,N_19949,N_19610);
and UO_2210 (O_2210,N_19654,N_19987);
or UO_2211 (O_2211,N_19697,N_19590);
and UO_2212 (O_2212,N_19681,N_19820);
nand UO_2213 (O_2213,N_19742,N_19986);
or UO_2214 (O_2214,N_19633,N_19690);
nand UO_2215 (O_2215,N_19769,N_19889);
or UO_2216 (O_2216,N_19626,N_19776);
xnor UO_2217 (O_2217,N_19564,N_19821);
or UO_2218 (O_2218,N_19786,N_19750);
xnor UO_2219 (O_2219,N_19756,N_19842);
xor UO_2220 (O_2220,N_19983,N_19543);
xor UO_2221 (O_2221,N_19838,N_19703);
and UO_2222 (O_2222,N_19600,N_19766);
nand UO_2223 (O_2223,N_19606,N_19974);
nand UO_2224 (O_2224,N_19583,N_19723);
nor UO_2225 (O_2225,N_19636,N_19677);
nand UO_2226 (O_2226,N_19770,N_19684);
or UO_2227 (O_2227,N_19804,N_19676);
xnor UO_2228 (O_2228,N_19924,N_19832);
or UO_2229 (O_2229,N_19644,N_19762);
xor UO_2230 (O_2230,N_19953,N_19903);
nand UO_2231 (O_2231,N_19681,N_19548);
nor UO_2232 (O_2232,N_19617,N_19852);
nand UO_2233 (O_2233,N_19747,N_19709);
xor UO_2234 (O_2234,N_19727,N_19920);
nor UO_2235 (O_2235,N_19532,N_19614);
nor UO_2236 (O_2236,N_19976,N_19923);
xor UO_2237 (O_2237,N_19722,N_19646);
xor UO_2238 (O_2238,N_19893,N_19553);
and UO_2239 (O_2239,N_19686,N_19502);
nor UO_2240 (O_2240,N_19954,N_19584);
nand UO_2241 (O_2241,N_19849,N_19569);
nand UO_2242 (O_2242,N_19905,N_19940);
nand UO_2243 (O_2243,N_19905,N_19735);
xor UO_2244 (O_2244,N_19767,N_19897);
or UO_2245 (O_2245,N_19983,N_19602);
and UO_2246 (O_2246,N_19546,N_19830);
or UO_2247 (O_2247,N_19706,N_19714);
nand UO_2248 (O_2248,N_19926,N_19903);
or UO_2249 (O_2249,N_19692,N_19997);
or UO_2250 (O_2250,N_19641,N_19817);
or UO_2251 (O_2251,N_19742,N_19977);
or UO_2252 (O_2252,N_19552,N_19891);
and UO_2253 (O_2253,N_19858,N_19731);
nand UO_2254 (O_2254,N_19989,N_19606);
nand UO_2255 (O_2255,N_19868,N_19549);
nor UO_2256 (O_2256,N_19631,N_19623);
or UO_2257 (O_2257,N_19817,N_19660);
nor UO_2258 (O_2258,N_19862,N_19898);
or UO_2259 (O_2259,N_19985,N_19936);
xor UO_2260 (O_2260,N_19744,N_19787);
or UO_2261 (O_2261,N_19881,N_19671);
nor UO_2262 (O_2262,N_19559,N_19642);
xor UO_2263 (O_2263,N_19977,N_19997);
and UO_2264 (O_2264,N_19928,N_19783);
or UO_2265 (O_2265,N_19886,N_19922);
xor UO_2266 (O_2266,N_19556,N_19805);
xnor UO_2267 (O_2267,N_19941,N_19754);
nand UO_2268 (O_2268,N_19699,N_19878);
xnor UO_2269 (O_2269,N_19728,N_19591);
nand UO_2270 (O_2270,N_19554,N_19870);
or UO_2271 (O_2271,N_19677,N_19652);
and UO_2272 (O_2272,N_19947,N_19656);
or UO_2273 (O_2273,N_19517,N_19749);
nand UO_2274 (O_2274,N_19524,N_19927);
or UO_2275 (O_2275,N_19811,N_19665);
nand UO_2276 (O_2276,N_19609,N_19803);
and UO_2277 (O_2277,N_19753,N_19697);
or UO_2278 (O_2278,N_19949,N_19534);
and UO_2279 (O_2279,N_19829,N_19551);
nand UO_2280 (O_2280,N_19843,N_19544);
or UO_2281 (O_2281,N_19671,N_19729);
and UO_2282 (O_2282,N_19552,N_19542);
xor UO_2283 (O_2283,N_19946,N_19656);
nand UO_2284 (O_2284,N_19886,N_19821);
and UO_2285 (O_2285,N_19801,N_19998);
xor UO_2286 (O_2286,N_19564,N_19625);
xor UO_2287 (O_2287,N_19823,N_19637);
and UO_2288 (O_2288,N_19830,N_19849);
xor UO_2289 (O_2289,N_19843,N_19666);
and UO_2290 (O_2290,N_19582,N_19994);
nor UO_2291 (O_2291,N_19632,N_19862);
xor UO_2292 (O_2292,N_19672,N_19948);
xnor UO_2293 (O_2293,N_19803,N_19794);
xor UO_2294 (O_2294,N_19946,N_19674);
xor UO_2295 (O_2295,N_19727,N_19553);
xor UO_2296 (O_2296,N_19847,N_19797);
nand UO_2297 (O_2297,N_19992,N_19777);
or UO_2298 (O_2298,N_19817,N_19899);
and UO_2299 (O_2299,N_19632,N_19829);
nor UO_2300 (O_2300,N_19702,N_19821);
nand UO_2301 (O_2301,N_19560,N_19772);
nand UO_2302 (O_2302,N_19867,N_19749);
and UO_2303 (O_2303,N_19807,N_19677);
and UO_2304 (O_2304,N_19598,N_19731);
nand UO_2305 (O_2305,N_19639,N_19901);
and UO_2306 (O_2306,N_19774,N_19771);
or UO_2307 (O_2307,N_19940,N_19852);
nand UO_2308 (O_2308,N_19514,N_19823);
and UO_2309 (O_2309,N_19969,N_19759);
nand UO_2310 (O_2310,N_19885,N_19571);
or UO_2311 (O_2311,N_19723,N_19746);
nand UO_2312 (O_2312,N_19618,N_19804);
nor UO_2313 (O_2313,N_19615,N_19670);
and UO_2314 (O_2314,N_19773,N_19947);
xnor UO_2315 (O_2315,N_19547,N_19595);
xnor UO_2316 (O_2316,N_19699,N_19553);
xor UO_2317 (O_2317,N_19987,N_19614);
and UO_2318 (O_2318,N_19668,N_19990);
nand UO_2319 (O_2319,N_19976,N_19526);
or UO_2320 (O_2320,N_19832,N_19856);
nand UO_2321 (O_2321,N_19651,N_19905);
and UO_2322 (O_2322,N_19720,N_19669);
xor UO_2323 (O_2323,N_19574,N_19528);
and UO_2324 (O_2324,N_19656,N_19838);
nand UO_2325 (O_2325,N_19501,N_19658);
and UO_2326 (O_2326,N_19881,N_19876);
nand UO_2327 (O_2327,N_19708,N_19940);
and UO_2328 (O_2328,N_19682,N_19572);
and UO_2329 (O_2329,N_19703,N_19749);
or UO_2330 (O_2330,N_19931,N_19832);
or UO_2331 (O_2331,N_19756,N_19874);
or UO_2332 (O_2332,N_19604,N_19814);
nand UO_2333 (O_2333,N_19761,N_19506);
nor UO_2334 (O_2334,N_19766,N_19877);
nor UO_2335 (O_2335,N_19914,N_19557);
and UO_2336 (O_2336,N_19851,N_19882);
nand UO_2337 (O_2337,N_19526,N_19678);
nor UO_2338 (O_2338,N_19670,N_19866);
nor UO_2339 (O_2339,N_19863,N_19874);
xor UO_2340 (O_2340,N_19825,N_19940);
xor UO_2341 (O_2341,N_19729,N_19745);
or UO_2342 (O_2342,N_19963,N_19748);
xnor UO_2343 (O_2343,N_19621,N_19683);
or UO_2344 (O_2344,N_19720,N_19921);
nor UO_2345 (O_2345,N_19812,N_19693);
nor UO_2346 (O_2346,N_19572,N_19603);
or UO_2347 (O_2347,N_19836,N_19537);
nor UO_2348 (O_2348,N_19844,N_19980);
xnor UO_2349 (O_2349,N_19687,N_19690);
xor UO_2350 (O_2350,N_19638,N_19522);
nand UO_2351 (O_2351,N_19861,N_19566);
nand UO_2352 (O_2352,N_19863,N_19972);
nand UO_2353 (O_2353,N_19684,N_19662);
and UO_2354 (O_2354,N_19785,N_19542);
or UO_2355 (O_2355,N_19949,N_19683);
nand UO_2356 (O_2356,N_19599,N_19752);
or UO_2357 (O_2357,N_19538,N_19803);
xor UO_2358 (O_2358,N_19590,N_19621);
xnor UO_2359 (O_2359,N_19993,N_19515);
and UO_2360 (O_2360,N_19711,N_19853);
xnor UO_2361 (O_2361,N_19585,N_19505);
nor UO_2362 (O_2362,N_19855,N_19604);
nor UO_2363 (O_2363,N_19567,N_19764);
nand UO_2364 (O_2364,N_19794,N_19808);
and UO_2365 (O_2365,N_19724,N_19791);
or UO_2366 (O_2366,N_19506,N_19639);
or UO_2367 (O_2367,N_19838,N_19623);
nand UO_2368 (O_2368,N_19918,N_19969);
or UO_2369 (O_2369,N_19552,N_19674);
xnor UO_2370 (O_2370,N_19568,N_19720);
and UO_2371 (O_2371,N_19801,N_19887);
and UO_2372 (O_2372,N_19617,N_19819);
or UO_2373 (O_2373,N_19714,N_19531);
or UO_2374 (O_2374,N_19868,N_19691);
xor UO_2375 (O_2375,N_19825,N_19551);
and UO_2376 (O_2376,N_19636,N_19608);
nor UO_2377 (O_2377,N_19544,N_19647);
xnor UO_2378 (O_2378,N_19617,N_19817);
nor UO_2379 (O_2379,N_19552,N_19566);
nor UO_2380 (O_2380,N_19570,N_19876);
nor UO_2381 (O_2381,N_19857,N_19751);
xnor UO_2382 (O_2382,N_19771,N_19602);
xnor UO_2383 (O_2383,N_19517,N_19683);
nor UO_2384 (O_2384,N_19853,N_19787);
nand UO_2385 (O_2385,N_19925,N_19999);
nand UO_2386 (O_2386,N_19660,N_19947);
nor UO_2387 (O_2387,N_19919,N_19746);
xor UO_2388 (O_2388,N_19780,N_19782);
and UO_2389 (O_2389,N_19527,N_19526);
and UO_2390 (O_2390,N_19634,N_19639);
xnor UO_2391 (O_2391,N_19578,N_19967);
nand UO_2392 (O_2392,N_19877,N_19800);
nor UO_2393 (O_2393,N_19853,N_19790);
or UO_2394 (O_2394,N_19892,N_19734);
and UO_2395 (O_2395,N_19750,N_19691);
nand UO_2396 (O_2396,N_19873,N_19727);
or UO_2397 (O_2397,N_19865,N_19591);
nand UO_2398 (O_2398,N_19869,N_19945);
xnor UO_2399 (O_2399,N_19880,N_19552);
and UO_2400 (O_2400,N_19741,N_19717);
and UO_2401 (O_2401,N_19779,N_19953);
nand UO_2402 (O_2402,N_19842,N_19964);
xor UO_2403 (O_2403,N_19844,N_19508);
or UO_2404 (O_2404,N_19872,N_19661);
xor UO_2405 (O_2405,N_19804,N_19716);
or UO_2406 (O_2406,N_19987,N_19721);
nand UO_2407 (O_2407,N_19817,N_19795);
nor UO_2408 (O_2408,N_19843,N_19583);
nand UO_2409 (O_2409,N_19718,N_19987);
nor UO_2410 (O_2410,N_19846,N_19632);
nand UO_2411 (O_2411,N_19747,N_19846);
or UO_2412 (O_2412,N_19730,N_19712);
nand UO_2413 (O_2413,N_19594,N_19561);
xnor UO_2414 (O_2414,N_19930,N_19520);
or UO_2415 (O_2415,N_19558,N_19639);
or UO_2416 (O_2416,N_19617,N_19672);
or UO_2417 (O_2417,N_19709,N_19810);
nand UO_2418 (O_2418,N_19630,N_19748);
nand UO_2419 (O_2419,N_19999,N_19867);
and UO_2420 (O_2420,N_19936,N_19904);
or UO_2421 (O_2421,N_19520,N_19782);
and UO_2422 (O_2422,N_19802,N_19609);
nor UO_2423 (O_2423,N_19639,N_19821);
nand UO_2424 (O_2424,N_19544,N_19618);
xnor UO_2425 (O_2425,N_19885,N_19905);
xnor UO_2426 (O_2426,N_19988,N_19573);
or UO_2427 (O_2427,N_19989,N_19579);
and UO_2428 (O_2428,N_19783,N_19588);
nor UO_2429 (O_2429,N_19981,N_19956);
xnor UO_2430 (O_2430,N_19569,N_19712);
nor UO_2431 (O_2431,N_19780,N_19820);
nand UO_2432 (O_2432,N_19530,N_19735);
nor UO_2433 (O_2433,N_19646,N_19512);
nor UO_2434 (O_2434,N_19668,N_19928);
xnor UO_2435 (O_2435,N_19706,N_19973);
and UO_2436 (O_2436,N_19847,N_19834);
and UO_2437 (O_2437,N_19661,N_19836);
or UO_2438 (O_2438,N_19921,N_19572);
or UO_2439 (O_2439,N_19794,N_19562);
nor UO_2440 (O_2440,N_19689,N_19815);
xor UO_2441 (O_2441,N_19776,N_19607);
nor UO_2442 (O_2442,N_19734,N_19944);
or UO_2443 (O_2443,N_19919,N_19776);
nor UO_2444 (O_2444,N_19628,N_19779);
xor UO_2445 (O_2445,N_19684,N_19915);
xor UO_2446 (O_2446,N_19746,N_19834);
and UO_2447 (O_2447,N_19860,N_19700);
xor UO_2448 (O_2448,N_19707,N_19628);
nand UO_2449 (O_2449,N_19833,N_19867);
nor UO_2450 (O_2450,N_19583,N_19558);
and UO_2451 (O_2451,N_19791,N_19655);
xnor UO_2452 (O_2452,N_19706,N_19741);
and UO_2453 (O_2453,N_19729,N_19541);
nor UO_2454 (O_2454,N_19687,N_19552);
nor UO_2455 (O_2455,N_19529,N_19629);
nand UO_2456 (O_2456,N_19651,N_19525);
nand UO_2457 (O_2457,N_19549,N_19891);
xnor UO_2458 (O_2458,N_19972,N_19646);
or UO_2459 (O_2459,N_19798,N_19626);
nor UO_2460 (O_2460,N_19861,N_19992);
nand UO_2461 (O_2461,N_19716,N_19666);
nor UO_2462 (O_2462,N_19976,N_19603);
or UO_2463 (O_2463,N_19593,N_19506);
nand UO_2464 (O_2464,N_19738,N_19715);
and UO_2465 (O_2465,N_19845,N_19627);
nand UO_2466 (O_2466,N_19602,N_19705);
or UO_2467 (O_2467,N_19826,N_19523);
xor UO_2468 (O_2468,N_19742,N_19990);
nor UO_2469 (O_2469,N_19550,N_19580);
nand UO_2470 (O_2470,N_19649,N_19674);
or UO_2471 (O_2471,N_19760,N_19958);
or UO_2472 (O_2472,N_19767,N_19598);
xnor UO_2473 (O_2473,N_19986,N_19881);
xor UO_2474 (O_2474,N_19702,N_19688);
xnor UO_2475 (O_2475,N_19501,N_19867);
and UO_2476 (O_2476,N_19979,N_19670);
nor UO_2477 (O_2477,N_19926,N_19598);
nor UO_2478 (O_2478,N_19831,N_19846);
and UO_2479 (O_2479,N_19823,N_19613);
and UO_2480 (O_2480,N_19572,N_19737);
or UO_2481 (O_2481,N_19968,N_19525);
nor UO_2482 (O_2482,N_19595,N_19631);
and UO_2483 (O_2483,N_19836,N_19549);
or UO_2484 (O_2484,N_19613,N_19903);
nor UO_2485 (O_2485,N_19532,N_19852);
nand UO_2486 (O_2486,N_19742,N_19598);
and UO_2487 (O_2487,N_19886,N_19687);
xnor UO_2488 (O_2488,N_19721,N_19937);
nand UO_2489 (O_2489,N_19930,N_19990);
or UO_2490 (O_2490,N_19985,N_19975);
xor UO_2491 (O_2491,N_19924,N_19535);
nand UO_2492 (O_2492,N_19735,N_19549);
or UO_2493 (O_2493,N_19664,N_19667);
nand UO_2494 (O_2494,N_19823,N_19970);
or UO_2495 (O_2495,N_19565,N_19746);
or UO_2496 (O_2496,N_19747,N_19651);
nand UO_2497 (O_2497,N_19553,N_19606);
nand UO_2498 (O_2498,N_19986,N_19632);
xnor UO_2499 (O_2499,N_19564,N_19531);
endmodule