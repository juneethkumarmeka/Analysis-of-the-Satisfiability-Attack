module basic_1500_15000_2000_120_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_658,In_6);
nor U1 (N_1,In_1398,In_613);
nor U2 (N_2,In_413,In_639);
nor U3 (N_3,In_683,In_330);
or U4 (N_4,In_163,In_1050);
and U5 (N_5,In_1300,In_696);
and U6 (N_6,In_1177,In_582);
nor U7 (N_7,In_853,In_1296);
xnor U8 (N_8,In_1170,In_1469);
nand U9 (N_9,In_626,In_579);
or U10 (N_10,In_248,In_1373);
nor U11 (N_11,In_642,In_146);
or U12 (N_12,In_158,In_1429);
and U13 (N_13,In_1353,In_621);
nand U14 (N_14,In_741,In_1079);
nand U15 (N_15,In_58,In_299);
xor U16 (N_16,In_598,In_95);
and U17 (N_17,In_392,In_1083);
xor U18 (N_18,In_960,In_1007);
nand U19 (N_19,In_860,In_959);
and U20 (N_20,In_249,In_793);
and U21 (N_21,In_1198,In_1244);
and U22 (N_22,In_819,In_270);
nor U23 (N_23,In_457,In_878);
or U24 (N_24,In_1403,In_225);
and U25 (N_25,In_1009,In_1231);
nand U26 (N_26,In_665,In_992);
nand U27 (N_27,In_482,In_1037);
nand U28 (N_28,In_756,In_1217);
nand U29 (N_29,In_214,In_1492);
xnor U30 (N_30,In_564,In_1111);
xnor U31 (N_31,In_804,In_129);
and U32 (N_32,In_999,In_572);
or U33 (N_33,In_983,In_806);
and U34 (N_34,In_628,In_1033);
nand U35 (N_35,In_38,In_595);
xnor U36 (N_36,In_332,In_141);
and U37 (N_37,In_1116,In_339);
or U38 (N_38,In_153,In_1242);
xnor U39 (N_39,In_1268,In_1408);
or U40 (N_40,In_916,In_17);
nor U41 (N_41,In_865,In_986);
nand U42 (N_42,In_821,In_679);
nand U43 (N_43,In_401,In_1057);
or U44 (N_44,In_279,In_97);
nor U45 (N_45,In_1061,In_354);
nor U46 (N_46,In_767,In_874);
nor U47 (N_47,In_882,In_929);
nand U48 (N_48,In_1308,In_91);
and U49 (N_49,In_615,In_479);
or U50 (N_50,In_638,In_1128);
and U51 (N_51,In_1312,In_1490);
and U52 (N_52,In_750,In_801);
xor U53 (N_53,In_1072,In_1415);
nand U54 (N_54,In_773,In_728);
xnor U55 (N_55,In_967,In_89);
xor U56 (N_56,In_1091,In_757);
nor U57 (N_57,In_1291,In_28);
xnor U58 (N_58,In_216,In_527);
xor U59 (N_59,In_1342,In_1440);
nor U60 (N_60,In_969,In_1012);
or U61 (N_61,In_701,In_597);
xor U62 (N_62,In_996,In_1327);
nor U63 (N_63,In_1136,In_981);
nor U64 (N_64,In_453,In_165);
xnor U65 (N_65,In_934,In_124);
nand U66 (N_66,In_964,In_1101);
nor U67 (N_67,In_765,In_544);
or U68 (N_68,In_494,In_1393);
and U69 (N_69,In_654,In_939);
nand U70 (N_70,In_723,In_475);
xnor U71 (N_71,In_243,In_301);
nand U72 (N_72,In_811,In_541);
or U73 (N_73,In_478,In_891);
or U74 (N_74,In_218,In_651);
or U75 (N_75,In_1424,In_787);
nor U76 (N_76,In_1160,In_1224);
nor U77 (N_77,In_1391,In_114);
nor U78 (N_78,In_647,In_837);
or U79 (N_79,In_1234,In_1135);
and U80 (N_80,In_606,In_752);
nand U81 (N_81,In_1474,In_50);
or U82 (N_82,In_1051,In_602);
nor U83 (N_83,In_1431,In_1099);
nor U84 (N_84,In_1154,In_173);
and U85 (N_85,In_396,In_761);
xor U86 (N_86,In_1064,In_23);
and U87 (N_87,In_438,In_1069);
or U88 (N_88,In_1229,In_943);
and U89 (N_89,In_545,In_716);
xor U90 (N_90,In_1321,In_283);
or U91 (N_91,In_1301,In_603);
xnor U92 (N_92,In_697,In_1476);
nand U93 (N_93,In_1416,In_502);
xor U94 (N_94,In_1378,In_167);
nand U95 (N_95,In_390,In_805);
and U96 (N_96,In_319,In_184);
nand U97 (N_97,In_858,In_1281);
or U98 (N_98,In_1106,In_281);
xor U99 (N_99,In_357,In_3);
nand U100 (N_100,In_1481,In_133);
xor U101 (N_101,In_818,In_1288);
nand U102 (N_102,In_1274,In_1248);
nand U103 (N_103,In_292,In_557);
and U104 (N_104,In_220,In_61);
nand U105 (N_105,In_12,In_901);
xnor U106 (N_106,In_1212,In_1131);
and U107 (N_107,In_1144,In_1376);
and U108 (N_108,In_1386,In_1112);
xnor U109 (N_109,In_1200,In_109);
nor U110 (N_110,In_331,In_103);
and U111 (N_111,In_7,In_1361);
and U112 (N_112,In_1280,In_508);
or U113 (N_113,In_927,In_1232);
and U114 (N_114,In_113,In_1210);
xor U115 (N_115,In_18,In_576);
or U116 (N_116,In_736,In_873);
nand U117 (N_117,In_1412,In_172);
and U118 (N_118,In_1038,In_329);
or U119 (N_119,In_1120,In_1040);
nor U120 (N_120,In_1117,In_1314);
and U121 (N_121,In_549,In_600);
or U122 (N_122,In_31,In_1467);
and U123 (N_123,In_727,In_136);
or U124 (N_124,In_1263,In_1086);
nand U125 (N_125,In_8,In_719);
or U126 (N_126,In_143,In_1203);
xor U127 (N_127,In_190,In_536);
nor U128 (N_128,In_671,In_646);
or U129 (N_129,In_180,N_60);
and U130 (N_130,In_1137,N_122);
nor U131 (N_131,In_42,In_64);
or U132 (N_132,In_66,In_238);
nand U133 (N_133,In_952,In_1145);
nand U134 (N_134,N_120,In_925);
or U135 (N_135,In_1381,N_48);
xor U136 (N_136,N_105,In_1031);
or U137 (N_137,In_1433,In_257);
nor U138 (N_138,In_1186,In_786);
xnor U139 (N_139,In_1324,In_295);
nor U140 (N_140,In_569,In_1097);
or U141 (N_141,In_310,In_490);
xnor U142 (N_142,In_643,In_680);
nand U143 (N_143,In_99,In_1284);
or U144 (N_144,In_90,In_49);
and U145 (N_145,In_1310,In_1077);
and U146 (N_146,In_1347,N_99);
and U147 (N_147,In_930,In_16);
nand U148 (N_148,In_624,In_152);
or U149 (N_149,In_868,In_1441);
nor U150 (N_150,In_78,In_1143);
nand U151 (N_151,In_970,In_21);
nand U152 (N_152,In_1294,In_459);
nand U153 (N_153,In_704,In_1426);
or U154 (N_154,In_915,In_754);
nand U155 (N_155,In_1205,In_935);
xnor U156 (N_156,In_1055,In_116);
xnor U157 (N_157,In_991,In_619);
nand U158 (N_158,In_524,N_51);
nor U159 (N_159,In_486,In_179);
xor U160 (N_160,In_1082,In_135);
xor U161 (N_161,In_1382,In_356);
and U162 (N_162,In_749,In_217);
xnor U163 (N_163,In_588,N_91);
xor U164 (N_164,In_1350,In_1236);
nor U165 (N_165,In_393,In_233);
xor U166 (N_166,In_127,In_107);
or U167 (N_167,In_869,In_1427);
xor U168 (N_168,In_327,In_1283);
or U169 (N_169,In_1161,In_1222);
xor U170 (N_170,In_487,In_1417);
nor U171 (N_171,In_239,In_1233);
xnor U172 (N_172,N_67,N_78);
xor U173 (N_173,N_92,N_79);
nor U174 (N_174,In_705,In_1275);
or U175 (N_175,In_556,In_192);
and U176 (N_176,In_34,In_269);
or U177 (N_177,In_976,In_795);
and U178 (N_178,In_779,N_36);
xnor U179 (N_179,In_790,In_1206);
or U180 (N_180,In_1325,In_601);
and U181 (N_181,In_1108,In_1109);
and U182 (N_182,N_101,In_698);
xor U183 (N_183,In_1435,In_1052);
xnor U184 (N_184,In_209,In_961);
xnor U185 (N_185,In_221,In_540);
or U186 (N_186,In_1346,In_825);
nand U187 (N_187,In_778,In_315);
or U188 (N_188,In_721,N_40);
nand U189 (N_189,In_594,In_1219);
or U190 (N_190,In_980,In_1389);
xor U191 (N_191,In_280,In_810);
nand U192 (N_192,In_692,N_44);
xor U193 (N_193,In_1022,In_1436);
xor U194 (N_194,In_1498,In_670);
nor U195 (N_195,In_1025,In_1479);
xnor U196 (N_196,In_1497,In_1228);
nor U197 (N_197,In_481,In_872);
nand U198 (N_198,In_1317,In_691);
xor U199 (N_199,In_590,In_896);
and U200 (N_200,In_1473,In_988);
xor U201 (N_201,In_84,In_1029);
and U202 (N_202,In_79,In_489);
or U203 (N_203,In_178,In_794);
nand U204 (N_204,In_379,In_561);
nor U205 (N_205,In_465,In_194);
nand U206 (N_206,In_436,In_1377);
or U207 (N_207,In_1085,In_971);
nand U208 (N_208,In_312,In_1053);
and U209 (N_209,In_11,In_206);
and U210 (N_210,In_13,In_592);
xor U211 (N_211,In_1194,In_875);
nor U212 (N_212,In_1460,N_115);
and U213 (N_213,In_1311,In_408);
and U214 (N_214,In_1100,In_372);
or U215 (N_215,In_797,In_854);
nand U216 (N_216,In_525,In_147);
or U217 (N_217,In_430,In_1295);
and U218 (N_218,In_318,In_1);
xnor U219 (N_219,In_110,In_1454);
xor U220 (N_220,In_429,In_965);
and U221 (N_221,In_844,In_1028);
nand U222 (N_222,In_325,In_1343);
nor U223 (N_223,In_231,In_566);
and U224 (N_224,In_448,N_56);
xnor U225 (N_225,In_345,In_1179);
or U226 (N_226,In_563,In_1098);
nor U227 (N_227,In_669,In_1258);
nor U228 (N_228,In_884,N_47);
xor U229 (N_229,In_958,In_899);
or U230 (N_230,In_1419,In_102);
nor U231 (N_231,In_87,N_106);
and U232 (N_232,In_689,In_953);
xor U233 (N_233,In_311,In_962);
and U234 (N_234,In_1046,In_195);
xnor U235 (N_235,In_1392,In_1169);
xnor U236 (N_236,In_1035,In_1306);
and U237 (N_237,In_738,In_883);
nand U238 (N_238,In_1036,N_22);
or U239 (N_239,In_1411,In_1193);
nand U240 (N_240,In_505,In_451);
nor U241 (N_241,In_843,In_725);
nor U242 (N_242,N_35,In_1148);
and U243 (N_243,In_522,In_904);
nand U244 (N_244,In_1013,In_321);
nor U245 (N_245,In_1142,In_575);
xor U246 (N_246,In_1304,In_1071);
or U247 (N_247,In_921,In_48);
nand U248 (N_248,In_788,In_998);
nand U249 (N_249,In_1379,In_1214);
nand U250 (N_250,N_80,In_517);
nor U251 (N_251,In_1450,N_82);
and U252 (N_252,In_931,In_973);
or U253 (N_253,In_352,In_1276);
or U254 (N_254,N_194,In_610);
xor U255 (N_255,In_52,In_1113);
nand U256 (N_256,In_63,In_1024);
or U257 (N_257,In_807,In_423);
xor U258 (N_258,In_403,In_75);
xnor U259 (N_259,In_397,In_866);
xor U260 (N_260,In_1124,In_622);
or U261 (N_261,In_497,N_141);
xor U262 (N_262,In_1430,In_1380);
and U263 (N_263,In_417,In_743);
xnor U264 (N_264,In_236,N_232);
and U265 (N_265,In_171,N_157);
and U266 (N_266,In_1059,In_1437);
and U267 (N_267,In_938,In_842);
nand U268 (N_268,In_630,In_956);
nor U269 (N_269,In_957,In_870);
and U270 (N_270,In_338,In_228);
nand U271 (N_271,In_1330,In_942);
and U272 (N_272,In_532,In_360);
nand U273 (N_273,N_153,In_1388);
or U274 (N_274,In_121,In_1063);
or U275 (N_275,In_997,In_302);
or U276 (N_276,In_745,In_2);
xnor U277 (N_277,In_1039,In_586);
or U278 (N_278,In_1484,N_202);
nand U279 (N_279,In_1404,In_1215);
nor U280 (N_280,In_1282,N_11);
nand U281 (N_281,In_1319,In_923);
and U282 (N_282,In_452,N_112);
nor U283 (N_283,In_1332,In_207);
nand U284 (N_284,In_1104,In_80);
or U285 (N_285,In_72,N_0);
and U286 (N_286,N_94,In_758);
or U287 (N_287,In_335,In_36);
or U288 (N_288,N_185,N_4);
nor U289 (N_289,In_1309,In_693);
nand U290 (N_290,In_568,In_333);
and U291 (N_291,N_224,In_1259);
nand U292 (N_292,In_782,In_104);
nor U293 (N_293,N_178,In_1463);
nand U294 (N_294,In_241,In_714);
nand U295 (N_295,In_1365,In_531);
or U296 (N_296,N_111,In_251);
nor U297 (N_297,N_162,In_898);
nor U298 (N_298,In_106,In_286);
nor U299 (N_299,In_1105,In_317);
nand U300 (N_300,N_179,In_373);
or U301 (N_301,N_192,N_170);
xor U302 (N_302,In_128,In_663);
nand U303 (N_303,In_1209,In_328);
nor U304 (N_304,In_294,In_1188);
or U305 (N_305,In_1394,N_93);
nor U306 (N_306,In_421,N_156);
and U307 (N_307,In_130,In_1181);
nor U308 (N_308,In_378,In_336);
nor U309 (N_309,In_746,In_368);
or U310 (N_310,In_1357,In_1223);
nor U311 (N_311,In_56,In_156);
and U312 (N_312,In_777,In_274);
xor U313 (N_313,In_140,In_924);
or U314 (N_314,In_1241,In_82);
and U315 (N_315,In_712,N_34);
xor U316 (N_316,N_88,In_644);
or U317 (N_317,N_247,In_289);
or U318 (N_318,In_781,In_1269);
and U319 (N_319,N_116,N_16);
nor U320 (N_320,In_911,In_1134);
or U321 (N_321,In_1164,In_96);
and U322 (N_322,N_113,In_968);
xnor U323 (N_323,In_1066,In_839);
or U324 (N_324,In_578,In_191);
nand U325 (N_325,In_445,N_37);
and U326 (N_326,In_1218,In_1151);
xnor U327 (N_327,In_1189,In_1487);
or U328 (N_328,In_1414,In_933);
and U329 (N_329,In_43,In_1102);
or U330 (N_330,In_1445,In_1413);
and U331 (N_331,In_537,N_72);
xor U332 (N_332,In_612,In_366);
or U333 (N_333,In_1466,In_1364);
or U334 (N_334,In_288,In_247);
or U335 (N_335,In_166,In_659);
nor U336 (N_336,In_1140,In_1010);
nor U337 (N_337,In_1251,In_304);
and U338 (N_338,In_1322,In_690);
and U339 (N_339,In_637,In_599);
nor U340 (N_340,In_1023,In_735);
nor U341 (N_341,In_1422,N_139);
xnor U342 (N_342,In_1340,In_162);
xor U343 (N_343,N_155,In_365);
nand U344 (N_344,In_155,In_941);
nor U345 (N_345,In_1348,In_1485);
nor U346 (N_346,In_272,In_1246);
or U347 (N_347,In_905,In_694);
or U348 (N_348,N_61,In_803);
nor U349 (N_349,N_96,N_30);
nor U350 (N_350,In_1183,In_1461);
nand U351 (N_351,In_908,N_239);
nand U352 (N_352,In_1420,In_1049);
nor U353 (N_353,N_241,In_33);
or U354 (N_354,In_1173,N_121);
nor U355 (N_355,N_89,In_1305);
and U356 (N_356,In_1434,In_1265);
nand U357 (N_357,In_616,N_210);
xor U358 (N_358,In_1355,In_261);
and U359 (N_359,In_729,In_1480);
nand U360 (N_360,In_1096,In_695);
or U361 (N_361,In_5,In_881);
xor U362 (N_362,In_850,In_9);
and U363 (N_363,N_223,In_341);
nor U364 (N_364,N_124,In_709);
nor U365 (N_365,N_6,In_142);
or U366 (N_366,In_554,N_46);
nor U367 (N_367,N_220,In_731);
xnor U368 (N_368,In_355,In_664);
nor U369 (N_369,In_343,In_168);
nand U370 (N_370,N_50,In_60);
xnor U371 (N_371,In_210,N_3);
nor U372 (N_372,In_203,In_149);
and U373 (N_373,In_204,In_1299);
and U374 (N_374,In_937,In_101);
nor U375 (N_375,In_47,In_230);
xor U376 (N_376,In_859,In_1146);
xor U377 (N_377,In_672,In_182);
xnor U378 (N_378,In_65,In_170);
nand U379 (N_379,In_657,In_1176);
nand U380 (N_380,N_309,In_383);
or U381 (N_381,In_1043,N_317);
and U382 (N_382,N_137,N_312);
xnor U383 (N_383,In_1180,In_1175);
or U384 (N_384,N_69,In_323);
or U385 (N_385,In_287,N_266);
xnor U386 (N_386,N_356,N_358);
nand U387 (N_387,In_558,N_38);
nand U388 (N_388,In_57,In_1192);
nor U389 (N_389,In_822,In_635);
or U390 (N_390,In_1432,In_836);
and U391 (N_391,In_528,In_668);
or U392 (N_392,N_74,In_951);
nand U393 (N_393,In_414,In_235);
nor U394 (N_394,In_268,In_450);
xnor U395 (N_395,In_1326,In_334);
nand U396 (N_396,In_151,In_1499);
nor U397 (N_397,N_372,In_1163);
xnor U398 (N_398,N_62,N_12);
xnor U399 (N_399,N_349,In_1323);
xor U400 (N_400,N_234,In_1115);
xnor U401 (N_401,In_1496,N_190);
xnor U402 (N_402,In_296,In_1338);
xor U403 (N_403,In_660,In_208);
nor U404 (N_404,In_1328,In_985);
nor U405 (N_405,In_254,In_812);
nor U406 (N_406,N_327,N_332);
and U407 (N_407,In_783,In_1008);
and U408 (N_408,N_254,In_92);
and U409 (N_409,In_174,In_666);
nand U410 (N_410,In_1453,In_420);
nand U411 (N_411,In_1132,In_1261);
nand U412 (N_412,In_1020,In_539);
and U413 (N_413,In_1399,N_117);
nand U414 (N_414,In_380,In_1447);
or U415 (N_415,N_291,N_201);
nor U416 (N_416,In_1087,In_1114);
and U417 (N_417,In_1088,In_1272);
or U418 (N_418,In_353,In_1019);
and U419 (N_419,In_538,In_340);
xor U420 (N_420,In_909,N_335);
nor U421 (N_421,N_322,In_205);
nor U422 (N_422,N_203,In_455);
xor U423 (N_423,In_1245,In_840);
nand U424 (N_424,In_677,N_213);
nor U425 (N_425,In_1307,In_1329);
nand U426 (N_426,In_1290,In_1092);
nor U427 (N_427,In_808,In_316);
nand U428 (N_428,In_369,In_351);
nor U429 (N_429,In_444,N_365);
nor U430 (N_430,In_662,In_838);
nor U431 (N_431,In_389,In_1237);
and U432 (N_432,In_447,In_890);
nand U433 (N_433,In_1093,In_201);
nor U434 (N_434,In_1253,In_722);
nand U435 (N_435,In_1138,N_215);
or U436 (N_436,In_226,N_21);
xor U437 (N_437,N_147,In_526);
nor U438 (N_438,In_1400,N_299);
and U439 (N_439,In_54,In_553);
nor U440 (N_440,In_100,N_20);
and U441 (N_441,In_1320,In_1375);
or U442 (N_442,In_181,In_1060);
nand U443 (N_443,In_887,N_175);
xor U444 (N_444,In_1358,N_166);
nand U445 (N_445,In_1333,In_77);
nor U446 (N_446,In_346,In_892);
nand U447 (N_447,In_880,In_25);
nor U448 (N_448,In_211,N_219);
or U449 (N_449,In_867,In_1211);
nand U450 (N_450,In_632,In_454);
and U451 (N_451,In_1153,In_720);
nand U452 (N_452,In_667,In_963);
xor U453 (N_453,N_136,In_744);
and U454 (N_454,In_88,In_337);
xnor U455 (N_455,In_1047,In_83);
nand U456 (N_456,In_894,In_1493);
and U457 (N_457,N_297,N_333);
xor U458 (N_458,In_1107,In_715);
nor U459 (N_459,In_1159,In_1452);
and U460 (N_460,In_1150,In_920);
or U461 (N_461,In_1383,In_548);
nand U462 (N_462,In_199,In_1407);
nand U463 (N_463,N_250,In_984);
or U464 (N_464,In_1011,In_223);
nor U465 (N_465,In_955,In_948);
xnor U466 (N_466,In_385,In_814);
or U467 (N_467,N_285,In_358);
and U468 (N_468,N_158,N_261);
xnor U469 (N_469,In_0,In_1345);
and U470 (N_470,N_143,In_753);
xor U471 (N_471,N_65,N_351);
nor U472 (N_472,In_1336,In_1001);
or U473 (N_473,In_717,In_1014);
and U474 (N_474,N_361,N_237);
or U475 (N_475,N_9,In_183);
and U476 (N_476,In_885,In_845);
or U477 (N_477,In_132,N_97);
xnor U478 (N_478,N_154,N_128);
nand U479 (N_479,In_416,In_51);
nand U480 (N_480,In_766,In_802);
xnor U481 (N_481,N_58,In_888);
xnor U482 (N_482,In_833,N_95);
or U483 (N_483,In_918,In_111);
nor U484 (N_484,N_330,In_222);
nand U485 (N_485,In_418,N_228);
xnor U486 (N_486,In_1235,In_219);
and U487 (N_487,In_907,In_1318);
xor U488 (N_488,In_462,In_398);
xor U489 (N_489,In_30,In_1225);
nand U490 (N_490,In_1352,In_134);
and U491 (N_491,In_409,N_264);
nor U492 (N_492,In_584,N_320);
nand U493 (N_493,In_580,In_1239);
and U494 (N_494,In_1483,N_318);
or U495 (N_495,In_405,In_1495);
nand U496 (N_496,In_824,In_510);
nor U497 (N_497,N_133,In_402);
xor U498 (N_498,In_857,In_22);
or U499 (N_499,In_1126,In_1185);
nor U500 (N_500,In_734,In_1468);
and U501 (N_501,N_464,N_319);
xor U502 (N_502,N_315,N_440);
xnor U503 (N_503,In_1162,In_625);
nor U504 (N_504,In_523,In_1368);
nand U505 (N_505,N_406,In_466);
and U506 (N_506,In_574,In_1339);
or U507 (N_507,In_125,In_687);
nand U508 (N_508,N_8,In_1015);
nor U509 (N_509,In_1006,N_480);
and U510 (N_510,N_403,N_290);
xor U511 (N_511,In_1397,In_45);
and U512 (N_512,N_359,In_760);
nor U513 (N_513,In_1062,In_587);
and U514 (N_514,In_186,In_1457);
nor U515 (N_515,N_212,N_103);
nand U516 (N_516,N_308,In_76);
and U517 (N_517,N_416,N_214);
nor U518 (N_518,In_108,N_422);
xnor U519 (N_519,In_1158,In_1488);
nor U520 (N_520,In_1075,N_476);
nand U521 (N_521,N_345,N_249);
xnor U522 (N_522,N_145,In_1298);
or U523 (N_523,In_177,N_126);
nand U524 (N_524,In_533,In_1448);
or U525 (N_525,N_53,N_395);
or U526 (N_526,N_364,In_276);
nor U527 (N_527,N_243,In_950);
nand U528 (N_528,In_370,In_258);
and U529 (N_529,N_230,In_460);
or U530 (N_530,N_32,In_498);
xnor U531 (N_531,In_796,In_145);
nand U532 (N_532,N_373,N_159);
xor U533 (N_533,In_1384,In_253);
or U534 (N_534,N_176,In_684);
nor U535 (N_535,In_1471,In_193);
and U536 (N_536,N_437,In_1313);
or U537 (N_537,In_1442,In_431);
nor U538 (N_538,N_468,N_174);
and U539 (N_539,N_397,N_90);
and U540 (N_540,In_303,In_994);
nor U541 (N_541,In_458,N_409);
nor U542 (N_542,N_251,N_235);
or U543 (N_543,N_54,In_1171);
nand U544 (N_544,In_1302,In_604);
nand U545 (N_545,N_13,In_1167);
nor U546 (N_546,In_1080,N_180);
nor U547 (N_547,In_188,In_1000);
and U548 (N_548,In_900,N_102);
and U549 (N_549,In_242,In_1270);
xnor U550 (N_550,In_39,N_483);
xor U551 (N_551,In_271,In_813);
or U552 (N_552,In_618,In_1199);
xor U553 (N_553,In_161,In_771);
nand U554 (N_554,N_191,In_856);
nor U555 (N_555,In_897,In_895);
nor U556 (N_556,N_370,In_267);
xnor U557 (N_557,N_281,In_1285);
and U558 (N_558,N_296,N_19);
nor U559 (N_559,In_1273,N_233);
xnor U560 (N_560,In_1267,In_1045);
nand U561 (N_561,In_435,In_196);
xor U562 (N_562,In_410,In_1152);
nor U563 (N_563,In_1425,In_1084);
nor U564 (N_564,In_424,In_426);
and U565 (N_565,In_1094,In_852);
nand U566 (N_566,N_336,In_1002);
and U567 (N_567,N_274,N_497);
xnor U568 (N_568,In_979,In_1456);
nor U569 (N_569,N_418,In_627);
or U570 (N_570,In_726,In_742);
or U571 (N_571,N_45,In_1250);
or U572 (N_572,In_641,In_1367);
or U573 (N_573,In_86,In_636);
nor U574 (N_574,N_490,N_119);
xor U575 (N_575,N_426,In_93);
or U576 (N_576,N_59,In_1195);
nor U577 (N_577,In_1477,N_184);
nor U578 (N_578,In_944,N_391);
nor U579 (N_579,In_367,N_301);
xnor U580 (N_580,N_189,N_377);
nand U581 (N_581,In_1279,In_138);
nand U582 (N_582,N_340,In_946);
nor U583 (N_583,In_648,In_617);
nand U584 (N_584,In_144,In_551);
or U585 (N_585,N_366,In_535);
or U586 (N_586,In_326,In_543);
or U587 (N_587,In_1410,In_608);
xor U588 (N_588,In_496,N_262);
or U589 (N_589,In_1459,N_458);
nor U590 (N_590,N_456,N_294);
xor U591 (N_591,In_449,In_987);
and U592 (N_592,N_27,In_1395);
nand U593 (N_593,In_798,In_581);
or U594 (N_594,In_686,In_94);
nor U595 (N_595,N_66,N_324);
or U596 (N_596,N_494,In_1074);
nor U597 (N_597,N_486,N_369);
nor U598 (N_598,In_425,In_491);
and U599 (N_599,In_768,In_966);
xor U600 (N_600,N_415,N_218);
and U601 (N_601,In_759,N_475);
or U602 (N_602,In_480,In_376);
nand U603 (N_603,In_262,In_772);
nand U604 (N_604,N_77,In_815);
xnor U605 (N_605,N_380,In_297);
or U606 (N_606,N_432,N_187);
or U607 (N_607,N_289,In_855);
xnor U608 (N_608,In_675,N_221);
or U609 (N_609,In_1182,N_360);
xor U610 (N_610,N_75,In_775);
xnor U611 (N_611,N_33,N_114);
or U612 (N_612,N_181,N_204);
or U613 (N_613,N_73,In_433);
nand U614 (N_614,In_730,In_1359);
nor U615 (N_615,N_407,N_2);
and U616 (N_616,In_1004,N_164);
and U617 (N_617,N_334,In_1125);
or U618 (N_618,In_849,In_309);
nand U619 (N_619,In_278,N_118);
nand U620 (N_620,In_513,N_492);
nor U621 (N_621,In_1402,N_193);
nor U622 (N_622,In_412,N_208);
and U623 (N_623,N_255,In_1127);
nand U624 (N_624,N_286,In_559);
nor U625 (N_625,In_1065,N_507);
nor U626 (N_626,N_502,N_580);
nand U627 (N_627,In_546,In_293);
nand U628 (N_628,In_650,In_347);
nor U629 (N_629,In_506,In_44);
nor U630 (N_630,In_263,N_487);
xnor U631 (N_631,N_561,In_893);
nor U632 (N_632,N_599,N_31);
nand U633 (N_633,N_229,In_1409);
and U634 (N_634,In_661,In_55);
xnor U635 (N_635,In_391,In_164);
xor U636 (N_636,In_977,N_347);
xnor U637 (N_637,In_917,In_831);
xor U638 (N_638,In_567,In_515);
and U639 (N_639,In_847,N_399);
and U640 (N_640,In_381,In_1252);
nor U641 (N_641,N_588,In_415);
nor U642 (N_642,In_774,In_154);
nand U643 (N_643,N_142,N_379);
or U644 (N_644,In_298,In_820);
nor U645 (N_645,N_248,In_947);
or U646 (N_646,In_1130,In_1216);
nor U647 (N_647,In_547,In_1129);
nor U648 (N_648,N_107,N_275);
nand U649 (N_649,In_562,N_410);
nand U650 (N_650,In_780,In_1354);
nand U651 (N_651,N_138,N_413);
nand U652 (N_652,N_18,N_443);
nor U653 (N_653,In_1254,In_1462);
and U654 (N_654,N_337,In_737);
nand U655 (N_655,N_169,N_591);
or U656 (N_656,N_477,In_1073);
xor U657 (N_657,In_240,In_711);
nand U658 (N_658,N_165,N_537);
xnor U659 (N_659,N_535,In_864);
and U660 (N_660,In_1118,In_1472);
xnor U661 (N_661,N_425,N_384);
nor U662 (N_662,In_792,N_402);
nand U663 (N_663,In_322,In_1190);
nor U664 (N_664,N_260,In_148);
nand U665 (N_665,In_583,N_421);
nand U666 (N_666,In_374,In_1451);
nand U667 (N_667,N_423,In_1048);
and U668 (N_668,In_1478,In_464);
xor U669 (N_669,In_364,N_198);
xor U670 (N_670,N_167,N_374);
nor U671 (N_671,N_196,In_359);
or U672 (N_672,N_355,In_1489);
and U673 (N_673,N_508,In_800);
and U674 (N_674,In_645,In_349);
or U675 (N_675,In_1271,In_1165);
and U676 (N_676,N_595,In_443);
or U677 (N_677,In_634,In_1221);
nand U678 (N_678,N_300,N_600);
xor U679 (N_679,In_542,N_527);
or U680 (N_680,In_629,In_876);
xnor U681 (N_681,In_256,In_406);
nand U682 (N_682,N_552,In_676);
nor U683 (N_683,In_1157,In_382);
and U684 (N_684,N_608,N_479);
and U685 (N_685,In_473,In_990);
and U686 (N_686,N_560,N_323);
or U687 (N_687,N_49,N_514);
and U688 (N_688,N_515,N_311);
or U689 (N_689,N_63,N_448);
xnor U690 (N_690,In_1089,In_1362);
or U691 (N_691,N_87,In_98);
and U692 (N_692,N_460,In_19);
or U693 (N_693,In_972,In_189);
nor U694 (N_694,In_1034,N_217);
nor U695 (N_695,N_550,In_555);
xnor U696 (N_696,In_700,In_620);
nand U697 (N_697,N_427,In_573);
or U698 (N_698,N_417,N_506);
nand U699 (N_699,N_467,N_23);
and U700 (N_700,In_1374,In_41);
nor U701 (N_701,In_591,In_685);
nor U702 (N_702,N_378,In_126);
xnor U703 (N_703,N_564,N_452);
nand U704 (N_704,N_368,In_1369);
nor U705 (N_705,N_433,In_265);
or U706 (N_706,In_259,N_123);
and U707 (N_707,In_1446,N_125);
nand U708 (N_708,N_522,In_308);
nand U709 (N_709,In_266,In_495);
xnor U710 (N_710,In_589,In_512);
or U711 (N_711,N_55,In_889);
nand U712 (N_712,In_740,In_1204);
nor U713 (N_713,N_270,In_1070);
and U714 (N_714,In_974,In_1444);
or U715 (N_715,In_785,In_863);
nor U716 (N_716,N_258,In_1372);
xnor U717 (N_717,In_260,In_120);
or U718 (N_718,N_496,In_910);
xnor U719 (N_719,In_518,N_617);
nor U720 (N_720,In_46,In_1486);
nand U721 (N_721,In_707,In_832);
nand U722 (N_722,N_404,N_576);
nand U723 (N_723,In_879,N_493);
nor U724 (N_724,N_543,In_234);
and U725 (N_725,In_74,N_615);
or U726 (N_726,N_41,In_1149);
or U727 (N_727,N_57,In_789);
and U728 (N_728,N_100,N_70);
xnor U729 (N_729,N_148,N_24);
and U730 (N_730,N_15,N_485);
xor U731 (N_731,In_1438,In_10);
nand U732 (N_732,N_548,N_259);
nor U733 (N_733,N_521,N_471);
nand U734 (N_734,N_435,In_1119);
and U735 (N_735,N_240,N_549);
or U736 (N_736,N_280,N_242);
and U737 (N_737,In_1191,N_499);
or U738 (N_738,N_400,In_485);
or U739 (N_739,In_399,N_144);
xor U740 (N_740,In_1041,N_593);
or U741 (N_741,In_593,N_444);
or U742 (N_742,In_68,In_1370);
xor U743 (N_743,In_476,In_428);
and U744 (N_744,In_131,In_1076);
xnor U745 (N_745,In_1187,In_229);
nor U746 (N_746,In_769,In_1405);
or U747 (N_747,In_1363,N_621);
and U748 (N_748,N_195,N_434);
nand U749 (N_749,In_688,N_350);
or U750 (N_750,N_713,N_287);
nand U751 (N_751,In_710,N_558);
nand U752 (N_752,In_1385,In_1390);
nand U753 (N_753,N_183,N_577);
and U754 (N_754,In_463,N_545);
nor U755 (N_755,In_1054,N_161);
or U756 (N_756,In_200,N_83);
nor U757 (N_757,In_1078,N_629);
and U758 (N_758,N_700,N_706);
xor U759 (N_759,N_282,In_112);
or U760 (N_760,N_446,N_721);
xor U761 (N_761,In_1044,N_689);
and U762 (N_762,N_455,In_273);
nor U763 (N_763,N_719,In_649);
or U764 (N_764,N_671,In_509);
or U765 (N_765,In_1418,In_15);
nand U766 (N_766,N_715,In_954);
nor U767 (N_767,In_791,N_517);
or U768 (N_768,N_424,N_728);
nor U769 (N_769,N_696,N_723);
and U770 (N_770,N_441,In_137);
and U771 (N_771,N_343,N_470);
and U772 (N_772,N_542,N_134);
or U773 (N_773,In_1166,N_694);
nand U774 (N_774,In_1032,N_466);
and U775 (N_775,N_386,In_1335);
xor U776 (N_776,In_848,N_619);
nand U777 (N_777,In_747,In_1255);
and U778 (N_778,In_71,N_495);
and U779 (N_779,In_1068,N_693);
nor U780 (N_780,N_565,In_936);
nor U781 (N_781,N_686,N_546);
or U782 (N_782,In_1421,N_581);
nand U783 (N_783,N_236,N_431);
nor U784 (N_784,N_705,N_626);
xor U785 (N_785,N_151,N_707);
nand U786 (N_786,N_303,N_643);
or U787 (N_787,N_573,N_246);
and U788 (N_788,In_724,In_255);
or U789 (N_789,N_271,In_400);
or U790 (N_790,In_81,N_459);
nor U791 (N_791,N_316,In_1016);
nor U792 (N_792,N_676,In_442);
nand U793 (N_793,In_411,In_115);
nor U794 (N_794,N_536,N_607);
and U795 (N_795,N_163,N_314);
and U796 (N_796,In_1387,In_27);
and U797 (N_797,In_784,In_232);
and U798 (N_798,N_457,N_729);
and U799 (N_799,N_520,In_290);
nor U800 (N_800,In_928,In_926);
and U801 (N_801,In_678,N_367);
nor U802 (N_802,In_1458,N_653);
or U803 (N_803,In_62,In_157);
or U804 (N_804,N_630,In_823);
and U805 (N_805,N_722,In_834);
or U806 (N_806,In_53,N_673);
nand U807 (N_807,N_108,N_748);
and U808 (N_808,N_265,In_1406);
or U809 (N_809,N_461,N_698);
or U810 (N_810,N_357,In_1331);
xor U811 (N_811,N_503,N_484);
nor U812 (N_812,N_257,N_478);
nor U813 (N_813,N_528,N_746);
xnor U814 (N_814,N_569,In_596);
xnor U815 (N_815,In_440,In_1133);
or U816 (N_816,In_456,In_1464);
or U817 (N_817,In_176,In_520);
nor U818 (N_818,In_762,In_565);
and U819 (N_819,In_1443,In_1201);
or U820 (N_820,In_982,N_669);
or U821 (N_821,N_375,In_732);
xor U822 (N_822,In_1156,N_633);
and U823 (N_823,N_346,In_653);
nand U824 (N_824,N_530,In_446);
and U825 (N_825,In_534,In_1018);
and U826 (N_826,In_488,N_329);
xor U827 (N_827,In_764,In_1396);
nor U828 (N_828,N_606,N_526);
and U829 (N_829,N_616,N_579);
and U830 (N_830,In_324,In_300);
or U831 (N_831,In_160,N_740);
nor U832 (N_832,N_640,N_587);
nor U833 (N_833,N_701,In_407);
nand U834 (N_834,In_978,N_547);
or U835 (N_835,In_529,N_389);
nor U836 (N_836,N_306,In_1207);
nor U837 (N_837,N_182,N_362);
and U838 (N_838,In_829,In_1026);
nor U839 (N_839,In_682,N_110);
nor U840 (N_840,In_1017,In_1103);
xnor U841 (N_841,N_625,N_313);
nand U842 (N_842,N_29,N_64);
and U843 (N_843,N_568,In_949);
and U844 (N_844,In_817,In_422);
or U845 (N_845,N_160,In_570);
nand U846 (N_846,N_430,In_1337);
nand U847 (N_847,In_871,N_197);
or U848 (N_848,N_186,In_24);
nand U849 (N_849,N_199,N_636);
nand U850 (N_850,N_252,In_1287);
and U851 (N_851,N_331,In_699);
nor U852 (N_852,N_661,In_187);
xnor U853 (N_853,N_670,In_250);
or U854 (N_854,In_1297,N_604);
or U855 (N_855,N_627,In_1262);
or U856 (N_856,In_419,In_1293);
and U857 (N_857,In_305,N_39);
and U858 (N_858,N_563,In_1292);
xor U859 (N_859,N_749,N_42);
or U860 (N_860,In_105,N_742);
nand U861 (N_861,In_1449,N_150);
nand U862 (N_862,In_472,N_743);
or U863 (N_863,N_703,In_227);
xor U864 (N_864,In_914,N_697);
xor U865 (N_865,In_477,In_493);
xor U866 (N_866,In_375,N_472);
nor U867 (N_867,N_277,N_735);
and U868 (N_868,In_175,N_645);
nor U869 (N_869,In_640,In_499);
or U870 (N_870,N_244,In_244);
nor U871 (N_871,In_1030,In_1465);
and U872 (N_872,N_269,N_278);
xnor U873 (N_873,N_152,In_1439);
nor U874 (N_874,N_207,N_473);
xor U875 (N_875,In_605,N_687);
xor U876 (N_876,N_750,In_67);
xor U877 (N_877,N_342,N_699);
and U878 (N_878,N_85,In_185);
nand U879 (N_879,N_772,In_1257);
and U880 (N_880,N_777,In_40);
and U881 (N_881,N_695,N_353);
and U882 (N_882,N_846,N_775);
and U883 (N_883,In_841,N_768);
or U884 (N_884,N_873,N_685);
xnor U885 (N_885,N_752,N_173);
xor U886 (N_886,In_673,N_648);
nor U887 (N_887,N_385,In_1316);
or U888 (N_888,N_412,In_344);
xor U889 (N_889,N_453,In_277);
xor U890 (N_890,N_463,N_767);
xnor U891 (N_891,N_654,N_792);
xor U892 (N_892,In_718,N_428);
and U893 (N_893,N_806,N_662);
nor U894 (N_894,N_328,N_830);
xor U895 (N_895,In_560,In_799);
or U896 (N_896,In_708,In_469);
and U897 (N_897,N_632,N_555);
nor U898 (N_898,N_575,N_821);
or U899 (N_899,N_684,N_302);
nor U900 (N_900,N_849,N_798);
xor U901 (N_901,In_995,N_26);
or U902 (N_902,N_225,N_567);
or U903 (N_903,In_1360,N_711);
and U904 (N_904,N_509,N_864);
xor U905 (N_905,In_237,N_531);
or U906 (N_906,N_321,N_758);
nor U907 (N_907,N_803,In_1428);
or U908 (N_908,N_238,N_810);
nor U909 (N_909,In_1475,N_582);
or U910 (N_910,N_510,In_123);
or U911 (N_911,N_852,N_341);
nand U912 (N_912,In_4,N_870);
nor U913 (N_913,N_833,N_598);
or U914 (N_914,In_246,N_819);
and U915 (N_915,N_841,N_794);
or U916 (N_916,In_514,N_556);
and U917 (N_917,In_1226,In_706);
and U918 (N_918,N_853,N_226);
nor U919 (N_919,In_1349,In_461);
nor U920 (N_920,In_224,In_1005);
and U921 (N_921,In_484,N_393);
nand U922 (N_922,In_1027,In_922);
xnor U923 (N_923,N_436,N_793);
nor U924 (N_924,In_32,In_1081);
nand U925 (N_925,N_488,In_776);
nor U926 (N_926,N_668,N_551);
xor U927 (N_927,N_518,N_611);
xor U928 (N_928,In_252,N_603);
or U929 (N_929,N_657,N_708);
nand U930 (N_930,N_352,N_716);
or U931 (N_931,N_200,N_489);
and U932 (N_932,In_1178,N_612);
nor U933 (N_933,In_827,N_188);
and U934 (N_934,N_52,N_557);
nor U935 (N_935,In_314,In_652);
nor U936 (N_936,In_674,N_651);
nor U937 (N_937,N_622,N_635);
nor U938 (N_938,In_1247,N_831);
xnor U939 (N_939,N_602,N_628);
nor U940 (N_940,N_408,In_139);
nand U941 (N_941,N_272,N_780);
nor U942 (N_942,N_127,In_713);
xor U943 (N_943,In_1334,In_919);
xnor U944 (N_944,In_1289,N_454);
nor U945 (N_945,N_268,N_675);
or U946 (N_946,N_815,In_577);
nor U947 (N_947,In_1277,N_760);
and U948 (N_948,In_903,In_85);
nand U949 (N_949,N_843,N_376);
nor U950 (N_950,N_649,In_37);
xnor U951 (N_951,In_1260,In_770);
nand U952 (N_952,N_848,N_354);
or U953 (N_953,In_202,N_84);
nand U954 (N_954,N_583,N_655);
nand U955 (N_955,N_720,N_790);
and U956 (N_956,N_856,In_913);
xor U957 (N_957,N_859,N_874);
nand U958 (N_958,N_730,In_59);
nand U959 (N_959,N_104,N_610);
nor U960 (N_960,N_725,In_739);
xor U961 (N_961,N_679,N_638);
or U962 (N_962,In_1278,In_1155);
and U963 (N_963,In_755,N_820);
nand U964 (N_964,N_753,N_825);
xor U965 (N_965,In_14,In_1264);
or U966 (N_966,N_338,N_761);
and U967 (N_967,N_81,In_1139);
nand U968 (N_968,In_118,In_1058);
xnor U969 (N_969,In_439,N_71);
nand U970 (N_970,In_388,In_511);
nand U971 (N_971,N_667,N_211);
xor U972 (N_972,N_414,In_275);
nor U973 (N_973,In_467,N_765);
nor U974 (N_974,N_339,In_1172);
xnor U975 (N_975,N_724,N_809);
nor U976 (N_976,N_146,N_709);
and U977 (N_977,N_666,N_267);
xnor U978 (N_978,N_620,N_245);
and U979 (N_979,In_748,N_129);
nor U980 (N_980,N_171,N_663);
xor U981 (N_981,N_511,N_469);
xnor U982 (N_982,N_131,N_500);
and U983 (N_983,In_245,N_525);
nand U984 (N_984,N_601,In_1315);
or U985 (N_985,N_745,In_886);
nand U986 (N_986,In_483,N_795);
or U987 (N_987,In_320,In_1042);
xor U988 (N_988,N_586,N_544);
xnor U989 (N_989,In_932,N_596);
nand U990 (N_990,N_597,N_283);
nor U991 (N_991,In_73,N_394);
nor U992 (N_992,In_1123,N_584);
nand U993 (N_993,N_738,N_585);
nor U994 (N_994,In_902,N_438);
and U995 (N_995,N_465,N_858);
xor U996 (N_996,N_276,N_295);
or U997 (N_997,N_498,N_98);
or U998 (N_998,N_634,In_386);
nand U999 (N_999,N_501,N_726);
and U1000 (N_1000,N_886,In_1303);
nor U1001 (N_1001,In_861,N_902);
nand U1002 (N_1002,N_947,N_572);
nor U1003 (N_1003,N_429,In_371);
or U1004 (N_1004,N_882,N_754);
and U1005 (N_1005,In_1196,N_885);
nand U1006 (N_1006,In_631,N_909);
and U1007 (N_1007,N_5,N_876);
nor U1008 (N_1008,In_940,N_881);
and U1009 (N_1009,N_688,N_952);
xnor U1010 (N_1010,N_439,In_851);
nor U1011 (N_1011,In_1423,In_507);
nor U1012 (N_1012,N_1,N_926);
nand U1013 (N_1013,In_633,In_1168);
xor U1014 (N_1014,N_298,N_578);
nand U1015 (N_1015,N_958,N_10);
xnor U1016 (N_1016,In_751,N_718);
nor U1017 (N_1017,In_835,N_862);
and U1018 (N_1018,N_811,In_1208);
or U1019 (N_1019,N_691,N_836);
xnor U1020 (N_1020,In_342,N_914);
and U1021 (N_1021,N_996,N_523);
and U1022 (N_1022,In_1240,In_846);
nor U1023 (N_1023,N_519,N_529);
nand U1024 (N_1024,N_714,N_936);
nor U1025 (N_1025,N_800,N_804);
and U1026 (N_1026,In_468,N_847);
xnor U1027 (N_1027,N_978,In_501);
xnor U1028 (N_1028,N_710,N_875);
nand U1029 (N_1029,N_293,In_702);
nor U1030 (N_1030,In_159,In_1286);
nor U1031 (N_1031,In_377,N_609);
or U1032 (N_1032,N_894,N_925);
nand U1033 (N_1033,N_305,In_733);
and U1034 (N_1034,In_404,N_906);
nand U1035 (N_1035,N_995,N_991);
nor U1036 (N_1036,N_371,N_860);
nand U1037 (N_1037,N_678,N_450);
or U1038 (N_1038,N_824,N_646);
or U1039 (N_1039,N_877,N_664);
or U1040 (N_1040,In_703,In_607);
and U1041 (N_1041,N_209,N_883);
or U1042 (N_1042,N_637,N_837);
xnor U1043 (N_1043,N_762,N_559);
or U1044 (N_1044,In_993,N_773);
and U1045 (N_1045,In_212,N_826);
nand U1046 (N_1046,N_916,N_801);
or U1047 (N_1047,N_972,N_680);
nand U1048 (N_1048,N_562,N_968);
or U1049 (N_1049,In_1371,N_690);
and U1050 (N_1050,In_975,N_442);
or U1051 (N_1051,In_614,N_168);
xor U1052 (N_1052,N_871,N_387);
xnor U1053 (N_1053,N_791,N_672);
or U1054 (N_1054,N_401,In_69);
nor U1055 (N_1055,N_932,In_519);
or U1056 (N_1056,In_264,N_764);
or U1057 (N_1057,N_822,In_362);
or U1058 (N_1058,In_197,N_963);
nand U1059 (N_1059,N_631,N_222);
and U1060 (N_1060,In_213,N_969);
xor U1061 (N_1061,N_570,N_924);
xor U1062 (N_1062,N_789,N_766);
or U1063 (N_1063,N_907,N_986);
xor U1064 (N_1064,N_918,In_611);
xor U1065 (N_1065,N_17,N_807);
nand U1066 (N_1066,N_960,In_516);
and U1067 (N_1067,N_917,N_900);
and U1068 (N_1068,N_839,N_832);
nor U1069 (N_1069,In_394,N_850);
and U1070 (N_1070,In_503,N_954);
nor U1071 (N_1071,N_481,In_35);
and U1072 (N_1072,N_344,N_660);
nor U1073 (N_1073,N_816,N_381);
nand U1074 (N_1074,In_1220,N_513);
nor U1075 (N_1075,N_845,In_384);
xor U1076 (N_1076,N_674,N_256);
xor U1077 (N_1077,N_644,N_965);
xor U1078 (N_1078,In_552,In_1121);
or U1079 (N_1079,In_284,N_774);
xnor U1080 (N_1080,N_989,N_979);
nor U1081 (N_1081,In_20,In_906);
xor U1082 (N_1082,In_816,N_86);
or U1083 (N_1083,N_624,N_903);
xor U1084 (N_1084,In_1197,N_592);
or U1085 (N_1085,In_1243,N_731);
nand U1086 (N_1086,N_747,In_609);
nand U1087 (N_1087,N_310,N_491);
nand U1088 (N_1088,In_521,N_992);
or U1089 (N_1089,In_387,In_530);
nor U1090 (N_1090,N_834,In_1266);
or U1091 (N_1091,In_169,N_348);
or U1092 (N_1092,N_956,N_993);
xor U1093 (N_1093,N_808,In_809);
nand U1094 (N_1094,N_445,In_307);
nor U1095 (N_1095,N_922,N_889);
xor U1096 (N_1096,In_350,In_1213);
xor U1097 (N_1097,N_966,N_984);
xnor U1098 (N_1098,N_911,N_842);
xnor U1099 (N_1099,N_890,In_623);
nor U1100 (N_1100,N_574,N_769);
nand U1101 (N_1101,N_538,N_505);
nor U1102 (N_1102,N_957,In_432);
xor U1103 (N_1103,N_945,N_553);
nand U1104 (N_1104,In_1147,N_411);
xor U1105 (N_1105,In_427,N_704);
and U1106 (N_1106,N_447,N_43);
nor U1107 (N_1107,In_313,N_971);
and U1108 (N_1108,N_639,In_492);
or U1109 (N_1109,N_744,N_942);
xor U1110 (N_1110,N_304,In_1366);
nor U1111 (N_1111,N_284,In_1356);
xnor U1112 (N_1112,In_29,N_613);
and U1113 (N_1113,N_908,N_231);
nand U1114 (N_1114,N_827,In_1341);
and U1115 (N_1115,In_1401,N_326);
nand U1116 (N_1116,N_878,N_887);
or U1117 (N_1117,N_999,N_149);
or U1118 (N_1118,N_68,N_420);
and U1119 (N_1119,N_28,N_650);
or U1120 (N_1120,N_532,N_796);
nor U1121 (N_1121,In_877,In_1056);
nor U1122 (N_1122,In_1021,In_1351);
nor U1123 (N_1123,N_390,N_534);
and U1124 (N_1124,N_135,N_788);
or U1125 (N_1125,N_642,N_915);
and U1126 (N_1126,N_1069,N_177);
xnor U1127 (N_1127,N_1012,In_1067);
nand U1128 (N_1128,N_647,N_683);
or U1129 (N_1129,N_1097,N_1035);
xnor U1130 (N_1130,N_307,N_953);
xnor U1131 (N_1131,N_927,In_945);
nor U1132 (N_1132,N_817,N_1122);
nand U1133 (N_1133,N_1054,N_1007);
or U1134 (N_1134,In_1470,N_943);
or U1135 (N_1135,In_348,N_897);
nand U1136 (N_1136,N_865,In_1122);
or U1137 (N_1137,N_1063,N_109);
and U1138 (N_1138,N_1100,N_799);
nor U1139 (N_1139,N_712,N_1031);
and U1140 (N_1140,N_784,N_1003);
or U1141 (N_1141,N_929,N_785);
and U1142 (N_1142,In_504,N_961);
and U1143 (N_1143,N_388,N_732);
or U1144 (N_1144,N_462,N_1049);
and U1145 (N_1145,N_1106,N_733);
nand U1146 (N_1146,N_778,N_1088);
and U1147 (N_1147,N_955,N_1094);
nor U1148 (N_1148,N_1101,N_1013);
or U1149 (N_1149,N_851,N_1025);
nand U1150 (N_1150,N_1040,N_681);
or U1151 (N_1151,N_482,In_585);
nor U1152 (N_1152,N_1037,N_891);
and U1153 (N_1153,N_288,N_206);
nor U1154 (N_1154,N_1053,N_504);
xnor U1155 (N_1155,N_861,In_437);
nand U1156 (N_1156,N_1010,N_823);
nand U1157 (N_1157,N_652,N_770);
or U1158 (N_1158,N_879,N_216);
xor U1159 (N_1159,N_896,N_951);
nand U1160 (N_1160,N_1047,N_1041);
nand U1161 (N_1161,N_854,N_829);
nand U1162 (N_1162,N_1030,N_895);
xnor U1163 (N_1163,N_1055,N_1109);
nand U1164 (N_1164,N_1115,In_117);
xnor U1165 (N_1165,N_921,N_985);
nand U1166 (N_1166,N_253,N_227);
and U1167 (N_1167,N_1064,N_641);
xor U1168 (N_1168,N_405,N_383);
and U1169 (N_1169,N_1065,N_757);
and U1170 (N_1170,N_1038,N_756);
xor U1171 (N_1171,N_1091,N_594);
nand U1172 (N_1172,N_863,In_395);
or U1173 (N_1173,In_830,In_70);
and U1174 (N_1174,N_1029,In_1174);
and U1175 (N_1175,In_1482,N_516);
nor U1176 (N_1176,N_759,N_1114);
xnor U1177 (N_1177,N_1066,In_550);
and U1178 (N_1178,N_1021,N_904);
xnor U1179 (N_1179,N_263,N_1068);
xnor U1180 (N_1180,N_755,N_931);
and U1181 (N_1181,N_665,N_1048);
xor U1182 (N_1182,N_1015,N_997);
or U1183 (N_1183,N_814,N_571);
nor U1184 (N_1184,N_867,N_786);
and U1185 (N_1185,N_1034,In_361);
and U1186 (N_1186,N_838,N_1020);
nand U1187 (N_1187,N_1105,N_959);
or U1188 (N_1188,In_198,In_912);
nand U1189 (N_1189,N_541,N_533);
or U1190 (N_1190,N_797,In_1227);
or U1191 (N_1191,N_899,N_893);
nand U1192 (N_1192,N_1078,N_1059);
nand U1193 (N_1193,N_392,N_1044);
nor U1194 (N_1194,N_928,N_1103);
xor U1195 (N_1195,N_776,In_363);
nand U1196 (N_1196,In_500,N_1077);
nand U1197 (N_1197,N_1024,N_974);
nand U1198 (N_1198,N_884,N_857);
nand U1199 (N_1199,N_1067,N_988);
or U1200 (N_1200,N_658,N_1061);
nand U1201 (N_1201,N_934,N_1080);
nand U1202 (N_1202,N_910,N_1014);
and U1203 (N_1203,N_905,N_1058);
and U1204 (N_1204,N_540,N_1000);
xor U1205 (N_1205,N_589,N_976);
nand U1206 (N_1206,N_977,N_990);
xor U1207 (N_1207,N_512,N_449);
xor U1208 (N_1208,In_306,N_913);
nand U1209 (N_1209,In_1230,N_14);
xor U1210 (N_1210,N_872,N_1002);
nand U1211 (N_1211,N_554,N_1076);
nand U1212 (N_1212,N_901,N_741);
nand U1213 (N_1213,N_1102,N_812);
or U1214 (N_1214,N_1107,In_1095);
nor U1215 (N_1215,N_1104,N_1011);
nand U1216 (N_1216,N_1095,N_692);
or U1217 (N_1217,In_989,N_659);
and U1218 (N_1218,N_1108,N_1045);
nor U1219 (N_1219,N_987,N_919);
and U1220 (N_1220,N_739,N_783);
nor U1221 (N_1221,N_998,N_132);
xor U1222 (N_1222,N_1073,In_291);
or U1223 (N_1223,N_1046,In_571);
or U1224 (N_1224,N_802,N_590);
or U1225 (N_1225,N_923,N_869);
xor U1226 (N_1226,N_828,N_172);
or U1227 (N_1227,N_938,N_944);
and U1228 (N_1228,N_1086,N_279);
nor U1229 (N_1229,In_1455,N_1090);
and U1230 (N_1230,N_618,N_941);
and U1231 (N_1231,N_930,N_868);
or U1232 (N_1232,N_866,In_828);
nand U1233 (N_1233,In_434,In_1110);
or U1234 (N_1234,In_282,N_1005);
nor U1235 (N_1235,N_363,N_1116);
and U1236 (N_1236,N_1039,In_122);
or U1237 (N_1237,N_1042,N_1009);
and U1238 (N_1238,N_566,N_1081);
and U1239 (N_1239,N_1056,In_1491);
and U1240 (N_1240,N_736,In_1238);
nor U1241 (N_1241,N_980,N_451);
or U1242 (N_1242,N_727,In_656);
or U1243 (N_1243,N_892,N_656);
xor U1244 (N_1244,N_1119,N_325);
nor U1245 (N_1245,N_973,N_763);
xor U1246 (N_1246,N_1032,N_734);
nor U1247 (N_1247,N_1098,N_948);
xnor U1248 (N_1248,N_623,N_1093);
nand U1249 (N_1249,N_818,In_1494);
or U1250 (N_1250,N_1178,N_1170);
and U1251 (N_1251,N_813,N_949);
or U1252 (N_1252,N_962,N_1192);
or U1253 (N_1253,In_1141,N_1175);
and U1254 (N_1254,N_130,N_1140);
nand U1255 (N_1255,N_1079,N_1022);
or U1256 (N_1256,N_205,N_1135);
and U1257 (N_1257,N_1043,N_1241);
or U1258 (N_1258,N_1139,N_1247);
nor U1259 (N_1259,N_1182,N_1083);
nor U1260 (N_1260,N_1228,In_1090);
xnor U1261 (N_1261,N_1205,N_940);
nand U1262 (N_1262,N_1209,N_1222);
nand U1263 (N_1263,N_1163,N_1166);
and U1264 (N_1264,N_1188,N_1017);
and U1265 (N_1265,N_1164,N_524);
and U1266 (N_1266,N_419,N_1173);
or U1267 (N_1267,In_862,N_1249);
and U1268 (N_1268,N_1123,N_840);
nand U1269 (N_1269,N_1131,N_855);
or U1270 (N_1270,N_880,N_1156);
nor U1271 (N_1271,N_1238,N_1153);
nand U1272 (N_1272,N_737,N_25);
xnor U1273 (N_1273,N_1019,N_1197);
nor U1274 (N_1274,N_1221,N_1125);
or U1275 (N_1275,In_1184,N_1240);
nand U1276 (N_1276,N_1171,N_1190);
xor U1277 (N_1277,N_398,N_677);
nand U1278 (N_1278,N_1074,N_1199);
nand U1279 (N_1279,In_763,N_1208);
xnor U1280 (N_1280,In_441,N_1231);
nor U1281 (N_1281,N_1145,N_1147);
or U1282 (N_1282,N_1210,N_1143);
and U1283 (N_1283,N_1087,N_1172);
nand U1284 (N_1284,N_1084,N_835);
nor U1285 (N_1285,N_994,N_898);
or U1286 (N_1286,N_751,N_983);
and U1287 (N_1287,N_1219,N_1174);
xnor U1288 (N_1288,N_1155,N_912);
or U1289 (N_1289,N_1198,N_140);
and U1290 (N_1290,N_920,N_1186);
and U1291 (N_1291,In_285,N_1132);
and U1292 (N_1292,N_982,N_1243);
and U1293 (N_1293,N_1023,N_975);
xnor U1294 (N_1294,N_1230,N_1144);
or U1295 (N_1295,N_1033,In_1344);
xnor U1296 (N_1296,N_1202,N_1124);
or U1297 (N_1297,N_1126,N_1235);
nand U1298 (N_1298,In_215,In_119);
xnor U1299 (N_1299,N_1207,N_946);
and U1300 (N_1300,N_539,N_1184);
nand U1301 (N_1301,In_26,N_1130);
nand U1302 (N_1302,N_844,N_1027);
or U1303 (N_1303,N_382,N_1121);
and U1304 (N_1304,N_1085,N_1008);
or U1305 (N_1305,N_1089,N_1236);
nor U1306 (N_1306,N_782,N_1134);
and U1307 (N_1307,N_1211,N_1214);
and U1308 (N_1308,N_888,N_1050);
nand U1309 (N_1309,N_1092,N_474);
nand U1310 (N_1310,In_1003,N_1072);
nand U1311 (N_1311,N_1196,N_1181);
xnor U1312 (N_1312,N_1176,N_1193);
or U1313 (N_1313,N_1191,N_1203);
nor U1314 (N_1314,N_682,N_1138);
nor U1315 (N_1315,N_1051,In_655);
nand U1316 (N_1316,N_970,N_1118);
nor U1317 (N_1317,N_1136,N_1150);
nor U1318 (N_1318,N_1148,N_1234);
xor U1319 (N_1319,N_1071,N_1133);
nand U1320 (N_1320,N_1162,N_1242);
nor U1321 (N_1321,In_1202,N_1001);
and U1322 (N_1322,N_1227,N_1112);
nor U1323 (N_1323,N_1159,N_1137);
nand U1324 (N_1324,N_1129,N_292);
nor U1325 (N_1325,In_474,N_1218);
and U1326 (N_1326,N_939,N_1111);
or U1327 (N_1327,N_1113,N_967);
xor U1328 (N_1328,N_1177,N_1004);
xnor U1329 (N_1329,N_1018,N_1195);
nand U1330 (N_1330,N_1215,N_614);
xnor U1331 (N_1331,N_1128,N_1070);
or U1332 (N_1332,N_787,N_1239);
nor U1333 (N_1333,N_1225,N_1149);
and U1334 (N_1334,N_1016,N_1180);
nor U1335 (N_1335,N_1194,N_1246);
nor U1336 (N_1336,In_1256,In_1249);
nor U1337 (N_1337,N_1142,N_1248);
xor U1338 (N_1338,N_1216,N_1244);
nor U1339 (N_1339,N_937,N_1062);
nand U1340 (N_1340,N_702,N_1226);
nand U1341 (N_1341,N_1185,N_1213);
nor U1342 (N_1342,N_1161,N_1158);
nand U1343 (N_1343,N_1165,N_1117);
nor U1344 (N_1344,N_1204,N_717);
or U1345 (N_1345,N_1187,In_826);
xor U1346 (N_1346,N_1057,N_1120);
nand U1347 (N_1347,In_681,N_1167);
nand U1348 (N_1348,N_1220,N_1036);
nor U1349 (N_1349,N_1169,In_150);
nor U1350 (N_1350,N_1157,N_1154);
nor U1351 (N_1351,N_1224,N_1075);
xor U1352 (N_1352,N_1160,N_1060);
and U1353 (N_1353,N_1179,N_1006);
nor U1354 (N_1354,N_1189,N_805);
and U1355 (N_1355,In_471,N_964);
nand U1356 (N_1356,N_1245,N_1099);
and U1357 (N_1357,N_1183,N_1229);
and U1358 (N_1358,N_1141,N_1201);
nand U1359 (N_1359,N_781,N_1237);
or U1360 (N_1360,N_1152,N_981);
xor U1361 (N_1361,N_1232,N_771);
or U1362 (N_1362,N_1206,N_1127);
and U1363 (N_1363,N_950,N_1212);
nand U1364 (N_1364,N_935,N_1052);
or U1365 (N_1365,N_605,N_7);
nor U1366 (N_1366,N_1217,N_76);
or U1367 (N_1367,N_1026,N_779);
nor U1368 (N_1368,N_1082,N_1146);
nor U1369 (N_1369,N_1028,N_396);
and U1370 (N_1370,N_1223,In_470);
nand U1371 (N_1371,N_1233,N_1200);
xor U1372 (N_1372,N_1168,N_1096);
nand U1373 (N_1373,N_1151,N_933);
or U1374 (N_1374,N_273,N_1110);
and U1375 (N_1375,N_1374,N_1294);
and U1376 (N_1376,N_1331,N_1313);
or U1377 (N_1377,N_1356,N_1314);
and U1378 (N_1378,N_1269,N_1365);
and U1379 (N_1379,N_1338,N_1251);
nor U1380 (N_1380,N_1296,N_1254);
xor U1381 (N_1381,N_1271,N_1362);
and U1382 (N_1382,N_1350,N_1343);
and U1383 (N_1383,N_1351,N_1308);
xnor U1384 (N_1384,N_1298,N_1359);
nor U1385 (N_1385,N_1299,N_1293);
and U1386 (N_1386,N_1274,N_1316);
nand U1387 (N_1387,N_1253,N_1360);
or U1388 (N_1388,N_1341,N_1267);
xor U1389 (N_1389,N_1326,N_1322);
nor U1390 (N_1390,N_1279,N_1371);
nor U1391 (N_1391,N_1345,N_1291);
nand U1392 (N_1392,N_1364,N_1281);
nor U1393 (N_1393,N_1252,N_1270);
xnor U1394 (N_1394,N_1318,N_1300);
xor U1395 (N_1395,N_1315,N_1335);
xnor U1396 (N_1396,N_1290,N_1334);
and U1397 (N_1397,N_1268,N_1255);
xor U1398 (N_1398,N_1366,N_1333);
nand U1399 (N_1399,N_1276,N_1280);
nand U1400 (N_1400,N_1321,N_1260);
or U1401 (N_1401,N_1325,N_1257);
xor U1402 (N_1402,N_1324,N_1263);
nor U1403 (N_1403,N_1285,N_1262);
xor U1404 (N_1404,N_1288,N_1311);
nor U1405 (N_1405,N_1354,N_1355);
nor U1406 (N_1406,N_1278,N_1340);
nor U1407 (N_1407,N_1317,N_1258);
or U1408 (N_1408,N_1358,N_1328);
and U1409 (N_1409,N_1273,N_1286);
nand U1410 (N_1410,N_1347,N_1370);
or U1411 (N_1411,N_1352,N_1272);
nor U1412 (N_1412,N_1301,N_1259);
nand U1413 (N_1413,N_1332,N_1289);
or U1414 (N_1414,N_1310,N_1336);
nand U1415 (N_1415,N_1361,N_1330);
or U1416 (N_1416,N_1329,N_1250);
nand U1417 (N_1417,N_1277,N_1348);
or U1418 (N_1418,N_1323,N_1287);
and U1419 (N_1419,N_1320,N_1302);
and U1420 (N_1420,N_1297,N_1363);
nand U1421 (N_1421,N_1368,N_1295);
xor U1422 (N_1422,N_1312,N_1357);
or U1423 (N_1423,N_1303,N_1282);
or U1424 (N_1424,N_1265,N_1327);
and U1425 (N_1425,N_1337,N_1266);
nand U1426 (N_1426,N_1372,N_1342);
nor U1427 (N_1427,N_1284,N_1346);
and U1428 (N_1428,N_1369,N_1373);
or U1429 (N_1429,N_1349,N_1339);
or U1430 (N_1430,N_1306,N_1261);
nor U1431 (N_1431,N_1344,N_1256);
nand U1432 (N_1432,N_1353,N_1319);
nand U1433 (N_1433,N_1307,N_1292);
xnor U1434 (N_1434,N_1305,N_1264);
nor U1435 (N_1435,N_1367,N_1283);
and U1436 (N_1436,N_1275,N_1309);
or U1437 (N_1437,N_1304,N_1319);
xnor U1438 (N_1438,N_1254,N_1304);
or U1439 (N_1439,N_1337,N_1348);
and U1440 (N_1440,N_1311,N_1294);
nand U1441 (N_1441,N_1255,N_1359);
nor U1442 (N_1442,N_1356,N_1362);
and U1443 (N_1443,N_1371,N_1298);
nor U1444 (N_1444,N_1264,N_1323);
or U1445 (N_1445,N_1339,N_1289);
nand U1446 (N_1446,N_1307,N_1261);
and U1447 (N_1447,N_1282,N_1275);
nor U1448 (N_1448,N_1347,N_1365);
xor U1449 (N_1449,N_1350,N_1273);
or U1450 (N_1450,N_1347,N_1288);
nand U1451 (N_1451,N_1298,N_1265);
or U1452 (N_1452,N_1347,N_1297);
nor U1453 (N_1453,N_1316,N_1317);
xnor U1454 (N_1454,N_1340,N_1366);
nand U1455 (N_1455,N_1371,N_1257);
nor U1456 (N_1456,N_1297,N_1278);
or U1457 (N_1457,N_1258,N_1266);
or U1458 (N_1458,N_1367,N_1341);
or U1459 (N_1459,N_1372,N_1355);
nor U1460 (N_1460,N_1260,N_1363);
nand U1461 (N_1461,N_1334,N_1339);
xnor U1462 (N_1462,N_1374,N_1330);
xor U1463 (N_1463,N_1274,N_1334);
or U1464 (N_1464,N_1294,N_1366);
and U1465 (N_1465,N_1297,N_1365);
nor U1466 (N_1466,N_1303,N_1369);
xnor U1467 (N_1467,N_1371,N_1313);
xnor U1468 (N_1468,N_1347,N_1337);
nor U1469 (N_1469,N_1327,N_1362);
or U1470 (N_1470,N_1258,N_1373);
nand U1471 (N_1471,N_1348,N_1289);
xor U1472 (N_1472,N_1317,N_1274);
xor U1473 (N_1473,N_1355,N_1305);
and U1474 (N_1474,N_1297,N_1292);
nand U1475 (N_1475,N_1358,N_1320);
and U1476 (N_1476,N_1278,N_1255);
or U1477 (N_1477,N_1370,N_1327);
or U1478 (N_1478,N_1259,N_1362);
nand U1479 (N_1479,N_1344,N_1334);
and U1480 (N_1480,N_1301,N_1342);
nand U1481 (N_1481,N_1342,N_1282);
and U1482 (N_1482,N_1252,N_1275);
xnor U1483 (N_1483,N_1323,N_1329);
nor U1484 (N_1484,N_1345,N_1262);
nor U1485 (N_1485,N_1330,N_1369);
and U1486 (N_1486,N_1344,N_1297);
xnor U1487 (N_1487,N_1291,N_1312);
or U1488 (N_1488,N_1312,N_1372);
or U1489 (N_1489,N_1293,N_1271);
xor U1490 (N_1490,N_1311,N_1352);
nand U1491 (N_1491,N_1320,N_1336);
xor U1492 (N_1492,N_1295,N_1252);
xnor U1493 (N_1493,N_1304,N_1311);
or U1494 (N_1494,N_1315,N_1297);
xor U1495 (N_1495,N_1293,N_1259);
nor U1496 (N_1496,N_1334,N_1335);
or U1497 (N_1497,N_1286,N_1271);
or U1498 (N_1498,N_1346,N_1296);
or U1499 (N_1499,N_1345,N_1280);
nand U1500 (N_1500,N_1395,N_1460);
or U1501 (N_1501,N_1450,N_1483);
and U1502 (N_1502,N_1498,N_1487);
xnor U1503 (N_1503,N_1390,N_1377);
or U1504 (N_1504,N_1429,N_1466);
and U1505 (N_1505,N_1431,N_1397);
or U1506 (N_1506,N_1447,N_1472);
xor U1507 (N_1507,N_1438,N_1391);
or U1508 (N_1508,N_1485,N_1441);
or U1509 (N_1509,N_1482,N_1401);
and U1510 (N_1510,N_1481,N_1459);
nor U1511 (N_1511,N_1495,N_1494);
xnor U1512 (N_1512,N_1497,N_1430);
xor U1513 (N_1513,N_1455,N_1415);
nand U1514 (N_1514,N_1427,N_1477);
nor U1515 (N_1515,N_1404,N_1436);
and U1516 (N_1516,N_1467,N_1428);
xnor U1517 (N_1517,N_1402,N_1463);
nand U1518 (N_1518,N_1442,N_1439);
and U1519 (N_1519,N_1408,N_1392);
xnor U1520 (N_1520,N_1376,N_1381);
or U1521 (N_1521,N_1416,N_1452);
nand U1522 (N_1522,N_1384,N_1480);
xor U1523 (N_1523,N_1453,N_1473);
and U1524 (N_1524,N_1488,N_1446);
or U1525 (N_1525,N_1440,N_1464);
and U1526 (N_1526,N_1417,N_1414);
nor U1527 (N_1527,N_1435,N_1424);
nor U1528 (N_1528,N_1432,N_1437);
nor U1529 (N_1529,N_1421,N_1405);
or U1530 (N_1530,N_1385,N_1496);
nand U1531 (N_1531,N_1470,N_1478);
nand U1532 (N_1532,N_1382,N_1490);
nand U1533 (N_1533,N_1389,N_1379);
or U1534 (N_1534,N_1469,N_1388);
nand U1535 (N_1535,N_1476,N_1474);
xor U1536 (N_1536,N_1465,N_1410);
and U1537 (N_1537,N_1449,N_1422);
nand U1538 (N_1538,N_1425,N_1468);
nand U1539 (N_1539,N_1454,N_1444);
nor U1540 (N_1540,N_1394,N_1406);
and U1541 (N_1541,N_1456,N_1409);
nor U1542 (N_1542,N_1443,N_1493);
nand U1543 (N_1543,N_1413,N_1378);
xnor U1544 (N_1544,N_1471,N_1492);
and U1545 (N_1545,N_1499,N_1491);
or U1546 (N_1546,N_1458,N_1380);
and U1547 (N_1547,N_1399,N_1387);
xor U1548 (N_1548,N_1393,N_1407);
and U1549 (N_1549,N_1375,N_1411);
nor U1550 (N_1550,N_1457,N_1461);
or U1551 (N_1551,N_1412,N_1484);
and U1552 (N_1552,N_1403,N_1419);
and U1553 (N_1553,N_1448,N_1396);
nor U1554 (N_1554,N_1489,N_1479);
nor U1555 (N_1555,N_1486,N_1433);
xor U1556 (N_1556,N_1434,N_1386);
and U1557 (N_1557,N_1420,N_1418);
nor U1558 (N_1558,N_1383,N_1423);
nand U1559 (N_1559,N_1445,N_1400);
xnor U1560 (N_1560,N_1462,N_1426);
nor U1561 (N_1561,N_1398,N_1475);
or U1562 (N_1562,N_1451,N_1425);
xor U1563 (N_1563,N_1383,N_1412);
xnor U1564 (N_1564,N_1483,N_1381);
nand U1565 (N_1565,N_1497,N_1414);
or U1566 (N_1566,N_1447,N_1484);
and U1567 (N_1567,N_1455,N_1432);
nor U1568 (N_1568,N_1472,N_1470);
xor U1569 (N_1569,N_1457,N_1416);
nand U1570 (N_1570,N_1387,N_1428);
or U1571 (N_1571,N_1469,N_1405);
xnor U1572 (N_1572,N_1404,N_1470);
or U1573 (N_1573,N_1396,N_1423);
and U1574 (N_1574,N_1382,N_1411);
and U1575 (N_1575,N_1473,N_1464);
and U1576 (N_1576,N_1491,N_1392);
xor U1577 (N_1577,N_1463,N_1380);
nor U1578 (N_1578,N_1429,N_1413);
xnor U1579 (N_1579,N_1465,N_1379);
nor U1580 (N_1580,N_1406,N_1471);
nand U1581 (N_1581,N_1488,N_1415);
nor U1582 (N_1582,N_1484,N_1487);
nand U1583 (N_1583,N_1469,N_1382);
xnor U1584 (N_1584,N_1385,N_1436);
and U1585 (N_1585,N_1392,N_1455);
and U1586 (N_1586,N_1496,N_1378);
nand U1587 (N_1587,N_1450,N_1404);
and U1588 (N_1588,N_1495,N_1464);
or U1589 (N_1589,N_1375,N_1482);
and U1590 (N_1590,N_1401,N_1464);
nor U1591 (N_1591,N_1467,N_1389);
xnor U1592 (N_1592,N_1399,N_1398);
nor U1593 (N_1593,N_1463,N_1429);
nand U1594 (N_1594,N_1497,N_1437);
xor U1595 (N_1595,N_1448,N_1425);
xnor U1596 (N_1596,N_1384,N_1424);
and U1597 (N_1597,N_1376,N_1488);
or U1598 (N_1598,N_1430,N_1457);
xor U1599 (N_1599,N_1408,N_1427);
xnor U1600 (N_1600,N_1478,N_1402);
nand U1601 (N_1601,N_1410,N_1453);
nor U1602 (N_1602,N_1389,N_1421);
and U1603 (N_1603,N_1422,N_1431);
xnor U1604 (N_1604,N_1463,N_1394);
xnor U1605 (N_1605,N_1468,N_1466);
and U1606 (N_1606,N_1451,N_1464);
nand U1607 (N_1607,N_1429,N_1412);
or U1608 (N_1608,N_1406,N_1479);
nor U1609 (N_1609,N_1439,N_1450);
and U1610 (N_1610,N_1385,N_1499);
and U1611 (N_1611,N_1494,N_1392);
xor U1612 (N_1612,N_1476,N_1424);
and U1613 (N_1613,N_1398,N_1424);
or U1614 (N_1614,N_1485,N_1398);
nor U1615 (N_1615,N_1418,N_1454);
or U1616 (N_1616,N_1493,N_1385);
nand U1617 (N_1617,N_1399,N_1422);
xnor U1618 (N_1618,N_1496,N_1493);
or U1619 (N_1619,N_1472,N_1384);
xor U1620 (N_1620,N_1408,N_1476);
or U1621 (N_1621,N_1473,N_1427);
nand U1622 (N_1622,N_1488,N_1487);
nor U1623 (N_1623,N_1442,N_1460);
xor U1624 (N_1624,N_1397,N_1473);
and U1625 (N_1625,N_1539,N_1601);
xnor U1626 (N_1626,N_1573,N_1595);
or U1627 (N_1627,N_1616,N_1510);
nand U1628 (N_1628,N_1588,N_1600);
or U1629 (N_1629,N_1624,N_1511);
nand U1630 (N_1630,N_1548,N_1506);
or U1631 (N_1631,N_1592,N_1551);
nor U1632 (N_1632,N_1515,N_1607);
nor U1633 (N_1633,N_1504,N_1554);
or U1634 (N_1634,N_1505,N_1596);
nand U1635 (N_1635,N_1550,N_1581);
or U1636 (N_1636,N_1599,N_1576);
or U1637 (N_1637,N_1609,N_1622);
xor U1638 (N_1638,N_1611,N_1545);
and U1639 (N_1639,N_1522,N_1559);
xor U1640 (N_1640,N_1568,N_1560);
and U1641 (N_1641,N_1602,N_1534);
and U1642 (N_1642,N_1575,N_1517);
and U1643 (N_1643,N_1586,N_1583);
nand U1644 (N_1644,N_1619,N_1514);
nand U1645 (N_1645,N_1540,N_1608);
nand U1646 (N_1646,N_1562,N_1530);
xor U1647 (N_1647,N_1566,N_1582);
and U1648 (N_1648,N_1523,N_1614);
or U1649 (N_1649,N_1598,N_1574);
and U1650 (N_1650,N_1590,N_1543);
or U1651 (N_1651,N_1584,N_1524);
and U1652 (N_1652,N_1557,N_1503);
or U1653 (N_1653,N_1558,N_1561);
and U1654 (N_1654,N_1501,N_1580);
nor U1655 (N_1655,N_1535,N_1553);
xnor U1656 (N_1656,N_1552,N_1519);
nor U1657 (N_1657,N_1536,N_1587);
or U1658 (N_1658,N_1508,N_1623);
and U1659 (N_1659,N_1620,N_1546);
or U1660 (N_1660,N_1529,N_1531);
or U1661 (N_1661,N_1578,N_1516);
xor U1662 (N_1662,N_1512,N_1605);
and U1663 (N_1663,N_1606,N_1610);
or U1664 (N_1664,N_1621,N_1533);
and U1665 (N_1665,N_1542,N_1537);
and U1666 (N_1666,N_1572,N_1538);
nand U1667 (N_1667,N_1544,N_1577);
or U1668 (N_1668,N_1597,N_1526);
nand U1669 (N_1669,N_1518,N_1604);
xor U1670 (N_1670,N_1520,N_1527);
nor U1671 (N_1671,N_1500,N_1556);
nor U1672 (N_1672,N_1612,N_1549);
nand U1673 (N_1673,N_1532,N_1509);
xnor U1674 (N_1674,N_1603,N_1507);
nand U1675 (N_1675,N_1569,N_1528);
xnor U1676 (N_1676,N_1593,N_1525);
and U1677 (N_1677,N_1617,N_1567);
xor U1678 (N_1678,N_1571,N_1565);
xnor U1679 (N_1679,N_1594,N_1547);
or U1680 (N_1680,N_1591,N_1555);
xnor U1681 (N_1681,N_1541,N_1513);
xnor U1682 (N_1682,N_1521,N_1613);
or U1683 (N_1683,N_1585,N_1502);
or U1684 (N_1684,N_1563,N_1570);
and U1685 (N_1685,N_1615,N_1579);
nand U1686 (N_1686,N_1618,N_1589);
and U1687 (N_1687,N_1564,N_1612);
and U1688 (N_1688,N_1513,N_1595);
nor U1689 (N_1689,N_1528,N_1501);
xor U1690 (N_1690,N_1529,N_1607);
nor U1691 (N_1691,N_1591,N_1618);
nand U1692 (N_1692,N_1538,N_1567);
or U1693 (N_1693,N_1545,N_1544);
and U1694 (N_1694,N_1558,N_1607);
nand U1695 (N_1695,N_1622,N_1517);
nand U1696 (N_1696,N_1575,N_1556);
nand U1697 (N_1697,N_1580,N_1567);
and U1698 (N_1698,N_1547,N_1560);
xnor U1699 (N_1699,N_1572,N_1567);
and U1700 (N_1700,N_1623,N_1566);
xor U1701 (N_1701,N_1624,N_1623);
nor U1702 (N_1702,N_1552,N_1597);
and U1703 (N_1703,N_1600,N_1573);
nand U1704 (N_1704,N_1532,N_1507);
nand U1705 (N_1705,N_1616,N_1555);
nand U1706 (N_1706,N_1582,N_1595);
and U1707 (N_1707,N_1534,N_1614);
xnor U1708 (N_1708,N_1507,N_1619);
and U1709 (N_1709,N_1608,N_1568);
and U1710 (N_1710,N_1510,N_1507);
and U1711 (N_1711,N_1584,N_1578);
and U1712 (N_1712,N_1555,N_1515);
and U1713 (N_1713,N_1617,N_1519);
nor U1714 (N_1714,N_1571,N_1584);
nor U1715 (N_1715,N_1586,N_1584);
or U1716 (N_1716,N_1524,N_1560);
and U1717 (N_1717,N_1546,N_1534);
or U1718 (N_1718,N_1573,N_1589);
nand U1719 (N_1719,N_1623,N_1583);
nor U1720 (N_1720,N_1604,N_1523);
xor U1721 (N_1721,N_1606,N_1516);
or U1722 (N_1722,N_1540,N_1551);
nand U1723 (N_1723,N_1615,N_1586);
and U1724 (N_1724,N_1550,N_1540);
xor U1725 (N_1725,N_1569,N_1624);
nor U1726 (N_1726,N_1581,N_1520);
and U1727 (N_1727,N_1579,N_1617);
nor U1728 (N_1728,N_1512,N_1501);
and U1729 (N_1729,N_1617,N_1561);
nor U1730 (N_1730,N_1530,N_1580);
and U1731 (N_1731,N_1596,N_1584);
or U1732 (N_1732,N_1563,N_1504);
xor U1733 (N_1733,N_1617,N_1594);
nor U1734 (N_1734,N_1516,N_1595);
nor U1735 (N_1735,N_1538,N_1581);
and U1736 (N_1736,N_1560,N_1569);
xor U1737 (N_1737,N_1522,N_1536);
nand U1738 (N_1738,N_1518,N_1564);
nor U1739 (N_1739,N_1576,N_1507);
or U1740 (N_1740,N_1507,N_1503);
xor U1741 (N_1741,N_1537,N_1610);
or U1742 (N_1742,N_1525,N_1528);
and U1743 (N_1743,N_1529,N_1527);
nor U1744 (N_1744,N_1553,N_1589);
or U1745 (N_1745,N_1613,N_1528);
and U1746 (N_1746,N_1599,N_1511);
nand U1747 (N_1747,N_1516,N_1545);
nor U1748 (N_1748,N_1591,N_1532);
nand U1749 (N_1749,N_1539,N_1618);
nor U1750 (N_1750,N_1674,N_1732);
nand U1751 (N_1751,N_1668,N_1725);
nor U1752 (N_1752,N_1741,N_1705);
and U1753 (N_1753,N_1697,N_1645);
xnor U1754 (N_1754,N_1662,N_1686);
and U1755 (N_1755,N_1634,N_1671);
xnor U1756 (N_1756,N_1726,N_1696);
nand U1757 (N_1757,N_1708,N_1707);
or U1758 (N_1758,N_1735,N_1684);
or U1759 (N_1759,N_1699,N_1712);
nand U1760 (N_1760,N_1689,N_1744);
xnor U1761 (N_1761,N_1737,N_1648);
xor U1762 (N_1762,N_1745,N_1639);
nor U1763 (N_1763,N_1703,N_1693);
and U1764 (N_1764,N_1672,N_1640);
nor U1765 (N_1765,N_1694,N_1638);
nand U1766 (N_1766,N_1675,N_1630);
or U1767 (N_1767,N_1743,N_1667);
xnor U1768 (N_1768,N_1649,N_1669);
nor U1769 (N_1769,N_1644,N_1720);
xnor U1770 (N_1770,N_1641,N_1651);
and U1771 (N_1771,N_1700,N_1633);
nand U1772 (N_1772,N_1663,N_1710);
xnor U1773 (N_1773,N_1747,N_1738);
xnor U1774 (N_1774,N_1742,N_1691);
and U1775 (N_1775,N_1647,N_1723);
nand U1776 (N_1776,N_1659,N_1701);
nor U1777 (N_1777,N_1660,N_1673);
or U1778 (N_1778,N_1724,N_1679);
or U1779 (N_1779,N_1736,N_1654);
and U1780 (N_1780,N_1714,N_1704);
nor U1781 (N_1781,N_1731,N_1653);
xor U1782 (N_1782,N_1698,N_1642);
nor U1783 (N_1783,N_1682,N_1678);
nand U1784 (N_1784,N_1690,N_1661);
and U1785 (N_1785,N_1695,N_1728);
and U1786 (N_1786,N_1727,N_1721);
nand U1787 (N_1787,N_1656,N_1713);
and U1788 (N_1788,N_1657,N_1650);
and U1789 (N_1789,N_1646,N_1665);
or U1790 (N_1790,N_1717,N_1680);
and U1791 (N_1791,N_1677,N_1637);
and U1792 (N_1792,N_1664,N_1719);
nand U1793 (N_1793,N_1636,N_1666);
xnor U1794 (N_1794,N_1715,N_1658);
xor U1795 (N_1795,N_1635,N_1652);
xor U1796 (N_1796,N_1722,N_1706);
nand U1797 (N_1797,N_1692,N_1670);
nand U1798 (N_1798,N_1716,N_1631);
nor U1799 (N_1799,N_1626,N_1629);
xnor U1800 (N_1800,N_1711,N_1709);
nor U1801 (N_1801,N_1632,N_1748);
xor U1802 (N_1802,N_1729,N_1687);
nand U1803 (N_1803,N_1749,N_1740);
or U1804 (N_1804,N_1746,N_1718);
nor U1805 (N_1805,N_1730,N_1734);
nor U1806 (N_1806,N_1655,N_1625);
nand U1807 (N_1807,N_1643,N_1688);
xnor U1808 (N_1808,N_1676,N_1628);
nand U1809 (N_1809,N_1627,N_1733);
xor U1810 (N_1810,N_1739,N_1685);
xnor U1811 (N_1811,N_1681,N_1702);
nand U1812 (N_1812,N_1683,N_1663);
and U1813 (N_1813,N_1735,N_1652);
or U1814 (N_1814,N_1654,N_1708);
and U1815 (N_1815,N_1627,N_1724);
or U1816 (N_1816,N_1707,N_1725);
xnor U1817 (N_1817,N_1647,N_1666);
or U1818 (N_1818,N_1732,N_1680);
nand U1819 (N_1819,N_1628,N_1631);
and U1820 (N_1820,N_1692,N_1627);
nand U1821 (N_1821,N_1664,N_1637);
nand U1822 (N_1822,N_1739,N_1625);
or U1823 (N_1823,N_1728,N_1732);
and U1824 (N_1824,N_1681,N_1663);
xnor U1825 (N_1825,N_1662,N_1706);
xor U1826 (N_1826,N_1749,N_1690);
nor U1827 (N_1827,N_1666,N_1659);
nand U1828 (N_1828,N_1652,N_1681);
or U1829 (N_1829,N_1698,N_1705);
nor U1830 (N_1830,N_1704,N_1686);
nand U1831 (N_1831,N_1736,N_1708);
nand U1832 (N_1832,N_1628,N_1699);
and U1833 (N_1833,N_1674,N_1659);
or U1834 (N_1834,N_1634,N_1644);
or U1835 (N_1835,N_1657,N_1634);
nand U1836 (N_1836,N_1715,N_1725);
nor U1837 (N_1837,N_1698,N_1665);
or U1838 (N_1838,N_1701,N_1738);
and U1839 (N_1839,N_1688,N_1714);
or U1840 (N_1840,N_1726,N_1674);
xor U1841 (N_1841,N_1716,N_1650);
nor U1842 (N_1842,N_1710,N_1743);
xnor U1843 (N_1843,N_1663,N_1735);
nor U1844 (N_1844,N_1677,N_1659);
nand U1845 (N_1845,N_1697,N_1659);
nor U1846 (N_1846,N_1714,N_1678);
xor U1847 (N_1847,N_1667,N_1718);
nand U1848 (N_1848,N_1655,N_1697);
nand U1849 (N_1849,N_1644,N_1652);
xor U1850 (N_1850,N_1720,N_1693);
or U1851 (N_1851,N_1657,N_1677);
and U1852 (N_1852,N_1643,N_1733);
or U1853 (N_1853,N_1739,N_1656);
nand U1854 (N_1854,N_1727,N_1674);
nor U1855 (N_1855,N_1697,N_1737);
nor U1856 (N_1856,N_1683,N_1667);
nand U1857 (N_1857,N_1629,N_1744);
or U1858 (N_1858,N_1731,N_1664);
xor U1859 (N_1859,N_1714,N_1682);
nor U1860 (N_1860,N_1685,N_1730);
or U1861 (N_1861,N_1726,N_1647);
xor U1862 (N_1862,N_1735,N_1699);
and U1863 (N_1863,N_1703,N_1653);
nand U1864 (N_1864,N_1717,N_1739);
nand U1865 (N_1865,N_1701,N_1631);
nor U1866 (N_1866,N_1747,N_1705);
nor U1867 (N_1867,N_1673,N_1690);
or U1868 (N_1868,N_1693,N_1741);
and U1869 (N_1869,N_1637,N_1634);
nor U1870 (N_1870,N_1702,N_1639);
or U1871 (N_1871,N_1747,N_1737);
or U1872 (N_1872,N_1643,N_1709);
xnor U1873 (N_1873,N_1661,N_1643);
nand U1874 (N_1874,N_1724,N_1680);
nor U1875 (N_1875,N_1863,N_1815);
nor U1876 (N_1876,N_1819,N_1867);
nor U1877 (N_1877,N_1825,N_1858);
xnor U1878 (N_1878,N_1790,N_1827);
xnor U1879 (N_1879,N_1857,N_1782);
nor U1880 (N_1880,N_1769,N_1835);
or U1881 (N_1881,N_1794,N_1795);
or U1882 (N_1882,N_1813,N_1850);
xor U1883 (N_1883,N_1823,N_1830);
nor U1884 (N_1884,N_1842,N_1818);
and U1885 (N_1885,N_1773,N_1768);
nand U1886 (N_1886,N_1821,N_1780);
xnor U1887 (N_1887,N_1873,N_1757);
nand U1888 (N_1888,N_1811,N_1854);
or U1889 (N_1889,N_1871,N_1855);
nor U1890 (N_1890,N_1844,N_1751);
or U1891 (N_1891,N_1846,N_1786);
and U1892 (N_1892,N_1781,N_1849);
or U1893 (N_1893,N_1851,N_1788);
and U1894 (N_1894,N_1829,N_1840);
nand U1895 (N_1895,N_1817,N_1859);
nand U1896 (N_1896,N_1755,N_1816);
nand U1897 (N_1897,N_1847,N_1787);
or U1898 (N_1898,N_1799,N_1804);
or U1899 (N_1899,N_1838,N_1831);
nor U1900 (N_1900,N_1868,N_1869);
nand U1901 (N_1901,N_1785,N_1792);
nor U1902 (N_1902,N_1798,N_1803);
or U1903 (N_1903,N_1865,N_1807);
xor U1904 (N_1904,N_1833,N_1828);
nor U1905 (N_1905,N_1845,N_1820);
and U1906 (N_1906,N_1856,N_1841);
nand U1907 (N_1907,N_1802,N_1784);
nor U1908 (N_1908,N_1767,N_1758);
nand U1909 (N_1909,N_1762,N_1824);
and U1910 (N_1910,N_1837,N_1753);
nor U1911 (N_1911,N_1832,N_1861);
and U1912 (N_1912,N_1772,N_1761);
xnor U1913 (N_1913,N_1853,N_1839);
and U1914 (N_1914,N_1754,N_1783);
xnor U1915 (N_1915,N_1796,N_1771);
xor U1916 (N_1916,N_1764,N_1759);
xor U1917 (N_1917,N_1812,N_1765);
nand U1918 (N_1918,N_1791,N_1822);
nor U1919 (N_1919,N_1874,N_1793);
or U1920 (N_1920,N_1805,N_1862);
nand U1921 (N_1921,N_1809,N_1843);
nand U1922 (N_1922,N_1870,N_1848);
and U1923 (N_1923,N_1760,N_1789);
xor U1924 (N_1924,N_1774,N_1806);
nor U1925 (N_1925,N_1826,N_1864);
nand U1926 (N_1926,N_1770,N_1756);
nand U1927 (N_1927,N_1836,N_1814);
and U1928 (N_1928,N_1752,N_1777);
nor U1929 (N_1929,N_1852,N_1776);
nor U1930 (N_1930,N_1766,N_1801);
xnor U1931 (N_1931,N_1834,N_1775);
and U1932 (N_1932,N_1860,N_1872);
nor U1933 (N_1933,N_1763,N_1808);
and U1934 (N_1934,N_1779,N_1866);
nand U1935 (N_1935,N_1778,N_1800);
or U1936 (N_1936,N_1810,N_1750);
or U1937 (N_1937,N_1797,N_1874);
or U1938 (N_1938,N_1818,N_1848);
or U1939 (N_1939,N_1768,N_1822);
nor U1940 (N_1940,N_1752,N_1837);
and U1941 (N_1941,N_1777,N_1849);
or U1942 (N_1942,N_1836,N_1764);
xor U1943 (N_1943,N_1799,N_1775);
and U1944 (N_1944,N_1764,N_1820);
nor U1945 (N_1945,N_1855,N_1805);
or U1946 (N_1946,N_1808,N_1804);
nor U1947 (N_1947,N_1796,N_1759);
nand U1948 (N_1948,N_1799,N_1785);
or U1949 (N_1949,N_1788,N_1803);
nor U1950 (N_1950,N_1814,N_1802);
or U1951 (N_1951,N_1790,N_1873);
and U1952 (N_1952,N_1781,N_1764);
xnor U1953 (N_1953,N_1768,N_1809);
xnor U1954 (N_1954,N_1750,N_1848);
and U1955 (N_1955,N_1822,N_1865);
nand U1956 (N_1956,N_1820,N_1763);
or U1957 (N_1957,N_1870,N_1867);
nand U1958 (N_1958,N_1760,N_1861);
nor U1959 (N_1959,N_1865,N_1754);
and U1960 (N_1960,N_1753,N_1754);
or U1961 (N_1961,N_1793,N_1779);
xor U1962 (N_1962,N_1752,N_1821);
nor U1963 (N_1963,N_1828,N_1826);
and U1964 (N_1964,N_1851,N_1761);
nor U1965 (N_1965,N_1776,N_1862);
xor U1966 (N_1966,N_1817,N_1839);
nor U1967 (N_1967,N_1781,N_1760);
nand U1968 (N_1968,N_1868,N_1762);
xnor U1969 (N_1969,N_1870,N_1864);
nor U1970 (N_1970,N_1780,N_1811);
xor U1971 (N_1971,N_1789,N_1786);
nor U1972 (N_1972,N_1766,N_1796);
nor U1973 (N_1973,N_1796,N_1861);
or U1974 (N_1974,N_1751,N_1750);
nor U1975 (N_1975,N_1867,N_1797);
and U1976 (N_1976,N_1771,N_1864);
and U1977 (N_1977,N_1856,N_1801);
nand U1978 (N_1978,N_1832,N_1766);
or U1979 (N_1979,N_1869,N_1836);
nor U1980 (N_1980,N_1829,N_1843);
nand U1981 (N_1981,N_1874,N_1757);
and U1982 (N_1982,N_1846,N_1807);
xor U1983 (N_1983,N_1817,N_1813);
nor U1984 (N_1984,N_1872,N_1841);
xnor U1985 (N_1985,N_1833,N_1862);
xor U1986 (N_1986,N_1853,N_1796);
or U1987 (N_1987,N_1822,N_1778);
or U1988 (N_1988,N_1833,N_1837);
or U1989 (N_1989,N_1797,N_1801);
or U1990 (N_1990,N_1787,N_1869);
nand U1991 (N_1991,N_1775,N_1866);
xnor U1992 (N_1992,N_1832,N_1847);
and U1993 (N_1993,N_1831,N_1853);
or U1994 (N_1994,N_1793,N_1797);
or U1995 (N_1995,N_1860,N_1858);
xor U1996 (N_1996,N_1871,N_1859);
nor U1997 (N_1997,N_1841,N_1816);
and U1998 (N_1998,N_1860,N_1760);
xor U1999 (N_1999,N_1818,N_1769);
nor U2000 (N_2000,N_1935,N_1931);
nor U2001 (N_2001,N_1995,N_1888);
or U2002 (N_2002,N_1998,N_1951);
nand U2003 (N_2003,N_1892,N_1906);
nand U2004 (N_2004,N_1945,N_1940);
nand U2005 (N_2005,N_1879,N_1944);
xor U2006 (N_2006,N_1908,N_1877);
nor U2007 (N_2007,N_1916,N_1894);
or U2008 (N_2008,N_1939,N_1974);
nor U2009 (N_2009,N_1925,N_1948);
and U2010 (N_2010,N_1878,N_1923);
xor U2011 (N_2011,N_1937,N_1913);
nand U2012 (N_2012,N_1900,N_1897);
or U2013 (N_2013,N_1926,N_1883);
nor U2014 (N_2014,N_1992,N_1968);
nor U2015 (N_2015,N_1952,N_1993);
nand U2016 (N_2016,N_1983,N_1958);
nand U2017 (N_2017,N_1895,N_1911);
or U2018 (N_2018,N_1941,N_1876);
nor U2019 (N_2019,N_1966,N_1943);
nand U2020 (N_2020,N_1936,N_1887);
and U2021 (N_2021,N_1927,N_1982);
xnor U2022 (N_2022,N_1909,N_1915);
nor U2023 (N_2023,N_1960,N_1956);
xor U2024 (N_2024,N_1976,N_1977);
or U2025 (N_2025,N_1996,N_1882);
nor U2026 (N_2026,N_1963,N_1890);
and U2027 (N_2027,N_1917,N_1919);
nand U2028 (N_2028,N_1928,N_1930);
nand U2029 (N_2029,N_1947,N_1886);
and U2030 (N_2030,N_1999,N_1924);
xor U2031 (N_2031,N_1921,N_1946);
nand U2032 (N_2032,N_1889,N_1975);
nand U2033 (N_2033,N_1972,N_1884);
xnor U2034 (N_2034,N_1875,N_1985);
xnor U2035 (N_2035,N_1962,N_1969);
or U2036 (N_2036,N_1904,N_1910);
nand U2037 (N_2037,N_1978,N_1899);
nor U2038 (N_2038,N_1989,N_1903);
and U2039 (N_2039,N_1964,N_1905);
and U2040 (N_2040,N_1934,N_1933);
or U2041 (N_2041,N_1885,N_1891);
nor U2042 (N_2042,N_1896,N_1953);
or U2043 (N_2043,N_1981,N_1942);
nor U2044 (N_2044,N_1918,N_1980);
nand U2045 (N_2045,N_1973,N_1970);
nand U2046 (N_2046,N_1965,N_1938);
xor U2047 (N_2047,N_1912,N_1914);
nand U2048 (N_2048,N_1957,N_1932);
nor U2049 (N_2049,N_1907,N_1898);
nand U2050 (N_2050,N_1880,N_1922);
and U2051 (N_2051,N_1902,N_1920);
nand U2052 (N_2052,N_1955,N_1991);
nor U2053 (N_2053,N_1893,N_1971);
xnor U2054 (N_2054,N_1979,N_1959);
nand U2055 (N_2055,N_1984,N_1967);
nor U2056 (N_2056,N_1961,N_1994);
or U2057 (N_2057,N_1949,N_1901);
or U2058 (N_2058,N_1881,N_1950);
xnor U2059 (N_2059,N_1954,N_1997);
nor U2060 (N_2060,N_1987,N_1929);
xor U2061 (N_2061,N_1986,N_1988);
or U2062 (N_2062,N_1990,N_1909);
nand U2063 (N_2063,N_1912,N_1945);
and U2064 (N_2064,N_1877,N_1891);
xor U2065 (N_2065,N_1909,N_1904);
or U2066 (N_2066,N_1958,N_1985);
nand U2067 (N_2067,N_1918,N_1884);
and U2068 (N_2068,N_1941,N_1908);
nor U2069 (N_2069,N_1972,N_1913);
or U2070 (N_2070,N_1950,N_1928);
and U2071 (N_2071,N_1958,N_1928);
nor U2072 (N_2072,N_1985,N_1880);
nor U2073 (N_2073,N_1907,N_1969);
nand U2074 (N_2074,N_1940,N_1898);
nor U2075 (N_2075,N_1899,N_1919);
or U2076 (N_2076,N_1937,N_1901);
and U2077 (N_2077,N_1907,N_1998);
and U2078 (N_2078,N_1972,N_1958);
nand U2079 (N_2079,N_1984,N_1929);
xor U2080 (N_2080,N_1901,N_1975);
and U2081 (N_2081,N_1972,N_1888);
and U2082 (N_2082,N_1970,N_1958);
nor U2083 (N_2083,N_1899,N_1972);
and U2084 (N_2084,N_1956,N_1925);
nand U2085 (N_2085,N_1962,N_1937);
or U2086 (N_2086,N_1944,N_1993);
nand U2087 (N_2087,N_1886,N_1884);
xnor U2088 (N_2088,N_1974,N_1994);
or U2089 (N_2089,N_1927,N_1905);
xor U2090 (N_2090,N_1949,N_1954);
and U2091 (N_2091,N_1924,N_1969);
or U2092 (N_2092,N_1964,N_1886);
nand U2093 (N_2093,N_1972,N_1944);
and U2094 (N_2094,N_1882,N_1876);
nand U2095 (N_2095,N_1986,N_1922);
xnor U2096 (N_2096,N_1993,N_1903);
or U2097 (N_2097,N_1888,N_1940);
xor U2098 (N_2098,N_1986,N_1930);
and U2099 (N_2099,N_1879,N_1907);
or U2100 (N_2100,N_1968,N_1875);
nand U2101 (N_2101,N_1919,N_1978);
xor U2102 (N_2102,N_1906,N_1876);
nand U2103 (N_2103,N_1899,N_1970);
and U2104 (N_2104,N_1935,N_1959);
nor U2105 (N_2105,N_1931,N_1943);
or U2106 (N_2106,N_1945,N_1959);
or U2107 (N_2107,N_1940,N_1982);
nand U2108 (N_2108,N_1897,N_1917);
or U2109 (N_2109,N_1890,N_1936);
and U2110 (N_2110,N_1942,N_1949);
nand U2111 (N_2111,N_1969,N_1938);
nand U2112 (N_2112,N_1913,N_1935);
or U2113 (N_2113,N_1948,N_1892);
xnor U2114 (N_2114,N_1931,N_1907);
or U2115 (N_2115,N_1914,N_1890);
nor U2116 (N_2116,N_1987,N_1934);
xnor U2117 (N_2117,N_1926,N_1927);
or U2118 (N_2118,N_1916,N_1884);
nor U2119 (N_2119,N_1883,N_1990);
or U2120 (N_2120,N_1998,N_1896);
nand U2121 (N_2121,N_1916,N_1957);
xor U2122 (N_2122,N_1938,N_1988);
nor U2123 (N_2123,N_1963,N_1902);
nand U2124 (N_2124,N_1979,N_1980);
xor U2125 (N_2125,N_2057,N_2117);
and U2126 (N_2126,N_2035,N_2038);
and U2127 (N_2127,N_2058,N_2104);
or U2128 (N_2128,N_2121,N_2073);
or U2129 (N_2129,N_2017,N_2026);
xor U2130 (N_2130,N_2048,N_2109);
nand U2131 (N_2131,N_2071,N_2068);
or U2132 (N_2132,N_2005,N_2074);
or U2133 (N_2133,N_2039,N_2041);
or U2134 (N_2134,N_2077,N_2010);
nor U2135 (N_2135,N_2037,N_2032);
and U2136 (N_2136,N_2042,N_2079);
and U2137 (N_2137,N_2021,N_2024);
xnor U2138 (N_2138,N_2007,N_2112);
nor U2139 (N_2139,N_2011,N_2034);
xnor U2140 (N_2140,N_2056,N_2108);
xor U2141 (N_2141,N_2008,N_2022);
nor U2142 (N_2142,N_2050,N_2031);
and U2143 (N_2143,N_2089,N_2070);
nand U2144 (N_2144,N_2098,N_2114);
or U2145 (N_2145,N_2009,N_2015);
or U2146 (N_2146,N_2036,N_2063);
nand U2147 (N_2147,N_2113,N_2023);
and U2148 (N_2148,N_2103,N_2019);
and U2149 (N_2149,N_2067,N_2069);
and U2150 (N_2150,N_2004,N_2027);
or U2151 (N_2151,N_2118,N_2093);
or U2152 (N_2152,N_2001,N_2072);
or U2153 (N_2153,N_2013,N_2096);
and U2154 (N_2154,N_2075,N_2055);
xor U2155 (N_2155,N_2030,N_2084);
xor U2156 (N_2156,N_2095,N_2020);
or U2157 (N_2157,N_2062,N_2124);
and U2158 (N_2158,N_2045,N_2101);
or U2159 (N_2159,N_2080,N_2086);
xor U2160 (N_2160,N_2082,N_2116);
or U2161 (N_2161,N_2060,N_2014);
nor U2162 (N_2162,N_2091,N_2046);
xor U2163 (N_2163,N_2043,N_2049);
nand U2164 (N_2164,N_2090,N_2000);
nor U2165 (N_2165,N_2025,N_2053);
and U2166 (N_2166,N_2081,N_2012);
and U2167 (N_2167,N_2065,N_2044);
or U2168 (N_2168,N_2115,N_2119);
nand U2169 (N_2169,N_2102,N_2106);
nand U2170 (N_2170,N_2123,N_2122);
and U2171 (N_2171,N_2110,N_2016);
nor U2172 (N_2172,N_2051,N_2052);
and U2173 (N_2173,N_2083,N_2054);
or U2174 (N_2174,N_2120,N_2100);
or U2175 (N_2175,N_2107,N_2087);
nor U2176 (N_2176,N_2040,N_2076);
xor U2177 (N_2177,N_2006,N_2111);
nand U2178 (N_2178,N_2059,N_2064);
xor U2179 (N_2179,N_2097,N_2094);
or U2180 (N_2180,N_2003,N_2061);
or U2181 (N_2181,N_2033,N_2018);
nor U2182 (N_2182,N_2099,N_2047);
and U2183 (N_2183,N_2105,N_2029);
xnor U2184 (N_2184,N_2085,N_2088);
nand U2185 (N_2185,N_2028,N_2092);
xnor U2186 (N_2186,N_2066,N_2078);
and U2187 (N_2187,N_2002,N_2085);
xnor U2188 (N_2188,N_2083,N_2110);
or U2189 (N_2189,N_2007,N_2074);
nor U2190 (N_2190,N_2068,N_2053);
nor U2191 (N_2191,N_2030,N_2044);
and U2192 (N_2192,N_2059,N_2022);
nor U2193 (N_2193,N_2085,N_2055);
or U2194 (N_2194,N_2118,N_2007);
nand U2195 (N_2195,N_2058,N_2091);
nor U2196 (N_2196,N_2031,N_2106);
nand U2197 (N_2197,N_2043,N_2067);
nor U2198 (N_2198,N_2119,N_2071);
or U2199 (N_2199,N_2016,N_2022);
or U2200 (N_2200,N_2083,N_2027);
and U2201 (N_2201,N_2019,N_2056);
and U2202 (N_2202,N_2119,N_2094);
or U2203 (N_2203,N_2067,N_2030);
xor U2204 (N_2204,N_2055,N_2106);
and U2205 (N_2205,N_2046,N_2064);
nand U2206 (N_2206,N_2039,N_2060);
or U2207 (N_2207,N_2007,N_2073);
nor U2208 (N_2208,N_2054,N_2096);
xor U2209 (N_2209,N_2052,N_2041);
or U2210 (N_2210,N_2030,N_2057);
nand U2211 (N_2211,N_2067,N_2105);
nand U2212 (N_2212,N_2039,N_2115);
and U2213 (N_2213,N_2075,N_2042);
nor U2214 (N_2214,N_2085,N_2036);
or U2215 (N_2215,N_2046,N_2045);
nand U2216 (N_2216,N_2113,N_2056);
nor U2217 (N_2217,N_2015,N_2083);
or U2218 (N_2218,N_2118,N_2016);
xor U2219 (N_2219,N_2118,N_2021);
nand U2220 (N_2220,N_2041,N_2048);
nand U2221 (N_2221,N_2015,N_2058);
xnor U2222 (N_2222,N_2091,N_2055);
and U2223 (N_2223,N_2006,N_2016);
and U2224 (N_2224,N_2028,N_2045);
xnor U2225 (N_2225,N_2116,N_2075);
nand U2226 (N_2226,N_2039,N_2069);
nor U2227 (N_2227,N_2042,N_2007);
or U2228 (N_2228,N_2050,N_2088);
nor U2229 (N_2229,N_2094,N_2046);
nand U2230 (N_2230,N_2096,N_2093);
and U2231 (N_2231,N_2003,N_2065);
xor U2232 (N_2232,N_2071,N_2016);
nor U2233 (N_2233,N_2081,N_2088);
and U2234 (N_2234,N_2095,N_2051);
and U2235 (N_2235,N_2087,N_2024);
nor U2236 (N_2236,N_2114,N_2011);
or U2237 (N_2237,N_2036,N_2031);
and U2238 (N_2238,N_2032,N_2014);
nand U2239 (N_2239,N_2089,N_2078);
nand U2240 (N_2240,N_2120,N_2028);
and U2241 (N_2241,N_2057,N_2001);
xnor U2242 (N_2242,N_2116,N_2016);
or U2243 (N_2243,N_2063,N_2062);
nand U2244 (N_2244,N_2118,N_2108);
or U2245 (N_2245,N_2073,N_2113);
nor U2246 (N_2246,N_2000,N_2066);
and U2247 (N_2247,N_2050,N_2097);
nand U2248 (N_2248,N_2041,N_2008);
or U2249 (N_2249,N_2057,N_2077);
nand U2250 (N_2250,N_2189,N_2242);
xnor U2251 (N_2251,N_2174,N_2218);
xor U2252 (N_2252,N_2248,N_2201);
xor U2253 (N_2253,N_2219,N_2136);
nand U2254 (N_2254,N_2147,N_2211);
nor U2255 (N_2255,N_2150,N_2169);
or U2256 (N_2256,N_2173,N_2246);
nand U2257 (N_2257,N_2153,N_2166);
nor U2258 (N_2258,N_2234,N_2209);
nand U2259 (N_2259,N_2133,N_2208);
nand U2260 (N_2260,N_2148,N_2142);
xnor U2261 (N_2261,N_2157,N_2229);
nand U2262 (N_2262,N_2156,N_2154);
nor U2263 (N_2263,N_2160,N_2212);
nor U2264 (N_2264,N_2214,N_2158);
nand U2265 (N_2265,N_2241,N_2193);
nand U2266 (N_2266,N_2195,N_2131);
xor U2267 (N_2267,N_2141,N_2237);
nor U2268 (N_2268,N_2197,N_2172);
nand U2269 (N_2269,N_2217,N_2177);
and U2270 (N_2270,N_2199,N_2170);
xor U2271 (N_2271,N_2162,N_2216);
nand U2272 (N_2272,N_2125,N_2227);
nand U2273 (N_2273,N_2207,N_2221);
nor U2274 (N_2274,N_2181,N_2178);
or U2275 (N_2275,N_2231,N_2192);
or U2276 (N_2276,N_2180,N_2206);
nor U2277 (N_2277,N_2130,N_2182);
and U2278 (N_2278,N_2168,N_2245);
and U2279 (N_2279,N_2188,N_2244);
and U2280 (N_2280,N_2224,N_2249);
xor U2281 (N_2281,N_2210,N_2196);
xnor U2282 (N_2282,N_2179,N_2235);
nor U2283 (N_2283,N_2167,N_2161);
and U2284 (N_2284,N_2146,N_2137);
and U2285 (N_2285,N_2190,N_2225);
and U2286 (N_2286,N_2238,N_2134);
nor U2287 (N_2287,N_2194,N_2232);
nand U2288 (N_2288,N_2139,N_2163);
or U2289 (N_2289,N_2215,N_2223);
or U2290 (N_2290,N_2191,N_2183);
nor U2291 (N_2291,N_2144,N_2220);
and U2292 (N_2292,N_2155,N_2203);
and U2293 (N_2293,N_2135,N_2205);
nor U2294 (N_2294,N_2247,N_2202);
or U2295 (N_2295,N_2151,N_2140);
and U2296 (N_2296,N_2222,N_2145);
nand U2297 (N_2297,N_2186,N_2236);
nor U2298 (N_2298,N_2226,N_2243);
and U2299 (N_2299,N_2176,N_2171);
nand U2300 (N_2300,N_2138,N_2230);
xor U2301 (N_2301,N_2187,N_2126);
or U2302 (N_2302,N_2184,N_2228);
or U2303 (N_2303,N_2233,N_2159);
xnor U2304 (N_2304,N_2127,N_2149);
xnor U2305 (N_2305,N_2239,N_2143);
xor U2306 (N_2306,N_2200,N_2240);
nor U2307 (N_2307,N_2204,N_2129);
nand U2308 (N_2308,N_2152,N_2175);
nor U2309 (N_2309,N_2128,N_2165);
nand U2310 (N_2310,N_2198,N_2213);
xnor U2311 (N_2311,N_2185,N_2132);
xnor U2312 (N_2312,N_2164,N_2246);
nand U2313 (N_2313,N_2159,N_2135);
and U2314 (N_2314,N_2228,N_2164);
nand U2315 (N_2315,N_2163,N_2136);
and U2316 (N_2316,N_2211,N_2197);
xor U2317 (N_2317,N_2160,N_2135);
or U2318 (N_2318,N_2203,N_2128);
or U2319 (N_2319,N_2206,N_2132);
nor U2320 (N_2320,N_2223,N_2246);
and U2321 (N_2321,N_2145,N_2237);
xnor U2322 (N_2322,N_2160,N_2174);
xor U2323 (N_2323,N_2218,N_2244);
and U2324 (N_2324,N_2194,N_2218);
or U2325 (N_2325,N_2221,N_2174);
and U2326 (N_2326,N_2171,N_2244);
nor U2327 (N_2327,N_2145,N_2133);
or U2328 (N_2328,N_2200,N_2131);
and U2329 (N_2329,N_2246,N_2155);
nand U2330 (N_2330,N_2216,N_2241);
nor U2331 (N_2331,N_2166,N_2133);
or U2332 (N_2332,N_2144,N_2234);
xor U2333 (N_2333,N_2146,N_2172);
and U2334 (N_2334,N_2153,N_2242);
and U2335 (N_2335,N_2239,N_2200);
xnor U2336 (N_2336,N_2156,N_2186);
nor U2337 (N_2337,N_2187,N_2199);
or U2338 (N_2338,N_2176,N_2136);
nand U2339 (N_2339,N_2159,N_2171);
nor U2340 (N_2340,N_2232,N_2156);
or U2341 (N_2341,N_2133,N_2148);
and U2342 (N_2342,N_2198,N_2212);
and U2343 (N_2343,N_2131,N_2213);
or U2344 (N_2344,N_2148,N_2245);
or U2345 (N_2345,N_2229,N_2239);
or U2346 (N_2346,N_2142,N_2140);
or U2347 (N_2347,N_2140,N_2138);
nor U2348 (N_2348,N_2213,N_2216);
or U2349 (N_2349,N_2228,N_2179);
and U2350 (N_2350,N_2125,N_2226);
and U2351 (N_2351,N_2198,N_2149);
xor U2352 (N_2352,N_2183,N_2149);
and U2353 (N_2353,N_2130,N_2240);
nor U2354 (N_2354,N_2202,N_2222);
nand U2355 (N_2355,N_2130,N_2165);
or U2356 (N_2356,N_2223,N_2179);
or U2357 (N_2357,N_2132,N_2187);
and U2358 (N_2358,N_2125,N_2190);
or U2359 (N_2359,N_2231,N_2223);
and U2360 (N_2360,N_2131,N_2228);
nand U2361 (N_2361,N_2222,N_2244);
nor U2362 (N_2362,N_2158,N_2204);
xor U2363 (N_2363,N_2241,N_2137);
or U2364 (N_2364,N_2239,N_2184);
xor U2365 (N_2365,N_2170,N_2157);
or U2366 (N_2366,N_2233,N_2169);
nand U2367 (N_2367,N_2186,N_2247);
xnor U2368 (N_2368,N_2157,N_2189);
nor U2369 (N_2369,N_2170,N_2126);
xor U2370 (N_2370,N_2203,N_2227);
nand U2371 (N_2371,N_2157,N_2135);
nor U2372 (N_2372,N_2178,N_2144);
xor U2373 (N_2373,N_2215,N_2184);
and U2374 (N_2374,N_2167,N_2173);
xor U2375 (N_2375,N_2261,N_2370);
or U2376 (N_2376,N_2311,N_2256);
and U2377 (N_2377,N_2282,N_2274);
xnor U2378 (N_2378,N_2342,N_2371);
nor U2379 (N_2379,N_2255,N_2362);
xor U2380 (N_2380,N_2366,N_2338);
nor U2381 (N_2381,N_2291,N_2333);
or U2382 (N_2382,N_2273,N_2324);
nand U2383 (N_2383,N_2331,N_2360);
nand U2384 (N_2384,N_2369,N_2262);
or U2385 (N_2385,N_2374,N_2251);
nand U2386 (N_2386,N_2301,N_2364);
nand U2387 (N_2387,N_2326,N_2264);
or U2388 (N_2388,N_2272,N_2271);
and U2389 (N_2389,N_2351,N_2354);
or U2390 (N_2390,N_2340,N_2295);
nor U2391 (N_2391,N_2277,N_2339);
nor U2392 (N_2392,N_2258,N_2266);
or U2393 (N_2393,N_2283,N_2313);
nor U2394 (N_2394,N_2315,N_2341);
nand U2395 (N_2395,N_2335,N_2267);
nor U2396 (N_2396,N_2358,N_2281);
nand U2397 (N_2397,N_2307,N_2353);
nand U2398 (N_2398,N_2348,N_2363);
nand U2399 (N_2399,N_2308,N_2280);
nor U2400 (N_2400,N_2328,N_2317);
or U2401 (N_2401,N_2349,N_2357);
or U2402 (N_2402,N_2293,N_2304);
xnor U2403 (N_2403,N_2289,N_2290);
nor U2404 (N_2404,N_2260,N_2329);
nor U2405 (N_2405,N_2323,N_2361);
nand U2406 (N_2406,N_2337,N_2309);
xor U2407 (N_2407,N_2316,N_2314);
nor U2408 (N_2408,N_2296,N_2327);
and U2409 (N_2409,N_2343,N_2318);
nor U2410 (N_2410,N_2285,N_2286);
or U2411 (N_2411,N_2284,N_2345);
or U2412 (N_2412,N_2250,N_2352);
xor U2413 (N_2413,N_2321,N_2319);
or U2414 (N_2414,N_2299,N_2263);
nand U2415 (N_2415,N_2330,N_2300);
or U2416 (N_2416,N_2305,N_2367);
or U2417 (N_2417,N_2275,N_2325);
nor U2418 (N_2418,N_2346,N_2372);
xnor U2419 (N_2419,N_2254,N_2334);
nor U2420 (N_2420,N_2297,N_2344);
xor U2421 (N_2421,N_2292,N_2332);
nor U2422 (N_2422,N_2310,N_2359);
nor U2423 (N_2423,N_2302,N_2350);
nand U2424 (N_2424,N_2355,N_2252);
or U2425 (N_2425,N_2253,N_2322);
nand U2426 (N_2426,N_2294,N_2312);
nand U2427 (N_2427,N_2270,N_2336);
nand U2428 (N_2428,N_2276,N_2320);
and U2429 (N_2429,N_2269,N_2265);
nor U2430 (N_2430,N_2303,N_2365);
and U2431 (N_2431,N_2356,N_2259);
or U2432 (N_2432,N_2298,N_2257);
xor U2433 (N_2433,N_2306,N_2268);
nand U2434 (N_2434,N_2278,N_2288);
xnor U2435 (N_2435,N_2368,N_2373);
or U2436 (N_2436,N_2287,N_2279);
and U2437 (N_2437,N_2347,N_2275);
nand U2438 (N_2438,N_2290,N_2311);
or U2439 (N_2439,N_2343,N_2322);
and U2440 (N_2440,N_2362,N_2329);
nand U2441 (N_2441,N_2254,N_2273);
xor U2442 (N_2442,N_2323,N_2304);
xnor U2443 (N_2443,N_2355,N_2259);
nor U2444 (N_2444,N_2264,N_2278);
and U2445 (N_2445,N_2270,N_2343);
xnor U2446 (N_2446,N_2365,N_2347);
nand U2447 (N_2447,N_2312,N_2297);
and U2448 (N_2448,N_2268,N_2355);
nor U2449 (N_2449,N_2319,N_2253);
or U2450 (N_2450,N_2359,N_2268);
nand U2451 (N_2451,N_2283,N_2360);
or U2452 (N_2452,N_2346,N_2352);
xnor U2453 (N_2453,N_2263,N_2296);
nor U2454 (N_2454,N_2339,N_2317);
and U2455 (N_2455,N_2334,N_2293);
nand U2456 (N_2456,N_2262,N_2294);
or U2457 (N_2457,N_2255,N_2299);
and U2458 (N_2458,N_2348,N_2271);
and U2459 (N_2459,N_2345,N_2279);
nand U2460 (N_2460,N_2293,N_2282);
nand U2461 (N_2461,N_2363,N_2342);
nand U2462 (N_2462,N_2314,N_2318);
xor U2463 (N_2463,N_2269,N_2261);
xor U2464 (N_2464,N_2250,N_2354);
nor U2465 (N_2465,N_2259,N_2335);
nand U2466 (N_2466,N_2284,N_2328);
xnor U2467 (N_2467,N_2271,N_2321);
nor U2468 (N_2468,N_2330,N_2253);
and U2469 (N_2469,N_2294,N_2339);
nor U2470 (N_2470,N_2292,N_2285);
or U2471 (N_2471,N_2292,N_2355);
nor U2472 (N_2472,N_2348,N_2280);
nor U2473 (N_2473,N_2279,N_2281);
and U2474 (N_2474,N_2269,N_2290);
nor U2475 (N_2475,N_2252,N_2342);
xnor U2476 (N_2476,N_2344,N_2260);
nor U2477 (N_2477,N_2352,N_2336);
nand U2478 (N_2478,N_2321,N_2348);
nor U2479 (N_2479,N_2272,N_2250);
nand U2480 (N_2480,N_2264,N_2287);
nand U2481 (N_2481,N_2366,N_2313);
xor U2482 (N_2482,N_2353,N_2283);
xor U2483 (N_2483,N_2250,N_2277);
nor U2484 (N_2484,N_2369,N_2312);
xor U2485 (N_2485,N_2358,N_2285);
and U2486 (N_2486,N_2354,N_2314);
xor U2487 (N_2487,N_2347,N_2364);
xor U2488 (N_2488,N_2337,N_2279);
and U2489 (N_2489,N_2285,N_2351);
nor U2490 (N_2490,N_2339,N_2333);
nand U2491 (N_2491,N_2264,N_2305);
xor U2492 (N_2492,N_2307,N_2332);
nor U2493 (N_2493,N_2349,N_2306);
nand U2494 (N_2494,N_2324,N_2325);
xnor U2495 (N_2495,N_2309,N_2308);
nand U2496 (N_2496,N_2304,N_2371);
xor U2497 (N_2497,N_2357,N_2256);
or U2498 (N_2498,N_2264,N_2355);
and U2499 (N_2499,N_2303,N_2255);
nand U2500 (N_2500,N_2400,N_2449);
or U2501 (N_2501,N_2393,N_2444);
and U2502 (N_2502,N_2466,N_2422);
and U2503 (N_2503,N_2440,N_2410);
nor U2504 (N_2504,N_2386,N_2487);
nor U2505 (N_2505,N_2488,N_2478);
and U2506 (N_2506,N_2416,N_2480);
nand U2507 (N_2507,N_2423,N_2497);
or U2508 (N_2508,N_2431,N_2407);
nand U2509 (N_2509,N_2476,N_2494);
xnor U2510 (N_2510,N_2404,N_2477);
or U2511 (N_2511,N_2489,N_2385);
nand U2512 (N_2512,N_2453,N_2443);
xor U2513 (N_2513,N_2455,N_2495);
xnor U2514 (N_2514,N_2415,N_2380);
or U2515 (N_2515,N_2481,N_2432);
and U2516 (N_2516,N_2475,N_2412);
or U2517 (N_2517,N_2389,N_2468);
xor U2518 (N_2518,N_2445,N_2448);
xor U2519 (N_2519,N_2474,N_2375);
or U2520 (N_2520,N_2485,N_2498);
xor U2521 (N_2521,N_2436,N_2403);
xor U2522 (N_2522,N_2376,N_2438);
xor U2523 (N_2523,N_2429,N_2387);
xnor U2524 (N_2524,N_2428,N_2381);
or U2525 (N_2525,N_2496,N_2461);
nand U2526 (N_2526,N_2441,N_2471);
nand U2527 (N_2527,N_2399,N_2435);
nand U2528 (N_2528,N_2484,N_2452);
or U2529 (N_2529,N_2450,N_2384);
and U2530 (N_2530,N_2382,N_2433);
or U2531 (N_2531,N_2464,N_2437);
nand U2532 (N_2532,N_2397,N_2447);
nand U2533 (N_2533,N_2390,N_2411);
nand U2534 (N_2534,N_2421,N_2413);
nand U2535 (N_2535,N_2420,N_2402);
xnor U2536 (N_2536,N_2378,N_2467);
and U2537 (N_2537,N_2458,N_2459);
xor U2538 (N_2538,N_2479,N_2442);
xor U2539 (N_2539,N_2396,N_2425);
nand U2540 (N_2540,N_2392,N_2388);
and U2541 (N_2541,N_2473,N_2401);
or U2542 (N_2542,N_2446,N_2451);
or U2543 (N_2543,N_2414,N_2398);
or U2544 (N_2544,N_2469,N_2439);
xnor U2545 (N_2545,N_2424,N_2465);
or U2546 (N_2546,N_2430,N_2405);
or U2547 (N_2547,N_2470,N_2492);
or U2548 (N_2548,N_2394,N_2491);
nor U2549 (N_2549,N_2418,N_2427);
nor U2550 (N_2550,N_2457,N_2395);
xnor U2551 (N_2551,N_2377,N_2463);
or U2552 (N_2552,N_2419,N_2462);
xnor U2553 (N_2553,N_2490,N_2472);
nor U2554 (N_2554,N_2456,N_2426);
and U2555 (N_2555,N_2499,N_2379);
or U2556 (N_2556,N_2391,N_2408);
nor U2557 (N_2557,N_2460,N_2482);
xnor U2558 (N_2558,N_2493,N_2486);
xor U2559 (N_2559,N_2383,N_2406);
and U2560 (N_2560,N_2454,N_2417);
and U2561 (N_2561,N_2434,N_2409);
or U2562 (N_2562,N_2483,N_2441);
or U2563 (N_2563,N_2402,N_2430);
nand U2564 (N_2564,N_2411,N_2394);
nand U2565 (N_2565,N_2437,N_2485);
and U2566 (N_2566,N_2445,N_2433);
xor U2567 (N_2567,N_2415,N_2418);
xor U2568 (N_2568,N_2467,N_2452);
xnor U2569 (N_2569,N_2444,N_2496);
nand U2570 (N_2570,N_2475,N_2446);
nor U2571 (N_2571,N_2418,N_2399);
or U2572 (N_2572,N_2394,N_2417);
and U2573 (N_2573,N_2447,N_2418);
xnor U2574 (N_2574,N_2432,N_2436);
xnor U2575 (N_2575,N_2416,N_2460);
xor U2576 (N_2576,N_2474,N_2493);
nand U2577 (N_2577,N_2434,N_2426);
nand U2578 (N_2578,N_2376,N_2403);
xor U2579 (N_2579,N_2469,N_2434);
or U2580 (N_2580,N_2415,N_2458);
nand U2581 (N_2581,N_2450,N_2490);
nand U2582 (N_2582,N_2386,N_2402);
xnor U2583 (N_2583,N_2485,N_2450);
and U2584 (N_2584,N_2463,N_2471);
xor U2585 (N_2585,N_2469,N_2405);
or U2586 (N_2586,N_2477,N_2426);
nand U2587 (N_2587,N_2441,N_2443);
nand U2588 (N_2588,N_2448,N_2489);
nand U2589 (N_2589,N_2460,N_2437);
and U2590 (N_2590,N_2426,N_2484);
or U2591 (N_2591,N_2397,N_2435);
or U2592 (N_2592,N_2383,N_2460);
nand U2593 (N_2593,N_2499,N_2451);
xnor U2594 (N_2594,N_2423,N_2481);
nor U2595 (N_2595,N_2479,N_2385);
or U2596 (N_2596,N_2447,N_2445);
and U2597 (N_2597,N_2408,N_2482);
nand U2598 (N_2598,N_2392,N_2382);
nor U2599 (N_2599,N_2489,N_2479);
xor U2600 (N_2600,N_2480,N_2497);
and U2601 (N_2601,N_2466,N_2393);
or U2602 (N_2602,N_2384,N_2436);
or U2603 (N_2603,N_2439,N_2479);
or U2604 (N_2604,N_2425,N_2397);
xor U2605 (N_2605,N_2434,N_2443);
or U2606 (N_2606,N_2416,N_2465);
nand U2607 (N_2607,N_2465,N_2406);
or U2608 (N_2608,N_2413,N_2455);
or U2609 (N_2609,N_2499,N_2402);
or U2610 (N_2610,N_2436,N_2491);
and U2611 (N_2611,N_2478,N_2494);
xnor U2612 (N_2612,N_2416,N_2466);
or U2613 (N_2613,N_2395,N_2384);
nand U2614 (N_2614,N_2433,N_2463);
nor U2615 (N_2615,N_2421,N_2396);
nand U2616 (N_2616,N_2425,N_2419);
xnor U2617 (N_2617,N_2421,N_2485);
xor U2618 (N_2618,N_2476,N_2433);
nor U2619 (N_2619,N_2454,N_2479);
nor U2620 (N_2620,N_2443,N_2401);
nand U2621 (N_2621,N_2406,N_2451);
nor U2622 (N_2622,N_2457,N_2491);
xor U2623 (N_2623,N_2493,N_2375);
or U2624 (N_2624,N_2411,N_2416);
nor U2625 (N_2625,N_2586,N_2624);
and U2626 (N_2626,N_2551,N_2530);
or U2627 (N_2627,N_2592,N_2547);
xnor U2628 (N_2628,N_2622,N_2503);
or U2629 (N_2629,N_2620,N_2544);
and U2630 (N_2630,N_2571,N_2507);
nor U2631 (N_2631,N_2593,N_2576);
nor U2632 (N_2632,N_2505,N_2603);
and U2633 (N_2633,N_2560,N_2584);
xor U2634 (N_2634,N_2556,N_2545);
or U2635 (N_2635,N_2578,N_2582);
and U2636 (N_2636,N_2595,N_2517);
nor U2637 (N_2637,N_2618,N_2526);
nand U2638 (N_2638,N_2581,N_2562);
or U2639 (N_2639,N_2588,N_2520);
or U2640 (N_2640,N_2510,N_2501);
or U2641 (N_2641,N_2539,N_2527);
or U2642 (N_2642,N_2594,N_2573);
nand U2643 (N_2643,N_2557,N_2522);
and U2644 (N_2644,N_2536,N_2508);
or U2645 (N_2645,N_2533,N_2608);
nor U2646 (N_2646,N_2565,N_2514);
and U2647 (N_2647,N_2612,N_2572);
or U2648 (N_2648,N_2542,N_2596);
xnor U2649 (N_2649,N_2511,N_2583);
nand U2650 (N_2650,N_2504,N_2518);
nor U2651 (N_2651,N_2569,N_2607);
nor U2652 (N_2652,N_2591,N_2552);
or U2653 (N_2653,N_2602,N_2506);
and U2654 (N_2654,N_2528,N_2516);
xor U2655 (N_2655,N_2615,N_2623);
xor U2656 (N_2656,N_2549,N_2609);
nand U2657 (N_2657,N_2540,N_2521);
nand U2658 (N_2658,N_2541,N_2567);
or U2659 (N_2659,N_2587,N_2553);
xnor U2660 (N_2660,N_2513,N_2598);
nand U2661 (N_2661,N_2525,N_2601);
nor U2662 (N_2662,N_2512,N_2577);
xor U2663 (N_2663,N_2606,N_2532);
or U2664 (N_2664,N_2617,N_2574);
nand U2665 (N_2665,N_2589,N_2564);
xnor U2666 (N_2666,N_2531,N_2590);
xnor U2667 (N_2667,N_2509,N_2561);
or U2668 (N_2668,N_2558,N_2563);
and U2669 (N_2669,N_2600,N_2515);
and U2670 (N_2670,N_2579,N_2555);
nand U2671 (N_2671,N_2502,N_2570);
and U2672 (N_2672,N_2604,N_2568);
xor U2673 (N_2673,N_2616,N_2605);
and U2674 (N_2674,N_2524,N_2621);
xor U2675 (N_2675,N_2611,N_2597);
nor U2676 (N_2676,N_2619,N_2566);
and U2677 (N_2677,N_2500,N_2538);
or U2678 (N_2678,N_2559,N_2537);
xor U2679 (N_2679,N_2529,N_2535);
xor U2680 (N_2680,N_2546,N_2523);
nand U2681 (N_2681,N_2534,N_2519);
nor U2682 (N_2682,N_2543,N_2554);
and U2683 (N_2683,N_2599,N_2550);
nor U2684 (N_2684,N_2610,N_2614);
nand U2685 (N_2685,N_2575,N_2580);
and U2686 (N_2686,N_2613,N_2548);
xor U2687 (N_2687,N_2585,N_2519);
or U2688 (N_2688,N_2604,N_2551);
xnor U2689 (N_2689,N_2583,N_2503);
or U2690 (N_2690,N_2540,N_2588);
xnor U2691 (N_2691,N_2525,N_2527);
nand U2692 (N_2692,N_2541,N_2509);
xnor U2693 (N_2693,N_2511,N_2610);
and U2694 (N_2694,N_2589,N_2599);
xor U2695 (N_2695,N_2571,N_2615);
nand U2696 (N_2696,N_2577,N_2599);
and U2697 (N_2697,N_2571,N_2588);
xor U2698 (N_2698,N_2507,N_2553);
and U2699 (N_2699,N_2511,N_2609);
and U2700 (N_2700,N_2515,N_2555);
nand U2701 (N_2701,N_2549,N_2597);
and U2702 (N_2702,N_2543,N_2501);
or U2703 (N_2703,N_2585,N_2522);
xor U2704 (N_2704,N_2511,N_2503);
nor U2705 (N_2705,N_2524,N_2519);
and U2706 (N_2706,N_2593,N_2583);
nand U2707 (N_2707,N_2578,N_2564);
xnor U2708 (N_2708,N_2570,N_2545);
nor U2709 (N_2709,N_2587,N_2610);
xnor U2710 (N_2710,N_2535,N_2528);
nand U2711 (N_2711,N_2588,N_2622);
and U2712 (N_2712,N_2602,N_2541);
xnor U2713 (N_2713,N_2602,N_2595);
nor U2714 (N_2714,N_2524,N_2536);
nor U2715 (N_2715,N_2546,N_2601);
nand U2716 (N_2716,N_2556,N_2608);
nand U2717 (N_2717,N_2557,N_2576);
or U2718 (N_2718,N_2584,N_2585);
and U2719 (N_2719,N_2555,N_2501);
and U2720 (N_2720,N_2538,N_2568);
xnor U2721 (N_2721,N_2522,N_2502);
or U2722 (N_2722,N_2619,N_2617);
and U2723 (N_2723,N_2620,N_2588);
or U2724 (N_2724,N_2575,N_2559);
or U2725 (N_2725,N_2515,N_2558);
nor U2726 (N_2726,N_2553,N_2508);
or U2727 (N_2727,N_2529,N_2554);
nand U2728 (N_2728,N_2558,N_2593);
or U2729 (N_2729,N_2599,N_2553);
xor U2730 (N_2730,N_2572,N_2527);
xor U2731 (N_2731,N_2526,N_2583);
or U2732 (N_2732,N_2586,N_2504);
nor U2733 (N_2733,N_2565,N_2550);
or U2734 (N_2734,N_2540,N_2589);
and U2735 (N_2735,N_2523,N_2500);
and U2736 (N_2736,N_2580,N_2613);
xor U2737 (N_2737,N_2557,N_2578);
nand U2738 (N_2738,N_2531,N_2514);
or U2739 (N_2739,N_2569,N_2553);
or U2740 (N_2740,N_2500,N_2531);
and U2741 (N_2741,N_2541,N_2521);
nor U2742 (N_2742,N_2540,N_2619);
xor U2743 (N_2743,N_2506,N_2594);
nor U2744 (N_2744,N_2581,N_2620);
nand U2745 (N_2745,N_2549,N_2538);
nand U2746 (N_2746,N_2535,N_2559);
and U2747 (N_2747,N_2580,N_2593);
or U2748 (N_2748,N_2503,N_2621);
xnor U2749 (N_2749,N_2593,N_2570);
and U2750 (N_2750,N_2735,N_2740);
nand U2751 (N_2751,N_2681,N_2637);
xor U2752 (N_2752,N_2744,N_2687);
xor U2753 (N_2753,N_2738,N_2633);
and U2754 (N_2754,N_2673,N_2666);
and U2755 (N_2755,N_2686,N_2685);
and U2756 (N_2756,N_2711,N_2705);
xnor U2757 (N_2757,N_2677,N_2627);
xnor U2758 (N_2758,N_2728,N_2638);
nand U2759 (N_2759,N_2642,N_2650);
nor U2760 (N_2760,N_2718,N_2732);
nand U2761 (N_2761,N_2653,N_2714);
nand U2762 (N_2762,N_2658,N_2631);
xnor U2763 (N_2763,N_2663,N_2662);
or U2764 (N_2764,N_2639,N_2668);
nand U2765 (N_2765,N_2641,N_2743);
nor U2766 (N_2766,N_2747,N_2645);
nor U2767 (N_2767,N_2630,N_2716);
xor U2768 (N_2768,N_2721,N_2731);
or U2769 (N_2769,N_2706,N_2659);
and U2770 (N_2770,N_2726,N_2691);
xor U2771 (N_2771,N_2665,N_2644);
and U2772 (N_2772,N_2676,N_2683);
xor U2773 (N_2773,N_2736,N_2719);
or U2774 (N_2774,N_2697,N_2727);
or U2775 (N_2775,N_2640,N_2748);
nor U2776 (N_2776,N_2674,N_2700);
nand U2777 (N_2777,N_2635,N_2724);
xor U2778 (N_2778,N_2657,N_2746);
nand U2779 (N_2779,N_2648,N_2712);
nand U2780 (N_2780,N_2670,N_2690);
nor U2781 (N_2781,N_2729,N_2698);
or U2782 (N_2782,N_2625,N_2632);
or U2783 (N_2783,N_2660,N_2628);
xor U2784 (N_2784,N_2655,N_2723);
nand U2785 (N_2785,N_2679,N_2694);
xnor U2786 (N_2786,N_2702,N_2634);
xor U2787 (N_2787,N_2717,N_2737);
nand U2788 (N_2788,N_2643,N_2722);
and U2789 (N_2789,N_2693,N_2654);
nand U2790 (N_2790,N_2667,N_2651);
nand U2791 (N_2791,N_2696,N_2739);
nor U2792 (N_2792,N_2725,N_2652);
xnor U2793 (N_2793,N_2675,N_2671);
and U2794 (N_2794,N_2742,N_2745);
nor U2795 (N_2795,N_2709,N_2749);
xnor U2796 (N_2796,N_2710,N_2664);
xor U2797 (N_2797,N_2661,N_2715);
nor U2798 (N_2798,N_2730,N_2741);
nor U2799 (N_2799,N_2636,N_2713);
nand U2800 (N_2800,N_2704,N_2695);
nand U2801 (N_2801,N_2626,N_2699);
nand U2802 (N_2802,N_2669,N_2720);
nor U2803 (N_2803,N_2707,N_2701);
nand U2804 (N_2804,N_2689,N_2649);
xnor U2805 (N_2805,N_2629,N_2733);
xor U2806 (N_2806,N_2672,N_2656);
nand U2807 (N_2807,N_2684,N_2646);
nor U2808 (N_2808,N_2680,N_2703);
xor U2809 (N_2809,N_2692,N_2647);
or U2810 (N_2810,N_2682,N_2678);
nor U2811 (N_2811,N_2708,N_2688);
nor U2812 (N_2812,N_2734,N_2705);
xor U2813 (N_2813,N_2744,N_2723);
or U2814 (N_2814,N_2705,N_2746);
nor U2815 (N_2815,N_2633,N_2707);
xor U2816 (N_2816,N_2625,N_2673);
nor U2817 (N_2817,N_2709,N_2716);
xor U2818 (N_2818,N_2666,N_2683);
nor U2819 (N_2819,N_2647,N_2698);
nand U2820 (N_2820,N_2708,N_2652);
nand U2821 (N_2821,N_2719,N_2639);
nand U2822 (N_2822,N_2731,N_2662);
nor U2823 (N_2823,N_2739,N_2676);
xnor U2824 (N_2824,N_2648,N_2690);
nand U2825 (N_2825,N_2671,N_2718);
or U2826 (N_2826,N_2650,N_2643);
xor U2827 (N_2827,N_2718,N_2692);
nand U2828 (N_2828,N_2661,N_2740);
or U2829 (N_2829,N_2717,N_2721);
nand U2830 (N_2830,N_2628,N_2671);
nand U2831 (N_2831,N_2626,N_2640);
and U2832 (N_2832,N_2721,N_2696);
nand U2833 (N_2833,N_2677,N_2685);
nor U2834 (N_2834,N_2689,N_2703);
xor U2835 (N_2835,N_2692,N_2737);
or U2836 (N_2836,N_2716,N_2654);
nor U2837 (N_2837,N_2737,N_2670);
xnor U2838 (N_2838,N_2659,N_2648);
or U2839 (N_2839,N_2652,N_2625);
and U2840 (N_2840,N_2718,N_2638);
nand U2841 (N_2841,N_2716,N_2635);
nand U2842 (N_2842,N_2677,N_2701);
xor U2843 (N_2843,N_2637,N_2641);
and U2844 (N_2844,N_2703,N_2668);
xnor U2845 (N_2845,N_2662,N_2656);
nand U2846 (N_2846,N_2703,N_2666);
nand U2847 (N_2847,N_2669,N_2667);
nor U2848 (N_2848,N_2729,N_2649);
or U2849 (N_2849,N_2678,N_2729);
and U2850 (N_2850,N_2730,N_2703);
and U2851 (N_2851,N_2693,N_2648);
nand U2852 (N_2852,N_2691,N_2727);
nor U2853 (N_2853,N_2745,N_2697);
nor U2854 (N_2854,N_2749,N_2641);
and U2855 (N_2855,N_2663,N_2669);
nor U2856 (N_2856,N_2664,N_2638);
and U2857 (N_2857,N_2740,N_2663);
nand U2858 (N_2858,N_2692,N_2676);
nor U2859 (N_2859,N_2651,N_2647);
and U2860 (N_2860,N_2749,N_2743);
nor U2861 (N_2861,N_2683,N_2634);
or U2862 (N_2862,N_2633,N_2644);
or U2863 (N_2863,N_2698,N_2742);
or U2864 (N_2864,N_2629,N_2699);
or U2865 (N_2865,N_2746,N_2667);
nor U2866 (N_2866,N_2706,N_2642);
nand U2867 (N_2867,N_2749,N_2715);
nor U2868 (N_2868,N_2639,N_2650);
nand U2869 (N_2869,N_2691,N_2677);
xnor U2870 (N_2870,N_2642,N_2713);
or U2871 (N_2871,N_2720,N_2738);
and U2872 (N_2872,N_2745,N_2645);
nor U2873 (N_2873,N_2694,N_2717);
or U2874 (N_2874,N_2684,N_2690);
and U2875 (N_2875,N_2774,N_2843);
xnor U2876 (N_2876,N_2861,N_2845);
or U2877 (N_2877,N_2814,N_2804);
and U2878 (N_2878,N_2852,N_2752);
nor U2879 (N_2879,N_2794,N_2805);
or U2880 (N_2880,N_2754,N_2821);
or U2881 (N_2881,N_2838,N_2820);
nand U2882 (N_2882,N_2818,N_2851);
xnor U2883 (N_2883,N_2860,N_2862);
or U2884 (N_2884,N_2767,N_2866);
nand U2885 (N_2885,N_2759,N_2809);
and U2886 (N_2886,N_2757,N_2783);
or U2887 (N_2887,N_2836,N_2828);
nand U2888 (N_2888,N_2787,N_2858);
xor U2889 (N_2889,N_2784,N_2786);
or U2890 (N_2890,N_2863,N_2793);
and U2891 (N_2891,N_2808,N_2856);
xor U2892 (N_2892,N_2773,N_2769);
or U2893 (N_2893,N_2825,N_2842);
or U2894 (N_2894,N_2768,N_2864);
xnor U2895 (N_2895,N_2796,N_2791);
and U2896 (N_2896,N_2833,N_2801);
xnor U2897 (N_2897,N_2841,N_2819);
xnor U2898 (N_2898,N_2874,N_2868);
xnor U2899 (N_2899,N_2853,N_2830);
nand U2900 (N_2900,N_2800,N_2849);
xor U2901 (N_2901,N_2857,N_2839);
nor U2902 (N_2902,N_2823,N_2778);
or U2903 (N_2903,N_2873,N_2846);
nor U2904 (N_2904,N_2770,N_2766);
xor U2905 (N_2905,N_2762,N_2835);
or U2906 (N_2906,N_2806,N_2832);
nor U2907 (N_2907,N_2850,N_2782);
and U2908 (N_2908,N_2771,N_2837);
nand U2909 (N_2909,N_2781,N_2798);
or U2910 (N_2910,N_2807,N_2865);
nand U2911 (N_2911,N_2854,N_2867);
and U2912 (N_2912,N_2790,N_2872);
nand U2913 (N_2913,N_2760,N_2789);
xor U2914 (N_2914,N_2755,N_2815);
or U2915 (N_2915,N_2812,N_2817);
or U2916 (N_2916,N_2871,N_2840);
or U2917 (N_2917,N_2855,N_2848);
xor U2918 (N_2918,N_2761,N_2772);
or U2919 (N_2919,N_2829,N_2826);
xnor U2920 (N_2920,N_2780,N_2816);
nand U2921 (N_2921,N_2803,N_2777);
nand U2922 (N_2922,N_2797,N_2870);
and U2923 (N_2923,N_2756,N_2810);
and U2924 (N_2924,N_2834,N_2824);
or U2925 (N_2925,N_2859,N_2822);
nor U2926 (N_2926,N_2827,N_2844);
nor U2927 (N_2927,N_2785,N_2847);
nor U2928 (N_2928,N_2802,N_2775);
xnor U2929 (N_2929,N_2750,N_2779);
or U2930 (N_2930,N_2765,N_2776);
nand U2931 (N_2931,N_2831,N_2788);
xor U2932 (N_2932,N_2795,N_2753);
xor U2933 (N_2933,N_2811,N_2869);
nor U2934 (N_2934,N_2763,N_2799);
xor U2935 (N_2935,N_2813,N_2758);
or U2936 (N_2936,N_2764,N_2792);
and U2937 (N_2937,N_2751,N_2773);
nor U2938 (N_2938,N_2752,N_2857);
nand U2939 (N_2939,N_2871,N_2854);
and U2940 (N_2940,N_2793,N_2812);
or U2941 (N_2941,N_2838,N_2789);
nand U2942 (N_2942,N_2830,N_2806);
nor U2943 (N_2943,N_2816,N_2840);
nor U2944 (N_2944,N_2802,N_2827);
nor U2945 (N_2945,N_2804,N_2841);
nand U2946 (N_2946,N_2813,N_2852);
xnor U2947 (N_2947,N_2756,N_2801);
nand U2948 (N_2948,N_2773,N_2758);
and U2949 (N_2949,N_2830,N_2804);
and U2950 (N_2950,N_2803,N_2805);
nand U2951 (N_2951,N_2773,N_2872);
and U2952 (N_2952,N_2848,N_2812);
nand U2953 (N_2953,N_2852,N_2807);
nor U2954 (N_2954,N_2852,N_2831);
xnor U2955 (N_2955,N_2777,N_2760);
and U2956 (N_2956,N_2815,N_2750);
or U2957 (N_2957,N_2869,N_2820);
and U2958 (N_2958,N_2801,N_2860);
nor U2959 (N_2959,N_2824,N_2868);
or U2960 (N_2960,N_2820,N_2871);
or U2961 (N_2961,N_2836,N_2799);
and U2962 (N_2962,N_2861,N_2841);
or U2963 (N_2963,N_2832,N_2758);
and U2964 (N_2964,N_2821,N_2778);
and U2965 (N_2965,N_2760,N_2758);
and U2966 (N_2966,N_2786,N_2761);
nand U2967 (N_2967,N_2855,N_2832);
nand U2968 (N_2968,N_2771,N_2770);
nand U2969 (N_2969,N_2836,N_2873);
xnor U2970 (N_2970,N_2840,N_2776);
or U2971 (N_2971,N_2801,N_2857);
and U2972 (N_2972,N_2812,N_2752);
and U2973 (N_2973,N_2783,N_2764);
or U2974 (N_2974,N_2792,N_2761);
nor U2975 (N_2975,N_2821,N_2869);
nor U2976 (N_2976,N_2827,N_2818);
nor U2977 (N_2977,N_2794,N_2799);
xor U2978 (N_2978,N_2803,N_2754);
and U2979 (N_2979,N_2792,N_2756);
xnor U2980 (N_2980,N_2832,N_2866);
and U2981 (N_2981,N_2820,N_2761);
nand U2982 (N_2982,N_2837,N_2814);
or U2983 (N_2983,N_2873,N_2796);
nand U2984 (N_2984,N_2824,N_2783);
and U2985 (N_2985,N_2831,N_2829);
or U2986 (N_2986,N_2778,N_2803);
or U2987 (N_2987,N_2846,N_2847);
or U2988 (N_2988,N_2761,N_2785);
nand U2989 (N_2989,N_2839,N_2830);
or U2990 (N_2990,N_2804,N_2845);
nor U2991 (N_2991,N_2792,N_2774);
nor U2992 (N_2992,N_2820,N_2822);
xor U2993 (N_2993,N_2765,N_2791);
or U2994 (N_2994,N_2847,N_2788);
xnor U2995 (N_2995,N_2750,N_2855);
or U2996 (N_2996,N_2765,N_2757);
xor U2997 (N_2997,N_2868,N_2775);
xor U2998 (N_2998,N_2808,N_2838);
nor U2999 (N_2999,N_2845,N_2859);
and U3000 (N_3000,N_2967,N_2896);
nor U3001 (N_3001,N_2897,N_2937);
nor U3002 (N_3002,N_2996,N_2916);
nor U3003 (N_3003,N_2905,N_2970);
nor U3004 (N_3004,N_2966,N_2955);
nand U3005 (N_3005,N_2975,N_2980);
and U3006 (N_3006,N_2973,N_2946);
nor U3007 (N_3007,N_2992,N_2998);
nand U3008 (N_3008,N_2910,N_2974);
nor U3009 (N_3009,N_2991,N_2927);
or U3010 (N_3010,N_2987,N_2887);
or U3011 (N_3011,N_2969,N_2986);
xor U3012 (N_3012,N_2961,N_2945);
and U3013 (N_3013,N_2957,N_2904);
xnor U3014 (N_3014,N_2911,N_2925);
or U3015 (N_3015,N_2940,N_2994);
xnor U3016 (N_3016,N_2939,N_2901);
nand U3017 (N_3017,N_2891,N_2875);
nor U3018 (N_3018,N_2968,N_2907);
or U3019 (N_3019,N_2963,N_2890);
nor U3020 (N_3020,N_2913,N_2922);
xnor U3021 (N_3021,N_2960,N_2964);
and U3022 (N_3022,N_2943,N_2976);
and U3023 (N_3023,N_2971,N_2944);
xnor U3024 (N_3024,N_2951,N_2886);
nand U3025 (N_3025,N_2878,N_2983);
or U3026 (N_3026,N_2898,N_2942);
nor U3027 (N_3027,N_2931,N_2936);
xor U3028 (N_3028,N_2906,N_2920);
xnor U3029 (N_3029,N_2934,N_2900);
nand U3030 (N_3030,N_2932,N_2972);
and U3031 (N_3031,N_2954,N_2885);
nor U3032 (N_3032,N_2930,N_2882);
nand U3033 (N_3033,N_2935,N_2877);
or U3034 (N_3034,N_2956,N_2921);
nand U3035 (N_3035,N_2929,N_2958);
nor U3036 (N_3036,N_2982,N_2953);
or U3037 (N_3037,N_2988,N_2962);
nor U3038 (N_3038,N_2924,N_2965);
nor U3039 (N_3039,N_2949,N_2879);
xor U3040 (N_3040,N_2908,N_2881);
nand U3041 (N_3041,N_2915,N_2948);
xnor U3042 (N_3042,N_2909,N_2993);
nand U3043 (N_3043,N_2959,N_2918);
and U3044 (N_3044,N_2893,N_2917);
or U3045 (N_3045,N_2926,N_2894);
or U3046 (N_3046,N_2895,N_2903);
nor U3047 (N_3047,N_2923,N_2884);
nand U3048 (N_3048,N_2977,N_2889);
or U3049 (N_3049,N_2888,N_2883);
or U3050 (N_3050,N_2952,N_2995);
or U3051 (N_3051,N_2880,N_2990);
nor U3052 (N_3052,N_2981,N_2933);
and U3053 (N_3053,N_2984,N_2912);
xor U3054 (N_3054,N_2979,N_2876);
and U3055 (N_3055,N_2999,N_2997);
or U3056 (N_3056,N_2947,N_2899);
nor U3057 (N_3057,N_2902,N_2941);
and U3058 (N_3058,N_2985,N_2914);
and U3059 (N_3059,N_2989,N_2950);
and U3060 (N_3060,N_2892,N_2919);
nor U3061 (N_3061,N_2938,N_2928);
nor U3062 (N_3062,N_2978,N_2936);
or U3063 (N_3063,N_2968,N_2996);
nand U3064 (N_3064,N_2976,N_2940);
or U3065 (N_3065,N_2890,N_2896);
or U3066 (N_3066,N_2878,N_2892);
or U3067 (N_3067,N_2919,N_2997);
xor U3068 (N_3068,N_2890,N_2956);
and U3069 (N_3069,N_2920,N_2954);
and U3070 (N_3070,N_2899,N_2982);
or U3071 (N_3071,N_2977,N_2944);
xnor U3072 (N_3072,N_2914,N_2931);
and U3073 (N_3073,N_2921,N_2948);
or U3074 (N_3074,N_2894,N_2941);
nand U3075 (N_3075,N_2956,N_2916);
nand U3076 (N_3076,N_2878,N_2885);
nor U3077 (N_3077,N_2939,N_2922);
and U3078 (N_3078,N_2909,N_2959);
or U3079 (N_3079,N_2906,N_2960);
xnor U3080 (N_3080,N_2931,N_2886);
nand U3081 (N_3081,N_2992,N_2906);
nand U3082 (N_3082,N_2906,N_2968);
and U3083 (N_3083,N_2910,N_2969);
nor U3084 (N_3084,N_2932,N_2878);
nand U3085 (N_3085,N_2939,N_2985);
or U3086 (N_3086,N_2894,N_2893);
xor U3087 (N_3087,N_2952,N_2944);
and U3088 (N_3088,N_2955,N_2968);
nor U3089 (N_3089,N_2909,N_2922);
and U3090 (N_3090,N_2926,N_2902);
nand U3091 (N_3091,N_2893,N_2999);
xor U3092 (N_3092,N_2978,N_2950);
xor U3093 (N_3093,N_2914,N_2898);
nor U3094 (N_3094,N_2919,N_2903);
or U3095 (N_3095,N_2885,N_2942);
xnor U3096 (N_3096,N_2906,N_2888);
or U3097 (N_3097,N_2930,N_2990);
xor U3098 (N_3098,N_2995,N_2965);
nor U3099 (N_3099,N_2905,N_2962);
and U3100 (N_3100,N_2960,N_2914);
nor U3101 (N_3101,N_2935,N_2895);
xor U3102 (N_3102,N_2932,N_2965);
or U3103 (N_3103,N_2988,N_2972);
xnor U3104 (N_3104,N_2937,N_2921);
nor U3105 (N_3105,N_2890,N_2969);
xnor U3106 (N_3106,N_2915,N_2962);
nor U3107 (N_3107,N_2895,N_2906);
nor U3108 (N_3108,N_2883,N_2991);
xor U3109 (N_3109,N_2992,N_2913);
xnor U3110 (N_3110,N_2965,N_2997);
nor U3111 (N_3111,N_2943,N_2898);
nand U3112 (N_3112,N_2885,N_2983);
or U3113 (N_3113,N_2929,N_2947);
and U3114 (N_3114,N_2923,N_2966);
nand U3115 (N_3115,N_2902,N_2904);
nand U3116 (N_3116,N_2960,N_2928);
and U3117 (N_3117,N_2925,N_2975);
and U3118 (N_3118,N_2877,N_2882);
xor U3119 (N_3119,N_2977,N_2999);
or U3120 (N_3120,N_2880,N_2903);
or U3121 (N_3121,N_2946,N_2894);
nand U3122 (N_3122,N_2908,N_2909);
nor U3123 (N_3123,N_2971,N_2892);
nor U3124 (N_3124,N_2989,N_2947);
and U3125 (N_3125,N_3124,N_3098);
nand U3126 (N_3126,N_3035,N_3063);
nor U3127 (N_3127,N_3105,N_3122);
and U3128 (N_3128,N_3000,N_3022);
xor U3129 (N_3129,N_3032,N_3060);
xor U3130 (N_3130,N_3059,N_3068);
nand U3131 (N_3131,N_3062,N_3077);
and U3132 (N_3132,N_3116,N_3016);
nor U3133 (N_3133,N_3054,N_3018);
or U3134 (N_3134,N_3101,N_3027);
nand U3135 (N_3135,N_3048,N_3046);
and U3136 (N_3136,N_3031,N_3041);
nor U3137 (N_3137,N_3121,N_3084);
and U3138 (N_3138,N_3023,N_3110);
nor U3139 (N_3139,N_3029,N_3038);
or U3140 (N_3140,N_3004,N_3028);
nor U3141 (N_3141,N_3024,N_3106);
xor U3142 (N_3142,N_3092,N_3025);
and U3143 (N_3143,N_3117,N_3011);
nand U3144 (N_3144,N_3019,N_3045);
xor U3145 (N_3145,N_3070,N_3073);
nand U3146 (N_3146,N_3093,N_3043);
and U3147 (N_3147,N_3079,N_3067);
and U3148 (N_3148,N_3088,N_3109);
and U3149 (N_3149,N_3107,N_3065);
nand U3150 (N_3150,N_3118,N_3072);
nand U3151 (N_3151,N_3040,N_3015);
xnor U3152 (N_3152,N_3007,N_3050);
or U3153 (N_3153,N_3100,N_3087);
or U3154 (N_3154,N_3086,N_3010);
nor U3155 (N_3155,N_3108,N_3044);
nor U3156 (N_3156,N_3094,N_3009);
and U3157 (N_3157,N_3013,N_3006);
or U3158 (N_3158,N_3052,N_3089);
and U3159 (N_3159,N_3069,N_3026);
and U3160 (N_3160,N_3014,N_3111);
nor U3161 (N_3161,N_3114,N_3104);
nor U3162 (N_3162,N_3064,N_3057);
nor U3163 (N_3163,N_3036,N_3058);
or U3164 (N_3164,N_3123,N_3039);
nand U3165 (N_3165,N_3055,N_3001);
xnor U3166 (N_3166,N_3034,N_3037);
or U3167 (N_3167,N_3103,N_3112);
or U3168 (N_3168,N_3071,N_3080);
nor U3169 (N_3169,N_3113,N_3049);
xor U3170 (N_3170,N_3119,N_3090);
nand U3171 (N_3171,N_3091,N_3081);
and U3172 (N_3172,N_3042,N_3033);
nand U3173 (N_3173,N_3115,N_3099);
xor U3174 (N_3174,N_3012,N_3020);
nor U3175 (N_3175,N_3061,N_3047);
xor U3176 (N_3176,N_3075,N_3076);
or U3177 (N_3177,N_3017,N_3120);
nor U3178 (N_3178,N_3066,N_3095);
nand U3179 (N_3179,N_3082,N_3008);
nand U3180 (N_3180,N_3030,N_3097);
or U3181 (N_3181,N_3083,N_3078);
xnor U3182 (N_3182,N_3074,N_3053);
nor U3183 (N_3183,N_3096,N_3002);
xnor U3184 (N_3184,N_3021,N_3003);
and U3185 (N_3185,N_3056,N_3005);
nand U3186 (N_3186,N_3085,N_3051);
xor U3187 (N_3187,N_3102,N_3043);
xnor U3188 (N_3188,N_3078,N_3117);
nand U3189 (N_3189,N_3087,N_3084);
or U3190 (N_3190,N_3053,N_3005);
xnor U3191 (N_3191,N_3115,N_3029);
or U3192 (N_3192,N_3011,N_3105);
and U3193 (N_3193,N_3025,N_3107);
and U3194 (N_3194,N_3105,N_3038);
nand U3195 (N_3195,N_3048,N_3011);
xnor U3196 (N_3196,N_3055,N_3016);
or U3197 (N_3197,N_3062,N_3061);
nand U3198 (N_3198,N_3055,N_3112);
and U3199 (N_3199,N_3087,N_3067);
or U3200 (N_3200,N_3020,N_3037);
nand U3201 (N_3201,N_3057,N_3059);
nand U3202 (N_3202,N_3018,N_3006);
xor U3203 (N_3203,N_3086,N_3124);
or U3204 (N_3204,N_3110,N_3005);
nor U3205 (N_3205,N_3041,N_3042);
nand U3206 (N_3206,N_3099,N_3088);
xnor U3207 (N_3207,N_3091,N_3099);
nand U3208 (N_3208,N_3092,N_3037);
or U3209 (N_3209,N_3101,N_3099);
nand U3210 (N_3210,N_3116,N_3047);
nor U3211 (N_3211,N_3073,N_3002);
and U3212 (N_3212,N_3008,N_3002);
xor U3213 (N_3213,N_3064,N_3049);
xor U3214 (N_3214,N_3002,N_3042);
or U3215 (N_3215,N_3119,N_3080);
nor U3216 (N_3216,N_3043,N_3029);
xor U3217 (N_3217,N_3037,N_3059);
xnor U3218 (N_3218,N_3117,N_3038);
nand U3219 (N_3219,N_3030,N_3057);
xor U3220 (N_3220,N_3049,N_3098);
nand U3221 (N_3221,N_3087,N_3058);
nor U3222 (N_3222,N_3002,N_3068);
nor U3223 (N_3223,N_3115,N_3065);
nand U3224 (N_3224,N_3015,N_3006);
nand U3225 (N_3225,N_3013,N_3074);
nand U3226 (N_3226,N_3039,N_3103);
nor U3227 (N_3227,N_3108,N_3115);
xor U3228 (N_3228,N_3005,N_3003);
nor U3229 (N_3229,N_3120,N_3106);
xnor U3230 (N_3230,N_3113,N_3098);
nand U3231 (N_3231,N_3074,N_3102);
nor U3232 (N_3232,N_3038,N_3101);
and U3233 (N_3233,N_3026,N_3064);
xor U3234 (N_3234,N_3009,N_3108);
nand U3235 (N_3235,N_3109,N_3113);
xor U3236 (N_3236,N_3061,N_3112);
nand U3237 (N_3237,N_3068,N_3017);
xor U3238 (N_3238,N_3104,N_3022);
xor U3239 (N_3239,N_3015,N_3078);
nor U3240 (N_3240,N_3050,N_3091);
xor U3241 (N_3241,N_3018,N_3085);
and U3242 (N_3242,N_3054,N_3122);
xnor U3243 (N_3243,N_3122,N_3117);
and U3244 (N_3244,N_3120,N_3124);
and U3245 (N_3245,N_3051,N_3056);
and U3246 (N_3246,N_3116,N_3004);
or U3247 (N_3247,N_3090,N_3102);
and U3248 (N_3248,N_3030,N_3041);
nand U3249 (N_3249,N_3015,N_3124);
xnor U3250 (N_3250,N_3129,N_3133);
nand U3251 (N_3251,N_3126,N_3213);
nor U3252 (N_3252,N_3236,N_3138);
and U3253 (N_3253,N_3243,N_3151);
and U3254 (N_3254,N_3128,N_3167);
xor U3255 (N_3255,N_3217,N_3234);
nand U3256 (N_3256,N_3184,N_3153);
or U3257 (N_3257,N_3211,N_3249);
nor U3258 (N_3258,N_3207,N_3210);
and U3259 (N_3259,N_3162,N_3175);
nor U3260 (N_3260,N_3161,N_3187);
xnor U3261 (N_3261,N_3208,N_3144);
or U3262 (N_3262,N_3188,N_3224);
xor U3263 (N_3263,N_3170,N_3156);
nand U3264 (N_3264,N_3185,N_3125);
xnor U3265 (N_3265,N_3163,N_3235);
nor U3266 (N_3266,N_3172,N_3171);
or U3267 (N_3267,N_3131,N_3215);
xor U3268 (N_3268,N_3149,N_3202);
nand U3269 (N_3269,N_3179,N_3242);
xnor U3270 (N_3270,N_3159,N_3228);
xor U3271 (N_3271,N_3189,N_3248);
xnor U3272 (N_3272,N_3160,N_3180);
or U3273 (N_3273,N_3177,N_3127);
and U3274 (N_3274,N_3196,N_3199);
nand U3275 (N_3275,N_3216,N_3173);
nand U3276 (N_3276,N_3176,N_3193);
and U3277 (N_3277,N_3247,N_3169);
and U3278 (N_3278,N_3142,N_3147);
or U3279 (N_3279,N_3137,N_3132);
nor U3280 (N_3280,N_3139,N_3214);
nor U3281 (N_3281,N_3182,N_3154);
nand U3282 (N_3282,N_3209,N_3135);
xor U3283 (N_3283,N_3158,N_3178);
nand U3284 (N_3284,N_3148,N_3227);
nand U3285 (N_3285,N_3230,N_3197);
and U3286 (N_3286,N_3246,N_3195);
nand U3287 (N_3287,N_3239,N_3223);
or U3288 (N_3288,N_3157,N_3231);
nand U3289 (N_3289,N_3130,N_3229);
nor U3290 (N_3290,N_3226,N_3198);
or U3291 (N_3291,N_3212,N_3241);
nand U3292 (N_3292,N_3221,N_3219);
or U3293 (N_3293,N_3174,N_3134);
and U3294 (N_3294,N_3136,N_3165);
nand U3295 (N_3295,N_3150,N_3205);
nand U3296 (N_3296,N_3181,N_3143);
nor U3297 (N_3297,N_3218,N_3200);
and U3298 (N_3298,N_3168,N_3203);
or U3299 (N_3299,N_3164,N_3194);
nand U3300 (N_3300,N_3140,N_3155);
nor U3301 (N_3301,N_3192,N_3146);
and U3302 (N_3302,N_3238,N_3225);
and U3303 (N_3303,N_3190,N_3240);
nor U3304 (N_3304,N_3166,N_3141);
xor U3305 (N_3305,N_3186,N_3201);
or U3306 (N_3306,N_3206,N_3191);
xor U3307 (N_3307,N_3232,N_3220);
xor U3308 (N_3308,N_3245,N_3152);
and U3309 (N_3309,N_3237,N_3204);
nand U3310 (N_3310,N_3233,N_3222);
nor U3311 (N_3311,N_3244,N_3183);
or U3312 (N_3312,N_3145,N_3214);
nand U3313 (N_3313,N_3238,N_3233);
and U3314 (N_3314,N_3204,N_3246);
or U3315 (N_3315,N_3248,N_3131);
xor U3316 (N_3316,N_3240,N_3236);
nor U3317 (N_3317,N_3212,N_3217);
or U3318 (N_3318,N_3178,N_3214);
nand U3319 (N_3319,N_3190,N_3180);
and U3320 (N_3320,N_3189,N_3243);
or U3321 (N_3321,N_3237,N_3244);
and U3322 (N_3322,N_3183,N_3179);
and U3323 (N_3323,N_3196,N_3217);
nand U3324 (N_3324,N_3171,N_3170);
xor U3325 (N_3325,N_3212,N_3216);
nor U3326 (N_3326,N_3129,N_3248);
nand U3327 (N_3327,N_3239,N_3192);
and U3328 (N_3328,N_3238,N_3152);
nor U3329 (N_3329,N_3151,N_3148);
nand U3330 (N_3330,N_3169,N_3151);
nand U3331 (N_3331,N_3227,N_3126);
nand U3332 (N_3332,N_3169,N_3239);
and U3333 (N_3333,N_3231,N_3196);
or U3334 (N_3334,N_3136,N_3239);
and U3335 (N_3335,N_3249,N_3128);
nor U3336 (N_3336,N_3190,N_3126);
nor U3337 (N_3337,N_3202,N_3140);
nor U3338 (N_3338,N_3187,N_3225);
nand U3339 (N_3339,N_3202,N_3173);
and U3340 (N_3340,N_3218,N_3189);
nor U3341 (N_3341,N_3191,N_3132);
nor U3342 (N_3342,N_3236,N_3221);
or U3343 (N_3343,N_3132,N_3243);
nand U3344 (N_3344,N_3154,N_3235);
xnor U3345 (N_3345,N_3228,N_3182);
nor U3346 (N_3346,N_3136,N_3142);
nand U3347 (N_3347,N_3221,N_3145);
nand U3348 (N_3348,N_3166,N_3150);
xor U3349 (N_3349,N_3242,N_3228);
xnor U3350 (N_3350,N_3224,N_3237);
nor U3351 (N_3351,N_3173,N_3215);
nand U3352 (N_3352,N_3220,N_3226);
nor U3353 (N_3353,N_3200,N_3246);
nor U3354 (N_3354,N_3202,N_3143);
nand U3355 (N_3355,N_3232,N_3142);
and U3356 (N_3356,N_3171,N_3140);
and U3357 (N_3357,N_3245,N_3222);
and U3358 (N_3358,N_3158,N_3169);
xnor U3359 (N_3359,N_3174,N_3166);
nor U3360 (N_3360,N_3193,N_3172);
and U3361 (N_3361,N_3170,N_3209);
or U3362 (N_3362,N_3230,N_3231);
xor U3363 (N_3363,N_3168,N_3164);
nor U3364 (N_3364,N_3248,N_3228);
or U3365 (N_3365,N_3164,N_3132);
xnor U3366 (N_3366,N_3227,N_3186);
or U3367 (N_3367,N_3186,N_3194);
and U3368 (N_3368,N_3172,N_3154);
nand U3369 (N_3369,N_3178,N_3189);
nand U3370 (N_3370,N_3185,N_3134);
xnor U3371 (N_3371,N_3188,N_3139);
or U3372 (N_3372,N_3241,N_3192);
and U3373 (N_3373,N_3146,N_3144);
xor U3374 (N_3374,N_3136,N_3235);
nand U3375 (N_3375,N_3324,N_3340);
nor U3376 (N_3376,N_3270,N_3320);
and U3377 (N_3377,N_3288,N_3346);
nor U3378 (N_3378,N_3341,N_3256);
nor U3379 (N_3379,N_3331,N_3300);
and U3380 (N_3380,N_3333,N_3301);
or U3381 (N_3381,N_3286,N_3322);
or U3382 (N_3382,N_3257,N_3302);
nor U3383 (N_3383,N_3303,N_3362);
nor U3384 (N_3384,N_3345,N_3293);
nand U3385 (N_3385,N_3268,N_3364);
nor U3386 (N_3386,N_3327,N_3369);
nor U3387 (N_3387,N_3285,N_3321);
and U3388 (N_3388,N_3307,N_3330);
and U3389 (N_3389,N_3308,N_3306);
xor U3390 (N_3390,N_3342,N_3292);
xnor U3391 (N_3391,N_3304,N_3277);
nand U3392 (N_3392,N_3252,N_3356);
or U3393 (N_3393,N_3314,N_3373);
or U3394 (N_3394,N_3262,N_3311);
nand U3395 (N_3395,N_3354,N_3275);
nand U3396 (N_3396,N_3317,N_3253);
xor U3397 (N_3397,N_3371,N_3325);
or U3398 (N_3398,N_3335,N_3296);
or U3399 (N_3399,N_3374,N_3282);
or U3400 (N_3400,N_3310,N_3348);
and U3401 (N_3401,N_3276,N_3336);
and U3402 (N_3402,N_3360,N_3349);
xnor U3403 (N_3403,N_3250,N_3290);
nand U3404 (N_3404,N_3326,N_3294);
or U3405 (N_3405,N_3339,N_3297);
nand U3406 (N_3406,N_3357,N_3278);
nor U3407 (N_3407,N_3267,N_3359);
nand U3408 (N_3408,N_3363,N_3284);
and U3409 (N_3409,N_3316,N_3351);
and U3410 (N_3410,N_3274,N_3312);
nor U3411 (N_3411,N_3319,N_3273);
and U3412 (N_3412,N_3298,N_3370);
and U3413 (N_3413,N_3280,N_3313);
or U3414 (N_3414,N_3259,N_3344);
xor U3415 (N_3415,N_3329,N_3338);
nor U3416 (N_3416,N_3366,N_3255);
nor U3417 (N_3417,N_3368,N_3372);
nand U3418 (N_3418,N_3365,N_3283);
nand U3419 (N_3419,N_3251,N_3361);
xnor U3420 (N_3420,N_3309,N_3350);
or U3421 (N_3421,N_3355,N_3343);
nand U3422 (N_3422,N_3295,N_3334);
nand U3423 (N_3423,N_3263,N_3279);
nand U3424 (N_3424,N_3323,N_3260);
xnor U3425 (N_3425,N_3367,N_3299);
nand U3426 (N_3426,N_3261,N_3358);
xnor U3427 (N_3427,N_3347,N_3353);
nor U3428 (N_3428,N_3289,N_3315);
nand U3429 (N_3429,N_3254,N_3264);
nand U3430 (N_3430,N_3269,N_3287);
xor U3431 (N_3431,N_3305,N_3265);
nand U3432 (N_3432,N_3281,N_3266);
xnor U3433 (N_3433,N_3258,N_3328);
xnor U3434 (N_3434,N_3332,N_3352);
xnor U3435 (N_3435,N_3291,N_3271);
nand U3436 (N_3436,N_3337,N_3272);
nor U3437 (N_3437,N_3318,N_3368);
and U3438 (N_3438,N_3369,N_3356);
nand U3439 (N_3439,N_3339,N_3255);
nand U3440 (N_3440,N_3271,N_3340);
nand U3441 (N_3441,N_3310,N_3251);
nand U3442 (N_3442,N_3289,N_3363);
and U3443 (N_3443,N_3360,N_3337);
nand U3444 (N_3444,N_3268,N_3262);
or U3445 (N_3445,N_3254,N_3335);
or U3446 (N_3446,N_3305,N_3278);
nand U3447 (N_3447,N_3263,N_3283);
or U3448 (N_3448,N_3357,N_3365);
nor U3449 (N_3449,N_3305,N_3318);
nor U3450 (N_3450,N_3343,N_3348);
and U3451 (N_3451,N_3335,N_3342);
xnor U3452 (N_3452,N_3366,N_3325);
nor U3453 (N_3453,N_3315,N_3356);
and U3454 (N_3454,N_3373,N_3324);
and U3455 (N_3455,N_3348,N_3295);
nand U3456 (N_3456,N_3300,N_3255);
nand U3457 (N_3457,N_3275,N_3260);
and U3458 (N_3458,N_3263,N_3293);
xnor U3459 (N_3459,N_3267,N_3284);
and U3460 (N_3460,N_3325,N_3322);
nand U3461 (N_3461,N_3351,N_3251);
and U3462 (N_3462,N_3292,N_3269);
and U3463 (N_3463,N_3266,N_3314);
or U3464 (N_3464,N_3325,N_3305);
xor U3465 (N_3465,N_3324,N_3261);
xor U3466 (N_3466,N_3303,N_3319);
nor U3467 (N_3467,N_3307,N_3327);
nand U3468 (N_3468,N_3356,N_3307);
nand U3469 (N_3469,N_3333,N_3277);
nand U3470 (N_3470,N_3307,N_3346);
or U3471 (N_3471,N_3370,N_3316);
nor U3472 (N_3472,N_3266,N_3260);
nor U3473 (N_3473,N_3347,N_3325);
xor U3474 (N_3474,N_3318,N_3369);
xnor U3475 (N_3475,N_3258,N_3297);
nand U3476 (N_3476,N_3307,N_3313);
and U3477 (N_3477,N_3282,N_3262);
or U3478 (N_3478,N_3290,N_3368);
nor U3479 (N_3479,N_3265,N_3347);
and U3480 (N_3480,N_3303,N_3280);
xnor U3481 (N_3481,N_3317,N_3323);
xor U3482 (N_3482,N_3319,N_3311);
or U3483 (N_3483,N_3340,N_3365);
and U3484 (N_3484,N_3335,N_3340);
nor U3485 (N_3485,N_3281,N_3283);
and U3486 (N_3486,N_3294,N_3338);
or U3487 (N_3487,N_3289,N_3307);
nand U3488 (N_3488,N_3326,N_3368);
nor U3489 (N_3489,N_3330,N_3298);
nand U3490 (N_3490,N_3253,N_3359);
xnor U3491 (N_3491,N_3321,N_3373);
or U3492 (N_3492,N_3338,N_3266);
and U3493 (N_3493,N_3323,N_3360);
and U3494 (N_3494,N_3374,N_3330);
nand U3495 (N_3495,N_3348,N_3340);
and U3496 (N_3496,N_3274,N_3320);
xor U3497 (N_3497,N_3330,N_3327);
xor U3498 (N_3498,N_3320,N_3345);
or U3499 (N_3499,N_3346,N_3331);
and U3500 (N_3500,N_3394,N_3498);
nand U3501 (N_3501,N_3469,N_3455);
or U3502 (N_3502,N_3376,N_3380);
or U3503 (N_3503,N_3417,N_3485);
xor U3504 (N_3504,N_3412,N_3442);
nor U3505 (N_3505,N_3416,N_3441);
xor U3506 (N_3506,N_3486,N_3425);
and U3507 (N_3507,N_3472,N_3451);
and U3508 (N_3508,N_3483,N_3439);
xnor U3509 (N_3509,N_3436,N_3420);
and U3510 (N_3510,N_3383,N_3461);
xor U3511 (N_3511,N_3445,N_3488);
and U3512 (N_3512,N_3395,N_3410);
or U3513 (N_3513,N_3386,N_3422);
xnor U3514 (N_3514,N_3392,N_3473);
xnor U3515 (N_3515,N_3490,N_3443);
nand U3516 (N_3516,N_3377,N_3448);
xnor U3517 (N_3517,N_3415,N_3474);
nand U3518 (N_3518,N_3418,N_3444);
nand U3519 (N_3519,N_3431,N_3426);
xnor U3520 (N_3520,N_3482,N_3449);
nand U3521 (N_3521,N_3432,N_3494);
and U3522 (N_3522,N_3497,N_3495);
nand U3523 (N_3523,N_3384,N_3391);
xor U3524 (N_3524,N_3411,N_3385);
and U3525 (N_3525,N_3475,N_3471);
or U3526 (N_3526,N_3479,N_3493);
and U3527 (N_3527,N_3446,N_3492);
xor U3528 (N_3528,N_3453,N_3387);
nor U3529 (N_3529,N_3419,N_3382);
and U3530 (N_3530,N_3435,N_3489);
xor U3531 (N_3531,N_3459,N_3400);
and U3532 (N_3532,N_3454,N_3465);
nand U3533 (N_3533,N_3478,N_3399);
and U3534 (N_3534,N_3393,N_3379);
nand U3535 (N_3535,N_3460,N_3428);
nor U3536 (N_3536,N_3476,N_3450);
nor U3537 (N_3537,N_3466,N_3447);
or U3538 (N_3538,N_3407,N_3440);
xor U3539 (N_3539,N_3467,N_3408);
or U3540 (N_3540,N_3452,N_3381);
nor U3541 (N_3541,N_3405,N_3421);
xnor U3542 (N_3542,N_3403,N_3481);
xor U3543 (N_3543,N_3375,N_3430);
nand U3544 (N_3544,N_3429,N_3477);
nand U3545 (N_3545,N_3427,N_3433);
nand U3546 (N_3546,N_3468,N_3404);
or U3547 (N_3547,N_3491,N_3496);
or U3548 (N_3548,N_3458,N_3423);
nand U3549 (N_3549,N_3438,N_3402);
nand U3550 (N_3550,N_3414,N_3378);
or U3551 (N_3551,N_3457,N_3437);
nor U3552 (N_3552,N_3389,N_3464);
nor U3553 (N_3553,N_3434,N_3424);
and U3554 (N_3554,N_3409,N_3463);
or U3555 (N_3555,N_3487,N_3396);
nor U3556 (N_3556,N_3397,N_3398);
nor U3557 (N_3557,N_3390,N_3470);
nor U3558 (N_3558,N_3462,N_3480);
and U3559 (N_3559,N_3413,N_3406);
and U3560 (N_3560,N_3401,N_3499);
xor U3561 (N_3561,N_3456,N_3388);
xnor U3562 (N_3562,N_3484,N_3395);
xor U3563 (N_3563,N_3446,N_3397);
or U3564 (N_3564,N_3494,N_3477);
nand U3565 (N_3565,N_3438,N_3445);
nor U3566 (N_3566,N_3378,N_3496);
or U3567 (N_3567,N_3466,N_3375);
nand U3568 (N_3568,N_3386,N_3476);
nor U3569 (N_3569,N_3489,N_3411);
nand U3570 (N_3570,N_3492,N_3416);
xnor U3571 (N_3571,N_3432,N_3406);
and U3572 (N_3572,N_3458,N_3424);
nand U3573 (N_3573,N_3423,N_3433);
and U3574 (N_3574,N_3383,N_3391);
xor U3575 (N_3575,N_3481,N_3442);
nand U3576 (N_3576,N_3424,N_3473);
nand U3577 (N_3577,N_3409,N_3491);
nor U3578 (N_3578,N_3460,N_3468);
or U3579 (N_3579,N_3417,N_3397);
xor U3580 (N_3580,N_3388,N_3442);
xor U3581 (N_3581,N_3472,N_3379);
nor U3582 (N_3582,N_3436,N_3395);
and U3583 (N_3583,N_3377,N_3481);
xor U3584 (N_3584,N_3492,N_3412);
nor U3585 (N_3585,N_3405,N_3451);
xnor U3586 (N_3586,N_3385,N_3446);
or U3587 (N_3587,N_3477,N_3464);
or U3588 (N_3588,N_3486,N_3462);
and U3589 (N_3589,N_3389,N_3484);
nor U3590 (N_3590,N_3429,N_3441);
and U3591 (N_3591,N_3413,N_3424);
nand U3592 (N_3592,N_3446,N_3395);
nor U3593 (N_3593,N_3481,N_3379);
or U3594 (N_3594,N_3381,N_3392);
nor U3595 (N_3595,N_3475,N_3408);
or U3596 (N_3596,N_3476,N_3459);
nand U3597 (N_3597,N_3444,N_3464);
or U3598 (N_3598,N_3421,N_3414);
xnor U3599 (N_3599,N_3476,N_3432);
nor U3600 (N_3600,N_3494,N_3391);
xnor U3601 (N_3601,N_3497,N_3474);
xor U3602 (N_3602,N_3486,N_3438);
nor U3603 (N_3603,N_3466,N_3384);
nor U3604 (N_3604,N_3402,N_3457);
nor U3605 (N_3605,N_3431,N_3485);
nor U3606 (N_3606,N_3484,N_3474);
or U3607 (N_3607,N_3439,N_3404);
xnor U3608 (N_3608,N_3491,N_3458);
nand U3609 (N_3609,N_3430,N_3466);
xnor U3610 (N_3610,N_3479,N_3408);
xor U3611 (N_3611,N_3382,N_3418);
and U3612 (N_3612,N_3412,N_3417);
and U3613 (N_3613,N_3444,N_3462);
or U3614 (N_3614,N_3387,N_3441);
nor U3615 (N_3615,N_3483,N_3478);
or U3616 (N_3616,N_3453,N_3461);
and U3617 (N_3617,N_3379,N_3430);
and U3618 (N_3618,N_3495,N_3465);
xnor U3619 (N_3619,N_3485,N_3453);
or U3620 (N_3620,N_3490,N_3385);
nand U3621 (N_3621,N_3436,N_3381);
xor U3622 (N_3622,N_3375,N_3438);
nand U3623 (N_3623,N_3402,N_3455);
nor U3624 (N_3624,N_3421,N_3492);
nor U3625 (N_3625,N_3583,N_3506);
or U3626 (N_3626,N_3561,N_3551);
nand U3627 (N_3627,N_3597,N_3622);
nor U3628 (N_3628,N_3563,N_3511);
and U3629 (N_3629,N_3607,N_3560);
xor U3630 (N_3630,N_3567,N_3547);
nand U3631 (N_3631,N_3591,N_3600);
and U3632 (N_3632,N_3574,N_3535);
and U3633 (N_3633,N_3604,N_3608);
nor U3634 (N_3634,N_3504,N_3501);
or U3635 (N_3635,N_3584,N_3508);
nand U3636 (N_3636,N_3530,N_3503);
or U3637 (N_3637,N_3569,N_3543);
nor U3638 (N_3638,N_3568,N_3595);
nand U3639 (N_3639,N_3515,N_3610);
nor U3640 (N_3640,N_3575,N_3572);
xor U3641 (N_3641,N_3510,N_3605);
and U3642 (N_3642,N_3520,N_3564);
and U3643 (N_3643,N_3514,N_3556);
nor U3644 (N_3644,N_3581,N_3621);
nand U3645 (N_3645,N_3537,N_3549);
nand U3646 (N_3646,N_3599,N_3500);
and U3647 (N_3647,N_3623,N_3580);
nand U3648 (N_3648,N_3523,N_3519);
and U3649 (N_3649,N_3539,N_3619);
nor U3650 (N_3650,N_3518,N_3606);
nor U3651 (N_3651,N_3544,N_3562);
or U3652 (N_3652,N_3579,N_3602);
xnor U3653 (N_3653,N_3578,N_3546);
and U3654 (N_3654,N_3582,N_3557);
xnor U3655 (N_3655,N_3612,N_3577);
or U3656 (N_3656,N_3538,N_3534);
or U3657 (N_3657,N_3529,N_3573);
xnor U3658 (N_3658,N_3541,N_3553);
xnor U3659 (N_3659,N_3526,N_3528);
nand U3660 (N_3660,N_3588,N_3586);
nor U3661 (N_3661,N_3509,N_3540);
and U3662 (N_3662,N_3590,N_3616);
xor U3663 (N_3663,N_3502,N_3542);
nand U3664 (N_3664,N_3613,N_3611);
nor U3665 (N_3665,N_3589,N_3524);
nor U3666 (N_3666,N_3614,N_3532);
nor U3667 (N_3667,N_3603,N_3565);
nand U3668 (N_3668,N_3555,N_3513);
and U3669 (N_3669,N_3571,N_3527);
and U3670 (N_3670,N_3609,N_3536);
and U3671 (N_3671,N_3516,N_3620);
and U3672 (N_3672,N_3552,N_3566);
or U3673 (N_3673,N_3585,N_3521);
and U3674 (N_3674,N_3505,N_3517);
or U3675 (N_3675,N_3576,N_3531);
and U3676 (N_3676,N_3548,N_3615);
xnor U3677 (N_3677,N_3587,N_3558);
nand U3678 (N_3678,N_3594,N_3512);
nor U3679 (N_3679,N_3593,N_3525);
and U3680 (N_3680,N_3545,N_3559);
nor U3681 (N_3681,N_3618,N_3598);
and U3682 (N_3682,N_3570,N_3592);
or U3683 (N_3683,N_3550,N_3533);
and U3684 (N_3684,N_3596,N_3601);
xnor U3685 (N_3685,N_3554,N_3507);
and U3686 (N_3686,N_3624,N_3522);
xnor U3687 (N_3687,N_3617,N_3582);
xor U3688 (N_3688,N_3591,N_3579);
nand U3689 (N_3689,N_3578,N_3601);
xnor U3690 (N_3690,N_3525,N_3538);
xor U3691 (N_3691,N_3555,N_3623);
or U3692 (N_3692,N_3545,N_3604);
and U3693 (N_3693,N_3582,N_3598);
nand U3694 (N_3694,N_3594,N_3522);
and U3695 (N_3695,N_3538,N_3510);
nand U3696 (N_3696,N_3505,N_3580);
xnor U3697 (N_3697,N_3509,N_3581);
xor U3698 (N_3698,N_3622,N_3596);
nand U3699 (N_3699,N_3563,N_3621);
xor U3700 (N_3700,N_3581,N_3602);
nand U3701 (N_3701,N_3577,N_3531);
and U3702 (N_3702,N_3562,N_3507);
nand U3703 (N_3703,N_3569,N_3546);
xnor U3704 (N_3704,N_3599,N_3519);
xor U3705 (N_3705,N_3579,N_3571);
xor U3706 (N_3706,N_3536,N_3551);
nor U3707 (N_3707,N_3569,N_3587);
and U3708 (N_3708,N_3593,N_3622);
or U3709 (N_3709,N_3580,N_3568);
xnor U3710 (N_3710,N_3609,N_3567);
nand U3711 (N_3711,N_3586,N_3568);
or U3712 (N_3712,N_3597,N_3572);
nand U3713 (N_3713,N_3580,N_3565);
nor U3714 (N_3714,N_3547,N_3539);
nand U3715 (N_3715,N_3594,N_3546);
and U3716 (N_3716,N_3563,N_3512);
and U3717 (N_3717,N_3612,N_3528);
nand U3718 (N_3718,N_3578,N_3528);
nor U3719 (N_3719,N_3509,N_3541);
xor U3720 (N_3720,N_3555,N_3514);
nand U3721 (N_3721,N_3500,N_3532);
nand U3722 (N_3722,N_3550,N_3554);
and U3723 (N_3723,N_3545,N_3565);
and U3724 (N_3724,N_3508,N_3510);
nor U3725 (N_3725,N_3556,N_3586);
xor U3726 (N_3726,N_3505,N_3613);
or U3727 (N_3727,N_3549,N_3571);
nand U3728 (N_3728,N_3500,N_3521);
or U3729 (N_3729,N_3575,N_3537);
or U3730 (N_3730,N_3552,N_3520);
xnor U3731 (N_3731,N_3608,N_3592);
and U3732 (N_3732,N_3565,N_3590);
and U3733 (N_3733,N_3582,N_3610);
nor U3734 (N_3734,N_3579,N_3583);
xor U3735 (N_3735,N_3604,N_3528);
xnor U3736 (N_3736,N_3565,N_3510);
nor U3737 (N_3737,N_3603,N_3623);
nand U3738 (N_3738,N_3505,N_3522);
nor U3739 (N_3739,N_3603,N_3518);
xor U3740 (N_3740,N_3587,N_3602);
xnor U3741 (N_3741,N_3521,N_3505);
and U3742 (N_3742,N_3587,N_3592);
nor U3743 (N_3743,N_3503,N_3522);
nand U3744 (N_3744,N_3559,N_3512);
xnor U3745 (N_3745,N_3579,N_3586);
nand U3746 (N_3746,N_3554,N_3541);
xor U3747 (N_3747,N_3545,N_3587);
nand U3748 (N_3748,N_3512,N_3589);
and U3749 (N_3749,N_3591,N_3577);
or U3750 (N_3750,N_3643,N_3706);
or U3751 (N_3751,N_3727,N_3686);
xnor U3752 (N_3752,N_3729,N_3733);
and U3753 (N_3753,N_3672,N_3677);
nor U3754 (N_3754,N_3687,N_3693);
and U3755 (N_3755,N_3713,N_3639);
nand U3756 (N_3756,N_3707,N_3670);
nand U3757 (N_3757,N_3647,N_3736);
or U3758 (N_3758,N_3685,N_3722);
nand U3759 (N_3759,N_3701,N_3746);
xor U3760 (N_3760,N_3721,N_3696);
nor U3761 (N_3761,N_3705,N_3709);
xnor U3762 (N_3762,N_3719,N_3718);
or U3763 (N_3763,N_3649,N_3749);
and U3764 (N_3764,N_3630,N_3742);
or U3765 (N_3765,N_3726,N_3720);
nand U3766 (N_3766,N_3651,N_3744);
or U3767 (N_3767,N_3673,N_3631);
xnor U3768 (N_3768,N_3711,N_3741);
nand U3769 (N_3769,N_3626,N_3732);
xnor U3770 (N_3770,N_3661,N_3634);
nand U3771 (N_3771,N_3728,N_3699);
xnor U3772 (N_3772,N_3735,N_3641);
nand U3773 (N_3773,N_3655,N_3738);
and U3774 (N_3774,N_3676,N_3652);
or U3775 (N_3775,N_3723,N_3646);
xor U3776 (N_3776,N_3692,N_3659);
and U3777 (N_3777,N_3637,N_3635);
nand U3778 (N_3778,N_3645,N_3747);
nor U3779 (N_3779,N_3683,N_3665);
nor U3780 (N_3780,N_3714,N_3704);
or U3781 (N_3781,N_3737,N_3648);
nand U3782 (N_3782,N_3684,N_3667);
xor U3783 (N_3783,N_3724,N_3653);
nand U3784 (N_3784,N_3663,N_3679);
xor U3785 (N_3785,N_3725,N_3712);
or U3786 (N_3786,N_3627,N_3632);
xnor U3787 (N_3787,N_3700,N_3695);
and U3788 (N_3788,N_3710,N_3708);
nand U3789 (N_3789,N_3668,N_3702);
and U3790 (N_3790,N_3629,N_3681);
xor U3791 (N_3791,N_3654,N_3644);
nor U3792 (N_3792,N_3745,N_3682);
nor U3793 (N_3793,N_3656,N_3642);
nor U3794 (N_3794,N_3657,N_3666);
or U3795 (N_3795,N_3697,N_3640);
nor U3796 (N_3796,N_3636,N_3689);
nand U3797 (N_3797,N_3633,N_3715);
nor U3798 (N_3798,N_3628,N_3675);
or U3799 (N_3799,N_3688,N_3658);
xor U3800 (N_3800,N_3716,N_3734);
nand U3801 (N_3801,N_3739,N_3748);
and U3802 (N_3802,N_3669,N_3662);
nor U3803 (N_3803,N_3730,N_3743);
or U3804 (N_3804,N_3678,N_3694);
or U3805 (N_3805,N_3625,N_3650);
xnor U3806 (N_3806,N_3691,N_3703);
and U3807 (N_3807,N_3717,N_3638);
nand U3808 (N_3808,N_3660,N_3680);
or U3809 (N_3809,N_3731,N_3664);
nand U3810 (N_3810,N_3690,N_3740);
or U3811 (N_3811,N_3698,N_3671);
or U3812 (N_3812,N_3674,N_3646);
nand U3813 (N_3813,N_3735,N_3670);
or U3814 (N_3814,N_3716,N_3637);
nand U3815 (N_3815,N_3657,N_3676);
nor U3816 (N_3816,N_3674,N_3671);
xor U3817 (N_3817,N_3665,N_3641);
xor U3818 (N_3818,N_3722,N_3663);
and U3819 (N_3819,N_3632,N_3697);
xnor U3820 (N_3820,N_3748,N_3684);
or U3821 (N_3821,N_3743,N_3709);
xnor U3822 (N_3822,N_3665,N_3707);
xor U3823 (N_3823,N_3705,N_3671);
nand U3824 (N_3824,N_3702,N_3675);
nor U3825 (N_3825,N_3674,N_3726);
xnor U3826 (N_3826,N_3648,N_3678);
nand U3827 (N_3827,N_3636,N_3700);
xor U3828 (N_3828,N_3667,N_3714);
xnor U3829 (N_3829,N_3688,N_3698);
and U3830 (N_3830,N_3699,N_3725);
nand U3831 (N_3831,N_3701,N_3637);
or U3832 (N_3832,N_3665,N_3715);
and U3833 (N_3833,N_3693,N_3683);
nand U3834 (N_3834,N_3683,N_3748);
nand U3835 (N_3835,N_3689,N_3670);
nand U3836 (N_3836,N_3743,N_3630);
xnor U3837 (N_3837,N_3648,N_3652);
nor U3838 (N_3838,N_3651,N_3641);
nand U3839 (N_3839,N_3633,N_3709);
and U3840 (N_3840,N_3722,N_3702);
xor U3841 (N_3841,N_3658,N_3711);
or U3842 (N_3842,N_3688,N_3692);
nor U3843 (N_3843,N_3698,N_3646);
nand U3844 (N_3844,N_3707,N_3741);
nor U3845 (N_3845,N_3702,N_3662);
nand U3846 (N_3846,N_3745,N_3633);
nand U3847 (N_3847,N_3700,N_3714);
and U3848 (N_3848,N_3678,N_3687);
xnor U3849 (N_3849,N_3696,N_3668);
nor U3850 (N_3850,N_3740,N_3706);
and U3851 (N_3851,N_3741,N_3659);
and U3852 (N_3852,N_3689,N_3650);
and U3853 (N_3853,N_3749,N_3641);
nand U3854 (N_3854,N_3736,N_3718);
nor U3855 (N_3855,N_3636,N_3718);
or U3856 (N_3856,N_3682,N_3698);
nor U3857 (N_3857,N_3686,N_3692);
and U3858 (N_3858,N_3634,N_3723);
or U3859 (N_3859,N_3727,N_3684);
nor U3860 (N_3860,N_3703,N_3732);
xnor U3861 (N_3861,N_3735,N_3697);
nand U3862 (N_3862,N_3638,N_3749);
nand U3863 (N_3863,N_3642,N_3677);
xnor U3864 (N_3864,N_3688,N_3720);
or U3865 (N_3865,N_3668,N_3739);
nor U3866 (N_3866,N_3663,N_3731);
xnor U3867 (N_3867,N_3710,N_3735);
nor U3868 (N_3868,N_3734,N_3640);
or U3869 (N_3869,N_3639,N_3651);
and U3870 (N_3870,N_3665,N_3690);
and U3871 (N_3871,N_3693,N_3701);
nand U3872 (N_3872,N_3659,N_3672);
nor U3873 (N_3873,N_3739,N_3629);
or U3874 (N_3874,N_3629,N_3666);
nor U3875 (N_3875,N_3867,N_3817);
xnor U3876 (N_3876,N_3862,N_3812);
and U3877 (N_3877,N_3821,N_3796);
nor U3878 (N_3878,N_3848,N_3835);
or U3879 (N_3879,N_3792,N_3807);
xnor U3880 (N_3880,N_3778,N_3776);
nor U3881 (N_3881,N_3836,N_3840);
and U3882 (N_3882,N_3762,N_3760);
nor U3883 (N_3883,N_3847,N_3874);
nand U3884 (N_3884,N_3756,N_3753);
nor U3885 (N_3885,N_3841,N_3786);
nand U3886 (N_3886,N_3782,N_3795);
nand U3887 (N_3887,N_3868,N_3755);
and U3888 (N_3888,N_3811,N_3774);
or U3889 (N_3889,N_3818,N_3783);
or U3890 (N_3890,N_3813,N_3777);
xor U3891 (N_3891,N_3788,N_3846);
and U3892 (N_3892,N_3838,N_3844);
nor U3893 (N_3893,N_3842,N_3827);
and U3894 (N_3894,N_3856,N_3767);
nor U3895 (N_3895,N_3804,N_3750);
and U3896 (N_3896,N_3873,N_3759);
and U3897 (N_3897,N_3771,N_3787);
nor U3898 (N_3898,N_3772,N_3822);
nor U3899 (N_3899,N_3843,N_3852);
nor U3900 (N_3900,N_3785,N_3870);
and U3901 (N_3901,N_3823,N_3851);
or U3902 (N_3902,N_3810,N_3808);
nand U3903 (N_3903,N_3806,N_3864);
and U3904 (N_3904,N_3849,N_3820);
nor U3905 (N_3905,N_3773,N_3809);
nor U3906 (N_3906,N_3832,N_3829);
nand U3907 (N_3907,N_3850,N_3859);
xnor U3908 (N_3908,N_3830,N_3805);
xnor U3909 (N_3909,N_3791,N_3781);
nor U3910 (N_3910,N_3831,N_3765);
nand U3911 (N_3911,N_3793,N_3866);
or U3912 (N_3912,N_3869,N_3789);
or U3913 (N_3913,N_3861,N_3854);
nor U3914 (N_3914,N_3815,N_3824);
nor U3915 (N_3915,N_3761,N_3872);
xnor U3916 (N_3916,N_3799,N_3775);
nor U3917 (N_3917,N_3770,N_3803);
nand U3918 (N_3918,N_3816,N_3751);
and U3919 (N_3919,N_3794,N_3828);
xor U3920 (N_3920,N_3754,N_3860);
nand U3921 (N_3921,N_3865,N_3752);
nor U3922 (N_3922,N_3801,N_3845);
xnor U3923 (N_3923,N_3784,N_3764);
or U3924 (N_3924,N_3855,N_3758);
nand U3925 (N_3925,N_3863,N_3819);
nand U3926 (N_3926,N_3853,N_3797);
or U3927 (N_3927,N_3834,N_3798);
and U3928 (N_3928,N_3790,N_3779);
xnor U3929 (N_3929,N_3768,N_3800);
and U3930 (N_3930,N_3802,N_3763);
and U3931 (N_3931,N_3766,N_3833);
or U3932 (N_3932,N_3780,N_3769);
and U3933 (N_3933,N_3837,N_3826);
nor U3934 (N_3934,N_3757,N_3871);
xnor U3935 (N_3935,N_3814,N_3839);
nor U3936 (N_3936,N_3857,N_3825);
nor U3937 (N_3937,N_3858,N_3857);
nand U3938 (N_3938,N_3847,N_3795);
or U3939 (N_3939,N_3780,N_3776);
and U3940 (N_3940,N_3828,N_3865);
nor U3941 (N_3941,N_3808,N_3768);
xnor U3942 (N_3942,N_3847,N_3818);
and U3943 (N_3943,N_3826,N_3821);
or U3944 (N_3944,N_3768,N_3816);
nor U3945 (N_3945,N_3857,N_3819);
nand U3946 (N_3946,N_3843,N_3815);
or U3947 (N_3947,N_3815,N_3755);
or U3948 (N_3948,N_3763,N_3865);
nor U3949 (N_3949,N_3861,N_3752);
or U3950 (N_3950,N_3790,N_3825);
xnor U3951 (N_3951,N_3818,N_3873);
nor U3952 (N_3952,N_3768,N_3829);
nand U3953 (N_3953,N_3759,N_3870);
nand U3954 (N_3954,N_3817,N_3803);
and U3955 (N_3955,N_3841,N_3771);
nand U3956 (N_3956,N_3758,N_3763);
nor U3957 (N_3957,N_3793,N_3794);
nand U3958 (N_3958,N_3763,N_3797);
nand U3959 (N_3959,N_3760,N_3787);
xnor U3960 (N_3960,N_3867,N_3826);
nor U3961 (N_3961,N_3772,N_3798);
or U3962 (N_3962,N_3792,N_3766);
xnor U3963 (N_3963,N_3767,N_3802);
and U3964 (N_3964,N_3818,N_3817);
and U3965 (N_3965,N_3832,N_3873);
xnor U3966 (N_3966,N_3864,N_3854);
nor U3967 (N_3967,N_3791,N_3816);
and U3968 (N_3968,N_3767,N_3791);
xor U3969 (N_3969,N_3871,N_3760);
or U3970 (N_3970,N_3828,N_3753);
nor U3971 (N_3971,N_3810,N_3799);
or U3972 (N_3972,N_3843,N_3854);
and U3973 (N_3973,N_3833,N_3866);
nand U3974 (N_3974,N_3838,N_3823);
xor U3975 (N_3975,N_3829,N_3837);
xnor U3976 (N_3976,N_3783,N_3780);
or U3977 (N_3977,N_3802,N_3852);
nand U3978 (N_3978,N_3851,N_3806);
nor U3979 (N_3979,N_3767,N_3826);
xnor U3980 (N_3980,N_3757,N_3829);
or U3981 (N_3981,N_3866,N_3803);
or U3982 (N_3982,N_3758,N_3838);
nor U3983 (N_3983,N_3824,N_3869);
or U3984 (N_3984,N_3824,N_3868);
and U3985 (N_3985,N_3762,N_3761);
xnor U3986 (N_3986,N_3750,N_3815);
nor U3987 (N_3987,N_3851,N_3750);
nand U3988 (N_3988,N_3823,N_3762);
xor U3989 (N_3989,N_3771,N_3799);
and U3990 (N_3990,N_3817,N_3830);
or U3991 (N_3991,N_3810,N_3781);
or U3992 (N_3992,N_3795,N_3805);
nand U3993 (N_3993,N_3792,N_3819);
nand U3994 (N_3994,N_3872,N_3801);
xor U3995 (N_3995,N_3824,N_3784);
nor U3996 (N_3996,N_3797,N_3794);
xor U3997 (N_3997,N_3756,N_3845);
nand U3998 (N_3998,N_3769,N_3869);
nand U3999 (N_3999,N_3854,N_3762);
and U4000 (N_4000,N_3888,N_3877);
xnor U4001 (N_4001,N_3905,N_3996);
and U4002 (N_4002,N_3897,N_3976);
or U4003 (N_4003,N_3960,N_3952);
and U4004 (N_4004,N_3999,N_3932);
and U4005 (N_4005,N_3938,N_3993);
and U4006 (N_4006,N_3891,N_3933);
and U4007 (N_4007,N_3934,N_3875);
and U4008 (N_4008,N_3882,N_3987);
or U4009 (N_4009,N_3921,N_3935);
nand U4010 (N_4010,N_3964,N_3945);
nor U4011 (N_4011,N_3928,N_3970);
and U4012 (N_4012,N_3948,N_3914);
xnor U4013 (N_4013,N_3925,N_3985);
xor U4014 (N_4014,N_3988,N_3876);
and U4015 (N_4015,N_3965,N_3994);
or U4016 (N_4016,N_3959,N_3881);
or U4017 (N_4017,N_3904,N_3909);
xor U4018 (N_4018,N_3893,N_3930);
nor U4019 (N_4019,N_3951,N_3975);
nor U4020 (N_4020,N_3878,N_3989);
or U4021 (N_4021,N_3941,N_3992);
xnor U4022 (N_4022,N_3957,N_3907);
xnor U4023 (N_4023,N_3984,N_3981);
nor U4024 (N_4024,N_3926,N_3971);
nor U4025 (N_4025,N_3880,N_3968);
nor U4026 (N_4026,N_3887,N_3911);
and U4027 (N_4027,N_3947,N_3885);
nor U4028 (N_4028,N_3943,N_3966);
nor U4029 (N_4029,N_3958,N_3899);
and U4030 (N_4030,N_3903,N_3927);
and U4031 (N_4031,N_3901,N_3922);
nand U4032 (N_4032,N_3955,N_3967);
and U4033 (N_4033,N_3982,N_3979);
nor U4034 (N_4034,N_3990,N_3936);
and U4035 (N_4035,N_3890,N_3913);
xor U4036 (N_4036,N_3961,N_3940);
xor U4037 (N_4037,N_3963,N_3883);
and U4038 (N_4038,N_3973,N_3902);
nand U4039 (N_4039,N_3986,N_3995);
or U4040 (N_4040,N_3910,N_3942);
nor U4041 (N_4041,N_3974,N_3998);
nand U4042 (N_4042,N_3906,N_3946);
and U4043 (N_4043,N_3969,N_3997);
xor U4044 (N_4044,N_3894,N_3962);
nor U4045 (N_4045,N_3953,N_3924);
and U4046 (N_4046,N_3908,N_3978);
and U4047 (N_4047,N_3937,N_3900);
and U4048 (N_4048,N_3949,N_3972);
nor U4049 (N_4049,N_3944,N_3983);
xor U4050 (N_4050,N_3917,N_3923);
and U4051 (N_4051,N_3980,N_3889);
or U4052 (N_4052,N_3954,N_3912);
nor U4053 (N_4053,N_3918,N_3896);
nand U4054 (N_4054,N_3977,N_3920);
xnor U4055 (N_4055,N_3929,N_3898);
xor U4056 (N_4056,N_3916,N_3956);
and U4057 (N_4057,N_3919,N_3886);
or U4058 (N_4058,N_3884,N_3892);
or U4059 (N_4059,N_3939,N_3915);
xor U4060 (N_4060,N_3931,N_3895);
xnor U4061 (N_4061,N_3950,N_3879);
xnor U4062 (N_4062,N_3991,N_3943);
and U4063 (N_4063,N_3976,N_3984);
nand U4064 (N_4064,N_3967,N_3916);
and U4065 (N_4065,N_3994,N_3927);
xnor U4066 (N_4066,N_3921,N_3973);
xor U4067 (N_4067,N_3944,N_3973);
and U4068 (N_4068,N_3999,N_3939);
and U4069 (N_4069,N_3918,N_3884);
nand U4070 (N_4070,N_3892,N_3888);
nor U4071 (N_4071,N_3948,N_3925);
or U4072 (N_4072,N_3995,N_3925);
nand U4073 (N_4073,N_3902,N_3986);
nand U4074 (N_4074,N_3937,N_3944);
nor U4075 (N_4075,N_3878,N_3929);
nor U4076 (N_4076,N_3993,N_3877);
and U4077 (N_4077,N_3960,N_3901);
or U4078 (N_4078,N_3949,N_3948);
nor U4079 (N_4079,N_3896,N_3968);
nor U4080 (N_4080,N_3896,N_3899);
nand U4081 (N_4081,N_3880,N_3910);
nor U4082 (N_4082,N_3930,N_3965);
nor U4083 (N_4083,N_3897,N_3905);
and U4084 (N_4084,N_3930,N_3911);
nand U4085 (N_4085,N_3997,N_3929);
xnor U4086 (N_4086,N_3875,N_3906);
nor U4087 (N_4087,N_3882,N_3909);
nor U4088 (N_4088,N_3890,N_3967);
or U4089 (N_4089,N_3936,N_3914);
nand U4090 (N_4090,N_3976,N_3982);
nand U4091 (N_4091,N_3975,N_3900);
or U4092 (N_4092,N_3886,N_3952);
nand U4093 (N_4093,N_3892,N_3937);
and U4094 (N_4094,N_3968,N_3924);
xor U4095 (N_4095,N_3906,N_3935);
nor U4096 (N_4096,N_3912,N_3905);
nor U4097 (N_4097,N_3993,N_3985);
nor U4098 (N_4098,N_3985,N_3930);
xor U4099 (N_4099,N_3993,N_3880);
or U4100 (N_4100,N_3908,N_3968);
or U4101 (N_4101,N_3928,N_3893);
nand U4102 (N_4102,N_3883,N_3934);
or U4103 (N_4103,N_3924,N_3879);
or U4104 (N_4104,N_3895,N_3939);
or U4105 (N_4105,N_3975,N_3904);
nor U4106 (N_4106,N_3949,N_3894);
nand U4107 (N_4107,N_3885,N_3990);
or U4108 (N_4108,N_3988,N_3894);
and U4109 (N_4109,N_3923,N_3910);
or U4110 (N_4110,N_3998,N_3955);
or U4111 (N_4111,N_3905,N_3941);
nor U4112 (N_4112,N_3893,N_3881);
nor U4113 (N_4113,N_3985,N_3931);
xor U4114 (N_4114,N_3941,N_3900);
nor U4115 (N_4115,N_3922,N_3963);
or U4116 (N_4116,N_3963,N_3994);
and U4117 (N_4117,N_3981,N_3888);
nand U4118 (N_4118,N_3921,N_3999);
nor U4119 (N_4119,N_3993,N_3947);
or U4120 (N_4120,N_3999,N_3916);
xnor U4121 (N_4121,N_3876,N_3986);
and U4122 (N_4122,N_3887,N_3971);
nand U4123 (N_4123,N_3966,N_3924);
and U4124 (N_4124,N_3999,N_3995);
xor U4125 (N_4125,N_4066,N_4001);
nand U4126 (N_4126,N_4079,N_4017);
nand U4127 (N_4127,N_4104,N_4043);
nand U4128 (N_4128,N_4050,N_4119);
nor U4129 (N_4129,N_4120,N_4039);
and U4130 (N_4130,N_4034,N_4071);
and U4131 (N_4131,N_4047,N_4008);
and U4132 (N_4132,N_4056,N_4122);
nand U4133 (N_4133,N_4112,N_4075);
nor U4134 (N_4134,N_4049,N_4085);
and U4135 (N_4135,N_4109,N_4055);
or U4136 (N_4136,N_4123,N_4021);
xor U4137 (N_4137,N_4116,N_4115);
nand U4138 (N_4138,N_4100,N_4087);
xor U4139 (N_4139,N_4108,N_4052);
and U4140 (N_4140,N_4103,N_4026);
nand U4141 (N_4141,N_4003,N_4064);
or U4142 (N_4142,N_4037,N_4076);
nor U4143 (N_4143,N_4083,N_4012);
nand U4144 (N_4144,N_4069,N_4113);
and U4145 (N_4145,N_4054,N_4090);
nand U4146 (N_4146,N_4036,N_4058);
or U4147 (N_4147,N_4009,N_4097);
and U4148 (N_4148,N_4074,N_4081);
or U4149 (N_4149,N_4059,N_4063);
xor U4150 (N_4150,N_4086,N_4088);
xor U4151 (N_4151,N_4073,N_4099);
xor U4152 (N_4152,N_4094,N_4051);
and U4153 (N_4153,N_4044,N_4018);
xor U4154 (N_4154,N_4106,N_4042);
or U4155 (N_4155,N_4060,N_4068);
nand U4156 (N_4156,N_4095,N_4067);
and U4157 (N_4157,N_4062,N_4098);
and U4158 (N_4158,N_4124,N_4048);
nand U4159 (N_4159,N_4031,N_4053);
and U4160 (N_4160,N_4082,N_4013);
nand U4161 (N_4161,N_4016,N_4025);
and U4162 (N_4162,N_4023,N_4107);
and U4163 (N_4163,N_4030,N_4093);
xnor U4164 (N_4164,N_4057,N_4011);
or U4165 (N_4165,N_4015,N_4084);
nand U4166 (N_4166,N_4041,N_4019);
nand U4167 (N_4167,N_4007,N_4061);
xor U4168 (N_4168,N_4070,N_4046);
or U4169 (N_4169,N_4020,N_4101);
and U4170 (N_4170,N_4024,N_4029);
or U4171 (N_4171,N_4027,N_4080);
nand U4172 (N_4172,N_4096,N_4110);
and U4173 (N_4173,N_4035,N_4014);
or U4174 (N_4174,N_4121,N_4072);
xor U4175 (N_4175,N_4102,N_4000);
nand U4176 (N_4176,N_4033,N_4077);
xor U4177 (N_4177,N_4022,N_4091);
or U4178 (N_4178,N_4032,N_4028);
nor U4179 (N_4179,N_4004,N_4114);
nand U4180 (N_4180,N_4089,N_4006);
and U4181 (N_4181,N_4045,N_4002);
nand U4182 (N_4182,N_4078,N_4005);
nand U4183 (N_4183,N_4092,N_4105);
xor U4184 (N_4184,N_4117,N_4038);
nor U4185 (N_4185,N_4111,N_4065);
xor U4186 (N_4186,N_4118,N_4010);
xor U4187 (N_4187,N_4040,N_4080);
and U4188 (N_4188,N_4037,N_4046);
nor U4189 (N_4189,N_4020,N_4016);
nand U4190 (N_4190,N_4085,N_4122);
or U4191 (N_4191,N_4035,N_4101);
and U4192 (N_4192,N_4075,N_4019);
or U4193 (N_4193,N_4073,N_4102);
and U4194 (N_4194,N_4087,N_4027);
xnor U4195 (N_4195,N_4033,N_4050);
nand U4196 (N_4196,N_4028,N_4020);
and U4197 (N_4197,N_4105,N_4029);
xnor U4198 (N_4198,N_4090,N_4062);
nor U4199 (N_4199,N_4114,N_4003);
and U4200 (N_4200,N_4006,N_4064);
xnor U4201 (N_4201,N_4123,N_4053);
xnor U4202 (N_4202,N_4082,N_4079);
nand U4203 (N_4203,N_4080,N_4033);
nor U4204 (N_4204,N_4033,N_4024);
nor U4205 (N_4205,N_4041,N_4040);
xnor U4206 (N_4206,N_4055,N_4078);
nand U4207 (N_4207,N_4036,N_4037);
xnor U4208 (N_4208,N_4038,N_4004);
nor U4209 (N_4209,N_4076,N_4053);
or U4210 (N_4210,N_4094,N_4015);
xnor U4211 (N_4211,N_4074,N_4032);
xor U4212 (N_4212,N_4067,N_4028);
nor U4213 (N_4213,N_4017,N_4004);
or U4214 (N_4214,N_4084,N_4016);
or U4215 (N_4215,N_4060,N_4066);
xor U4216 (N_4216,N_4051,N_4027);
nor U4217 (N_4217,N_4088,N_4066);
nor U4218 (N_4218,N_4099,N_4107);
or U4219 (N_4219,N_4068,N_4045);
or U4220 (N_4220,N_4062,N_4032);
and U4221 (N_4221,N_4086,N_4006);
nand U4222 (N_4222,N_4116,N_4104);
or U4223 (N_4223,N_4019,N_4033);
xnor U4224 (N_4224,N_4029,N_4037);
or U4225 (N_4225,N_4058,N_4008);
and U4226 (N_4226,N_4051,N_4095);
xor U4227 (N_4227,N_4077,N_4090);
and U4228 (N_4228,N_4065,N_4054);
nand U4229 (N_4229,N_4010,N_4043);
nand U4230 (N_4230,N_4080,N_4078);
nand U4231 (N_4231,N_4116,N_4085);
nor U4232 (N_4232,N_4120,N_4109);
and U4233 (N_4233,N_4111,N_4105);
nor U4234 (N_4234,N_4100,N_4023);
nand U4235 (N_4235,N_4026,N_4099);
nand U4236 (N_4236,N_4033,N_4032);
nand U4237 (N_4237,N_4019,N_4083);
xor U4238 (N_4238,N_4007,N_4099);
nor U4239 (N_4239,N_4035,N_4048);
or U4240 (N_4240,N_4104,N_4014);
or U4241 (N_4241,N_4112,N_4015);
nor U4242 (N_4242,N_4005,N_4063);
and U4243 (N_4243,N_4012,N_4018);
nand U4244 (N_4244,N_4004,N_4071);
xnor U4245 (N_4245,N_4059,N_4000);
nor U4246 (N_4246,N_4024,N_4079);
nand U4247 (N_4247,N_4107,N_4003);
nor U4248 (N_4248,N_4001,N_4082);
or U4249 (N_4249,N_4050,N_4003);
or U4250 (N_4250,N_4160,N_4135);
nor U4251 (N_4251,N_4150,N_4221);
and U4252 (N_4252,N_4175,N_4225);
nor U4253 (N_4253,N_4181,N_4220);
nand U4254 (N_4254,N_4137,N_4178);
or U4255 (N_4255,N_4177,N_4223);
and U4256 (N_4256,N_4172,N_4134);
and U4257 (N_4257,N_4179,N_4141);
nor U4258 (N_4258,N_4170,N_4180);
nor U4259 (N_4259,N_4226,N_4143);
or U4260 (N_4260,N_4227,N_4207);
nand U4261 (N_4261,N_4230,N_4128);
xor U4262 (N_4262,N_4197,N_4176);
or U4263 (N_4263,N_4191,N_4182);
nand U4264 (N_4264,N_4156,N_4151);
and U4265 (N_4265,N_4200,N_4140);
xor U4266 (N_4266,N_4217,N_4146);
or U4267 (N_4267,N_4149,N_4167);
nand U4268 (N_4268,N_4171,N_4231);
nor U4269 (N_4269,N_4145,N_4130);
nor U4270 (N_4270,N_4211,N_4152);
xnor U4271 (N_4271,N_4154,N_4189);
or U4272 (N_4272,N_4193,N_4188);
nand U4273 (N_4273,N_4209,N_4237);
and U4274 (N_4274,N_4210,N_4132);
nand U4275 (N_4275,N_4185,N_4214);
nand U4276 (N_4276,N_4184,N_4192);
xor U4277 (N_4277,N_4241,N_4245);
nor U4278 (N_4278,N_4183,N_4224);
or U4279 (N_4279,N_4125,N_4247);
or U4280 (N_4280,N_4163,N_4206);
and U4281 (N_4281,N_4142,N_4239);
xor U4282 (N_4282,N_4153,N_4235);
nand U4283 (N_4283,N_4218,N_4203);
xnor U4284 (N_4284,N_4136,N_4244);
nor U4285 (N_4285,N_4144,N_4169);
nand U4286 (N_4286,N_4139,N_4159);
nand U4287 (N_4287,N_4166,N_4186);
or U4288 (N_4288,N_4155,N_4204);
nor U4289 (N_4289,N_4127,N_4236);
or U4290 (N_4290,N_4162,N_4205);
nor U4291 (N_4291,N_4195,N_4147);
or U4292 (N_4292,N_4165,N_4248);
xnor U4293 (N_4293,N_4238,N_4187);
nor U4294 (N_4294,N_4243,N_4213);
and U4295 (N_4295,N_4229,N_4199);
nor U4296 (N_4296,N_4129,N_4174);
or U4297 (N_4297,N_4158,N_4161);
or U4298 (N_4298,N_4194,N_4131);
xor U4299 (N_4299,N_4126,N_4157);
and U4300 (N_4300,N_4222,N_4198);
and U4301 (N_4301,N_4232,N_4190);
nand U4302 (N_4302,N_4234,N_4216);
and U4303 (N_4303,N_4212,N_4215);
or U4304 (N_4304,N_4240,N_4219);
xor U4305 (N_4305,N_4208,N_4242);
or U4306 (N_4306,N_4228,N_4246);
and U4307 (N_4307,N_4138,N_4133);
nor U4308 (N_4308,N_4233,N_4164);
nor U4309 (N_4309,N_4168,N_4202);
and U4310 (N_4310,N_4196,N_4201);
and U4311 (N_4311,N_4148,N_4173);
xor U4312 (N_4312,N_4249,N_4131);
xnor U4313 (N_4313,N_4246,N_4215);
or U4314 (N_4314,N_4188,N_4186);
xor U4315 (N_4315,N_4214,N_4164);
nand U4316 (N_4316,N_4192,N_4150);
nand U4317 (N_4317,N_4216,N_4164);
nor U4318 (N_4318,N_4202,N_4170);
nor U4319 (N_4319,N_4176,N_4220);
nor U4320 (N_4320,N_4211,N_4214);
xnor U4321 (N_4321,N_4175,N_4239);
or U4322 (N_4322,N_4236,N_4174);
nand U4323 (N_4323,N_4151,N_4228);
or U4324 (N_4324,N_4219,N_4233);
and U4325 (N_4325,N_4240,N_4155);
and U4326 (N_4326,N_4144,N_4175);
and U4327 (N_4327,N_4128,N_4176);
and U4328 (N_4328,N_4191,N_4156);
xor U4329 (N_4329,N_4232,N_4195);
and U4330 (N_4330,N_4162,N_4126);
nor U4331 (N_4331,N_4164,N_4131);
and U4332 (N_4332,N_4151,N_4134);
nor U4333 (N_4333,N_4166,N_4184);
xnor U4334 (N_4334,N_4157,N_4162);
xor U4335 (N_4335,N_4182,N_4248);
xor U4336 (N_4336,N_4181,N_4132);
and U4337 (N_4337,N_4162,N_4227);
nand U4338 (N_4338,N_4144,N_4137);
nor U4339 (N_4339,N_4235,N_4222);
or U4340 (N_4340,N_4172,N_4238);
nand U4341 (N_4341,N_4237,N_4158);
nor U4342 (N_4342,N_4149,N_4248);
xnor U4343 (N_4343,N_4219,N_4191);
xor U4344 (N_4344,N_4164,N_4172);
xnor U4345 (N_4345,N_4167,N_4247);
xor U4346 (N_4346,N_4163,N_4166);
nor U4347 (N_4347,N_4244,N_4220);
nand U4348 (N_4348,N_4176,N_4226);
xnor U4349 (N_4349,N_4216,N_4212);
or U4350 (N_4350,N_4154,N_4131);
nand U4351 (N_4351,N_4185,N_4136);
and U4352 (N_4352,N_4220,N_4141);
xor U4353 (N_4353,N_4190,N_4243);
xor U4354 (N_4354,N_4152,N_4136);
or U4355 (N_4355,N_4137,N_4126);
or U4356 (N_4356,N_4208,N_4151);
nand U4357 (N_4357,N_4215,N_4167);
nor U4358 (N_4358,N_4179,N_4126);
nand U4359 (N_4359,N_4217,N_4232);
xor U4360 (N_4360,N_4199,N_4140);
and U4361 (N_4361,N_4171,N_4162);
nor U4362 (N_4362,N_4209,N_4155);
nand U4363 (N_4363,N_4131,N_4130);
or U4364 (N_4364,N_4219,N_4159);
xnor U4365 (N_4365,N_4205,N_4240);
nor U4366 (N_4366,N_4245,N_4216);
and U4367 (N_4367,N_4206,N_4142);
or U4368 (N_4368,N_4212,N_4170);
xnor U4369 (N_4369,N_4182,N_4152);
or U4370 (N_4370,N_4128,N_4158);
xnor U4371 (N_4371,N_4154,N_4229);
nand U4372 (N_4372,N_4132,N_4208);
and U4373 (N_4373,N_4125,N_4175);
xnor U4374 (N_4374,N_4193,N_4205);
or U4375 (N_4375,N_4267,N_4303);
or U4376 (N_4376,N_4328,N_4312);
xor U4377 (N_4377,N_4313,N_4250);
and U4378 (N_4378,N_4337,N_4289);
xnor U4379 (N_4379,N_4268,N_4264);
and U4380 (N_4380,N_4360,N_4251);
nor U4381 (N_4381,N_4286,N_4342);
nor U4382 (N_4382,N_4253,N_4256);
xnor U4383 (N_4383,N_4353,N_4266);
or U4384 (N_4384,N_4371,N_4295);
xor U4385 (N_4385,N_4316,N_4325);
and U4386 (N_4386,N_4301,N_4284);
nand U4387 (N_4387,N_4338,N_4335);
nand U4388 (N_4388,N_4293,N_4324);
and U4389 (N_4389,N_4346,N_4279);
nand U4390 (N_4390,N_4296,N_4285);
xor U4391 (N_4391,N_4307,N_4300);
nor U4392 (N_4392,N_4321,N_4275);
or U4393 (N_4393,N_4257,N_4314);
nand U4394 (N_4394,N_4323,N_4372);
nand U4395 (N_4395,N_4259,N_4332);
nor U4396 (N_4396,N_4345,N_4298);
nand U4397 (N_4397,N_4356,N_4358);
and U4398 (N_4398,N_4291,N_4331);
nor U4399 (N_4399,N_4344,N_4288);
nor U4400 (N_4400,N_4363,N_4272);
nor U4401 (N_4401,N_4339,N_4359);
and U4402 (N_4402,N_4310,N_4343);
and U4403 (N_4403,N_4355,N_4290);
xor U4404 (N_4404,N_4283,N_4322);
xor U4405 (N_4405,N_4364,N_4333);
nor U4406 (N_4406,N_4281,N_4341);
or U4407 (N_4407,N_4351,N_4287);
xor U4408 (N_4408,N_4318,N_4354);
nand U4409 (N_4409,N_4278,N_4368);
nand U4410 (N_4410,N_4319,N_4302);
xnor U4411 (N_4411,N_4270,N_4326);
nand U4412 (N_4412,N_4265,N_4292);
nor U4413 (N_4413,N_4254,N_4299);
nor U4414 (N_4414,N_4361,N_4304);
and U4415 (N_4415,N_4365,N_4327);
or U4416 (N_4416,N_4306,N_4276);
nor U4417 (N_4417,N_4308,N_4320);
and U4418 (N_4418,N_4374,N_4317);
xnor U4419 (N_4419,N_4309,N_4329);
nand U4420 (N_4420,N_4262,N_4297);
nand U4421 (N_4421,N_4294,N_4357);
nand U4422 (N_4422,N_4271,N_4370);
nand U4423 (N_4423,N_4263,N_4369);
nand U4424 (N_4424,N_4340,N_4269);
or U4425 (N_4425,N_4258,N_4347);
and U4426 (N_4426,N_4311,N_4255);
and U4427 (N_4427,N_4260,N_4273);
nand U4428 (N_4428,N_4362,N_4348);
nand U4429 (N_4429,N_4373,N_4282);
nand U4430 (N_4430,N_4350,N_4261);
nor U4431 (N_4431,N_4367,N_4336);
nand U4432 (N_4432,N_4334,N_4352);
nand U4433 (N_4433,N_4274,N_4330);
and U4434 (N_4434,N_4277,N_4349);
and U4435 (N_4435,N_4366,N_4305);
and U4436 (N_4436,N_4280,N_4252);
nand U4437 (N_4437,N_4315,N_4298);
and U4438 (N_4438,N_4338,N_4332);
or U4439 (N_4439,N_4350,N_4331);
or U4440 (N_4440,N_4317,N_4278);
nand U4441 (N_4441,N_4257,N_4285);
nand U4442 (N_4442,N_4272,N_4296);
xor U4443 (N_4443,N_4269,N_4267);
nand U4444 (N_4444,N_4357,N_4365);
or U4445 (N_4445,N_4359,N_4259);
and U4446 (N_4446,N_4340,N_4359);
and U4447 (N_4447,N_4250,N_4274);
nand U4448 (N_4448,N_4304,N_4253);
and U4449 (N_4449,N_4288,N_4255);
nor U4450 (N_4450,N_4323,N_4359);
nand U4451 (N_4451,N_4290,N_4332);
nand U4452 (N_4452,N_4263,N_4356);
and U4453 (N_4453,N_4294,N_4303);
xor U4454 (N_4454,N_4278,N_4323);
nor U4455 (N_4455,N_4264,N_4273);
and U4456 (N_4456,N_4308,N_4330);
and U4457 (N_4457,N_4270,N_4311);
nor U4458 (N_4458,N_4325,N_4311);
and U4459 (N_4459,N_4282,N_4312);
xor U4460 (N_4460,N_4339,N_4318);
nor U4461 (N_4461,N_4343,N_4251);
nor U4462 (N_4462,N_4348,N_4342);
nor U4463 (N_4463,N_4304,N_4346);
nor U4464 (N_4464,N_4368,N_4294);
and U4465 (N_4465,N_4353,N_4282);
xor U4466 (N_4466,N_4317,N_4333);
xor U4467 (N_4467,N_4365,N_4309);
and U4468 (N_4468,N_4307,N_4263);
xor U4469 (N_4469,N_4282,N_4332);
or U4470 (N_4470,N_4353,N_4325);
and U4471 (N_4471,N_4257,N_4256);
or U4472 (N_4472,N_4280,N_4273);
or U4473 (N_4473,N_4271,N_4266);
and U4474 (N_4474,N_4371,N_4360);
nor U4475 (N_4475,N_4297,N_4320);
and U4476 (N_4476,N_4319,N_4296);
and U4477 (N_4477,N_4332,N_4286);
nand U4478 (N_4478,N_4366,N_4270);
nand U4479 (N_4479,N_4270,N_4342);
nand U4480 (N_4480,N_4370,N_4321);
xor U4481 (N_4481,N_4330,N_4300);
nand U4482 (N_4482,N_4282,N_4306);
xor U4483 (N_4483,N_4317,N_4327);
nand U4484 (N_4484,N_4316,N_4250);
xnor U4485 (N_4485,N_4283,N_4278);
or U4486 (N_4486,N_4349,N_4357);
and U4487 (N_4487,N_4309,N_4314);
or U4488 (N_4488,N_4307,N_4295);
xnor U4489 (N_4489,N_4342,N_4287);
or U4490 (N_4490,N_4296,N_4259);
xor U4491 (N_4491,N_4343,N_4322);
nor U4492 (N_4492,N_4361,N_4294);
and U4493 (N_4493,N_4276,N_4264);
and U4494 (N_4494,N_4327,N_4345);
or U4495 (N_4495,N_4316,N_4313);
nand U4496 (N_4496,N_4274,N_4296);
nor U4497 (N_4497,N_4324,N_4276);
and U4498 (N_4498,N_4284,N_4293);
xnor U4499 (N_4499,N_4349,N_4340);
and U4500 (N_4500,N_4414,N_4413);
and U4501 (N_4501,N_4480,N_4479);
nor U4502 (N_4502,N_4440,N_4443);
xor U4503 (N_4503,N_4395,N_4436);
nand U4504 (N_4504,N_4494,N_4489);
nand U4505 (N_4505,N_4411,N_4486);
or U4506 (N_4506,N_4406,N_4426);
xnor U4507 (N_4507,N_4447,N_4485);
nor U4508 (N_4508,N_4460,N_4476);
nand U4509 (N_4509,N_4498,N_4427);
nor U4510 (N_4510,N_4449,N_4496);
nor U4511 (N_4511,N_4439,N_4474);
or U4512 (N_4512,N_4483,N_4448);
xor U4513 (N_4513,N_4451,N_4377);
nand U4514 (N_4514,N_4499,N_4469);
nand U4515 (N_4515,N_4487,N_4401);
xnor U4516 (N_4516,N_4432,N_4456);
nor U4517 (N_4517,N_4417,N_4389);
or U4518 (N_4518,N_4492,N_4379);
nor U4519 (N_4519,N_4415,N_4420);
xnor U4520 (N_4520,N_4402,N_4382);
or U4521 (N_4521,N_4444,N_4429);
and U4522 (N_4522,N_4386,N_4446);
xnor U4523 (N_4523,N_4468,N_4385);
nor U4524 (N_4524,N_4473,N_4454);
xnor U4525 (N_4525,N_4418,N_4384);
nand U4526 (N_4526,N_4438,N_4394);
nand U4527 (N_4527,N_4428,N_4422);
or U4528 (N_4528,N_4416,N_4390);
nor U4529 (N_4529,N_4441,N_4431);
xor U4530 (N_4530,N_4419,N_4388);
xor U4531 (N_4531,N_4392,N_4435);
and U4532 (N_4532,N_4430,N_4493);
nand U4533 (N_4533,N_4387,N_4465);
nor U4534 (N_4534,N_4397,N_4378);
nand U4535 (N_4535,N_4490,N_4433);
and U4536 (N_4536,N_4405,N_4455);
and U4537 (N_4537,N_4457,N_4407);
and U4538 (N_4538,N_4412,N_4408);
nand U4539 (N_4539,N_4383,N_4409);
nand U4540 (N_4540,N_4396,N_4475);
xor U4541 (N_4541,N_4458,N_4434);
and U4542 (N_4542,N_4467,N_4404);
or U4543 (N_4543,N_4495,N_4453);
xor U4544 (N_4544,N_4472,N_4464);
nand U4545 (N_4545,N_4463,N_4452);
xnor U4546 (N_4546,N_4484,N_4471);
or U4547 (N_4547,N_4425,N_4470);
nand U4548 (N_4548,N_4375,N_4400);
nand U4549 (N_4549,N_4466,N_4477);
or U4550 (N_4550,N_4421,N_4393);
xor U4551 (N_4551,N_4437,N_4423);
nand U4552 (N_4552,N_4461,N_4462);
or U4553 (N_4553,N_4399,N_4478);
nand U4554 (N_4554,N_4445,N_4424);
nor U4555 (N_4555,N_4491,N_4376);
and U4556 (N_4556,N_4391,N_4497);
and U4557 (N_4557,N_4482,N_4481);
nor U4558 (N_4558,N_4459,N_4380);
and U4559 (N_4559,N_4410,N_4381);
nand U4560 (N_4560,N_4442,N_4488);
or U4561 (N_4561,N_4398,N_4403);
or U4562 (N_4562,N_4450,N_4398);
xnor U4563 (N_4563,N_4463,N_4455);
xor U4564 (N_4564,N_4481,N_4499);
xnor U4565 (N_4565,N_4483,N_4379);
or U4566 (N_4566,N_4409,N_4447);
nand U4567 (N_4567,N_4479,N_4381);
and U4568 (N_4568,N_4495,N_4446);
xor U4569 (N_4569,N_4484,N_4470);
and U4570 (N_4570,N_4416,N_4387);
xor U4571 (N_4571,N_4497,N_4459);
or U4572 (N_4572,N_4383,N_4480);
xor U4573 (N_4573,N_4379,N_4403);
xor U4574 (N_4574,N_4484,N_4431);
or U4575 (N_4575,N_4480,N_4394);
nand U4576 (N_4576,N_4485,N_4475);
nand U4577 (N_4577,N_4453,N_4416);
or U4578 (N_4578,N_4401,N_4407);
or U4579 (N_4579,N_4479,N_4448);
xor U4580 (N_4580,N_4407,N_4438);
xor U4581 (N_4581,N_4435,N_4465);
nand U4582 (N_4582,N_4388,N_4440);
xnor U4583 (N_4583,N_4452,N_4494);
or U4584 (N_4584,N_4422,N_4444);
or U4585 (N_4585,N_4438,N_4442);
nor U4586 (N_4586,N_4442,N_4454);
xnor U4587 (N_4587,N_4421,N_4377);
and U4588 (N_4588,N_4423,N_4493);
nand U4589 (N_4589,N_4438,N_4401);
xnor U4590 (N_4590,N_4477,N_4420);
xnor U4591 (N_4591,N_4480,N_4417);
or U4592 (N_4592,N_4379,N_4490);
or U4593 (N_4593,N_4466,N_4487);
nor U4594 (N_4594,N_4417,N_4423);
or U4595 (N_4595,N_4378,N_4398);
or U4596 (N_4596,N_4480,N_4495);
xnor U4597 (N_4597,N_4397,N_4431);
nand U4598 (N_4598,N_4389,N_4439);
and U4599 (N_4599,N_4418,N_4455);
nor U4600 (N_4600,N_4484,N_4377);
nor U4601 (N_4601,N_4424,N_4411);
nand U4602 (N_4602,N_4410,N_4434);
or U4603 (N_4603,N_4445,N_4406);
nor U4604 (N_4604,N_4496,N_4473);
or U4605 (N_4605,N_4454,N_4477);
nand U4606 (N_4606,N_4462,N_4493);
nand U4607 (N_4607,N_4494,N_4388);
nand U4608 (N_4608,N_4480,N_4400);
nor U4609 (N_4609,N_4457,N_4428);
and U4610 (N_4610,N_4396,N_4491);
xnor U4611 (N_4611,N_4498,N_4429);
nor U4612 (N_4612,N_4461,N_4385);
and U4613 (N_4613,N_4382,N_4447);
and U4614 (N_4614,N_4454,N_4381);
nor U4615 (N_4615,N_4473,N_4468);
nand U4616 (N_4616,N_4455,N_4430);
or U4617 (N_4617,N_4436,N_4406);
nand U4618 (N_4618,N_4391,N_4385);
nor U4619 (N_4619,N_4484,N_4442);
xnor U4620 (N_4620,N_4490,N_4436);
xnor U4621 (N_4621,N_4493,N_4401);
nand U4622 (N_4622,N_4455,N_4382);
or U4623 (N_4623,N_4395,N_4378);
or U4624 (N_4624,N_4460,N_4445);
or U4625 (N_4625,N_4565,N_4526);
nand U4626 (N_4626,N_4621,N_4588);
nand U4627 (N_4627,N_4522,N_4551);
and U4628 (N_4628,N_4513,N_4545);
nor U4629 (N_4629,N_4530,N_4519);
nand U4630 (N_4630,N_4556,N_4546);
xor U4631 (N_4631,N_4575,N_4554);
and U4632 (N_4632,N_4523,N_4533);
xor U4633 (N_4633,N_4518,N_4517);
nand U4634 (N_4634,N_4599,N_4548);
nand U4635 (N_4635,N_4547,N_4514);
nand U4636 (N_4636,N_4613,N_4574);
nand U4637 (N_4637,N_4578,N_4550);
nor U4638 (N_4638,N_4531,N_4596);
or U4639 (N_4639,N_4540,N_4535);
or U4640 (N_4640,N_4584,N_4507);
nor U4641 (N_4641,N_4541,N_4515);
nor U4642 (N_4642,N_4615,N_4538);
xnor U4643 (N_4643,N_4608,N_4604);
xnor U4644 (N_4644,N_4509,N_4580);
and U4645 (N_4645,N_4516,N_4528);
nand U4646 (N_4646,N_4624,N_4500);
nor U4647 (N_4647,N_4563,N_4597);
xnor U4648 (N_4648,N_4567,N_4562);
nor U4649 (N_4649,N_4544,N_4585);
nand U4650 (N_4650,N_4503,N_4537);
xnor U4651 (N_4651,N_4582,N_4594);
nor U4652 (N_4652,N_4549,N_4520);
and U4653 (N_4653,N_4579,N_4610);
nand U4654 (N_4654,N_4502,N_4504);
xor U4655 (N_4655,N_4616,N_4571);
nor U4656 (N_4656,N_4561,N_4570);
xor U4657 (N_4657,N_4501,N_4573);
nand U4658 (N_4658,N_4564,N_4527);
or U4659 (N_4659,N_4593,N_4552);
nor U4660 (N_4660,N_4587,N_4601);
nor U4661 (N_4661,N_4524,N_4569);
xor U4662 (N_4662,N_4622,N_4589);
nor U4663 (N_4663,N_4568,N_4592);
and U4664 (N_4664,N_4559,N_4577);
nand U4665 (N_4665,N_4553,N_4560);
nor U4666 (N_4666,N_4576,N_4521);
or U4667 (N_4667,N_4623,N_4505);
and U4668 (N_4668,N_4572,N_4606);
xnor U4669 (N_4669,N_4591,N_4536);
nor U4670 (N_4670,N_4581,N_4539);
xor U4671 (N_4671,N_4506,N_4590);
nand U4672 (N_4672,N_4614,N_4510);
nand U4673 (N_4673,N_4532,N_4534);
or U4674 (N_4674,N_4609,N_4602);
or U4675 (N_4675,N_4611,N_4583);
nand U4676 (N_4676,N_4620,N_4603);
nand U4677 (N_4677,N_4558,N_4525);
nor U4678 (N_4678,N_4511,N_4607);
and U4679 (N_4679,N_4595,N_4605);
or U4680 (N_4680,N_4566,N_4598);
nor U4681 (N_4681,N_4512,N_4619);
or U4682 (N_4682,N_4586,N_4557);
or U4683 (N_4683,N_4543,N_4618);
nor U4684 (N_4684,N_4529,N_4600);
nand U4685 (N_4685,N_4555,N_4542);
or U4686 (N_4686,N_4508,N_4617);
and U4687 (N_4687,N_4612,N_4504);
nor U4688 (N_4688,N_4523,N_4603);
nand U4689 (N_4689,N_4529,N_4585);
or U4690 (N_4690,N_4579,N_4556);
nand U4691 (N_4691,N_4609,N_4591);
and U4692 (N_4692,N_4522,N_4532);
nor U4693 (N_4693,N_4588,N_4527);
nor U4694 (N_4694,N_4566,N_4537);
nor U4695 (N_4695,N_4592,N_4591);
or U4696 (N_4696,N_4570,N_4539);
and U4697 (N_4697,N_4533,N_4503);
or U4698 (N_4698,N_4510,N_4591);
nand U4699 (N_4699,N_4501,N_4509);
and U4700 (N_4700,N_4619,N_4501);
nor U4701 (N_4701,N_4511,N_4532);
or U4702 (N_4702,N_4553,N_4608);
nor U4703 (N_4703,N_4537,N_4519);
xnor U4704 (N_4704,N_4593,N_4535);
and U4705 (N_4705,N_4580,N_4515);
xnor U4706 (N_4706,N_4560,N_4575);
and U4707 (N_4707,N_4509,N_4505);
or U4708 (N_4708,N_4562,N_4591);
xnor U4709 (N_4709,N_4550,N_4500);
or U4710 (N_4710,N_4604,N_4520);
nor U4711 (N_4711,N_4578,N_4607);
nand U4712 (N_4712,N_4554,N_4590);
or U4713 (N_4713,N_4585,N_4564);
or U4714 (N_4714,N_4555,N_4601);
nand U4715 (N_4715,N_4575,N_4613);
and U4716 (N_4716,N_4542,N_4514);
nand U4717 (N_4717,N_4621,N_4607);
nand U4718 (N_4718,N_4559,N_4580);
nand U4719 (N_4719,N_4567,N_4570);
or U4720 (N_4720,N_4610,N_4544);
or U4721 (N_4721,N_4526,N_4502);
xor U4722 (N_4722,N_4569,N_4592);
xor U4723 (N_4723,N_4543,N_4616);
and U4724 (N_4724,N_4588,N_4614);
or U4725 (N_4725,N_4524,N_4549);
nand U4726 (N_4726,N_4538,N_4561);
xnor U4727 (N_4727,N_4560,N_4597);
and U4728 (N_4728,N_4598,N_4590);
or U4729 (N_4729,N_4614,N_4619);
or U4730 (N_4730,N_4531,N_4569);
and U4731 (N_4731,N_4524,N_4555);
or U4732 (N_4732,N_4553,N_4554);
or U4733 (N_4733,N_4535,N_4577);
nand U4734 (N_4734,N_4536,N_4595);
or U4735 (N_4735,N_4575,N_4604);
or U4736 (N_4736,N_4622,N_4553);
nor U4737 (N_4737,N_4564,N_4513);
and U4738 (N_4738,N_4609,N_4505);
and U4739 (N_4739,N_4522,N_4546);
or U4740 (N_4740,N_4582,N_4612);
nor U4741 (N_4741,N_4510,N_4602);
nand U4742 (N_4742,N_4536,N_4557);
xor U4743 (N_4743,N_4568,N_4527);
xnor U4744 (N_4744,N_4550,N_4621);
or U4745 (N_4745,N_4576,N_4593);
xor U4746 (N_4746,N_4551,N_4513);
or U4747 (N_4747,N_4591,N_4551);
or U4748 (N_4748,N_4609,N_4513);
nor U4749 (N_4749,N_4585,N_4569);
or U4750 (N_4750,N_4636,N_4670);
or U4751 (N_4751,N_4679,N_4699);
or U4752 (N_4752,N_4633,N_4680);
or U4753 (N_4753,N_4732,N_4738);
nor U4754 (N_4754,N_4712,N_4646);
nand U4755 (N_4755,N_4725,N_4627);
and U4756 (N_4756,N_4630,N_4683);
xor U4757 (N_4757,N_4705,N_4717);
nor U4758 (N_4758,N_4746,N_4673);
nand U4759 (N_4759,N_4688,N_4745);
nor U4760 (N_4760,N_4628,N_4710);
xnor U4761 (N_4761,N_4719,N_4643);
nand U4762 (N_4762,N_4690,N_4713);
or U4763 (N_4763,N_4653,N_4703);
nand U4764 (N_4764,N_4720,N_4747);
nand U4765 (N_4765,N_4728,N_4744);
xor U4766 (N_4766,N_4685,N_4651);
nor U4767 (N_4767,N_4635,N_4715);
xnor U4768 (N_4768,N_4639,N_4693);
nor U4769 (N_4769,N_4748,N_4743);
nor U4770 (N_4770,N_4659,N_4649);
and U4771 (N_4771,N_4727,N_4644);
nand U4772 (N_4772,N_4736,N_4637);
or U4773 (N_4773,N_4626,N_4678);
nand U4774 (N_4774,N_4682,N_4657);
nor U4775 (N_4775,N_4625,N_4714);
and U4776 (N_4776,N_4739,N_4735);
or U4777 (N_4777,N_4629,N_4648);
or U4778 (N_4778,N_4675,N_4691);
xor U4779 (N_4779,N_4642,N_4668);
xnor U4780 (N_4780,N_4737,N_4672);
and U4781 (N_4781,N_4734,N_4687);
nand U4782 (N_4782,N_4632,N_4671);
and U4783 (N_4783,N_4650,N_4658);
xor U4784 (N_4784,N_4723,N_4697);
or U4785 (N_4785,N_4711,N_4689);
nor U4786 (N_4786,N_4665,N_4662);
nor U4787 (N_4787,N_4702,N_4647);
or U4788 (N_4788,N_4641,N_4656);
and U4789 (N_4789,N_4631,N_4716);
or U4790 (N_4790,N_4726,N_4700);
xnor U4791 (N_4791,N_4664,N_4718);
or U4792 (N_4792,N_4684,N_4731);
xor U4793 (N_4793,N_4701,N_4749);
nor U4794 (N_4794,N_4645,N_4741);
or U4795 (N_4795,N_4655,N_4709);
and U4796 (N_4796,N_4695,N_4694);
nand U4797 (N_4797,N_4707,N_4706);
xnor U4798 (N_4798,N_4724,N_4667);
nor U4799 (N_4799,N_4661,N_4704);
nand U4800 (N_4800,N_4674,N_4742);
nand U4801 (N_4801,N_4652,N_4696);
nand U4802 (N_4802,N_4666,N_4676);
xor U4803 (N_4803,N_4660,N_4686);
nor U4804 (N_4804,N_4634,N_4708);
or U4805 (N_4805,N_4698,N_4729);
nor U4806 (N_4806,N_4677,N_4740);
or U4807 (N_4807,N_4669,N_4638);
nor U4808 (N_4808,N_4721,N_4722);
xor U4809 (N_4809,N_4730,N_4640);
nand U4810 (N_4810,N_4654,N_4692);
or U4811 (N_4811,N_4663,N_4681);
and U4812 (N_4812,N_4733,N_4674);
nand U4813 (N_4813,N_4626,N_4664);
nor U4814 (N_4814,N_4686,N_4695);
nor U4815 (N_4815,N_4654,N_4718);
nand U4816 (N_4816,N_4632,N_4670);
xor U4817 (N_4817,N_4664,N_4650);
and U4818 (N_4818,N_4737,N_4708);
or U4819 (N_4819,N_4743,N_4707);
and U4820 (N_4820,N_4725,N_4723);
nand U4821 (N_4821,N_4672,N_4630);
xor U4822 (N_4822,N_4696,N_4638);
nor U4823 (N_4823,N_4664,N_4737);
and U4824 (N_4824,N_4735,N_4665);
xnor U4825 (N_4825,N_4729,N_4661);
nor U4826 (N_4826,N_4734,N_4717);
and U4827 (N_4827,N_4690,N_4701);
nor U4828 (N_4828,N_4664,N_4742);
and U4829 (N_4829,N_4748,N_4679);
or U4830 (N_4830,N_4714,N_4709);
and U4831 (N_4831,N_4640,N_4637);
or U4832 (N_4832,N_4681,N_4643);
nand U4833 (N_4833,N_4658,N_4690);
xor U4834 (N_4834,N_4689,N_4714);
and U4835 (N_4835,N_4629,N_4683);
and U4836 (N_4836,N_4634,N_4646);
and U4837 (N_4837,N_4657,N_4669);
xnor U4838 (N_4838,N_4655,N_4734);
nand U4839 (N_4839,N_4719,N_4683);
and U4840 (N_4840,N_4694,N_4741);
xnor U4841 (N_4841,N_4679,N_4648);
nand U4842 (N_4842,N_4701,N_4683);
nand U4843 (N_4843,N_4639,N_4687);
or U4844 (N_4844,N_4637,N_4691);
xnor U4845 (N_4845,N_4734,N_4657);
nand U4846 (N_4846,N_4744,N_4647);
or U4847 (N_4847,N_4743,N_4686);
xor U4848 (N_4848,N_4664,N_4700);
nor U4849 (N_4849,N_4696,N_4671);
xnor U4850 (N_4850,N_4749,N_4696);
nand U4851 (N_4851,N_4682,N_4702);
or U4852 (N_4852,N_4744,N_4638);
or U4853 (N_4853,N_4749,N_4726);
or U4854 (N_4854,N_4717,N_4670);
xnor U4855 (N_4855,N_4686,N_4634);
xor U4856 (N_4856,N_4696,N_4692);
or U4857 (N_4857,N_4719,N_4663);
xnor U4858 (N_4858,N_4668,N_4721);
nor U4859 (N_4859,N_4636,N_4658);
and U4860 (N_4860,N_4703,N_4727);
and U4861 (N_4861,N_4652,N_4628);
xnor U4862 (N_4862,N_4637,N_4704);
and U4863 (N_4863,N_4748,N_4683);
and U4864 (N_4864,N_4681,N_4653);
and U4865 (N_4865,N_4713,N_4665);
and U4866 (N_4866,N_4657,N_4647);
and U4867 (N_4867,N_4725,N_4669);
and U4868 (N_4868,N_4649,N_4663);
xnor U4869 (N_4869,N_4745,N_4723);
nor U4870 (N_4870,N_4656,N_4646);
and U4871 (N_4871,N_4716,N_4693);
nand U4872 (N_4872,N_4739,N_4749);
and U4873 (N_4873,N_4704,N_4641);
nand U4874 (N_4874,N_4635,N_4723);
and U4875 (N_4875,N_4799,N_4797);
nand U4876 (N_4876,N_4778,N_4828);
and U4877 (N_4877,N_4761,N_4763);
nand U4878 (N_4878,N_4870,N_4768);
nand U4879 (N_4879,N_4845,N_4758);
xor U4880 (N_4880,N_4848,N_4788);
and U4881 (N_4881,N_4809,N_4847);
and U4882 (N_4882,N_4813,N_4834);
or U4883 (N_4883,N_4760,N_4868);
and U4884 (N_4884,N_4772,N_4825);
and U4885 (N_4885,N_4829,N_4766);
or U4886 (N_4886,N_4754,N_4780);
nand U4887 (N_4887,N_4789,N_4863);
or U4888 (N_4888,N_4805,N_4846);
or U4889 (N_4889,N_4802,N_4785);
nand U4890 (N_4890,N_4762,N_4752);
or U4891 (N_4891,N_4804,N_4801);
nand U4892 (N_4892,N_4832,N_4798);
and U4893 (N_4893,N_4755,N_4751);
xor U4894 (N_4894,N_4810,N_4874);
nand U4895 (N_4895,N_4857,N_4869);
nor U4896 (N_4896,N_4855,N_4854);
or U4897 (N_4897,N_4753,N_4796);
or U4898 (N_4898,N_4795,N_4820);
or U4899 (N_4899,N_4865,N_4871);
and U4900 (N_4900,N_4836,N_4843);
nor U4901 (N_4901,N_4852,N_4819);
and U4902 (N_4902,N_4759,N_4812);
and U4903 (N_4903,N_4841,N_4849);
and U4904 (N_4904,N_4850,N_4764);
nor U4905 (N_4905,N_4833,N_4784);
or U4906 (N_4906,N_4757,N_4858);
or U4907 (N_4907,N_4864,N_4808);
xnor U4908 (N_4908,N_4866,N_4774);
nand U4909 (N_4909,N_4822,N_4816);
xnor U4910 (N_4910,N_4779,N_4769);
or U4911 (N_4911,N_4830,N_4826);
nor U4912 (N_4912,N_4790,N_4807);
xor U4913 (N_4913,N_4803,N_4842);
nand U4914 (N_4914,N_4853,N_4838);
and U4915 (N_4915,N_4765,N_4787);
nand U4916 (N_4916,N_4756,N_4811);
nor U4917 (N_4917,N_4775,N_4851);
or U4918 (N_4918,N_4792,N_4835);
xor U4919 (N_4919,N_4817,N_4873);
or U4920 (N_4920,N_4860,N_4859);
nor U4921 (N_4921,N_4861,N_4862);
and U4922 (N_4922,N_4791,N_4773);
nor U4923 (N_4923,N_4793,N_4837);
and U4924 (N_4924,N_4786,N_4794);
nand U4925 (N_4925,N_4839,N_4777);
nor U4926 (N_4926,N_4783,N_4831);
nand U4927 (N_4927,N_4776,N_4815);
xor U4928 (N_4928,N_4840,N_4806);
and U4929 (N_4929,N_4821,N_4771);
and U4930 (N_4930,N_4823,N_4750);
nor U4931 (N_4931,N_4856,N_4827);
and U4932 (N_4932,N_4814,N_4818);
nor U4933 (N_4933,N_4767,N_4781);
nor U4934 (N_4934,N_4844,N_4782);
and U4935 (N_4935,N_4800,N_4770);
and U4936 (N_4936,N_4824,N_4867);
or U4937 (N_4937,N_4872,N_4764);
xnor U4938 (N_4938,N_4866,N_4773);
or U4939 (N_4939,N_4799,N_4856);
and U4940 (N_4940,N_4792,N_4782);
and U4941 (N_4941,N_4757,N_4754);
xor U4942 (N_4942,N_4834,N_4755);
or U4943 (N_4943,N_4835,N_4827);
xnor U4944 (N_4944,N_4854,N_4813);
xnor U4945 (N_4945,N_4831,N_4778);
xnor U4946 (N_4946,N_4768,N_4833);
nand U4947 (N_4947,N_4775,N_4792);
and U4948 (N_4948,N_4861,N_4769);
nand U4949 (N_4949,N_4860,N_4805);
nand U4950 (N_4950,N_4825,N_4805);
or U4951 (N_4951,N_4756,N_4834);
nor U4952 (N_4952,N_4835,N_4791);
or U4953 (N_4953,N_4758,N_4869);
nand U4954 (N_4954,N_4803,N_4825);
nand U4955 (N_4955,N_4835,N_4755);
or U4956 (N_4956,N_4851,N_4760);
nand U4957 (N_4957,N_4820,N_4857);
nor U4958 (N_4958,N_4791,N_4758);
xnor U4959 (N_4959,N_4808,N_4816);
xor U4960 (N_4960,N_4804,N_4768);
nor U4961 (N_4961,N_4849,N_4809);
or U4962 (N_4962,N_4751,N_4778);
nor U4963 (N_4963,N_4834,N_4838);
nand U4964 (N_4964,N_4759,N_4860);
and U4965 (N_4965,N_4832,N_4828);
or U4966 (N_4966,N_4763,N_4870);
and U4967 (N_4967,N_4785,N_4796);
nor U4968 (N_4968,N_4760,N_4805);
nand U4969 (N_4969,N_4764,N_4754);
nand U4970 (N_4970,N_4847,N_4806);
and U4971 (N_4971,N_4796,N_4823);
or U4972 (N_4972,N_4779,N_4832);
or U4973 (N_4973,N_4825,N_4830);
or U4974 (N_4974,N_4855,N_4753);
nand U4975 (N_4975,N_4816,N_4832);
nor U4976 (N_4976,N_4850,N_4871);
xor U4977 (N_4977,N_4759,N_4874);
nand U4978 (N_4978,N_4797,N_4802);
xnor U4979 (N_4979,N_4756,N_4812);
or U4980 (N_4980,N_4829,N_4857);
or U4981 (N_4981,N_4865,N_4838);
and U4982 (N_4982,N_4806,N_4823);
nor U4983 (N_4983,N_4830,N_4842);
or U4984 (N_4984,N_4855,N_4800);
xnor U4985 (N_4985,N_4829,N_4826);
nand U4986 (N_4986,N_4824,N_4792);
xor U4987 (N_4987,N_4840,N_4773);
nor U4988 (N_4988,N_4783,N_4757);
or U4989 (N_4989,N_4783,N_4756);
xor U4990 (N_4990,N_4824,N_4815);
or U4991 (N_4991,N_4826,N_4835);
or U4992 (N_4992,N_4835,N_4846);
or U4993 (N_4993,N_4856,N_4835);
xor U4994 (N_4994,N_4818,N_4831);
nor U4995 (N_4995,N_4792,N_4856);
xor U4996 (N_4996,N_4809,N_4755);
nand U4997 (N_4997,N_4828,N_4823);
nand U4998 (N_4998,N_4825,N_4841);
or U4999 (N_4999,N_4818,N_4777);
xnor U5000 (N_5000,N_4947,N_4987);
and U5001 (N_5001,N_4950,N_4961);
nand U5002 (N_5002,N_4995,N_4893);
nand U5003 (N_5003,N_4967,N_4907);
nand U5004 (N_5004,N_4891,N_4926);
xnor U5005 (N_5005,N_4953,N_4906);
and U5006 (N_5006,N_4973,N_4899);
xor U5007 (N_5007,N_4978,N_4990);
xor U5008 (N_5008,N_4911,N_4902);
and U5009 (N_5009,N_4933,N_4974);
nand U5010 (N_5010,N_4915,N_4940);
nand U5011 (N_5011,N_4979,N_4981);
nand U5012 (N_5012,N_4875,N_4991);
nor U5013 (N_5013,N_4901,N_4890);
nand U5014 (N_5014,N_4900,N_4957);
and U5015 (N_5015,N_4916,N_4912);
nor U5016 (N_5016,N_4887,N_4898);
or U5017 (N_5017,N_4982,N_4993);
xor U5018 (N_5018,N_4892,N_4980);
nand U5019 (N_5019,N_4983,N_4876);
or U5020 (N_5020,N_4917,N_4884);
xnor U5021 (N_5021,N_4942,N_4975);
xor U5022 (N_5022,N_4971,N_4963);
and U5023 (N_5023,N_4996,N_4938);
and U5024 (N_5024,N_4896,N_4984);
nand U5025 (N_5025,N_4989,N_4885);
and U5026 (N_5026,N_4986,N_4949);
xnor U5027 (N_5027,N_4925,N_4994);
xnor U5028 (N_5028,N_4970,N_4913);
nand U5029 (N_5029,N_4932,N_4905);
xor U5030 (N_5030,N_4934,N_4877);
xnor U5031 (N_5031,N_4883,N_4965);
xnor U5032 (N_5032,N_4927,N_4960);
xnor U5033 (N_5033,N_4923,N_4937);
nor U5034 (N_5034,N_4886,N_4944);
nor U5035 (N_5035,N_4954,N_4945);
and U5036 (N_5036,N_4959,N_4968);
nor U5037 (N_5037,N_4956,N_4952);
and U5038 (N_5038,N_4939,N_4999);
and U5039 (N_5039,N_4977,N_4921);
nor U5040 (N_5040,N_4879,N_4951);
and U5041 (N_5041,N_4918,N_4880);
or U5042 (N_5042,N_4929,N_4888);
and U5043 (N_5043,N_4988,N_4969);
xor U5044 (N_5044,N_4928,N_4962);
nand U5045 (N_5045,N_4935,N_4936);
or U5046 (N_5046,N_4976,N_4895);
nand U5047 (N_5047,N_4903,N_4943);
nand U5048 (N_5048,N_4958,N_4992);
nand U5049 (N_5049,N_4998,N_4919);
nand U5050 (N_5050,N_4972,N_4908);
nand U5051 (N_5051,N_4966,N_4897);
nand U5052 (N_5052,N_4920,N_4955);
and U5053 (N_5053,N_4997,N_4881);
and U5054 (N_5054,N_4985,N_4930);
nand U5055 (N_5055,N_4922,N_4931);
and U5056 (N_5056,N_4946,N_4894);
nand U5057 (N_5057,N_4948,N_4941);
nor U5058 (N_5058,N_4924,N_4964);
or U5059 (N_5059,N_4914,N_4889);
xor U5060 (N_5060,N_4909,N_4910);
or U5061 (N_5061,N_4904,N_4878);
nor U5062 (N_5062,N_4882,N_4912);
and U5063 (N_5063,N_4910,N_4991);
or U5064 (N_5064,N_4922,N_4888);
nand U5065 (N_5065,N_4929,N_4913);
xnor U5066 (N_5066,N_4879,N_4977);
or U5067 (N_5067,N_4956,N_4898);
nand U5068 (N_5068,N_4991,N_4946);
nand U5069 (N_5069,N_4950,N_4936);
and U5070 (N_5070,N_4901,N_4907);
nand U5071 (N_5071,N_4984,N_4915);
and U5072 (N_5072,N_4928,N_4939);
nand U5073 (N_5073,N_4987,N_4974);
or U5074 (N_5074,N_4964,N_4916);
xnor U5075 (N_5075,N_4936,N_4998);
nor U5076 (N_5076,N_4955,N_4974);
xnor U5077 (N_5077,N_4954,N_4916);
xnor U5078 (N_5078,N_4940,N_4963);
nand U5079 (N_5079,N_4974,N_4914);
or U5080 (N_5080,N_4907,N_4936);
xnor U5081 (N_5081,N_4905,N_4890);
nor U5082 (N_5082,N_4917,N_4977);
nor U5083 (N_5083,N_4935,N_4998);
xor U5084 (N_5084,N_4903,N_4966);
nor U5085 (N_5085,N_4878,N_4933);
and U5086 (N_5086,N_4952,N_4897);
and U5087 (N_5087,N_4980,N_4930);
nand U5088 (N_5088,N_4892,N_4946);
or U5089 (N_5089,N_4989,N_4877);
xnor U5090 (N_5090,N_4969,N_4942);
or U5091 (N_5091,N_4909,N_4943);
xor U5092 (N_5092,N_4890,N_4886);
and U5093 (N_5093,N_4970,N_4976);
nand U5094 (N_5094,N_4962,N_4989);
or U5095 (N_5095,N_4913,N_4927);
or U5096 (N_5096,N_4878,N_4930);
or U5097 (N_5097,N_4899,N_4993);
nand U5098 (N_5098,N_4934,N_4908);
nor U5099 (N_5099,N_4964,N_4900);
xor U5100 (N_5100,N_4932,N_4972);
and U5101 (N_5101,N_4933,N_4965);
and U5102 (N_5102,N_4957,N_4967);
nand U5103 (N_5103,N_4938,N_4890);
nand U5104 (N_5104,N_4967,N_4996);
or U5105 (N_5105,N_4888,N_4954);
xor U5106 (N_5106,N_4881,N_4889);
and U5107 (N_5107,N_4886,N_4989);
and U5108 (N_5108,N_4983,N_4911);
nor U5109 (N_5109,N_4899,N_4924);
nand U5110 (N_5110,N_4947,N_4876);
nor U5111 (N_5111,N_4982,N_4919);
nand U5112 (N_5112,N_4916,N_4968);
or U5113 (N_5113,N_4977,N_4899);
xor U5114 (N_5114,N_4988,N_4940);
or U5115 (N_5115,N_4922,N_4976);
nand U5116 (N_5116,N_4919,N_4898);
or U5117 (N_5117,N_4931,N_4936);
nand U5118 (N_5118,N_4916,N_4927);
and U5119 (N_5119,N_4880,N_4973);
or U5120 (N_5120,N_4915,N_4952);
nor U5121 (N_5121,N_4932,N_4916);
nor U5122 (N_5122,N_4953,N_4917);
nand U5123 (N_5123,N_4903,N_4902);
nor U5124 (N_5124,N_4912,N_4990);
or U5125 (N_5125,N_5098,N_5082);
nand U5126 (N_5126,N_5010,N_5099);
xor U5127 (N_5127,N_5122,N_5119);
xnor U5128 (N_5128,N_5035,N_5034);
or U5129 (N_5129,N_5039,N_5014);
and U5130 (N_5130,N_5065,N_5053);
or U5131 (N_5131,N_5118,N_5021);
or U5132 (N_5132,N_5005,N_5025);
or U5133 (N_5133,N_5093,N_5070);
and U5134 (N_5134,N_5064,N_5109);
nor U5135 (N_5135,N_5084,N_5113);
or U5136 (N_5136,N_5016,N_5024);
or U5137 (N_5137,N_5031,N_5003);
nor U5138 (N_5138,N_5043,N_5061);
xnor U5139 (N_5139,N_5076,N_5048);
xor U5140 (N_5140,N_5063,N_5011);
and U5141 (N_5141,N_5067,N_5046);
xor U5142 (N_5142,N_5094,N_5042);
or U5143 (N_5143,N_5085,N_5102);
nor U5144 (N_5144,N_5000,N_5121);
and U5145 (N_5145,N_5090,N_5086);
nor U5146 (N_5146,N_5092,N_5052);
nor U5147 (N_5147,N_5038,N_5020);
and U5148 (N_5148,N_5032,N_5103);
or U5149 (N_5149,N_5105,N_5058);
and U5150 (N_5150,N_5080,N_5059);
xnor U5151 (N_5151,N_5047,N_5002);
xnor U5152 (N_5152,N_5041,N_5069);
nor U5153 (N_5153,N_5012,N_5120);
or U5154 (N_5154,N_5007,N_5115);
xnor U5155 (N_5155,N_5029,N_5072);
or U5156 (N_5156,N_5106,N_5017);
nand U5157 (N_5157,N_5123,N_5107);
nor U5158 (N_5158,N_5050,N_5027);
xor U5159 (N_5159,N_5019,N_5079);
and U5160 (N_5160,N_5112,N_5101);
nor U5161 (N_5161,N_5008,N_5028);
nand U5162 (N_5162,N_5051,N_5055);
nand U5163 (N_5163,N_5104,N_5088);
or U5164 (N_5164,N_5036,N_5004);
nand U5165 (N_5165,N_5013,N_5081);
and U5166 (N_5166,N_5030,N_5040);
xor U5167 (N_5167,N_5056,N_5097);
xor U5168 (N_5168,N_5015,N_5111);
nand U5169 (N_5169,N_5057,N_5033);
and U5170 (N_5170,N_5117,N_5062);
nor U5171 (N_5171,N_5116,N_5108);
or U5172 (N_5172,N_5073,N_5006);
xnor U5173 (N_5173,N_5078,N_5083);
and U5174 (N_5174,N_5018,N_5110);
and U5175 (N_5175,N_5044,N_5068);
nor U5176 (N_5176,N_5074,N_5100);
nand U5177 (N_5177,N_5049,N_5095);
nor U5178 (N_5178,N_5077,N_5023);
xnor U5179 (N_5179,N_5045,N_5001);
and U5180 (N_5180,N_5054,N_5114);
nand U5181 (N_5181,N_5066,N_5089);
xnor U5182 (N_5182,N_5124,N_5091);
or U5183 (N_5183,N_5026,N_5022);
xor U5184 (N_5184,N_5060,N_5096);
nor U5185 (N_5185,N_5075,N_5087);
or U5186 (N_5186,N_5009,N_5037);
nor U5187 (N_5187,N_5071,N_5003);
and U5188 (N_5188,N_5057,N_5094);
and U5189 (N_5189,N_5058,N_5076);
and U5190 (N_5190,N_5008,N_5116);
or U5191 (N_5191,N_5046,N_5095);
xor U5192 (N_5192,N_5077,N_5033);
xnor U5193 (N_5193,N_5077,N_5117);
and U5194 (N_5194,N_5032,N_5096);
or U5195 (N_5195,N_5078,N_5029);
xnor U5196 (N_5196,N_5015,N_5100);
nor U5197 (N_5197,N_5078,N_5034);
and U5198 (N_5198,N_5094,N_5010);
and U5199 (N_5199,N_5028,N_5093);
nor U5200 (N_5200,N_5069,N_5076);
nand U5201 (N_5201,N_5118,N_5060);
nand U5202 (N_5202,N_5043,N_5050);
nand U5203 (N_5203,N_5006,N_5054);
and U5204 (N_5204,N_5082,N_5095);
nor U5205 (N_5205,N_5116,N_5009);
and U5206 (N_5206,N_5015,N_5106);
or U5207 (N_5207,N_5079,N_5062);
nor U5208 (N_5208,N_5094,N_5055);
and U5209 (N_5209,N_5020,N_5025);
and U5210 (N_5210,N_5105,N_5121);
or U5211 (N_5211,N_5060,N_5093);
nor U5212 (N_5212,N_5083,N_5055);
and U5213 (N_5213,N_5021,N_5049);
nor U5214 (N_5214,N_5047,N_5059);
nand U5215 (N_5215,N_5032,N_5120);
or U5216 (N_5216,N_5040,N_5078);
xor U5217 (N_5217,N_5093,N_5029);
or U5218 (N_5218,N_5076,N_5026);
or U5219 (N_5219,N_5018,N_5081);
or U5220 (N_5220,N_5026,N_5017);
nand U5221 (N_5221,N_5054,N_5115);
xor U5222 (N_5222,N_5120,N_5074);
and U5223 (N_5223,N_5041,N_5025);
xnor U5224 (N_5224,N_5092,N_5097);
or U5225 (N_5225,N_5120,N_5001);
nor U5226 (N_5226,N_5010,N_5021);
or U5227 (N_5227,N_5001,N_5052);
nor U5228 (N_5228,N_5106,N_5120);
and U5229 (N_5229,N_5089,N_5059);
or U5230 (N_5230,N_5089,N_5036);
nand U5231 (N_5231,N_5089,N_5099);
or U5232 (N_5232,N_5038,N_5111);
nor U5233 (N_5233,N_5124,N_5023);
or U5234 (N_5234,N_5022,N_5102);
nor U5235 (N_5235,N_5073,N_5051);
and U5236 (N_5236,N_5005,N_5120);
or U5237 (N_5237,N_5092,N_5018);
and U5238 (N_5238,N_5121,N_5099);
nor U5239 (N_5239,N_5040,N_5008);
and U5240 (N_5240,N_5075,N_5059);
nor U5241 (N_5241,N_5124,N_5107);
nand U5242 (N_5242,N_5000,N_5098);
xor U5243 (N_5243,N_5097,N_5086);
nand U5244 (N_5244,N_5048,N_5016);
nand U5245 (N_5245,N_5027,N_5040);
and U5246 (N_5246,N_5106,N_5119);
nor U5247 (N_5247,N_5107,N_5009);
nand U5248 (N_5248,N_5085,N_5046);
nor U5249 (N_5249,N_5055,N_5082);
or U5250 (N_5250,N_5207,N_5178);
and U5251 (N_5251,N_5172,N_5232);
and U5252 (N_5252,N_5198,N_5127);
xor U5253 (N_5253,N_5163,N_5228);
xnor U5254 (N_5254,N_5249,N_5225);
nand U5255 (N_5255,N_5210,N_5181);
and U5256 (N_5256,N_5151,N_5153);
and U5257 (N_5257,N_5234,N_5141);
nand U5258 (N_5258,N_5128,N_5227);
or U5259 (N_5259,N_5165,N_5169);
or U5260 (N_5260,N_5215,N_5138);
xor U5261 (N_5261,N_5241,N_5132);
nor U5262 (N_5262,N_5230,N_5161);
xor U5263 (N_5263,N_5221,N_5223);
nand U5264 (N_5264,N_5219,N_5177);
xnor U5265 (N_5265,N_5203,N_5222);
xor U5266 (N_5266,N_5139,N_5231);
and U5267 (N_5267,N_5170,N_5196);
nor U5268 (N_5268,N_5147,N_5125);
nand U5269 (N_5269,N_5166,N_5235);
nor U5270 (N_5270,N_5224,N_5199);
or U5271 (N_5271,N_5173,N_5188);
and U5272 (N_5272,N_5154,N_5145);
and U5273 (N_5273,N_5143,N_5242);
xnor U5274 (N_5274,N_5208,N_5213);
and U5275 (N_5275,N_5229,N_5200);
xor U5276 (N_5276,N_5204,N_5247);
nor U5277 (N_5277,N_5205,N_5137);
nand U5278 (N_5278,N_5244,N_5193);
xnor U5279 (N_5279,N_5136,N_5150);
nor U5280 (N_5280,N_5133,N_5160);
or U5281 (N_5281,N_5212,N_5156);
xnor U5282 (N_5282,N_5202,N_5168);
and U5283 (N_5283,N_5190,N_5246);
or U5284 (N_5284,N_5149,N_5176);
nor U5285 (N_5285,N_5214,N_5233);
nand U5286 (N_5286,N_5201,N_5216);
xnor U5287 (N_5287,N_5180,N_5189);
nand U5288 (N_5288,N_5236,N_5140);
or U5289 (N_5289,N_5146,N_5187);
and U5290 (N_5290,N_5217,N_5148);
or U5291 (N_5291,N_5179,N_5174);
nor U5292 (N_5292,N_5129,N_5182);
and U5293 (N_5293,N_5220,N_5159);
xor U5294 (N_5294,N_5131,N_5183);
xor U5295 (N_5295,N_5164,N_5155);
nand U5296 (N_5296,N_5239,N_5197);
nor U5297 (N_5297,N_5130,N_5237);
xor U5298 (N_5298,N_5175,N_5209);
and U5299 (N_5299,N_5248,N_5195);
and U5300 (N_5300,N_5240,N_5245);
xnor U5301 (N_5301,N_5162,N_5186);
xnor U5302 (N_5302,N_5206,N_5192);
or U5303 (N_5303,N_5218,N_5144);
nand U5304 (N_5304,N_5243,N_5134);
nand U5305 (N_5305,N_5126,N_5158);
xnor U5306 (N_5306,N_5157,N_5184);
nand U5307 (N_5307,N_5211,N_5152);
nand U5308 (N_5308,N_5142,N_5171);
or U5309 (N_5309,N_5191,N_5238);
or U5310 (N_5310,N_5167,N_5226);
nand U5311 (N_5311,N_5194,N_5135);
and U5312 (N_5312,N_5185,N_5202);
and U5313 (N_5313,N_5161,N_5246);
xnor U5314 (N_5314,N_5224,N_5206);
nor U5315 (N_5315,N_5206,N_5191);
xor U5316 (N_5316,N_5146,N_5170);
nand U5317 (N_5317,N_5239,N_5170);
or U5318 (N_5318,N_5187,N_5149);
nor U5319 (N_5319,N_5139,N_5143);
nand U5320 (N_5320,N_5135,N_5236);
nor U5321 (N_5321,N_5211,N_5156);
and U5322 (N_5322,N_5192,N_5169);
nand U5323 (N_5323,N_5138,N_5241);
and U5324 (N_5324,N_5163,N_5227);
or U5325 (N_5325,N_5193,N_5228);
or U5326 (N_5326,N_5193,N_5187);
xor U5327 (N_5327,N_5193,N_5137);
xnor U5328 (N_5328,N_5200,N_5186);
xnor U5329 (N_5329,N_5182,N_5173);
nor U5330 (N_5330,N_5192,N_5185);
or U5331 (N_5331,N_5172,N_5220);
nor U5332 (N_5332,N_5225,N_5179);
nor U5333 (N_5333,N_5169,N_5141);
xnor U5334 (N_5334,N_5150,N_5217);
or U5335 (N_5335,N_5227,N_5218);
nor U5336 (N_5336,N_5210,N_5237);
and U5337 (N_5337,N_5235,N_5128);
xor U5338 (N_5338,N_5148,N_5180);
and U5339 (N_5339,N_5177,N_5154);
or U5340 (N_5340,N_5143,N_5149);
and U5341 (N_5341,N_5240,N_5193);
and U5342 (N_5342,N_5180,N_5221);
or U5343 (N_5343,N_5132,N_5171);
and U5344 (N_5344,N_5158,N_5183);
xnor U5345 (N_5345,N_5176,N_5209);
and U5346 (N_5346,N_5191,N_5165);
xnor U5347 (N_5347,N_5213,N_5196);
nor U5348 (N_5348,N_5186,N_5203);
nand U5349 (N_5349,N_5169,N_5204);
nand U5350 (N_5350,N_5205,N_5191);
xor U5351 (N_5351,N_5152,N_5182);
nand U5352 (N_5352,N_5142,N_5239);
nor U5353 (N_5353,N_5128,N_5145);
nor U5354 (N_5354,N_5222,N_5179);
nand U5355 (N_5355,N_5210,N_5140);
nand U5356 (N_5356,N_5202,N_5178);
nor U5357 (N_5357,N_5202,N_5221);
nand U5358 (N_5358,N_5159,N_5179);
and U5359 (N_5359,N_5204,N_5239);
and U5360 (N_5360,N_5181,N_5139);
or U5361 (N_5361,N_5211,N_5231);
nor U5362 (N_5362,N_5133,N_5154);
nor U5363 (N_5363,N_5203,N_5153);
nand U5364 (N_5364,N_5231,N_5195);
and U5365 (N_5365,N_5128,N_5240);
nor U5366 (N_5366,N_5238,N_5224);
and U5367 (N_5367,N_5235,N_5237);
nor U5368 (N_5368,N_5205,N_5230);
or U5369 (N_5369,N_5169,N_5187);
xnor U5370 (N_5370,N_5207,N_5241);
xnor U5371 (N_5371,N_5229,N_5175);
or U5372 (N_5372,N_5191,N_5181);
and U5373 (N_5373,N_5189,N_5175);
xor U5374 (N_5374,N_5183,N_5221);
xor U5375 (N_5375,N_5303,N_5270);
or U5376 (N_5376,N_5284,N_5291);
or U5377 (N_5377,N_5344,N_5302);
nor U5378 (N_5378,N_5252,N_5363);
nand U5379 (N_5379,N_5317,N_5359);
and U5380 (N_5380,N_5339,N_5301);
or U5381 (N_5381,N_5258,N_5282);
nand U5382 (N_5382,N_5260,N_5369);
and U5383 (N_5383,N_5274,N_5316);
and U5384 (N_5384,N_5309,N_5355);
nor U5385 (N_5385,N_5275,N_5279);
xor U5386 (N_5386,N_5334,N_5333);
or U5387 (N_5387,N_5314,N_5372);
nor U5388 (N_5388,N_5269,N_5323);
nor U5389 (N_5389,N_5352,N_5288);
nor U5390 (N_5390,N_5304,N_5261);
or U5391 (N_5391,N_5307,N_5330);
or U5392 (N_5392,N_5338,N_5366);
nor U5393 (N_5393,N_5370,N_5364);
and U5394 (N_5394,N_5285,N_5297);
and U5395 (N_5395,N_5340,N_5310);
or U5396 (N_5396,N_5327,N_5328);
nor U5397 (N_5397,N_5337,N_5273);
nor U5398 (N_5398,N_5374,N_5313);
nor U5399 (N_5399,N_5335,N_5332);
xnor U5400 (N_5400,N_5259,N_5349);
or U5401 (N_5401,N_5351,N_5371);
xnor U5402 (N_5402,N_5287,N_5250);
nor U5403 (N_5403,N_5368,N_5253);
nand U5404 (N_5404,N_5357,N_5331);
and U5405 (N_5405,N_5283,N_5295);
xnor U5406 (N_5406,N_5360,N_5311);
or U5407 (N_5407,N_5315,N_5348);
nor U5408 (N_5408,N_5264,N_5256);
xor U5409 (N_5409,N_5280,N_5353);
nor U5410 (N_5410,N_5361,N_5277);
xnor U5411 (N_5411,N_5267,N_5346);
nand U5412 (N_5412,N_5362,N_5324);
and U5413 (N_5413,N_5254,N_5300);
nand U5414 (N_5414,N_5266,N_5354);
nor U5415 (N_5415,N_5341,N_5292);
and U5416 (N_5416,N_5320,N_5358);
xor U5417 (N_5417,N_5262,N_5306);
or U5418 (N_5418,N_5325,N_5281);
nand U5419 (N_5419,N_5276,N_5336);
and U5420 (N_5420,N_5293,N_5299);
xor U5421 (N_5421,N_5272,N_5290);
nand U5422 (N_5422,N_5318,N_5342);
nand U5423 (N_5423,N_5305,N_5294);
nand U5424 (N_5424,N_5286,N_5312);
or U5425 (N_5425,N_5319,N_5278);
and U5426 (N_5426,N_5321,N_5367);
and U5427 (N_5427,N_5257,N_5308);
and U5428 (N_5428,N_5356,N_5365);
nand U5429 (N_5429,N_5322,N_5255);
nand U5430 (N_5430,N_5263,N_5350);
xnor U5431 (N_5431,N_5347,N_5251);
and U5432 (N_5432,N_5345,N_5289);
nand U5433 (N_5433,N_5271,N_5329);
or U5434 (N_5434,N_5373,N_5343);
xor U5435 (N_5435,N_5268,N_5296);
nand U5436 (N_5436,N_5265,N_5326);
nand U5437 (N_5437,N_5298,N_5293);
xnor U5438 (N_5438,N_5257,N_5315);
nor U5439 (N_5439,N_5309,N_5274);
or U5440 (N_5440,N_5264,N_5255);
nand U5441 (N_5441,N_5317,N_5289);
nor U5442 (N_5442,N_5319,N_5306);
nand U5443 (N_5443,N_5308,N_5291);
and U5444 (N_5444,N_5369,N_5299);
and U5445 (N_5445,N_5279,N_5348);
xor U5446 (N_5446,N_5314,N_5266);
or U5447 (N_5447,N_5328,N_5264);
nor U5448 (N_5448,N_5286,N_5333);
nor U5449 (N_5449,N_5357,N_5365);
and U5450 (N_5450,N_5344,N_5351);
nor U5451 (N_5451,N_5263,N_5364);
xor U5452 (N_5452,N_5274,N_5357);
or U5453 (N_5453,N_5321,N_5299);
and U5454 (N_5454,N_5366,N_5265);
xnor U5455 (N_5455,N_5274,N_5338);
xor U5456 (N_5456,N_5337,N_5370);
nand U5457 (N_5457,N_5273,N_5250);
and U5458 (N_5458,N_5300,N_5332);
xor U5459 (N_5459,N_5366,N_5328);
and U5460 (N_5460,N_5323,N_5317);
nand U5461 (N_5461,N_5276,N_5356);
nand U5462 (N_5462,N_5327,N_5346);
and U5463 (N_5463,N_5287,N_5264);
xnor U5464 (N_5464,N_5334,N_5357);
nor U5465 (N_5465,N_5325,N_5330);
or U5466 (N_5466,N_5278,N_5373);
and U5467 (N_5467,N_5365,N_5362);
nor U5468 (N_5468,N_5258,N_5259);
or U5469 (N_5469,N_5319,N_5347);
or U5470 (N_5470,N_5344,N_5309);
or U5471 (N_5471,N_5363,N_5361);
nand U5472 (N_5472,N_5316,N_5298);
and U5473 (N_5473,N_5256,N_5266);
nor U5474 (N_5474,N_5259,N_5363);
nor U5475 (N_5475,N_5257,N_5373);
or U5476 (N_5476,N_5300,N_5275);
nand U5477 (N_5477,N_5308,N_5320);
or U5478 (N_5478,N_5288,N_5322);
nand U5479 (N_5479,N_5277,N_5307);
xor U5480 (N_5480,N_5365,N_5264);
and U5481 (N_5481,N_5356,N_5295);
or U5482 (N_5482,N_5324,N_5250);
or U5483 (N_5483,N_5330,N_5303);
or U5484 (N_5484,N_5296,N_5357);
nand U5485 (N_5485,N_5275,N_5362);
xor U5486 (N_5486,N_5357,N_5366);
nand U5487 (N_5487,N_5273,N_5306);
nand U5488 (N_5488,N_5266,N_5352);
and U5489 (N_5489,N_5316,N_5277);
xor U5490 (N_5490,N_5316,N_5292);
nor U5491 (N_5491,N_5256,N_5325);
or U5492 (N_5492,N_5292,N_5333);
xnor U5493 (N_5493,N_5304,N_5299);
and U5494 (N_5494,N_5372,N_5269);
nor U5495 (N_5495,N_5359,N_5354);
or U5496 (N_5496,N_5274,N_5337);
xnor U5497 (N_5497,N_5312,N_5372);
xnor U5498 (N_5498,N_5313,N_5343);
xnor U5499 (N_5499,N_5297,N_5251);
xor U5500 (N_5500,N_5428,N_5420);
xnor U5501 (N_5501,N_5485,N_5459);
nand U5502 (N_5502,N_5449,N_5457);
and U5503 (N_5503,N_5477,N_5376);
or U5504 (N_5504,N_5495,N_5433);
nand U5505 (N_5505,N_5389,N_5481);
xnor U5506 (N_5506,N_5473,N_5474);
xor U5507 (N_5507,N_5483,N_5465);
and U5508 (N_5508,N_5448,N_5498);
or U5509 (N_5509,N_5416,N_5445);
or U5510 (N_5510,N_5400,N_5430);
xor U5511 (N_5511,N_5440,N_5419);
or U5512 (N_5512,N_5493,N_5476);
xor U5513 (N_5513,N_5432,N_5393);
xor U5514 (N_5514,N_5480,N_5439);
nand U5515 (N_5515,N_5409,N_5499);
nor U5516 (N_5516,N_5414,N_5461);
and U5517 (N_5517,N_5404,N_5438);
and U5518 (N_5518,N_5383,N_5434);
xor U5519 (N_5519,N_5444,N_5381);
and U5520 (N_5520,N_5468,N_5467);
nor U5521 (N_5521,N_5469,N_5379);
nand U5522 (N_5522,N_5472,N_5463);
and U5523 (N_5523,N_5447,N_5446);
or U5524 (N_5524,N_5391,N_5489);
nand U5525 (N_5525,N_5421,N_5406);
and U5526 (N_5526,N_5410,N_5494);
or U5527 (N_5527,N_5375,N_5385);
xnor U5528 (N_5528,N_5442,N_5423);
nor U5529 (N_5529,N_5466,N_5488);
nor U5530 (N_5530,N_5425,N_5491);
and U5531 (N_5531,N_5453,N_5396);
xor U5532 (N_5532,N_5386,N_5412);
xor U5533 (N_5533,N_5487,N_5486);
xnor U5534 (N_5534,N_5462,N_5451);
nand U5535 (N_5535,N_5417,N_5454);
or U5536 (N_5536,N_5455,N_5378);
and U5537 (N_5537,N_5443,N_5395);
or U5538 (N_5538,N_5398,N_5464);
nand U5539 (N_5539,N_5380,N_5415);
nor U5540 (N_5540,N_5418,N_5456);
or U5541 (N_5541,N_5413,N_5490);
or U5542 (N_5542,N_5422,N_5424);
or U5543 (N_5543,N_5479,N_5387);
or U5544 (N_5544,N_5496,N_5377);
nor U5545 (N_5545,N_5401,N_5458);
and U5546 (N_5546,N_5460,N_5407);
and U5547 (N_5547,N_5482,N_5452);
and U5548 (N_5548,N_5397,N_5478);
nor U5549 (N_5549,N_5475,N_5437);
nand U5550 (N_5550,N_5384,N_5399);
and U5551 (N_5551,N_5471,N_5450);
nor U5552 (N_5552,N_5470,N_5441);
and U5553 (N_5553,N_5435,N_5382);
or U5554 (N_5554,N_5484,N_5390);
or U5555 (N_5555,N_5492,N_5411);
nor U5556 (N_5556,N_5402,N_5394);
nor U5557 (N_5557,N_5431,N_5405);
or U5558 (N_5558,N_5388,N_5426);
xnor U5559 (N_5559,N_5429,N_5392);
nor U5560 (N_5560,N_5408,N_5497);
nor U5561 (N_5561,N_5427,N_5403);
and U5562 (N_5562,N_5436,N_5460);
or U5563 (N_5563,N_5424,N_5381);
and U5564 (N_5564,N_5470,N_5473);
or U5565 (N_5565,N_5380,N_5498);
nor U5566 (N_5566,N_5419,N_5436);
and U5567 (N_5567,N_5375,N_5456);
xnor U5568 (N_5568,N_5391,N_5496);
xor U5569 (N_5569,N_5457,N_5425);
nor U5570 (N_5570,N_5382,N_5394);
and U5571 (N_5571,N_5440,N_5411);
and U5572 (N_5572,N_5482,N_5440);
and U5573 (N_5573,N_5432,N_5487);
nor U5574 (N_5574,N_5410,N_5445);
xnor U5575 (N_5575,N_5415,N_5408);
nor U5576 (N_5576,N_5460,N_5423);
and U5577 (N_5577,N_5494,N_5481);
and U5578 (N_5578,N_5495,N_5496);
xnor U5579 (N_5579,N_5421,N_5423);
xnor U5580 (N_5580,N_5494,N_5439);
or U5581 (N_5581,N_5448,N_5475);
and U5582 (N_5582,N_5406,N_5436);
xnor U5583 (N_5583,N_5446,N_5379);
and U5584 (N_5584,N_5476,N_5416);
nand U5585 (N_5585,N_5462,N_5485);
xnor U5586 (N_5586,N_5486,N_5489);
and U5587 (N_5587,N_5439,N_5420);
or U5588 (N_5588,N_5389,N_5391);
nor U5589 (N_5589,N_5441,N_5476);
nand U5590 (N_5590,N_5431,N_5481);
nand U5591 (N_5591,N_5466,N_5486);
or U5592 (N_5592,N_5427,N_5447);
or U5593 (N_5593,N_5424,N_5404);
or U5594 (N_5594,N_5460,N_5440);
nand U5595 (N_5595,N_5478,N_5434);
xnor U5596 (N_5596,N_5407,N_5429);
and U5597 (N_5597,N_5481,N_5474);
or U5598 (N_5598,N_5459,N_5476);
or U5599 (N_5599,N_5468,N_5421);
xor U5600 (N_5600,N_5412,N_5488);
nor U5601 (N_5601,N_5414,N_5389);
nand U5602 (N_5602,N_5414,N_5427);
nor U5603 (N_5603,N_5490,N_5466);
xor U5604 (N_5604,N_5400,N_5442);
or U5605 (N_5605,N_5377,N_5456);
xnor U5606 (N_5606,N_5409,N_5420);
or U5607 (N_5607,N_5416,N_5422);
xor U5608 (N_5608,N_5451,N_5426);
nor U5609 (N_5609,N_5461,N_5476);
and U5610 (N_5610,N_5395,N_5393);
xor U5611 (N_5611,N_5420,N_5462);
and U5612 (N_5612,N_5389,N_5403);
and U5613 (N_5613,N_5375,N_5430);
and U5614 (N_5614,N_5489,N_5430);
or U5615 (N_5615,N_5447,N_5425);
and U5616 (N_5616,N_5397,N_5427);
nand U5617 (N_5617,N_5390,N_5406);
and U5618 (N_5618,N_5467,N_5483);
and U5619 (N_5619,N_5390,N_5442);
nand U5620 (N_5620,N_5400,N_5481);
nand U5621 (N_5621,N_5456,N_5469);
and U5622 (N_5622,N_5474,N_5466);
nor U5623 (N_5623,N_5393,N_5383);
xor U5624 (N_5624,N_5433,N_5383);
xor U5625 (N_5625,N_5591,N_5619);
nor U5626 (N_5626,N_5560,N_5509);
nand U5627 (N_5627,N_5511,N_5578);
xor U5628 (N_5628,N_5530,N_5592);
xnor U5629 (N_5629,N_5519,N_5501);
or U5630 (N_5630,N_5609,N_5512);
nand U5631 (N_5631,N_5617,N_5540);
and U5632 (N_5632,N_5620,N_5614);
xor U5633 (N_5633,N_5582,N_5577);
xor U5634 (N_5634,N_5550,N_5599);
nand U5635 (N_5635,N_5600,N_5587);
xor U5636 (N_5636,N_5537,N_5580);
xor U5637 (N_5637,N_5543,N_5548);
or U5638 (N_5638,N_5613,N_5558);
and U5639 (N_5639,N_5597,N_5534);
xnor U5640 (N_5640,N_5552,N_5621);
and U5641 (N_5641,N_5536,N_5611);
xnor U5642 (N_5642,N_5615,N_5573);
xnor U5643 (N_5643,N_5516,N_5583);
nand U5644 (N_5644,N_5612,N_5546);
nand U5645 (N_5645,N_5527,N_5595);
nand U5646 (N_5646,N_5571,N_5603);
nor U5647 (N_5647,N_5594,N_5596);
and U5648 (N_5648,N_5556,N_5508);
and U5649 (N_5649,N_5525,N_5576);
nand U5650 (N_5650,N_5601,N_5542);
nand U5651 (N_5651,N_5557,N_5555);
or U5652 (N_5652,N_5507,N_5549);
xor U5653 (N_5653,N_5514,N_5570);
xor U5654 (N_5654,N_5526,N_5579);
or U5655 (N_5655,N_5503,N_5544);
or U5656 (N_5656,N_5623,N_5554);
or U5657 (N_5657,N_5553,N_5510);
nand U5658 (N_5658,N_5585,N_5622);
xnor U5659 (N_5659,N_5605,N_5547);
nand U5660 (N_5660,N_5520,N_5567);
and U5661 (N_5661,N_5610,N_5535);
and U5662 (N_5662,N_5517,N_5589);
and U5663 (N_5663,N_5564,N_5523);
nand U5664 (N_5664,N_5531,N_5565);
and U5665 (N_5665,N_5541,N_5513);
xor U5666 (N_5666,N_5581,N_5604);
and U5667 (N_5667,N_5521,N_5588);
nor U5668 (N_5668,N_5598,N_5568);
and U5669 (N_5669,N_5533,N_5545);
and U5670 (N_5670,N_5559,N_5569);
and U5671 (N_5671,N_5572,N_5528);
nor U5672 (N_5672,N_5574,N_5562);
nor U5673 (N_5673,N_5616,N_5593);
xor U5674 (N_5674,N_5539,N_5590);
nor U5675 (N_5675,N_5624,N_5505);
nand U5676 (N_5676,N_5575,N_5506);
nand U5677 (N_5677,N_5524,N_5518);
nand U5678 (N_5678,N_5563,N_5566);
nor U5679 (N_5679,N_5504,N_5586);
or U5680 (N_5680,N_5607,N_5515);
nand U5681 (N_5681,N_5606,N_5500);
nand U5682 (N_5682,N_5551,N_5602);
xnor U5683 (N_5683,N_5561,N_5608);
nor U5684 (N_5684,N_5618,N_5502);
and U5685 (N_5685,N_5522,N_5538);
nand U5686 (N_5686,N_5584,N_5529);
nand U5687 (N_5687,N_5532,N_5511);
or U5688 (N_5688,N_5611,N_5526);
nor U5689 (N_5689,N_5510,N_5511);
and U5690 (N_5690,N_5607,N_5597);
nand U5691 (N_5691,N_5558,N_5539);
nand U5692 (N_5692,N_5614,N_5599);
and U5693 (N_5693,N_5574,N_5556);
and U5694 (N_5694,N_5580,N_5500);
and U5695 (N_5695,N_5582,N_5502);
nand U5696 (N_5696,N_5622,N_5588);
nand U5697 (N_5697,N_5520,N_5580);
nor U5698 (N_5698,N_5512,N_5559);
xnor U5699 (N_5699,N_5533,N_5603);
xnor U5700 (N_5700,N_5540,N_5512);
and U5701 (N_5701,N_5591,N_5577);
or U5702 (N_5702,N_5503,N_5549);
xor U5703 (N_5703,N_5611,N_5514);
and U5704 (N_5704,N_5537,N_5591);
nand U5705 (N_5705,N_5562,N_5505);
nor U5706 (N_5706,N_5504,N_5549);
nor U5707 (N_5707,N_5516,N_5569);
and U5708 (N_5708,N_5602,N_5591);
and U5709 (N_5709,N_5593,N_5505);
and U5710 (N_5710,N_5512,N_5508);
or U5711 (N_5711,N_5511,N_5601);
and U5712 (N_5712,N_5507,N_5517);
nor U5713 (N_5713,N_5571,N_5618);
or U5714 (N_5714,N_5613,N_5526);
and U5715 (N_5715,N_5556,N_5612);
nor U5716 (N_5716,N_5605,N_5528);
nor U5717 (N_5717,N_5594,N_5534);
and U5718 (N_5718,N_5504,N_5607);
or U5719 (N_5719,N_5595,N_5594);
or U5720 (N_5720,N_5531,N_5560);
nand U5721 (N_5721,N_5604,N_5572);
xor U5722 (N_5722,N_5548,N_5542);
nand U5723 (N_5723,N_5521,N_5518);
or U5724 (N_5724,N_5557,N_5613);
nor U5725 (N_5725,N_5593,N_5512);
nand U5726 (N_5726,N_5551,N_5558);
nand U5727 (N_5727,N_5531,N_5587);
or U5728 (N_5728,N_5523,N_5542);
xor U5729 (N_5729,N_5571,N_5509);
nor U5730 (N_5730,N_5527,N_5608);
or U5731 (N_5731,N_5504,N_5581);
or U5732 (N_5732,N_5544,N_5574);
and U5733 (N_5733,N_5512,N_5584);
xnor U5734 (N_5734,N_5514,N_5540);
nor U5735 (N_5735,N_5525,N_5506);
or U5736 (N_5736,N_5522,N_5620);
xor U5737 (N_5737,N_5548,N_5560);
xnor U5738 (N_5738,N_5504,N_5617);
or U5739 (N_5739,N_5564,N_5541);
nor U5740 (N_5740,N_5509,N_5565);
and U5741 (N_5741,N_5577,N_5588);
xnor U5742 (N_5742,N_5620,N_5624);
xnor U5743 (N_5743,N_5530,N_5600);
xnor U5744 (N_5744,N_5513,N_5579);
xor U5745 (N_5745,N_5602,N_5542);
and U5746 (N_5746,N_5587,N_5591);
and U5747 (N_5747,N_5536,N_5554);
nor U5748 (N_5748,N_5612,N_5565);
and U5749 (N_5749,N_5507,N_5513);
or U5750 (N_5750,N_5728,N_5625);
nand U5751 (N_5751,N_5670,N_5749);
xnor U5752 (N_5752,N_5705,N_5642);
nor U5753 (N_5753,N_5736,N_5686);
nand U5754 (N_5754,N_5661,N_5746);
xor U5755 (N_5755,N_5710,N_5687);
or U5756 (N_5756,N_5726,N_5641);
or U5757 (N_5757,N_5692,N_5640);
nand U5758 (N_5758,N_5743,N_5645);
xor U5759 (N_5759,N_5740,N_5682);
nand U5760 (N_5760,N_5721,N_5694);
and U5761 (N_5761,N_5724,N_5725);
xnor U5762 (N_5762,N_5685,N_5660);
or U5763 (N_5763,N_5739,N_5708);
and U5764 (N_5764,N_5693,N_5709);
nor U5765 (N_5765,N_5690,N_5712);
nand U5766 (N_5766,N_5632,N_5679);
nand U5767 (N_5767,N_5695,N_5733);
nor U5768 (N_5768,N_5648,N_5707);
xnor U5769 (N_5769,N_5706,N_5681);
and U5770 (N_5770,N_5714,N_5701);
xor U5771 (N_5771,N_5629,N_5664);
or U5772 (N_5772,N_5689,N_5672);
and U5773 (N_5773,N_5631,N_5634);
and U5774 (N_5774,N_5730,N_5633);
xnor U5775 (N_5775,N_5678,N_5723);
xnor U5776 (N_5776,N_5718,N_5744);
nand U5777 (N_5777,N_5674,N_5655);
nand U5778 (N_5778,N_5650,N_5643);
nor U5779 (N_5779,N_5627,N_5704);
xor U5780 (N_5780,N_5666,N_5684);
or U5781 (N_5781,N_5741,N_5702);
and U5782 (N_5782,N_5656,N_5665);
nand U5783 (N_5783,N_5698,N_5683);
nor U5784 (N_5784,N_5716,N_5748);
xor U5785 (N_5785,N_5638,N_5699);
xnor U5786 (N_5786,N_5659,N_5646);
and U5787 (N_5787,N_5667,N_5700);
xor U5788 (N_5788,N_5658,N_5668);
or U5789 (N_5789,N_5717,N_5688);
or U5790 (N_5790,N_5735,N_5680);
xnor U5791 (N_5791,N_5647,N_5731);
xor U5792 (N_5792,N_5654,N_5727);
nand U5793 (N_5793,N_5734,N_5677);
nor U5794 (N_5794,N_5711,N_5671);
nor U5795 (N_5795,N_5732,N_5696);
and U5796 (N_5796,N_5738,N_5676);
and U5797 (N_5797,N_5652,N_5628);
nand U5798 (N_5798,N_5657,N_5747);
nand U5799 (N_5799,N_5722,N_5745);
and U5800 (N_5800,N_5644,N_5663);
nand U5801 (N_5801,N_5649,N_5697);
nand U5802 (N_5802,N_5703,N_5651);
nand U5803 (N_5803,N_5729,N_5639);
nor U5804 (N_5804,N_5713,N_5662);
xnor U5805 (N_5805,N_5635,N_5715);
xor U5806 (N_5806,N_5720,N_5742);
and U5807 (N_5807,N_5719,N_5737);
or U5808 (N_5808,N_5669,N_5691);
xnor U5809 (N_5809,N_5626,N_5637);
xor U5810 (N_5810,N_5673,N_5636);
and U5811 (N_5811,N_5675,N_5630);
or U5812 (N_5812,N_5653,N_5697);
xor U5813 (N_5813,N_5659,N_5708);
nand U5814 (N_5814,N_5698,N_5695);
xor U5815 (N_5815,N_5663,N_5704);
or U5816 (N_5816,N_5692,N_5636);
nand U5817 (N_5817,N_5666,N_5664);
and U5818 (N_5818,N_5679,N_5744);
nor U5819 (N_5819,N_5712,N_5667);
nand U5820 (N_5820,N_5700,N_5730);
and U5821 (N_5821,N_5678,N_5692);
and U5822 (N_5822,N_5680,N_5674);
xor U5823 (N_5823,N_5686,N_5747);
or U5824 (N_5824,N_5735,N_5700);
xor U5825 (N_5825,N_5705,N_5743);
and U5826 (N_5826,N_5725,N_5712);
xnor U5827 (N_5827,N_5731,N_5667);
nand U5828 (N_5828,N_5649,N_5646);
xor U5829 (N_5829,N_5713,N_5741);
and U5830 (N_5830,N_5689,N_5738);
xor U5831 (N_5831,N_5736,N_5669);
nand U5832 (N_5832,N_5700,N_5744);
nor U5833 (N_5833,N_5666,N_5668);
nor U5834 (N_5834,N_5700,N_5734);
and U5835 (N_5835,N_5733,N_5746);
or U5836 (N_5836,N_5659,N_5695);
or U5837 (N_5837,N_5725,N_5664);
or U5838 (N_5838,N_5628,N_5735);
xnor U5839 (N_5839,N_5640,N_5709);
nor U5840 (N_5840,N_5688,N_5712);
and U5841 (N_5841,N_5740,N_5667);
or U5842 (N_5842,N_5640,N_5701);
nor U5843 (N_5843,N_5625,N_5679);
or U5844 (N_5844,N_5713,N_5738);
nand U5845 (N_5845,N_5649,N_5679);
xnor U5846 (N_5846,N_5717,N_5708);
or U5847 (N_5847,N_5661,N_5652);
nand U5848 (N_5848,N_5627,N_5630);
xor U5849 (N_5849,N_5642,N_5692);
nor U5850 (N_5850,N_5699,N_5702);
and U5851 (N_5851,N_5663,N_5706);
or U5852 (N_5852,N_5737,N_5665);
or U5853 (N_5853,N_5737,N_5747);
and U5854 (N_5854,N_5659,N_5694);
or U5855 (N_5855,N_5667,N_5699);
nor U5856 (N_5856,N_5730,N_5644);
and U5857 (N_5857,N_5636,N_5664);
nor U5858 (N_5858,N_5678,N_5704);
nand U5859 (N_5859,N_5714,N_5657);
xor U5860 (N_5860,N_5677,N_5681);
nand U5861 (N_5861,N_5652,N_5707);
nand U5862 (N_5862,N_5728,N_5650);
and U5863 (N_5863,N_5728,N_5729);
nand U5864 (N_5864,N_5710,N_5628);
nor U5865 (N_5865,N_5684,N_5726);
xor U5866 (N_5866,N_5689,N_5647);
or U5867 (N_5867,N_5655,N_5736);
xnor U5868 (N_5868,N_5667,N_5702);
xnor U5869 (N_5869,N_5726,N_5693);
nor U5870 (N_5870,N_5670,N_5659);
and U5871 (N_5871,N_5670,N_5745);
nand U5872 (N_5872,N_5749,N_5698);
nand U5873 (N_5873,N_5714,N_5720);
nor U5874 (N_5874,N_5714,N_5682);
xnor U5875 (N_5875,N_5755,N_5801);
xnor U5876 (N_5876,N_5831,N_5842);
nand U5877 (N_5877,N_5791,N_5818);
xnor U5878 (N_5878,N_5870,N_5823);
and U5879 (N_5879,N_5798,N_5787);
xor U5880 (N_5880,N_5835,N_5789);
nor U5881 (N_5881,N_5825,N_5782);
nand U5882 (N_5882,N_5866,N_5804);
nand U5883 (N_5883,N_5802,N_5771);
nand U5884 (N_5884,N_5869,N_5872);
nand U5885 (N_5885,N_5873,N_5843);
xnor U5886 (N_5886,N_5847,N_5779);
xor U5887 (N_5887,N_5816,N_5809);
xor U5888 (N_5888,N_5751,N_5810);
nand U5889 (N_5889,N_5793,N_5833);
or U5890 (N_5890,N_5837,N_5851);
nand U5891 (N_5891,N_5777,N_5774);
nand U5892 (N_5892,N_5836,N_5838);
and U5893 (N_5893,N_5757,N_5813);
nor U5894 (N_5894,N_5859,N_5828);
nor U5895 (N_5895,N_5790,N_5753);
or U5896 (N_5896,N_5857,N_5849);
nor U5897 (N_5897,N_5780,N_5764);
or U5898 (N_5898,N_5766,N_5820);
nor U5899 (N_5899,N_5803,N_5811);
nor U5900 (N_5900,N_5846,N_5808);
xor U5901 (N_5901,N_5758,N_5750);
and U5902 (N_5902,N_5840,N_5867);
nor U5903 (N_5903,N_5827,N_5844);
xnor U5904 (N_5904,N_5776,N_5795);
nand U5905 (N_5905,N_5772,N_5863);
nand U5906 (N_5906,N_5819,N_5868);
and U5907 (N_5907,N_5762,N_5799);
or U5908 (N_5908,N_5845,N_5781);
nor U5909 (N_5909,N_5858,N_5770);
xnor U5910 (N_5910,N_5815,N_5822);
and U5911 (N_5911,N_5788,N_5761);
xnor U5912 (N_5912,N_5767,N_5853);
nand U5913 (N_5913,N_5850,N_5784);
nor U5914 (N_5914,N_5861,N_5814);
and U5915 (N_5915,N_5800,N_5864);
or U5916 (N_5916,N_5783,N_5865);
and U5917 (N_5917,N_5768,N_5778);
nor U5918 (N_5918,N_5769,N_5796);
nor U5919 (N_5919,N_5812,N_5830);
nor U5920 (N_5920,N_5860,N_5759);
nor U5921 (N_5921,N_5839,N_5785);
nand U5922 (N_5922,N_5832,N_5752);
nor U5923 (N_5923,N_5807,N_5806);
xor U5924 (N_5924,N_5874,N_5852);
or U5925 (N_5925,N_5854,N_5773);
nor U5926 (N_5926,N_5765,N_5824);
or U5927 (N_5927,N_5821,N_5805);
nor U5928 (N_5928,N_5826,N_5841);
and U5929 (N_5929,N_5754,N_5848);
and U5930 (N_5930,N_5862,N_5797);
nand U5931 (N_5931,N_5775,N_5786);
nand U5932 (N_5932,N_5760,N_5855);
or U5933 (N_5933,N_5794,N_5871);
nand U5934 (N_5934,N_5763,N_5856);
or U5935 (N_5935,N_5829,N_5834);
and U5936 (N_5936,N_5817,N_5792);
and U5937 (N_5937,N_5756,N_5830);
xor U5938 (N_5938,N_5814,N_5870);
nor U5939 (N_5939,N_5838,N_5830);
nand U5940 (N_5940,N_5752,N_5858);
or U5941 (N_5941,N_5843,N_5805);
nand U5942 (N_5942,N_5794,N_5785);
and U5943 (N_5943,N_5761,N_5844);
nor U5944 (N_5944,N_5832,N_5821);
nor U5945 (N_5945,N_5761,N_5838);
nor U5946 (N_5946,N_5775,N_5857);
nand U5947 (N_5947,N_5757,N_5864);
nand U5948 (N_5948,N_5831,N_5755);
xnor U5949 (N_5949,N_5808,N_5847);
xnor U5950 (N_5950,N_5776,N_5807);
xnor U5951 (N_5951,N_5751,N_5779);
nor U5952 (N_5952,N_5837,N_5768);
xor U5953 (N_5953,N_5829,N_5751);
or U5954 (N_5954,N_5835,N_5806);
nor U5955 (N_5955,N_5777,N_5766);
nor U5956 (N_5956,N_5824,N_5794);
xnor U5957 (N_5957,N_5800,N_5794);
nor U5958 (N_5958,N_5843,N_5844);
and U5959 (N_5959,N_5856,N_5788);
nor U5960 (N_5960,N_5866,N_5826);
nor U5961 (N_5961,N_5760,N_5788);
nand U5962 (N_5962,N_5871,N_5832);
nor U5963 (N_5963,N_5782,N_5762);
and U5964 (N_5964,N_5758,N_5769);
xnor U5965 (N_5965,N_5869,N_5826);
nand U5966 (N_5966,N_5860,N_5836);
and U5967 (N_5967,N_5835,N_5824);
or U5968 (N_5968,N_5829,N_5782);
xnor U5969 (N_5969,N_5783,N_5775);
nor U5970 (N_5970,N_5777,N_5759);
and U5971 (N_5971,N_5768,N_5751);
xor U5972 (N_5972,N_5827,N_5806);
nand U5973 (N_5973,N_5778,N_5783);
xnor U5974 (N_5974,N_5870,N_5802);
nor U5975 (N_5975,N_5753,N_5826);
xnor U5976 (N_5976,N_5806,N_5774);
nor U5977 (N_5977,N_5767,N_5832);
and U5978 (N_5978,N_5783,N_5769);
nand U5979 (N_5979,N_5818,N_5769);
xnor U5980 (N_5980,N_5839,N_5812);
nor U5981 (N_5981,N_5809,N_5871);
xor U5982 (N_5982,N_5845,N_5790);
xnor U5983 (N_5983,N_5870,N_5776);
or U5984 (N_5984,N_5797,N_5838);
and U5985 (N_5985,N_5828,N_5858);
xnor U5986 (N_5986,N_5796,N_5791);
nor U5987 (N_5987,N_5752,N_5853);
nand U5988 (N_5988,N_5831,N_5816);
nand U5989 (N_5989,N_5825,N_5862);
nand U5990 (N_5990,N_5841,N_5865);
and U5991 (N_5991,N_5835,N_5762);
nand U5992 (N_5992,N_5765,N_5802);
or U5993 (N_5993,N_5800,N_5792);
or U5994 (N_5994,N_5803,N_5857);
and U5995 (N_5995,N_5824,N_5761);
nand U5996 (N_5996,N_5791,N_5805);
or U5997 (N_5997,N_5762,N_5853);
and U5998 (N_5998,N_5784,N_5854);
nor U5999 (N_5999,N_5794,N_5802);
and U6000 (N_6000,N_5911,N_5965);
nor U6001 (N_6001,N_5990,N_5967);
nand U6002 (N_6002,N_5887,N_5986);
and U6003 (N_6003,N_5904,N_5975);
nand U6004 (N_6004,N_5999,N_5906);
xnor U6005 (N_6005,N_5993,N_5957);
and U6006 (N_6006,N_5976,N_5886);
nor U6007 (N_6007,N_5881,N_5956);
and U6008 (N_6008,N_5934,N_5893);
or U6009 (N_6009,N_5978,N_5878);
and U6010 (N_6010,N_5917,N_5876);
nand U6011 (N_6011,N_5949,N_5875);
nand U6012 (N_6012,N_5979,N_5924);
and U6013 (N_6013,N_5970,N_5931);
and U6014 (N_6014,N_5900,N_5929);
and U6015 (N_6015,N_5888,N_5884);
and U6016 (N_6016,N_5921,N_5960);
and U6017 (N_6017,N_5923,N_5895);
nand U6018 (N_6018,N_5963,N_5971);
nor U6019 (N_6019,N_5995,N_5938);
xor U6020 (N_6020,N_5985,N_5890);
nor U6021 (N_6021,N_5959,N_5901);
or U6022 (N_6022,N_5925,N_5977);
nor U6023 (N_6023,N_5943,N_5973);
nand U6024 (N_6024,N_5932,N_5937);
xnor U6025 (N_6025,N_5992,N_5915);
and U6026 (N_6026,N_5982,N_5951);
nor U6027 (N_6027,N_5958,N_5945);
nor U6028 (N_6028,N_5913,N_5946);
nor U6029 (N_6029,N_5998,N_5966);
xor U6030 (N_6030,N_5892,N_5983);
nand U6031 (N_6031,N_5972,N_5910);
nor U6032 (N_6032,N_5939,N_5920);
or U6033 (N_6033,N_5896,N_5882);
nand U6034 (N_6034,N_5914,N_5980);
or U6035 (N_6035,N_5961,N_5935);
nor U6036 (N_6036,N_5930,N_5974);
or U6037 (N_6037,N_5889,N_5950);
nor U6038 (N_6038,N_5996,N_5987);
nor U6039 (N_6039,N_5905,N_5964);
xnor U6040 (N_6040,N_5948,N_5912);
nor U6041 (N_6041,N_5955,N_5994);
nand U6042 (N_6042,N_5897,N_5879);
or U6043 (N_6043,N_5936,N_5940);
and U6044 (N_6044,N_5880,N_5933);
nand U6045 (N_6045,N_5907,N_5927);
and U6046 (N_6046,N_5922,N_5926);
or U6047 (N_6047,N_5899,N_5954);
and U6048 (N_6048,N_5953,N_5919);
xnor U6049 (N_6049,N_5942,N_5883);
nor U6050 (N_6050,N_5988,N_5903);
nand U6051 (N_6051,N_5928,N_5944);
nand U6052 (N_6052,N_5885,N_5894);
xor U6053 (N_6053,N_5952,N_5908);
and U6054 (N_6054,N_5909,N_5902);
and U6055 (N_6055,N_5991,N_5989);
xor U6056 (N_6056,N_5898,N_5981);
nand U6057 (N_6057,N_5969,N_5877);
or U6058 (N_6058,N_5968,N_5918);
or U6059 (N_6059,N_5997,N_5984);
nor U6060 (N_6060,N_5947,N_5941);
nor U6061 (N_6061,N_5891,N_5916);
or U6062 (N_6062,N_5962,N_5998);
or U6063 (N_6063,N_5998,N_5910);
or U6064 (N_6064,N_5955,N_5894);
and U6065 (N_6065,N_5886,N_5986);
xnor U6066 (N_6066,N_5961,N_5954);
nor U6067 (N_6067,N_5906,N_5908);
nand U6068 (N_6068,N_5927,N_5926);
or U6069 (N_6069,N_5899,N_5993);
and U6070 (N_6070,N_5968,N_5949);
xor U6071 (N_6071,N_5924,N_5943);
nor U6072 (N_6072,N_5899,N_5934);
xnor U6073 (N_6073,N_5954,N_5892);
and U6074 (N_6074,N_5986,N_5962);
xor U6075 (N_6075,N_5882,N_5914);
and U6076 (N_6076,N_5968,N_5888);
nand U6077 (N_6077,N_5994,N_5913);
xor U6078 (N_6078,N_5953,N_5913);
nand U6079 (N_6079,N_5961,N_5992);
and U6080 (N_6080,N_5947,N_5909);
xnor U6081 (N_6081,N_5878,N_5914);
nand U6082 (N_6082,N_5970,N_5999);
nand U6083 (N_6083,N_5978,N_5984);
nor U6084 (N_6084,N_5919,N_5917);
xor U6085 (N_6085,N_5962,N_5969);
nor U6086 (N_6086,N_5894,N_5891);
and U6087 (N_6087,N_5896,N_5936);
nor U6088 (N_6088,N_5980,N_5893);
and U6089 (N_6089,N_5927,N_5901);
xor U6090 (N_6090,N_5923,N_5986);
or U6091 (N_6091,N_5902,N_5955);
or U6092 (N_6092,N_5914,N_5915);
nand U6093 (N_6093,N_5933,N_5892);
xnor U6094 (N_6094,N_5897,N_5998);
or U6095 (N_6095,N_5888,N_5899);
nor U6096 (N_6096,N_5999,N_5958);
nor U6097 (N_6097,N_5992,N_5925);
xor U6098 (N_6098,N_5949,N_5967);
and U6099 (N_6099,N_5968,N_5905);
nor U6100 (N_6100,N_5929,N_5980);
and U6101 (N_6101,N_5954,N_5881);
nor U6102 (N_6102,N_5922,N_5990);
or U6103 (N_6103,N_5941,N_5952);
or U6104 (N_6104,N_5894,N_5931);
or U6105 (N_6105,N_5962,N_5922);
or U6106 (N_6106,N_5999,N_5927);
nand U6107 (N_6107,N_5892,N_5926);
xor U6108 (N_6108,N_5896,N_5897);
xor U6109 (N_6109,N_5907,N_5899);
xor U6110 (N_6110,N_5886,N_5965);
nand U6111 (N_6111,N_5964,N_5934);
nor U6112 (N_6112,N_5903,N_5992);
nand U6113 (N_6113,N_5913,N_5956);
or U6114 (N_6114,N_5875,N_5927);
xor U6115 (N_6115,N_5875,N_5915);
and U6116 (N_6116,N_5968,N_5939);
or U6117 (N_6117,N_5915,N_5966);
and U6118 (N_6118,N_5912,N_5876);
nand U6119 (N_6119,N_5936,N_5911);
xnor U6120 (N_6120,N_5956,N_5906);
and U6121 (N_6121,N_5957,N_5939);
nand U6122 (N_6122,N_5970,N_5909);
or U6123 (N_6123,N_5940,N_5880);
xnor U6124 (N_6124,N_5967,N_5928);
and U6125 (N_6125,N_6050,N_6124);
xnor U6126 (N_6126,N_6087,N_6116);
nand U6127 (N_6127,N_6035,N_6048);
nor U6128 (N_6128,N_6106,N_6043);
nand U6129 (N_6129,N_6041,N_6097);
and U6130 (N_6130,N_6021,N_6069);
xor U6131 (N_6131,N_6107,N_6037);
nor U6132 (N_6132,N_6018,N_6091);
or U6133 (N_6133,N_6066,N_6044);
xor U6134 (N_6134,N_6098,N_6019);
nor U6135 (N_6135,N_6002,N_6024);
and U6136 (N_6136,N_6084,N_6022);
or U6137 (N_6137,N_6046,N_6023);
nor U6138 (N_6138,N_6072,N_6061);
xor U6139 (N_6139,N_6085,N_6003);
xnor U6140 (N_6140,N_6082,N_6052);
or U6141 (N_6141,N_6014,N_6123);
or U6142 (N_6142,N_6103,N_6067);
nor U6143 (N_6143,N_6031,N_6054);
nand U6144 (N_6144,N_6032,N_6068);
and U6145 (N_6145,N_6039,N_6077);
and U6146 (N_6146,N_6001,N_6029);
nor U6147 (N_6147,N_6057,N_6114);
or U6148 (N_6148,N_6100,N_6120);
nand U6149 (N_6149,N_6081,N_6034);
or U6150 (N_6150,N_6010,N_6015);
and U6151 (N_6151,N_6013,N_6033);
nor U6152 (N_6152,N_6083,N_6086);
nor U6153 (N_6153,N_6025,N_6093);
xor U6154 (N_6154,N_6005,N_6062);
xnor U6155 (N_6155,N_6102,N_6076);
or U6156 (N_6156,N_6101,N_6070);
and U6157 (N_6157,N_6099,N_6027);
and U6158 (N_6158,N_6079,N_6105);
or U6159 (N_6159,N_6008,N_6051);
nand U6160 (N_6160,N_6089,N_6115);
and U6161 (N_6161,N_6080,N_6007);
and U6162 (N_6162,N_6119,N_6055);
and U6163 (N_6163,N_6121,N_6017);
nand U6164 (N_6164,N_6110,N_6112);
and U6165 (N_6165,N_6004,N_6096);
and U6166 (N_6166,N_6078,N_6012);
and U6167 (N_6167,N_6006,N_6026);
and U6168 (N_6168,N_6108,N_6056);
or U6169 (N_6169,N_6047,N_6040);
xor U6170 (N_6170,N_6020,N_6117);
and U6171 (N_6171,N_6088,N_6073);
and U6172 (N_6172,N_6038,N_6049);
xor U6173 (N_6173,N_6028,N_6113);
and U6174 (N_6174,N_6074,N_6111);
nor U6175 (N_6175,N_6016,N_6065);
xor U6176 (N_6176,N_6058,N_6042);
xnor U6177 (N_6177,N_6064,N_6118);
or U6178 (N_6178,N_6122,N_6075);
or U6179 (N_6179,N_6063,N_6090);
or U6180 (N_6180,N_6094,N_6104);
and U6181 (N_6181,N_6000,N_6009);
nor U6182 (N_6182,N_6011,N_6053);
and U6183 (N_6183,N_6092,N_6109);
and U6184 (N_6184,N_6045,N_6036);
nand U6185 (N_6185,N_6059,N_6060);
nor U6186 (N_6186,N_6030,N_6071);
or U6187 (N_6187,N_6095,N_6109);
and U6188 (N_6188,N_6017,N_6056);
nor U6189 (N_6189,N_6056,N_6105);
or U6190 (N_6190,N_6032,N_6063);
nor U6191 (N_6191,N_6083,N_6088);
and U6192 (N_6192,N_6048,N_6005);
or U6193 (N_6193,N_6009,N_6090);
nand U6194 (N_6194,N_6109,N_6045);
or U6195 (N_6195,N_6072,N_6092);
or U6196 (N_6196,N_6056,N_6071);
xnor U6197 (N_6197,N_6090,N_6029);
or U6198 (N_6198,N_6038,N_6022);
nor U6199 (N_6199,N_6087,N_6048);
and U6200 (N_6200,N_6089,N_6071);
nand U6201 (N_6201,N_6045,N_6059);
and U6202 (N_6202,N_6078,N_6025);
and U6203 (N_6203,N_6066,N_6092);
and U6204 (N_6204,N_6067,N_6007);
or U6205 (N_6205,N_6069,N_6123);
and U6206 (N_6206,N_6049,N_6066);
nor U6207 (N_6207,N_6067,N_6016);
and U6208 (N_6208,N_6119,N_6072);
and U6209 (N_6209,N_6062,N_6000);
and U6210 (N_6210,N_6039,N_6033);
and U6211 (N_6211,N_6036,N_6000);
nand U6212 (N_6212,N_6091,N_6114);
xnor U6213 (N_6213,N_6099,N_6102);
or U6214 (N_6214,N_6055,N_6104);
nand U6215 (N_6215,N_6035,N_6084);
nand U6216 (N_6216,N_6033,N_6093);
xnor U6217 (N_6217,N_6023,N_6000);
and U6218 (N_6218,N_6018,N_6021);
xnor U6219 (N_6219,N_6076,N_6117);
nand U6220 (N_6220,N_6058,N_6103);
and U6221 (N_6221,N_6076,N_6052);
and U6222 (N_6222,N_6070,N_6066);
xnor U6223 (N_6223,N_6105,N_6046);
or U6224 (N_6224,N_6024,N_6029);
or U6225 (N_6225,N_6111,N_6116);
nor U6226 (N_6226,N_6056,N_6061);
nand U6227 (N_6227,N_6029,N_6048);
nand U6228 (N_6228,N_6068,N_6058);
nand U6229 (N_6229,N_6067,N_6008);
nand U6230 (N_6230,N_6003,N_6014);
nand U6231 (N_6231,N_6065,N_6050);
nor U6232 (N_6232,N_6053,N_6100);
xnor U6233 (N_6233,N_6059,N_6095);
nand U6234 (N_6234,N_6084,N_6082);
and U6235 (N_6235,N_6113,N_6065);
nand U6236 (N_6236,N_6080,N_6119);
and U6237 (N_6237,N_6010,N_6056);
and U6238 (N_6238,N_6084,N_6002);
nor U6239 (N_6239,N_6083,N_6050);
nor U6240 (N_6240,N_6060,N_6095);
and U6241 (N_6241,N_6086,N_6006);
or U6242 (N_6242,N_6059,N_6006);
xnor U6243 (N_6243,N_6120,N_6048);
or U6244 (N_6244,N_6122,N_6063);
xor U6245 (N_6245,N_6008,N_6019);
nand U6246 (N_6246,N_6052,N_6054);
nor U6247 (N_6247,N_6086,N_6104);
nor U6248 (N_6248,N_6117,N_6105);
nand U6249 (N_6249,N_6068,N_6094);
and U6250 (N_6250,N_6234,N_6231);
or U6251 (N_6251,N_6228,N_6232);
and U6252 (N_6252,N_6140,N_6248);
and U6253 (N_6253,N_6155,N_6213);
and U6254 (N_6254,N_6217,N_6147);
and U6255 (N_6255,N_6163,N_6190);
xor U6256 (N_6256,N_6168,N_6177);
and U6257 (N_6257,N_6199,N_6161);
and U6258 (N_6258,N_6186,N_6221);
nand U6259 (N_6259,N_6200,N_6205);
and U6260 (N_6260,N_6125,N_6194);
nor U6261 (N_6261,N_6238,N_6152);
and U6262 (N_6262,N_6160,N_6171);
or U6263 (N_6263,N_6178,N_6151);
nor U6264 (N_6264,N_6153,N_6249);
or U6265 (N_6265,N_6220,N_6214);
xor U6266 (N_6266,N_6130,N_6240);
xor U6267 (N_6267,N_6196,N_6154);
nand U6268 (N_6268,N_6237,N_6129);
xnor U6269 (N_6269,N_6243,N_6165);
and U6270 (N_6270,N_6224,N_6164);
or U6271 (N_6271,N_6150,N_6172);
or U6272 (N_6272,N_6158,N_6169);
nor U6273 (N_6273,N_6184,N_6204);
or U6274 (N_6274,N_6219,N_6187);
or U6275 (N_6275,N_6195,N_6182);
nand U6276 (N_6276,N_6247,N_6183);
nand U6277 (N_6277,N_6162,N_6142);
or U6278 (N_6278,N_6226,N_6156);
nor U6279 (N_6279,N_6180,N_6201);
xnor U6280 (N_6280,N_6227,N_6235);
and U6281 (N_6281,N_6207,N_6145);
nand U6282 (N_6282,N_6212,N_6135);
nand U6283 (N_6283,N_6244,N_6136);
or U6284 (N_6284,N_6157,N_6132);
nand U6285 (N_6285,N_6167,N_6185);
or U6286 (N_6286,N_6233,N_6126);
and U6287 (N_6287,N_6188,N_6192);
or U6288 (N_6288,N_6149,N_6137);
and U6289 (N_6289,N_6203,N_6176);
nand U6290 (N_6290,N_6242,N_6191);
or U6291 (N_6291,N_6133,N_6215);
nor U6292 (N_6292,N_6210,N_6128);
and U6293 (N_6293,N_6141,N_6179);
xnor U6294 (N_6294,N_6181,N_6206);
or U6295 (N_6295,N_6241,N_6131);
nor U6296 (N_6296,N_6189,N_6225);
or U6297 (N_6297,N_6170,N_6146);
or U6298 (N_6298,N_6175,N_6193);
and U6299 (N_6299,N_6138,N_6208);
xnor U6300 (N_6300,N_6246,N_6236);
nand U6301 (N_6301,N_6134,N_6198);
nand U6302 (N_6302,N_6166,N_6218);
and U6303 (N_6303,N_6143,N_6223);
xor U6304 (N_6304,N_6197,N_6229);
and U6305 (N_6305,N_6239,N_6202);
and U6306 (N_6306,N_6148,N_6209);
nor U6307 (N_6307,N_6127,N_6222);
nor U6308 (N_6308,N_6139,N_6144);
and U6309 (N_6309,N_6216,N_6245);
nand U6310 (N_6310,N_6211,N_6230);
xor U6311 (N_6311,N_6173,N_6174);
or U6312 (N_6312,N_6159,N_6208);
nor U6313 (N_6313,N_6184,N_6233);
and U6314 (N_6314,N_6235,N_6164);
nor U6315 (N_6315,N_6186,N_6138);
xnor U6316 (N_6316,N_6214,N_6226);
and U6317 (N_6317,N_6199,N_6249);
or U6318 (N_6318,N_6189,N_6238);
xor U6319 (N_6319,N_6210,N_6163);
or U6320 (N_6320,N_6155,N_6169);
or U6321 (N_6321,N_6135,N_6160);
or U6322 (N_6322,N_6224,N_6233);
or U6323 (N_6323,N_6201,N_6157);
or U6324 (N_6324,N_6247,N_6161);
nor U6325 (N_6325,N_6125,N_6238);
or U6326 (N_6326,N_6133,N_6236);
xnor U6327 (N_6327,N_6134,N_6126);
and U6328 (N_6328,N_6220,N_6213);
and U6329 (N_6329,N_6206,N_6238);
and U6330 (N_6330,N_6202,N_6184);
nor U6331 (N_6331,N_6228,N_6150);
or U6332 (N_6332,N_6205,N_6188);
xnor U6333 (N_6333,N_6185,N_6125);
nand U6334 (N_6334,N_6210,N_6144);
xnor U6335 (N_6335,N_6179,N_6160);
nand U6336 (N_6336,N_6236,N_6197);
or U6337 (N_6337,N_6245,N_6127);
nor U6338 (N_6338,N_6228,N_6169);
and U6339 (N_6339,N_6144,N_6190);
and U6340 (N_6340,N_6152,N_6142);
nand U6341 (N_6341,N_6158,N_6204);
xor U6342 (N_6342,N_6166,N_6148);
nor U6343 (N_6343,N_6135,N_6181);
or U6344 (N_6344,N_6137,N_6204);
xor U6345 (N_6345,N_6216,N_6135);
nand U6346 (N_6346,N_6185,N_6222);
nor U6347 (N_6347,N_6183,N_6226);
nand U6348 (N_6348,N_6183,N_6132);
nand U6349 (N_6349,N_6154,N_6234);
nor U6350 (N_6350,N_6178,N_6206);
nand U6351 (N_6351,N_6204,N_6156);
xor U6352 (N_6352,N_6230,N_6181);
nand U6353 (N_6353,N_6198,N_6130);
nand U6354 (N_6354,N_6239,N_6146);
nor U6355 (N_6355,N_6158,N_6209);
nor U6356 (N_6356,N_6169,N_6161);
xnor U6357 (N_6357,N_6179,N_6180);
or U6358 (N_6358,N_6171,N_6239);
or U6359 (N_6359,N_6212,N_6234);
or U6360 (N_6360,N_6213,N_6171);
nor U6361 (N_6361,N_6153,N_6198);
nand U6362 (N_6362,N_6146,N_6216);
xor U6363 (N_6363,N_6219,N_6175);
nand U6364 (N_6364,N_6237,N_6174);
or U6365 (N_6365,N_6247,N_6235);
or U6366 (N_6366,N_6151,N_6221);
and U6367 (N_6367,N_6184,N_6236);
nand U6368 (N_6368,N_6147,N_6135);
nand U6369 (N_6369,N_6138,N_6130);
or U6370 (N_6370,N_6172,N_6211);
or U6371 (N_6371,N_6204,N_6225);
nand U6372 (N_6372,N_6166,N_6191);
xnor U6373 (N_6373,N_6229,N_6204);
or U6374 (N_6374,N_6125,N_6179);
and U6375 (N_6375,N_6328,N_6294);
or U6376 (N_6376,N_6364,N_6301);
nand U6377 (N_6377,N_6289,N_6281);
xnor U6378 (N_6378,N_6285,N_6312);
nand U6379 (N_6379,N_6359,N_6324);
and U6380 (N_6380,N_6332,N_6365);
or U6381 (N_6381,N_6373,N_6251);
and U6382 (N_6382,N_6260,N_6310);
nor U6383 (N_6383,N_6330,N_6327);
xnor U6384 (N_6384,N_6348,N_6299);
nor U6385 (N_6385,N_6368,N_6267);
or U6386 (N_6386,N_6269,N_6313);
nand U6387 (N_6387,N_6263,N_6314);
nor U6388 (N_6388,N_6266,N_6356);
or U6389 (N_6389,N_6300,N_6268);
nand U6390 (N_6390,N_6253,N_6369);
nor U6391 (N_6391,N_6320,N_6259);
nand U6392 (N_6392,N_6340,N_6350);
nor U6393 (N_6393,N_6345,N_6349);
or U6394 (N_6394,N_6297,N_6338);
nand U6395 (N_6395,N_6309,N_6347);
nand U6396 (N_6396,N_6270,N_6296);
nand U6397 (N_6397,N_6370,N_6308);
nor U6398 (N_6398,N_6293,N_6288);
nand U6399 (N_6399,N_6272,N_6306);
nor U6400 (N_6400,N_6331,N_6276);
or U6401 (N_6401,N_6252,N_6361);
and U6402 (N_6402,N_6292,N_6358);
or U6403 (N_6403,N_6357,N_6280);
and U6404 (N_6404,N_6273,N_6321);
xor U6405 (N_6405,N_6334,N_6353);
or U6406 (N_6406,N_6274,N_6304);
nor U6407 (N_6407,N_6278,N_6352);
or U6408 (N_6408,N_6290,N_6360);
or U6409 (N_6409,N_6311,N_6250);
nor U6410 (N_6410,N_6343,N_6265);
or U6411 (N_6411,N_6333,N_6302);
nand U6412 (N_6412,N_6319,N_6355);
nand U6413 (N_6413,N_6336,N_6363);
nor U6414 (N_6414,N_6258,N_6287);
nand U6415 (N_6415,N_6329,N_6335);
nor U6416 (N_6416,N_6255,N_6362);
and U6417 (N_6417,N_6339,N_6291);
nand U6418 (N_6418,N_6371,N_6284);
or U6419 (N_6419,N_6307,N_6374);
nand U6420 (N_6420,N_6271,N_6286);
and U6421 (N_6421,N_6305,N_6275);
and U6422 (N_6422,N_6264,N_6316);
and U6423 (N_6423,N_6317,N_6318);
xor U6424 (N_6424,N_6337,N_6261);
and U6425 (N_6425,N_6372,N_6277);
and U6426 (N_6426,N_6315,N_6325);
nor U6427 (N_6427,N_6342,N_6326);
xor U6428 (N_6428,N_6295,N_6303);
nor U6429 (N_6429,N_6254,N_6283);
or U6430 (N_6430,N_6351,N_6323);
xnor U6431 (N_6431,N_6346,N_6366);
nor U6432 (N_6432,N_6257,N_6367);
nand U6433 (N_6433,N_6341,N_6322);
nor U6434 (N_6434,N_6262,N_6282);
and U6435 (N_6435,N_6279,N_6354);
xor U6436 (N_6436,N_6256,N_6344);
or U6437 (N_6437,N_6298,N_6287);
or U6438 (N_6438,N_6371,N_6361);
and U6439 (N_6439,N_6300,N_6290);
or U6440 (N_6440,N_6320,N_6329);
nand U6441 (N_6441,N_6347,N_6332);
nand U6442 (N_6442,N_6307,N_6292);
and U6443 (N_6443,N_6357,N_6255);
or U6444 (N_6444,N_6357,N_6354);
xor U6445 (N_6445,N_6257,N_6297);
nand U6446 (N_6446,N_6252,N_6258);
and U6447 (N_6447,N_6292,N_6301);
and U6448 (N_6448,N_6301,N_6367);
nor U6449 (N_6449,N_6318,N_6314);
and U6450 (N_6450,N_6287,N_6281);
xor U6451 (N_6451,N_6300,N_6372);
nand U6452 (N_6452,N_6339,N_6336);
nand U6453 (N_6453,N_6356,N_6311);
or U6454 (N_6454,N_6352,N_6315);
xnor U6455 (N_6455,N_6323,N_6340);
or U6456 (N_6456,N_6274,N_6285);
nor U6457 (N_6457,N_6367,N_6364);
or U6458 (N_6458,N_6272,N_6291);
or U6459 (N_6459,N_6311,N_6303);
nor U6460 (N_6460,N_6252,N_6307);
or U6461 (N_6461,N_6323,N_6303);
nor U6462 (N_6462,N_6263,N_6324);
nor U6463 (N_6463,N_6320,N_6324);
and U6464 (N_6464,N_6322,N_6324);
and U6465 (N_6465,N_6323,N_6309);
nor U6466 (N_6466,N_6345,N_6342);
nor U6467 (N_6467,N_6300,N_6296);
xor U6468 (N_6468,N_6342,N_6321);
xor U6469 (N_6469,N_6299,N_6363);
and U6470 (N_6470,N_6361,N_6285);
or U6471 (N_6471,N_6279,N_6309);
nand U6472 (N_6472,N_6271,N_6268);
nor U6473 (N_6473,N_6356,N_6280);
or U6474 (N_6474,N_6330,N_6320);
and U6475 (N_6475,N_6265,N_6267);
nor U6476 (N_6476,N_6254,N_6366);
nor U6477 (N_6477,N_6291,N_6279);
and U6478 (N_6478,N_6309,N_6322);
xor U6479 (N_6479,N_6338,N_6294);
and U6480 (N_6480,N_6319,N_6296);
or U6481 (N_6481,N_6305,N_6370);
xnor U6482 (N_6482,N_6278,N_6314);
nand U6483 (N_6483,N_6371,N_6362);
nor U6484 (N_6484,N_6308,N_6298);
or U6485 (N_6485,N_6252,N_6354);
or U6486 (N_6486,N_6253,N_6265);
or U6487 (N_6487,N_6323,N_6271);
nand U6488 (N_6488,N_6305,N_6312);
and U6489 (N_6489,N_6282,N_6272);
nand U6490 (N_6490,N_6354,N_6287);
xor U6491 (N_6491,N_6363,N_6335);
xnor U6492 (N_6492,N_6288,N_6321);
or U6493 (N_6493,N_6350,N_6320);
xnor U6494 (N_6494,N_6320,N_6282);
xor U6495 (N_6495,N_6325,N_6267);
or U6496 (N_6496,N_6321,N_6296);
nand U6497 (N_6497,N_6346,N_6270);
or U6498 (N_6498,N_6251,N_6366);
or U6499 (N_6499,N_6250,N_6307);
nand U6500 (N_6500,N_6459,N_6450);
nand U6501 (N_6501,N_6378,N_6413);
and U6502 (N_6502,N_6469,N_6488);
and U6503 (N_6503,N_6412,N_6449);
and U6504 (N_6504,N_6434,N_6441);
nor U6505 (N_6505,N_6415,N_6462);
and U6506 (N_6506,N_6425,N_6394);
nor U6507 (N_6507,N_6417,N_6382);
and U6508 (N_6508,N_6446,N_6409);
nor U6509 (N_6509,N_6426,N_6397);
xor U6510 (N_6510,N_6401,N_6388);
or U6511 (N_6511,N_6439,N_6411);
nand U6512 (N_6512,N_6489,N_6435);
xor U6513 (N_6513,N_6437,N_6438);
xnor U6514 (N_6514,N_6460,N_6393);
nand U6515 (N_6515,N_6499,N_6475);
nor U6516 (N_6516,N_6482,N_6457);
xor U6517 (N_6517,N_6497,N_6456);
or U6518 (N_6518,N_6410,N_6395);
and U6519 (N_6519,N_6443,N_6420);
and U6520 (N_6520,N_6383,N_6491);
xnor U6521 (N_6521,N_6442,N_6405);
or U6522 (N_6522,N_6452,N_6471);
or U6523 (N_6523,N_6422,N_6483);
nor U6524 (N_6524,N_6468,N_6448);
or U6525 (N_6525,N_6432,N_6464);
nand U6526 (N_6526,N_6377,N_6403);
or U6527 (N_6527,N_6453,N_6381);
nand U6528 (N_6528,N_6474,N_6375);
xnor U6529 (N_6529,N_6428,N_6386);
nor U6530 (N_6530,N_6487,N_6385);
and U6531 (N_6531,N_6436,N_6376);
or U6532 (N_6532,N_6494,N_6472);
nor U6533 (N_6533,N_6465,N_6485);
or U6534 (N_6534,N_6414,N_6467);
and U6535 (N_6535,N_6379,N_6498);
xnor U6536 (N_6536,N_6444,N_6387);
and U6537 (N_6537,N_6479,N_6427);
nor U6538 (N_6538,N_6486,N_6389);
and U6539 (N_6539,N_6418,N_6447);
or U6540 (N_6540,N_6440,N_6454);
nand U6541 (N_6541,N_6476,N_6398);
and U6542 (N_6542,N_6391,N_6430);
xnor U6543 (N_6543,N_6392,N_6493);
xor U6544 (N_6544,N_6495,N_6380);
nand U6545 (N_6545,N_6419,N_6484);
or U6546 (N_6546,N_6463,N_6451);
nor U6547 (N_6547,N_6429,N_6384);
or U6548 (N_6548,N_6423,N_6470);
and U6549 (N_6549,N_6406,N_6396);
nor U6550 (N_6550,N_6416,N_6492);
nand U6551 (N_6551,N_6466,N_6496);
and U6552 (N_6552,N_6478,N_6455);
or U6553 (N_6553,N_6424,N_6473);
nand U6554 (N_6554,N_6407,N_6404);
and U6555 (N_6555,N_6408,N_6490);
nand U6556 (N_6556,N_6461,N_6399);
xor U6557 (N_6557,N_6402,N_6400);
xnor U6558 (N_6558,N_6421,N_6481);
xor U6559 (N_6559,N_6480,N_6431);
nor U6560 (N_6560,N_6390,N_6458);
nand U6561 (N_6561,N_6445,N_6433);
nand U6562 (N_6562,N_6477,N_6427);
and U6563 (N_6563,N_6441,N_6388);
and U6564 (N_6564,N_6406,N_6496);
and U6565 (N_6565,N_6377,N_6482);
or U6566 (N_6566,N_6417,N_6489);
and U6567 (N_6567,N_6497,N_6428);
nand U6568 (N_6568,N_6466,N_6498);
nand U6569 (N_6569,N_6478,N_6458);
nand U6570 (N_6570,N_6421,N_6461);
nand U6571 (N_6571,N_6481,N_6476);
xnor U6572 (N_6572,N_6481,N_6439);
and U6573 (N_6573,N_6462,N_6437);
and U6574 (N_6574,N_6430,N_6386);
or U6575 (N_6575,N_6483,N_6403);
nand U6576 (N_6576,N_6460,N_6383);
or U6577 (N_6577,N_6376,N_6400);
nand U6578 (N_6578,N_6484,N_6478);
nor U6579 (N_6579,N_6465,N_6434);
nor U6580 (N_6580,N_6430,N_6447);
and U6581 (N_6581,N_6393,N_6439);
xnor U6582 (N_6582,N_6413,N_6447);
and U6583 (N_6583,N_6495,N_6456);
or U6584 (N_6584,N_6436,N_6419);
nand U6585 (N_6585,N_6376,N_6417);
nor U6586 (N_6586,N_6411,N_6400);
nor U6587 (N_6587,N_6406,N_6408);
xor U6588 (N_6588,N_6376,N_6454);
nor U6589 (N_6589,N_6390,N_6431);
or U6590 (N_6590,N_6491,N_6453);
nor U6591 (N_6591,N_6421,N_6378);
xnor U6592 (N_6592,N_6492,N_6440);
and U6593 (N_6593,N_6389,N_6455);
xor U6594 (N_6594,N_6403,N_6486);
nand U6595 (N_6595,N_6395,N_6461);
xor U6596 (N_6596,N_6493,N_6410);
xor U6597 (N_6597,N_6447,N_6412);
nor U6598 (N_6598,N_6494,N_6429);
nor U6599 (N_6599,N_6491,N_6411);
and U6600 (N_6600,N_6395,N_6486);
and U6601 (N_6601,N_6416,N_6451);
xnor U6602 (N_6602,N_6462,N_6489);
or U6603 (N_6603,N_6499,N_6411);
xor U6604 (N_6604,N_6467,N_6494);
nor U6605 (N_6605,N_6402,N_6418);
nand U6606 (N_6606,N_6492,N_6395);
or U6607 (N_6607,N_6398,N_6408);
nor U6608 (N_6608,N_6465,N_6407);
xor U6609 (N_6609,N_6379,N_6490);
and U6610 (N_6610,N_6476,N_6377);
or U6611 (N_6611,N_6470,N_6375);
and U6612 (N_6612,N_6488,N_6415);
nor U6613 (N_6613,N_6386,N_6405);
xor U6614 (N_6614,N_6458,N_6468);
and U6615 (N_6615,N_6460,N_6426);
nor U6616 (N_6616,N_6392,N_6435);
xnor U6617 (N_6617,N_6388,N_6453);
nor U6618 (N_6618,N_6471,N_6396);
nand U6619 (N_6619,N_6497,N_6495);
nor U6620 (N_6620,N_6487,N_6429);
nor U6621 (N_6621,N_6411,N_6383);
or U6622 (N_6622,N_6382,N_6377);
or U6623 (N_6623,N_6460,N_6407);
xor U6624 (N_6624,N_6481,N_6400);
and U6625 (N_6625,N_6605,N_6602);
and U6626 (N_6626,N_6561,N_6621);
xnor U6627 (N_6627,N_6547,N_6564);
xor U6628 (N_6628,N_6592,N_6523);
xnor U6629 (N_6629,N_6565,N_6617);
xnor U6630 (N_6630,N_6591,N_6593);
and U6631 (N_6631,N_6512,N_6580);
or U6632 (N_6632,N_6571,N_6520);
or U6633 (N_6633,N_6532,N_6609);
and U6634 (N_6634,N_6536,N_6587);
nor U6635 (N_6635,N_6503,N_6502);
nor U6636 (N_6636,N_6508,N_6515);
nor U6637 (N_6637,N_6516,N_6509);
nor U6638 (N_6638,N_6539,N_6511);
nor U6639 (N_6639,N_6537,N_6500);
nor U6640 (N_6640,N_6541,N_6519);
or U6641 (N_6641,N_6535,N_6599);
nand U6642 (N_6642,N_6606,N_6607);
nor U6643 (N_6643,N_6595,N_6575);
nand U6644 (N_6644,N_6522,N_6619);
xor U6645 (N_6645,N_6563,N_6558);
or U6646 (N_6646,N_6578,N_6501);
and U6647 (N_6647,N_6514,N_6585);
and U6648 (N_6648,N_6560,N_6618);
nand U6649 (N_6649,N_6555,N_6588);
xnor U6650 (N_6650,N_6528,N_6584);
or U6651 (N_6651,N_6566,N_6548);
nor U6652 (N_6652,N_6505,N_6562);
xnor U6653 (N_6653,N_6554,N_6567);
nand U6654 (N_6654,N_6612,N_6596);
or U6655 (N_6655,N_6524,N_6576);
xnor U6656 (N_6656,N_6594,N_6569);
nor U6657 (N_6657,N_6615,N_6597);
nand U6658 (N_6658,N_6538,N_6624);
xor U6659 (N_6659,N_6623,N_6543);
xnor U6660 (N_6660,N_6544,N_6603);
nand U6661 (N_6661,N_6550,N_6573);
and U6662 (N_6662,N_6521,N_6542);
or U6663 (N_6663,N_6530,N_6582);
xnor U6664 (N_6664,N_6556,N_6526);
and U6665 (N_6665,N_6586,N_6589);
xnor U6666 (N_6666,N_6570,N_6527);
and U6667 (N_6667,N_6545,N_6518);
nand U6668 (N_6668,N_6513,N_6551);
nand U6669 (N_6669,N_6590,N_6506);
and U6670 (N_6670,N_6507,N_6600);
nor U6671 (N_6671,N_6557,N_6549);
nand U6672 (N_6672,N_6577,N_6525);
xnor U6673 (N_6673,N_6598,N_6529);
xnor U6674 (N_6674,N_6601,N_6614);
nor U6675 (N_6675,N_6534,N_6581);
or U6676 (N_6676,N_6574,N_6620);
nor U6677 (N_6677,N_6552,N_6616);
nor U6678 (N_6678,N_6613,N_6622);
nand U6679 (N_6679,N_6572,N_6568);
nor U6680 (N_6680,N_6546,N_6553);
xor U6681 (N_6681,N_6608,N_6540);
nand U6682 (N_6682,N_6559,N_6604);
xor U6683 (N_6683,N_6510,N_6611);
xor U6684 (N_6684,N_6504,N_6517);
xor U6685 (N_6685,N_6579,N_6610);
nor U6686 (N_6686,N_6531,N_6533);
nor U6687 (N_6687,N_6583,N_6510);
or U6688 (N_6688,N_6598,N_6600);
nand U6689 (N_6689,N_6526,N_6559);
xor U6690 (N_6690,N_6535,N_6547);
or U6691 (N_6691,N_6514,N_6552);
or U6692 (N_6692,N_6525,N_6596);
and U6693 (N_6693,N_6531,N_6554);
nand U6694 (N_6694,N_6520,N_6547);
and U6695 (N_6695,N_6528,N_6617);
or U6696 (N_6696,N_6557,N_6501);
nand U6697 (N_6697,N_6581,N_6510);
and U6698 (N_6698,N_6543,N_6618);
nand U6699 (N_6699,N_6556,N_6603);
or U6700 (N_6700,N_6518,N_6549);
nor U6701 (N_6701,N_6514,N_6546);
or U6702 (N_6702,N_6550,N_6590);
and U6703 (N_6703,N_6579,N_6620);
and U6704 (N_6704,N_6610,N_6619);
and U6705 (N_6705,N_6506,N_6578);
nand U6706 (N_6706,N_6613,N_6562);
xnor U6707 (N_6707,N_6517,N_6506);
or U6708 (N_6708,N_6513,N_6529);
nor U6709 (N_6709,N_6501,N_6526);
and U6710 (N_6710,N_6562,N_6581);
or U6711 (N_6711,N_6517,N_6595);
nand U6712 (N_6712,N_6518,N_6522);
or U6713 (N_6713,N_6543,N_6608);
xnor U6714 (N_6714,N_6570,N_6602);
and U6715 (N_6715,N_6614,N_6538);
nor U6716 (N_6716,N_6613,N_6502);
nand U6717 (N_6717,N_6529,N_6549);
xnor U6718 (N_6718,N_6554,N_6583);
and U6719 (N_6719,N_6547,N_6569);
nand U6720 (N_6720,N_6594,N_6621);
and U6721 (N_6721,N_6553,N_6520);
and U6722 (N_6722,N_6602,N_6606);
and U6723 (N_6723,N_6566,N_6593);
or U6724 (N_6724,N_6530,N_6547);
nor U6725 (N_6725,N_6520,N_6600);
xnor U6726 (N_6726,N_6505,N_6545);
or U6727 (N_6727,N_6541,N_6618);
or U6728 (N_6728,N_6623,N_6510);
or U6729 (N_6729,N_6502,N_6509);
nand U6730 (N_6730,N_6577,N_6544);
and U6731 (N_6731,N_6604,N_6560);
xor U6732 (N_6732,N_6582,N_6598);
xor U6733 (N_6733,N_6574,N_6566);
xnor U6734 (N_6734,N_6623,N_6551);
and U6735 (N_6735,N_6592,N_6594);
or U6736 (N_6736,N_6525,N_6503);
nor U6737 (N_6737,N_6500,N_6508);
nand U6738 (N_6738,N_6607,N_6536);
and U6739 (N_6739,N_6555,N_6505);
or U6740 (N_6740,N_6554,N_6581);
or U6741 (N_6741,N_6594,N_6515);
nand U6742 (N_6742,N_6572,N_6570);
nor U6743 (N_6743,N_6613,N_6555);
xor U6744 (N_6744,N_6532,N_6506);
or U6745 (N_6745,N_6577,N_6538);
or U6746 (N_6746,N_6603,N_6505);
nand U6747 (N_6747,N_6604,N_6523);
nor U6748 (N_6748,N_6520,N_6550);
nand U6749 (N_6749,N_6531,N_6561);
xor U6750 (N_6750,N_6744,N_6654);
or U6751 (N_6751,N_6626,N_6668);
or U6752 (N_6752,N_6628,N_6680);
xnor U6753 (N_6753,N_6659,N_6676);
nor U6754 (N_6754,N_6660,N_6655);
nor U6755 (N_6755,N_6672,N_6749);
nor U6756 (N_6756,N_6636,N_6707);
xnor U6757 (N_6757,N_6737,N_6631);
nand U6758 (N_6758,N_6716,N_6641);
nor U6759 (N_6759,N_6667,N_6688);
xnor U6760 (N_6760,N_6698,N_6703);
xnor U6761 (N_6761,N_6692,N_6651);
or U6762 (N_6762,N_6644,N_6646);
nand U6763 (N_6763,N_6743,N_6695);
nor U6764 (N_6764,N_6671,N_6694);
nand U6765 (N_6765,N_6693,N_6685);
and U6766 (N_6766,N_6720,N_6734);
and U6767 (N_6767,N_6648,N_6745);
nand U6768 (N_6768,N_6632,N_6658);
nor U6769 (N_6769,N_6709,N_6679);
and U6770 (N_6770,N_6645,N_6643);
xnor U6771 (N_6771,N_6724,N_6711);
or U6772 (N_6772,N_6706,N_6735);
and U6773 (N_6773,N_6691,N_6687);
or U6774 (N_6774,N_6725,N_6666);
and U6775 (N_6775,N_6686,N_6683);
nand U6776 (N_6776,N_6670,N_6682);
or U6777 (N_6777,N_6718,N_6663);
nor U6778 (N_6778,N_6649,N_6717);
nand U6779 (N_6779,N_6705,N_6675);
xnor U6780 (N_6780,N_6640,N_6731);
xor U6781 (N_6781,N_6684,N_6678);
nor U6782 (N_6782,N_6637,N_6677);
or U6783 (N_6783,N_6652,N_6738);
xor U6784 (N_6784,N_6722,N_6748);
nand U6785 (N_6785,N_6697,N_6723);
nand U6786 (N_6786,N_6736,N_6712);
and U6787 (N_6787,N_6719,N_6661);
nand U6788 (N_6788,N_6689,N_6729);
or U6789 (N_6789,N_6710,N_6733);
and U6790 (N_6790,N_6635,N_6625);
and U6791 (N_6791,N_6638,N_6681);
nand U6792 (N_6792,N_6740,N_6642);
and U6793 (N_6793,N_6739,N_6630);
xor U6794 (N_6794,N_6732,N_6700);
nand U6795 (N_6795,N_6704,N_6662);
nor U6796 (N_6796,N_6714,N_6639);
xor U6797 (N_6797,N_6726,N_6728);
nand U6798 (N_6798,N_6657,N_6664);
or U6799 (N_6799,N_6741,N_6673);
or U6800 (N_6800,N_6634,N_6715);
nor U6801 (N_6801,N_6730,N_6702);
and U6802 (N_6802,N_6665,N_6742);
or U6803 (N_6803,N_6721,N_6627);
or U6804 (N_6804,N_6633,N_6708);
and U6805 (N_6805,N_6674,N_6747);
and U6806 (N_6806,N_6653,N_6669);
xnor U6807 (N_6807,N_6746,N_6656);
and U6808 (N_6808,N_6727,N_6696);
nor U6809 (N_6809,N_6699,N_6647);
xnor U6810 (N_6810,N_6629,N_6701);
or U6811 (N_6811,N_6713,N_6650);
nand U6812 (N_6812,N_6690,N_6675);
or U6813 (N_6813,N_6667,N_6676);
and U6814 (N_6814,N_6717,N_6658);
and U6815 (N_6815,N_6662,N_6681);
xnor U6816 (N_6816,N_6674,N_6735);
and U6817 (N_6817,N_6713,N_6707);
nor U6818 (N_6818,N_6693,N_6634);
nor U6819 (N_6819,N_6633,N_6701);
xnor U6820 (N_6820,N_6738,N_6654);
or U6821 (N_6821,N_6731,N_6659);
and U6822 (N_6822,N_6739,N_6696);
xnor U6823 (N_6823,N_6694,N_6657);
and U6824 (N_6824,N_6700,N_6661);
and U6825 (N_6825,N_6695,N_6716);
and U6826 (N_6826,N_6629,N_6732);
or U6827 (N_6827,N_6735,N_6673);
and U6828 (N_6828,N_6732,N_6660);
nor U6829 (N_6829,N_6648,N_6707);
nor U6830 (N_6830,N_6625,N_6691);
or U6831 (N_6831,N_6691,N_6747);
nand U6832 (N_6832,N_6628,N_6685);
nor U6833 (N_6833,N_6710,N_6650);
xor U6834 (N_6834,N_6636,N_6632);
or U6835 (N_6835,N_6685,N_6640);
nand U6836 (N_6836,N_6660,N_6713);
or U6837 (N_6837,N_6738,N_6742);
xor U6838 (N_6838,N_6647,N_6747);
and U6839 (N_6839,N_6675,N_6736);
nor U6840 (N_6840,N_6739,N_6659);
nand U6841 (N_6841,N_6741,N_6716);
nor U6842 (N_6842,N_6660,N_6702);
xnor U6843 (N_6843,N_6638,N_6747);
and U6844 (N_6844,N_6668,N_6724);
xor U6845 (N_6845,N_6705,N_6704);
or U6846 (N_6846,N_6637,N_6702);
or U6847 (N_6847,N_6632,N_6660);
nand U6848 (N_6848,N_6625,N_6709);
nor U6849 (N_6849,N_6641,N_6647);
nor U6850 (N_6850,N_6740,N_6736);
nand U6851 (N_6851,N_6663,N_6659);
nor U6852 (N_6852,N_6662,N_6650);
nor U6853 (N_6853,N_6667,N_6745);
and U6854 (N_6854,N_6697,N_6712);
xnor U6855 (N_6855,N_6628,N_6674);
or U6856 (N_6856,N_6639,N_6635);
xor U6857 (N_6857,N_6721,N_6636);
nor U6858 (N_6858,N_6681,N_6722);
and U6859 (N_6859,N_6737,N_6739);
or U6860 (N_6860,N_6639,N_6735);
nor U6861 (N_6861,N_6664,N_6697);
or U6862 (N_6862,N_6729,N_6716);
or U6863 (N_6863,N_6686,N_6653);
or U6864 (N_6864,N_6657,N_6699);
or U6865 (N_6865,N_6714,N_6725);
or U6866 (N_6866,N_6681,N_6710);
and U6867 (N_6867,N_6713,N_6683);
nand U6868 (N_6868,N_6682,N_6698);
or U6869 (N_6869,N_6629,N_6746);
nor U6870 (N_6870,N_6656,N_6651);
and U6871 (N_6871,N_6688,N_6747);
or U6872 (N_6872,N_6684,N_6667);
nor U6873 (N_6873,N_6719,N_6690);
nor U6874 (N_6874,N_6740,N_6643);
xnor U6875 (N_6875,N_6762,N_6844);
nand U6876 (N_6876,N_6767,N_6754);
nor U6877 (N_6877,N_6752,N_6814);
xnor U6878 (N_6878,N_6856,N_6755);
nor U6879 (N_6879,N_6774,N_6863);
and U6880 (N_6880,N_6772,N_6837);
nand U6881 (N_6881,N_6853,N_6847);
and U6882 (N_6882,N_6764,N_6768);
or U6883 (N_6883,N_6843,N_6776);
nand U6884 (N_6884,N_6798,N_6832);
nor U6885 (N_6885,N_6806,N_6804);
nor U6886 (N_6886,N_6873,N_6820);
and U6887 (N_6887,N_6807,N_6791);
or U6888 (N_6888,N_6846,N_6835);
xor U6889 (N_6889,N_6860,N_6780);
nor U6890 (N_6890,N_6855,N_6809);
nor U6891 (N_6891,N_6784,N_6833);
nor U6892 (N_6892,N_6818,N_6808);
and U6893 (N_6893,N_6852,N_6848);
xor U6894 (N_6894,N_6757,N_6777);
nand U6895 (N_6895,N_6822,N_6865);
or U6896 (N_6896,N_6816,N_6786);
or U6897 (N_6897,N_6828,N_6795);
or U6898 (N_6898,N_6851,N_6758);
nand U6899 (N_6899,N_6773,N_6838);
nor U6900 (N_6900,N_6766,N_6760);
xor U6901 (N_6901,N_6858,N_6765);
nor U6902 (N_6902,N_6836,N_6783);
nand U6903 (N_6903,N_6779,N_6870);
and U6904 (N_6904,N_6854,N_6845);
and U6905 (N_6905,N_6785,N_6792);
or U6906 (N_6906,N_6841,N_6793);
xnor U6907 (N_6907,N_6866,N_6874);
nand U6908 (N_6908,N_6787,N_6790);
or U6909 (N_6909,N_6799,N_6829);
nor U6910 (N_6910,N_6810,N_6794);
and U6911 (N_6911,N_6868,N_6782);
and U6912 (N_6912,N_6797,N_6827);
or U6913 (N_6913,N_6857,N_6769);
nand U6914 (N_6914,N_6761,N_6824);
xor U6915 (N_6915,N_6763,N_6819);
nand U6916 (N_6916,N_6778,N_6840);
and U6917 (N_6917,N_6753,N_6770);
and U6918 (N_6918,N_6796,N_6812);
nor U6919 (N_6919,N_6759,N_6788);
xor U6920 (N_6920,N_6849,N_6869);
xnor U6921 (N_6921,N_6803,N_6756);
nor U6922 (N_6922,N_6821,N_6789);
and U6923 (N_6923,N_6861,N_6815);
xnor U6924 (N_6924,N_6862,N_6867);
or U6925 (N_6925,N_6805,N_6802);
xor U6926 (N_6926,N_6830,N_6825);
nand U6927 (N_6927,N_6811,N_6842);
nor U6928 (N_6928,N_6775,N_6823);
and U6929 (N_6929,N_6750,N_6813);
nand U6930 (N_6930,N_6834,N_6801);
xnor U6931 (N_6931,N_6831,N_6850);
nand U6932 (N_6932,N_6839,N_6800);
nor U6933 (N_6933,N_6826,N_6817);
xnor U6934 (N_6934,N_6781,N_6771);
or U6935 (N_6935,N_6859,N_6864);
and U6936 (N_6936,N_6872,N_6751);
xor U6937 (N_6937,N_6871,N_6827);
nand U6938 (N_6938,N_6851,N_6757);
nand U6939 (N_6939,N_6775,N_6848);
or U6940 (N_6940,N_6787,N_6770);
or U6941 (N_6941,N_6855,N_6833);
or U6942 (N_6942,N_6824,N_6817);
and U6943 (N_6943,N_6778,N_6802);
xor U6944 (N_6944,N_6774,N_6810);
xor U6945 (N_6945,N_6846,N_6872);
and U6946 (N_6946,N_6755,N_6813);
nor U6947 (N_6947,N_6775,N_6753);
nor U6948 (N_6948,N_6873,N_6855);
or U6949 (N_6949,N_6786,N_6806);
nor U6950 (N_6950,N_6851,N_6804);
xor U6951 (N_6951,N_6838,N_6776);
or U6952 (N_6952,N_6794,N_6823);
and U6953 (N_6953,N_6862,N_6760);
or U6954 (N_6954,N_6792,N_6811);
xor U6955 (N_6955,N_6846,N_6818);
nor U6956 (N_6956,N_6825,N_6761);
or U6957 (N_6957,N_6861,N_6843);
or U6958 (N_6958,N_6782,N_6806);
and U6959 (N_6959,N_6805,N_6796);
xnor U6960 (N_6960,N_6823,N_6873);
nand U6961 (N_6961,N_6841,N_6826);
or U6962 (N_6962,N_6839,N_6824);
or U6963 (N_6963,N_6789,N_6802);
and U6964 (N_6964,N_6774,N_6791);
nor U6965 (N_6965,N_6766,N_6843);
and U6966 (N_6966,N_6810,N_6765);
nand U6967 (N_6967,N_6776,N_6804);
nand U6968 (N_6968,N_6834,N_6804);
or U6969 (N_6969,N_6810,N_6760);
xnor U6970 (N_6970,N_6778,N_6780);
nand U6971 (N_6971,N_6761,N_6860);
xnor U6972 (N_6972,N_6759,N_6864);
nand U6973 (N_6973,N_6831,N_6839);
and U6974 (N_6974,N_6823,N_6780);
nand U6975 (N_6975,N_6863,N_6837);
nand U6976 (N_6976,N_6829,N_6859);
nand U6977 (N_6977,N_6800,N_6788);
nor U6978 (N_6978,N_6764,N_6806);
nor U6979 (N_6979,N_6828,N_6779);
and U6980 (N_6980,N_6829,N_6763);
nor U6981 (N_6981,N_6790,N_6756);
xnor U6982 (N_6982,N_6773,N_6845);
or U6983 (N_6983,N_6836,N_6857);
and U6984 (N_6984,N_6820,N_6816);
nand U6985 (N_6985,N_6753,N_6802);
and U6986 (N_6986,N_6784,N_6756);
xor U6987 (N_6987,N_6854,N_6767);
or U6988 (N_6988,N_6870,N_6798);
xor U6989 (N_6989,N_6848,N_6794);
nor U6990 (N_6990,N_6756,N_6802);
nor U6991 (N_6991,N_6837,N_6801);
nand U6992 (N_6992,N_6814,N_6846);
nor U6993 (N_6993,N_6790,N_6834);
or U6994 (N_6994,N_6751,N_6835);
or U6995 (N_6995,N_6820,N_6791);
or U6996 (N_6996,N_6850,N_6871);
or U6997 (N_6997,N_6787,N_6868);
and U6998 (N_6998,N_6854,N_6844);
nand U6999 (N_6999,N_6831,N_6802);
nor U7000 (N_7000,N_6996,N_6912);
or U7001 (N_7001,N_6900,N_6885);
and U7002 (N_7002,N_6894,N_6896);
nor U7003 (N_7003,N_6969,N_6929);
xor U7004 (N_7004,N_6962,N_6977);
and U7005 (N_7005,N_6907,N_6940);
and U7006 (N_7006,N_6902,N_6998);
xnor U7007 (N_7007,N_6987,N_6892);
or U7008 (N_7008,N_6948,N_6972);
or U7009 (N_7009,N_6978,N_6931);
and U7010 (N_7010,N_6952,N_6963);
nand U7011 (N_7011,N_6986,N_6895);
nor U7012 (N_7012,N_6964,N_6932);
and U7013 (N_7013,N_6997,N_6889);
nor U7014 (N_7014,N_6893,N_6985);
nand U7015 (N_7015,N_6949,N_6946);
xnor U7016 (N_7016,N_6890,N_6981);
xor U7017 (N_7017,N_6908,N_6957);
nor U7018 (N_7018,N_6924,N_6980);
nor U7019 (N_7019,N_6875,N_6923);
nand U7020 (N_7020,N_6994,N_6979);
or U7021 (N_7021,N_6999,N_6915);
and U7022 (N_7022,N_6877,N_6958);
and U7023 (N_7023,N_6939,N_6909);
and U7024 (N_7024,N_6956,N_6911);
and U7025 (N_7025,N_6955,N_6961);
xnor U7026 (N_7026,N_6930,N_6886);
and U7027 (N_7027,N_6888,N_6954);
or U7028 (N_7028,N_6920,N_6941);
xnor U7029 (N_7029,N_6950,N_6995);
nand U7030 (N_7030,N_6910,N_6938);
nand U7031 (N_7031,N_6988,N_6934);
nand U7032 (N_7032,N_6984,N_6951);
and U7033 (N_7033,N_6913,N_6966);
nor U7034 (N_7034,N_6947,N_6901);
nand U7035 (N_7035,N_6959,N_6906);
or U7036 (N_7036,N_6925,N_6918);
nand U7037 (N_7037,N_6876,N_6968);
nor U7038 (N_7038,N_6971,N_6904);
nor U7039 (N_7039,N_6897,N_6975);
and U7040 (N_7040,N_6914,N_6973);
and U7041 (N_7041,N_6992,N_6935);
nand U7042 (N_7042,N_6945,N_6917);
nand U7043 (N_7043,N_6944,N_6960);
and U7044 (N_7044,N_6953,N_6974);
xor U7045 (N_7045,N_6905,N_6967);
nand U7046 (N_7046,N_6982,N_6899);
xor U7047 (N_7047,N_6880,N_6922);
xor U7048 (N_7048,N_6879,N_6916);
nand U7049 (N_7049,N_6993,N_6926);
and U7050 (N_7050,N_6881,N_6943);
nor U7051 (N_7051,N_6884,N_6983);
nor U7052 (N_7052,N_6898,N_6942);
xor U7053 (N_7053,N_6928,N_6882);
xor U7054 (N_7054,N_6933,N_6878);
xor U7055 (N_7055,N_6936,N_6970);
xor U7056 (N_7056,N_6919,N_6887);
nor U7057 (N_7057,N_6989,N_6937);
nor U7058 (N_7058,N_6976,N_6891);
or U7059 (N_7059,N_6921,N_6883);
nor U7060 (N_7060,N_6990,N_6991);
nor U7061 (N_7061,N_6965,N_6927);
or U7062 (N_7062,N_6903,N_6899);
nor U7063 (N_7063,N_6978,N_6941);
nand U7064 (N_7064,N_6931,N_6914);
nor U7065 (N_7065,N_6928,N_6898);
nor U7066 (N_7066,N_6895,N_6881);
xor U7067 (N_7067,N_6917,N_6978);
nor U7068 (N_7068,N_6959,N_6903);
nor U7069 (N_7069,N_6943,N_6899);
or U7070 (N_7070,N_6919,N_6929);
or U7071 (N_7071,N_6915,N_6945);
xor U7072 (N_7072,N_6983,N_6918);
nand U7073 (N_7073,N_6934,N_6946);
and U7074 (N_7074,N_6992,N_6910);
xnor U7075 (N_7075,N_6920,N_6958);
nor U7076 (N_7076,N_6889,N_6959);
and U7077 (N_7077,N_6981,N_6968);
nor U7078 (N_7078,N_6983,N_6893);
or U7079 (N_7079,N_6886,N_6997);
xor U7080 (N_7080,N_6990,N_6903);
nor U7081 (N_7081,N_6923,N_6926);
and U7082 (N_7082,N_6986,N_6953);
or U7083 (N_7083,N_6995,N_6956);
xor U7084 (N_7084,N_6899,N_6958);
nand U7085 (N_7085,N_6969,N_6962);
nor U7086 (N_7086,N_6922,N_6988);
nand U7087 (N_7087,N_6966,N_6892);
nor U7088 (N_7088,N_6905,N_6906);
or U7089 (N_7089,N_6995,N_6914);
or U7090 (N_7090,N_6906,N_6984);
nor U7091 (N_7091,N_6964,N_6988);
or U7092 (N_7092,N_6961,N_6926);
nor U7093 (N_7093,N_6971,N_6920);
or U7094 (N_7094,N_6914,N_6963);
or U7095 (N_7095,N_6987,N_6907);
nand U7096 (N_7096,N_6893,N_6957);
nor U7097 (N_7097,N_6981,N_6879);
or U7098 (N_7098,N_6887,N_6959);
xnor U7099 (N_7099,N_6908,N_6962);
xor U7100 (N_7100,N_6917,N_6922);
or U7101 (N_7101,N_6966,N_6911);
nor U7102 (N_7102,N_6957,N_6876);
nand U7103 (N_7103,N_6883,N_6971);
and U7104 (N_7104,N_6876,N_6932);
nand U7105 (N_7105,N_6951,N_6939);
and U7106 (N_7106,N_6883,N_6988);
nor U7107 (N_7107,N_6887,N_6977);
nand U7108 (N_7108,N_6882,N_6978);
and U7109 (N_7109,N_6999,N_6925);
and U7110 (N_7110,N_6987,N_6953);
and U7111 (N_7111,N_6949,N_6905);
and U7112 (N_7112,N_6915,N_6970);
nor U7113 (N_7113,N_6938,N_6878);
and U7114 (N_7114,N_6967,N_6993);
nand U7115 (N_7115,N_6952,N_6949);
and U7116 (N_7116,N_6964,N_6919);
and U7117 (N_7117,N_6955,N_6962);
nor U7118 (N_7118,N_6886,N_6943);
nor U7119 (N_7119,N_6876,N_6901);
nand U7120 (N_7120,N_6996,N_6949);
nand U7121 (N_7121,N_6939,N_6988);
and U7122 (N_7122,N_6888,N_6894);
nand U7123 (N_7123,N_6942,N_6988);
or U7124 (N_7124,N_6966,N_6998);
nor U7125 (N_7125,N_7115,N_7093);
nand U7126 (N_7126,N_7103,N_7005);
nor U7127 (N_7127,N_7025,N_7104);
and U7128 (N_7128,N_7033,N_7030);
nand U7129 (N_7129,N_7042,N_7015);
nor U7130 (N_7130,N_7088,N_7054);
nor U7131 (N_7131,N_7019,N_7056);
nor U7132 (N_7132,N_7045,N_7009);
nand U7133 (N_7133,N_7047,N_7026);
nor U7134 (N_7134,N_7077,N_7073);
nand U7135 (N_7135,N_7024,N_7041);
or U7136 (N_7136,N_7086,N_7096);
xnor U7137 (N_7137,N_7043,N_7117);
nor U7138 (N_7138,N_7010,N_7106);
nand U7139 (N_7139,N_7051,N_7050);
nor U7140 (N_7140,N_7062,N_7023);
nor U7141 (N_7141,N_7018,N_7089);
xnor U7142 (N_7142,N_7074,N_7065);
nor U7143 (N_7143,N_7122,N_7003);
nand U7144 (N_7144,N_7108,N_7100);
nor U7145 (N_7145,N_7070,N_7111);
nand U7146 (N_7146,N_7032,N_7022);
or U7147 (N_7147,N_7069,N_7071);
xor U7148 (N_7148,N_7028,N_7078);
nor U7149 (N_7149,N_7094,N_7034);
and U7150 (N_7150,N_7000,N_7004);
or U7151 (N_7151,N_7040,N_7080);
xor U7152 (N_7152,N_7085,N_7013);
nand U7153 (N_7153,N_7014,N_7002);
nand U7154 (N_7154,N_7113,N_7012);
nor U7155 (N_7155,N_7101,N_7064);
nor U7156 (N_7156,N_7055,N_7109);
nand U7157 (N_7157,N_7123,N_7027);
nor U7158 (N_7158,N_7059,N_7039);
or U7159 (N_7159,N_7107,N_7006);
xnor U7160 (N_7160,N_7017,N_7110);
nand U7161 (N_7161,N_7057,N_7008);
nor U7162 (N_7162,N_7066,N_7099);
xnor U7163 (N_7163,N_7046,N_7083);
nor U7164 (N_7164,N_7098,N_7067);
nor U7165 (N_7165,N_7095,N_7036);
or U7166 (N_7166,N_7081,N_7116);
nand U7167 (N_7167,N_7052,N_7114);
xnor U7168 (N_7168,N_7038,N_7090);
and U7169 (N_7169,N_7020,N_7091);
nand U7170 (N_7170,N_7044,N_7082);
and U7171 (N_7171,N_7124,N_7021);
and U7172 (N_7172,N_7118,N_7037);
xor U7173 (N_7173,N_7053,N_7076);
xnor U7174 (N_7174,N_7011,N_7119);
and U7175 (N_7175,N_7084,N_7058);
nand U7176 (N_7176,N_7097,N_7007);
or U7177 (N_7177,N_7121,N_7048);
xor U7178 (N_7178,N_7087,N_7112);
xor U7179 (N_7179,N_7049,N_7016);
or U7180 (N_7180,N_7031,N_7072);
and U7181 (N_7181,N_7105,N_7001);
xor U7182 (N_7182,N_7120,N_7092);
nor U7183 (N_7183,N_7063,N_7102);
and U7184 (N_7184,N_7029,N_7061);
and U7185 (N_7185,N_7079,N_7068);
nand U7186 (N_7186,N_7075,N_7060);
nor U7187 (N_7187,N_7035,N_7094);
nand U7188 (N_7188,N_7121,N_7106);
nand U7189 (N_7189,N_7062,N_7014);
xnor U7190 (N_7190,N_7098,N_7030);
nor U7191 (N_7191,N_7011,N_7061);
and U7192 (N_7192,N_7094,N_7058);
xnor U7193 (N_7193,N_7121,N_7006);
and U7194 (N_7194,N_7024,N_7025);
or U7195 (N_7195,N_7025,N_7082);
and U7196 (N_7196,N_7095,N_7117);
xnor U7197 (N_7197,N_7075,N_7089);
xor U7198 (N_7198,N_7047,N_7032);
nand U7199 (N_7199,N_7045,N_7096);
or U7200 (N_7200,N_7068,N_7110);
and U7201 (N_7201,N_7112,N_7109);
or U7202 (N_7202,N_7029,N_7098);
nor U7203 (N_7203,N_7046,N_7119);
nand U7204 (N_7204,N_7050,N_7036);
xnor U7205 (N_7205,N_7093,N_7008);
nand U7206 (N_7206,N_7055,N_7006);
and U7207 (N_7207,N_7031,N_7034);
nor U7208 (N_7208,N_7008,N_7007);
or U7209 (N_7209,N_7109,N_7100);
and U7210 (N_7210,N_7063,N_7006);
nor U7211 (N_7211,N_7007,N_7059);
or U7212 (N_7212,N_7104,N_7046);
or U7213 (N_7213,N_7050,N_7018);
xnor U7214 (N_7214,N_7099,N_7028);
nor U7215 (N_7215,N_7107,N_7109);
nor U7216 (N_7216,N_7064,N_7086);
xnor U7217 (N_7217,N_7057,N_7047);
nand U7218 (N_7218,N_7038,N_7011);
and U7219 (N_7219,N_7031,N_7071);
nor U7220 (N_7220,N_7011,N_7084);
nand U7221 (N_7221,N_7122,N_7054);
and U7222 (N_7222,N_7064,N_7045);
or U7223 (N_7223,N_7015,N_7082);
and U7224 (N_7224,N_7076,N_7095);
nand U7225 (N_7225,N_7010,N_7110);
and U7226 (N_7226,N_7095,N_7054);
nor U7227 (N_7227,N_7042,N_7054);
or U7228 (N_7228,N_7080,N_7069);
or U7229 (N_7229,N_7080,N_7053);
and U7230 (N_7230,N_7027,N_7017);
nor U7231 (N_7231,N_7097,N_7030);
or U7232 (N_7232,N_7088,N_7079);
nor U7233 (N_7233,N_7051,N_7109);
nand U7234 (N_7234,N_7059,N_7024);
and U7235 (N_7235,N_7056,N_7070);
xor U7236 (N_7236,N_7080,N_7086);
xnor U7237 (N_7237,N_7004,N_7120);
nand U7238 (N_7238,N_7024,N_7049);
and U7239 (N_7239,N_7058,N_7101);
or U7240 (N_7240,N_7015,N_7035);
xor U7241 (N_7241,N_7056,N_7049);
nand U7242 (N_7242,N_7068,N_7011);
and U7243 (N_7243,N_7001,N_7104);
and U7244 (N_7244,N_7105,N_7046);
or U7245 (N_7245,N_7034,N_7083);
nor U7246 (N_7246,N_7046,N_7055);
nor U7247 (N_7247,N_7005,N_7007);
and U7248 (N_7248,N_7000,N_7070);
nor U7249 (N_7249,N_7020,N_7110);
nand U7250 (N_7250,N_7239,N_7151);
nand U7251 (N_7251,N_7242,N_7173);
and U7252 (N_7252,N_7229,N_7194);
xnor U7253 (N_7253,N_7230,N_7231);
nand U7254 (N_7254,N_7244,N_7171);
nor U7255 (N_7255,N_7204,N_7165);
nor U7256 (N_7256,N_7218,N_7129);
or U7257 (N_7257,N_7226,N_7178);
and U7258 (N_7258,N_7128,N_7156);
nor U7259 (N_7259,N_7217,N_7132);
and U7260 (N_7260,N_7130,N_7201);
nor U7261 (N_7261,N_7220,N_7147);
xnor U7262 (N_7262,N_7237,N_7160);
and U7263 (N_7263,N_7248,N_7233);
nand U7264 (N_7264,N_7227,N_7197);
or U7265 (N_7265,N_7145,N_7247);
nand U7266 (N_7266,N_7140,N_7219);
nand U7267 (N_7267,N_7190,N_7174);
and U7268 (N_7268,N_7136,N_7192);
or U7269 (N_7269,N_7170,N_7223);
and U7270 (N_7270,N_7161,N_7141);
and U7271 (N_7271,N_7216,N_7168);
xnor U7272 (N_7272,N_7137,N_7207);
nand U7273 (N_7273,N_7172,N_7222);
nor U7274 (N_7274,N_7184,N_7187);
nor U7275 (N_7275,N_7221,N_7144);
and U7276 (N_7276,N_7238,N_7155);
or U7277 (N_7277,N_7153,N_7143);
and U7278 (N_7278,N_7146,N_7162);
nor U7279 (N_7279,N_7181,N_7131);
or U7280 (N_7280,N_7126,N_7127);
xor U7281 (N_7281,N_7245,N_7240);
nor U7282 (N_7282,N_7182,N_7209);
nand U7283 (N_7283,N_7183,N_7203);
xor U7284 (N_7284,N_7125,N_7166);
or U7285 (N_7285,N_7133,N_7212);
nor U7286 (N_7286,N_7185,N_7224);
nor U7287 (N_7287,N_7234,N_7195);
or U7288 (N_7288,N_7198,N_7193);
and U7289 (N_7289,N_7164,N_7243);
xnor U7290 (N_7290,N_7152,N_7228);
and U7291 (N_7291,N_7169,N_7189);
xnor U7292 (N_7292,N_7236,N_7180);
xnor U7293 (N_7293,N_7232,N_7139);
or U7294 (N_7294,N_7211,N_7138);
and U7295 (N_7295,N_7213,N_7225);
and U7296 (N_7296,N_7191,N_7199);
or U7297 (N_7297,N_7150,N_7135);
nor U7298 (N_7298,N_7246,N_7167);
xor U7299 (N_7299,N_7158,N_7142);
nand U7300 (N_7300,N_7241,N_7175);
nor U7301 (N_7301,N_7159,N_7200);
nand U7302 (N_7302,N_7215,N_7206);
or U7303 (N_7303,N_7179,N_7134);
nor U7304 (N_7304,N_7214,N_7177);
and U7305 (N_7305,N_7163,N_7157);
nand U7306 (N_7306,N_7210,N_7235);
nor U7307 (N_7307,N_7249,N_7205);
or U7308 (N_7308,N_7176,N_7208);
or U7309 (N_7309,N_7149,N_7196);
and U7310 (N_7310,N_7148,N_7202);
and U7311 (N_7311,N_7154,N_7186);
and U7312 (N_7312,N_7188,N_7248);
nand U7313 (N_7313,N_7210,N_7204);
and U7314 (N_7314,N_7132,N_7215);
nand U7315 (N_7315,N_7229,N_7143);
nand U7316 (N_7316,N_7174,N_7165);
and U7317 (N_7317,N_7173,N_7158);
or U7318 (N_7318,N_7209,N_7187);
and U7319 (N_7319,N_7204,N_7143);
nand U7320 (N_7320,N_7209,N_7151);
and U7321 (N_7321,N_7136,N_7210);
xnor U7322 (N_7322,N_7138,N_7161);
or U7323 (N_7323,N_7127,N_7206);
and U7324 (N_7324,N_7232,N_7177);
and U7325 (N_7325,N_7195,N_7224);
and U7326 (N_7326,N_7160,N_7127);
nand U7327 (N_7327,N_7242,N_7150);
nand U7328 (N_7328,N_7184,N_7140);
nor U7329 (N_7329,N_7247,N_7208);
or U7330 (N_7330,N_7127,N_7230);
xnor U7331 (N_7331,N_7176,N_7131);
or U7332 (N_7332,N_7241,N_7240);
or U7333 (N_7333,N_7160,N_7242);
nand U7334 (N_7334,N_7217,N_7177);
nor U7335 (N_7335,N_7180,N_7204);
xnor U7336 (N_7336,N_7158,N_7213);
xor U7337 (N_7337,N_7235,N_7230);
nor U7338 (N_7338,N_7212,N_7189);
and U7339 (N_7339,N_7248,N_7227);
and U7340 (N_7340,N_7176,N_7227);
nor U7341 (N_7341,N_7217,N_7135);
xor U7342 (N_7342,N_7220,N_7170);
xnor U7343 (N_7343,N_7126,N_7173);
nand U7344 (N_7344,N_7246,N_7171);
and U7345 (N_7345,N_7153,N_7195);
and U7346 (N_7346,N_7186,N_7134);
nor U7347 (N_7347,N_7143,N_7242);
nor U7348 (N_7348,N_7240,N_7180);
nand U7349 (N_7349,N_7234,N_7181);
xor U7350 (N_7350,N_7233,N_7153);
or U7351 (N_7351,N_7129,N_7184);
nor U7352 (N_7352,N_7163,N_7236);
xnor U7353 (N_7353,N_7201,N_7220);
or U7354 (N_7354,N_7235,N_7222);
nand U7355 (N_7355,N_7188,N_7212);
nand U7356 (N_7356,N_7139,N_7215);
nor U7357 (N_7357,N_7161,N_7214);
nand U7358 (N_7358,N_7236,N_7137);
or U7359 (N_7359,N_7223,N_7228);
nand U7360 (N_7360,N_7186,N_7213);
and U7361 (N_7361,N_7187,N_7127);
xor U7362 (N_7362,N_7169,N_7180);
nor U7363 (N_7363,N_7231,N_7174);
nor U7364 (N_7364,N_7148,N_7182);
nor U7365 (N_7365,N_7185,N_7234);
nor U7366 (N_7366,N_7131,N_7224);
xor U7367 (N_7367,N_7230,N_7217);
or U7368 (N_7368,N_7202,N_7236);
nor U7369 (N_7369,N_7126,N_7174);
or U7370 (N_7370,N_7131,N_7142);
and U7371 (N_7371,N_7143,N_7176);
or U7372 (N_7372,N_7249,N_7182);
xor U7373 (N_7373,N_7217,N_7141);
nor U7374 (N_7374,N_7249,N_7185);
or U7375 (N_7375,N_7252,N_7286);
or U7376 (N_7376,N_7330,N_7335);
nand U7377 (N_7377,N_7292,N_7271);
and U7378 (N_7378,N_7349,N_7348);
and U7379 (N_7379,N_7284,N_7304);
nor U7380 (N_7380,N_7363,N_7297);
xnor U7381 (N_7381,N_7360,N_7352);
or U7382 (N_7382,N_7298,N_7257);
xor U7383 (N_7383,N_7322,N_7269);
or U7384 (N_7384,N_7255,N_7366);
nor U7385 (N_7385,N_7343,N_7256);
nand U7386 (N_7386,N_7274,N_7287);
nor U7387 (N_7387,N_7361,N_7370);
and U7388 (N_7388,N_7344,N_7268);
and U7389 (N_7389,N_7267,N_7368);
and U7390 (N_7390,N_7356,N_7329);
or U7391 (N_7391,N_7310,N_7263);
xnor U7392 (N_7392,N_7306,N_7296);
or U7393 (N_7393,N_7328,N_7320);
nand U7394 (N_7394,N_7293,N_7357);
xnor U7395 (N_7395,N_7270,N_7290);
or U7396 (N_7396,N_7326,N_7280);
or U7397 (N_7397,N_7325,N_7253);
and U7398 (N_7398,N_7331,N_7313);
xor U7399 (N_7399,N_7303,N_7373);
and U7400 (N_7400,N_7288,N_7333);
nor U7401 (N_7401,N_7334,N_7327);
nand U7402 (N_7402,N_7277,N_7354);
nor U7403 (N_7403,N_7300,N_7314);
and U7404 (N_7404,N_7351,N_7340);
and U7405 (N_7405,N_7346,N_7259);
xor U7406 (N_7406,N_7342,N_7260);
and U7407 (N_7407,N_7347,N_7324);
nand U7408 (N_7408,N_7371,N_7367);
xor U7409 (N_7409,N_7299,N_7285);
or U7410 (N_7410,N_7369,N_7372);
or U7411 (N_7411,N_7359,N_7281);
nor U7412 (N_7412,N_7339,N_7291);
or U7413 (N_7413,N_7266,N_7278);
nand U7414 (N_7414,N_7282,N_7251);
xor U7415 (N_7415,N_7301,N_7350);
or U7416 (N_7416,N_7345,N_7353);
or U7417 (N_7417,N_7258,N_7272);
xnor U7418 (N_7418,N_7355,N_7261);
nor U7419 (N_7419,N_7358,N_7311);
and U7420 (N_7420,N_7283,N_7312);
xor U7421 (N_7421,N_7365,N_7295);
nand U7422 (N_7422,N_7307,N_7294);
or U7423 (N_7423,N_7321,N_7315);
and U7424 (N_7424,N_7289,N_7319);
xnor U7425 (N_7425,N_7374,N_7332);
nand U7426 (N_7426,N_7275,N_7341);
or U7427 (N_7427,N_7276,N_7316);
and U7428 (N_7428,N_7337,N_7250);
xnor U7429 (N_7429,N_7262,N_7338);
nor U7430 (N_7430,N_7308,N_7336);
nand U7431 (N_7431,N_7265,N_7273);
and U7432 (N_7432,N_7309,N_7264);
or U7433 (N_7433,N_7305,N_7362);
nand U7434 (N_7434,N_7302,N_7323);
or U7435 (N_7435,N_7318,N_7279);
or U7436 (N_7436,N_7254,N_7317);
xnor U7437 (N_7437,N_7364,N_7341);
or U7438 (N_7438,N_7359,N_7301);
or U7439 (N_7439,N_7332,N_7355);
and U7440 (N_7440,N_7263,N_7297);
xor U7441 (N_7441,N_7269,N_7321);
and U7442 (N_7442,N_7348,N_7324);
nand U7443 (N_7443,N_7279,N_7255);
nand U7444 (N_7444,N_7318,N_7335);
and U7445 (N_7445,N_7261,N_7336);
nor U7446 (N_7446,N_7251,N_7270);
xor U7447 (N_7447,N_7299,N_7282);
nor U7448 (N_7448,N_7349,N_7309);
or U7449 (N_7449,N_7368,N_7254);
xor U7450 (N_7450,N_7371,N_7368);
nor U7451 (N_7451,N_7273,N_7299);
xor U7452 (N_7452,N_7259,N_7307);
nand U7453 (N_7453,N_7291,N_7318);
and U7454 (N_7454,N_7344,N_7259);
nor U7455 (N_7455,N_7358,N_7300);
or U7456 (N_7456,N_7264,N_7326);
or U7457 (N_7457,N_7316,N_7296);
xor U7458 (N_7458,N_7267,N_7372);
nand U7459 (N_7459,N_7310,N_7363);
xnor U7460 (N_7460,N_7253,N_7299);
or U7461 (N_7461,N_7360,N_7362);
and U7462 (N_7462,N_7358,N_7374);
and U7463 (N_7463,N_7279,N_7344);
or U7464 (N_7464,N_7354,N_7323);
nor U7465 (N_7465,N_7262,N_7318);
nor U7466 (N_7466,N_7312,N_7355);
xor U7467 (N_7467,N_7276,N_7325);
nor U7468 (N_7468,N_7371,N_7337);
xnor U7469 (N_7469,N_7320,N_7342);
and U7470 (N_7470,N_7258,N_7313);
xor U7471 (N_7471,N_7251,N_7345);
nor U7472 (N_7472,N_7342,N_7352);
nor U7473 (N_7473,N_7252,N_7261);
or U7474 (N_7474,N_7323,N_7306);
nor U7475 (N_7475,N_7290,N_7316);
nor U7476 (N_7476,N_7327,N_7332);
or U7477 (N_7477,N_7308,N_7292);
and U7478 (N_7478,N_7336,N_7341);
xor U7479 (N_7479,N_7371,N_7308);
xor U7480 (N_7480,N_7262,N_7304);
and U7481 (N_7481,N_7327,N_7279);
and U7482 (N_7482,N_7265,N_7339);
or U7483 (N_7483,N_7287,N_7277);
xnor U7484 (N_7484,N_7255,N_7321);
or U7485 (N_7485,N_7257,N_7278);
or U7486 (N_7486,N_7315,N_7340);
nor U7487 (N_7487,N_7369,N_7255);
nand U7488 (N_7488,N_7266,N_7370);
and U7489 (N_7489,N_7272,N_7295);
and U7490 (N_7490,N_7303,N_7311);
xnor U7491 (N_7491,N_7280,N_7282);
and U7492 (N_7492,N_7349,N_7316);
or U7493 (N_7493,N_7288,N_7255);
nand U7494 (N_7494,N_7298,N_7348);
or U7495 (N_7495,N_7300,N_7273);
and U7496 (N_7496,N_7324,N_7287);
nand U7497 (N_7497,N_7348,N_7326);
nor U7498 (N_7498,N_7299,N_7303);
or U7499 (N_7499,N_7345,N_7279);
nor U7500 (N_7500,N_7436,N_7424);
or U7501 (N_7501,N_7490,N_7413);
and U7502 (N_7502,N_7399,N_7492);
and U7503 (N_7503,N_7486,N_7402);
or U7504 (N_7504,N_7400,N_7396);
nand U7505 (N_7505,N_7426,N_7385);
nor U7506 (N_7506,N_7473,N_7480);
xnor U7507 (N_7507,N_7420,N_7487);
or U7508 (N_7508,N_7472,N_7414);
or U7509 (N_7509,N_7438,N_7388);
or U7510 (N_7510,N_7491,N_7478);
and U7511 (N_7511,N_7379,N_7457);
nor U7512 (N_7512,N_7409,N_7430);
or U7513 (N_7513,N_7466,N_7483);
nand U7514 (N_7514,N_7471,N_7435);
xor U7515 (N_7515,N_7411,N_7497);
and U7516 (N_7516,N_7493,N_7439);
nor U7517 (N_7517,N_7458,N_7432);
xor U7518 (N_7518,N_7499,N_7383);
or U7519 (N_7519,N_7442,N_7431);
nor U7520 (N_7520,N_7444,N_7421);
nor U7521 (N_7521,N_7474,N_7477);
and U7522 (N_7522,N_7455,N_7453);
or U7523 (N_7523,N_7460,N_7429);
xnor U7524 (N_7524,N_7407,N_7387);
nand U7525 (N_7525,N_7397,N_7498);
xnor U7526 (N_7526,N_7449,N_7494);
or U7527 (N_7527,N_7440,N_7404);
nor U7528 (N_7528,N_7450,N_7376);
and U7529 (N_7529,N_7390,N_7398);
or U7530 (N_7530,N_7456,N_7465);
xnor U7531 (N_7531,N_7467,N_7386);
nor U7532 (N_7532,N_7384,N_7475);
or U7533 (N_7533,N_7375,N_7496);
nand U7534 (N_7534,N_7481,N_7451);
or U7535 (N_7535,N_7415,N_7406);
nand U7536 (N_7536,N_7392,N_7378);
xor U7537 (N_7537,N_7403,N_7470);
xor U7538 (N_7538,N_7462,N_7476);
nor U7539 (N_7539,N_7408,N_7445);
or U7540 (N_7540,N_7464,N_7393);
nand U7541 (N_7541,N_7454,N_7484);
and U7542 (N_7542,N_7437,N_7433);
nand U7543 (N_7543,N_7377,N_7485);
or U7544 (N_7544,N_7419,N_7425);
or U7545 (N_7545,N_7427,N_7482);
and U7546 (N_7546,N_7479,N_7495);
or U7547 (N_7547,N_7428,N_7469);
and U7548 (N_7548,N_7446,N_7423);
or U7549 (N_7549,N_7394,N_7461);
nor U7550 (N_7550,N_7381,N_7418);
nand U7551 (N_7551,N_7463,N_7412);
nand U7552 (N_7552,N_7391,N_7441);
nand U7553 (N_7553,N_7380,N_7459);
xnor U7554 (N_7554,N_7401,N_7422);
and U7555 (N_7555,N_7452,N_7489);
nor U7556 (N_7556,N_7395,N_7417);
and U7557 (N_7557,N_7410,N_7447);
and U7558 (N_7558,N_7405,N_7443);
xnor U7559 (N_7559,N_7416,N_7448);
and U7560 (N_7560,N_7434,N_7389);
or U7561 (N_7561,N_7382,N_7468);
nor U7562 (N_7562,N_7488,N_7456);
and U7563 (N_7563,N_7378,N_7474);
xor U7564 (N_7564,N_7413,N_7387);
and U7565 (N_7565,N_7420,N_7385);
nand U7566 (N_7566,N_7412,N_7466);
nor U7567 (N_7567,N_7412,N_7454);
xor U7568 (N_7568,N_7437,N_7460);
xnor U7569 (N_7569,N_7413,N_7474);
nand U7570 (N_7570,N_7392,N_7474);
nor U7571 (N_7571,N_7492,N_7448);
or U7572 (N_7572,N_7416,N_7459);
nand U7573 (N_7573,N_7406,N_7457);
xor U7574 (N_7574,N_7442,N_7454);
nand U7575 (N_7575,N_7499,N_7412);
nor U7576 (N_7576,N_7436,N_7450);
nand U7577 (N_7577,N_7393,N_7420);
xnor U7578 (N_7578,N_7445,N_7393);
and U7579 (N_7579,N_7451,N_7405);
nand U7580 (N_7580,N_7487,N_7386);
xor U7581 (N_7581,N_7464,N_7489);
xor U7582 (N_7582,N_7495,N_7397);
nand U7583 (N_7583,N_7450,N_7476);
nand U7584 (N_7584,N_7496,N_7442);
or U7585 (N_7585,N_7425,N_7383);
nand U7586 (N_7586,N_7455,N_7486);
nor U7587 (N_7587,N_7429,N_7499);
or U7588 (N_7588,N_7383,N_7420);
and U7589 (N_7589,N_7457,N_7439);
nand U7590 (N_7590,N_7455,N_7413);
nor U7591 (N_7591,N_7409,N_7451);
nand U7592 (N_7592,N_7483,N_7412);
nand U7593 (N_7593,N_7473,N_7462);
or U7594 (N_7594,N_7473,N_7481);
or U7595 (N_7595,N_7432,N_7491);
and U7596 (N_7596,N_7404,N_7401);
and U7597 (N_7597,N_7482,N_7407);
nor U7598 (N_7598,N_7421,N_7488);
nand U7599 (N_7599,N_7486,N_7487);
nor U7600 (N_7600,N_7407,N_7472);
nand U7601 (N_7601,N_7481,N_7478);
xnor U7602 (N_7602,N_7439,N_7376);
nor U7603 (N_7603,N_7387,N_7494);
nor U7604 (N_7604,N_7386,N_7446);
xnor U7605 (N_7605,N_7408,N_7470);
or U7606 (N_7606,N_7487,N_7494);
xor U7607 (N_7607,N_7427,N_7451);
or U7608 (N_7608,N_7451,N_7425);
nor U7609 (N_7609,N_7495,N_7399);
or U7610 (N_7610,N_7451,N_7492);
or U7611 (N_7611,N_7399,N_7381);
or U7612 (N_7612,N_7455,N_7399);
nand U7613 (N_7613,N_7447,N_7431);
nor U7614 (N_7614,N_7494,N_7376);
nor U7615 (N_7615,N_7430,N_7477);
xnor U7616 (N_7616,N_7450,N_7383);
and U7617 (N_7617,N_7425,N_7435);
nand U7618 (N_7618,N_7475,N_7404);
xor U7619 (N_7619,N_7460,N_7377);
nand U7620 (N_7620,N_7391,N_7497);
xnor U7621 (N_7621,N_7393,N_7383);
xor U7622 (N_7622,N_7442,N_7497);
nand U7623 (N_7623,N_7409,N_7444);
nand U7624 (N_7624,N_7461,N_7410);
xnor U7625 (N_7625,N_7528,N_7501);
nand U7626 (N_7626,N_7504,N_7613);
nor U7627 (N_7627,N_7596,N_7529);
and U7628 (N_7628,N_7589,N_7610);
or U7629 (N_7629,N_7520,N_7536);
xnor U7630 (N_7630,N_7604,N_7560);
and U7631 (N_7631,N_7518,N_7576);
xnor U7632 (N_7632,N_7592,N_7551);
nor U7633 (N_7633,N_7523,N_7575);
and U7634 (N_7634,N_7602,N_7619);
nor U7635 (N_7635,N_7597,N_7525);
or U7636 (N_7636,N_7583,N_7508);
or U7637 (N_7637,N_7517,N_7535);
nand U7638 (N_7638,N_7611,N_7624);
nand U7639 (N_7639,N_7516,N_7585);
xor U7640 (N_7640,N_7569,N_7537);
and U7641 (N_7641,N_7521,N_7621);
or U7642 (N_7642,N_7522,N_7500);
nor U7643 (N_7643,N_7590,N_7614);
xnor U7644 (N_7644,N_7538,N_7507);
xnor U7645 (N_7645,N_7598,N_7509);
nand U7646 (N_7646,N_7513,N_7591);
nand U7647 (N_7647,N_7555,N_7616);
nand U7648 (N_7648,N_7570,N_7548);
or U7649 (N_7649,N_7600,N_7549);
nor U7650 (N_7650,N_7587,N_7505);
and U7651 (N_7651,N_7568,N_7622);
nor U7652 (N_7652,N_7553,N_7562);
nor U7653 (N_7653,N_7581,N_7558);
nor U7654 (N_7654,N_7543,N_7612);
or U7655 (N_7655,N_7615,N_7554);
and U7656 (N_7656,N_7510,N_7512);
nor U7657 (N_7657,N_7546,N_7605);
nand U7658 (N_7658,N_7544,N_7606);
and U7659 (N_7659,N_7565,N_7524);
and U7660 (N_7660,N_7533,N_7593);
xor U7661 (N_7661,N_7572,N_7577);
or U7662 (N_7662,N_7563,N_7620);
xnor U7663 (N_7663,N_7511,N_7540);
or U7664 (N_7664,N_7547,N_7567);
and U7665 (N_7665,N_7519,N_7515);
nor U7666 (N_7666,N_7566,N_7617);
xor U7667 (N_7667,N_7545,N_7618);
nand U7668 (N_7668,N_7503,N_7582);
xnor U7669 (N_7669,N_7571,N_7608);
and U7670 (N_7670,N_7601,N_7603);
and U7671 (N_7671,N_7561,N_7623);
xnor U7672 (N_7672,N_7539,N_7574);
nand U7673 (N_7673,N_7530,N_7552);
and U7674 (N_7674,N_7586,N_7502);
nand U7675 (N_7675,N_7557,N_7526);
nor U7676 (N_7676,N_7534,N_7573);
and U7677 (N_7677,N_7514,N_7607);
xnor U7678 (N_7678,N_7541,N_7588);
nor U7679 (N_7679,N_7506,N_7532);
nor U7680 (N_7680,N_7527,N_7578);
or U7681 (N_7681,N_7564,N_7595);
xor U7682 (N_7682,N_7550,N_7542);
xor U7683 (N_7683,N_7579,N_7609);
or U7684 (N_7684,N_7580,N_7559);
nor U7685 (N_7685,N_7584,N_7556);
nor U7686 (N_7686,N_7531,N_7594);
or U7687 (N_7687,N_7599,N_7522);
or U7688 (N_7688,N_7590,N_7617);
nand U7689 (N_7689,N_7503,N_7520);
nor U7690 (N_7690,N_7534,N_7568);
nand U7691 (N_7691,N_7544,N_7552);
nor U7692 (N_7692,N_7550,N_7611);
nand U7693 (N_7693,N_7578,N_7579);
nand U7694 (N_7694,N_7586,N_7618);
nor U7695 (N_7695,N_7515,N_7590);
nor U7696 (N_7696,N_7555,N_7539);
and U7697 (N_7697,N_7623,N_7624);
nor U7698 (N_7698,N_7607,N_7581);
and U7699 (N_7699,N_7606,N_7527);
or U7700 (N_7700,N_7577,N_7583);
xnor U7701 (N_7701,N_7595,N_7532);
xnor U7702 (N_7702,N_7568,N_7536);
and U7703 (N_7703,N_7562,N_7518);
nand U7704 (N_7704,N_7551,N_7589);
or U7705 (N_7705,N_7531,N_7617);
nor U7706 (N_7706,N_7511,N_7504);
xor U7707 (N_7707,N_7558,N_7579);
xnor U7708 (N_7708,N_7537,N_7579);
nand U7709 (N_7709,N_7539,N_7580);
and U7710 (N_7710,N_7598,N_7548);
nand U7711 (N_7711,N_7569,N_7579);
nand U7712 (N_7712,N_7532,N_7509);
and U7713 (N_7713,N_7508,N_7541);
nand U7714 (N_7714,N_7567,N_7612);
and U7715 (N_7715,N_7566,N_7606);
or U7716 (N_7716,N_7522,N_7514);
or U7717 (N_7717,N_7593,N_7557);
xor U7718 (N_7718,N_7571,N_7543);
and U7719 (N_7719,N_7510,N_7558);
nor U7720 (N_7720,N_7544,N_7506);
xor U7721 (N_7721,N_7578,N_7565);
xor U7722 (N_7722,N_7592,N_7536);
or U7723 (N_7723,N_7558,N_7617);
xor U7724 (N_7724,N_7540,N_7544);
nor U7725 (N_7725,N_7623,N_7533);
and U7726 (N_7726,N_7611,N_7573);
xnor U7727 (N_7727,N_7515,N_7511);
or U7728 (N_7728,N_7532,N_7621);
and U7729 (N_7729,N_7569,N_7614);
and U7730 (N_7730,N_7545,N_7590);
nand U7731 (N_7731,N_7528,N_7527);
or U7732 (N_7732,N_7622,N_7588);
xnor U7733 (N_7733,N_7505,N_7543);
nand U7734 (N_7734,N_7543,N_7561);
xnor U7735 (N_7735,N_7608,N_7554);
or U7736 (N_7736,N_7564,N_7558);
xnor U7737 (N_7737,N_7600,N_7545);
and U7738 (N_7738,N_7578,N_7575);
nand U7739 (N_7739,N_7546,N_7573);
and U7740 (N_7740,N_7557,N_7545);
xnor U7741 (N_7741,N_7515,N_7565);
xnor U7742 (N_7742,N_7621,N_7587);
xor U7743 (N_7743,N_7520,N_7602);
or U7744 (N_7744,N_7526,N_7542);
or U7745 (N_7745,N_7538,N_7612);
or U7746 (N_7746,N_7599,N_7533);
or U7747 (N_7747,N_7522,N_7502);
or U7748 (N_7748,N_7607,N_7559);
nand U7749 (N_7749,N_7543,N_7526);
or U7750 (N_7750,N_7709,N_7667);
nand U7751 (N_7751,N_7661,N_7645);
nor U7752 (N_7752,N_7672,N_7713);
nand U7753 (N_7753,N_7666,N_7731);
nand U7754 (N_7754,N_7714,N_7735);
or U7755 (N_7755,N_7649,N_7700);
nor U7756 (N_7756,N_7745,N_7670);
or U7757 (N_7757,N_7646,N_7728);
xnor U7758 (N_7758,N_7685,N_7648);
or U7759 (N_7759,N_7651,N_7638);
or U7760 (N_7760,N_7725,N_7699);
nor U7761 (N_7761,N_7657,N_7695);
nand U7762 (N_7762,N_7629,N_7655);
nor U7763 (N_7763,N_7718,N_7644);
xnor U7764 (N_7764,N_7634,N_7710);
or U7765 (N_7765,N_7664,N_7741);
nor U7766 (N_7766,N_7678,N_7717);
and U7767 (N_7767,N_7688,N_7631);
xor U7768 (N_7768,N_7673,N_7668);
nand U7769 (N_7769,N_7722,N_7641);
nand U7770 (N_7770,N_7737,N_7742);
or U7771 (N_7771,N_7703,N_7652);
nor U7772 (N_7772,N_7724,N_7704);
or U7773 (N_7773,N_7654,N_7702);
and U7774 (N_7774,N_7719,N_7708);
nand U7775 (N_7775,N_7687,N_7726);
and U7776 (N_7776,N_7686,N_7697);
nor U7777 (N_7777,N_7716,N_7739);
nor U7778 (N_7778,N_7749,N_7727);
and U7779 (N_7779,N_7663,N_7658);
or U7780 (N_7780,N_7676,N_7682);
xnor U7781 (N_7781,N_7690,N_7626);
nand U7782 (N_7782,N_7642,N_7694);
and U7783 (N_7783,N_7691,N_7689);
and U7784 (N_7784,N_7732,N_7677);
nand U7785 (N_7785,N_7692,N_7653);
nand U7786 (N_7786,N_7679,N_7684);
or U7787 (N_7787,N_7660,N_7643);
nand U7788 (N_7788,N_7711,N_7681);
xor U7789 (N_7789,N_7705,N_7665);
or U7790 (N_7790,N_7747,N_7656);
nand U7791 (N_7791,N_7712,N_7733);
xnor U7792 (N_7792,N_7639,N_7693);
or U7793 (N_7793,N_7723,N_7637);
or U7794 (N_7794,N_7650,N_7630);
or U7795 (N_7795,N_7706,N_7627);
xor U7796 (N_7796,N_7736,N_7659);
and U7797 (N_7797,N_7698,N_7720);
nand U7798 (N_7798,N_7635,N_7715);
nor U7799 (N_7799,N_7740,N_7674);
nand U7800 (N_7800,N_7662,N_7738);
nor U7801 (N_7801,N_7707,N_7683);
and U7802 (N_7802,N_7636,N_7744);
or U7803 (N_7803,N_7721,N_7640);
and U7804 (N_7804,N_7680,N_7746);
nor U7805 (N_7805,N_7729,N_7632);
nor U7806 (N_7806,N_7743,N_7734);
and U7807 (N_7807,N_7633,N_7696);
and U7808 (N_7808,N_7671,N_7647);
xor U7809 (N_7809,N_7675,N_7701);
xnor U7810 (N_7810,N_7628,N_7625);
nor U7811 (N_7811,N_7730,N_7748);
and U7812 (N_7812,N_7669,N_7660);
or U7813 (N_7813,N_7639,N_7670);
nor U7814 (N_7814,N_7721,N_7706);
nor U7815 (N_7815,N_7723,N_7683);
or U7816 (N_7816,N_7657,N_7639);
xor U7817 (N_7817,N_7645,N_7634);
xor U7818 (N_7818,N_7654,N_7664);
or U7819 (N_7819,N_7696,N_7692);
xnor U7820 (N_7820,N_7713,N_7642);
or U7821 (N_7821,N_7633,N_7671);
and U7822 (N_7822,N_7656,N_7717);
nand U7823 (N_7823,N_7632,N_7683);
nor U7824 (N_7824,N_7685,N_7642);
nor U7825 (N_7825,N_7648,N_7743);
nor U7826 (N_7826,N_7729,N_7660);
nor U7827 (N_7827,N_7658,N_7666);
nor U7828 (N_7828,N_7692,N_7670);
or U7829 (N_7829,N_7658,N_7717);
and U7830 (N_7830,N_7686,N_7656);
nor U7831 (N_7831,N_7745,N_7719);
xor U7832 (N_7832,N_7670,N_7746);
xor U7833 (N_7833,N_7701,N_7711);
xnor U7834 (N_7834,N_7653,N_7721);
and U7835 (N_7835,N_7707,N_7686);
nor U7836 (N_7836,N_7659,N_7726);
or U7837 (N_7837,N_7676,N_7731);
xnor U7838 (N_7838,N_7647,N_7711);
nor U7839 (N_7839,N_7746,N_7634);
and U7840 (N_7840,N_7645,N_7699);
nand U7841 (N_7841,N_7717,N_7729);
and U7842 (N_7842,N_7736,N_7747);
or U7843 (N_7843,N_7730,N_7720);
nor U7844 (N_7844,N_7684,N_7656);
nand U7845 (N_7845,N_7659,N_7740);
and U7846 (N_7846,N_7724,N_7684);
and U7847 (N_7847,N_7733,N_7672);
xnor U7848 (N_7848,N_7674,N_7713);
nand U7849 (N_7849,N_7665,N_7650);
nor U7850 (N_7850,N_7659,N_7634);
and U7851 (N_7851,N_7666,N_7631);
nor U7852 (N_7852,N_7691,N_7663);
and U7853 (N_7853,N_7681,N_7677);
nand U7854 (N_7854,N_7629,N_7735);
nand U7855 (N_7855,N_7683,N_7656);
nand U7856 (N_7856,N_7653,N_7665);
nand U7857 (N_7857,N_7664,N_7631);
and U7858 (N_7858,N_7712,N_7732);
nand U7859 (N_7859,N_7734,N_7674);
nand U7860 (N_7860,N_7677,N_7679);
xnor U7861 (N_7861,N_7630,N_7671);
nor U7862 (N_7862,N_7629,N_7747);
xor U7863 (N_7863,N_7676,N_7679);
nor U7864 (N_7864,N_7742,N_7679);
and U7865 (N_7865,N_7657,N_7686);
or U7866 (N_7866,N_7658,N_7724);
nor U7867 (N_7867,N_7701,N_7632);
xor U7868 (N_7868,N_7749,N_7743);
and U7869 (N_7869,N_7653,N_7690);
nand U7870 (N_7870,N_7693,N_7665);
xor U7871 (N_7871,N_7704,N_7691);
nand U7872 (N_7872,N_7689,N_7704);
and U7873 (N_7873,N_7659,N_7663);
nor U7874 (N_7874,N_7702,N_7696);
or U7875 (N_7875,N_7759,N_7751);
and U7876 (N_7876,N_7866,N_7811);
or U7877 (N_7877,N_7753,N_7874);
nor U7878 (N_7878,N_7826,N_7834);
and U7879 (N_7879,N_7858,N_7755);
xnor U7880 (N_7880,N_7768,N_7829);
xor U7881 (N_7881,N_7788,N_7773);
nor U7882 (N_7882,N_7842,N_7831);
and U7883 (N_7883,N_7765,N_7841);
xnor U7884 (N_7884,N_7793,N_7849);
xnor U7885 (N_7885,N_7861,N_7810);
xnor U7886 (N_7886,N_7830,N_7776);
xnor U7887 (N_7887,N_7848,N_7772);
nor U7888 (N_7888,N_7795,N_7813);
nor U7889 (N_7889,N_7868,N_7796);
or U7890 (N_7890,N_7856,N_7786);
or U7891 (N_7891,N_7843,N_7869);
and U7892 (N_7892,N_7802,N_7803);
or U7893 (N_7893,N_7844,N_7839);
and U7894 (N_7894,N_7754,N_7764);
or U7895 (N_7895,N_7867,N_7827);
nor U7896 (N_7896,N_7758,N_7791);
nor U7897 (N_7897,N_7770,N_7860);
xor U7898 (N_7898,N_7821,N_7822);
nor U7899 (N_7899,N_7823,N_7854);
nor U7900 (N_7900,N_7851,N_7815);
or U7901 (N_7901,N_7846,N_7852);
nand U7902 (N_7902,N_7807,N_7820);
nand U7903 (N_7903,N_7836,N_7814);
nor U7904 (N_7904,N_7799,N_7789);
xnor U7905 (N_7905,N_7857,N_7855);
and U7906 (N_7906,N_7862,N_7804);
or U7907 (N_7907,N_7805,N_7824);
nor U7908 (N_7908,N_7850,N_7840);
and U7909 (N_7909,N_7864,N_7787);
nor U7910 (N_7910,N_7792,N_7812);
nor U7911 (N_7911,N_7769,N_7817);
or U7912 (N_7912,N_7835,N_7816);
nor U7913 (N_7913,N_7870,N_7771);
or U7914 (N_7914,N_7800,N_7766);
nor U7915 (N_7915,N_7794,N_7845);
xor U7916 (N_7916,N_7853,N_7798);
or U7917 (N_7917,N_7801,N_7762);
and U7918 (N_7918,N_7847,N_7782);
nand U7919 (N_7919,N_7763,N_7828);
or U7920 (N_7920,N_7760,N_7777);
xnor U7921 (N_7921,N_7832,N_7781);
xnor U7922 (N_7922,N_7797,N_7825);
or U7923 (N_7923,N_7784,N_7750);
nand U7924 (N_7924,N_7863,N_7757);
xor U7925 (N_7925,N_7790,N_7774);
nor U7926 (N_7926,N_7838,N_7785);
xnor U7927 (N_7927,N_7752,N_7833);
and U7928 (N_7928,N_7780,N_7767);
and U7929 (N_7929,N_7775,N_7865);
nand U7930 (N_7930,N_7808,N_7859);
or U7931 (N_7931,N_7818,N_7873);
nand U7932 (N_7932,N_7809,N_7779);
and U7933 (N_7933,N_7778,N_7871);
or U7934 (N_7934,N_7837,N_7783);
xor U7935 (N_7935,N_7806,N_7756);
nand U7936 (N_7936,N_7761,N_7819);
and U7937 (N_7937,N_7872,N_7861);
nand U7938 (N_7938,N_7764,N_7816);
xor U7939 (N_7939,N_7816,N_7821);
nor U7940 (N_7940,N_7795,N_7796);
xor U7941 (N_7941,N_7753,N_7805);
and U7942 (N_7942,N_7806,N_7797);
xnor U7943 (N_7943,N_7856,N_7845);
xnor U7944 (N_7944,N_7757,N_7815);
xor U7945 (N_7945,N_7859,N_7837);
or U7946 (N_7946,N_7805,N_7833);
nor U7947 (N_7947,N_7750,N_7825);
nand U7948 (N_7948,N_7796,N_7870);
nor U7949 (N_7949,N_7750,N_7792);
and U7950 (N_7950,N_7859,N_7858);
and U7951 (N_7951,N_7834,N_7844);
xnor U7952 (N_7952,N_7812,N_7837);
xor U7953 (N_7953,N_7760,N_7752);
xnor U7954 (N_7954,N_7782,N_7850);
and U7955 (N_7955,N_7849,N_7842);
or U7956 (N_7956,N_7798,N_7768);
or U7957 (N_7957,N_7853,N_7846);
nand U7958 (N_7958,N_7791,N_7752);
and U7959 (N_7959,N_7758,N_7785);
and U7960 (N_7960,N_7861,N_7753);
or U7961 (N_7961,N_7810,N_7843);
or U7962 (N_7962,N_7855,N_7870);
and U7963 (N_7963,N_7822,N_7817);
nor U7964 (N_7964,N_7824,N_7851);
nor U7965 (N_7965,N_7823,N_7874);
nor U7966 (N_7966,N_7755,N_7751);
nand U7967 (N_7967,N_7847,N_7833);
or U7968 (N_7968,N_7789,N_7812);
or U7969 (N_7969,N_7801,N_7796);
nand U7970 (N_7970,N_7756,N_7851);
and U7971 (N_7971,N_7851,N_7862);
nand U7972 (N_7972,N_7819,N_7845);
nor U7973 (N_7973,N_7752,N_7827);
and U7974 (N_7974,N_7822,N_7802);
or U7975 (N_7975,N_7769,N_7853);
nand U7976 (N_7976,N_7824,N_7791);
nand U7977 (N_7977,N_7757,N_7752);
nor U7978 (N_7978,N_7858,N_7851);
xnor U7979 (N_7979,N_7777,N_7765);
nand U7980 (N_7980,N_7835,N_7772);
or U7981 (N_7981,N_7797,N_7789);
nor U7982 (N_7982,N_7828,N_7764);
xor U7983 (N_7983,N_7837,N_7842);
nand U7984 (N_7984,N_7761,N_7769);
nor U7985 (N_7985,N_7771,N_7861);
nand U7986 (N_7986,N_7814,N_7793);
nor U7987 (N_7987,N_7760,N_7792);
xor U7988 (N_7988,N_7821,N_7870);
or U7989 (N_7989,N_7819,N_7791);
or U7990 (N_7990,N_7834,N_7835);
nor U7991 (N_7991,N_7782,N_7834);
nor U7992 (N_7992,N_7759,N_7819);
and U7993 (N_7993,N_7796,N_7822);
and U7994 (N_7994,N_7772,N_7854);
nand U7995 (N_7995,N_7826,N_7862);
or U7996 (N_7996,N_7830,N_7846);
nor U7997 (N_7997,N_7834,N_7855);
nor U7998 (N_7998,N_7802,N_7798);
nor U7999 (N_7999,N_7864,N_7846);
or U8000 (N_8000,N_7943,N_7973);
nor U8001 (N_8001,N_7900,N_7894);
xnor U8002 (N_8002,N_7998,N_7954);
nor U8003 (N_8003,N_7968,N_7901);
and U8004 (N_8004,N_7982,N_7990);
nand U8005 (N_8005,N_7893,N_7922);
and U8006 (N_8006,N_7975,N_7963);
or U8007 (N_8007,N_7936,N_7976);
nor U8008 (N_8008,N_7918,N_7925);
xor U8009 (N_8009,N_7964,N_7938);
or U8010 (N_8010,N_7881,N_7940);
and U8011 (N_8011,N_7986,N_7890);
nor U8012 (N_8012,N_7930,N_7927);
xor U8013 (N_8013,N_7958,N_7966);
nor U8014 (N_8014,N_7993,N_7935);
xnor U8015 (N_8015,N_7889,N_7908);
nand U8016 (N_8016,N_7884,N_7933);
or U8017 (N_8017,N_7997,N_7952);
and U8018 (N_8018,N_7907,N_7981);
and U8019 (N_8019,N_7920,N_7934);
or U8020 (N_8020,N_7899,N_7882);
nand U8021 (N_8021,N_7953,N_7887);
or U8022 (N_8022,N_7992,N_7942);
and U8023 (N_8023,N_7886,N_7983);
xor U8024 (N_8024,N_7949,N_7959);
or U8025 (N_8025,N_7980,N_7923);
nand U8026 (N_8026,N_7909,N_7921);
and U8027 (N_8027,N_7906,N_7944);
nor U8028 (N_8028,N_7913,N_7891);
or U8029 (N_8029,N_7994,N_7883);
nor U8030 (N_8030,N_7941,N_7965);
xor U8031 (N_8031,N_7987,N_7905);
xnor U8032 (N_8032,N_7903,N_7957);
or U8033 (N_8033,N_7946,N_7974);
nand U8034 (N_8034,N_7879,N_7904);
or U8035 (N_8035,N_7996,N_7960);
and U8036 (N_8036,N_7924,N_7915);
or U8037 (N_8037,N_7937,N_7948);
nor U8038 (N_8038,N_7977,N_7876);
nor U8039 (N_8039,N_7911,N_7931);
xor U8040 (N_8040,N_7962,N_7945);
or U8041 (N_8041,N_7912,N_7979);
or U8042 (N_8042,N_7929,N_7897);
or U8043 (N_8043,N_7932,N_7951);
or U8044 (N_8044,N_7999,N_7888);
xnor U8045 (N_8045,N_7895,N_7961);
and U8046 (N_8046,N_7875,N_7939);
or U8047 (N_8047,N_7956,N_7919);
and U8048 (N_8048,N_7896,N_7878);
xor U8049 (N_8049,N_7910,N_7969);
nand U8050 (N_8050,N_7988,N_7955);
nor U8051 (N_8051,N_7902,N_7892);
xor U8052 (N_8052,N_7880,N_7967);
or U8053 (N_8053,N_7950,N_7995);
and U8054 (N_8054,N_7985,N_7898);
and U8055 (N_8055,N_7947,N_7970);
nor U8056 (N_8056,N_7991,N_7928);
nand U8057 (N_8057,N_7916,N_7971);
and U8058 (N_8058,N_7978,N_7926);
nor U8059 (N_8059,N_7917,N_7984);
xnor U8060 (N_8060,N_7972,N_7885);
nor U8061 (N_8061,N_7877,N_7914);
and U8062 (N_8062,N_7989,N_7950);
and U8063 (N_8063,N_7931,N_7898);
nor U8064 (N_8064,N_7933,N_7892);
or U8065 (N_8065,N_7932,N_7877);
nand U8066 (N_8066,N_7979,N_7968);
and U8067 (N_8067,N_7986,N_7903);
or U8068 (N_8068,N_7988,N_7966);
or U8069 (N_8069,N_7964,N_7934);
nand U8070 (N_8070,N_7947,N_7926);
and U8071 (N_8071,N_7971,N_7958);
and U8072 (N_8072,N_7976,N_7878);
nor U8073 (N_8073,N_7900,N_7891);
nand U8074 (N_8074,N_7898,N_7882);
or U8075 (N_8075,N_7938,N_7982);
xnor U8076 (N_8076,N_7889,N_7986);
nor U8077 (N_8077,N_7926,N_7946);
nor U8078 (N_8078,N_7914,N_7950);
nor U8079 (N_8079,N_7977,N_7985);
and U8080 (N_8080,N_7983,N_7885);
nor U8081 (N_8081,N_7967,N_7935);
and U8082 (N_8082,N_7924,N_7965);
xor U8083 (N_8083,N_7993,N_7879);
and U8084 (N_8084,N_7899,N_7939);
nor U8085 (N_8085,N_7924,N_7952);
nand U8086 (N_8086,N_7891,N_7935);
xnor U8087 (N_8087,N_7946,N_7891);
nor U8088 (N_8088,N_7977,N_7944);
nand U8089 (N_8089,N_7935,N_7978);
xnor U8090 (N_8090,N_7939,N_7993);
xor U8091 (N_8091,N_7977,N_7900);
nand U8092 (N_8092,N_7980,N_7965);
or U8093 (N_8093,N_7899,N_7958);
or U8094 (N_8094,N_7938,N_7923);
xor U8095 (N_8095,N_7971,N_7986);
nand U8096 (N_8096,N_7932,N_7999);
nand U8097 (N_8097,N_7911,N_7882);
or U8098 (N_8098,N_7900,N_7881);
and U8099 (N_8099,N_7984,N_7902);
nor U8100 (N_8100,N_7910,N_7933);
and U8101 (N_8101,N_7981,N_7875);
and U8102 (N_8102,N_7921,N_7949);
nand U8103 (N_8103,N_7922,N_7911);
or U8104 (N_8104,N_7877,N_7906);
nand U8105 (N_8105,N_7890,N_7959);
nor U8106 (N_8106,N_7985,N_7946);
nor U8107 (N_8107,N_7993,N_7969);
nor U8108 (N_8108,N_7998,N_7946);
and U8109 (N_8109,N_7945,N_7995);
xor U8110 (N_8110,N_7976,N_7882);
or U8111 (N_8111,N_7971,N_7951);
and U8112 (N_8112,N_7897,N_7938);
nand U8113 (N_8113,N_7945,N_7982);
or U8114 (N_8114,N_7886,N_7883);
and U8115 (N_8115,N_7923,N_7915);
and U8116 (N_8116,N_7922,N_7993);
or U8117 (N_8117,N_7957,N_7938);
and U8118 (N_8118,N_7971,N_7966);
or U8119 (N_8119,N_7996,N_7881);
xnor U8120 (N_8120,N_7957,N_7879);
nor U8121 (N_8121,N_7888,N_7899);
and U8122 (N_8122,N_7931,N_7881);
or U8123 (N_8123,N_7980,N_7921);
and U8124 (N_8124,N_7994,N_7951);
xor U8125 (N_8125,N_8080,N_8051);
or U8126 (N_8126,N_8019,N_8123);
nand U8127 (N_8127,N_8086,N_8020);
nor U8128 (N_8128,N_8031,N_8069);
or U8129 (N_8129,N_8038,N_8098);
nand U8130 (N_8130,N_8057,N_8044);
xnor U8131 (N_8131,N_8056,N_8091);
or U8132 (N_8132,N_8035,N_8111);
xor U8133 (N_8133,N_8063,N_8117);
nor U8134 (N_8134,N_8062,N_8054);
nand U8135 (N_8135,N_8087,N_8033);
and U8136 (N_8136,N_8079,N_8088);
nor U8137 (N_8137,N_8042,N_8028);
nand U8138 (N_8138,N_8082,N_8084);
or U8139 (N_8139,N_8094,N_8003);
or U8140 (N_8140,N_8099,N_8022);
nand U8141 (N_8141,N_8012,N_8093);
and U8142 (N_8142,N_8114,N_8004);
or U8143 (N_8143,N_8014,N_8050);
and U8144 (N_8144,N_8041,N_8073);
nor U8145 (N_8145,N_8013,N_8018);
nor U8146 (N_8146,N_8124,N_8053);
or U8147 (N_8147,N_8074,N_8016);
or U8148 (N_8148,N_8008,N_8120);
xor U8149 (N_8149,N_8011,N_8045);
nand U8150 (N_8150,N_8026,N_8059);
or U8151 (N_8151,N_8017,N_8009);
nor U8152 (N_8152,N_8113,N_8060);
nand U8153 (N_8153,N_8110,N_8036);
xnor U8154 (N_8154,N_8048,N_8058);
and U8155 (N_8155,N_8081,N_8005);
or U8156 (N_8156,N_8000,N_8105);
and U8157 (N_8157,N_8116,N_8040);
or U8158 (N_8158,N_8072,N_8039);
and U8159 (N_8159,N_8108,N_8052);
and U8160 (N_8160,N_8015,N_8100);
nand U8161 (N_8161,N_8029,N_8067);
and U8162 (N_8162,N_8066,N_8001);
xnor U8163 (N_8163,N_8043,N_8024);
or U8164 (N_8164,N_8119,N_8075);
and U8165 (N_8165,N_8092,N_8077);
nand U8166 (N_8166,N_8032,N_8021);
nor U8167 (N_8167,N_8025,N_8096);
nand U8168 (N_8168,N_8007,N_8061);
and U8169 (N_8169,N_8101,N_8102);
nor U8170 (N_8170,N_8112,N_8064);
xor U8171 (N_8171,N_8010,N_8106);
nand U8172 (N_8172,N_8115,N_8070);
xnor U8173 (N_8173,N_8095,N_8037);
and U8174 (N_8174,N_8055,N_8089);
nor U8175 (N_8175,N_8006,N_8085);
nand U8176 (N_8176,N_8122,N_8046);
xnor U8177 (N_8177,N_8027,N_8047);
nor U8178 (N_8178,N_8083,N_8107);
or U8179 (N_8179,N_8049,N_8118);
xnor U8180 (N_8180,N_8076,N_8109);
nor U8181 (N_8181,N_8002,N_8121);
xor U8182 (N_8182,N_8090,N_8071);
nand U8183 (N_8183,N_8097,N_8068);
xor U8184 (N_8184,N_8065,N_8023);
and U8185 (N_8185,N_8030,N_8103);
and U8186 (N_8186,N_8078,N_8104);
xnor U8187 (N_8187,N_8034,N_8116);
or U8188 (N_8188,N_8058,N_8091);
xnor U8189 (N_8189,N_8082,N_8046);
nor U8190 (N_8190,N_8036,N_8055);
xnor U8191 (N_8191,N_8084,N_8045);
nand U8192 (N_8192,N_8119,N_8025);
xnor U8193 (N_8193,N_8076,N_8043);
xnor U8194 (N_8194,N_8009,N_8116);
xnor U8195 (N_8195,N_8097,N_8072);
xnor U8196 (N_8196,N_8060,N_8015);
nand U8197 (N_8197,N_8005,N_8122);
xor U8198 (N_8198,N_8009,N_8121);
or U8199 (N_8199,N_8071,N_8108);
and U8200 (N_8200,N_8001,N_8062);
nand U8201 (N_8201,N_8081,N_8087);
nor U8202 (N_8202,N_8082,N_8070);
or U8203 (N_8203,N_8032,N_8117);
and U8204 (N_8204,N_8034,N_8035);
and U8205 (N_8205,N_8022,N_8024);
nor U8206 (N_8206,N_8059,N_8088);
or U8207 (N_8207,N_8117,N_8026);
or U8208 (N_8208,N_8096,N_8094);
or U8209 (N_8209,N_8063,N_8084);
xnor U8210 (N_8210,N_8111,N_8051);
xor U8211 (N_8211,N_8001,N_8064);
xor U8212 (N_8212,N_8048,N_8037);
nor U8213 (N_8213,N_8030,N_8118);
xnor U8214 (N_8214,N_8093,N_8017);
nand U8215 (N_8215,N_8078,N_8047);
or U8216 (N_8216,N_8055,N_8097);
or U8217 (N_8217,N_8060,N_8123);
xor U8218 (N_8218,N_8117,N_8111);
or U8219 (N_8219,N_8005,N_8021);
nor U8220 (N_8220,N_8023,N_8046);
nand U8221 (N_8221,N_8032,N_8033);
or U8222 (N_8222,N_8038,N_8063);
and U8223 (N_8223,N_8004,N_8068);
and U8224 (N_8224,N_8112,N_8099);
or U8225 (N_8225,N_8097,N_8109);
nand U8226 (N_8226,N_8084,N_8079);
xor U8227 (N_8227,N_8038,N_8078);
nor U8228 (N_8228,N_8074,N_8099);
or U8229 (N_8229,N_8034,N_8012);
and U8230 (N_8230,N_8057,N_8116);
nor U8231 (N_8231,N_8052,N_8120);
or U8232 (N_8232,N_8094,N_8075);
xor U8233 (N_8233,N_8030,N_8013);
xor U8234 (N_8234,N_8082,N_8008);
nand U8235 (N_8235,N_8050,N_8039);
or U8236 (N_8236,N_8041,N_8007);
nand U8237 (N_8237,N_8077,N_8101);
nor U8238 (N_8238,N_8018,N_8054);
and U8239 (N_8239,N_8037,N_8035);
and U8240 (N_8240,N_8089,N_8042);
nand U8241 (N_8241,N_8052,N_8090);
or U8242 (N_8242,N_8082,N_8104);
or U8243 (N_8243,N_8062,N_8097);
and U8244 (N_8244,N_8053,N_8003);
and U8245 (N_8245,N_8037,N_8104);
nand U8246 (N_8246,N_8068,N_8041);
or U8247 (N_8247,N_8104,N_8027);
nor U8248 (N_8248,N_8015,N_8044);
xor U8249 (N_8249,N_8022,N_8033);
nand U8250 (N_8250,N_8208,N_8205);
nand U8251 (N_8251,N_8136,N_8202);
nand U8252 (N_8252,N_8160,N_8232);
or U8253 (N_8253,N_8156,N_8129);
nand U8254 (N_8254,N_8192,N_8183);
or U8255 (N_8255,N_8128,N_8155);
nand U8256 (N_8256,N_8228,N_8167);
nor U8257 (N_8257,N_8153,N_8206);
and U8258 (N_8258,N_8143,N_8236);
nor U8259 (N_8259,N_8180,N_8223);
or U8260 (N_8260,N_8164,N_8209);
nand U8261 (N_8261,N_8159,N_8157);
xor U8262 (N_8262,N_8218,N_8234);
or U8263 (N_8263,N_8217,N_8229);
nor U8264 (N_8264,N_8178,N_8174);
nand U8265 (N_8265,N_8235,N_8158);
or U8266 (N_8266,N_8127,N_8233);
or U8267 (N_8267,N_8165,N_8193);
and U8268 (N_8268,N_8220,N_8249);
or U8269 (N_8269,N_8133,N_8248);
and U8270 (N_8270,N_8181,N_8207);
nor U8271 (N_8271,N_8175,N_8179);
nor U8272 (N_8272,N_8242,N_8146);
or U8273 (N_8273,N_8201,N_8142);
and U8274 (N_8274,N_8169,N_8141);
nand U8275 (N_8275,N_8211,N_8162);
or U8276 (N_8276,N_8161,N_8238);
or U8277 (N_8277,N_8198,N_8219);
nor U8278 (N_8278,N_8147,N_8152);
xor U8279 (N_8279,N_8177,N_8195);
and U8280 (N_8280,N_8170,N_8171);
xor U8281 (N_8281,N_8213,N_8196);
nand U8282 (N_8282,N_8163,N_8227);
or U8283 (N_8283,N_8246,N_8215);
and U8284 (N_8284,N_8189,N_8139);
nand U8285 (N_8285,N_8204,N_8140);
nor U8286 (N_8286,N_8125,N_8214);
xor U8287 (N_8287,N_8212,N_8166);
nand U8288 (N_8288,N_8226,N_8200);
nand U8289 (N_8289,N_8225,N_8245);
or U8290 (N_8290,N_8186,N_8190);
nor U8291 (N_8291,N_8210,N_8241);
or U8292 (N_8292,N_8172,N_8188);
and U8293 (N_8293,N_8237,N_8150);
nor U8294 (N_8294,N_8194,N_8176);
nand U8295 (N_8295,N_8231,N_8187);
and U8296 (N_8296,N_8247,N_8224);
and U8297 (N_8297,N_8239,N_8130);
xnor U8298 (N_8298,N_8138,N_8132);
and U8299 (N_8299,N_8199,N_8216);
nor U8300 (N_8300,N_8131,N_8243);
nand U8301 (N_8301,N_8168,N_8173);
nand U8302 (N_8302,N_8135,N_8151);
nand U8303 (N_8303,N_8221,N_8149);
and U8304 (N_8304,N_8230,N_8222);
or U8305 (N_8305,N_8154,N_8184);
xor U8306 (N_8306,N_8148,N_8191);
xor U8307 (N_8307,N_8144,N_8197);
xor U8308 (N_8308,N_8134,N_8240);
nor U8309 (N_8309,N_8244,N_8185);
or U8310 (N_8310,N_8145,N_8126);
or U8311 (N_8311,N_8137,N_8203);
or U8312 (N_8312,N_8182,N_8185);
xor U8313 (N_8313,N_8157,N_8197);
or U8314 (N_8314,N_8133,N_8231);
nor U8315 (N_8315,N_8220,N_8186);
nand U8316 (N_8316,N_8130,N_8218);
and U8317 (N_8317,N_8212,N_8207);
xnor U8318 (N_8318,N_8246,N_8168);
nor U8319 (N_8319,N_8158,N_8219);
nand U8320 (N_8320,N_8196,N_8180);
nor U8321 (N_8321,N_8160,N_8170);
nand U8322 (N_8322,N_8198,N_8140);
xnor U8323 (N_8323,N_8236,N_8146);
nand U8324 (N_8324,N_8153,N_8154);
and U8325 (N_8325,N_8128,N_8132);
nand U8326 (N_8326,N_8226,N_8231);
xnor U8327 (N_8327,N_8139,N_8215);
and U8328 (N_8328,N_8234,N_8158);
and U8329 (N_8329,N_8141,N_8172);
nor U8330 (N_8330,N_8165,N_8216);
and U8331 (N_8331,N_8226,N_8162);
or U8332 (N_8332,N_8232,N_8246);
or U8333 (N_8333,N_8154,N_8236);
nor U8334 (N_8334,N_8191,N_8154);
nand U8335 (N_8335,N_8232,N_8208);
xnor U8336 (N_8336,N_8156,N_8172);
nor U8337 (N_8337,N_8142,N_8157);
xnor U8338 (N_8338,N_8242,N_8194);
nor U8339 (N_8339,N_8227,N_8238);
nand U8340 (N_8340,N_8188,N_8169);
or U8341 (N_8341,N_8157,N_8153);
nor U8342 (N_8342,N_8160,N_8229);
or U8343 (N_8343,N_8151,N_8159);
xor U8344 (N_8344,N_8245,N_8171);
or U8345 (N_8345,N_8194,N_8155);
or U8346 (N_8346,N_8190,N_8206);
nand U8347 (N_8347,N_8221,N_8214);
or U8348 (N_8348,N_8228,N_8151);
xnor U8349 (N_8349,N_8197,N_8132);
or U8350 (N_8350,N_8146,N_8147);
nor U8351 (N_8351,N_8182,N_8163);
and U8352 (N_8352,N_8193,N_8125);
nand U8353 (N_8353,N_8212,N_8240);
and U8354 (N_8354,N_8149,N_8183);
nand U8355 (N_8355,N_8224,N_8207);
and U8356 (N_8356,N_8211,N_8241);
or U8357 (N_8357,N_8176,N_8156);
or U8358 (N_8358,N_8186,N_8242);
nor U8359 (N_8359,N_8185,N_8174);
xor U8360 (N_8360,N_8242,N_8217);
and U8361 (N_8361,N_8147,N_8200);
and U8362 (N_8362,N_8178,N_8230);
and U8363 (N_8363,N_8162,N_8210);
nand U8364 (N_8364,N_8172,N_8178);
and U8365 (N_8365,N_8229,N_8206);
and U8366 (N_8366,N_8162,N_8151);
xnor U8367 (N_8367,N_8208,N_8195);
and U8368 (N_8368,N_8205,N_8195);
or U8369 (N_8369,N_8213,N_8139);
and U8370 (N_8370,N_8146,N_8249);
xor U8371 (N_8371,N_8164,N_8175);
nor U8372 (N_8372,N_8190,N_8233);
and U8373 (N_8373,N_8175,N_8168);
and U8374 (N_8374,N_8191,N_8134);
xor U8375 (N_8375,N_8347,N_8317);
nor U8376 (N_8376,N_8255,N_8333);
xor U8377 (N_8377,N_8284,N_8359);
nand U8378 (N_8378,N_8292,N_8308);
and U8379 (N_8379,N_8288,N_8315);
nor U8380 (N_8380,N_8342,N_8295);
xnor U8381 (N_8381,N_8251,N_8293);
nor U8382 (N_8382,N_8286,N_8257);
or U8383 (N_8383,N_8358,N_8312);
or U8384 (N_8384,N_8351,N_8332);
nor U8385 (N_8385,N_8353,N_8373);
xor U8386 (N_8386,N_8275,N_8321);
and U8387 (N_8387,N_8285,N_8303);
nor U8388 (N_8388,N_8368,N_8304);
xnor U8389 (N_8389,N_8331,N_8302);
or U8390 (N_8390,N_8326,N_8299);
xor U8391 (N_8391,N_8276,N_8372);
xnor U8392 (N_8392,N_8282,N_8340);
xnor U8393 (N_8393,N_8328,N_8357);
and U8394 (N_8394,N_8280,N_8278);
nand U8395 (N_8395,N_8313,N_8283);
nand U8396 (N_8396,N_8269,N_8291);
xnor U8397 (N_8397,N_8352,N_8290);
nor U8398 (N_8398,N_8272,N_8365);
nand U8399 (N_8399,N_8330,N_8256);
xnor U8400 (N_8400,N_8329,N_8287);
nand U8401 (N_8401,N_8298,N_8319);
nand U8402 (N_8402,N_8311,N_8289);
xor U8403 (N_8403,N_8254,N_8363);
nor U8404 (N_8404,N_8345,N_8250);
or U8405 (N_8405,N_8361,N_8274);
xor U8406 (N_8406,N_8266,N_8273);
nor U8407 (N_8407,N_8300,N_8354);
nor U8408 (N_8408,N_8355,N_8264);
or U8409 (N_8409,N_8267,N_8296);
or U8410 (N_8410,N_8271,N_8258);
xnor U8411 (N_8411,N_8366,N_8263);
nand U8412 (N_8412,N_8259,N_8348);
nand U8413 (N_8413,N_8322,N_8318);
nor U8414 (N_8414,N_8360,N_8305);
nand U8415 (N_8415,N_8335,N_8309);
or U8416 (N_8416,N_8344,N_8320);
and U8417 (N_8417,N_8306,N_8371);
xor U8418 (N_8418,N_8277,N_8323);
xnor U8419 (N_8419,N_8297,N_8279);
and U8420 (N_8420,N_8252,N_8339);
or U8421 (N_8421,N_8324,N_8374);
and U8422 (N_8422,N_8336,N_8307);
or U8423 (N_8423,N_8310,N_8265);
nor U8424 (N_8424,N_8367,N_8370);
or U8425 (N_8425,N_8268,N_8314);
xor U8426 (N_8426,N_8301,N_8260);
nor U8427 (N_8427,N_8341,N_8316);
nand U8428 (N_8428,N_8337,N_8253);
or U8429 (N_8429,N_8364,N_8325);
xnor U8430 (N_8430,N_8327,N_8270);
or U8431 (N_8431,N_8349,N_8262);
or U8432 (N_8432,N_8356,N_8294);
nand U8433 (N_8433,N_8350,N_8362);
or U8434 (N_8434,N_8281,N_8346);
nor U8435 (N_8435,N_8338,N_8369);
nand U8436 (N_8436,N_8261,N_8343);
xnor U8437 (N_8437,N_8334,N_8311);
nand U8438 (N_8438,N_8263,N_8347);
and U8439 (N_8439,N_8370,N_8321);
nand U8440 (N_8440,N_8305,N_8274);
or U8441 (N_8441,N_8323,N_8371);
or U8442 (N_8442,N_8368,N_8360);
nand U8443 (N_8443,N_8329,N_8343);
nand U8444 (N_8444,N_8300,N_8320);
nor U8445 (N_8445,N_8315,N_8279);
nor U8446 (N_8446,N_8262,N_8324);
nor U8447 (N_8447,N_8364,N_8261);
or U8448 (N_8448,N_8334,N_8272);
xor U8449 (N_8449,N_8278,N_8292);
and U8450 (N_8450,N_8360,N_8329);
nor U8451 (N_8451,N_8329,N_8345);
and U8452 (N_8452,N_8351,N_8314);
and U8453 (N_8453,N_8293,N_8289);
or U8454 (N_8454,N_8261,N_8258);
xor U8455 (N_8455,N_8280,N_8368);
or U8456 (N_8456,N_8284,N_8310);
nor U8457 (N_8457,N_8274,N_8340);
and U8458 (N_8458,N_8333,N_8287);
nor U8459 (N_8459,N_8272,N_8280);
or U8460 (N_8460,N_8300,N_8255);
xor U8461 (N_8461,N_8259,N_8337);
nand U8462 (N_8462,N_8326,N_8366);
and U8463 (N_8463,N_8271,N_8299);
or U8464 (N_8464,N_8276,N_8307);
xnor U8465 (N_8465,N_8344,N_8346);
or U8466 (N_8466,N_8368,N_8256);
nor U8467 (N_8467,N_8299,N_8256);
nor U8468 (N_8468,N_8263,N_8364);
or U8469 (N_8469,N_8366,N_8340);
and U8470 (N_8470,N_8299,N_8303);
and U8471 (N_8471,N_8267,N_8294);
xnor U8472 (N_8472,N_8281,N_8354);
nor U8473 (N_8473,N_8347,N_8331);
nand U8474 (N_8474,N_8360,N_8346);
xor U8475 (N_8475,N_8312,N_8266);
nor U8476 (N_8476,N_8368,N_8319);
and U8477 (N_8477,N_8352,N_8270);
and U8478 (N_8478,N_8351,N_8347);
nor U8479 (N_8479,N_8364,N_8327);
nor U8480 (N_8480,N_8265,N_8295);
nor U8481 (N_8481,N_8339,N_8334);
nand U8482 (N_8482,N_8342,N_8296);
xor U8483 (N_8483,N_8263,N_8297);
nor U8484 (N_8484,N_8365,N_8367);
or U8485 (N_8485,N_8313,N_8266);
xor U8486 (N_8486,N_8361,N_8352);
nor U8487 (N_8487,N_8364,N_8256);
or U8488 (N_8488,N_8295,N_8299);
and U8489 (N_8489,N_8293,N_8262);
nor U8490 (N_8490,N_8299,N_8360);
or U8491 (N_8491,N_8251,N_8315);
xnor U8492 (N_8492,N_8285,N_8294);
and U8493 (N_8493,N_8325,N_8321);
nand U8494 (N_8494,N_8360,N_8336);
xor U8495 (N_8495,N_8355,N_8359);
xor U8496 (N_8496,N_8283,N_8287);
nand U8497 (N_8497,N_8330,N_8265);
xnor U8498 (N_8498,N_8263,N_8282);
nand U8499 (N_8499,N_8303,N_8290);
nor U8500 (N_8500,N_8389,N_8481);
nand U8501 (N_8501,N_8384,N_8431);
and U8502 (N_8502,N_8432,N_8464);
nor U8503 (N_8503,N_8450,N_8472);
and U8504 (N_8504,N_8385,N_8415);
or U8505 (N_8505,N_8493,N_8383);
or U8506 (N_8506,N_8486,N_8410);
or U8507 (N_8507,N_8488,N_8465);
and U8508 (N_8508,N_8406,N_8490);
nor U8509 (N_8509,N_8427,N_8416);
nand U8510 (N_8510,N_8394,N_8392);
nor U8511 (N_8511,N_8459,N_8435);
nand U8512 (N_8512,N_8401,N_8471);
nand U8513 (N_8513,N_8379,N_8420);
nand U8514 (N_8514,N_8386,N_8381);
xor U8515 (N_8515,N_8495,N_8390);
or U8516 (N_8516,N_8437,N_8395);
or U8517 (N_8517,N_8455,N_8463);
nand U8518 (N_8518,N_8398,N_8447);
and U8519 (N_8519,N_8461,N_8428);
nor U8520 (N_8520,N_8439,N_8440);
and U8521 (N_8521,N_8470,N_8388);
nand U8522 (N_8522,N_8499,N_8396);
nand U8523 (N_8523,N_8422,N_8438);
and U8524 (N_8524,N_8482,N_8491);
or U8525 (N_8525,N_8419,N_8442);
or U8526 (N_8526,N_8407,N_8479);
xnor U8527 (N_8527,N_8475,N_8494);
or U8528 (N_8528,N_8484,N_8468);
nand U8529 (N_8529,N_8391,N_8466);
nor U8530 (N_8530,N_8453,N_8400);
and U8531 (N_8531,N_8476,N_8405);
or U8532 (N_8532,N_8380,N_8397);
and U8533 (N_8533,N_8451,N_8497);
nand U8534 (N_8534,N_8393,N_8378);
nand U8535 (N_8535,N_8460,N_8408);
or U8536 (N_8536,N_8403,N_8489);
xnor U8537 (N_8537,N_8458,N_8480);
and U8538 (N_8538,N_8377,N_8433);
or U8539 (N_8539,N_8376,N_8424);
nand U8540 (N_8540,N_8412,N_8402);
and U8541 (N_8541,N_8448,N_8473);
nor U8542 (N_8542,N_8444,N_8425);
xnor U8543 (N_8543,N_8436,N_8382);
nand U8544 (N_8544,N_8485,N_8387);
or U8545 (N_8545,N_8457,N_8483);
or U8546 (N_8546,N_8409,N_8449);
nand U8547 (N_8547,N_8430,N_8434);
nand U8548 (N_8548,N_8404,N_8467);
nand U8549 (N_8549,N_8456,N_8487);
nand U8550 (N_8550,N_8462,N_8429);
nand U8551 (N_8551,N_8426,N_8446);
nand U8552 (N_8552,N_8417,N_8414);
and U8553 (N_8553,N_8413,N_8399);
nor U8554 (N_8554,N_8477,N_8443);
nor U8555 (N_8555,N_8496,N_8423);
and U8556 (N_8556,N_8498,N_8421);
nor U8557 (N_8557,N_8474,N_8411);
or U8558 (N_8558,N_8492,N_8478);
nand U8559 (N_8559,N_8445,N_8469);
or U8560 (N_8560,N_8418,N_8452);
nor U8561 (N_8561,N_8375,N_8441);
or U8562 (N_8562,N_8454,N_8463);
and U8563 (N_8563,N_8396,N_8454);
nor U8564 (N_8564,N_8446,N_8465);
nor U8565 (N_8565,N_8474,N_8454);
nor U8566 (N_8566,N_8420,N_8482);
xor U8567 (N_8567,N_8464,N_8417);
or U8568 (N_8568,N_8411,N_8454);
nand U8569 (N_8569,N_8449,N_8437);
and U8570 (N_8570,N_8455,N_8490);
nand U8571 (N_8571,N_8407,N_8463);
xnor U8572 (N_8572,N_8414,N_8496);
and U8573 (N_8573,N_8493,N_8417);
xnor U8574 (N_8574,N_8491,N_8448);
xor U8575 (N_8575,N_8433,N_8469);
xor U8576 (N_8576,N_8440,N_8498);
nor U8577 (N_8577,N_8455,N_8472);
nor U8578 (N_8578,N_8418,N_8450);
and U8579 (N_8579,N_8428,N_8485);
xnor U8580 (N_8580,N_8398,N_8383);
nand U8581 (N_8581,N_8464,N_8412);
or U8582 (N_8582,N_8455,N_8406);
xnor U8583 (N_8583,N_8419,N_8409);
nor U8584 (N_8584,N_8452,N_8404);
nand U8585 (N_8585,N_8407,N_8448);
nor U8586 (N_8586,N_8402,N_8478);
nor U8587 (N_8587,N_8465,N_8472);
nand U8588 (N_8588,N_8441,N_8475);
and U8589 (N_8589,N_8455,N_8487);
nor U8590 (N_8590,N_8456,N_8377);
and U8591 (N_8591,N_8484,N_8428);
xnor U8592 (N_8592,N_8485,N_8436);
or U8593 (N_8593,N_8483,N_8443);
or U8594 (N_8594,N_8398,N_8449);
or U8595 (N_8595,N_8411,N_8451);
nor U8596 (N_8596,N_8472,N_8399);
and U8597 (N_8597,N_8403,N_8442);
and U8598 (N_8598,N_8388,N_8456);
xor U8599 (N_8599,N_8469,N_8375);
xnor U8600 (N_8600,N_8456,N_8432);
nor U8601 (N_8601,N_8492,N_8416);
nand U8602 (N_8602,N_8453,N_8385);
nand U8603 (N_8603,N_8424,N_8404);
nor U8604 (N_8604,N_8420,N_8382);
nand U8605 (N_8605,N_8478,N_8399);
nor U8606 (N_8606,N_8395,N_8470);
xnor U8607 (N_8607,N_8396,N_8447);
xnor U8608 (N_8608,N_8396,N_8464);
nor U8609 (N_8609,N_8448,N_8428);
xor U8610 (N_8610,N_8420,N_8397);
and U8611 (N_8611,N_8383,N_8439);
or U8612 (N_8612,N_8437,N_8452);
and U8613 (N_8613,N_8476,N_8470);
nand U8614 (N_8614,N_8431,N_8427);
xnor U8615 (N_8615,N_8417,N_8457);
and U8616 (N_8616,N_8453,N_8454);
nand U8617 (N_8617,N_8468,N_8404);
nand U8618 (N_8618,N_8412,N_8377);
xor U8619 (N_8619,N_8390,N_8383);
or U8620 (N_8620,N_8409,N_8434);
nor U8621 (N_8621,N_8444,N_8441);
xor U8622 (N_8622,N_8484,N_8447);
and U8623 (N_8623,N_8393,N_8409);
xor U8624 (N_8624,N_8381,N_8447);
and U8625 (N_8625,N_8531,N_8505);
nor U8626 (N_8626,N_8502,N_8500);
nor U8627 (N_8627,N_8567,N_8508);
xnor U8628 (N_8628,N_8592,N_8525);
and U8629 (N_8629,N_8591,N_8614);
and U8630 (N_8630,N_8545,N_8609);
or U8631 (N_8631,N_8564,N_8586);
nand U8632 (N_8632,N_8528,N_8590);
xnor U8633 (N_8633,N_8541,N_8555);
nand U8634 (N_8634,N_8540,N_8549);
xor U8635 (N_8635,N_8529,N_8518);
nand U8636 (N_8636,N_8559,N_8560);
and U8637 (N_8637,N_8580,N_8503);
nand U8638 (N_8638,N_8527,N_8579);
nor U8639 (N_8639,N_8601,N_8556);
and U8640 (N_8640,N_8513,N_8512);
and U8641 (N_8641,N_8557,N_8603);
nand U8642 (N_8642,N_8514,N_8618);
nand U8643 (N_8643,N_8551,N_8552);
nand U8644 (N_8644,N_8621,N_8602);
xor U8645 (N_8645,N_8605,N_8569);
and U8646 (N_8646,N_8516,N_8538);
xor U8647 (N_8647,N_8574,N_8517);
xnor U8648 (N_8648,N_8611,N_8617);
and U8649 (N_8649,N_8534,N_8604);
xnor U8650 (N_8650,N_8571,N_8526);
or U8651 (N_8651,N_8565,N_8568);
and U8652 (N_8652,N_8544,N_8577);
and U8653 (N_8653,N_8535,N_8519);
xnor U8654 (N_8654,N_8520,N_8588);
nor U8655 (N_8655,N_8561,N_8523);
xnor U8656 (N_8656,N_8533,N_8606);
or U8657 (N_8657,N_8610,N_8548);
or U8658 (N_8658,N_8537,N_8532);
or U8659 (N_8659,N_8598,N_8554);
xor U8660 (N_8660,N_8585,N_8619);
and U8661 (N_8661,N_8511,N_8543);
and U8662 (N_8662,N_8524,N_8595);
or U8663 (N_8663,N_8607,N_8563);
or U8664 (N_8664,N_8573,N_8558);
nand U8665 (N_8665,N_8624,N_8608);
and U8666 (N_8666,N_8570,N_8509);
or U8667 (N_8667,N_8597,N_8510);
and U8668 (N_8668,N_8521,N_8596);
and U8669 (N_8669,N_8504,N_8550);
xor U8670 (N_8670,N_8622,N_8581);
or U8671 (N_8671,N_8522,N_8566);
nor U8672 (N_8672,N_8612,N_8547);
nor U8673 (N_8673,N_8553,N_8536);
or U8674 (N_8674,N_8507,N_8515);
and U8675 (N_8675,N_8539,N_8599);
nand U8676 (N_8676,N_8616,N_8600);
or U8677 (N_8677,N_8615,N_8584);
and U8678 (N_8678,N_8576,N_8542);
nor U8679 (N_8679,N_8623,N_8613);
or U8680 (N_8680,N_8575,N_8583);
nand U8681 (N_8681,N_8578,N_8582);
xor U8682 (N_8682,N_8593,N_8589);
and U8683 (N_8683,N_8506,N_8501);
and U8684 (N_8684,N_8587,N_8572);
and U8685 (N_8685,N_8620,N_8546);
xnor U8686 (N_8686,N_8594,N_8530);
and U8687 (N_8687,N_8562,N_8503);
or U8688 (N_8688,N_8581,N_8600);
nand U8689 (N_8689,N_8586,N_8524);
xor U8690 (N_8690,N_8616,N_8554);
nand U8691 (N_8691,N_8593,N_8545);
xor U8692 (N_8692,N_8565,N_8518);
nor U8693 (N_8693,N_8503,N_8526);
xor U8694 (N_8694,N_8587,N_8575);
xor U8695 (N_8695,N_8603,N_8612);
or U8696 (N_8696,N_8602,N_8520);
xor U8697 (N_8697,N_8611,N_8534);
nand U8698 (N_8698,N_8504,N_8573);
or U8699 (N_8699,N_8525,N_8596);
xnor U8700 (N_8700,N_8607,N_8525);
or U8701 (N_8701,N_8515,N_8578);
nand U8702 (N_8702,N_8540,N_8591);
xnor U8703 (N_8703,N_8569,N_8506);
xnor U8704 (N_8704,N_8617,N_8570);
nor U8705 (N_8705,N_8507,N_8523);
xor U8706 (N_8706,N_8603,N_8528);
nand U8707 (N_8707,N_8620,N_8618);
nor U8708 (N_8708,N_8530,N_8506);
or U8709 (N_8709,N_8548,N_8517);
nor U8710 (N_8710,N_8536,N_8504);
and U8711 (N_8711,N_8506,N_8604);
xnor U8712 (N_8712,N_8623,N_8606);
xor U8713 (N_8713,N_8613,N_8508);
and U8714 (N_8714,N_8519,N_8595);
or U8715 (N_8715,N_8585,N_8571);
nor U8716 (N_8716,N_8576,N_8621);
and U8717 (N_8717,N_8571,N_8539);
nor U8718 (N_8718,N_8507,N_8578);
xnor U8719 (N_8719,N_8558,N_8577);
or U8720 (N_8720,N_8542,N_8613);
nor U8721 (N_8721,N_8561,N_8601);
and U8722 (N_8722,N_8544,N_8550);
and U8723 (N_8723,N_8572,N_8576);
nand U8724 (N_8724,N_8550,N_8562);
or U8725 (N_8725,N_8611,N_8580);
nand U8726 (N_8726,N_8542,N_8567);
nor U8727 (N_8727,N_8505,N_8620);
and U8728 (N_8728,N_8612,N_8551);
nor U8729 (N_8729,N_8562,N_8596);
or U8730 (N_8730,N_8601,N_8510);
and U8731 (N_8731,N_8618,N_8587);
xnor U8732 (N_8732,N_8620,N_8523);
nor U8733 (N_8733,N_8551,N_8522);
nor U8734 (N_8734,N_8584,N_8564);
nor U8735 (N_8735,N_8579,N_8576);
xor U8736 (N_8736,N_8617,N_8562);
and U8737 (N_8737,N_8578,N_8592);
and U8738 (N_8738,N_8557,N_8520);
or U8739 (N_8739,N_8615,N_8548);
and U8740 (N_8740,N_8616,N_8559);
or U8741 (N_8741,N_8503,N_8579);
xor U8742 (N_8742,N_8500,N_8542);
nand U8743 (N_8743,N_8523,N_8519);
nor U8744 (N_8744,N_8541,N_8619);
and U8745 (N_8745,N_8622,N_8598);
nor U8746 (N_8746,N_8600,N_8539);
nor U8747 (N_8747,N_8507,N_8541);
or U8748 (N_8748,N_8556,N_8534);
xor U8749 (N_8749,N_8576,N_8624);
and U8750 (N_8750,N_8717,N_8736);
xor U8751 (N_8751,N_8699,N_8692);
nor U8752 (N_8752,N_8653,N_8731);
xnor U8753 (N_8753,N_8660,N_8687);
nor U8754 (N_8754,N_8688,N_8684);
and U8755 (N_8755,N_8715,N_8719);
nor U8756 (N_8756,N_8672,N_8658);
or U8757 (N_8757,N_8635,N_8727);
and U8758 (N_8758,N_8649,N_8666);
xnor U8759 (N_8759,N_8633,N_8686);
nor U8760 (N_8760,N_8728,N_8740);
or U8761 (N_8761,N_8721,N_8663);
nand U8762 (N_8762,N_8657,N_8701);
nand U8763 (N_8763,N_8675,N_8691);
and U8764 (N_8764,N_8748,N_8638);
xor U8765 (N_8765,N_8646,N_8669);
xnor U8766 (N_8766,N_8704,N_8706);
or U8767 (N_8767,N_8739,N_8634);
nor U8768 (N_8768,N_8738,N_8735);
xor U8769 (N_8769,N_8673,N_8671);
and U8770 (N_8770,N_8723,N_8641);
nand U8771 (N_8771,N_8667,N_8733);
nor U8772 (N_8772,N_8674,N_8726);
or U8773 (N_8773,N_8690,N_8722);
xor U8774 (N_8774,N_8689,N_8696);
and U8775 (N_8775,N_8642,N_8631);
or U8776 (N_8776,N_8645,N_8713);
and U8777 (N_8777,N_8716,N_8743);
nand U8778 (N_8778,N_8680,N_8654);
and U8779 (N_8779,N_8681,N_8676);
and U8780 (N_8780,N_8714,N_8747);
or U8781 (N_8781,N_8685,N_8712);
xor U8782 (N_8782,N_8682,N_8678);
nor U8783 (N_8783,N_8625,N_8630);
nor U8784 (N_8784,N_8711,N_8640);
nor U8785 (N_8785,N_8742,N_8724);
xnor U8786 (N_8786,N_8632,N_8734);
nor U8787 (N_8787,N_8697,N_8695);
and U8788 (N_8788,N_8679,N_8677);
nor U8789 (N_8789,N_8656,N_8650);
nor U8790 (N_8790,N_8629,N_8749);
or U8791 (N_8791,N_8705,N_8737);
nor U8792 (N_8792,N_8700,N_8718);
and U8793 (N_8793,N_8683,N_8647);
nand U8794 (N_8794,N_8698,N_8746);
xor U8795 (N_8795,N_8707,N_8626);
nor U8796 (N_8796,N_8648,N_8741);
and U8797 (N_8797,N_8708,N_8745);
and U8798 (N_8798,N_8643,N_8668);
nor U8799 (N_8799,N_8644,N_8659);
and U8800 (N_8800,N_8725,N_8732);
nand U8801 (N_8801,N_8710,N_8652);
or U8802 (N_8802,N_8628,N_8661);
xor U8803 (N_8803,N_8651,N_8636);
xnor U8804 (N_8804,N_8639,N_8693);
xnor U8805 (N_8805,N_8665,N_8670);
or U8806 (N_8806,N_8655,N_8709);
xor U8807 (N_8807,N_8730,N_8702);
or U8808 (N_8808,N_8694,N_8703);
and U8809 (N_8809,N_8729,N_8637);
or U8810 (N_8810,N_8664,N_8662);
or U8811 (N_8811,N_8627,N_8744);
nand U8812 (N_8812,N_8720,N_8694);
nor U8813 (N_8813,N_8697,N_8694);
nor U8814 (N_8814,N_8644,N_8648);
nand U8815 (N_8815,N_8627,N_8679);
nor U8816 (N_8816,N_8630,N_8648);
nand U8817 (N_8817,N_8667,N_8675);
or U8818 (N_8818,N_8630,N_8669);
nand U8819 (N_8819,N_8677,N_8632);
xor U8820 (N_8820,N_8713,N_8736);
xor U8821 (N_8821,N_8657,N_8684);
or U8822 (N_8822,N_8635,N_8665);
or U8823 (N_8823,N_8732,N_8641);
nor U8824 (N_8824,N_8730,N_8712);
xnor U8825 (N_8825,N_8639,N_8728);
and U8826 (N_8826,N_8707,N_8710);
and U8827 (N_8827,N_8651,N_8701);
or U8828 (N_8828,N_8738,N_8727);
nor U8829 (N_8829,N_8748,N_8664);
xnor U8830 (N_8830,N_8646,N_8683);
nand U8831 (N_8831,N_8631,N_8744);
xor U8832 (N_8832,N_8672,N_8696);
xor U8833 (N_8833,N_8703,N_8717);
xnor U8834 (N_8834,N_8653,N_8746);
xnor U8835 (N_8835,N_8716,N_8748);
nand U8836 (N_8836,N_8666,N_8690);
nor U8837 (N_8837,N_8721,N_8633);
xor U8838 (N_8838,N_8746,N_8740);
nor U8839 (N_8839,N_8669,N_8717);
nand U8840 (N_8840,N_8625,N_8747);
xnor U8841 (N_8841,N_8746,N_8733);
xnor U8842 (N_8842,N_8652,N_8701);
and U8843 (N_8843,N_8746,N_8691);
xor U8844 (N_8844,N_8699,N_8724);
and U8845 (N_8845,N_8694,N_8690);
nor U8846 (N_8846,N_8689,N_8749);
or U8847 (N_8847,N_8722,N_8636);
xnor U8848 (N_8848,N_8711,N_8709);
xor U8849 (N_8849,N_8666,N_8709);
and U8850 (N_8850,N_8711,N_8744);
nor U8851 (N_8851,N_8717,N_8655);
and U8852 (N_8852,N_8638,N_8744);
nor U8853 (N_8853,N_8676,N_8639);
or U8854 (N_8854,N_8637,N_8640);
and U8855 (N_8855,N_8711,N_8645);
nor U8856 (N_8856,N_8700,N_8735);
or U8857 (N_8857,N_8626,N_8639);
nor U8858 (N_8858,N_8685,N_8732);
or U8859 (N_8859,N_8721,N_8627);
nor U8860 (N_8860,N_8643,N_8697);
or U8861 (N_8861,N_8691,N_8672);
nand U8862 (N_8862,N_8656,N_8726);
xnor U8863 (N_8863,N_8629,N_8736);
xnor U8864 (N_8864,N_8691,N_8650);
nor U8865 (N_8865,N_8743,N_8701);
or U8866 (N_8866,N_8700,N_8742);
and U8867 (N_8867,N_8638,N_8715);
and U8868 (N_8868,N_8699,N_8638);
nor U8869 (N_8869,N_8630,N_8711);
xnor U8870 (N_8870,N_8636,N_8698);
and U8871 (N_8871,N_8637,N_8722);
xor U8872 (N_8872,N_8689,N_8646);
xnor U8873 (N_8873,N_8679,N_8660);
or U8874 (N_8874,N_8634,N_8650);
and U8875 (N_8875,N_8847,N_8773);
xor U8876 (N_8876,N_8801,N_8792);
or U8877 (N_8877,N_8826,N_8760);
nand U8878 (N_8878,N_8779,N_8818);
and U8879 (N_8879,N_8859,N_8821);
and U8880 (N_8880,N_8820,N_8813);
or U8881 (N_8881,N_8823,N_8803);
or U8882 (N_8882,N_8804,N_8854);
nand U8883 (N_8883,N_8758,N_8829);
xor U8884 (N_8884,N_8782,N_8832);
or U8885 (N_8885,N_8831,N_8750);
nor U8886 (N_8886,N_8849,N_8767);
nand U8887 (N_8887,N_8762,N_8855);
nor U8888 (N_8888,N_8771,N_8787);
and U8889 (N_8889,N_8822,N_8825);
or U8890 (N_8890,N_8751,N_8786);
xnor U8891 (N_8891,N_8754,N_8815);
or U8892 (N_8892,N_8863,N_8796);
xor U8893 (N_8893,N_8862,N_8761);
nand U8894 (N_8894,N_8840,N_8851);
and U8895 (N_8895,N_8830,N_8770);
nor U8896 (N_8896,N_8763,N_8841);
and U8897 (N_8897,N_8802,N_8811);
nor U8898 (N_8898,N_8853,N_8867);
nand U8899 (N_8899,N_8809,N_8864);
or U8900 (N_8900,N_8785,N_8874);
or U8901 (N_8901,N_8807,N_8780);
nand U8902 (N_8902,N_8752,N_8790);
xnor U8903 (N_8903,N_8837,N_8795);
nand U8904 (N_8904,N_8778,N_8846);
nand U8905 (N_8905,N_8810,N_8806);
xor U8906 (N_8906,N_8860,N_8756);
xor U8907 (N_8907,N_8852,N_8857);
nor U8908 (N_8908,N_8794,N_8793);
and U8909 (N_8909,N_8868,N_8819);
nand U8910 (N_8910,N_8799,N_8757);
xnor U8911 (N_8911,N_8856,N_8845);
xnor U8912 (N_8912,N_8842,N_8850);
nor U8913 (N_8913,N_8844,N_8866);
and U8914 (N_8914,N_8768,N_8776);
xnor U8915 (N_8915,N_8766,N_8765);
xnor U8916 (N_8916,N_8753,N_8775);
nor U8917 (N_8917,N_8817,N_8788);
nor U8918 (N_8918,N_8861,N_8784);
nor U8919 (N_8919,N_8789,N_8828);
nand U8920 (N_8920,N_8759,N_8777);
and U8921 (N_8921,N_8836,N_8865);
xnor U8922 (N_8922,N_8800,N_8772);
nor U8923 (N_8923,N_8869,N_8827);
or U8924 (N_8924,N_8764,N_8838);
nor U8925 (N_8925,N_8798,N_8835);
and U8926 (N_8926,N_8833,N_8769);
and U8927 (N_8927,N_8848,N_8814);
nand U8928 (N_8928,N_8870,N_8781);
and U8929 (N_8929,N_8839,N_8774);
nor U8930 (N_8930,N_8812,N_8755);
and U8931 (N_8931,N_8791,N_8805);
nand U8932 (N_8932,N_8816,N_8808);
nor U8933 (N_8933,N_8783,N_8858);
nand U8934 (N_8934,N_8834,N_8871);
and U8935 (N_8935,N_8843,N_8873);
nand U8936 (N_8936,N_8824,N_8872);
nor U8937 (N_8937,N_8797,N_8839);
nand U8938 (N_8938,N_8838,N_8807);
and U8939 (N_8939,N_8827,N_8873);
nor U8940 (N_8940,N_8851,N_8784);
nor U8941 (N_8941,N_8835,N_8829);
xnor U8942 (N_8942,N_8795,N_8871);
nor U8943 (N_8943,N_8844,N_8839);
nor U8944 (N_8944,N_8815,N_8858);
or U8945 (N_8945,N_8854,N_8768);
xnor U8946 (N_8946,N_8804,N_8789);
nand U8947 (N_8947,N_8808,N_8788);
or U8948 (N_8948,N_8820,N_8771);
xnor U8949 (N_8949,N_8799,N_8856);
or U8950 (N_8950,N_8768,N_8763);
nand U8951 (N_8951,N_8826,N_8824);
nor U8952 (N_8952,N_8849,N_8780);
nor U8953 (N_8953,N_8820,N_8750);
and U8954 (N_8954,N_8865,N_8768);
nand U8955 (N_8955,N_8815,N_8753);
nand U8956 (N_8956,N_8841,N_8812);
nand U8957 (N_8957,N_8839,N_8820);
xnor U8958 (N_8958,N_8864,N_8779);
and U8959 (N_8959,N_8800,N_8783);
nor U8960 (N_8960,N_8794,N_8838);
xor U8961 (N_8961,N_8806,N_8838);
nor U8962 (N_8962,N_8843,N_8810);
and U8963 (N_8963,N_8827,N_8842);
or U8964 (N_8964,N_8768,N_8873);
xor U8965 (N_8965,N_8768,N_8833);
or U8966 (N_8966,N_8814,N_8821);
nor U8967 (N_8967,N_8822,N_8832);
or U8968 (N_8968,N_8764,N_8793);
nand U8969 (N_8969,N_8794,N_8870);
and U8970 (N_8970,N_8795,N_8857);
nor U8971 (N_8971,N_8782,N_8780);
and U8972 (N_8972,N_8833,N_8818);
and U8973 (N_8973,N_8822,N_8827);
xor U8974 (N_8974,N_8871,N_8850);
and U8975 (N_8975,N_8751,N_8777);
nand U8976 (N_8976,N_8776,N_8864);
nand U8977 (N_8977,N_8838,N_8789);
and U8978 (N_8978,N_8843,N_8766);
or U8979 (N_8979,N_8829,N_8839);
nand U8980 (N_8980,N_8773,N_8767);
and U8981 (N_8981,N_8831,N_8754);
nand U8982 (N_8982,N_8842,N_8755);
nand U8983 (N_8983,N_8773,N_8835);
nand U8984 (N_8984,N_8778,N_8764);
or U8985 (N_8985,N_8855,N_8836);
or U8986 (N_8986,N_8819,N_8797);
nor U8987 (N_8987,N_8856,N_8789);
xor U8988 (N_8988,N_8786,N_8874);
or U8989 (N_8989,N_8871,N_8793);
nand U8990 (N_8990,N_8813,N_8858);
nor U8991 (N_8991,N_8822,N_8826);
nor U8992 (N_8992,N_8792,N_8869);
nor U8993 (N_8993,N_8819,N_8822);
nand U8994 (N_8994,N_8847,N_8775);
nor U8995 (N_8995,N_8838,N_8791);
nand U8996 (N_8996,N_8804,N_8756);
nand U8997 (N_8997,N_8787,N_8807);
or U8998 (N_8998,N_8860,N_8813);
xor U8999 (N_8999,N_8751,N_8753);
xor U9000 (N_9000,N_8894,N_8994);
and U9001 (N_9001,N_8920,N_8931);
nor U9002 (N_9002,N_8905,N_8917);
nand U9003 (N_9003,N_8963,N_8875);
or U9004 (N_9004,N_8982,N_8906);
nand U9005 (N_9005,N_8925,N_8964);
nand U9006 (N_9006,N_8888,N_8961);
xnor U9007 (N_9007,N_8885,N_8900);
nand U9008 (N_9008,N_8895,N_8914);
xor U9009 (N_9009,N_8876,N_8977);
xor U9010 (N_9010,N_8921,N_8949);
and U9011 (N_9011,N_8992,N_8986);
and U9012 (N_9012,N_8922,N_8946);
or U9013 (N_9013,N_8918,N_8954);
xnor U9014 (N_9014,N_8934,N_8939);
and U9015 (N_9015,N_8912,N_8987);
or U9016 (N_9016,N_8877,N_8995);
nand U9017 (N_9017,N_8990,N_8965);
xnor U9018 (N_9018,N_8923,N_8969);
nand U9019 (N_9019,N_8952,N_8883);
nand U9020 (N_9020,N_8878,N_8936);
and U9021 (N_9021,N_8893,N_8950);
xnor U9022 (N_9022,N_8926,N_8983);
and U9023 (N_9023,N_8901,N_8968);
or U9024 (N_9024,N_8972,N_8966);
or U9025 (N_9025,N_8919,N_8997);
nand U9026 (N_9026,N_8907,N_8970);
or U9027 (N_9027,N_8882,N_8890);
and U9028 (N_9028,N_8929,N_8889);
xor U9029 (N_9029,N_8957,N_8951);
nand U9030 (N_9030,N_8979,N_8967);
and U9031 (N_9031,N_8910,N_8935);
or U9032 (N_9032,N_8909,N_8980);
and U9033 (N_9033,N_8903,N_8948);
xnor U9034 (N_9034,N_8928,N_8973);
or U9035 (N_9035,N_8911,N_8940);
or U9036 (N_9036,N_8924,N_8993);
nand U9037 (N_9037,N_8974,N_8879);
or U9038 (N_9038,N_8908,N_8981);
and U9039 (N_9039,N_8988,N_8959);
nor U9040 (N_9040,N_8886,N_8880);
and U9041 (N_9041,N_8943,N_8976);
nor U9042 (N_9042,N_8941,N_8932);
or U9043 (N_9043,N_8953,N_8930);
and U9044 (N_9044,N_8984,N_8915);
and U9045 (N_9045,N_8971,N_8942);
or U9046 (N_9046,N_8887,N_8891);
nand U9047 (N_9047,N_8945,N_8996);
nor U9048 (N_9048,N_8999,N_8978);
nor U9049 (N_9049,N_8937,N_8938);
or U9050 (N_9050,N_8884,N_8956);
nor U9051 (N_9051,N_8904,N_8896);
and U9052 (N_9052,N_8962,N_8960);
nand U9053 (N_9053,N_8989,N_8998);
xor U9054 (N_9054,N_8881,N_8944);
nand U9055 (N_9055,N_8897,N_8916);
xnor U9056 (N_9056,N_8947,N_8955);
and U9057 (N_9057,N_8898,N_8958);
nor U9058 (N_9058,N_8985,N_8899);
xor U9059 (N_9059,N_8975,N_8991);
xor U9060 (N_9060,N_8913,N_8927);
and U9061 (N_9061,N_8892,N_8933);
or U9062 (N_9062,N_8902,N_8909);
xor U9063 (N_9063,N_8898,N_8949);
nand U9064 (N_9064,N_8974,N_8969);
nor U9065 (N_9065,N_8952,N_8949);
xor U9066 (N_9066,N_8932,N_8965);
xnor U9067 (N_9067,N_8994,N_8954);
or U9068 (N_9068,N_8953,N_8994);
or U9069 (N_9069,N_8992,N_8958);
and U9070 (N_9070,N_8923,N_8994);
nand U9071 (N_9071,N_8894,N_8946);
nand U9072 (N_9072,N_8878,N_8973);
nand U9073 (N_9073,N_8896,N_8917);
nor U9074 (N_9074,N_8922,N_8947);
or U9075 (N_9075,N_8926,N_8945);
nand U9076 (N_9076,N_8906,N_8938);
or U9077 (N_9077,N_8933,N_8957);
or U9078 (N_9078,N_8893,N_8961);
nor U9079 (N_9079,N_8955,N_8886);
or U9080 (N_9080,N_8939,N_8904);
or U9081 (N_9081,N_8978,N_8900);
xnor U9082 (N_9082,N_8936,N_8998);
nand U9083 (N_9083,N_8918,N_8983);
and U9084 (N_9084,N_8903,N_8966);
nand U9085 (N_9085,N_8970,N_8985);
nor U9086 (N_9086,N_8940,N_8993);
nand U9087 (N_9087,N_8887,N_8925);
nor U9088 (N_9088,N_8978,N_8895);
nor U9089 (N_9089,N_8918,N_8923);
nand U9090 (N_9090,N_8897,N_8929);
nand U9091 (N_9091,N_8986,N_8906);
nand U9092 (N_9092,N_8948,N_8880);
nand U9093 (N_9093,N_8968,N_8949);
nand U9094 (N_9094,N_8957,N_8947);
nor U9095 (N_9095,N_8967,N_8906);
and U9096 (N_9096,N_8886,N_8891);
nor U9097 (N_9097,N_8907,N_8949);
nor U9098 (N_9098,N_8885,N_8879);
nor U9099 (N_9099,N_8881,N_8992);
xor U9100 (N_9100,N_8998,N_8963);
nor U9101 (N_9101,N_8958,N_8882);
nor U9102 (N_9102,N_8993,N_8969);
nand U9103 (N_9103,N_8932,N_8907);
or U9104 (N_9104,N_8920,N_8921);
nand U9105 (N_9105,N_8915,N_8898);
nand U9106 (N_9106,N_8928,N_8888);
nor U9107 (N_9107,N_8988,N_8965);
or U9108 (N_9108,N_8877,N_8907);
xnor U9109 (N_9109,N_8922,N_8897);
xor U9110 (N_9110,N_8950,N_8905);
or U9111 (N_9111,N_8960,N_8946);
and U9112 (N_9112,N_8892,N_8945);
nor U9113 (N_9113,N_8996,N_8955);
and U9114 (N_9114,N_8994,N_8903);
xnor U9115 (N_9115,N_8963,N_8895);
or U9116 (N_9116,N_8904,N_8903);
nor U9117 (N_9117,N_8902,N_8894);
nand U9118 (N_9118,N_8967,N_8897);
nor U9119 (N_9119,N_8953,N_8911);
nand U9120 (N_9120,N_8954,N_8944);
nand U9121 (N_9121,N_8954,N_8890);
and U9122 (N_9122,N_8961,N_8875);
xnor U9123 (N_9123,N_8886,N_8956);
and U9124 (N_9124,N_8988,N_8912);
nor U9125 (N_9125,N_9088,N_9005);
or U9126 (N_9126,N_9118,N_9122);
or U9127 (N_9127,N_9067,N_9042);
nand U9128 (N_9128,N_9079,N_9048);
xor U9129 (N_9129,N_9041,N_9040);
or U9130 (N_9130,N_9068,N_9020);
xor U9131 (N_9131,N_9097,N_9013);
xnor U9132 (N_9132,N_9000,N_9085);
or U9133 (N_9133,N_9065,N_9110);
and U9134 (N_9134,N_9109,N_9124);
nor U9135 (N_9135,N_9116,N_9015);
nand U9136 (N_9136,N_9036,N_9078);
xor U9137 (N_9137,N_9034,N_9007);
nand U9138 (N_9138,N_9012,N_9086);
nor U9139 (N_9139,N_9084,N_9063);
xnor U9140 (N_9140,N_9003,N_9031);
xnor U9141 (N_9141,N_9108,N_9098);
xnor U9142 (N_9142,N_9073,N_9083);
and U9143 (N_9143,N_9001,N_9014);
or U9144 (N_9144,N_9062,N_9071);
nand U9145 (N_9145,N_9103,N_9018);
or U9146 (N_9146,N_9044,N_9053);
nand U9147 (N_9147,N_9093,N_9120);
nor U9148 (N_9148,N_9050,N_9107);
xor U9149 (N_9149,N_9035,N_9056);
xnor U9150 (N_9150,N_9002,N_9119);
nor U9151 (N_9151,N_9057,N_9029);
and U9152 (N_9152,N_9046,N_9096);
nor U9153 (N_9153,N_9037,N_9010);
and U9154 (N_9154,N_9087,N_9076);
nand U9155 (N_9155,N_9023,N_9106);
nand U9156 (N_9156,N_9069,N_9028);
or U9157 (N_9157,N_9082,N_9099);
nand U9158 (N_9158,N_9021,N_9101);
nand U9159 (N_9159,N_9077,N_9055);
xnor U9160 (N_9160,N_9016,N_9009);
and U9161 (N_9161,N_9052,N_9033);
xor U9162 (N_9162,N_9072,N_9112);
xnor U9163 (N_9163,N_9080,N_9094);
nand U9164 (N_9164,N_9022,N_9051);
and U9165 (N_9165,N_9039,N_9017);
nor U9166 (N_9166,N_9117,N_9090);
or U9167 (N_9167,N_9089,N_9030);
xnor U9168 (N_9168,N_9043,N_9004);
xnor U9169 (N_9169,N_9074,N_9049);
nor U9170 (N_9170,N_9111,N_9027);
or U9171 (N_9171,N_9121,N_9105);
nor U9172 (N_9172,N_9081,N_9113);
nor U9173 (N_9173,N_9019,N_9092);
and U9174 (N_9174,N_9006,N_9114);
nor U9175 (N_9175,N_9058,N_9070);
xor U9176 (N_9176,N_9045,N_9032);
nor U9177 (N_9177,N_9038,N_9100);
xor U9178 (N_9178,N_9061,N_9054);
or U9179 (N_9179,N_9008,N_9104);
and U9180 (N_9180,N_9047,N_9060);
and U9181 (N_9181,N_9026,N_9064);
nand U9182 (N_9182,N_9095,N_9025);
and U9183 (N_9183,N_9075,N_9123);
nor U9184 (N_9184,N_9024,N_9066);
nand U9185 (N_9185,N_9011,N_9091);
or U9186 (N_9186,N_9115,N_9059);
xnor U9187 (N_9187,N_9102,N_9013);
or U9188 (N_9188,N_9116,N_9098);
or U9189 (N_9189,N_9024,N_9027);
or U9190 (N_9190,N_9003,N_9085);
nor U9191 (N_9191,N_9112,N_9102);
and U9192 (N_9192,N_9056,N_9111);
xor U9193 (N_9193,N_9031,N_9032);
nand U9194 (N_9194,N_9066,N_9003);
nand U9195 (N_9195,N_9104,N_9001);
xor U9196 (N_9196,N_9036,N_9064);
or U9197 (N_9197,N_9058,N_9019);
nand U9198 (N_9198,N_9060,N_9085);
and U9199 (N_9199,N_9074,N_9080);
xor U9200 (N_9200,N_9088,N_9006);
nand U9201 (N_9201,N_9078,N_9122);
and U9202 (N_9202,N_9079,N_9124);
or U9203 (N_9203,N_9106,N_9042);
or U9204 (N_9204,N_9056,N_9052);
or U9205 (N_9205,N_9053,N_9113);
nand U9206 (N_9206,N_9084,N_9082);
xnor U9207 (N_9207,N_9053,N_9105);
and U9208 (N_9208,N_9085,N_9062);
xor U9209 (N_9209,N_9010,N_9114);
xnor U9210 (N_9210,N_9060,N_9044);
and U9211 (N_9211,N_9014,N_9037);
or U9212 (N_9212,N_9101,N_9117);
or U9213 (N_9213,N_9102,N_9032);
and U9214 (N_9214,N_9118,N_9073);
and U9215 (N_9215,N_9124,N_9104);
xor U9216 (N_9216,N_9041,N_9102);
and U9217 (N_9217,N_9092,N_9088);
nor U9218 (N_9218,N_9024,N_9090);
xnor U9219 (N_9219,N_9031,N_9044);
or U9220 (N_9220,N_9080,N_9076);
xor U9221 (N_9221,N_9003,N_9093);
nand U9222 (N_9222,N_9100,N_9005);
nor U9223 (N_9223,N_9010,N_9017);
xor U9224 (N_9224,N_9009,N_9038);
nor U9225 (N_9225,N_9005,N_9071);
or U9226 (N_9226,N_9025,N_9102);
or U9227 (N_9227,N_9066,N_9068);
nor U9228 (N_9228,N_9117,N_9069);
and U9229 (N_9229,N_9048,N_9021);
nor U9230 (N_9230,N_9035,N_9097);
xor U9231 (N_9231,N_9065,N_9090);
nor U9232 (N_9232,N_9027,N_9045);
and U9233 (N_9233,N_9085,N_9046);
nand U9234 (N_9234,N_9121,N_9050);
nor U9235 (N_9235,N_9062,N_9024);
nor U9236 (N_9236,N_9033,N_9070);
or U9237 (N_9237,N_9090,N_9084);
nor U9238 (N_9238,N_9035,N_9123);
nand U9239 (N_9239,N_9056,N_9037);
and U9240 (N_9240,N_9067,N_9066);
and U9241 (N_9241,N_9000,N_9119);
nand U9242 (N_9242,N_9063,N_9021);
nand U9243 (N_9243,N_9031,N_9091);
xor U9244 (N_9244,N_9123,N_9006);
xor U9245 (N_9245,N_9016,N_9105);
xnor U9246 (N_9246,N_9055,N_9078);
xor U9247 (N_9247,N_9107,N_9017);
or U9248 (N_9248,N_9021,N_9016);
nand U9249 (N_9249,N_9107,N_9086);
nor U9250 (N_9250,N_9246,N_9236);
nand U9251 (N_9251,N_9132,N_9160);
or U9252 (N_9252,N_9149,N_9181);
xor U9253 (N_9253,N_9226,N_9135);
nor U9254 (N_9254,N_9139,N_9245);
nor U9255 (N_9255,N_9205,N_9158);
xnor U9256 (N_9256,N_9168,N_9189);
xnor U9257 (N_9257,N_9224,N_9147);
and U9258 (N_9258,N_9161,N_9238);
xnor U9259 (N_9259,N_9131,N_9156);
and U9260 (N_9260,N_9174,N_9231);
and U9261 (N_9261,N_9130,N_9159);
xnor U9262 (N_9262,N_9235,N_9134);
or U9263 (N_9263,N_9170,N_9210);
xnor U9264 (N_9264,N_9162,N_9143);
nor U9265 (N_9265,N_9186,N_9171);
or U9266 (N_9266,N_9185,N_9216);
and U9267 (N_9267,N_9145,N_9165);
and U9268 (N_9268,N_9196,N_9163);
xor U9269 (N_9269,N_9191,N_9142);
and U9270 (N_9270,N_9232,N_9207);
nor U9271 (N_9271,N_9199,N_9244);
nor U9272 (N_9272,N_9234,N_9180);
or U9273 (N_9273,N_9177,N_9169);
nor U9274 (N_9274,N_9128,N_9194);
nor U9275 (N_9275,N_9184,N_9173);
xnor U9276 (N_9276,N_9146,N_9230);
and U9277 (N_9277,N_9195,N_9175);
and U9278 (N_9278,N_9140,N_9187);
and U9279 (N_9279,N_9206,N_9212);
and U9280 (N_9280,N_9138,N_9249);
or U9281 (N_9281,N_9198,N_9141);
nand U9282 (N_9282,N_9125,N_9136);
nor U9283 (N_9283,N_9126,N_9201);
nand U9284 (N_9284,N_9144,N_9127);
xor U9285 (N_9285,N_9157,N_9179);
nor U9286 (N_9286,N_9208,N_9167);
xnor U9287 (N_9287,N_9225,N_9222);
and U9288 (N_9288,N_9193,N_9237);
nor U9289 (N_9289,N_9202,N_9211);
nand U9290 (N_9290,N_9220,N_9248);
xnor U9291 (N_9291,N_9213,N_9183);
or U9292 (N_9292,N_9241,N_9150);
or U9293 (N_9293,N_9239,N_9227);
xnor U9294 (N_9294,N_9154,N_9190);
nor U9295 (N_9295,N_9242,N_9219);
nor U9296 (N_9296,N_9233,N_9172);
nor U9297 (N_9297,N_9137,N_9155);
or U9298 (N_9298,N_9182,N_9133);
and U9299 (N_9299,N_9228,N_9218);
xor U9300 (N_9300,N_9176,N_9164);
xnor U9301 (N_9301,N_9153,N_9148);
or U9302 (N_9302,N_9178,N_9214);
nand U9303 (N_9303,N_9209,N_9200);
xor U9304 (N_9304,N_9151,N_9221);
nor U9305 (N_9305,N_9152,N_9203);
and U9306 (N_9306,N_9247,N_9240);
nor U9307 (N_9307,N_9243,N_9197);
nand U9308 (N_9308,N_9223,N_9229);
nor U9309 (N_9309,N_9192,N_9204);
and U9310 (N_9310,N_9215,N_9217);
xor U9311 (N_9311,N_9166,N_9129);
or U9312 (N_9312,N_9188,N_9220);
and U9313 (N_9313,N_9174,N_9214);
nor U9314 (N_9314,N_9184,N_9148);
or U9315 (N_9315,N_9157,N_9226);
nand U9316 (N_9316,N_9190,N_9225);
or U9317 (N_9317,N_9133,N_9221);
or U9318 (N_9318,N_9239,N_9153);
and U9319 (N_9319,N_9159,N_9244);
xor U9320 (N_9320,N_9187,N_9214);
nor U9321 (N_9321,N_9128,N_9224);
and U9322 (N_9322,N_9175,N_9232);
or U9323 (N_9323,N_9128,N_9231);
xnor U9324 (N_9324,N_9138,N_9185);
or U9325 (N_9325,N_9212,N_9211);
xnor U9326 (N_9326,N_9139,N_9248);
or U9327 (N_9327,N_9244,N_9149);
xor U9328 (N_9328,N_9215,N_9165);
nand U9329 (N_9329,N_9239,N_9234);
nand U9330 (N_9330,N_9198,N_9248);
nand U9331 (N_9331,N_9185,N_9128);
nor U9332 (N_9332,N_9187,N_9240);
and U9333 (N_9333,N_9190,N_9180);
and U9334 (N_9334,N_9215,N_9170);
and U9335 (N_9335,N_9229,N_9237);
nor U9336 (N_9336,N_9229,N_9233);
nor U9337 (N_9337,N_9131,N_9128);
or U9338 (N_9338,N_9145,N_9218);
and U9339 (N_9339,N_9138,N_9154);
nor U9340 (N_9340,N_9180,N_9164);
nor U9341 (N_9341,N_9129,N_9153);
or U9342 (N_9342,N_9215,N_9141);
and U9343 (N_9343,N_9228,N_9194);
or U9344 (N_9344,N_9193,N_9217);
and U9345 (N_9345,N_9205,N_9195);
or U9346 (N_9346,N_9168,N_9204);
and U9347 (N_9347,N_9180,N_9193);
nor U9348 (N_9348,N_9222,N_9160);
xor U9349 (N_9349,N_9182,N_9125);
nor U9350 (N_9350,N_9190,N_9179);
and U9351 (N_9351,N_9138,N_9163);
and U9352 (N_9352,N_9245,N_9169);
or U9353 (N_9353,N_9238,N_9219);
nand U9354 (N_9354,N_9176,N_9184);
or U9355 (N_9355,N_9200,N_9195);
nor U9356 (N_9356,N_9210,N_9174);
nand U9357 (N_9357,N_9219,N_9163);
xnor U9358 (N_9358,N_9153,N_9170);
nor U9359 (N_9359,N_9239,N_9150);
and U9360 (N_9360,N_9243,N_9167);
xnor U9361 (N_9361,N_9159,N_9144);
nor U9362 (N_9362,N_9183,N_9138);
nor U9363 (N_9363,N_9133,N_9194);
nand U9364 (N_9364,N_9196,N_9221);
nand U9365 (N_9365,N_9163,N_9221);
nand U9366 (N_9366,N_9162,N_9140);
nor U9367 (N_9367,N_9188,N_9215);
nor U9368 (N_9368,N_9208,N_9192);
or U9369 (N_9369,N_9229,N_9202);
nor U9370 (N_9370,N_9212,N_9161);
or U9371 (N_9371,N_9173,N_9229);
or U9372 (N_9372,N_9182,N_9191);
nor U9373 (N_9373,N_9171,N_9163);
nor U9374 (N_9374,N_9204,N_9129);
and U9375 (N_9375,N_9335,N_9250);
and U9376 (N_9376,N_9357,N_9346);
or U9377 (N_9377,N_9366,N_9292);
or U9378 (N_9378,N_9362,N_9337);
xnor U9379 (N_9379,N_9350,N_9321);
nor U9380 (N_9380,N_9274,N_9275);
or U9381 (N_9381,N_9301,N_9320);
nor U9382 (N_9382,N_9259,N_9291);
nand U9383 (N_9383,N_9279,N_9343);
and U9384 (N_9384,N_9367,N_9373);
nor U9385 (N_9385,N_9358,N_9371);
or U9386 (N_9386,N_9348,N_9338);
xnor U9387 (N_9387,N_9297,N_9272);
xnor U9388 (N_9388,N_9334,N_9340);
nand U9389 (N_9389,N_9363,N_9264);
nand U9390 (N_9390,N_9290,N_9322);
nand U9391 (N_9391,N_9296,N_9261);
xnor U9392 (N_9392,N_9333,N_9351);
nand U9393 (N_9393,N_9332,N_9323);
and U9394 (N_9394,N_9278,N_9265);
xnor U9395 (N_9395,N_9298,N_9282);
nor U9396 (N_9396,N_9271,N_9276);
and U9397 (N_9397,N_9372,N_9353);
nor U9398 (N_9398,N_9280,N_9328);
nand U9399 (N_9399,N_9314,N_9289);
or U9400 (N_9400,N_9254,N_9303);
or U9401 (N_9401,N_9317,N_9266);
and U9402 (N_9402,N_9341,N_9256);
nor U9403 (N_9403,N_9319,N_9313);
or U9404 (N_9404,N_9326,N_9316);
or U9405 (N_9405,N_9255,N_9309);
and U9406 (N_9406,N_9251,N_9293);
nand U9407 (N_9407,N_9352,N_9349);
or U9408 (N_9408,N_9342,N_9356);
nand U9409 (N_9409,N_9281,N_9252);
xnor U9410 (N_9410,N_9286,N_9325);
xnor U9411 (N_9411,N_9329,N_9263);
nand U9412 (N_9412,N_9344,N_9315);
xor U9413 (N_9413,N_9302,N_9370);
nor U9414 (N_9414,N_9361,N_9300);
or U9415 (N_9415,N_9258,N_9257);
xnor U9416 (N_9416,N_9339,N_9270);
nor U9417 (N_9417,N_9374,N_9304);
or U9418 (N_9418,N_9360,N_9305);
nand U9419 (N_9419,N_9283,N_9308);
and U9420 (N_9420,N_9336,N_9364);
nor U9421 (N_9421,N_9285,N_9307);
nand U9422 (N_9422,N_9354,N_9365);
xnor U9423 (N_9423,N_9345,N_9312);
and U9424 (N_9424,N_9288,N_9273);
nor U9425 (N_9425,N_9347,N_9324);
or U9426 (N_9426,N_9318,N_9355);
xor U9427 (N_9427,N_9369,N_9260);
nor U9428 (N_9428,N_9269,N_9311);
xor U9429 (N_9429,N_9262,N_9287);
and U9430 (N_9430,N_9359,N_9268);
xnor U9431 (N_9431,N_9331,N_9284);
or U9432 (N_9432,N_9327,N_9277);
nand U9433 (N_9433,N_9310,N_9267);
nor U9434 (N_9434,N_9299,N_9294);
xnor U9435 (N_9435,N_9368,N_9306);
and U9436 (N_9436,N_9295,N_9330);
nor U9437 (N_9437,N_9253,N_9313);
and U9438 (N_9438,N_9266,N_9359);
xor U9439 (N_9439,N_9342,N_9276);
or U9440 (N_9440,N_9373,N_9256);
nand U9441 (N_9441,N_9271,N_9315);
or U9442 (N_9442,N_9338,N_9306);
nand U9443 (N_9443,N_9373,N_9291);
nor U9444 (N_9444,N_9252,N_9354);
nand U9445 (N_9445,N_9287,N_9340);
xnor U9446 (N_9446,N_9274,N_9345);
or U9447 (N_9447,N_9314,N_9256);
xor U9448 (N_9448,N_9281,N_9267);
or U9449 (N_9449,N_9333,N_9256);
nand U9450 (N_9450,N_9318,N_9356);
nor U9451 (N_9451,N_9331,N_9369);
or U9452 (N_9452,N_9300,N_9285);
and U9453 (N_9453,N_9275,N_9325);
nor U9454 (N_9454,N_9296,N_9354);
nand U9455 (N_9455,N_9256,N_9285);
and U9456 (N_9456,N_9347,N_9369);
nand U9457 (N_9457,N_9270,N_9304);
or U9458 (N_9458,N_9271,N_9331);
nor U9459 (N_9459,N_9294,N_9373);
nand U9460 (N_9460,N_9282,N_9284);
nand U9461 (N_9461,N_9328,N_9372);
nand U9462 (N_9462,N_9290,N_9294);
or U9463 (N_9463,N_9322,N_9357);
or U9464 (N_9464,N_9263,N_9366);
xor U9465 (N_9465,N_9313,N_9267);
nor U9466 (N_9466,N_9265,N_9306);
nor U9467 (N_9467,N_9277,N_9326);
xnor U9468 (N_9468,N_9259,N_9322);
nand U9469 (N_9469,N_9373,N_9331);
and U9470 (N_9470,N_9287,N_9318);
nor U9471 (N_9471,N_9291,N_9355);
xnor U9472 (N_9472,N_9292,N_9329);
or U9473 (N_9473,N_9313,N_9252);
xor U9474 (N_9474,N_9365,N_9309);
or U9475 (N_9475,N_9301,N_9280);
nand U9476 (N_9476,N_9324,N_9359);
and U9477 (N_9477,N_9360,N_9366);
nand U9478 (N_9478,N_9270,N_9281);
nor U9479 (N_9479,N_9291,N_9334);
nand U9480 (N_9480,N_9340,N_9367);
xor U9481 (N_9481,N_9292,N_9266);
nor U9482 (N_9482,N_9278,N_9293);
xnor U9483 (N_9483,N_9294,N_9301);
nand U9484 (N_9484,N_9343,N_9335);
xor U9485 (N_9485,N_9319,N_9274);
nor U9486 (N_9486,N_9306,N_9333);
nor U9487 (N_9487,N_9336,N_9343);
nand U9488 (N_9488,N_9365,N_9352);
nand U9489 (N_9489,N_9280,N_9286);
or U9490 (N_9490,N_9252,N_9314);
or U9491 (N_9491,N_9339,N_9353);
and U9492 (N_9492,N_9282,N_9320);
or U9493 (N_9493,N_9320,N_9276);
xor U9494 (N_9494,N_9344,N_9368);
and U9495 (N_9495,N_9281,N_9303);
nand U9496 (N_9496,N_9353,N_9290);
or U9497 (N_9497,N_9304,N_9348);
nor U9498 (N_9498,N_9292,N_9323);
nand U9499 (N_9499,N_9276,N_9273);
and U9500 (N_9500,N_9387,N_9410);
xor U9501 (N_9501,N_9375,N_9391);
and U9502 (N_9502,N_9488,N_9386);
or U9503 (N_9503,N_9457,N_9487);
or U9504 (N_9504,N_9443,N_9390);
xor U9505 (N_9505,N_9485,N_9405);
or U9506 (N_9506,N_9409,N_9420);
nand U9507 (N_9507,N_9422,N_9393);
nor U9508 (N_9508,N_9432,N_9465);
nand U9509 (N_9509,N_9445,N_9448);
xor U9510 (N_9510,N_9415,N_9382);
nand U9511 (N_9511,N_9394,N_9392);
nand U9512 (N_9512,N_9498,N_9384);
nor U9513 (N_9513,N_9449,N_9430);
or U9514 (N_9514,N_9404,N_9439);
nand U9515 (N_9515,N_9462,N_9416);
nand U9516 (N_9516,N_9380,N_9414);
and U9517 (N_9517,N_9455,N_9473);
xnor U9518 (N_9518,N_9471,N_9397);
and U9519 (N_9519,N_9381,N_9442);
and U9520 (N_9520,N_9434,N_9383);
nor U9521 (N_9521,N_9427,N_9425);
xor U9522 (N_9522,N_9428,N_9378);
nand U9523 (N_9523,N_9483,N_9472);
xor U9524 (N_9524,N_9419,N_9494);
or U9525 (N_9525,N_9424,N_9401);
nor U9526 (N_9526,N_9389,N_9490);
or U9527 (N_9527,N_9496,N_9499);
and U9528 (N_9528,N_9398,N_9377);
xnor U9529 (N_9529,N_9468,N_9441);
xnor U9530 (N_9530,N_9429,N_9412);
and U9531 (N_9531,N_9385,N_9431);
nand U9532 (N_9532,N_9399,N_9435);
nand U9533 (N_9533,N_9388,N_9453);
xnor U9534 (N_9534,N_9486,N_9406);
xor U9535 (N_9535,N_9400,N_9408);
nor U9536 (N_9536,N_9440,N_9411);
xor U9537 (N_9537,N_9452,N_9477);
xor U9538 (N_9538,N_9493,N_9478);
and U9539 (N_9539,N_9407,N_9470);
or U9540 (N_9540,N_9418,N_9417);
and U9541 (N_9541,N_9451,N_9396);
xor U9542 (N_9542,N_9474,N_9421);
nor U9543 (N_9543,N_9447,N_9479);
or U9544 (N_9544,N_9489,N_9460);
and U9545 (N_9545,N_9454,N_9438);
or U9546 (N_9546,N_9469,N_9463);
nand U9547 (N_9547,N_9459,N_9482);
nor U9548 (N_9548,N_9437,N_9458);
nor U9549 (N_9549,N_9475,N_9402);
xor U9550 (N_9550,N_9395,N_9413);
or U9551 (N_9551,N_9484,N_9497);
and U9552 (N_9552,N_9492,N_9433);
xnor U9553 (N_9553,N_9423,N_9379);
xnor U9554 (N_9554,N_9376,N_9466);
and U9555 (N_9555,N_9456,N_9491);
and U9556 (N_9556,N_9467,N_9444);
nand U9557 (N_9557,N_9450,N_9426);
and U9558 (N_9558,N_9480,N_9481);
and U9559 (N_9559,N_9464,N_9403);
nand U9560 (N_9560,N_9461,N_9495);
or U9561 (N_9561,N_9476,N_9436);
nor U9562 (N_9562,N_9446,N_9487);
or U9563 (N_9563,N_9389,N_9464);
xnor U9564 (N_9564,N_9438,N_9400);
nand U9565 (N_9565,N_9403,N_9491);
xnor U9566 (N_9566,N_9381,N_9499);
nor U9567 (N_9567,N_9421,N_9426);
nand U9568 (N_9568,N_9487,N_9473);
nor U9569 (N_9569,N_9399,N_9455);
and U9570 (N_9570,N_9477,N_9430);
and U9571 (N_9571,N_9492,N_9498);
nand U9572 (N_9572,N_9480,N_9389);
nor U9573 (N_9573,N_9484,N_9399);
and U9574 (N_9574,N_9405,N_9449);
and U9575 (N_9575,N_9478,N_9482);
nor U9576 (N_9576,N_9423,N_9452);
and U9577 (N_9577,N_9403,N_9377);
xor U9578 (N_9578,N_9476,N_9405);
nand U9579 (N_9579,N_9412,N_9463);
nand U9580 (N_9580,N_9378,N_9434);
nor U9581 (N_9581,N_9376,N_9432);
or U9582 (N_9582,N_9385,N_9478);
or U9583 (N_9583,N_9488,N_9485);
nor U9584 (N_9584,N_9459,N_9486);
or U9585 (N_9585,N_9416,N_9433);
and U9586 (N_9586,N_9496,N_9488);
nor U9587 (N_9587,N_9497,N_9481);
or U9588 (N_9588,N_9404,N_9388);
nor U9589 (N_9589,N_9428,N_9418);
xor U9590 (N_9590,N_9453,N_9460);
nand U9591 (N_9591,N_9462,N_9484);
nor U9592 (N_9592,N_9433,N_9423);
nor U9593 (N_9593,N_9377,N_9494);
nor U9594 (N_9594,N_9447,N_9413);
or U9595 (N_9595,N_9453,N_9447);
nand U9596 (N_9596,N_9377,N_9435);
and U9597 (N_9597,N_9439,N_9396);
nor U9598 (N_9598,N_9407,N_9386);
xor U9599 (N_9599,N_9383,N_9381);
nand U9600 (N_9600,N_9387,N_9431);
and U9601 (N_9601,N_9381,N_9385);
and U9602 (N_9602,N_9437,N_9479);
nor U9603 (N_9603,N_9479,N_9481);
nand U9604 (N_9604,N_9480,N_9399);
xnor U9605 (N_9605,N_9481,N_9468);
nor U9606 (N_9606,N_9466,N_9377);
nor U9607 (N_9607,N_9485,N_9402);
or U9608 (N_9608,N_9380,N_9433);
nor U9609 (N_9609,N_9396,N_9436);
xor U9610 (N_9610,N_9416,N_9450);
nor U9611 (N_9611,N_9479,N_9470);
nand U9612 (N_9612,N_9380,N_9401);
or U9613 (N_9613,N_9443,N_9427);
and U9614 (N_9614,N_9417,N_9486);
xnor U9615 (N_9615,N_9389,N_9482);
xor U9616 (N_9616,N_9451,N_9397);
and U9617 (N_9617,N_9424,N_9415);
nand U9618 (N_9618,N_9412,N_9413);
xnor U9619 (N_9619,N_9438,N_9399);
nor U9620 (N_9620,N_9457,N_9471);
nor U9621 (N_9621,N_9396,N_9393);
and U9622 (N_9622,N_9396,N_9435);
and U9623 (N_9623,N_9451,N_9467);
and U9624 (N_9624,N_9448,N_9439);
nand U9625 (N_9625,N_9520,N_9570);
nand U9626 (N_9626,N_9557,N_9586);
nor U9627 (N_9627,N_9555,N_9554);
nand U9628 (N_9628,N_9556,N_9532);
and U9629 (N_9629,N_9596,N_9622);
or U9630 (N_9630,N_9528,N_9572);
xnor U9631 (N_9631,N_9542,N_9519);
and U9632 (N_9632,N_9538,N_9609);
xnor U9633 (N_9633,N_9619,N_9585);
nor U9634 (N_9634,N_9512,N_9503);
nand U9635 (N_9635,N_9568,N_9523);
nand U9636 (N_9636,N_9518,N_9613);
nand U9637 (N_9637,N_9514,N_9560);
nand U9638 (N_9638,N_9620,N_9574);
xor U9639 (N_9639,N_9602,N_9500);
and U9640 (N_9640,N_9505,N_9563);
or U9641 (N_9641,N_9603,N_9534);
xor U9642 (N_9642,N_9616,N_9511);
and U9643 (N_9643,N_9608,N_9583);
xnor U9644 (N_9644,N_9578,N_9584);
nand U9645 (N_9645,N_9546,N_9624);
and U9646 (N_9646,N_9529,N_9567);
xnor U9647 (N_9647,N_9548,N_9615);
xor U9648 (N_9648,N_9604,N_9576);
nor U9649 (N_9649,N_9515,N_9588);
nor U9650 (N_9650,N_9577,N_9531);
nor U9651 (N_9651,N_9595,N_9530);
nor U9652 (N_9652,N_9527,N_9502);
xor U9653 (N_9653,N_9592,N_9552);
nand U9654 (N_9654,N_9564,N_9513);
xor U9655 (N_9655,N_9533,N_9587);
nand U9656 (N_9656,N_9598,N_9593);
or U9657 (N_9657,N_9535,N_9606);
nand U9658 (N_9658,N_9621,N_9580);
nand U9659 (N_9659,N_9521,N_9569);
and U9660 (N_9660,N_9551,N_9575);
nand U9661 (N_9661,N_9562,N_9550);
or U9662 (N_9662,N_9599,N_9507);
nor U9663 (N_9663,N_9510,N_9524);
nand U9664 (N_9664,N_9539,N_9509);
nor U9665 (N_9665,N_9612,N_9571);
or U9666 (N_9666,N_9579,N_9594);
or U9667 (N_9667,N_9541,N_9517);
nor U9668 (N_9668,N_9591,N_9597);
and U9669 (N_9669,N_9544,N_9516);
nand U9670 (N_9670,N_9525,N_9590);
xnor U9671 (N_9671,N_9558,N_9565);
nor U9672 (N_9672,N_9547,N_9566);
nand U9673 (N_9673,N_9553,N_9506);
or U9674 (N_9674,N_9581,N_9561);
and U9675 (N_9675,N_9537,N_9549);
nor U9676 (N_9676,N_9617,N_9508);
or U9677 (N_9677,N_9618,N_9614);
nor U9678 (N_9678,N_9540,N_9589);
nand U9679 (N_9679,N_9543,N_9573);
xor U9680 (N_9680,N_9559,N_9610);
nor U9681 (N_9681,N_9582,N_9607);
xnor U9682 (N_9682,N_9545,N_9526);
and U9683 (N_9683,N_9605,N_9601);
nor U9684 (N_9684,N_9501,N_9600);
nor U9685 (N_9685,N_9522,N_9504);
xnor U9686 (N_9686,N_9611,N_9536);
nand U9687 (N_9687,N_9623,N_9542);
xnor U9688 (N_9688,N_9593,N_9524);
nor U9689 (N_9689,N_9598,N_9564);
xor U9690 (N_9690,N_9587,N_9597);
xor U9691 (N_9691,N_9541,N_9529);
nor U9692 (N_9692,N_9502,N_9523);
nor U9693 (N_9693,N_9521,N_9543);
or U9694 (N_9694,N_9567,N_9621);
xor U9695 (N_9695,N_9623,N_9594);
nand U9696 (N_9696,N_9512,N_9560);
xnor U9697 (N_9697,N_9543,N_9592);
nand U9698 (N_9698,N_9558,N_9614);
nor U9699 (N_9699,N_9504,N_9521);
and U9700 (N_9700,N_9548,N_9533);
or U9701 (N_9701,N_9610,N_9547);
nand U9702 (N_9702,N_9616,N_9572);
nor U9703 (N_9703,N_9525,N_9522);
nand U9704 (N_9704,N_9619,N_9563);
nor U9705 (N_9705,N_9584,N_9527);
or U9706 (N_9706,N_9539,N_9595);
or U9707 (N_9707,N_9517,N_9505);
xnor U9708 (N_9708,N_9554,N_9609);
xnor U9709 (N_9709,N_9607,N_9572);
xor U9710 (N_9710,N_9564,N_9581);
or U9711 (N_9711,N_9509,N_9607);
nand U9712 (N_9712,N_9575,N_9522);
and U9713 (N_9713,N_9507,N_9613);
and U9714 (N_9714,N_9602,N_9522);
or U9715 (N_9715,N_9597,N_9598);
and U9716 (N_9716,N_9527,N_9531);
xor U9717 (N_9717,N_9514,N_9572);
xor U9718 (N_9718,N_9571,N_9509);
or U9719 (N_9719,N_9516,N_9592);
or U9720 (N_9720,N_9587,N_9510);
and U9721 (N_9721,N_9529,N_9615);
nor U9722 (N_9722,N_9590,N_9605);
xor U9723 (N_9723,N_9571,N_9564);
nor U9724 (N_9724,N_9537,N_9525);
nor U9725 (N_9725,N_9585,N_9616);
nor U9726 (N_9726,N_9526,N_9539);
nor U9727 (N_9727,N_9544,N_9530);
nor U9728 (N_9728,N_9505,N_9522);
or U9729 (N_9729,N_9601,N_9602);
nand U9730 (N_9730,N_9543,N_9615);
nor U9731 (N_9731,N_9605,N_9594);
and U9732 (N_9732,N_9549,N_9513);
xor U9733 (N_9733,N_9515,N_9508);
and U9734 (N_9734,N_9500,N_9623);
or U9735 (N_9735,N_9548,N_9513);
xor U9736 (N_9736,N_9579,N_9597);
nand U9737 (N_9737,N_9527,N_9603);
or U9738 (N_9738,N_9593,N_9605);
nor U9739 (N_9739,N_9557,N_9560);
xnor U9740 (N_9740,N_9539,N_9591);
nor U9741 (N_9741,N_9605,N_9521);
nand U9742 (N_9742,N_9520,N_9512);
nor U9743 (N_9743,N_9570,N_9525);
nor U9744 (N_9744,N_9563,N_9503);
or U9745 (N_9745,N_9504,N_9517);
nor U9746 (N_9746,N_9563,N_9564);
nor U9747 (N_9747,N_9560,N_9584);
nor U9748 (N_9748,N_9528,N_9535);
nor U9749 (N_9749,N_9576,N_9536);
nor U9750 (N_9750,N_9660,N_9655);
nand U9751 (N_9751,N_9714,N_9695);
nand U9752 (N_9752,N_9739,N_9653);
xnor U9753 (N_9753,N_9729,N_9633);
or U9754 (N_9754,N_9689,N_9683);
or U9755 (N_9755,N_9646,N_9726);
xnor U9756 (N_9756,N_9686,N_9728);
and U9757 (N_9757,N_9738,N_9740);
nor U9758 (N_9758,N_9648,N_9703);
and U9759 (N_9759,N_9702,N_9743);
xor U9760 (N_9760,N_9654,N_9746);
nor U9761 (N_9761,N_9712,N_9668);
and U9762 (N_9762,N_9667,N_9676);
xnor U9763 (N_9763,N_9677,N_9671);
nor U9764 (N_9764,N_9741,N_9697);
and U9765 (N_9765,N_9720,N_9685);
nor U9766 (N_9766,N_9682,N_9744);
xor U9767 (N_9767,N_9707,N_9625);
or U9768 (N_9768,N_9688,N_9629);
xnor U9769 (N_9769,N_9638,N_9665);
xnor U9770 (N_9770,N_9673,N_9723);
xor U9771 (N_9771,N_9733,N_9631);
nand U9772 (N_9772,N_9672,N_9651);
nand U9773 (N_9773,N_9644,N_9694);
xor U9774 (N_9774,N_9664,N_9642);
and U9775 (N_9775,N_9709,N_9725);
nand U9776 (N_9776,N_9700,N_9663);
nand U9777 (N_9777,N_9630,N_9711);
nor U9778 (N_9778,N_9649,N_9675);
nand U9779 (N_9779,N_9666,N_9734);
xor U9780 (N_9780,N_9639,N_9716);
nand U9781 (N_9781,N_9724,N_9742);
nor U9782 (N_9782,N_9730,N_9745);
xnor U9783 (N_9783,N_9628,N_9719);
and U9784 (N_9784,N_9731,N_9636);
nor U9785 (N_9785,N_9627,N_9735);
and U9786 (N_9786,N_9749,N_9705);
or U9787 (N_9787,N_9715,N_9698);
xnor U9788 (N_9788,N_9737,N_9732);
or U9789 (N_9789,N_9662,N_9658);
and U9790 (N_9790,N_9652,N_9722);
or U9791 (N_9791,N_9647,N_9721);
xnor U9792 (N_9792,N_9659,N_9706);
nand U9793 (N_9793,N_9693,N_9661);
nand U9794 (N_9794,N_9708,N_9637);
or U9795 (N_9795,N_9687,N_9670);
nand U9796 (N_9796,N_9710,N_9684);
and U9797 (N_9797,N_9690,N_9680);
nand U9798 (N_9798,N_9643,N_9634);
xnor U9799 (N_9799,N_9645,N_9713);
and U9800 (N_9800,N_9626,N_9747);
or U9801 (N_9801,N_9656,N_9704);
or U9802 (N_9802,N_9635,N_9679);
and U9803 (N_9803,N_9692,N_9727);
nand U9804 (N_9804,N_9641,N_9736);
xnor U9805 (N_9805,N_9640,N_9650);
and U9806 (N_9806,N_9669,N_9699);
nand U9807 (N_9807,N_9674,N_9678);
or U9808 (N_9808,N_9748,N_9632);
and U9809 (N_9809,N_9696,N_9701);
nor U9810 (N_9810,N_9691,N_9717);
nor U9811 (N_9811,N_9681,N_9657);
and U9812 (N_9812,N_9718,N_9673);
or U9813 (N_9813,N_9699,N_9650);
and U9814 (N_9814,N_9725,N_9683);
nand U9815 (N_9815,N_9713,N_9741);
or U9816 (N_9816,N_9727,N_9653);
nor U9817 (N_9817,N_9743,N_9691);
and U9818 (N_9818,N_9663,N_9708);
xor U9819 (N_9819,N_9722,N_9651);
and U9820 (N_9820,N_9731,N_9720);
and U9821 (N_9821,N_9749,N_9746);
or U9822 (N_9822,N_9726,N_9747);
and U9823 (N_9823,N_9644,N_9654);
xnor U9824 (N_9824,N_9643,N_9693);
and U9825 (N_9825,N_9627,N_9730);
and U9826 (N_9826,N_9706,N_9735);
or U9827 (N_9827,N_9665,N_9673);
nor U9828 (N_9828,N_9688,N_9656);
and U9829 (N_9829,N_9670,N_9714);
nand U9830 (N_9830,N_9733,N_9728);
nor U9831 (N_9831,N_9748,N_9695);
nand U9832 (N_9832,N_9656,N_9662);
nor U9833 (N_9833,N_9653,N_9661);
nand U9834 (N_9834,N_9651,N_9731);
nor U9835 (N_9835,N_9715,N_9631);
xnor U9836 (N_9836,N_9667,N_9652);
xor U9837 (N_9837,N_9741,N_9677);
and U9838 (N_9838,N_9743,N_9687);
or U9839 (N_9839,N_9747,N_9638);
nor U9840 (N_9840,N_9659,N_9745);
xnor U9841 (N_9841,N_9662,N_9645);
nand U9842 (N_9842,N_9731,N_9724);
nand U9843 (N_9843,N_9720,N_9710);
xor U9844 (N_9844,N_9674,N_9676);
xnor U9845 (N_9845,N_9705,N_9681);
xnor U9846 (N_9846,N_9629,N_9685);
and U9847 (N_9847,N_9689,N_9679);
nand U9848 (N_9848,N_9628,N_9635);
or U9849 (N_9849,N_9733,N_9674);
nor U9850 (N_9850,N_9714,N_9653);
xor U9851 (N_9851,N_9662,N_9698);
xor U9852 (N_9852,N_9687,N_9634);
nor U9853 (N_9853,N_9714,N_9657);
or U9854 (N_9854,N_9706,N_9670);
xor U9855 (N_9855,N_9719,N_9731);
xnor U9856 (N_9856,N_9664,N_9676);
xor U9857 (N_9857,N_9739,N_9738);
and U9858 (N_9858,N_9686,N_9707);
or U9859 (N_9859,N_9644,N_9735);
or U9860 (N_9860,N_9748,N_9746);
and U9861 (N_9861,N_9703,N_9733);
nand U9862 (N_9862,N_9662,N_9744);
nor U9863 (N_9863,N_9658,N_9737);
and U9864 (N_9864,N_9639,N_9737);
xnor U9865 (N_9865,N_9724,N_9713);
or U9866 (N_9866,N_9739,N_9704);
nand U9867 (N_9867,N_9641,N_9651);
xor U9868 (N_9868,N_9672,N_9734);
nand U9869 (N_9869,N_9693,N_9732);
xor U9870 (N_9870,N_9738,N_9638);
nor U9871 (N_9871,N_9706,N_9679);
xnor U9872 (N_9872,N_9657,N_9697);
nor U9873 (N_9873,N_9676,N_9703);
or U9874 (N_9874,N_9669,N_9704);
nand U9875 (N_9875,N_9838,N_9835);
xnor U9876 (N_9876,N_9834,N_9827);
and U9877 (N_9877,N_9792,N_9860);
xor U9878 (N_9878,N_9820,N_9762);
xnor U9879 (N_9879,N_9751,N_9794);
nor U9880 (N_9880,N_9787,N_9760);
nor U9881 (N_9881,N_9874,N_9831);
nor U9882 (N_9882,N_9757,N_9821);
nand U9883 (N_9883,N_9864,N_9829);
or U9884 (N_9884,N_9815,N_9856);
or U9885 (N_9885,N_9858,N_9778);
xor U9886 (N_9886,N_9795,N_9768);
xnor U9887 (N_9887,N_9853,N_9840);
xnor U9888 (N_9888,N_9847,N_9799);
nor U9889 (N_9889,N_9818,N_9822);
nand U9890 (N_9890,N_9784,N_9788);
and U9891 (N_9891,N_9803,N_9791);
xor U9892 (N_9892,N_9767,N_9810);
and U9893 (N_9893,N_9753,N_9766);
xor U9894 (N_9894,N_9872,N_9867);
nand U9895 (N_9895,N_9841,N_9845);
nand U9896 (N_9896,N_9801,N_9846);
or U9897 (N_9897,N_9862,N_9855);
or U9898 (N_9898,N_9804,N_9756);
nand U9899 (N_9899,N_9851,N_9837);
nor U9900 (N_9900,N_9871,N_9844);
nand U9901 (N_9901,N_9849,N_9780);
nor U9902 (N_9902,N_9868,N_9836);
nor U9903 (N_9903,N_9785,N_9824);
nor U9904 (N_9904,N_9873,N_9865);
nand U9905 (N_9905,N_9802,N_9832);
xnor U9906 (N_9906,N_9752,N_9777);
nand U9907 (N_9907,N_9839,N_9786);
or U9908 (N_9908,N_9861,N_9796);
nor U9909 (N_9909,N_9869,N_9814);
or U9910 (N_9910,N_9826,N_9859);
xor U9911 (N_9911,N_9812,N_9819);
nand U9912 (N_9912,N_9800,N_9805);
and U9913 (N_9913,N_9789,N_9825);
nor U9914 (N_9914,N_9809,N_9823);
nand U9915 (N_9915,N_9807,N_9813);
xnor U9916 (N_9916,N_9830,N_9770);
nor U9917 (N_9917,N_9764,N_9863);
xnor U9918 (N_9918,N_9772,N_9776);
xnor U9919 (N_9919,N_9833,N_9828);
nand U9920 (N_9920,N_9870,N_9866);
nand U9921 (N_9921,N_9852,N_9843);
or U9922 (N_9922,N_9765,N_9816);
xnor U9923 (N_9923,N_9793,N_9771);
and U9924 (N_9924,N_9783,N_9779);
nand U9925 (N_9925,N_9842,N_9782);
nand U9926 (N_9926,N_9773,N_9769);
and U9927 (N_9927,N_9754,N_9857);
or U9928 (N_9928,N_9798,N_9755);
or U9929 (N_9929,N_9758,N_9817);
xor U9930 (N_9930,N_9811,N_9774);
nand U9931 (N_9931,N_9759,N_9808);
xor U9932 (N_9932,N_9781,N_9790);
xnor U9933 (N_9933,N_9848,N_9806);
nor U9934 (N_9934,N_9775,N_9750);
nor U9935 (N_9935,N_9763,N_9854);
xor U9936 (N_9936,N_9761,N_9797);
or U9937 (N_9937,N_9850,N_9756);
nand U9938 (N_9938,N_9815,N_9760);
xor U9939 (N_9939,N_9771,N_9807);
or U9940 (N_9940,N_9833,N_9836);
or U9941 (N_9941,N_9833,N_9819);
nor U9942 (N_9942,N_9838,N_9822);
nor U9943 (N_9943,N_9798,N_9825);
or U9944 (N_9944,N_9769,N_9834);
and U9945 (N_9945,N_9826,N_9872);
nor U9946 (N_9946,N_9783,N_9825);
xnor U9947 (N_9947,N_9838,N_9761);
nand U9948 (N_9948,N_9814,N_9808);
xnor U9949 (N_9949,N_9788,N_9807);
nand U9950 (N_9950,N_9822,N_9849);
and U9951 (N_9951,N_9753,N_9760);
and U9952 (N_9952,N_9795,N_9857);
and U9953 (N_9953,N_9789,N_9872);
xor U9954 (N_9954,N_9764,N_9835);
nand U9955 (N_9955,N_9781,N_9842);
nor U9956 (N_9956,N_9837,N_9865);
nor U9957 (N_9957,N_9829,N_9839);
nor U9958 (N_9958,N_9770,N_9834);
nand U9959 (N_9959,N_9799,N_9831);
xnor U9960 (N_9960,N_9850,N_9817);
or U9961 (N_9961,N_9870,N_9804);
and U9962 (N_9962,N_9760,N_9755);
nand U9963 (N_9963,N_9861,N_9841);
nor U9964 (N_9964,N_9862,N_9763);
nor U9965 (N_9965,N_9854,N_9820);
nor U9966 (N_9966,N_9847,N_9806);
or U9967 (N_9967,N_9868,N_9841);
or U9968 (N_9968,N_9830,N_9779);
nand U9969 (N_9969,N_9795,N_9834);
and U9970 (N_9970,N_9769,N_9850);
nand U9971 (N_9971,N_9796,N_9791);
or U9972 (N_9972,N_9811,N_9760);
nand U9973 (N_9973,N_9853,N_9813);
or U9974 (N_9974,N_9789,N_9807);
or U9975 (N_9975,N_9775,N_9838);
nor U9976 (N_9976,N_9868,N_9780);
or U9977 (N_9977,N_9827,N_9840);
or U9978 (N_9978,N_9791,N_9857);
nand U9979 (N_9979,N_9781,N_9843);
nand U9980 (N_9980,N_9832,N_9792);
and U9981 (N_9981,N_9795,N_9757);
nand U9982 (N_9982,N_9758,N_9812);
xnor U9983 (N_9983,N_9795,N_9784);
xnor U9984 (N_9984,N_9787,N_9757);
or U9985 (N_9985,N_9783,N_9808);
and U9986 (N_9986,N_9845,N_9820);
and U9987 (N_9987,N_9798,N_9838);
and U9988 (N_9988,N_9872,N_9821);
xnor U9989 (N_9989,N_9838,N_9795);
and U9990 (N_9990,N_9854,N_9764);
or U9991 (N_9991,N_9869,N_9806);
nor U9992 (N_9992,N_9829,N_9788);
nor U9993 (N_9993,N_9827,N_9832);
xnor U9994 (N_9994,N_9755,N_9873);
xnor U9995 (N_9995,N_9788,N_9772);
nor U9996 (N_9996,N_9777,N_9859);
nand U9997 (N_9997,N_9771,N_9861);
xnor U9998 (N_9998,N_9818,N_9838);
or U9999 (N_9999,N_9794,N_9874);
and U10000 (N_10000,N_9910,N_9891);
xor U10001 (N_10001,N_9917,N_9977);
and U10002 (N_10002,N_9897,N_9954);
and U10003 (N_10003,N_9972,N_9939);
and U10004 (N_10004,N_9936,N_9992);
xor U10005 (N_10005,N_9906,N_9945);
or U10006 (N_10006,N_9919,N_9914);
and U10007 (N_10007,N_9997,N_9928);
nand U10008 (N_10008,N_9985,N_9941);
or U10009 (N_10009,N_9990,N_9920);
or U10010 (N_10010,N_9966,N_9973);
and U10011 (N_10011,N_9896,N_9912);
and U10012 (N_10012,N_9884,N_9958);
and U10013 (N_10013,N_9875,N_9882);
and U10014 (N_10014,N_9894,N_9902);
nand U10015 (N_10015,N_9916,N_9994);
nor U10016 (N_10016,N_9984,N_9976);
nor U10017 (N_10017,N_9993,N_9921);
nor U10018 (N_10018,N_9981,N_9944);
nand U10019 (N_10019,N_9938,N_9932);
and U10020 (N_10020,N_9978,N_9905);
or U10021 (N_10021,N_9886,N_9948);
xor U10022 (N_10022,N_9898,N_9927);
and U10023 (N_10023,N_9946,N_9960);
xnor U10024 (N_10024,N_9970,N_9949);
nand U10025 (N_10025,N_9913,N_9965);
and U10026 (N_10026,N_9943,N_9934);
xor U10027 (N_10027,N_9952,N_9893);
or U10028 (N_10028,N_9933,N_9961);
and U10029 (N_10029,N_9989,N_9996);
or U10030 (N_10030,N_9879,N_9881);
nand U10031 (N_10031,N_9931,N_9940);
and U10032 (N_10032,N_9876,N_9889);
xnor U10033 (N_10033,N_9963,N_9915);
xor U10034 (N_10034,N_9979,N_9967);
nand U10035 (N_10035,N_9959,N_9903);
nor U10036 (N_10036,N_9877,N_9987);
nand U10037 (N_10037,N_9901,N_9925);
and U10038 (N_10038,N_9974,N_9899);
and U10039 (N_10039,N_9995,N_9924);
or U10040 (N_10040,N_9922,N_9918);
xor U10041 (N_10041,N_9892,N_9956);
xor U10042 (N_10042,N_9982,N_9980);
xor U10043 (N_10043,N_9937,N_9975);
nor U10044 (N_10044,N_9929,N_9880);
or U10045 (N_10045,N_9986,N_9900);
or U10046 (N_10046,N_9999,N_9926);
and U10047 (N_10047,N_9878,N_9907);
nor U10048 (N_10048,N_9935,N_9955);
or U10049 (N_10049,N_9968,N_9950);
nor U10050 (N_10050,N_9953,N_9969);
xnor U10051 (N_10051,N_9883,N_9962);
or U10052 (N_10052,N_9942,N_9887);
or U10053 (N_10053,N_9923,N_9983);
or U10054 (N_10054,N_9911,N_9988);
xnor U10055 (N_10055,N_9971,N_9904);
xor U10056 (N_10056,N_9947,N_9964);
xor U10057 (N_10057,N_9890,N_9957);
xnor U10058 (N_10058,N_9909,N_9908);
or U10059 (N_10059,N_9885,N_9930);
and U10060 (N_10060,N_9888,N_9895);
and U10061 (N_10061,N_9951,N_9991);
and U10062 (N_10062,N_9998,N_9962);
nor U10063 (N_10063,N_9885,N_9923);
nand U10064 (N_10064,N_9967,N_9880);
and U10065 (N_10065,N_9991,N_9973);
nand U10066 (N_10066,N_9985,N_9957);
or U10067 (N_10067,N_9964,N_9999);
and U10068 (N_10068,N_9932,N_9877);
xor U10069 (N_10069,N_9973,N_9889);
xor U10070 (N_10070,N_9950,N_9991);
nor U10071 (N_10071,N_9954,N_9927);
and U10072 (N_10072,N_9959,N_9905);
and U10073 (N_10073,N_9967,N_9894);
and U10074 (N_10074,N_9934,N_9965);
and U10075 (N_10075,N_9912,N_9994);
and U10076 (N_10076,N_9937,N_9881);
xor U10077 (N_10077,N_9964,N_9986);
and U10078 (N_10078,N_9946,N_9931);
nand U10079 (N_10079,N_9963,N_9999);
xor U10080 (N_10080,N_9984,N_9971);
and U10081 (N_10081,N_9879,N_9989);
or U10082 (N_10082,N_9994,N_9998);
xor U10083 (N_10083,N_9998,N_9984);
and U10084 (N_10084,N_9943,N_9968);
nand U10085 (N_10085,N_9889,N_9927);
nor U10086 (N_10086,N_9896,N_9964);
nor U10087 (N_10087,N_9950,N_9898);
nor U10088 (N_10088,N_9910,N_9965);
nor U10089 (N_10089,N_9875,N_9957);
xor U10090 (N_10090,N_9969,N_9975);
and U10091 (N_10091,N_9952,N_9915);
and U10092 (N_10092,N_9941,N_9971);
and U10093 (N_10093,N_9935,N_9975);
nor U10094 (N_10094,N_9978,N_9903);
nand U10095 (N_10095,N_9919,N_9963);
nand U10096 (N_10096,N_9963,N_9883);
nor U10097 (N_10097,N_9975,N_9972);
nor U10098 (N_10098,N_9956,N_9879);
nand U10099 (N_10099,N_9939,N_9982);
or U10100 (N_10100,N_9936,N_9895);
or U10101 (N_10101,N_9990,N_9966);
and U10102 (N_10102,N_9964,N_9886);
nor U10103 (N_10103,N_9953,N_9908);
nand U10104 (N_10104,N_9889,N_9911);
nor U10105 (N_10105,N_9918,N_9958);
nor U10106 (N_10106,N_9970,N_9969);
or U10107 (N_10107,N_9994,N_9933);
xnor U10108 (N_10108,N_9958,N_9910);
and U10109 (N_10109,N_9918,N_9952);
xor U10110 (N_10110,N_9944,N_9887);
nor U10111 (N_10111,N_9948,N_9913);
xor U10112 (N_10112,N_9950,N_9980);
or U10113 (N_10113,N_9931,N_9995);
xor U10114 (N_10114,N_9951,N_9998);
nor U10115 (N_10115,N_9972,N_9876);
xor U10116 (N_10116,N_9947,N_9924);
nand U10117 (N_10117,N_9959,N_9955);
or U10118 (N_10118,N_9941,N_9899);
xor U10119 (N_10119,N_9946,N_9948);
nor U10120 (N_10120,N_9948,N_9878);
nand U10121 (N_10121,N_9992,N_9977);
xor U10122 (N_10122,N_9978,N_9990);
nand U10123 (N_10123,N_9968,N_9915);
and U10124 (N_10124,N_9980,N_9898);
nor U10125 (N_10125,N_10117,N_10053);
or U10126 (N_10126,N_10064,N_10045);
or U10127 (N_10127,N_10021,N_10005);
xnor U10128 (N_10128,N_10088,N_10016);
and U10129 (N_10129,N_10107,N_10037);
nand U10130 (N_10130,N_10119,N_10039);
and U10131 (N_10131,N_10050,N_10017);
nand U10132 (N_10132,N_10000,N_10028);
xnor U10133 (N_10133,N_10108,N_10047);
nand U10134 (N_10134,N_10043,N_10111);
xor U10135 (N_10135,N_10094,N_10054);
and U10136 (N_10136,N_10058,N_10080);
or U10137 (N_10137,N_10076,N_10085);
and U10138 (N_10138,N_10022,N_10015);
nand U10139 (N_10139,N_10035,N_10074);
or U10140 (N_10140,N_10031,N_10065);
and U10141 (N_10141,N_10072,N_10120);
nand U10142 (N_10142,N_10046,N_10038);
or U10143 (N_10143,N_10008,N_10036);
nand U10144 (N_10144,N_10123,N_10096);
xor U10145 (N_10145,N_10114,N_10098);
nand U10146 (N_10146,N_10004,N_10118);
nand U10147 (N_10147,N_10124,N_10082);
xnor U10148 (N_10148,N_10025,N_10026);
nand U10149 (N_10149,N_10056,N_10112);
or U10150 (N_10150,N_10014,N_10121);
and U10151 (N_10151,N_10027,N_10049);
xnor U10152 (N_10152,N_10048,N_10079);
nor U10153 (N_10153,N_10100,N_10083);
xnor U10154 (N_10154,N_10044,N_10009);
nor U10155 (N_10155,N_10067,N_10069);
nand U10156 (N_10156,N_10062,N_10059);
nor U10157 (N_10157,N_10023,N_10055);
or U10158 (N_10158,N_10078,N_10024);
xor U10159 (N_10159,N_10066,N_10018);
xnor U10160 (N_10160,N_10075,N_10093);
nand U10161 (N_10161,N_10020,N_10040);
nand U10162 (N_10162,N_10113,N_10051);
nand U10163 (N_10163,N_10104,N_10095);
xor U10164 (N_10164,N_10092,N_10010);
xnor U10165 (N_10165,N_10032,N_10068);
nor U10166 (N_10166,N_10102,N_10110);
nor U10167 (N_10167,N_10077,N_10073);
nand U10168 (N_10168,N_10070,N_10099);
and U10169 (N_10169,N_10097,N_10030);
nand U10170 (N_10170,N_10116,N_10029);
and U10171 (N_10171,N_10071,N_10101);
nand U10172 (N_10172,N_10081,N_10011);
or U10173 (N_10173,N_10061,N_10003);
xor U10174 (N_10174,N_10091,N_10105);
xor U10175 (N_10175,N_10109,N_10013);
or U10176 (N_10176,N_10103,N_10052);
nor U10177 (N_10177,N_10019,N_10122);
and U10178 (N_10178,N_10041,N_10002);
nand U10179 (N_10179,N_10090,N_10060);
nor U10180 (N_10180,N_10042,N_10033);
xor U10181 (N_10181,N_10084,N_10086);
or U10182 (N_10182,N_10115,N_10007);
or U10183 (N_10183,N_10057,N_10034);
nand U10184 (N_10184,N_10089,N_10106);
and U10185 (N_10185,N_10087,N_10012);
nor U10186 (N_10186,N_10006,N_10001);
or U10187 (N_10187,N_10063,N_10023);
xor U10188 (N_10188,N_10062,N_10029);
or U10189 (N_10189,N_10037,N_10115);
and U10190 (N_10190,N_10089,N_10097);
xor U10191 (N_10191,N_10100,N_10017);
nor U10192 (N_10192,N_10072,N_10117);
and U10193 (N_10193,N_10060,N_10100);
and U10194 (N_10194,N_10086,N_10026);
nand U10195 (N_10195,N_10087,N_10088);
nand U10196 (N_10196,N_10106,N_10042);
or U10197 (N_10197,N_10013,N_10085);
or U10198 (N_10198,N_10052,N_10034);
and U10199 (N_10199,N_10003,N_10031);
or U10200 (N_10200,N_10119,N_10005);
and U10201 (N_10201,N_10100,N_10028);
nand U10202 (N_10202,N_10033,N_10080);
and U10203 (N_10203,N_10106,N_10061);
or U10204 (N_10204,N_10067,N_10052);
nor U10205 (N_10205,N_10121,N_10089);
nand U10206 (N_10206,N_10116,N_10028);
nand U10207 (N_10207,N_10015,N_10063);
and U10208 (N_10208,N_10087,N_10024);
and U10209 (N_10209,N_10031,N_10053);
xnor U10210 (N_10210,N_10053,N_10050);
and U10211 (N_10211,N_10004,N_10079);
nor U10212 (N_10212,N_10020,N_10012);
nor U10213 (N_10213,N_10086,N_10115);
or U10214 (N_10214,N_10055,N_10066);
xor U10215 (N_10215,N_10081,N_10031);
nor U10216 (N_10216,N_10108,N_10016);
xor U10217 (N_10217,N_10073,N_10011);
nor U10218 (N_10218,N_10115,N_10033);
or U10219 (N_10219,N_10115,N_10103);
and U10220 (N_10220,N_10113,N_10021);
and U10221 (N_10221,N_10077,N_10005);
nor U10222 (N_10222,N_10105,N_10044);
and U10223 (N_10223,N_10105,N_10040);
or U10224 (N_10224,N_10049,N_10020);
xor U10225 (N_10225,N_10058,N_10049);
xnor U10226 (N_10226,N_10038,N_10007);
and U10227 (N_10227,N_10046,N_10052);
or U10228 (N_10228,N_10096,N_10114);
nand U10229 (N_10229,N_10022,N_10098);
xnor U10230 (N_10230,N_10087,N_10031);
nor U10231 (N_10231,N_10074,N_10007);
and U10232 (N_10232,N_10089,N_10044);
nor U10233 (N_10233,N_10102,N_10029);
xnor U10234 (N_10234,N_10074,N_10121);
xnor U10235 (N_10235,N_10118,N_10030);
nor U10236 (N_10236,N_10062,N_10016);
and U10237 (N_10237,N_10088,N_10009);
and U10238 (N_10238,N_10051,N_10073);
and U10239 (N_10239,N_10084,N_10096);
xnor U10240 (N_10240,N_10004,N_10092);
and U10241 (N_10241,N_10113,N_10042);
nor U10242 (N_10242,N_10081,N_10088);
nor U10243 (N_10243,N_10096,N_10016);
or U10244 (N_10244,N_10045,N_10099);
xor U10245 (N_10245,N_10037,N_10108);
or U10246 (N_10246,N_10034,N_10061);
and U10247 (N_10247,N_10095,N_10079);
xnor U10248 (N_10248,N_10013,N_10006);
xor U10249 (N_10249,N_10064,N_10081);
or U10250 (N_10250,N_10216,N_10125);
and U10251 (N_10251,N_10209,N_10208);
xor U10252 (N_10252,N_10132,N_10186);
nor U10253 (N_10253,N_10225,N_10135);
and U10254 (N_10254,N_10196,N_10138);
nand U10255 (N_10255,N_10232,N_10222);
or U10256 (N_10256,N_10139,N_10183);
and U10257 (N_10257,N_10218,N_10205);
or U10258 (N_10258,N_10238,N_10167);
nor U10259 (N_10259,N_10174,N_10243);
or U10260 (N_10260,N_10226,N_10145);
and U10261 (N_10261,N_10236,N_10131);
xnor U10262 (N_10262,N_10199,N_10206);
nor U10263 (N_10263,N_10239,N_10136);
nor U10264 (N_10264,N_10134,N_10237);
nand U10265 (N_10265,N_10152,N_10148);
or U10266 (N_10266,N_10143,N_10129);
nor U10267 (N_10267,N_10172,N_10140);
xor U10268 (N_10268,N_10191,N_10149);
and U10269 (N_10269,N_10197,N_10128);
or U10270 (N_10270,N_10188,N_10221);
and U10271 (N_10271,N_10171,N_10185);
and U10272 (N_10272,N_10173,N_10126);
nand U10273 (N_10273,N_10200,N_10224);
or U10274 (N_10274,N_10147,N_10141);
nand U10275 (N_10275,N_10195,N_10157);
or U10276 (N_10276,N_10220,N_10207);
nor U10277 (N_10277,N_10144,N_10151);
xnor U10278 (N_10278,N_10214,N_10210);
nor U10279 (N_10279,N_10170,N_10158);
xor U10280 (N_10280,N_10219,N_10211);
and U10281 (N_10281,N_10166,N_10180);
xor U10282 (N_10282,N_10212,N_10228);
nand U10283 (N_10283,N_10181,N_10182);
and U10284 (N_10284,N_10241,N_10202);
or U10285 (N_10285,N_10246,N_10133);
xnor U10286 (N_10286,N_10184,N_10130);
nor U10287 (N_10287,N_10194,N_10189);
nand U10288 (N_10288,N_10233,N_10137);
and U10289 (N_10289,N_10192,N_10235);
xnor U10290 (N_10290,N_10244,N_10247);
nand U10291 (N_10291,N_10150,N_10154);
nor U10292 (N_10292,N_10201,N_10217);
nor U10293 (N_10293,N_10160,N_10142);
and U10294 (N_10294,N_10156,N_10175);
nand U10295 (N_10295,N_10234,N_10155);
xnor U10296 (N_10296,N_10146,N_10163);
nand U10297 (N_10297,N_10168,N_10153);
nor U10298 (N_10298,N_10162,N_10230);
xnor U10299 (N_10299,N_10240,N_10213);
and U10300 (N_10300,N_10215,N_10178);
xnor U10301 (N_10301,N_10245,N_10193);
or U10302 (N_10302,N_10165,N_10229);
xor U10303 (N_10303,N_10176,N_10190);
or U10304 (N_10304,N_10127,N_10204);
nor U10305 (N_10305,N_10248,N_10187);
or U10306 (N_10306,N_10161,N_10198);
nand U10307 (N_10307,N_10223,N_10179);
nand U10308 (N_10308,N_10249,N_10231);
nand U10309 (N_10309,N_10159,N_10169);
nand U10310 (N_10310,N_10227,N_10177);
or U10311 (N_10311,N_10164,N_10242);
nor U10312 (N_10312,N_10203,N_10179);
or U10313 (N_10313,N_10145,N_10204);
xor U10314 (N_10314,N_10192,N_10169);
and U10315 (N_10315,N_10203,N_10197);
nor U10316 (N_10316,N_10136,N_10225);
nor U10317 (N_10317,N_10217,N_10157);
nor U10318 (N_10318,N_10136,N_10200);
nand U10319 (N_10319,N_10175,N_10165);
nand U10320 (N_10320,N_10225,N_10189);
or U10321 (N_10321,N_10195,N_10193);
xor U10322 (N_10322,N_10240,N_10243);
nor U10323 (N_10323,N_10221,N_10174);
nand U10324 (N_10324,N_10135,N_10159);
nand U10325 (N_10325,N_10205,N_10193);
nand U10326 (N_10326,N_10144,N_10231);
nand U10327 (N_10327,N_10134,N_10239);
or U10328 (N_10328,N_10136,N_10145);
and U10329 (N_10329,N_10200,N_10245);
or U10330 (N_10330,N_10245,N_10218);
or U10331 (N_10331,N_10174,N_10135);
xor U10332 (N_10332,N_10135,N_10217);
or U10333 (N_10333,N_10226,N_10187);
and U10334 (N_10334,N_10145,N_10191);
nor U10335 (N_10335,N_10148,N_10206);
xor U10336 (N_10336,N_10198,N_10195);
xnor U10337 (N_10337,N_10135,N_10145);
xnor U10338 (N_10338,N_10150,N_10237);
and U10339 (N_10339,N_10237,N_10169);
or U10340 (N_10340,N_10236,N_10238);
nand U10341 (N_10341,N_10196,N_10218);
nor U10342 (N_10342,N_10233,N_10147);
and U10343 (N_10343,N_10219,N_10161);
and U10344 (N_10344,N_10233,N_10190);
nand U10345 (N_10345,N_10133,N_10126);
and U10346 (N_10346,N_10226,N_10199);
nor U10347 (N_10347,N_10156,N_10212);
xor U10348 (N_10348,N_10157,N_10186);
nor U10349 (N_10349,N_10129,N_10145);
or U10350 (N_10350,N_10152,N_10169);
and U10351 (N_10351,N_10195,N_10148);
and U10352 (N_10352,N_10150,N_10232);
xnor U10353 (N_10353,N_10232,N_10212);
nor U10354 (N_10354,N_10233,N_10192);
and U10355 (N_10355,N_10202,N_10159);
nand U10356 (N_10356,N_10128,N_10167);
or U10357 (N_10357,N_10217,N_10125);
or U10358 (N_10358,N_10222,N_10236);
xnor U10359 (N_10359,N_10235,N_10147);
and U10360 (N_10360,N_10151,N_10142);
nor U10361 (N_10361,N_10220,N_10174);
or U10362 (N_10362,N_10202,N_10207);
or U10363 (N_10363,N_10159,N_10179);
or U10364 (N_10364,N_10182,N_10242);
and U10365 (N_10365,N_10163,N_10248);
and U10366 (N_10366,N_10140,N_10165);
nor U10367 (N_10367,N_10176,N_10130);
or U10368 (N_10368,N_10229,N_10146);
xnor U10369 (N_10369,N_10127,N_10191);
xor U10370 (N_10370,N_10199,N_10245);
or U10371 (N_10371,N_10161,N_10169);
nand U10372 (N_10372,N_10202,N_10201);
or U10373 (N_10373,N_10127,N_10209);
nand U10374 (N_10374,N_10231,N_10155);
nand U10375 (N_10375,N_10302,N_10295);
xnor U10376 (N_10376,N_10284,N_10271);
and U10377 (N_10377,N_10371,N_10286);
or U10378 (N_10378,N_10283,N_10277);
nor U10379 (N_10379,N_10255,N_10280);
or U10380 (N_10380,N_10330,N_10344);
or U10381 (N_10381,N_10287,N_10362);
nor U10382 (N_10382,N_10356,N_10257);
xnor U10383 (N_10383,N_10253,N_10372);
nor U10384 (N_10384,N_10279,N_10296);
or U10385 (N_10385,N_10343,N_10348);
nand U10386 (N_10386,N_10363,N_10359);
and U10387 (N_10387,N_10297,N_10350);
nor U10388 (N_10388,N_10336,N_10335);
and U10389 (N_10389,N_10264,N_10262);
nand U10390 (N_10390,N_10346,N_10364);
nor U10391 (N_10391,N_10258,N_10339);
nand U10392 (N_10392,N_10268,N_10265);
or U10393 (N_10393,N_10261,N_10332);
and U10394 (N_10394,N_10345,N_10254);
xnor U10395 (N_10395,N_10360,N_10349);
and U10396 (N_10396,N_10316,N_10355);
and U10397 (N_10397,N_10294,N_10338);
nand U10398 (N_10398,N_10317,N_10278);
and U10399 (N_10399,N_10337,N_10276);
nand U10400 (N_10400,N_10370,N_10329);
nor U10401 (N_10401,N_10299,N_10288);
xnor U10402 (N_10402,N_10351,N_10366);
nand U10403 (N_10403,N_10301,N_10291);
or U10404 (N_10404,N_10310,N_10365);
and U10405 (N_10405,N_10320,N_10334);
or U10406 (N_10406,N_10282,N_10252);
or U10407 (N_10407,N_10314,N_10303);
xnor U10408 (N_10408,N_10260,N_10251);
or U10409 (N_10409,N_10324,N_10298);
nor U10410 (N_10410,N_10321,N_10341);
and U10411 (N_10411,N_10367,N_10275);
nor U10412 (N_10412,N_10318,N_10269);
and U10413 (N_10413,N_10358,N_10309);
or U10414 (N_10414,N_10290,N_10289);
or U10415 (N_10415,N_10304,N_10307);
nor U10416 (N_10416,N_10313,N_10326);
or U10417 (N_10417,N_10273,N_10259);
or U10418 (N_10418,N_10342,N_10266);
nand U10419 (N_10419,N_10267,N_10270);
or U10420 (N_10420,N_10272,N_10256);
nand U10421 (N_10421,N_10323,N_10306);
nor U10422 (N_10422,N_10347,N_10352);
nor U10423 (N_10423,N_10308,N_10285);
and U10424 (N_10424,N_10327,N_10300);
and U10425 (N_10425,N_10325,N_10293);
and U10426 (N_10426,N_10368,N_10315);
nor U10427 (N_10427,N_10311,N_10373);
nand U10428 (N_10428,N_10281,N_10322);
nor U10429 (N_10429,N_10250,N_10312);
or U10430 (N_10430,N_10328,N_10333);
and U10431 (N_10431,N_10263,N_10353);
or U10432 (N_10432,N_10357,N_10340);
nand U10433 (N_10433,N_10369,N_10361);
xor U10434 (N_10434,N_10319,N_10274);
or U10435 (N_10435,N_10292,N_10331);
nand U10436 (N_10436,N_10374,N_10354);
nand U10437 (N_10437,N_10305,N_10341);
xnor U10438 (N_10438,N_10287,N_10282);
nand U10439 (N_10439,N_10264,N_10332);
and U10440 (N_10440,N_10371,N_10342);
or U10441 (N_10441,N_10291,N_10373);
xnor U10442 (N_10442,N_10270,N_10356);
xnor U10443 (N_10443,N_10359,N_10279);
and U10444 (N_10444,N_10340,N_10354);
xnor U10445 (N_10445,N_10339,N_10266);
and U10446 (N_10446,N_10258,N_10268);
or U10447 (N_10447,N_10370,N_10291);
nor U10448 (N_10448,N_10369,N_10288);
and U10449 (N_10449,N_10373,N_10281);
nor U10450 (N_10450,N_10310,N_10345);
xnor U10451 (N_10451,N_10339,N_10306);
xor U10452 (N_10452,N_10282,N_10348);
xnor U10453 (N_10453,N_10332,N_10346);
or U10454 (N_10454,N_10255,N_10260);
nand U10455 (N_10455,N_10357,N_10275);
xor U10456 (N_10456,N_10327,N_10297);
and U10457 (N_10457,N_10310,N_10368);
nand U10458 (N_10458,N_10349,N_10297);
or U10459 (N_10459,N_10299,N_10356);
or U10460 (N_10460,N_10374,N_10272);
and U10461 (N_10461,N_10328,N_10282);
and U10462 (N_10462,N_10271,N_10337);
nor U10463 (N_10463,N_10360,N_10336);
or U10464 (N_10464,N_10273,N_10276);
xor U10465 (N_10465,N_10300,N_10276);
and U10466 (N_10466,N_10353,N_10354);
xor U10467 (N_10467,N_10351,N_10288);
nor U10468 (N_10468,N_10318,N_10272);
xnor U10469 (N_10469,N_10284,N_10291);
nand U10470 (N_10470,N_10252,N_10333);
nor U10471 (N_10471,N_10292,N_10259);
nand U10472 (N_10472,N_10327,N_10320);
or U10473 (N_10473,N_10290,N_10321);
nor U10474 (N_10474,N_10319,N_10345);
nor U10475 (N_10475,N_10266,N_10366);
nor U10476 (N_10476,N_10314,N_10283);
nand U10477 (N_10477,N_10290,N_10313);
xnor U10478 (N_10478,N_10344,N_10329);
or U10479 (N_10479,N_10327,N_10331);
and U10480 (N_10480,N_10318,N_10283);
or U10481 (N_10481,N_10349,N_10257);
nor U10482 (N_10482,N_10272,N_10277);
or U10483 (N_10483,N_10356,N_10269);
and U10484 (N_10484,N_10330,N_10360);
nand U10485 (N_10485,N_10350,N_10253);
xor U10486 (N_10486,N_10323,N_10357);
or U10487 (N_10487,N_10276,N_10286);
and U10488 (N_10488,N_10264,N_10269);
xnor U10489 (N_10489,N_10364,N_10347);
and U10490 (N_10490,N_10306,N_10358);
or U10491 (N_10491,N_10308,N_10263);
or U10492 (N_10492,N_10261,N_10275);
and U10493 (N_10493,N_10293,N_10306);
nand U10494 (N_10494,N_10372,N_10321);
nor U10495 (N_10495,N_10327,N_10257);
and U10496 (N_10496,N_10327,N_10336);
nor U10497 (N_10497,N_10333,N_10363);
nand U10498 (N_10498,N_10278,N_10372);
nand U10499 (N_10499,N_10287,N_10304);
nand U10500 (N_10500,N_10436,N_10488);
or U10501 (N_10501,N_10398,N_10412);
nor U10502 (N_10502,N_10425,N_10413);
xor U10503 (N_10503,N_10460,N_10416);
nand U10504 (N_10504,N_10457,N_10447);
nor U10505 (N_10505,N_10395,N_10442);
and U10506 (N_10506,N_10379,N_10487);
xnor U10507 (N_10507,N_10478,N_10411);
xnor U10508 (N_10508,N_10470,N_10437);
nor U10509 (N_10509,N_10464,N_10491);
and U10510 (N_10510,N_10454,N_10396);
xnor U10511 (N_10511,N_10484,N_10378);
or U10512 (N_10512,N_10439,N_10384);
and U10513 (N_10513,N_10419,N_10463);
or U10514 (N_10514,N_10399,N_10486);
or U10515 (N_10515,N_10446,N_10381);
nor U10516 (N_10516,N_10498,N_10405);
and U10517 (N_10517,N_10462,N_10389);
or U10518 (N_10518,N_10472,N_10474);
and U10519 (N_10519,N_10489,N_10451);
nand U10520 (N_10520,N_10404,N_10387);
nor U10521 (N_10521,N_10476,N_10469);
or U10522 (N_10522,N_10417,N_10438);
and U10523 (N_10523,N_10440,N_10499);
nand U10524 (N_10524,N_10432,N_10377);
xor U10525 (N_10525,N_10456,N_10408);
or U10526 (N_10526,N_10473,N_10435);
and U10527 (N_10527,N_10394,N_10376);
and U10528 (N_10528,N_10492,N_10388);
nor U10529 (N_10529,N_10490,N_10433);
xnor U10530 (N_10530,N_10481,N_10430);
nor U10531 (N_10531,N_10386,N_10449);
or U10532 (N_10532,N_10483,N_10467);
or U10533 (N_10533,N_10482,N_10431);
nor U10534 (N_10534,N_10402,N_10390);
xor U10535 (N_10535,N_10496,N_10448);
or U10536 (N_10536,N_10434,N_10495);
xor U10537 (N_10537,N_10480,N_10424);
nand U10538 (N_10538,N_10423,N_10497);
and U10539 (N_10539,N_10409,N_10380);
nor U10540 (N_10540,N_10494,N_10418);
xnor U10541 (N_10541,N_10392,N_10466);
xnor U10542 (N_10542,N_10385,N_10428);
xor U10543 (N_10543,N_10403,N_10468);
and U10544 (N_10544,N_10427,N_10393);
xor U10545 (N_10545,N_10445,N_10475);
xnor U10546 (N_10546,N_10452,N_10401);
nand U10547 (N_10547,N_10391,N_10450);
or U10548 (N_10548,N_10400,N_10461);
nor U10549 (N_10549,N_10479,N_10383);
xnor U10550 (N_10550,N_10397,N_10455);
or U10551 (N_10551,N_10407,N_10375);
xnor U10552 (N_10552,N_10485,N_10453);
or U10553 (N_10553,N_10465,N_10444);
nor U10554 (N_10554,N_10493,N_10471);
xor U10555 (N_10555,N_10477,N_10441);
xnor U10556 (N_10556,N_10422,N_10459);
nor U10557 (N_10557,N_10421,N_10458);
or U10558 (N_10558,N_10443,N_10429);
and U10559 (N_10559,N_10410,N_10415);
xnor U10560 (N_10560,N_10420,N_10426);
nor U10561 (N_10561,N_10406,N_10382);
nand U10562 (N_10562,N_10414,N_10389);
xor U10563 (N_10563,N_10417,N_10485);
or U10564 (N_10564,N_10487,N_10425);
or U10565 (N_10565,N_10404,N_10402);
or U10566 (N_10566,N_10402,N_10469);
nand U10567 (N_10567,N_10384,N_10443);
or U10568 (N_10568,N_10463,N_10437);
nand U10569 (N_10569,N_10494,N_10430);
nand U10570 (N_10570,N_10418,N_10437);
or U10571 (N_10571,N_10426,N_10459);
nor U10572 (N_10572,N_10379,N_10381);
nor U10573 (N_10573,N_10485,N_10463);
nand U10574 (N_10574,N_10458,N_10415);
nand U10575 (N_10575,N_10405,N_10441);
and U10576 (N_10576,N_10380,N_10451);
nand U10577 (N_10577,N_10379,N_10495);
and U10578 (N_10578,N_10395,N_10469);
nand U10579 (N_10579,N_10495,N_10475);
or U10580 (N_10580,N_10444,N_10458);
nand U10581 (N_10581,N_10466,N_10475);
or U10582 (N_10582,N_10485,N_10474);
and U10583 (N_10583,N_10438,N_10478);
or U10584 (N_10584,N_10438,N_10411);
nor U10585 (N_10585,N_10412,N_10469);
and U10586 (N_10586,N_10464,N_10431);
nor U10587 (N_10587,N_10468,N_10479);
xnor U10588 (N_10588,N_10488,N_10442);
nand U10589 (N_10589,N_10475,N_10446);
nor U10590 (N_10590,N_10409,N_10466);
nor U10591 (N_10591,N_10456,N_10391);
nand U10592 (N_10592,N_10487,N_10491);
and U10593 (N_10593,N_10399,N_10383);
nor U10594 (N_10594,N_10401,N_10433);
or U10595 (N_10595,N_10484,N_10482);
or U10596 (N_10596,N_10440,N_10389);
nor U10597 (N_10597,N_10475,N_10455);
nor U10598 (N_10598,N_10485,N_10473);
nor U10599 (N_10599,N_10426,N_10487);
nor U10600 (N_10600,N_10379,N_10417);
and U10601 (N_10601,N_10409,N_10427);
or U10602 (N_10602,N_10456,N_10381);
nor U10603 (N_10603,N_10459,N_10438);
nand U10604 (N_10604,N_10484,N_10441);
and U10605 (N_10605,N_10485,N_10383);
nand U10606 (N_10606,N_10455,N_10424);
or U10607 (N_10607,N_10398,N_10442);
or U10608 (N_10608,N_10415,N_10417);
or U10609 (N_10609,N_10441,N_10480);
xnor U10610 (N_10610,N_10460,N_10395);
or U10611 (N_10611,N_10446,N_10434);
xor U10612 (N_10612,N_10379,N_10430);
nor U10613 (N_10613,N_10388,N_10480);
or U10614 (N_10614,N_10445,N_10408);
or U10615 (N_10615,N_10396,N_10481);
and U10616 (N_10616,N_10497,N_10494);
and U10617 (N_10617,N_10422,N_10452);
xor U10618 (N_10618,N_10458,N_10481);
and U10619 (N_10619,N_10392,N_10493);
or U10620 (N_10620,N_10432,N_10499);
nor U10621 (N_10621,N_10404,N_10492);
nor U10622 (N_10622,N_10403,N_10448);
xor U10623 (N_10623,N_10385,N_10431);
xnor U10624 (N_10624,N_10453,N_10404);
xor U10625 (N_10625,N_10556,N_10601);
xor U10626 (N_10626,N_10565,N_10557);
and U10627 (N_10627,N_10569,N_10539);
nor U10628 (N_10628,N_10593,N_10617);
and U10629 (N_10629,N_10577,N_10551);
nor U10630 (N_10630,N_10583,N_10506);
xnor U10631 (N_10631,N_10597,N_10530);
nor U10632 (N_10632,N_10526,N_10540);
nor U10633 (N_10633,N_10541,N_10591);
xnor U10634 (N_10634,N_10575,N_10513);
nor U10635 (N_10635,N_10502,N_10618);
nand U10636 (N_10636,N_10598,N_10611);
and U10637 (N_10637,N_10614,N_10579);
xor U10638 (N_10638,N_10596,N_10525);
xnor U10639 (N_10639,N_10501,N_10534);
and U10640 (N_10640,N_10550,N_10582);
nand U10641 (N_10641,N_10615,N_10572);
xor U10642 (N_10642,N_10578,N_10524);
nand U10643 (N_10643,N_10561,N_10573);
and U10644 (N_10644,N_10503,N_10544);
and U10645 (N_10645,N_10620,N_10543);
nand U10646 (N_10646,N_10511,N_10531);
or U10647 (N_10647,N_10545,N_10547);
and U10648 (N_10648,N_10624,N_10554);
or U10649 (N_10649,N_10616,N_10564);
nand U10650 (N_10650,N_10562,N_10535);
or U10651 (N_10651,N_10538,N_10603);
nor U10652 (N_10652,N_10553,N_10527);
or U10653 (N_10653,N_10500,N_10552);
and U10654 (N_10654,N_10505,N_10515);
xnor U10655 (N_10655,N_10520,N_10558);
nand U10656 (N_10656,N_10519,N_10522);
xnor U10657 (N_10657,N_10589,N_10602);
xnor U10658 (N_10658,N_10549,N_10510);
and U10659 (N_10659,N_10518,N_10621);
or U10660 (N_10660,N_10533,N_10507);
xnor U10661 (N_10661,N_10560,N_10588);
nor U10662 (N_10662,N_10570,N_10581);
or U10663 (N_10663,N_10532,N_10607);
xnor U10664 (N_10664,N_10566,N_10609);
and U10665 (N_10665,N_10585,N_10604);
nand U10666 (N_10666,N_10584,N_10563);
and U10667 (N_10667,N_10504,N_10542);
nand U10668 (N_10668,N_10623,N_10600);
nor U10669 (N_10669,N_10592,N_10610);
nand U10670 (N_10670,N_10605,N_10568);
or U10671 (N_10671,N_10508,N_10521);
or U10672 (N_10672,N_10613,N_10509);
nor U10673 (N_10673,N_10576,N_10619);
or U10674 (N_10674,N_10523,N_10595);
or U10675 (N_10675,N_10516,N_10528);
or U10676 (N_10676,N_10512,N_10517);
or U10677 (N_10677,N_10612,N_10580);
xnor U10678 (N_10678,N_10546,N_10537);
and U10679 (N_10679,N_10574,N_10514);
nor U10680 (N_10680,N_10622,N_10529);
nor U10681 (N_10681,N_10586,N_10548);
nor U10682 (N_10682,N_10599,N_10587);
or U10683 (N_10683,N_10555,N_10590);
xnor U10684 (N_10684,N_10608,N_10567);
or U10685 (N_10685,N_10606,N_10571);
xor U10686 (N_10686,N_10594,N_10536);
nand U10687 (N_10687,N_10559,N_10519);
and U10688 (N_10688,N_10549,N_10618);
nand U10689 (N_10689,N_10583,N_10511);
or U10690 (N_10690,N_10534,N_10590);
xnor U10691 (N_10691,N_10617,N_10586);
or U10692 (N_10692,N_10607,N_10573);
nor U10693 (N_10693,N_10546,N_10598);
xnor U10694 (N_10694,N_10579,N_10567);
nand U10695 (N_10695,N_10595,N_10556);
nor U10696 (N_10696,N_10601,N_10530);
xnor U10697 (N_10697,N_10624,N_10572);
nor U10698 (N_10698,N_10586,N_10505);
nand U10699 (N_10699,N_10538,N_10520);
xnor U10700 (N_10700,N_10528,N_10538);
xor U10701 (N_10701,N_10520,N_10616);
nand U10702 (N_10702,N_10609,N_10544);
nand U10703 (N_10703,N_10590,N_10533);
nand U10704 (N_10704,N_10550,N_10518);
nand U10705 (N_10705,N_10599,N_10543);
xor U10706 (N_10706,N_10588,N_10601);
and U10707 (N_10707,N_10501,N_10509);
nand U10708 (N_10708,N_10503,N_10583);
nand U10709 (N_10709,N_10570,N_10599);
nor U10710 (N_10710,N_10599,N_10579);
or U10711 (N_10711,N_10574,N_10581);
or U10712 (N_10712,N_10518,N_10570);
or U10713 (N_10713,N_10610,N_10620);
nor U10714 (N_10714,N_10500,N_10620);
nand U10715 (N_10715,N_10618,N_10534);
nand U10716 (N_10716,N_10588,N_10600);
xnor U10717 (N_10717,N_10544,N_10584);
and U10718 (N_10718,N_10591,N_10593);
and U10719 (N_10719,N_10566,N_10591);
nor U10720 (N_10720,N_10597,N_10601);
or U10721 (N_10721,N_10508,N_10563);
nand U10722 (N_10722,N_10526,N_10589);
xor U10723 (N_10723,N_10620,N_10518);
or U10724 (N_10724,N_10591,N_10592);
and U10725 (N_10725,N_10567,N_10535);
xnor U10726 (N_10726,N_10511,N_10580);
or U10727 (N_10727,N_10586,N_10603);
nor U10728 (N_10728,N_10549,N_10538);
nor U10729 (N_10729,N_10513,N_10564);
and U10730 (N_10730,N_10501,N_10560);
or U10731 (N_10731,N_10550,N_10505);
and U10732 (N_10732,N_10617,N_10530);
nor U10733 (N_10733,N_10579,N_10541);
and U10734 (N_10734,N_10522,N_10622);
and U10735 (N_10735,N_10547,N_10615);
and U10736 (N_10736,N_10537,N_10553);
xnor U10737 (N_10737,N_10587,N_10557);
xnor U10738 (N_10738,N_10526,N_10584);
and U10739 (N_10739,N_10574,N_10618);
nor U10740 (N_10740,N_10555,N_10610);
xor U10741 (N_10741,N_10520,N_10553);
nor U10742 (N_10742,N_10594,N_10584);
nand U10743 (N_10743,N_10501,N_10510);
nand U10744 (N_10744,N_10540,N_10546);
nand U10745 (N_10745,N_10517,N_10581);
nand U10746 (N_10746,N_10568,N_10517);
xnor U10747 (N_10747,N_10568,N_10513);
and U10748 (N_10748,N_10555,N_10611);
nand U10749 (N_10749,N_10584,N_10608);
nand U10750 (N_10750,N_10699,N_10717);
or U10751 (N_10751,N_10724,N_10642);
xnor U10752 (N_10752,N_10627,N_10628);
nor U10753 (N_10753,N_10708,N_10701);
nand U10754 (N_10754,N_10677,N_10661);
and U10755 (N_10755,N_10695,N_10691);
xor U10756 (N_10756,N_10680,N_10703);
or U10757 (N_10757,N_10650,N_10637);
xor U10758 (N_10758,N_10736,N_10660);
nand U10759 (N_10759,N_10714,N_10726);
and U10760 (N_10760,N_10686,N_10641);
xnor U10761 (N_10761,N_10681,N_10716);
nand U10762 (N_10762,N_10630,N_10697);
and U10763 (N_10763,N_10672,N_10662);
nand U10764 (N_10764,N_10734,N_10636);
or U10765 (N_10765,N_10656,N_10725);
or U10766 (N_10766,N_10711,N_10676);
and U10767 (N_10767,N_10705,N_10635);
nand U10768 (N_10768,N_10668,N_10658);
xor U10769 (N_10769,N_10744,N_10729);
or U10770 (N_10770,N_10745,N_10679);
or U10771 (N_10771,N_10692,N_10738);
or U10772 (N_10772,N_10663,N_10626);
or U10773 (N_10773,N_10706,N_10733);
xnor U10774 (N_10774,N_10739,N_10749);
and U10775 (N_10775,N_10712,N_10657);
and U10776 (N_10776,N_10727,N_10640);
nand U10777 (N_10777,N_10685,N_10673);
and U10778 (N_10778,N_10732,N_10666);
and U10779 (N_10779,N_10633,N_10690);
xnor U10780 (N_10780,N_10747,N_10655);
nand U10781 (N_10781,N_10647,N_10728);
nor U10782 (N_10782,N_10671,N_10735);
nor U10783 (N_10783,N_10674,N_10629);
and U10784 (N_10784,N_10731,N_10667);
and U10785 (N_10785,N_10722,N_10748);
or U10786 (N_10786,N_10632,N_10664);
nor U10787 (N_10787,N_10652,N_10720);
nor U10788 (N_10788,N_10742,N_10710);
nand U10789 (N_10789,N_10719,N_10688);
nand U10790 (N_10790,N_10723,N_10631);
or U10791 (N_10791,N_10693,N_10665);
nor U10792 (N_10792,N_10645,N_10700);
nand U10793 (N_10793,N_10678,N_10653);
nor U10794 (N_10794,N_10670,N_10687);
xor U10795 (N_10795,N_10737,N_10689);
or U10796 (N_10796,N_10715,N_10709);
nand U10797 (N_10797,N_10718,N_10644);
or U10798 (N_10798,N_10659,N_10654);
and U10799 (N_10799,N_10638,N_10634);
or U10800 (N_10800,N_10643,N_10669);
or U10801 (N_10801,N_10625,N_10698);
nand U10802 (N_10802,N_10743,N_10648);
nor U10803 (N_10803,N_10649,N_10730);
and U10804 (N_10804,N_10702,N_10639);
nor U10805 (N_10805,N_10683,N_10651);
nand U10806 (N_10806,N_10675,N_10721);
and U10807 (N_10807,N_10713,N_10646);
nor U10808 (N_10808,N_10696,N_10704);
or U10809 (N_10809,N_10684,N_10707);
nand U10810 (N_10810,N_10682,N_10694);
or U10811 (N_10811,N_10740,N_10741);
or U10812 (N_10812,N_10746,N_10722);
xnor U10813 (N_10813,N_10680,N_10743);
or U10814 (N_10814,N_10690,N_10740);
nand U10815 (N_10815,N_10633,N_10630);
nand U10816 (N_10816,N_10643,N_10701);
nor U10817 (N_10817,N_10671,N_10650);
and U10818 (N_10818,N_10734,N_10718);
nand U10819 (N_10819,N_10716,N_10704);
nor U10820 (N_10820,N_10649,N_10665);
xnor U10821 (N_10821,N_10685,N_10707);
nor U10822 (N_10822,N_10737,N_10702);
xor U10823 (N_10823,N_10638,N_10708);
nand U10824 (N_10824,N_10672,N_10748);
nor U10825 (N_10825,N_10694,N_10631);
nand U10826 (N_10826,N_10683,N_10674);
or U10827 (N_10827,N_10694,N_10747);
xnor U10828 (N_10828,N_10688,N_10723);
or U10829 (N_10829,N_10746,N_10720);
nor U10830 (N_10830,N_10678,N_10721);
or U10831 (N_10831,N_10625,N_10720);
nor U10832 (N_10832,N_10666,N_10698);
and U10833 (N_10833,N_10664,N_10655);
nor U10834 (N_10834,N_10626,N_10748);
nor U10835 (N_10835,N_10627,N_10688);
xor U10836 (N_10836,N_10708,N_10678);
or U10837 (N_10837,N_10736,N_10711);
nor U10838 (N_10838,N_10709,N_10742);
or U10839 (N_10839,N_10625,N_10714);
and U10840 (N_10840,N_10650,N_10694);
or U10841 (N_10841,N_10640,N_10668);
xor U10842 (N_10842,N_10646,N_10726);
nand U10843 (N_10843,N_10684,N_10742);
nor U10844 (N_10844,N_10719,N_10632);
nand U10845 (N_10845,N_10705,N_10678);
nand U10846 (N_10846,N_10744,N_10687);
xnor U10847 (N_10847,N_10712,N_10653);
nand U10848 (N_10848,N_10726,N_10690);
nand U10849 (N_10849,N_10690,N_10653);
nor U10850 (N_10850,N_10722,N_10733);
nor U10851 (N_10851,N_10732,N_10654);
and U10852 (N_10852,N_10741,N_10642);
and U10853 (N_10853,N_10655,N_10732);
and U10854 (N_10854,N_10643,N_10691);
or U10855 (N_10855,N_10676,N_10633);
xor U10856 (N_10856,N_10639,N_10732);
xor U10857 (N_10857,N_10716,N_10708);
or U10858 (N_10858,N_10652,N_10673);
and U10859 (N_10859,N_10676,N_10657);
nand U10860 (N_10860,N_10650,N_10707);
nand U10861 (N_10861,N_10724,N_10712);
xnor U10862 (N_10862,N_10731,N_10706);
nor U10863 (N_10863,N_10663,N_10725);
and U10864 (N_10864,N_10739,N_10733);
nand U10865 (N_10865,N_10646,N_10650);
and U10866 (N_10866,N_10673,N_10720);
nor U10867 (N_10867,N_10721,N_10726);
xnor U10868 (N_10868,N_10739,N_10640);
and U10869 (N_10869,N_10681,N_10626);
and U10870 (N_10870,N_10679,N_10629);
or U10871 (N_10871,N_10680,N_10723);
xnor U10872 (N_10872,N_10748,N_10741);
xnor U10873 (N_10873,N_10687,N_10648);
or U10874 (N_10874,N_10649,N_10726);
or U10875 (N_10875,N_10836,N_10857);
nor U10876 (N_10876,N_10803,N_10807);
or U10877 (N_10877,N_10793,N_10843);
or U10878 (N_10878,N_10789,N_10778);
and U10879 (N_10879,N_10819,N_10828);
and U10880 (N_10880,N_10791,N_10862);
nor U10881 (N_10881,N_10774,N_10794);
and U10882 (N_10882,N_10814,N_10804);
or U10883 (N_10883,N_10754,N_10813);
or U10884 (N_10884,N_10801,N_10760);
nor U10885 (N_10885,N_10782,N_10765);
and U10886 (N_10886,N_10816,N_10859);
nor U10887 (N_10887,N_10802,N_10792);
or U10888 (N_10888,N_10856,N_10773);
xnor U10889 (N_10889,N_10776,N_10870);
nand U10890 (N_10890,N_10783,N_10799);
nor U10891 (N_10891,N_10757,N_10833);
nor U10892 (N_10892,N_10798,N_10835);
or U10893 (N_10893,N_10840,N_10824);
nor U10894 (N_10894,N_10821,N_10815);
or U10895 (N_10895,N_10787,N_10817);
or U10896 (N_10896,N_10796,N_10855);
xor U10897 (N_10897,N_10753,N_10854);
xnor U10898 (N_10898,N_10800,N_10845);
nor U10899 (N_10899,N_10844,N_10829);
nor U10900 (N_10900,N_10838,N_10756);
and U10901 (N_10901,N_10759,N_10849);
nand U10902 (N_10902,N_10809,N_10818);
or U10903 (N_10903,N_10861,N_10781);
nor U10904 (N_10904,N_10769,N_10755);
and U10905 (N_10905,N_10866,N_10750);
nand U10906 (N_10906,N_10810,N_10806);
nor U10907 (N_10907,N_10871,N_10839);
nor U10908 (N_10908,N_10860,N_10863);
nor U10909 (N_10909,N_10846,N_10762);
and U10910 (N_10910,N_10851,N_10869);
xnor U10911 (N_10911,N_10853,N_10784);
nor U10912 (N_10912,N_10751,N_10758);
and U10913 (N_10913,N_10842,N_10822);
or U10914 (N_10914,N_10823,N_10805);
and U10915 (N_10915,N_10777,N_10858);
or U10916 (N_10916,N_10852,N_10780);
xnor U10917 (N_10917,N_10864,N_10868);
nor U10918 (N_10918,N_10848,N_10761);
nand U10919 (N_10919,N_10785,N_10831);
nor U10920 (N_10920,N_10797,N_10811);
nor U10921 (N_10921,N_10775,N_10768);
nand U10922 (N_10922,N_10837,N_10841);
nor U10923 (N_10923,N_10772,N_10847);
xor U10924 (N_10924,N_10767,N_10752);
nor U10925 (N_10925,N_10779,N_10788);
or U10926 (N_10926,N_10790,N_10865);
or U10927 (N_10927,N_10826,N_10830);
nor U10928 (N_10928,N_10832,N_10850);
xor U10929 (N_10929,N_10771,N_10874);
xnor U10930 (N_10930,N_10872,N_10795);
xnor U10931 (N_10931,N_10770,N_10766);
nor U10932 (N_10932,N_10764,N_10786);
and U10933 (N_10933,N_10834,N_10763);
nand U10934 (N_10934,N_10825,N_10820);
nand U10935 (N_10935,N_10873,N_10808);
nand U10936 (N_10936,N_10812,N_10827);
xnor U10937 (N_10937,N_10867,N_10770);
nor U10938 (N_10938,N_10781,N_10774);
nor U10939 (N_10939,N_10816,N_10785);
xnor U10940 (N_10940,N_10759,N_10850);
nand U10941 (N_10941,N_10834,N_10777);
nand U10942 (N_10942,N_10776,N_10752);
and U10943 (N_10943,N_10873,N_10766);
xor U10944 (N_10944,N_10760,N_10831);
or U10945 (N_10945,N_10778,N_10777);
and U10946 (N_10946,N_10784,N_10814);
nand U10947 (N_10947,N_10767,N_10783);
nand U10948 (N_10948,N_10809,N_10813);
xnor U10949 (N_10949,N_10823,N_10752);
nor U10950 (N_10950,N_10789,N_10781);
xor U10951 (N_10951,N_10848,N_10809);
nor U10952 (N_10952,N_10854,N_10797);
or U10953 (N_10953,N_10800,N_10831);
and U10954 (N_10954,N_10873,N_10805);
nand U10955 (N_10955,N_10840,N_10772);
nor U10956 (N_10956,N_10805,N_10835);
nand U10957 (N_10957,N_10754,N_10780);
nor U10958 (N_10958,N_10828,N_10791);
or U10959 (N_10959,N_10756,N_10832);
nand U10960 (N_10960,N_10757,N_10856);
and U10961 (N_10961,N_10781,N_10823);
and U10962 (N_10962,N_10825,N_10842);
and U10963 (N_10963,N_10791,N_10838);
nand U10964 (N_10964,N_10834,N_10839);
nor U10965 (N_10965,N_10801,N_10839);
and U10966 (N_10966,N_10834,N_10757);
xor U10967 (N_10967,N_10786,N_10761);
or U10968 (N_10968,N_10856,N_10837);
nor U10969 (N_10969,N_10844,N_10820);
nor U10970 (N_10970,N_10874,N_10750);
nor U10971 (N_10971,N_10822,N_10777);
nor U10972 (N_10972,N_10800,N_10865);
and U10973 (N_10973,N_10821,N_10873);
xnor U10974 (N_10974,N_10754,N_10785);
nor U10975 (N_10975,N_10786,N_10837);
nor U10976 (N_10976,N_10753,N_10860);
nand U10977 (N_10977,N_10806,N_10779);
or U10978 (N_10978,N_10821,N_10759);
and U10979 (N_10979,N_10848,N_10788);
and U10980 (N_10980,N_10778,N_10868);
xor U10981 (N_10981,N_10846,N_10856);
nor U10982 (N_10982,N_10820,N_10780);
nand U10983 (N_10983,N_10852,N_10796);
xor U10984 (N_10984,N_10755,N_10786);
nor U10985 (N_10985,N_10771,N_10801);
nor U10986 (N_10986,N_10856,N_10850);
or U10987 (N_10987,N_10772,N_10766);
nor U10988 (N_10988,N_10822,N_10827);
or U10989 (N_10989,N_10850,N_10871);
and U10990 (N_10990,N_10820,N_10835);
xnor U10991 (N_10991,N_10808,N_10799);
nor U10992 (N_10992,N_10803,N_10845);
or U10993 (N_10993,N_10822,N_10756);
nor U10994 (N_10994,N_10874,N_10763);
or U10995 (N_10995,N_10819,N_10803);
nor U10996 (N_10996,N_10825,N_10828);
and U10997 (N_10997,N_10814,N_10854);
and U10998 (N_10998,N_10756,N_10779);
nor U10999 (N_10999,N_10772,N_10811);
nor U11000 (N_11000,N_10922,N_10952);
xnor U11001 (N_11001,N_10984,N_10911);
and U11002 (N_11002,N_10997,N_10978);
nor U11003 (N_11003,N_10889,N_10973);
nand U11004 (N_11004,N_10919,N_10954);
nor U11005 (N_11005,N_10914,N_10963);
xnor U11006 (N_11006,N_10920,N_10981);
or U11007 (N_11007,N_10902,N_10953);
or U11008 (N_11008,N_10966,N_10888);
and U11009 (N_11009,N_10968,N_10937);
or U11010 (N_11010,N_10908,N_10886);
and U11011 (N_11011,N_10992,N_10928);
nor U11012 (N_11012,N_10875,N_10942);
or U11013 (N_11013,N_10967,N_10974);
and U11014 (N_11014,N_10925,N_10995);
xor U11015 (N_11015,N_10927,N_10989);
nand U11016 (N_11016,N_10941,N_10957);
nor U11017 (N_11017,N_10980,N_10970);
xor U11018 (N_11018,N_10934,N_10881);
or U11019 (N_11019,N_10938,N_10936);
nand U11020 (N_11020,N_10944,N_10926);
nor U11021 (N_11021,N_10985,N_10901);
nor U11022 (N_11022,N_10895,N_10988);
and U11023 (N_11023,N_10918,N_10929);
and U11024 (N_11024,N_10964,N_10962);
and U11025 (N_11025,N_10876,N_10961);
nor U11026 (N_11026,N_10882,N_10894);
xor U11027 (N_11027,N_10982,N_10933);
and U11028 (N_11028,N_10899,N_10924);
or U11029 (N_11029,N_10987,N_10931);
xor U11030 (N_11030,N_10946,N_10892);
nand U11031 (N_11031,N_10935,N_10905);
or U11032 (N_11032,N_10877,N_10948);
nand U11033 (N_11033,N_10959,N_10913);
nor U11034 (N_11034,N_10878,N_10951);
or U11035 (N_11035,N_10972,N_10999);
and U11036 (N_11036,N_10956,N_10916);
nor U11037 (N_11037,N_10904,N_10880);
nand U11038 (N_11038,N_10955,N_10940);
nor U11039 (N_11039,N_10912,N_10943);
nand U11040 (N_11040,N_10896,N_10923);
nor U11041 (N_11041,N_10979,N_10887);
xor U11042 (N_11042,N_10969,N_10893);
xor U11043 (N_11043,N_10879,N_10915);
nor U11044 (N_11044,N_10890,N_10958);
nor U11045 (N_11045,N_10906,N_10990);
or U11046 (N_11046,N_10884,N_10909);
xor U11047 (N_11047,N_10986,N_10947);
xnor U11048 (N_11048,N_10976,N_10917);
and U11049 (N_11049,N_10897,N_10921);
or U11050 (N_11050,N_10945,N_10932);
xor U11051 (N_11051,N_10991,N_10971);
nand U11052 (N_11052,N_10949,N_10903);
nand U11053 (N_11053,N_10977,N_10996);
and U11054 (N_11054,N_10950,N_10998);
nor U11055 (N_11055,N_10930,N_10883);
or U11056 (N_11056,N_10993,N_10960);
or U11057 (N_11057,N_10939,N_10900);
nor U11058 (N_11058,N_10975,N_10965);
xor U11059 (N_11059,N_10983,N_10994);
or U11060 (N_11060,N_10910,N_10891);
and U11061 (N_11061,N_10885,N_10907);
and U11062 (N_11062,N_10898,N_10937);
nand U11063 (N_11063,N_10901,N_10881);
and U11064 (N_11064,N_10886,N_10940);
nand U11065 (N_11065,N_10934,N_10910);
and U11066 (N_11066,N_10966,N_10955);
or U11067 (N_11067,N_10969,N_10967);
or U11068 (N_11068,N_10897,N_10923);
xor U11069 (N_11069,N_10960,N_10908);
nand U11070 (N_11070,N_10954,N_10893);
or U11071 (N_11071,N_10895,N_10930);
xnor U11072 (N_11072,N_10919,N_10964);
and U11073 (N_11073,N_10978,N_10911);
or U11074 (N_11074,N_10989,N_10895);
nor U11075 (N_11075,N_10939,N_10974);
xnor U11076 (N_11076,N_10977,N_10894);
and U11077 (N_11077,N_10959,N_10923);
nor U11078 (N_11078,N_10966,N_10936);
xor U11079 (N_11079,N_10919,N_10913);
xor U11080 (N_11080,N_10991,N_10920);
nand U11081 (N_11081,N_10991,N_10907);
and U11082 (N_11082,N_10913,N_10944);
nand U11083 (N_11083,N_10917,N_10935);
xnor U11084 (N_11084,N_10927,N_10919);
nor U11085 (N_11085,N_10885,N_10949);
nor U11086 (N_11086,N_10967,N_10908);
xnor U11087 (N_11087,N_10930,N_10981);
xnor U11088 (N_11088,N_10899,N_10928);
xor U11089 (N_11089,N_10959,N_10963);
xor U11090 (N_11090,N_10995,N_10882);
nand U11091 (N_11091,N_10943,N_10986);
nand U11092 (N_11092,N_10904,N_10987);
nor U11093 (N_11093,N_10973,N_10961);
nand U11094 (N_11094,N_10928,N_10960);
or U11095 (N_11095,N_10956,N_10955);
nor U11096 (N_11096,N_10899,N_10960);
nand U11097 (N_11097,N_10929,N_10999);
and U11098 (N_11098,N_10896,N_10900);
nand U11099 (N_11099,N_10885,N_10928);
nand U11100 (N_11100,N_10966,N_10900);
and U11101 (N_11101,N_10875,N_10941);
nor U11102 (N_11102,N_10969,N_10877);
and U11103 (N_11103,N_10983,N_10950);
xor U11104 (N_11104,N_10901,N_10910);
and U11105 (N_11105,N_10876,N_10889);
or U11106 (N_11106,N_10893,N_10930);
or U11107 (N_11107,N_10906,N_10967);
xnor U11108 (N_11108,N_10959,N_10928);
nand U11109 (N_11109,N_10899,N_10895);
or U11110 (N_11110,N_10897,N_10885);
or U11111 (N_11111,N_10877,N_10932);
and U11112 (N_11112,N_10879,N_10937);
and U11113 (N_11113,N_10995,N_10881);
nand U11114 (N_11114,N_10951,N_10974);
or U11115 (N_11115,N_10985,N_10953);
and U11116 (N_11116,N_10942,N_10876);
xor U11117 (N_11117,N_10950,N_10935);
nand U11118 (N_11118,N_10931,N_10957);
nand U11119 (N_11119,N_10943,N_10901);
nand U11120 (N_11120,N_10919,N_10936);
nor U11121 (N_11121,N_10962,N_10923);
nor U11122 (N_11122,N_10946,N_10907);
nand U11123 (N_11123,N_10991,N_10890);
and U11124 (N_11124,N_10921,N_10912);
nor U11125 (N_11125,N_11003,N_11118);
xor U11126 (N_11126,N_11106,N_11117);
and U11127 (N_11127,N_11014,N_11087);
or U11128 (N_11128,N_11010,N_11051);
xor U11129 (N_11129,N_11083,N_11045);
nor U11130 (N_11130,N_11078,N_11025);
nand U11131 (N_11131,N_11031,N_11054);
nand U11132 (N_11132,N_11041,N_11017);
nand U11133 (N_11133,N_11084,N_11103);
nand U11134 (N_11134,N_11015,N_11086);
nor U11135 (N_11135,N_11043,N_11047);
or U11136 (N_11136,N_11001,N_11119);
and U11137 (N_11137,N_11077,N_11122);
nor U11138 (N_11138,N_11082,N_11089);
xnor U11139 (N_11139,N_11061,N_11069);
xnor U11140 (N_11140,N_11072,N_11062);
and U11141 (N_11141,N_11006,N_11064);
nand U11142 (N_11142,N_11097,N_11018);
xnor U11143 (N_11143,N_11071,N_11095);
nor U11144 (N_11144,N_11088,N_11034);
and U11145 (N_11145,N_11079,N_11112);
or U11146 (N_11146,N_11081,N_11055);
nand U11147 (N_11147,N_11029,N_11000);
nand U11148 (N_11148,N_11113,N_11105);
or U11149 (N_11149,N_11104,N_11021);
or U11150 (N_11150,N_11060,N_11074);
and U11151 (N_11151,N_11050,N_11035);
and U11152 (N_11152,N_11109,N_11100);
nor U11153 (N_11153,N_11028,N_11065);
and U11154 (N_11154,N_11005,N_11019);
xor U11155 (N_11155,N_11026,N_11066);
xnor U11156 (N_11156,N_11110,N_11108);
nor U11157 (N_11157,N_11053,N_11124);
nor U11158 (N_11158,N_11030,N_11057);
xnor U11159 (N_11159,N_11002,N_11012);
nor U11160 (N_11160,N_11009,N_11052);
nor U11161 (N_11161,N_11091,N_11044);
nor U11162 (N_11162,N_11056,N_11020);
nor U11163 (N_11163,N_11039,N_11076);
xnor U11164 (N_11164,N_11085,N_11036);
and U11165 (N_11165,N_11068,N_11115);
nor U11166 (N_11166,N_11011,N_11033);
nand U11167 (N_11167,N_11067,N_11046);
and U11168 (N_11168,N_11027,N_11023);
or U11169 (N_11169,N_11123,N_11016);
nor U11170 (N_11170,N_11008,N_11096);
or U11171 (N_11171,N_11032,N_11075);
nor U11172 (N_11172,N_11092,N_11120);
nand U11173 (N_11173,N_11059,N_11098);
nand U11174 (N_11174,N_11070,N_11024);
or U11175 (N_11175,N_11114,N_11107);
nor U11176 (N_11176,N_11101,N_11093);
or U11177 (N_11177,N_11094,N_11073);
and U11178 (N_11178,N_11080,N_11048);
xnor U11179 (N_11179,N_11037,N_11090);
or U11180 (N_11180,N_11063,N_11116);
xor U11181 (N_11181,N_11121,N_11099);
xnor U11182 (N_11182,N_11038,N_11042);
xor U11183 (N_11183,N_11007,N_11013);
nand U11184 (N_11184,N_11040,N_11049);
nor U11185 (N_11185,N_11058,N_11111);
or U11186 (N_11186,N_11004,N_11022);
nand U11187 (N_11187,N_11102,N_11111);
and U11188 (N_11188,N_11106,N_11095);
xor U11189 (N_11189,N_11090,N_11112);
or U11190 (N_11190,N_11070,N_11014);
or U11191 (N_11191,N_11030,N_11065);
and U11192 (N_11192,N_11095,N_11122);
nand U11193 (N_11193,N_11017,N_11103);
or U11194 (N_11194,N_11058,N_11088);
xor U11195 (N_11195,N_11035,N_11075);
or U11196 (N_11196,N_11036,N_11038);
or U11197 (N_11197,N_11023,N_11073);
xor U11198 (N_11198,N_11110,N_11104);
or U11199 (N_11199,N_11056,N_11073);
nand U11200 (N_11200,N_11006,N_11076);
xor U11201 (N_11201,N_11009,N_11061);
or U11202 (N_11202,N_11070,N_11049);
nor U11203 (N_11203,N_11057,N_11006);
xor U11204 (N_11204,N_11103,N_11036);
nor U11205 (N_11205,N_11096,N_11077);
nand U11206 (N_11206,N_11081,N_11090);
nor U11207 (N_11207,N_11092,N_11098);
or U11208 (N_11208,N_11086,N_11035);
nor U11209 (N_11209,N_11020,N_11014);
nand U11210 (N_11210,N_11043,N_11031);
xor U11211 (N_11211,N_11020,N_11070);
and U11212 (N_11212,N_11029,N_11050);
xor U11213 (N_11213,N_11000,N_11112);
and U11214 (N_11214,N_11047,N_11110);
nor U11215 (N_11215,N_11013,N_11033);
nor U11216 (N_11216,N_11093,N_11086);
nand U11217 (N_11217,N_11071,N_11102);
and U11218 (N_11218,N_11019,N_11112);
and U11219 (N_11219,N_11085,N_11076);
xnor U11220 (N_11220,N_11015,N_11085);
nor U11221 (N_11221,N_11089,N_11013);
nor U11222 (N_11222,N_11035,N_11016);
xnor U11223 (N_11223,N_11067,N_11065);
xor U11224 (N_11224,N_11118,N_11028);
and U11225 (N_11225,N_11020,N_11001);
and U11226 (N_11226,N_11035,N_11083);
xor U11227 (N_11227,N_11032,N_11065);
xnor U11228 (N_11228,N_11122,N_11121);
and U11229 (N_11229,N_11108,N_11103);
and U11230 (N_11230,N_11113,N_11065);
or U11231 (N_11231,N_11049,N_11116);
nor U11232 (N_11232,N_11033,N_11060);
nor U11233 (N_11233,N_11122,N_11012);
nor U11234 (N_11234,N_11052,N_11097);
and U11235 (N_11235,N_11022,N_11100);
nor U11236 (N_11236,N_11032,N_11084);
nor U11237 (N_11237,N_11085,N_11010);
nor U11238 (N_11238,N_11069,N_11008);
xnor U11239 (N_11239,N_11043,N_11106);
and U11240 (N_11240,N_11109,N_11111);
or U11241 (N_11241,N_11015,N_11102);
nand U11242 (N_11242,N_11037,N_11073);
nor U11243 (N_11243,N_11092,N_11034);
or U11244 (N_11244,N_11038,N_11037);
xor U11245 (N_11245,N_11103,N_11053);
or U11246 (N_11246,N_11042,N_11053);
and U11247 (N_11247,N_11075,N_11008);
and U11248 (N_11248,N_11108,N_11058);
or U11249 (N_11249,N_11095,N_11090);
and U11250 (N_11250,N_11237,N_11136);
or U11251 (N_11251,N_11225,N_11179);
xor U11252 (N_11252,N_11242,N_11191);
nand U11253 (N_11253,N_11217,N_11125);
or U11254 (N_11254,N_11233,N_11226);
and U11255 (N_11255,N_11134,N_11206);
nor U11256 (N_11256,N_11159,N_11224);
and U11257 (N_11257,N_11216,N_11249);
nor U11258 (N_11258,N_11205,N_11239);
xnor U11259 (N_11259,N_11201,N_11197);
nor U11260 (N_11260,N_11174,N_11194);
xor U11261 (N_11261,N_11208,N_11177);
and U11262 (N_11262,N_11240,N_11202);
or U11263 (N_11263,N_11199,N_11246);
nor U11264 (N_11264,N_11223,N_11207);
xnor U11265 (N_11265,N_11243,N_11234);
or U11266 (N_11266,N_11165,N_11198);
and U11267 (N_11267,N_11245,N_11143);
xnor U11268 (N_11268,N_11169,N_11154);
and U11269 (N_11269,N_11204,N_11135);
and U11270 (N_11270,N_11141,N_11166);
or U11271 (N_11271,N_11146,N_11190);
nand U11272 (N_11272,N_11138,N_11130);
or U11273 (N_11273,N_11212,N_11248);
and U11274 (N_11274,N_11144,N_11200);
nand U11275 (N_11275,N_11171,N_11232);
nand U11276 (N_11276,N_11195,N_11210);
nand U11277 (N_11277,N_11151,N_11167);
or U11278 (N_11278,N_11149,N_11222);
and U11279 (N_11279,N_11192,N_11238);
xor U11280 (N_11280,N_11140,N_11181);
xnor U11281 (N_11281,N_11126,N_11187);
nor U11282 (N_11282,N_11153,N_11132);
nand U11283 (N_11283,N_11158,N_11175);
nand U11284 (N_11284,N_11178,N_11230);
nand U11285 (N_11285,N_11186,N_11183);
nand U11286 (N_11286,N_11228,N_11247);
xor U11287 (N_11287,N_11173,N_11127);
or U11288 (N_11288,N_11157,N_11170);
nor U11289 (N_11289,N_11209,N_11231);
nor U11290 (N_11290,N_11160,N_11155);
nand U11291 (N_11291,N_11227,N_11182);
nor U11292 (N_11292,N_11131,N_11211);
nand U11293 (N_11293,N_11163,N_11129);
or U11294 (N_11294,N_11133,N_11203);
xor U11295 (N_11295,N_11172,N_11188);
or U11296 (N_11296,N_11168,N_11142);
nor U11297 (N_11297,N_11215,N_11162);
nand U11298 (N_11298,N_11147,N_11241);
or U11299 (N_11299,N_11176,N_11150);
or U11300 (N_11300,N_11219,N_11220);
or U11301 (N_11301,N_11196,N_11185);
nand U11302 (N_11302,N_11189,N_11244);
and U11303 (N_11303,N_11148,N_11145);
and U11304 (N_11304,N_11218,N_11156);
nand U11305 (N_11305,N_11213,N_11214);
nor U11306 (N_11306,N_11137,N_11236);
nor U11307 (N_11307,N_11139,N_11128);
xnor U11308 (N_11308,N_11184,N_11221);
xnor U11309 (N_11309,N_11161,N_11152);
nand U11310 (N_11310,N_11193,N_11235);
and U11311 (N_11311,N_11180,N_11164);
xnor U11312 (N_11312,N_11229,N_11183);
and U11313 (N_11313,N_11162,N_11182);
or U11314 (N_11314,N_11193,N_11141);
nor U11315 (N_11315,N_11216,N_11233);
nand U11316 (N_11316,N_11226,N_11178);
xnor U11317 (N_11317,N_11126,N_11125);
xnor U11318 (N_11318,N_11181,N_11142);
and U11319 (N_11319,N_11133,N_11216);
nor U11320 (N_11320,N_11223,N_11227);
nor U11321 (N_11321,N_11132,N_11145);
nor U11322 (N_11322,N_11217,N_11225);
xnor U11323 (N_11323,N_11152,N_11248);
xor U11324 (N_11324,N_11211,N_11244);
nor U11325 (N_11325,N_11216,N_11212);
xor U11326 (N_11326,N_11211,N_11177);
nor U11327 (N_11327,N_11236,N_11181);
nand U11328 (N_11328,N_11154,N_11203);
and U11329 (N_11329,N_11223,N_11205);
nand U11330 (N_11330,N_11131,N_11224);
nand U11331 (N_11331,N_11207,N_11211);
xnor U11332 (N_11332,N_11137,N_11218);
xnor U11333 (N_11333,N_11169,N_11160);
xor U11334 (N_11334,N_11238,N_11207);
and U11335 (N_11335,N_11184,N_11180);
and U11336 (N_11336,N_11237,N_11248);
or U11337 (N_11337,N_11127,N_11176);
or U11338 (N_11338,N_11142,N_11192);
xor U11339 (N_11339,N_11159,N_11192);
and U11340 (N_11340,N_11190,N_11205);
or U11341 (N_11341,N_11191,N_11245);
nor U11342 (N_11342,N_11201,N_11193);
and U11343 (N_11343,N_11202,N_11208);
and U11344 (N_11344,N_11133,N_11248);
or U11345 (N_11345,N_11174,N_11198);
or U11346 (N_11346,N_11139,N_11236);
xor U11347 (N_11347,N_11230,N_11204);
and U11348 (N_11348,N_11210,N_11221);
xor U11349 (N_11349,N_11194,N_11223);
or U11350 (N_11350,N_11200,N_11173);
xor U11351 (N_11351,N_11168,N_11149);
nand U11352 (N_11352,N_11143,N_11125);
nor U11353 (N_11353,N_11165,N_11206);
or U11354 (N_11354,N_11140,N_11233);
or U11355 (N_11355,N_11170,N_11237);
xnor U11356 (N_11356,N_11136,N_11223);
nand U11357 (N_11357,N_11172,N_11178);
xnor U11358 (N_11358,N_11174,N_11157);
xor U11359 (N_11359,N_11249,N_11224);
or U11360 (N_11360,N_11165,N_11180);
nand U11361 (N_11361,N_11215,N_11187);
and U11362 (N_11362,N_11160,N_11214);
or U11363 (N_11363,N_11149,N_11196);
and U11364 (N_11364,N_11132,N_11166);
xor U11365 (N_11365,N_11212,N_11217);
nor U11366 (N_11366,N_11233,N_11137);
nor U11367 (N_11367,N_11212,N_11148);
and U11368 (N_11368,N_11176,N_11173);
and U11369 (N_11369,N_11222,N_11153);
or U11370 (N_11370,N_11207,N_11133);
and U11371 (N_11371,N_11137,N_11232);
xnor U11372 (N_11372,N_11248,N_11150);
nand U11373 (N_11373,N_11129,N_11151);
and U11374 (N_11374,N_11233,N_11144);
and U11375 (N_11375,N_11339,N_11315);
nand U11376 (N_11376,N_11306,N_11278);
nand U11377 (N_11377,N_11302,N_11312);
nand U11378 (N_11378,N_11256,N_11348);
nand U11379 (N_11379,N_11360,N_11307);
nor U11380 (N_11380,N_11314,N_11296);
nor U11381 (N_11381,N_11265,N_11253);
xnor U11382 (N_11382,N_11250,N_11344);
nand U11383 (N_11383,N_11317,N_11354);
nor U11384 (N_11384,N_11311,N_11345);
and U11385 (N_11385,N_11292,N_11293);
and U11386 (N_11386,N_11341,N_11266);
and U11387 (N_11387,N_11300,N_11269);
xnor U11388 (N_11388,N_11324,N_11329);
or U11389 (N_11389,N_11335,N_11251);
nand U11390 (N_11390,N_11349,N_11343);
xor U11391 (N_11391,N_11267,N_11257);
nor U11392 (N_11392,N_11361,N_11350);
or U11393 (N_11393,N_11330,N_11325);
nand U11394 (N_11394,N_11298,N_11274);
xnor U11395 (N_11395,N_11337,N_11346);
nand U11396 (N_11396,N_11322,N_11270);
or U11397 (N_11397,N_11364,N_11370);
or U11398 (N_11398,N_11333,N_11371);
nor U11399 (N_11399,N_11310,N_11366);
nor U11400 (N_11400,N_11286,N_11297);
and U11401 (N_11401,N_11332,N_11359);
nor U11402 (N_11402,N_11363,N_11342);
xor U11403 (N_11403,N_11355,N_11316);
nor U11404 (N_11404,N_11323,N_11368);
or U11405 (N_11405,N_11261,N_11291);
nor U11406 (N_11406,N_11352,N_11294);
or U11407 (N_11407,N_11275,N_11367);
or U11408 (N_11408,N_11336,N_11334);
nand U11409 (N_11409,N_11271,N_11281);
nand U11410 (N_11410,N_11268,N_11347);
nor U11411 (N_11411,N_11258,N_11303);
and U11412 (N_11412,N_11340,N_11319);
nor U11413 (N_11413,N_11299,N_11369);
or U11414 (N_11414,N_11357,N_11260);
xor U11415 (N_11415,N_11264,N_11255);
xnor U11416 (N_11416,N_11326,N_11313);
or U11417 (N_11417,N_11280,N_11290);
and U11418 (N_11418,N_11277,N_11338);
nand U11419 (N_11419,N_11356,N_11263);
or U11420 (N_11420,N_11321,N_11305);
and U11421 (N_11421,N_11373,N_11331);
nor U11422 (N_11422,N_11276,N_11295);
nand U11423 (N_11423,N_11259,N_11358);
xor U11424 (N_11424,N_11372,N_11328);
and U11425 (N_11425,N_11318,N_11289);
nand U11426 (N_11426,N_11284,N_11252);
or U11427 (N_11427,N_11309,N_11351);
nand U11428 (N_11428,N_11285,N_11362);
nand U11429 (N_11429,N_11262,N_11308);
or U11430 (N_11430,N_11279,N_11301);
nand U11431 (N_11431,N_11374,N_11353);
xnor U11432 (N_11432,N_11273,N_11304);
nand U11433 (N_11433,N_11254,N_11272);
and U11434 (N_11434,N_11282,N_11320);
and U11435 (N_11435,N_11287,N_11288);
nor U11436 (N_11436,N_11327,N_11283);
nand U11437 (N_11437,N_11365,N_11361);
and U11438 (N_11438,N_11313,N_11276);
xnor U11439 (N_11439,N_11318,N_11338);
nand U11440 (N_11440,N_11264,N_11298);
or U11441 (N_11441,N_11352,N_11251);
xnor U11442 (N_11442,N_11274,N_11318);
xor U11443 (N_11443,N_11369,N_11300);
and U11444 (N_11444,N_11316,N_11364);
and U11445 (N_11445,N_11314,N_11276);
nand U11446 (N_11446,N_11310,N_11351);
or U11447 (N_11447,N_11355,N_11368);
nor U11448 (N_11448,N_11257,N_11322);
or U11449 (N_11449,N_11276,N_11329);
nor U11450 (N_11450,N_11294,N_11260);
nand U11451 (N_11451,N_11333,N_11355);
or U11452 (N_11452,N_11333,N_11269);
xor U11453 (N_11453,N_11324,N_11319);
and U11454 (N_11454,N_11254,N_11311);
nor U11455 (N_11455,N_11288,N_11313);
nand U11456 (N_11456,N_11289,N_11294);
xor U11457 (N_11457,N_11305,N_11277);
xor U11458 (N_11458,N_11254,N_11342);
nand U11459 (N_11459,N_11274,N_11342);
xor U11460 (N_11460,N_11279,N_11256);
or U11461 (N_11461,N_11289,N_11295);
or U11462 (N_11462,N_11340,N_11333);
or U11463 (N_11463,N_11312,N_11318);
xnor U11464 (N_11464,N_11315,N_11360);
xnor U11465 (N_11465,N_11277,N_11359);
or U11466 (N_11466,N_11264,N_11365);
or U11467 (N_11467,N_11373,N_11281);
xnor U11468 (N_11468,N_11256,N_11301);
nand U11469 (N_11469,N_11340,N_11250);
and U11470 (N_11470,N_11315,N_11350);
nand U11471 (N_11471,N_11316,N_11341);
xor U11472 (N_11472,N_11291,N_11332);
or U11473 (N_11473,N_11355,N_11258);
nor U11474 (N_11474,N_11281,N_11313);
nand U11475 (N_11475,N_11269,N_11311);
xnor U11476 (N_11476,N_11328,N_11351);
nand U11477 (N_11477,N_11366,N_11343);
or U11478 (N_11478,N_11366,N_11338);
xor U11479 (N_11479,N_11349,N_11260);
and U11480 (N_11480,N_11368,N_11335);
and U11481 (N_11481,N_11332,N_11317);
and U11482 (N_11482,N_11255,N_11296);
xnor U11483 (N_11483,N_11347,N_11266);
nor U11484 (N_11484,N_11374,N_11275);
and U11485 (N_11485,N_11369,N_11277);
xor U11486 (N_11486,N_11276,N_11335);
and U11487 (N_11487,N_11362,N_11289);
nand U11488 (N_11488,N_11305,N_11292);
nand U11489 (N_11489,N_11278,N_11335);
nor U11490 (N_11490,N_11337,N_11256);
and U11491 (N_11491,N_11365,N_11349);
and U11492 (N_11492,N_11254,N_11303);
nand U11493 (N_11493,N_11337,N_11269);
nor U11494 (N_11494,N_11262,N_11313);
and U11495 (N_11495,N_11255,N_11363);
nand U11496 (N_11496,N_11357,N_11331);
and U11497 (N_11497,N_11342,N_11273);
and U11498 (N_11498,N_11274,N_11253);
or U11499 (N_11499,N_11266,N_11290);
xnor U11500 (N_11500,N_11410,N_11396);
and U11501 (N_11501,N_11399,N_11402);
or U11502 (N_11502,N_11401,N_11450);
nand U11503 (N_11503,N_11407,N_11383);
nand U11504 (N_11504,N_11420,N_11385);
xor U11505 (N_11505,N_11446,N_11429);
xor U11506 (N_11506,N_11496,N_11418);
nor U11507 (N_11507,N_11438,N_11481);
xor U11508 (N_11508,N_11379,N_11455);
nor U11509 (N_11509,N_11463,N_11492);
and U11510 (N_11510,N_11472,N_11457);
nand U11511 (N_11511,N_11482,N_11431);
xnor U11512 (N_11512,N_11378,N_11416);
or U11513 (N_11513,N_11494,N_11493);
nand U11514 (N_11514,N_11439,N_11488);
nand U11515 (N_11515,N_11409,N_11419);
or U11516 (N_11516,N_11468,N_11461);
nand U11517 (N_11517,N_11456,N_11445);
and U11518 (N_11518,N_11454,N_11473);
nor U11519 (N_11519,N_11467,N_11380);
and U11520 (N_11520,N_11483,N_11478);
or U11521 (N_11521,N_11394,N_11412);
nor U11522 (N_11522,N_11442,N_11400);
nor U11523 (N_11523,N_11423,N_11435);
nand U11524 (N_11524,N_11425,N_11477);
and U11525 (N_11525,N_11484,N_11405);
xnor U11526 (N_11526,N_11444,N_11465);
and U11527 (N_11527,N_11430,N_11479);
nand U11528 (N_11528,N_11411,N_11397);
nor U11529 (N_11529,N_11475,N_11464);
xnor U11530 (N_11530,N_11462,N_11436);
xor U11531 (N_11531,N_11387,N_11422);
nor U11532 (N_11532,N_11485,N_11375);
or U11533 (N_11533,N_11443,N_11469);
nand U11534 (N_11534,N_11389,N_11459);
nand U11535 (N_11535,N_11393,N_11386);
xor U11536 (N_11536,N_11424,N_11384);
xor U11537 (N_11537,N_11381,N_11452);
nor U11538 (N_11538,N_11470,N_11406);
nand U11539 (N_11539,N_11433,N_11447);
xnor U11540 (N_11540,N_11487,N_11392);
nand U11541 (N_11541,N_11499,N_11458);
nor U11542 (N_11542,N_11421,N_11474);
or U11543 (N_11543,N_11497,N_11414);
xnor U11544 (N_11544,N_11434,N_11398);
nand U11545 (N_11545,N_11460,N_11377);
nor U11546 (N_11546,N_11440,N_11426);
or U11547 (N_11547,N_11491,N_11437);
or U11548 (N_11548,N_11415,N_11376);
nor U11549 (N_11549,N_11476,N_11441);
or U11550 (N_11550,N_11489,N_11404);
and U11551 (N_11551,N_11449,N_11480);
nor U11552 (N_11552,N_11417,N_11495);
and U11553 (N_11553,N_11408,N_11486);
nand U11554 (N_11554,N_11428,N_11453);
and U11555 (N_11555,N_11382,N_11498);
or U11556 (N_11556,N_11413,N_11432);
nor U11557 (N_11557,N_11448,N_11466);
or U11558 (N_11558,N_11490,N_11451);
nand U11559 (N_11559,N_11427,N_11471);
xnor U11560 (N_11560,N_11395,N_11403);
xor U11561 (N_11561,N_11390,N_11388);
xnor U11562 (N_11562,N_11391,N_11397);
and U11563 (N_11563,N_11387,N_11482);
nor U11564 (N_11564,N_11406,N_11491);
nand U11565 (N_11565,N_11418,N_11467);
nand U11566 (N_11566,N_11442,N_11427);
and U11567 (N_11567,N_11495,N_11471);
nand U11568 (N_11568,N_11457,N_11425);
nand U11569 (N_11569,N_11403,N_11454);
and U11570 (N_11570,N_11461,N_11436);
and U11571 (N_11571,N_11417,N_11484);
and U11572 (N_11572,N_11383,N_11483);
nor U11573 (N_11573,N_11460,N_11418);
and U11574 (N_11574,N_11442,N_11406);
nand U11575 (N_11575,N_11409,N_11399);
xnor U11576 (N_11576,N_11494,N_11484);
and U11577 (N_11577,N_11473,N_11397);
and U11578 (N_11578,N_11449,N_11476);
nand U11579 (N_11579,N_11396,N_11453);
nand U11580 (N_11580,N_11497,N_11464);
nand U11581 (N_11581,N_11426,N_11421);
nand U11582 (N_11582,N_11412,N_11484);
nand U11583 (N_11583,N_11472,N_11456);
nor U11584 (N_11584,N_11482,N_11443);
or U11585 (N_11585,N_11478,N_11375);
or U11586 (N_11586,N_11462,N_11379);
or U11587 (N_11587,N_11431,N_11401);
nand U11588 (N_11588,N_11423,N_11416);
and U11589 (N_11589,N_11400,N_11452);
or U11590 (N_11590,N_11442,N_11468);
xor U11591 (N_11591,N_11398,N_11427);
xnor U11592 (N_11592,N_11401,N_11416);
or U11593 (N_11593,N_11383,N_11393);
or U11594 (N_11594,N_11479,N_11462);
nor U11595 (N_11595,N_11391,N_11496);
nand U11596 (N_11596,N_11493,N_11473);
or U11597 (N_11597,N_11454,N_11375);
nor U11598 (N_11598,N_11488,N_11404);
xnor U11599 (N_11599,N_11466,N_11493);
or U11600 (N_11600,N_11400,N_11428);
xnor U11601 (N_11601,N_11409,N_11468);
xnor U11602 (N_11602,N_11459,N_11478);
and U11603 (N_11603,N_11469,N_11477);
or U11604 (N_11604,N_11397,N_11487);
xnor U11605 (N_11605,N_11381,N_11427);
nor U11606 (N_11606,N_11484,N_11438);
or U11607 (N_11607,N_11392,N_11385);
nand U11608 (N_11608,N_11393,N_11472);
nor U11609 (N_11609,N_11484,N_11451);
or U11610 (N_11610,N_11411,N_11467);
and U11611 (N_11611,N_11461,N_11431);
or U11612 (N_11612,N_11461,N_11406);
or U11613 (N_11613,N_11385,N_11400);
nor U11614 (N_11614,N_11412,N_11495);
xnor U11615 (N_11615,N_11428,N_11435);
and U11616 (N_11616,N_11399,N_11458);
xor U11617 (N_11617,N_11417,N_11446);
or U11618 (N_11618,N_11456,N_11418);
or U11619 (N_11619,N_11471,N_11451);
or U11620 (N_11620,N_11378,N_11447);
or U11621 (N_11621,N_11441,N_11395);
or U11622 (N_11622,N_11425,N_11471);
xor U11623 (N_11623,N_11390,N_11405);
xor U11624 (N_11624,N_11442,N_11404);
or U11625 (N_11625,N_11545,N_11513);
and U11626 (N_11626,N_11624,N_11510);
and U11627 (N_11627,N_11581,N_11597);
nand U11628 (N_11628,N_11580,N_11544);
xnor U11629 (N_11629,N_11570,N_11563);
xnor U11630 (N_11630,N_11520,N_11515);
nand U11631 (N_11631,N_11532,N_11548);
nand U11632 (N_11632,N_11576,N_11584);
nor U11633 (N_11633,N_11621,N_11539);
or U11634 (N_11634,N_11534,N_11573);
or U11635 (N_11635,N_11587,N_11586);
and U11636 (N_11636,N_11519,N_11610);
xnor U11637 (N_11637,N_11528,N_11589);
nor U11638 (N_11638,N_11522,N_11620);
xor U11639 (N_11639,N_11507,N_11619);
nand U11640 (N_11640,N_11523,N_11529);
nor U11641 (N_11641,N_11617,N_11598);
and U11642 (N_11642,N_11551,N_11601);
or U11643 (N_11643,N_11611,N_11595);
and U11644 (N_11644,N_11574,N_11540);
nand U11645 (N_11645,N_11547,N_11527);
xnor U11646 (N_11646,N_11613,N_11509);
xor U11647 (N_11647,N_11511,N_11596);
and U11648 (N_11648,N_11530,N_11622);
nand U11649 (N_11649,N_11546,N_11550);
nand U11650 (N_11650,N_11556,N_11555);
nand U11651 (N_11651,N_11602,N_11594);
or U11652 (N_11652,N_11582,N_11514);
or U11653 (N_11653,N_11525,N_11506);
xnor U11654 (N_11654,N_11500,N_11502);
nor U11655 (N_11655,N_11590,N_11614);
nor U11656 (N_11656,N_11568,N_11554);
xnor U11657 (N_11657,N_11577,N_11549);
or U11658 (N_11658,N_11615,N_11538);
xor U11659 (N_11659,N_11557,N_11560);
or U11660 (N_11660,N_11536,N_11605);
xor U11661 (N_11661,N_11541,N_11564);
and U11662 (N_11662,N_11535,N_11608);
and U11663 (N_11663,N_11518,N_11592);
or U11664 (N_11664,N_11609,N_11585);
and U11665 (N_11665,N_11607,N_11512);
nor U11666 (N_11666,N_11575,N_11504);
or U11667 (N_11667,N_11583,N_11591);
or U11668 (N_11668,N_11524,N_11526);
nor U11669 (N_11669,N_11618,N_11508);
nand U11670 (N_11670,N_11565,N_11566);
nand U11671 (N_11671,N_11537,N_11558);
and U11672 (N_11672,N_11578,N_11505);
or U11673 (N_11673,N_11603,N_11579);
xnor U11674 (N_11674,N_11521,N_11559);
nor U11675 (N_11675,N_11553,N_11562);
xnor U11676 (N_11676,N_11503,N_11571);
nor U11677 (N_11677,N_11516,N_11606);
nand U11678 (N_11678,N_11612,N_11588);
or U11679 (N_11679,N_11604,N_11593);
or U11680 (N_11680,N_11542,N_11533);
xor U11681 (N_11681,N_11572,N_11616);
nor U11682 (N_11682,N_11561,N_11623);
and U11683 (N_11683,N_11501,N_11552);
xnor U11684 (N_11684,N_11531,N_11600);
nor U11685 (N_11685,N_11517,N_11569);
xnor U11686 (N_11686,N_11599,N_11567);
xor U11687 (N_11687,N_11543,N_11597);
and U11688 (N_11688,N_11593,N_11554);
xnor U11689 (N_11689,N_11594,N_11533);
nand U11690 (N_11690,N_11521,N_11564);
or U11691 (N_11691,N_11609,N_11580);
xor U11692 (N_11692,N_11562,N_11595);
nand U11693 (N_11693,N_11561,N_11572);
or U11694 (N_11694,N_11592,N_11622);
or U11695 (N_11695,N_11553,N_11598);
nand U11696 (N_11696,N_11582,N_11545);
and U11697 (N_11697,N_11520,N_11576);
or U11698 (N_11698,N_11503,N_11506);
or U11699 (N_11699,N_11600,N_11512);
nor U11700 (N_11700,N_11583,N_11534);
xnor U11701 (N_11701,N_11551,N_11521);
and U11702 (N_11702,N_11524,N_11544);
nand U11703 (N_11703,N_11548,N_11513);
xnor U11704 (N_11704,N_11527,N_11507);
xnor U11705 (N_11705,N_11601,N_11527);
or U11706 (N_11706,N_11562,N_11563);
and U11707 (N_11707,N_11588,N_11559);
or U11708 (N_11708,N_11538,N_11521);
nand U11709 (N_11709,N_11506,N_11554);
and U11710 (N_11710,N_11612,N_11564);
and U11711 (N_11711,N_11528,N_11523);
and U11712 (N_11712,N_11551,N_11560);
nand U11713 (N_11713,N_11544,N_11534);
and U11714 (N_11714,N_11505,N_11621);
nor U11715 (N_11715,N_11571,N_11560);
and U11716 (N_11716,N_11508,N_11519);
and U11717 (N_11717,N_11613,N_11545);
xnor U11718 (N_11718,N_11553,N_11617);
nor U11719 (N_11719,N_11615,N_11590);
xor U11720 (N_11720,N_11594,N_11541);
and U11721 (N_11721,N_11595,N_11621);
and U11722 (N_11722,N_11502,N_11578);
and U11723 (N_11723,N_11545,N_11615);
nand U11724 (N_11724,N_11606,N_11523);
and U11725 (N_11725,N_11561,N_11552);
nand U11726 (N_11726,N_11577,N_11528);
nor U11727 (N_11727,N_11588,N_11561);
xnor U11728 (N_11728,N_11578,N_11527);
nor U11729 (N_11729,N_11547,N_11569);
nand U11730 (N_11730,N_11602,N_11560);
nand U11731 (N_11731,N_11560,N_11620);
nand U11732 (N_11732,N_11527,N_11598);
nor U11733 (N_11733,N_11618,N_11592);
xor U11734 (N_11734,N_11616,N_11533);
xor U11735 (N_11735,N_11534,N_11509);
nand U11736 (N_11736,N_11566,N_11545);
nor U11737 (N_11737,N_11617,N_11508);
and U11738 (N_11738,N_11526,N_11528);
or U11739 (N_11739,N_11609,N_11539);
or U11740 (N_11740,N_11530,N_11571);
or U11741 (N_11741,N_11518,N_11539);
and U11742 (N_11742,N_11540,N_11603);
or U11743 (N_11743,N_11558,N_11514);
nand U11744 (N_11744,N_11611,N_11525);
xor U11745 (N_11745,N_11531,N_11579);
xor U11746 (N_11746,N_11528,N_11606);
and U11747 (N_11747,N_11538,N_11509);
and U11748 (N_11748,N_11537,N_11585);
nor U11749 (N_11749,N_11615,N_11570);
nand U11750 (N_11750,N_11703,N_11741);
and U11751 (N_11751,N_11700,N_11677);
nand U11752 (N_11752,N_11654,N_11744);
nand U11753 (N_11753,N_11743,N_11647);
or U11754 (N_11754,N_11712,N_11684);
or U11755 (N_11755,N_11749,N_11731);
and U11756 (N_11756,N_11704,N_11717);
or U11757 (N_11757,N_11739,N_11695);
xor U11758 (N_11758,N_11676,N_11683);
and U11759 (N_11759,N_11646,N_11691);
or U11760 (N_11760,N_11655,N_11656);
nor U11761 (N_11761,N_11726,N_11682);
nand U11762 (N_11762,N_11679,N_11665);
and U11763 (N_11763,N_11742,N_11658);
nand U11764 (N_11764,N_11663,N_11625);
nand U11765 (N_11765,N_11667,N_11713);
nor U11766 (N_11766,N_11687,N_11664);
nor U11767 (N_11767,N_11748,N_11697);
xor U11768 (N_11768,N_11738,N_11633);
or U11769 (N_11769,N_11634,N_11629);
nor U11770 (N_11770,N_11626,N_11668);
nor U11771 (N_11771,N_11644,N_11734);
or U11772 (N_11772,N_11724,N_11688);
xnor U11773 (N_11773,N_11685,N_11696);
xnor U11774 (N_11774,N_11694,N_11672);
and U11775 (N_11775,N_11740,N_11701);
or U11776 (N_11776,N_11640,N_11678);
nand U11777 (N_11777,N_11666,N_11635);
xnor U11778 (N_11778,N_11718,N_11639);
xnor U11779 (N_11779,N_11730,N_11659);
nor U11780 (N_11780,N_11661,N_11652);
and U11781 (N_11781,N_11746,N_11637);
and U11782 (N_11782,N_11627,N_11725);
or U11783 (N_11783,N_11680,N_11693);
nor U11784 (N_11784,N_11715,N_11708);
nand U11785 (N_11785,N_11648,N_11705);
xnor U11786 (N_11786,N_11643,N_11711);
nor U11787 (N_11787,N_11669,N_11657);
nor U11788 (N_11788,N_11706,N_11729);
xnor U11789 (N_11789,N_11745,N_11707);
xnor U11790 (N_11790,N_11714,N_11660);
nor U11791 (N_11791,N_11689,N_11735);
or U11792 (N_11792,N_11736,N_11702);
xor U11793 (N_11793,N_11699,N_11719);
or U11794 (N_11794,N_11631,N_11638);
nor U11795 (N_11795,N_11681,N_11716);
nor U11796 (N_11796,N_11642,N_11662);
and U11797 (N_11797,N_11649,N_11709);
xnor U11798 (N_11798,N_11670,N_11632);
nand U11799 (N_11799,N_11651,N_11692);
or U11800 (N_11800,N_11650,N_11727);
nor U11801 (N_11801,N_11698,N_11674);
and U11802 (N_11802,N_11721,N_11653);
or U11803 (N_11803,N_11733,N_11723);
or U11804 (N_11804,N_11645,N_11628);
nand U11805 (N_11805,N_11737,N_11630);
nor U11806 (N_11806,N_11686,N_11728);
or U11807 (N_11807,N_11710,N_11675);
or U11808 (N_11808,N_11690,N_11747);
and U11809 (N_11809,N_11673,N_11641);
xnor U11810 (N_11810,N_11732,N_11636);
or U11811 (N_11811,N_11671,N_11722);
nor U11812 (N_11812,N_11720,N_11635);
nor U11813 (N_11813,N_11650,N_11749);
nor U11814 (N_11814,N_11661,N_11664);
nor U11815 (N_11815,N_11716,N_11663);
nor U11816 (N_11816,N_11649,N_11636);
xor U11817 (N_11817,N_11744,N_11637);
and U11818 (N_11818,N_11652,N_11680);
nor U11819 (N_11819,N_11705,N_11656);
or U11820 (N_11820,N_11669,N_11729);
xnor U11821 (N_11821,N_11686,N_11627);
nand U11822 (N_11822,N_11737,N_11720);
nor U11823 (N_11823,N_11727,N_11730);
or U11824 (N_11824,N_11690,N_11714);
nand U11825 (N_11825,N_11690,N_11650);
or U11826 (N_11826,N_11681,N_11678);
nand U11827 (N_11827,N_11637,N_11732);
nor U11828 (N_11828,N_11629,N_11745);
xor U11829 (N_11829,N_11626,N_11726);
nor U11830 (N_11830,N_11717,N_11653);
xnor U11831 (N_11831,N_11743,N_11700);
xnor U11832 (N_11832,N_11688,N_11639);
or U11833 (N_11833,N_11674,N_11723);
nor U11834 (N_11834,N_11669,N_11733);
or U11835 (N_11835,N_11703,N_11733);
or U11836 (N_11836,N_11664,N_11672);
and U11837 (N_11837,N_11644,N_11732);
nand U11838 (N_11838,N_11739,N_11671);
or U11839 (N_11839,N_11698,N_11712);
nor U11840 (N_11840,N_11689,N_11652);
nor U11841 (N_11841,N_11635,N_11690);
and U11842 (N_11842,N_11677,N_11689);
xor U11843 (N_11843,N_11700,N_11665);
xor U11844 (N_11844,N_11653,N_11683);
nand U11845 (N_11845,N_11695,N_11631);
xnor U11846 (N_11846,N_11657,N_11700);
and U11847 (N_11847,N_11734,N_11742);
nand U11848 (N_11848,N_11736,N_11748);
or U11849 (N_11849,N_11653,N_11647);
nand U11850 (N_11850,N_11680,N_11644);
and U11851 (N_11851,N_11676,N_11678);
or U11852 (N_11852,N_11636,N_11700);
xnor U11853 (N_11853,N_11741,N_11636);
nand U11854 (N_11854,N_11667,N_11741);
nand U11855 (N_11855,N_11715,N_11725);
nor U11856 (N_11856,N_11661,N_11679);
xnor U11857 (N_11857,N_11703,N_11640);
nand U11858 (N_11858,N_11676,N_11699);
or U11859 (N_11859,N_11741,N_11716);
nand U11860 (N_11860,N_11742,N_11741);
and U11861 (N_11861,N_11638,N_11693);
and U11862 (N_11862,N_11716,N_11721);
nor U11863 (N_11863,N_11644,N_11687);
nand U11864 (N_11864,N_11733,N_11683);
and U11865 (N_11865,N_11659,N_11747);
nor U11866 (N_11866,N_11663,N_11748);
and U11867 (N_11867,N_11735,N_11668);
xnor U11868 (N_11868,N_11742,N_11728);
xnor U11869 (N_11869,N_11653,N_11642);
or U11870 (N_11870,N_11746,N_11693);
xnor U11871 (N_11871,N_11660,N_11684);
xnor U11872 (N_11872,N_11646,N_11641);
xnor U11873 (N_11873,N_11748,N_11696);
and U11874 (N_11874,N_11704,N_11703);
and U11875 (N_11875,N_11760,N_11794);
nand U11876 (N_11876,N_11751,N_11812);
xnor U11877 (N_11877,N_11795,N_11790);
xnor U11878 (N_11878,N_11852,N_11857);
nor U11879 (N_11879,N_11769,N_11842);
xnor U11880 (N_11880,N_11797,N_11858);
xor U11881 (N_11881,N_11800,N_11785);
or U11882 (N_11882,N_11856,N_11758);
nand U11883 (N_11883,N_11796,N_11848);
xor U11884 (N_11884,N_11819,N_11825);
and U11885 (N_11885,N_11777,N_11839);
nand U11886 (N_11886,N_11836,N_11844);
nand U11887 (N_11887,N_11798,N_11754);
nand U11888 (N_11888,N_11768,N_11780);
xnor U11889 (N_11889,N_11789,N_11764);
xnor U11890 (N_11890,N_11775,N_11772);
and U11891 (N_11891,N_11787,N_11820);
or U11892 (N_11892,N_11869,N_11784);
and U11893 (N_11893,N_11763,N_11770);
or U11894 (N_11894,N_11782,N_11791);
xnor U11895 (N_11895,N_11783,N_11823);
xnor U11896 (N_11896,N_11854,N_11843);
xnor U11897 (N_11897,N_11830,N_11771);
nor U11898 (N_11898,N_11805,N_11828);
nand U11899 (N_11899,N_11861,N_11774);
or U11900 (N_11900,N_11827,N_11803);
nor U11901 (N_11901,N_11855,N_11753);
and U11902 (N_11902,N_11809,N_11851);
or U11903 (N_11903,N_11865,N_11802);
and U11904 (N_11904,N_11792,N_11807);
nor U11905 (N_11905,N_11831,N_11871);
nand U11906 (N_11906,N_11817,N_11847);
or U11907 (N_11907,N_11779,N_11860);
and U11908 (N_11908,N_11850,N_11821);
or U11909 (N_11909,N_11873,N_11818);
nor U11910 (N_11910,N_11813,N_11845);
and U11911 (N_11911,N_11755,N_11781);
nor U11912 (N_11912,N_11824,N_11838);
and U11913 (N_11913,N_11799,N_11846);
xor U11914 (N_11914,N_11756,N_11810);
nor U11915 (N_11915,N_11866,N_11833);
nor U11916 (N_11916,N_11766,N_11867);
or U11917 (N_11917,N_11874,N_11868);
nand U11918 (N_11918,N_11816,N_11829);
and U11919 (N_11919,N_11822,N_11804);
and U11920 (N_11920,N_11835,N_11761);
and U11921 (N_11921,N_11837,N_11786);
nor U11922 (N_11922,N_11862,N_11808);
or U11923 (N_11923,N_11849,N_11759);
xnor U11924 (N_11924,N_11757,N_11870);
nor U11925 (N_11925,N_11864,N_11762);
nand U11926 (N_11926,N_11752,N_11788);
or U11927 (N_11927,N_11801,N_11765);
or U11928 (N_11928,N_11853,N_11834);
and U11929 (N_11929,N_11832,N_11841);
nand U11930 (N_11930,N_11814,N_11859);
and U11931 (N_11931,N_11840,N_11806);
or U11932 (N_11932,N_11826,N_11767);
xnor U11933 (N_11933,N_11750,N_11778);
or U11934 (N_11934,N_11872,N_11863);
or U11935 (N_11935,N_11773,N_11815);
nor U11936 (N_11936,N_11793,N_11776);
nor U11937 (N_11937,N_11811,N_11858);
nand U11938 (N_11938,N_11782,N_11832);
or U11939 (N_11939,N_11823,N_11770);
and U11940 (N_11940,N_11777,N_11836);
xnor U11941 (N_11941,N_11788,N_11842);
nor U11942 (N_11942,N_11818,N_11824);
nor U11943 (N_11943,N_11833,N_11854);
xor U11944 (N_11944,N_11841,N_11795);
nand U11945 (N_11945,N_11797,N_11783);
xnor U11946 (N_11946,N_11793,N_11853);
nand U11947 (N_11947,N_11777,N_11811);
xor U11948 (N_11948,N_11795,N_11755);
nand U11949 (N_11949,N_11751,N_11774);
and U11950 (N_11950,N_11851,N_11861);
xnor U11951 (N_11951,N_11863,N_11822);
nand U11952 (N_11952,N_11849,N_11826);
xnor U11953 (N_11953,N_11851,N_11813);
nand U11954 (N_11954,N_11840,N_11809);
or U11955 (N_11955,N_11753,N_11754);
or U11956 (N_11956,N_11806,N_11780);
or U11957 (N_11957,N_11810,N_11787);
xor U11958 (N_11958,N_11786,N_11799);
and U11959 (N_11959,N_11799,N_11866);
and U11960 (N_11960,N_11785,N_11862);
or U11961 (N_11961,N_11790,N_11775);
nand U11962 (N_11962,N_11801,N_11779);
or U11963 (N_11963,N_11755,N_11863);
or U11964 (N_11964,N_11758,N_11771);
and U11965 (N_11965,N_11800,N_11828);
xor U11966 (N_11966,N_11803,N_11871);
or U11967 (N_11967,N_11811,N_11790);
nand U11968 (N_11968,N_11823,N_11763);
or U11969 (N_11969,N_11766,N_11767);
or U11970 (N_11970,N_11782,N_11779);
and U11971 (N_11971,N_11774,N_11755);
and U11972 (N_11972,N_11861,N_11776);
and U11973 (N_11973,N_11753,N_11826);
nand U11974 (N_11974,N_11761,N_11845);
nand U11975 (N_11975,N_11785,N_11767);
or U11976 (N_11976,N_11816,N_11848);
and U11977 (N_11977,N_11780,N_11751);
xor U11978 (N_11978,N_11871,N_11816);
and U11979 (N_11979,N_11867,N_11751);
nor U11980 (N_11980,N_11791,N_11825);
and U11981 (N_11981,N_11790,N_11802);
or U11982 (N_11982,N_11837,N_11838);
nand U11983 (N_11983,N_11790,N_11808);
or U11984 (N_11984,N_11758,N_11843);
and U11985 (N_11985,N_11817,N_11759);
and U11986 (N_11986,N_11856,N_11771);
or U11987 (N_11987,N_11817,N_11778);
and U11988 (N_11988,N_11777,N_11874);
xor U11989 (N_11989,N_11764,N_11750);
nand U11990 (N_11990,N_11800,N_11752);
or U11991 (N_11991,N_11872,N_11768);
or U11992 (N_11992,N_11756,N_11803);
and U11993 (N_11993,N_11850,N_11866);
xor U11994 (N_11994,N_11772,N_11820);
or U11995 (N_11995,N_11841,N_11783);
or U11996 (N_11996,N_11854,N_11828);
and U11997 (N_11997,N_11807,N_11797);
and U11998 (N_11998,N_11846,N_11838);
xnor U11999 (N_11999,N_11796,N_11852);
nand U12000 (N_12000,N_11909,N_11884);
and U12001 (N_12001,N_11919,N_11902);
or U12002 (N_12002,N_11979,N_11876);
or U12003 (N_12003,N_11958,N_11956);
nor U12004 (N_12004,N_11947,N_11999);
nor U12005 (N_12005,N_11975,N_11997);
nand U12006 (N_12006,N_11966,N_11996);
or U12007 (N_12007,N_11901,N_11887);
or U12008 (N_12008,N_11922,N_11913);
nor U12009 (N_12009,N_11886,N_11904);
nor U12010 (N_12010,N_11993,N_11944);
nand U12011 (N_12011,N_11957,N_11916);
nor U12012 (N_12012,N_11936,N_11917);
or U12013 (N_12013,N_11959,N_11881);
or U12014 (N_12014,N_11991,N_11908);
and U12015 (N_12015,N_11998,N_11896);
or U12016 (N_12016,N_11970,N_11923);
or U12017 (N_12017,N_11903,N_11983);
or U12018 (N_12018,N_11973,N_11948);
and U12019 (N_12019,N_11920,N_11927);
nor U12020 (N_12020,N_11945,N_11971);
or U12021 (N_12021,N_11982,N_11985);
and U12022 (N_12022,N_11955,N_11926);
nor U12023 (N_12023,N_11931,N_11933);
nand U12024 (N_12024,N_11967,N_11883);
nor U12025 (N_12025,N_11877,N_11937);
and U12026 (N_12026,N_11925,N_11914);
nand U12027 (N_12027,N_11885,N_11981);
nor U12028 (N_12028,N_11964,N_11974);
and U12029 (N_12029,N_11978,N_11995);
or U12030 (N_12030,N_11895,N_11953);
nor U12031 (N_12031,N_11880,N_11907);
nand U12032 (N_12032,N_11889,N_11992);
xnor U12033 (N_12033,N_11888,N_11951);
xor U12034 (N_12034,N_11977,N_11911);
or U12035 (N_12035,N_11934,N_11952);
xor U12036 (N_12036,N_11879,N_11950);
and U12037 (N_12037,N_11900,N_11891);
nand U12038 (N_12038,N_11980,N_11898);
xor U12039 (N_12039,N_11930,N_11939);
nor U12040 (N_12040,N_11942,N_11924);
nor U12041 (N_12041,N_11882,N_11962);
xor U12042 (N_12042,N_11943,N_11986);
xor U12043 (N_12043,N_11935,N_11938);
nor U12044 (N_12044,N_11912,N_11890);
and U12045 (N_12045,N_11893,N_11961);
nand U12046 (N_12046,N_11894,N_11954);
nand U12047 (N_12047,N_11932,N_11892);
nor U12048 (N_12048,N_11960,N_11940);
xor U12049 (N_12049,N_11918,N_11878);
nand U12050 (N_12050,N_11910,N_11928);
and U12051 (N_12051,N_11941,N_11915);
or U12052 (N_12052,N_11875,N_11929);
nor U12053 (N_12053,N_11976,N_11989);
and U12054 (N_12054,N_11990,N_11899);
and U12055 (N_12055,N_11963,N_11946);
xor U12056 (N_12056,N_11905,N_11972);
nor U12057 (N_12057,N_11987,N_11984);
and U12058 (N_12058,N_11897,N_11906);
nor U12059 (N_12059,N_11969,N_11994);
or U12060 (N_12060,N_11988,N_11921);
or U12061 (N_12061,N_11965,N_11949);
nor U12062 (N_12062,N_11968,N_11915);
or U12063 (N_12063,N_11978,N_11964);
nand U12064 (N_12064,N_11968,N_11913);
or U12065 (N_12065,N_11954,N_11920);
xor U12066 (N_12066,N_11971,N_11979);
and U12067 (N_12067,N_11912,N_11937);
or U12068 (N_12068,N_11972,N_11932);
xor U12069 (N_12069,N_11984,N_11897);
nor U12070 (N_12070,N_11939,N_11997);
nand U12071 (N_12071,N_11993,N_11987);
or U12072 (N_12072,N_11886,N_11939);
nand U12073 (N_12073,N_11931,N_11875);
nor U12074 (N_12074,N_11940,N_11963);
nand U12075 (N_12075,N_11917,N_11909);
nor U12076 (N_12076,N_11907,N_11925);
and U12077 (N_12077,N_11998,N_11918);
nor U12078 (N_12078,N_11918,N_11993);
and U12079 (N_12079,N_11953,N_11987);
or U12080 (N_12080,N_11902,N_11927);
xnor U12081 (N_12081,N_11969,N_11989);
or U12082 (N_12082,N_11884,N_11951);
nand U12083 (N_12083,N_11958,N_11924);
nand U12084 (N_12084,N_11975,N_11906);
and U12085 (N_12085,N_11998,N_11913);
nor U12086 (N_12086,N_11887,N_11943);
xor U12087 (N_12087,N_11975,N_11880);
nor U12088 (N_12088,N_11887,N_11998);
or U12089 (N_12089,N_11883,N_11953);
or U12090 (N_12090,N_11891,N_11964);
and U12091 (N_12091,N_11923,N_11969);
xnor U12092 (N_12092,N_11934,N_11975);
or U12093 (N_12093,N_11907,N_11875);
nor U12094 (N_12094,N_11951,N_11892);
xor U12095 (N_12095,N_11929,N_11993);
nand U12096 (N_12096,N_11986,N_11909);
nor U12097 (N_12097,N_11991,N_11914);
and U12098 (N_12098,N_11991,N_11898);
or U12099 (N_12099,N_11906,N_11928);
nand U12100 (N_12100,N_11963,N_11947);
and U12101 (N_12101,N_11913,N_11941);
nand U12102 (N_12102,N_11923,N_11966);
xnor U12103 (N_12103,N_11905,N_11983);
xor U12104 (N_12104,N_11985,N_11973);
nand U12105 (N_12105,N_11880,N_11928);
nand U12106 (N_12106,N_11958,N_11977);
and U12107 (N_12107,N_11932,N_11920);
or U12108 (N_12108,N_11905,N_11932);
or U12109 (N_12109,N_11926,N_11911);
or U12110 (N_12110,N_11932,N_11965);
xor U12111 (N_12111,N_11960,N_11876);
xor U12112 (N_12112,N_11880,N_11990);
nand U12113 (N_12113,N_11967,N_11943);
and U12114 (N_12114,N_11971,N_11884);
nand U12115 (N_12115,N_11924,N_11899);
nor U12116 (N_12116,N_11919,N_11896);
nand U12117 (N_12117,N_11905,N_11920);
nand U12118 (N_12118,N_11883,N_11943);
nor U12119 (N_12119,N_11908,N_11945);
nor U12120 (N_12120,N_11879,N_11985);
and U12121 (N_12121,N_11908,N_11990);
nand U12122 (N_12122,N_11924,N_11969);
and U12123 (N_12123,N_11998,N_11934);
and U12124 (N_12124,N_11984,N_11875);
nand U12125 (N_12125,N_12034,N_12022);
nor U12126 (N_12126,N_12026,N_12063);
or U12127 (N_12127,N_12083,N_12005);
xor U12128 (N_12128,N_12077,N_12082);
nand U12129 (N_12129,N_12067,N_12046);
nand U12130 (N_12130,N_12015,N_12049);
nand U12131 (N_12131,N_12110,N_12021);
and U12132 (N_12132,N_12091,N_12070);
or U12133 (N_12133,N_12030,N_12045);
and U12134 (N_12134,N_12039,N_12016);
nor U12135 (N_12135,N_12102,N_12087);
and U12136 (N_12136,N_12074,N_12117);
and U12137 (N_12137,N_12081,N_12120);
or U12138 (N_12138,N_12088,N_12001);
and U12139 (N_12139,N_12116,N_12057);
xnor U12140 (N_12140,N_12024,N_12047);
or U12141 (N_12141,N_12095,N_12111);
xor U12142 (N_12142,N_12031,N_12028);
or U12143 (N_12143,N_12094,N_12037);
nand U12144 (N_12144,N_12086,N_12056);
and U12145 (N_12145,N_12112,N_12059);
xor U12146 (N_12146,N_12084,N_12004);
and U12147 (N_12147,N_12010,N_12002);
nand U12148 (N_12148,N_12055,N_12052);
xor U12149 (N_12149,N_12012,N_12007);
nand U12150 (N_12150,N_12044,N_12036);
nor U12151 (N_12151,N_12108,N_12043);
nand U12152 (N_12152,N_12068,N_12027);
or U12153 (N_12153,N_12103,N_12064);
nor U12154 (N_12154,N_12080,N_12060);
xnor U12155 (N_12155,N_12113,N_12033);
nor U12156 (N_12156,N_12109,N_12053);
nand U12157 (N_12157,N_12099,N_12079);
nand U12158 (N_12158,N_12029,N_12096);
xnor U12159 (N_12159,N_12025,N_12048);
xor U12160 (N_12160,N_12051,N_12011);
and U12161 (N_12161,N_12089,N_12090);
and U12162 (N_12162,N_12062,N_12115);
nor U12163 (N_12163,N_12013,N_12042);
nand U12164 (N_12164,N_12100,N_12009);
and U12165 (N_12165,N_12014,N_12019);
or U12166 (N_12166,N_12093,N_12040);
nand U12167 (N_12167,N_12085,N_12000);
or U12168 (N_12168,N_12071,N_12023);
and U12169 (N_12169,N_12114,N_12078);
nand U12170 (N_12170,N_12038,N_12020);
and U12171 (N_12171,N_12050,N_12107);
or U12172 (N_12172,N_12101,N_12121);
and U12173 (N_12173,N_12123,N_12092);
nand U12174 (N_12174,N_12003,N_12097);
nand U12175 (N_12175,N_12076,N_12069);
or U12176 (N_12176,N_12072,N_12054);
and U12177 (N_12177,N_12008,N_12118);
and U12178 (N_12178,N_12018,N_12006);
nand U12179 (N_12179,N_12041,N_12106);
nand U12180 (N_12180,N_12032,N_12075);
nor U12181 (N_12181,N_12058,N_12104);
xor U12182 (N_12182,N_12066,N_12061);
nand U12183 (N_12183,N_12035,N_12124);
xnor U12184 (N_12184,N_12017,N_12119);
nand U12185 (N_12185,N_12105,N_12065);
xor U12186 (N_12186,N_12122,N_12073);
xor U12187 (N_12187,N_12098,N_12050);
nor U12188 (N_12188,N_12015,N_12095);
xnor U12189 (N_12189,N_12009,N_12084);
nor U12190 (N_12190,N_12096,N_12054);
or U12191 (N_12191,N_12078,N_12034);
or U12192 (N_12192,N_12002,N_12085);
xor U12193 (N_12193,N_12113,N_12089);
nand U12194 (N_12194,N_12015,N_12119);
or U12195 (N_12195,N_12107,N_12059);
or U12196 (N_12196,N_12124,N_12009);
xor U12197 (N_12197,N_12042,N_12000);
and U12198 (N_12198,N_12106,N_12085);
and U12199 (N_12199,N_12122,N_12124);
xor U12200 (N_12200,N_12083,N_12034);
and U12201 (N_12201,N_12118,N_12089);
and U12202 (N_12202,N_12040,N_12103);
nor U12203 (N_12203,N_12031,N_12112);
nand U12204 (N_12204,N_12028,N_12020);
nor U12205 (N_12205,N_12018,N_12031);
nand U12206 (N_12206,N_12078,N_12076);
xnor U12207 (N_12207,N_12044,N_12089);
xnor U12208 (N_12208,N_12060,N_12112);
or U12209 (N_12209,N_12121,N_12053);
nand U12210 (N_12210,N_12083,N_12101);
or U12211 (N_12211,N_12119,N_12090);
and U12212 (N_12212,N_12008,N_12102);
nor U12213 (N_12213,N_12121,N_12071);
nand U12214 (N_12214,N_12031,N_12115);
xor U12215 (N_12215,N_12004,N_12022);
nand U12216 (N_12216,N_12009,N_12034);
xnor U12217 (N_12217,N_12064,N_12049);
or U12218 (N_12218,N_12085,N_12105);
nor U12219 (N_12219,N_12057,N_12051);
nand U12220 (N_12220,N_12017,N_12065);
or U12221 (N_12221,N_12000,N_12064);
nand U12222 (N_12222,N_12063,N_12116);
nand U12223 (N_12223,N_12016,N_12070);
nand U12224 (N_12224,N_12044,N_12033);
or U12225 (N_12225,N_12085,N_12046);
nand U12226 (N_12226,N_12124,N_12034);
nand U12227 (N_12227,N_12070,N_12046);
nand U12228 (N_12228,N_12099,N_12094);
or U12229 (N_12229,N_12068,N_12070);
nand U12230 (N_12230,N_12009,N_12071);
and U12231 (N_12231,N_12117,N_12065);
xor U12232 (N_12232,N_12115,N_12105);
and U12233 (N_12233,N_12061,N_12037);
nor U12234 (N_12234,N_12118,N_12098);
xnor U12235 (N_12235,N_12123,N_12030);
nor U12236 (N_12236,N_12019,N_12053);
nand U12237 (N_12237,N_12013,N_12085);
nand U12238 (N_12238,N_12010,N_12112);
or U12239 (N_12239,N_12063,N_12095);
or U12240 (N_12240,N_12042,N_12014);
or U12241 (N_12241,N_12017,N_12046);
nand U12242 (N_12242,N_12124,N_12060);
xor U12243 (N_12243,N_12107,N_12067);
xor U12244 (N_12244,N_12094,N_12075);
nor U12245 (N_12245,N_12019,N_12067);
or U12246 (N_12246,N_12023,N_12115);
xor U12247 (N_12247,N_12123,N_12020);
or U12248 (N_12248,N_12051,N_12113);
or U12249 (N_12249,N_12040,N_12000);
or U12250 (N_12250,N_12188,N_12139);
nand U12251 (N_12251,N_12222,N_12191);
xnor U12252 (N_12252,N_12136,N_12155);
and U12253 (N_12253,N_12169,N_12197);
nand U12254 (N_12254,N_12225,N_12140);
xnor U12255 (N_12255,N_12152,N_12162);
nand U12256 (N_12256,N_12132,N_12219);
nor U12257 (N_12257,N_12226,N_12161);
nor U12258 (N_12258,N_12189,N_12202);
xor U12259 (N_12259,N_12224,N_12168);
or U12260 (N_12260,N_12178,N_12244);
and U12261 (N_12261,N_12235,N_12154);
and U12262 (N_12262,N_12172,N_12199);
nand U12263 (N_12263,N_12184,N_12227);
xnor U12264 (N_12264,N_12137,N_12249);
or U12265 (N_12265,N_12180,N_12130);
or U12266 (N_12266,N_12207,N_12181);
nor U12267 (N_12267,N_12194,N_12187);
nand U12268 (N_12268,N_12151,N_12216);
nor U12269 (N_12269,N_12241,N_12133);
xor U12270 (N_12270,N_12135,N_12170);
or U12271 (N_12271,N_12157,N_12240);
or U12272 (N_12272,N_12242,N_12159);
and U12273 (N_12273,N_12128,N_12248);
nand U12274 (N_12274,N_12156,N_12230);
nand U12275 (N_12275,N_12148,N_12210);
or U12276 (N_12276,N_12141,N_12206);
nor U12277 (N_12277,N_12218,N_12126);
nand U12278 (N_12278,N_12166,N_12174);
nand U12279 (N_12279,N_12173,N_12229);
xor U12280 (N_12280,N_12233,N_12163);
nor U12281 (N_12281,N_12131,N_12165);
nor U12282 (N_12282,N_12215,N_12238);
nand U12283 (N_12283,N_12185,N_12211);
and U12284 (N_12284,N_12196,N_12220);
xnor U12285 (N_12285,N_12212,N_12203);
nor U12286 (N_12286,N_12209,N_12147);
nand U12287 (N_12287,N_12146,N_12144);
nor U12288 (N_12288,N_12204,N_12179);
xor U12289 (N_12289,N_12205,N_12236);
xnor U12290 (N_12290,N_12186,N_12171);
and U12291 (N_12291,N_12223,N_12164);
nand U12292 (N_12292,N_12142,N_12176);
xor U12293 (N_12293,N_12198,N_12134);
or U12294 (N_12294,N_12246,N_12150);
nor U12295 (N_12295,N_12239,N_12125);
or U12296 (N_12296,N_12200,N_12231);
or U12297 (N_12297,N_12192,N_12127);
or U12298 (N_12298,N_12237,N_12217);
or U12299 (N_12299,N_12232,N_12245);
xor U12300 (N_12300,N_12149,N_12190);
and U12301 (N_12301,N_12138,N_12193);
nor U12302 (N_12302,N_12195,N_12182);
xnor U12303 (N_12303,N_12175,N_12167);
nand U12304 (N_12304,N_12234,N_12183);
nand U12305 (N_12305,N_12221,N_12208);
or U12306 (N_12306,N_12129,N_12247);
or U12307 (N_12307,N_12160,N_12201);
and U12308 (N_12308,N_12153,N_12214);
xor U12309 (N_12309,N_12145,N_12228);
or U12310 (N_12310,N_12243,N_12213);
nand U12311 (N_12311,N_12158,N_12143);
nor U12312 (N_12312,N_12177,N_12196);
or U12313 (N_12313,N_12172,N_12126);
nor U12314 (N_12314,N_12219,N_12201);
nand U12315 (N_12315,N_12236,N_12174);
nor U12316 (N_12316,N_12169,N_12227);
nor U12317 (N_12317,N_12154,N_12211);
xnor U12318 (N_12318,N_12170,N_12219);
nand U12319 (N_12319,N_12139,N_12138);
nand U12320 (N_12320,N_12168,N_12140);
or U12321 (N_12321,N_12210,N_12132);
nand U12322 (N_12322,N_12239,N_12238);
xor U12323 (N_12323,N_12240,N_12221);
nand U12324 (N_12324,N_12241,N_12196);
and U12325 (N_12325,N_12210,N_12246);
nor U12326 (N_12326,N_12200,N_12169);
xor U12327 (N_12327,N_12135,N_12236);
nand U12328 (N_12328,N_12232,N_12218);
nor U12329 (N_12329,N_12167,N_12143);
nor U12330 (N_12330,N_12138,N_12187);
nand U12331 (N_12331,N_12236,N_12211);
xnor U12332 (N_12332,N_12164,N_12239);
or U12333 (N_12333,N_12125,N_12155);
xnor U12334 (N_12334,N_12181,N_12184);
or U12335 (N_12335,N_12200,N_12235);
xor U12336 (N_12336,N_12246,N_12226);
and U12337 (N_12337,N_12144,N_12205);
and U12338 (N_12338,N_12198,N_12242);
and U12339 (N_12339,N_12210,N_12137);
xor U12340 (N_12340,N_12203,N_12137);
and U12341 (N_12341,N_12178,N_12196);
nand U12342 (N_12342,N_12233,N_12193);
or U12343 (N_12343,N_12219,N_12156);
and U12344 (N_12344,N_12157,N_12243);
or U12345 (N_12345,N_12165,N_12222);
xnor U12346 (N_12346,N_12232,N_12187);
nor U12347 (N_12347,N_12179,N_12249);
or U12348 (N_12348,N_12193,N_12174);
nand U12349 (N_12349,N_12248,N_12161);
nand U12350 (N_12350,N_12150,N_12199);
xnor U12351 (N_12351,N_12136,N_12232);
nand U12352 (N_12352,N_12183,N_12166);
nor U12353 (N_12353,N_12245,N_12125);
or U12354 (N_12354,N_12140,N_12196);
nor U12355 (N_12355,N_12145,N_12216);
xor U12356 (N_12356,N_12185,N_12133);
nand U12357 (N_12357,N_12229,N_12226);
or U12358 (N_12358,N_12203,N_12133);
nor U12359 (N_12359,N_12214,N_12142);
or U12360 (N_12360,N_12126,N_12221);
nand U12361 (N_12361,N_12247,N_12145);
nor U12362 (N_12362,N_12175,N_12215);
nor U12363 (N_12363,N_12179,N_12169);
or U12364 (N_12364,N_12186,N_12202);
nor U12365 (N_12365,N_12175,N_12176);
or U12366 (N_12366,N_12226,N_12201);
and U12367 (N_12367,N_12130,N_12155);
nor U12368 (N_12368,N_12235,N_12191);
nand U12369 (N_12369,N_12235,N_12219);
xor U12370 (N_12370,N_12194,N_12236);
nand U12371 (N_12371,N_12205,N_12187);
nor U12372 (N_12372,N_12144,N_12180);
xnor U12373 (N_12373,N_12156,N_12200);
nor U12374 (N_12374,N_12234,N_12246);
or U12375 (N_12375,N_12372,N_12367);
and U12376 (N_12376,N_12337,N_12250);
and U12377 (N_12377,N_12345,N_12319);
and U12378 (N_12378,N_12346,N_12290);
nor U12379 (N_12379,N_12327,N_12351);
or U12380 (N_12380,N_12282,N_12342);
xnor U12381 (N_12381,N_12276,N_12285);
or U12382 (N_12382,N_12353,N_12279);
and U12383 (N_12383,N_12366,N_12274);
nand U12384 (N_12384,N_12317,N_12266);
and U12385 (N_12385,N_12368,N_12336);
nor U12386 (N_12386,N_12303,N_12340);
or U12387 (N_12387,N_12326,N_12309);
nand U12388 (N_12388,N_12289,N_12257);
nor U12389 (N_12389,N_12329,N_12272);
and U12390 (N_12390,N_12271,N_12305);
or U12391 (N_12391,N_12341,N_12295);
nor U12392 (N_12392,N_12347,N_12297);
and U12393 (N_12393,N_12253,N_12314);
nor U12394 (N_12394,N_12362,N_12334);
and U12395 (N_12395,N_12356,N_12322);
xor U12396 (N_12396,N_12361,N_12269);
nand U12397 (N_12397,N_12335,N_12344);
and U12398 (N_12398,N_12275,N_12306);
or U12399 (N_12399,N_12291,N_12267);
xnor U12400 (N_12400,N_12312,N_12350);
and U12401 (N_12401,N_12251,N_12349);
or U12402 (N_12402,N_12281,N_12254);
nor U12403 (N_12403,N_12352,N_12287);
and U12404 (N_12404,N_12359,N_12308);
and U12405 (N_12405,N_12283,N_12354);
nor U12406 (N_12406,N_12262,N_12311);
and U12407 (N_12407,N_12255,N_12265);
or U12408 (N_12408,N_12363,N_12333);
and U12409 (N_12409,N_12286,N_12320);
nor U12410 (N_12410,N_12364,N_12302);
nand U12411 (N_12411,N_12338,N_12298);
nand U12412 (N_12412,N_12261,N_12256);
or U12413 (N_12413,N_12260,N_12316);
nand U12414 (N_12414,N_12371,N_12370);
and U12415 (N_12415,N_12277,N_12328);
nand U12416 (N_12416,N_12358,N_12325);
nor U12417 (N_12417,N_12284,N_12264);
nand U12418 (N_12418,N_12296,N_12331);
or U12419 (N_12419,N_12357,N_12343);
and U12420 (N_12420,N_12365,N_12373);
nand U12421 (N_12421,N_12330,N_12355);
nand U12422 (N_12422,N_12299,N_12307);
nand U12423 (N_12423,N_12324,N_12263);
nand U12424 (N_12424,N_12339,N_12252);
nand U12425 (N_12425,N_12323,N_12360);
or U12426 (N_12426,N_12374,N_12258);
and U12427 (N_12427,N_12369,N_12313);
or U12428 (N_12428,N_12273,N_12301);
nor U12429 (N_12429,N_12315,N_12318);
or U12430 (N_12430,N_12332,N_12292);
or U12431 (N_12431,N_12278,N_12304);
nor U12432 (N_12432,N_12321,N_12270);
and U12433 (N_12433,N_12294,N_12288);
nor U12434 (N_12434,N_12259,N_12280);
xnor U12435 (N_12435,N_12300,N_12293);
and U12436 (N_12436,N_12268,N_12310);
nor U12437 (N_12437,N_12348,N_12260);
and U12438 (N_12438,N_12325,N_12364);
xnor U12439 (N_12439,N_12364,N_12313);
and U12440 (N_12440,N_12253,N_12313);
xor U12441 (N_12441,N_12352,N_12253);
or U12442 (N_12442,N_12348,N_12330);
or U12443 (N_12443,N_12293,N_12312);
and U12444 (N_12444,N_12334,N_12298);
xnor U12445 (N_12445,N_12265,N_12256);
xnor U12446 (N_12446,N_12347,N_12336);
nand U12447 (N_12447,N_12261,N_12268);
and U12448 (N_12448,N_12363,N_12338);
and U12449 (N_12449,N_12360,N_12365);
xor U12450 (N_12450,N_12334,N_12363);
nor U12451 (N_12451,N_12357,N_12335);
nand U12452 (N_12452,N_12271,N_12350);
nor U12453 (N_12453,N_12266,N_12371);
xnor U12454 (N_12454,N_12343,N_12262);
nand U12455 (N_12455,N_12255,N_12341);
or U12456 (N_12456,N_12284,N_12285);
nand U12457 (N_12457,N_12258,N_12312);
and U12458 (N_12458,N_12253,N_12284);
nand U12459 (N_12459,N_12357,N_12344);
xor U12460 (N_12460,N_12277,N_12326);
nand U12461 (N_12461,N_12270,N_12361);
xor U12462 (N_12462,N_12268,N_12329);
nor U12463 (N_12463,N_12373,N_12320);
or U12464 (N_12464,N_12361,N_12333);
xor U12465 (N_12465,N_12274,N_12291);
nor U12466 (N_12466,N_12365,N_12361);
and U12467 (N_12467,N_12276,N_12250);
xnor U12468 (N_12468,N_12295,N_12314);
or U12469 (N_12469,N_12279,N_12286);
or U12470 (N_12470,N_12308,N_12258);
nand U12471 (N_12471,N_12332,N_12341);
nand U12472 (N_12472,N_12368,N_12293);
and U12473 (N_12473,N_12318,N_12356);
xnor U12474 (N_12474,N_12330,N_12285);
nand U12475 (N_12475,N_12330,N_12278);
nor U12476 (N_12476,N_12281,N_12373);
and U12477 (N_12477,N_12367,N_12276);
nand U12478 (N_12478,N_12285,N_12257);
and U12479 (N_12479,N_12321,N_12343);
and U12480 (N_12480,N_12343,N_12273);
or U12481 (N_12481,N_12289,N_12356);
and U12482 (N_12482,N_12280,N_12284);
xor U12483 (N_12483,N_12300,N_12321);
or U12484 (N_12484,N_12310,N_12307);
nor U12485 (N_12485,N_12312,N_12328);
and U12486 (N_12486,N_12333,N_12264);
or U12487 (N_12487,N_12274,N_12364);
and U12488 (N_12488,N_12285,N_12299);
or U12489 (N_12489,N_12349,N_12275);
nand U12490 (N_12490,N_12320,N_12307);
nor U12491 (N_12491,N_12367,N_12340);
xor U12492 (N_12492,N_12280,N_12252);
xor U12493 (N_12493,N_12364,N_12320);
xnor U12494 (N_12494,N_12353,N_12372);
and U12495 (N_12495,N_12350,N_12258);
or U12496 (N_12496,N_12354,N_12351);
and U12497 (N_12497,N_12303,N_12278);
xor U12498 (N_12498,N_12266,N_12285);
nor U12499 (N_12499,N_12373,N_12250);
nand U12500 (N_12500,N_12495,N_12375);
or U12501 (N_12501,N_12425,N_12427);
nor U12502 (N_12502,N_12485,N_12451);
or U12503 (N_12503,N_12464,N_12419);
or U12504 (N_12504,N_12394,N_12407);
or U12505 (N_12505,N_12404,N_12458);
xnor U12506 (N_12506,N_12418,N_12491);
and U12507 (N_12507,N_12460,N_12376);
or U12508 (N_12508,N_12417,N_12456);
or U12509 (N_12509,N_12490,N_12442);
nand U12510 (N_12510,N_12423,N_12479);
xor U12511 (N_12511,N_12422,N_12496);
or U12512 (N_12512,N_12401,N_12467);
and U12513 (N_12513,N_12444,N_12489);
nand U12514 (N_12514,N_12432,N_12492);
or U12515 (N_12515,N_12465,N_12424);
nor U12516 (N_12516,N_12450,N_12409);
and U12517 (N_12517,N_12435,N_12383);
or U12518 (N_12518,N_12457,N_12421);
and U12519 (N_12519,N_12471,N_12437);
nor U12520 (N_12520,N_12381,N_12411);
and U12521 (N_12521,N_12389,N_12396);
or U12522 (N_12522,N_12412,N_12483);
and U12523 (N_12523,N_12388,N_12497);
or U12524 (N_12524,N_12448,N_12436);
xnor U12525 (N_12525,N_12480,N_12482);
xor U12526 (N_12526,N_12443,N_12378);
or U12527 (N_12527,N_12433,N_12452);
or U12528 (N_12528,N_12453,N_12481);
nor U12529 (N_12529,N_12430,N_12382);
and U12530 (N_12530,N_12385,N_12473);
nor U12531 (N_12531,N_12403,N_12488);
and U12532 (N_12532,N_12470,N_12402);
xor U12533 (N_12533,N_12494,N_12393);
nand U12534 (N_12534,N_12397,N_12487);
nand U12535 (N_12535,N_12474,N_12416);
xnor U12536 (N_12536,N_12461,N_12472);
nand U12537 (N_12537,N_12398,N_12438);
nor U12538 (N_12538,N_12459,N_12410);
nor U12539 (N_12539,N_12447,N_12428);
nand U12540 (N_12540,N_12431,N_12399);
or U12541 (N_12541,N_12493,N_12408);
nor U12542 (N_12542,N_12420,N_12391);
xor U12543 (N_12543,N_12445,N_12414);
xor U12544 (N_12544,N_12462,N_12449);
nand U12545 (N_12545,N_12498,N_12439);
or U12546 (N_12546,N_12384,N_12466);
and U12547 (N_12547,N_12454,N_12386);
or U12548 (N_12548,N_12429,N_12406);
nor U12549 (N_12549,N_12484,N_12395);
nand U12550 (N_12550,N_12415,N_12392);
nand U12551 (N_12551,N_12468,N_12499);
nand U12552 (N_12552,N_12379,N_12387);
and U12553 (N_12553,N_12380,N_12426);
nand U12554 (N_12554,N_12469,N_12486);
xor U12555 (N_12555,N_12475,N_12377);
and U12556 (N_12556,N_12477,N_12434);
nor U12557 (N_12557,N_12476,N_12405);
nor U12558 (N_12558,N_12413,N_12400);
and U12559 (N_12559,N_12463,N_12440);
nor U12560 (N_12560,N_12455,N_12478);
and U12561 (N_12561,N_12441,N_12390);
nand U12562 (N_12562,N_12446,N_12420);
nor U12563 (N_12563,N_12395,N_12402);
or U12564 (N_12564,N_12441,N_12487);
nor U12565 (N_12565,N_12481,N_12432);
nand U12566 (N_12566,N_12440,N_12491);
xor U12567 (N_12567,N_12401,N_12431);
nand U12568 (N_12568,N_12441,N_12399);
or U12569 (N_12569,N_12427,N_12421);
or U12570 (N_12570,N_12422,N_12454);
nor U12571 (N_12571,N_12488,N_12450);
nor U12572 (N_12572,N_12425,N_12449);
xnor U12573 (N_12573,N_12425,N_12393);
nand U12574 (N_12574,N_12455,N_12399);
or U12575 (N_12575,N_12390,N_12497);
and U12576 (N_12576,N_12395,N_12453);
nand U12577 (N_12577,N_12379,N_12375);
and U12578 (N_12578,N_12426,N_12379);
nor U12579 (N_12579,N_12486,N_12480);
nand U12580 (N_12580,N_12486,N_12376);
and U12581 (N_12581,N_12416,N_12422);
nor U12582 (N_12582,N_12470,N_12399);
nand U12583 (N_12583,N_12415,N_12443);
or U12584 (N_12584,N_12441,N_12444);
xnor U12585 (N_12585,N_12480,N_12424);
and U12586 (N_12586,N_12439,N_12430);
nand U12587 (N_12587,N_12404,N_12482);
xnor U12588 (N_12588,N_12447,N_12380);
xnor U12589 (N_12589,N_12392,N_12457);
nor U12590 (N_12590,N_12408,N_12438);
and U12591 (N_12591,N_12384,N_12468);
and U12592 (N_12592,N_12375,N_12479);
nand U12593 (N_12593,N_12432,N_12448);
or U12594 (N_12594,N_12381,N_12460);
xnor U12595 (N_12595,N_12421,N_12479);
nor U12596 (N_12596,N_12406,N_12440);
nor U12597 (N_12597,N_12431,N_12440);
or U12598 (N_12598,N_12435,N_12480);
or U12599 (N_12599,N_12405,N_12443);
and U12600 (N_12600,N_12394,N_12424);
xnor U12601 (N_12601,N_12411,N_12450);
and U12602 (N_12602,N_12411,N_12460);
nor U12603 (N_12603,N_12391,N_12465);
nand U12604 (N_12604,N_12453,N_12472);
or U12605 (N_12605,N_12474,N_12464);
and U12606 (N_12606,N_12467,N_12453);
nor U12607 (N_12607,N_12491,N_12376);
nand U12608 (N_12608,N_12456,N_12459);
nor U12609 (N_12609,N_12411,N_12382);
and U12610 (N_12610,N_12477,N_12383);
xor U12611 (N_12611,N_12473,N_12438);
nor U12612 (N_12612,N_12439,N_12494);
or U12613 (N_12613,N_12456,N_12391);
xor U12614 (N_12614,N_12462,N_12400);
nand U12615 (N_12615,N_12473,N_12485);
nor U12616 (N_12616,N_12375,N_12434);
nand U12617 (N_12617,N_12416,N_12430);
nand U12618 (N_12618,N_12426,N_12425);
or U12619 (N_12619,N_12428,N_12467);
xor U12620 (N_12620,N_12499,N_12423);
xor U12621 (N_12621,N_12482,N_12486);
and U12622 (N_12622,N_12463,N_12404);
nand U12623 (N_12623,N_12413,N_12497);
nand U12624 (N_12624,N_12405,N_12468);
or U12625 (N_12625,N_12597,N_12572);
and U12626 (N_12626,N_12592,N_12599);
or U12627 (N_12627,N_12523,N_12508);
and U12628 (N_12628,N_12566,N_12500);
and U12629 (N_12629,N_12542,N_12539);
and U12630 (N_12630,N_12620,N_12547);
or U12631 (N_12631,N_12548,N_12578);
or U12632 (N_12632,N_12573,N_12504);
or U12633 (N_12633,N_12540,N_12612);
xor U12634 (N_12634,N_12513,N_12577);
nand U12635 (N_12635,N_12607,N_12619);
or U12636 (N_12636,N_12524,N_12530);
xor U12637 (N_12637,N_12502,N_12535);
nor U12638 (N_12638,N_12532,N_12518);
nor U12639 (N_12639,N_12516,N_12511);
or U12640 (N_12640,N_12580,N_12598);
and U12641 (N_12641,N_12603,N_12608);
nor U12642 (N_12642,N_12602,N_12560);
nor U12643 (N_12643,N_12503,N_12596);
nor U12644 (N_12644,N_12613,N_12550);
and U12645 (N_12645,N_12584,N_12582);
or U12646 (N_12646,N_12622,N_12543);
nor U12647 (N_12647,N_12564,N_12525);
xor U12648 (N_12648,N_12545,N_12544);
xnor U12649 (N_12649,N_12590,N_12567);
nand U12650 (N_12650,N_12534,N_12594);
xnor U12651 (N_12651,N_12616,N_12571);
nor U12652 (N_12652,N_12617,N_12521);
or U12653 (N_12653,N_12533,N_12505);
nor U12654 (N_12654,N_12558,N_12538);
xnor U12655 (N_12655,N_12606,N_12575);
or U12656 (N_12656,N_12537,N_12555);
xor U12657 (N_12657,N_12517,N_12559);
and U12658 (N_12658,N_12561,N_12589);
nand U12659 (N_12659,N_12610,N_12624);
nor U12660 (N_12660,N_12587,N_12527);
and U12661 (N_12661,N_12586,N_12552);
xnor U12662 (N_12662,N_12591,N_12536);
xnor U12663 (N_12663,N_12506,N_12614);
nor U12664 (N_12664,N_12568,N_12510);
nor U12665 (N_12665,N_12583,N_12515);
or U12666 (N_12666,N_12570,N_12593);
nand U12667 (N_12667,N_12576,N_12541);
or U12668 (N_12668,N_12512,N_12562);
nor U12669 (N_12669,N_12588,N_12509);
or U12670 (N_12670,N_12553,N_12600);
xor U12671 (N_12671,N_12531,N_12585);
nand U12672 (N_12672,N_12623,N_12581);
and U12673 (N_12673,N_12563,N_12528);
nor U12674 (N_12674,N_12569,N_12618);
xnor U12675 (N_12675,N_12615,N_12549);
and U12676 (N_12676,N_12546,N_12526);
or U12677 (N_12677,N_12514,N_12574);
nor U12678 (N_12678,N_12507,N_12557);
and U12679 (N_12679,N_12522,N_12519);
and U12680 (N_12680,N_12501,N_12565);
or U12681 (N_12681,N_12556,N_12579);
and U12682 (N_12682,N_12529,N_12601);
or U12683 (N_12683,N_12520,N_12551);
xnor U12684 (N_12684,N_12621,N_12611);
or U12685 (N_12685,N_12604,N_12554);
and U12686 (N_12686,N_12595,N_12609);
nand U12687 (N_12687,N_12605,N_12507);
or U12688 (N_12688,N_12607,N_12606);
and U12689 (N_12689,N_12616,N_12575);
xor U12690 (N_12690,N_12528,N_12598);
xor U12691 (N_12691,N_12552,N_12563);
nand U12692 (N_12692,N_12620,N_12559);
nand U12693 (N_12693,N_12617,N_12532);
and U12694 (N_12694,N_12615,N_12507);
or U12695 (N_12695,N_12570,N_12581);
nand U12696 (N_12696,N_12614,N_12513);
or U12697 (N_12697,N_12563,N_12565);
xor U12698 (N_12698,N_12588,N_12552);
nor U12699 (N_12699,N_12573,N_12549);
xor U12700 (N_12700,N_12514,N_12607);
nand U12701 (N_12701,N_12551,N_12559);
nor U12702 (N_12702,N_12603,N_12529);
nand U12703 (N_12703,N_12520,N_12576);
xnor U12704 (N_12704,N_12548,N_12505);
nor U12705 (N_12705,N_12543,N_12602);
and U12706 (N_12706,N_12605,N_12576);
nand U12707 (N_12707,N_12621,N_12574);
or U12708 (N_12708,N_12546,N_12509);
or U12709 (N_12709,N_12501,N_12530);
or U12710 (N_12710,N_12572,N_12524);
nor U12711 (N_12711,N_12572,N_12556);
or U12712 (N_12712,N_12614,N_12574);
and U12713 (N_12713,N_12605,N_12571);
nand U12714 (N_12714,N_12544,N_12595);
or U12715 (N_12715,N_12534,N_12566);
xor U12716 (N_12716,N_12534,N_12547);
nor U12717 (N_12717,N_12554,N_12579);
xor U12718 (N_12718,N_12558,N_12502);
nand U12719 (N_12719,N_12621,N_12576);
nand U12720 (N_12720,N_12620,N_12554);
xor U12721 (N_12721,N_12605,N_12564);
nor U12722 (N_12722,N_12619,N_12567);
nor U12723 (N_12723,N_12501,N_12622);
nor U12724 (N_12724,N_12527,N_12510);
nand U12725 (N_12725,N_12562,N_12593);
xnor U12726 (N_12726,N_12552,N_12619);
or U12727 (N_12727,N_12542,N_12606);
nor U12728 (N_12728,N_12517,N_12570);
nand U12729 (N_12729,N_12620,N_12577);
or U12730 (N_12730,N_12573,N_12544);
nor U12731 (N_12731,N_12542,N_12552);
and U12732 (N_12732,N_12598,N_12574);
nand U12733 (N_12733,N_12613,N_12581);
nor U12734 (N_12734,N_12533,N_12548);
and U12735 (N_12735,N_12612,N_12592);
xnor U12736 (N_12736,N_12602,N_12518);
nor U12737 (N_12737,N_12514,N_12516);
and U12738 (N_12738,N_12587,N_12574);
or U12739 (N_12739,N_12585,N_12558);
xor U12740 (N_12740,N_12560,N_12549);
or U12741 (N_12741,N_12525,N_12589);
or U12742 (N_12742,N_12533,N_12578);
or U12743 (N_12743,N_12616,N_12536);
nand U12744 (N_12744,N_12568,N_12564);
nor U12745 (N_12745,N_12507,N_12525);
nor U12746 (N_12746,N_12623,N_12562);
nand U12747 (N_12747,N_12534,N_12535);
nand U12748 (N_12748,N_12590,N_12605);
xor U12749 (N_12749,N_12572,N_12619);
nor U12750 (N_12750,N_12672,N_12735);
and U12751 (N_12751,N_12670,N_12696);
or U12752 (N_12752,N_12733,N_12652);
nor U12753 (N_12753,N_12689,N_12642);
nand U12754 (N_12754,N_12635,N_12686);
nand U12755 (N_12755,N_12747,N_12687);
xor U12756 (N_12756,N_12712,N_12692);
and U12757 (N_12757,N_12698,N_12676);
nand U12758 (N_12758,N_12721,N_12740);
xor U12759 (N_12759,N_12636,N_12629);
and U12760 (N_12760,N_12655,N_12668);
or U12761 (N_12761,N_12639,N_12677);
nand U12762 (N_12762,N_12679,N_12654);
nand U12763 (N_12763,N_12715,N_12731);
and U12764 (N_12764,N_12722,N_12660);
xnor U12765 (N_12765,N_12658,N_12625);
nor U12766 (N_12766,N_12633,N_12728);
xnor U12767 (N_12767,N_12665,N_12673);
nand U12768 (N_12768,N_12699,N_12719);
nand U12769 (N_12769,N_12709,N_12648);
xnor U12770 (N_12770,N_12637,N_12681);
and U12771 (N_12771,N_12663,N_12729);
and U12772 (N_12772,N_12697,N_12634);
and U12773 (N_12773,N_12651,N_12690);
nor U12774 (N_12774,N_12626,N_12632);
nor U12775 (N_12775,N_12678,N_12720);
and U12776 (N_12776,N_12706,N_12664);
or U12777 (N_12777,N_12666,N_12713);
nor U12778 (N_12778,N_12691,N_12630);
xor U12779 (N_12779,N_12705,N_12737);
nor U12780 (N_12780,N_12717,N_12646);
and U12781 (N_12781,N_12746,N_12742);
nor U12782 (N_12782,N_12656,N_12700);
or U12783 (N_12783,N_12744,N_12685);
or U12784 (N_12784,N_12701,N_12710);
nor U12785 (N_12785,N_12628,N_12695);
or U12786 (N_12786,N_12661,N_12640);
nand U12787 (N_12787,N_12716,N_12725);
and U12788 (N_12788,N_12743,N_12688);
and U12789 (N_12789,N_12649,N_12657);
nand U12790 (N_12790,N_12718,N_12707);
xnor U12791 (N_12791,N_12727,N_12671);
xor U12792 (N_12792,N_12683,N_12693);
xnor U12793 (N_12793,N_12674,N_12645);
xor U12794 (N_12794,N_12704,N_12730);
and U12795 (N_12795,N_12741,N_12680);
xnor U12796 (N_12796,N_12708,N_12647);
nor U12797 (N_12797,N_12749,N_12659);
nor U12798 (N_12798,N_12643,N_12662);
nand U12799 (N_12799,N_12641,N_12667);
or U12800 (N_12800,N_12711,N_12650);
xor U12801 (N_12801,N_12644,N_12702);
nor U12802 (N_12802,N_12703,N_12736);
and U12803 (N_12803,N_12675,N_12726);
or U12804 (N_12804,N_12748,N_12723);
nand U12805 (N_12805,N_12738,N_12684);
nand U12806 (N_12806,N_12653,N_12682);
nand U12807 (N_12807,N_12739,N_12745);
and U12808 (N_12808,N_12714,N_12734);
or U12809 (N_12809,N_12724,N_12669);
and U12810 (N_12810,N_12694,N_12631);
nor U12811 (N_12811,N_12638,N_12627);
nand U12812 (N_12812,N_12732,N_12712);
and U12813 (N_12813,N_12691,N_12722);
or U12814 (N_12814,N_12682,N_12736);
nor U12815 (N_12815,N_12640,N_12679);
nor U12816 (N_12816,N_12633,N_12721);
or U12817 (N_12817,N_12673,N_12630);
or U12818 (N_12818,N_12686,N_12671);
xor U12819 (N_12819,N_12665,N_12732);
nand U12820 (N_12820,N_12660,N_12748);
nor U12821 (N_12821,N_12644,N_12646);
xnor U12822 (N_12822,N_12638,N_12677);
and U12823 (N_12823,N_12637,N_12626);
nand U12824 (N_12824,N_12724,N_12691);
or U12825 (N_12825,N_12748,N_12647);
and U12826 (N_12826,N_12717,N_12737);
nor U12827 (N_12827,N_12710,N_12694);
and U12828 (N_12828,N_12701,N_12714);
nand U12829 (N_12829,N_12738,N_12743);
nand U12830 (N_12830,N_12731,N_12625);
xor U12831 (N_12831,N_12737,N_12744);
nand U12832 (N_12832,N_12732,N_12667);
or U12833 (N_12833,N_12740,N_12677);
or U12834 (N_12834,N_12730,N_12666);
or U12835 (N_12835,N_12646,N_12696);
and U12836 (N_12836,N_12633,N_12727);
and U12837 (N_12837,N_12717,N_12638);
nor U12838 (N_12838,N_12686,N_12740);
and U12839 (N_12839,N_12646,N_12733);
xnor U12840 (N_12840,N_12655,N_12635);
or U12841 (N_12841,N_12695,N_12702);
or U12842 (N_12842,N_12691,N_12685);
nand U12843 (N_12843,N_12704,N_12720);
xnor U12844 (N_12844,N_12721,N_12698);
nor U12845 (N_12845,N_12708,N_12721);
and U12846 (N_12846,N_12681,N_12679);
nand U12847 (N_12847,N_12652,N_12684);
nand U12848 (N_12848,N_12666,N_12688);
or U12849 (N_12849,N_12702,N_12736);
xor U12850 (N_12850,N_12655,N_12682);
or U12851 (N_12851,N_12654,N_12631);
xor U12852 (N_12852,N_12668,N_12705);
nor U12853 (N_12853,N_12740,N_12712);
xor U12854 (N_12854,N_12630,N_12715);
nand U12855 (N_12855,N_12709,N_12645);
and U12856 (N_12856,N_12712,N_12655);
nand U12857 (N_12857,N_12650,N_12669);
xnor U12858 (N_12858,N_12735,N_12712);
nor U12859 (N_12859,N_12717,N_12671);
xor U12860 (N_12860,N_12635,N_12700);
nor U12861 (N_12861,N_12629,N_12660);
and U12862 (N_12862,N_12749,N_12696);
nand U12863 (N_12863,N_12746,N_12636);
xnor U12864 (N_12864,N_12663,N_12725);
and U12865 (N_12865,N_12657,N_12728);
nand U12866 (N_12866,N_12669,N_12694);
nor U12867 (N_12867,N_12720,N_12723);
nor U12868 (N_12868,N_12663,N_12673);
or U12869 (N_12869,N_12704,N_12693);
nor U12870 (N_12870,N_12681,N_12661);
xor U12871 (N_12871,N_12646,N_12697);
xnor U12872 (N_12872,N_12630,N_12694);
xnor U12873 (N_12873,N_12730,N_12640);
and U12874 (N_12874,N_12628,N_12657);
nor U12875 (N_12875,N_12820,N_12851);
and U12876 (N_12876,N_12765,N_12773);
nor U12877 (N_12877,N_12796,N_12756);
xnor U12878 (N_12878,N_12757,N_12872);
nand U12879 (N_12879,N_12811,N_12784);
and U12880 (N_12880,N_12809,N_12845);
and U12881 (N_12881,N_12803,N_12831);
or U12882 (N_12882,N_12868,N_12846);
or U12883 (N_12883,N_12821,N_12825);
nor U12884 (N_12884,N_12813,N_12838);
or U12885 (N_12885,N_12830,N_12865);
and U12886 (N_12886,N_12815,N_12869);
nor U12887 (N_12887,N_12853,N_12754);
nor U12888 (N_12888,N_12807,N_12769);
nand U12889 (N_12889,N_12871,N_12836);
xnor U12890 (N_12890,N_12782,N_12789);
nand U12891 (N_12891,N_12827,N_12823);
or U12892 (N_12892,N_12844,N_12818);
xor U12893 (N_12893,N_12839,N_12849);
or U12894 (N_12894,N_12814,N_12762);
and U12895 (N_12895,N_12800,N_12771);
nor U12896 (N_12896,N_12842,N_12753);
nor U12897 (N_12897,N_12874,N_12778);
xor U12898 (N_12898,N_12774,N_12794);
nor U12899 (N_12899,N_12755,N_12834);
and U12900 (N_12900,N_12768,N_12828);
or U12901 (N_12901,N_12788,N_12858);
nand U12902 (N_12902,N_12783,N_12867);
or U12903 (N_12903,N_12801,N_12819);
nand U12904 (N_12904,N_12856,N_12799);
nand U12905 (N_12905,N_12781,N_12824);
nor U12906 (N_12906,N_12861,N_12862);
nand U12907 (N_12907,N_12841,N_12863);
nand U12908 (N_12908,N_12837,N_12776);
nand U12909 (N_12909,N_12750,N_12751);
and U12910 (N_12910,N_12767,N_12864);
nand U12911 (N_12911,N_12848,N_12805);
nor U12912 (N_12912,N_12840,N_12835);
xnor U12913 (N_12913,N_12760,N_12772);
nor U12914 (N_12914,N_12870,N_12787);
nand U12915 (N_12915,N_12855,N_12764);
nand U12916 (N_12916,N_12822,N_12775);
nand U12917 (N_12917,N_12866,N_12804);
or U12918 (N_12918,N_12843,N_12857);
or U12919 (N_12919,N_12790,N_12797);
or U12920 (N_12920,N_12816,N_12763);
xnor U12921 (N_12921,N_12829,N_12770);
nand U12922 (N_12922,N_12817,N_12798);
xnor U12923 (N_12923,N_12810,N_12854);
or U12924 (N_12924,N_12780,N_12777);
or U12925 (N_12925,N_12832,N_12766);
or U12926 (N_12926,N_12850,N_12873);
or U12927 (N_12927,N_12759,N_12852);
and U12928 (N_12928,N_12808,N_12758);
nor U12929 (N_12929,N_12793,N_12826);
nor U12930 (N_12930,N_12792,N_12761);
or U12931 (N_12931,N_12785,N_12779);
or U12932 (N_12932,N_12791,N_12833);
nand U12933 (N_12933,N_12786,N_12752);
and U12934 (N_12934,N_12806,N_12860);
or U12935 (N_12935,N_12859,N_12795);
nand U12936 (N_12936,N_12812,N_12847);
nand U12937 (N_12937,N_12802,N_12850);
or U12938 (N_12938,N_12837,N_12845);
nor U12939 (N_12939,N_12823,N_12764);
xor U12940 (N_12940,N_12751,N_12767);
nor U12941 (N_12941,N_12818,N_12767);
and U12942 (N_12942,N_12785,N_12788);
and U12943 (N_12943,N_12853,N_12864);
nor U12944 (N_12944,N_12822,N_12752);
nand U12945 (N_12945,N_12786,N_12811);
and U12946 (N_12946,N_12872,N_12814);
xnor U12947 (N_12947,N_12848,N_12811);
nor U12948 (N_12948,N_12833,N_12766);
nor U12949 (N_12949,N_12757,N_12816);
and U12950 (N_12950,N_12760,N_12854);
nand U12951 (N_12951,N_12841,N_12750);
and U12952 (N_12952,N_12775,N_12806);
xor U12953 (N_12953,N_12851,N_12871);
or U12954 (N_12954,N_12873,N_12817);
and U12955 (N_12955,N_12793,N_12817);
nor U12956 (N_12956,N_12800,N_12837);
or U12957 (N_12957,N_12771,N_12798);
or U12958 (N_12958,N_12839,N_12793);
xor U12959 (N_12959,N_12836,N_12866);
xnor U12960 (N_12960,N_12796,N_12853);
nor U12961 (N_12961,N_12772,N_12823);
nor U12962 (N_12962,N_12758,N_12771);
and U12963 (N_12963,N_12860,N_12847);
nor U12964 (N_12964,N_12814,N_12764);
and U12965 (N_12965,N_12774,N_12779);
xnor U12966 (N_12966,N_12822,N_12757);
and U12967 (N_12967,N_12817,N_12770);
and U12968 (N_12968,N_12821,N_12790);
or U12969 (N_12969,N_12782,N_12832);
or U12970 (N_12970,N_12817,N_12804);
or U12971 (N_12971,N_12779,N_12769);
nand U12972 (N_12972,N_12797,N_12769);
nand U12973 (N_12973,N_12864,N_12872);
nor U12974 (N_12974,N_12797,N_12860);
nor U12975 (N_12975,N_12798,N_12763);
xor U12976 (N_12976,N_12864,N_12762);
nand U12977 (N_12977,N_12830,N_12797);
nor U12978 (N_12978,N_12867,N_12842);
or U12979 (N_12979,N_12763,N_12874);
and U12980 (N_12980,N_12843,N_12872);
nor U12981 (N_12981,N_12780,N_12791);
nor U12982 (N_12982,N_12806,N_12851);
xor U12983 (N_12983,N_12792,N_12846);
xor U12984 (N_12984,N_12758,N_12869);
nand U12985 (N_12985,N_12765,N_12786);
xnor U12986 (N_12986,N_12806,N_12804);
and U12987 (N_12987,N_12768,N_12750);
or U12988 (N_12988,N_12867,N_12836);
and U12989 (N_12989,N_12844,N_12848);
and U12990 (N_12990,N_12821,N_12812);
and U12991 (N_12991,N_12834,N_12830);
xnor U12992 (N_12992,N_12842,N_12854);
nor U12993 (N_12993,N_12809,N_12769);
xor U12994 (N_12994,N_12837,N_12868);
xnor U12995 (N_12995,N_12848,N_12769);
nand U12996 (N_12996,N_12757,N_12835);
and U12997 (N_12997,N_12790,N_12835);
or U12998 (N_12998,N_12783,N_12750);
xnor U12999 (N_12999,N_12865,N_12798);
nor U13000 (N_13000,N_12955,N_12897);
nand U13001 (N_13001,N_12941,N_12981);
nand U13002 (N_13002,N_12902,N_12893);
and U13003 (N_13003,N_12961,N_12914);
nor U13004 (N_13004,N_12948,N_12950);
or U13005 (N_13005,N_12886,N_12970);
xor U13006 (N_13006,N_12993,N_12924);
xor U13007 (N_13007,N_12982,N_12963);
or U13008 (N_13008,N_12942,N_12999);
nand U13009 (N_13009,N_12960,N_12947);
and U13010 (N_13010,N_12906,N_12883);
or U13011 (N_13011,N_12911,N_12973);
xnor U13012 (N_13012,N_12899,N_12895);
xnor U13013 (N_13013,N_12926,N_12969);
nand U13014 (N_13014,N_12908,N_12956);
or U13015 (N_13015,N_12918,N_12991);
or U13016 (N_13016,N_12916,N_12954);
nor U13017 (N_13017,N_12933,N_12976);
xor U13018 (N_13018,N_12882,N_12974);
nand U13019 (N_13019,N_12898,N_12896);
nand U13020 (N_13020,N_12940,N_12975);
xor U13021 (N_13021,N_12876,N_12998);
or U13022 (N_13022,N_12952,N_12986);
xnor U13023 (N_13023,N_12875,N_12980);
and U13024 (N_13024,N_12953,N_12965);
and U13025 (N_13025,N_12946,N_12978);
xnor U13026 (N_13026,N_12992,N_12936);
nand U13027 (N_13027,N_12892,N_12985);
nor U13028 (N_13028,N_12907,N_12909);
and U13029 (N_13029,N_12894,N_12984);
nand U13030 (N_13030,N_12905,N_12881);
nor U13031 (N_13031,N_12878,N_12917);
nand U13032 (N_13032,N_12910,N_12903);
or U13033 (N_13033,N_12901,N_12913);
nor U13034 (N_13034,N_12949,N_12915);
or U13035 (N_13035,N_12922,N_12885);
or U13036 (N_13036,N_12877,N_12925);
nand U13037 (N_13037,N_12966,N_12935);
and U13038 (N_13038,N_12964,N_12921);
and U13039 (N_13039,N_12880,N_12967);
nand U13040 (N_13040,N_12890,N_12929);
and U13041 (N_13041,N_12944,N_12928);
or U13042 (N_13042,N_12887,N_12983);
xor U13043 (N_13043,N_12962,N_12879);
and U13044 (N_13044,N_12943,N_12891);
xnor U13045 (N_13045,N_12888,N_12990);
nand U13046 (N_13046,N_12938,N_12959);
or U13047 (N_13047,N_12971,N_12932);
and U13048 (N_13048,N_12919,N_12968);
nand U13049 (N_13049,N_12937,N_12945);
nor U13050 (N_13050,N_12951,N_12997);
and U13051 (N_13051,N_12994,N_12995);
and U13052 (N_13052,N_12923,N_12934);
or U13053 (N_13053,N_12987,N_12912);
and U13054 (N_13054,N_12958,N_12957);
and U13055 (N_13055,N_12996,N_12989);
or U13056 (N_13056,N_12972,N_12977);
and U13057 (N_13057,N_12931,N_12939);
or U13058 (N_13058,N_12927,N_12889);
xnor U13059 (N_13059,N_12979,N_12884);
xor U13060 (N_13060,N_12920,N_12904);
xnor U13061 (N_13061,N_12900,N_12988);
nand U13062 (N_13062,N_12930,N_12917);
xnor U13063 (N_13063,N_12964,N_12917);
and U13064 (N_13064,N_12925,N_12989);
nor U13065 (N_13065,N_12959,N_12899);
and U13066 (N_13066,N_12984,N_12990);
nand U13067 (N_13067,N_12945,N_12995);
and U13068 (N_13068,N_12898,N_12997);
nand U13069 (N_13069,N_12900,N_12930);
nand U13070 (N_13070,N_12982,N_12936);
nor U13071 (N_13071,N_12937,N_12939);
and U13072 (N_13072,N_12949,N_12943);
or U13073 (N_13073,N_12925,N_12914);
or U13074 (N_13074,N_12943,N_12984);
or U13075 (N_13075,N_12941,N_12959);
or U13076 (N_13076,N_12899,N_12951);
and U13077 (N_13077,N_12929,N_12952);
or U13078 (N_13078,N_12911,N_12886);
nor U13079 (N_13079,N_12968,N_12897);
xnor U13080 (N_13080,N_12960,N_12951);
or U13081 (N_13081,N_12879,N_12886);
xor U13082 (N_13082,N_12993,N_12941);
and U13083 (N_13083,N_12936,N_12962);
and U13084 (N_13084,N_12898,N_12973);
nand U13085 (N_13085,N_12929,N_12990);
xor U13086 (N_13086,N_12890,N_12941);
and U13087 (N_13087,N_12944,N_12950);
xnor U13088 (N_13088,N_12883,N_12995);
or U13089 (N_13089,N_12913,N_12972);
nor U13090 (N_13090,N_12892,N_12953);
nand U13091 (N_13091,N_12939,N_12890);
nor U13092 (N_13092,N_12991,N_12946);
or U13093 (N_13093,N_12906,N_12921);
or U13094 (N_13094,N_12905,N_12922);
and U13095 (N_13095,N_12964,N_12915);
xor U13096 (N_13096,N_12979,N_12878);
nand U13097 (N_13097,N_12913,N_12965);
xnor U13098 (N_13098,N_12940,N_12976);
and U13099 (N_13099,N_12943,N_12988);
or U13100 (N_13100,N_12876,N_12886);
or U13101 (N_13101,N_12883,N_12893);
nand U13102 (N_13102,N_12913,N_12896);
xnor U13103 (N_13103,N_12912,N_12969);
xor U13104 (N_13104,N_12960,N_12918);
xnor U13105 (N_13105,N_12976,N_12968);
nor U13106 (N_13106,N_12884,N_12960);
and U13107 (N_13107,N_12928,N_12992);
nor U13108 (N_13108,N_12945,N_12943);
nor U13109 (N_13109,N_12930,N_12943);
xor U13110 (N_13110,N_12920,N_12905);
nor U13111 (N_13111,N_12895,N_12950);
and U13112 (N_13112,N_12904,N_12929);
nor U13113 (N_13113,N_12989,N_12959);
nor U13114 (N_13114,N_12958,N_12998);
nand U13115 (N_13115,N_12989,N_12926);
nor U13116 (N_13116,N_12911,N_12889);
and U13117 (N_13117,N_12926,N_12886);
and U13118 (N_13118,N_12958,N_12929);
xor U13119 (N_13119,N_12953,N_12941);
and U13120 (N_13120,N_12954,N_12904);
and U13121 (N_13121,N_12938,N_12897);
nand U13122 (N_13122,N_12876,N_12971);
nand U13123 (N_13123,N_12930,N_12905);
xor U13124 (N_13124,N_12948,N_12912);
nand U13125 (N_13125,N_13001,N_13048);
xor U13126 (N_13126,N_13116,N_13089);
nor U13127 (N_13127,N_13092,N_13099);
and U13128 (N_13128,N_13014,N_13054);
nand U13129 (N_13129,N_13007,N_13060);
nor U13130 (N_13130,N_13055,N_13062);
nand U13131 (N_13131,N_13073,N_13041);
nand U13132 (N_13132,N_13098,N_13011);
nor U13133 (N_13133,N_13086,N_13074);
nor U13134 (N_13134,N_13077,N_13102);
or U13135 (N_13135,N_13115,N_13120);
nand U13136 (N_13136,N_13069,N_13021);
and U13137 (N_13137,N_13076,N_13033);
and U13138 (N_13138,N_13121,N_13008);
or U13139 (N_13139,N_13078,N_13020);
and U13140 (N_13140,N_13068,N_13064);
and U13141 (N_13141,N_13080,N_13058);
or U13142 (N_13142,N_13079,N_13043);
nor U13143 (N_13143,N_13059,N_13034);
nand U13144 (N_13144,N_13053,N_13114);
nor U13145 (N_13145,N_13025,N_13083);
nand U13146 (N_13146,N_13107,N_13036);
nor U13147 (N_13147,N_13090,N_13104);
and U13148 (N_13148,N_13013,N_13061);
or U13149 (N_13149,N_13087,N_13122);
nand U13150 (N_13150,N_13113,N_13112);
xnor U13151 (N_13151,N_13109,N_13091);
or U13152 (N_13152,N_13035,N_13031);
xor U13153 (N_13153,N_13046,N_13117);
nand U13154 (N_13154,N_13019,N_13032);
nand U13155 (N_13155,N_13094,N_13015);
nor U13156 (N_13156,N_13005,N_13123);
or U13157 (N_13157,N_13023,N_13044);
nor U13158 (N_13158,N_13071,N_13016);
xor U13159 (N_13159,N_13045,N_13118);
and U13160 (N_13160,N_13108,N_13063);
and U13161 (N_13161,N_13124,N_13065);
and U13162 (N_13162,N_13072,N_13085);
nor U13163 (N_13163,N_13056,N_13037);
or U13164 (N_13164,N_13017,N_13003);
nand U13165 (N_13165,N_13101,N_13002);
nand U13166 (N_13166,N_13088,N_13038);
or U13167 (N_13167,N_13051,N_13057);
or U13168 (N_13168,N_13029,N_13075);
and U13169 (N_13169,N_13027,N_13111);
xor U13170 (N_13170,N_13084,N_13040);
nand U13171 (N_13171,N_13039,N_13103);
xnor U13172 (N_13172,N_13082,N_13042);
nor U13173 (N_13173,N_13006,N_13022);
or U13174 (N_13174,N_13095,N_13018);
or U13175 (N_13175,N_13097,N_13000);
xor U13176 (N_13176,N_13047,N_13024);
nand U13177 (N_13177,N_13010,N_13067);
and U13178 (N_13178,N_13119,N_13009);
or U13179 (N_13179,N_13030,N_13106);
or U13180 (N_13180,N_13028,N_13093);
or U13181 (N_13181,N_13081,N_13012);
nor U13182 (N_13182,N_13070,N_13066);
xnor U13183 (N_13183,N_13050,N_13100);
nor U13184 (N_13184,N_13049,N_13052);
xnor U13185 (N_13185,N_13105,N_13026);
nor U13186 (N_13186,N_13110,N_13004);
or U13187 (N_13187,N_13096,N_13112);
xnor U13188 (N_13188,N_13039,N_13118);
xnor U13189 (N_13189,N_13075,N_13021);
nor U13190 (N_13190,N_13064,N_13043);
or U13191 (N_13191,N_13117,N_13110);
nand U13192 (N_13192,N_13003,N_13075);
xnor U13193 (N_13193,N_13066,N_13043);
and U13194 (N_13194,N_13094,N_13049);
xor U13195 (N_13195,N_13039,N_13116);
nor U13196 (N_13196,N_13019,N_13078);
or U13197 (N_13197,N_13106,N_13064);
xnor U13198 (N_13198,N_13017,N_13013);
and U13199 (N_13199,N_13078,N_13011);
xor U13200 (N_13200,N_13069,N_13096);
nand U13201 (N_13201,N_13048,N_13007);
and U13202 (N_13202,N_13007,N_13106);
or U13203 (N_13203,N_13035,N_13050);
nor U13204 (N_13204,N_13098,N_13073);
nor U13205 (N_13205,N_13119,N_13104);
and U13206 (N_13206,N_13084,N_13077);
xnor U13207 (N_13207,N_13075,N_13080);
and U13208 (N_13208,N_13043,N_13004);
xnor U13209 (N_13209,N_13024,N_13030);
nand U13210 (N_13210,N_13118,N_13103);
nor U13211 (N_13211,N_13014,N_13059);
nand U13212 (N_13212,N_13124,N_13009);
nand U13213 (N_13213,N_13017,N_13064);
nor U13214 (N_13214,N_13063,N_13081);
or U13215 (N_13215,N_13091,N_13061);
xor U13216 (N_13216,N_13111,N_13079);
nor U13217 (N_13217,N_13004,N_13065);
or U13218 (N_13218,N_13007,N_13088);
nor U13219 (N_13219,N_13105,N_13080);
and U13220 (N_13220,N_13123,N_13088);
nor U13221 (N_13221,N_13113,N_13067);
nor U13222 (N_13222,N_13029,N_13002);
and U13223 (N_13223,N_13026,N_13098);
nor U13224 (N_13224,N_13003,N_13065);
nand U13225 (N_13225,N_13064,N_13076);
nor U13226 (N_13226,N_13051,N_13004);
nor U13227 (N_13227,N_13068,N_13033);
or U13228 (N_13228,N_13038,N_13114);
xnor U13229 (N_13229,N_13118,N_13046);
xor U13230 (N_13230,N_13016,N_13057);
and U13231 (N_13231,N_13008,N_13054);
xor U13232 (N_13232,N_13077,N_13023);
xnor U13233 (N_13233,N_13085,N_13070);
nand U13234 (N_13234,N_13021,N_13025);
and U13235 (N_13235,N_13028,N_13099);
xnor U13236 (N_13236,N_13062,N_13032);
nor U13237 (N_13237,N_13050,N_13066);
and U13238 (N_13238,N_13123,N_13028);
and U13239 (N_13239,N_13116,N_13063);
nand U13240 (N_13240,N_13084,N_13041);
and U13241 (N_13241,N_13077,N_13049);
and U13242 (N_13242,N_13118,N_13107);
nand U13243 (N_13243,N_13081,N_13073);
and U13244 (N_13244,N_13062,N_13049);
nand U13245 (N_13245,N_13054,N_13121);
xor U13246 (N_13246,N_13088,N_13084);
or U13247 (N_13247,N_13119,N_13045);
or U13248 (N_13248,N_13092,N_13044);
or U13249 (N_13249,N_13037,N_13024);
and U13250 (N_13250,N_13213,N_13197);
and U13251 (N_13251,N_13130,N_13184);
or U13252 (N_13252,N_13149,N_13135);
nor U13253 (N_13253,N_13217,N_13139);
and U13254 (N_13254,N_13142,N_13216);
nor U13255 (N_13255,N_13179,N_13195);
and U13256 (N_13256,N_13237,N_13227);
or U13257 (N_13257,N_13206,N_13168);
and U13258 (N_13258,N_13243,N_13145);
and U13259 (N_13259,N_13157,N_13172);
nor U13260 (N_13260,N_13182,N_13245);
and U13261 (N_13261,N_13137,N_13154);
nand U13262 (N_13262,N_13189,N_13233);
nand U13263 (N_13263,N_13208,N_13235);
nor U13264 (N_13264,N_13187,N_13223);
xor U13265 (N_13265,N_13191,N_13193);
and U13266 (N_13266,N_13158,N_13221);
nor U13267 (N_13267,N_13247,N_13226);
and U13268 (N_13268,N_13238,N_13127);
and U13269 (N_13269,N_13128,N_13162);
xnor U13270 (N_13270,N_13167,N_13246);
xor U13271 (N_13271,N_13141,N_13224);
nor U13272 (N_13272,N_13210,N_13133);
nand U13273 (N_13273,N_13170,N_13180);
nand U13274 (N_13274,N_13240,N_13181);
nand U13275 (N_13275,N_13231,N_13215);
nand U13276 (N_13276,N_13196,N_13131);
or U13277 (N_13277,N_13171,N_13200);
xor U13278 (N_13278,N_13161,N_13209);
or U13279 (N_13279,N_13146,N_13136);
and U13280 (N_13280,N_13204,N_13176);
and U13281 (N_13281,N_13153,N_13165);
or U13282 (N_13282,N_13160,N_13132);
nor U13283 (N_13283,N_13152,N_13129);
nand U13284 (N_13284,N_13125,N_13178);
xor U13285 (N_13285,N_13219,N_13202);
xor U13286 (N_13286,N_13159,N_13249);
and U13287 (N_13287,N_13201,N_13232);
nor U13288 (N_13288,N_13198,N_13150);
nor U13289 (N_13289,N_13205,N_13194);
nand U13290 (N_13290,N_13175,N_13173);
or U13291 (N_13291,N_13248,N_13188);
nand U13292 (N_13292,N_13230,N_13185);
or U13293 (N_13293,N_13186,N_13163);
nor U13294 (N_13294,N_13241,N_13138);
nor U13295 (N_13295,N_13214,N_13174);
nand U13296 (N_13296,N_13242,N_13140);
nand U13297 (N_13297,N_13148,N_13164);
and U13298 (N_13298,N_13244,N_13212);
nand U13299 (N_13299,N_13151,N_13166);
xnor U13300 (N_13300,N_13218,N_13177);
nor U13301 (N_13301,N_13199,N_13239);
or U13302 (N_13302,N_13190,N_13225);
xor U13303 (N_13303,N_13222,N_13126);
or U13304 (N_13304,N_13183,N_13134);
nand U13305 (N_13305,N_13169,N_13229);
nand U13306 (N_13306,N_13228,N_13144);
or U13307 (N_13307,N_13211,N_13156);
xnor U13308 (N_13308,N_13155,N_13207);
xnor U13309 (N_13309,N_13220,N_13147);
or U13310 (N_13310,N_13234,N_13192);
and U13311 (N_13311,N_13203,N_13236);
or U13312 (N_13312,N_13143,N_13125);
nor U13313 (N_13313,N_13237,N_13166);
xnor U13314 (N_13314,N_13228,N_13158);
nor U13315 (N_13315,N_13198,N_13165);
or U13316 (N_13316,N_13176,N_13132);
and U13317 (N_13317,N_13185,N_13176);
nand U13318 (N_13318,N_13159,N_13176);
nand U13319 (N_13319,N_13246,N_13131);
nor U13320 (N_13320,N_13180,N_13213);
xnor U13321 (N_13321,N_13211,N_13179);
xnor U13322 (N_13322,N_13137,N_13155);
nor U13323 (N_13323,N_13237,N_13141);
or U13324 (N_13324,N_13160,N_13183);
xnor U13325 (N_13325,N_13157,N_13164);
nand U13326 (N_13326,N_13200,N_13151);
nor U13327 (N_13327,N_13215,N_13131);
nor U13328 (N_13328,N_13158,N_13212);
xor U13329 (N_13329,N_13134,N_13226);
or U13330 (N_13330,N_13214,N_13216);
nor U13331 (N_13331,N_13148,N_13182);
xnor U13332 (N_13332,N_13141,N_13168);
and U13333 (N_13333,N_13151,N_13131);
xor U13334 (N_13334,N_13136,N_13131);
nand U13335 (N_13335,N_13208,N_13150);
xor U13336 (N_13336,N_13209,N_13149);
or U13337 (N_13337,N_13240,N_13173);
xnor U13338 (N_13338,N_13208,N_13157);
nand U13339 (N_13339,N_13142,N_13230);
nand U13340 (N_13340,N_13206,N_13215);
and U13341 (N_13341,N_13137,N_13179);
nand U13342 (N_13342,N_13154,N_13240);
and U13343 (N_13343,N_13223,N_13135);
nand U13344 (N_13344,N_13163,N_13246);
xor U13345 (N_13345,N_13192,N_13223);
nor U13346 (N_13346,N_13135,N_13178);
and U13347 (N_13347,N_13242,N_13182);
nor U13348 (N_13348,N_13165,N_13203);
nand U13349 (N_13349,N_13203,N_13138);
nor U13350 (N_13350,N_13187,N_13243);
nand U13351 (N_13351,N_13230,N_13166);
xnor U13352 (N_13352,N_13205,N_13234);
xnor U13353 (N_13353,N_13134,N_13193);
xor U13354 (N_13354,N_13154,N_13179);
and U13355 (N_13355,N_13175,N_13169);
nand U13356 (N_13356,N_13132,N_13137);
nor U13357 (N_13357,N_13205,N_13199);
or U13358 (N_13358,N_13221,N_13229);
nor U13359 (N_13359,N_13215,N_13227);
and U13360 (N_13360,N_13230,N_13176);
nor U13361 (N_13361,N_13202,N_13128);
nand U13362 (N_13362,N_13229,N_13138);
or U13363 (N_13363,N_13150,N_13201);
xnor U13364 (N_13364,N_13238,N_13148);
or U13365 (N_13365,N_13179,N_13146);
nand U13366 (N_13366,N_13188,N_13131);
xnor U13367 (N_13367,N_13126,N_13211);
and U13368 (N_13368,N_13222,N_13152);
or U13369 (N_13369,N_13152,N_13133);
or U13370 (N_13370,N_13159,N_13138);
or U13371 (N_13371,N_13167,N_13180);
or U13372 (N_13372,N_13192,N_13189);
or U13373 (N_13373,N_13208,N_13234);
nand U13374 (N_13374,N_13144,N_13160);
xnor U13375 (N_13375,N_13354,N_13312);
nor U13376 (N_13376,N_13257,N_13347);
or U13377 (N_13377,N_13309,N_13284);
nor U13378 (N_13378,N_13315,N_13343);
or U13379 (N_13379,N_13294,N_13271);
nor U13380 (N_13380,N_13368,N_13254);
nand U13381 (N_13381,N_13326,N_13251);
and U13382 (N_13382,N_13258,N_13338);
nor U13383 (N_13383,N_13275,N_13336);
nor U13384 (N_13384,N_13290,N_13255);
xnor U13385 (N_13385,N_13277,N_13263);
nand U13386 (N_13386,N_13373,N_13328);
xor U13387 (N_13387,N_13367,N_13289);
or U13388 (N_13388,N_13305,N_13352);
and U13389 (N_13389,N_13359,N_13298);
xor U13390 (N_13390,N_13331,N_13340);
nand U13391 (N_13391,N_13348,N_13295);
xor U13392 (N_13392,N_13316,N_13268);
or U13393 (N_13393,N_13288,N_13319);
nand U13394 (N_13394,N_13308,N_13310);
nand U13395 (N_13395,N_13318,N_13353);
and U13396 (N_13396,N_13317,N_13270);
and U13397 (N_13397,N_13302,N_13321);
nor U13398 (N_13398,N_13286,N_13269);
or U13399 (N_13399,N_13346,N_13283);
and U13400 (N_13400,N_13370,N_13260);
or U13401 (N_13401,N_13363,N_13306);
and U13402 (N_13402,N_13278,N_13362);
or U13403 (N_13403,N_13261,N_13337);
nor U13404 (N_13404,N_13274,N_13273);
nand U13405 (N_13405,N_13372,N_13279);
xor U13406 (N_13406,N_13323,N_13272);
nand U13407 (N_13407,N_13369,N_13314);
or U13408 (N_13408,N_13360,N_13335);
xnor U13409 (N_13409,N_13262,N_13253);
nor U13410 (N_13410,N_13324,N_13357);
nor U13411 (N_13411,N_13264,N_13265);
xor U13412 (N_13412,N_13355,N_13320);
nor U13413 (N_13413,N_13332,N_13329);
and U13414 (N_13414,N_13304,N_13311);
nor U13415 (N_13415,N_13322,N_13349);
nand U13416 (N_13416,N_13361,N_13344);
nor U13417 (N_13417,N_13350,N_13291);
nand U13418 (N_13418,N_13281,N_13333);
nand U13419 (N_13419,N_13292,N_13280);
or U13420 (N_13420,N_13296,N_13299);
nand U13421 (N_13421,N_13259,N_13351);
xnor U13422 (N_13422,N_13293,N_13313);
nor U13423 (N_13423,N_13339,N_13342);
nor U13424 (N_13424,N_13256,N_13356);
and U13425 (N_13425,N_13325,N_13364);
nand U13426 (N_13426,N_13341,N_13301);
and U13427 (N_13427,N_13266,N_13297);
xnor U13428 (N_13428,N_13303,N_13358);
nor U13429 (N_13429,N_13330,N_13371);
nand U13430 (N_13430,N_13345,N_13307);
nand U13431 (N_13431,N_13334,N_13252);
or U13432 (N_13432,N_13276,N_13365);
and U13433 (N_13433,N_13300,N_13250);
xnor U13434 (N_13434,N_13366,N_13267);
nor U13435 (N_13435,N_13374,N_13282);
or U13436 (N_13436,N_13287,N_13285);
nor U13437 (N_13437,N_13327,N_13349);
and U13438 (N_13438,N_13263,N_13352);
nor U13439 (N_13439,N_13372,N_13273);
nand U13440 (N_13440,N_13276,N_13350);
xor U13441 (N_13441,N_13327,N_13284);
and U13442 (N_13442,N_13290,N_13362);
nor U13443 (N_13443,N_13332,N_13361);
or U13444 (N_13444,N_13262,N_13353);
nand U13445 (N_13445,N_13363,N_13366);
xnor U13446 (N_13446,N_13287,N_13272);
xor U13447 (N_13447,N_13351,N_13287);
nor U13448 (N_13448,N_13315,N_13373);
nand U13449 (N_13449,N_13309,N_13300);
nor U13450 (N_13450,N_13294,N_13274);
and U13451 (N_13451,N_13295,N_13277);
and U13452 (N_13452,N_13321,N_13331);
xor U13453 (N_13453,N_13300,N_13257);
xor U13454 (N_13454,N_13266,N_13271);
nor U13455 (N_13455,N_13296,N_13292);
and U13456 (N_13456,N_13296,N_13291);
and U13457 (N_13457,N_13320,N_13316);
nand U13458 (N_13458,N_13281,N_13346);
or U13459 (N_13459,N_13292,N_13328);
nor U13460 (N_13460,N_13362,N_13269);
xor U13461 (N_13461,N_13274,N_13285);
nor U13462 (N_13462,N_13268,N_13319);
or U13463 (N_13463,N_13303,N_13265);
nor U13464 (N_13464,N_13363,N_13360);
or U13465 (N_13465,N_13265,N_13327);
and U13466 (N_13466,N_13294,N_13267);
or U13467 (N_13467,N_13335,N_13346);
or U13468 (N_13468,N_13296,N_13285);
nor U13469 (N_13469,N_13264,N_13308);
and U13470 (N_13470,N_13370,N_13278);
xnor U13471 (N_13471,N_13370,N_13345);
or U13472 (N_13472,N_13263,N_13367);
and U13473 (N_13473,N_13284,N_13261);
or U13474 (N_13474,N_13258,N_13269);
and U13475 (N_13475,N_13278,N_13343);
or U13476 (N_13476,N_13285,N_13351);
nand U13477 (N_13477,N_13336,N_13265);
or U13478 (N_13478,N_13355,N_13257);
or U13479 (N_13479,N_13371,N_13270);
nor U13480 (N_13480,N_13281,N_13342);
and U13481 (N_13481,N_13358,N_13319);
xor U13482 (N_13482,N_13331,N_13301);
xnor U13483 (N_13483,N_13258,N_13286);
xnor U13484 (N_13484,N_13309,N_13335);
or U13485 (N_13485,N_13298,N_13266);
nand U13486 (N_13486,N_13302,N_13251);
nor U13487 (N_13487,N_13373,N_13285);
xor U13488 (N_13488,N_13262,N_13292);
xor U13489 (N_13489,N_13348,N_13265);
or U13490 (N_13490,N_13328,N_13285);
and U13491 (N_13491,N_13333,N_13352);
or U13492 (N_13492,N_13323,N_13274);
or U13493 (N_13493,N_13257,N_13374);
xnor U13494 (N_13494,N_13283,N_13352);
or U13495 (N_13495,N_13295,N_13290);
or U13496 (N_13496,N_13311,N_13275);
xnor U13497 (N_13497,N_13333,N_13339);
xor U13498 (N_13498,N_13271,N_13262);
xor U13499 (N_13499,N_13284,N_13267);
xnor U13500 (N_13500,N_13468,N_13442);
or U13501 (N_13501,N_13400,N_13377);
nand U13502 (N_13502,N_13436,N_13376);
and U13503 (N_13503,N_13453,N_13391);
nor U13504 (N_13504,N_13483,N_13439);
or U13505 (N_13505,N_13454,N_13497);
or U13506 (N_13506,N_13437,N_13462);
xnor U13507 (N_13507,N_13478,N_13499);
xnor U13508 (N_13508,N_13484,N_13491);
xnor U13509 (N_13509,N_13445,N_13395);
xnor U13510 (N_13510,N_13429,N_13455);
nand U13511 (N_13511,N_13496,N_13414);
nor U13512 (N_13512,N_13413,N_13404);
nor U13513 (N_13513,N_13440,N_13427);
nand U13514 (N_13514,N_13379,N_13441);
and U13515 (N_13515,N_13443,N_13435);
or U13516 (N_13516,N_13412,N_13488);
and U13517 (N_13517,N_13428,N_13493);
nor U13518 (N_13518,N_13424,N_13457);
xor U13519 (N_13519,N_13482,N_13464);
nor U13520 (N_13520,N_13422,N_13420);
nand U13521 (N_13521,N_13382,N_13430);
or U13522 (N_13522,N_13438,N_13381);
or U13523 (N_13523,N_13444,N_13383);
nand U13524 (N_13524,N_13397,N_13388);
or U13525 (N_13525,N_13416,N_13418);
xnor U13526 (N_13526,N_13449,N_13474);
nor U13527 (N_13527,N_13476,N_13450);
nand U13528 (N_13528,N_13398,N_13481);
xor U13529 (N_13529,N_13495,N_13434);
nand U13530 (N_13530,N_13385,N_13380);
nand U13531 (N_13531,N_13456,N_13394);
nand U13532 (N_13532,N_13415,N_13465);
nor U13533 (N_13533,N_13460,N_13426);
xor U13534 (N_13534,N_13410,N_13469);
xor U13535 (N_13535,N_13399,N_13378);
nand U13536 (N_13536,N_13390,N_13473);
and U13537 (N_13537,N_13492,N_13490);
nor U13538 (N_13538,N_13433,N_13423);
or U13539 (N_13539,N_13451,N_13396);
nand U13540 (N_13540,N_13421,N_13461);
nor U13541 (N_13541,N_13479,N_13386);
or U13542 (N_13542,N_13419,N_13459);
xor U13543 (N_13543,N_13480,N_13466);
xnor U13544 (N_13544,N_13485,N_13417);
and U13545 (N_13545,N_13463,N_13432);
xnor U13546 (N_13546,N_13402,N_13494);
xnor U13547 (N_13547,N_13467,N_13477);
nor U13548 (N_13548,N_13408,N_13431);
nor U13549 (N_13549,N_13403,N_13486);
and U13550 (N_13550,N_13471,N_13389);
nor U13551 (N_13551,N_13392,N_13487);
xnor U13552 (N_13552,N_13425,N_13401);
or U13553 (N_13553,N_13452,N_13406);
nand U13554 (N_13554,N_13375,N_13475);
and U13555 (N_13555,N_13407,N_13446);
or U13556 (N_13556,N_13393,N_13458);
or U13557 (N_13557,N_13387,N_13470);
nor U13558 (N_13558,N_13411,N_13489);
nand U13559 (N_13559,N_13384,N_13498);
xnor U13560 (N_13560,N_13409,N_13472);
xnor U13561 (N_13561,N_13448,N_13447);
xnor U13562 (N_13562,N_13405,N_13489);
nor U13563 (N_13563,N_13407,N_13415);
or U13564 (N_13564,N_13463,N_13405);
or U13565 (N_13565,N_13412,N_13446);
and U13566 (N_13566,N_13418,N_13382);
nand U13567 (N_13567,N_13442,N_13477);
or U13568 (N_13568,N_13455,N_13441);
or U13569 (N_13569,N_13486,N_13412);
and U13570 (N_13570,N_13498,N_13425);
nand U13571 (N_13571,N_13499,N_13498);
and U13572 (N_13572,N_13408,N_13468);
or U13573 (N_13573,N_13438,N_13379);
nor U13574 (N_13574,N_13395,N_13387);
or U13575 (N_13575,N_13470,N_13479);
nand U13576 (N_13576,N_13459,N_13436);
and U13577 (N_13577,N_13484,N_13470);
and U13578 (N_13578,N_13480,N_13462);
nand U13579 (N_13579,N_13446,N_13408);
and U13580 (N_13580,N_13468,N_13495);
nor U13581 (N_13581,N_13389,N_13376);
xnor U13582 (N_13582,N_13434,N_13411);
xnor U13583 (N_13583,N_13414,N_13419);
xor U13584 (N_13584,N_13382,N_13435);
and U13585 (N_13585,N_13377,N_13435);
nand U13586 (N_13586,N_13429,N_13424);
nor U13587 (N_13587,N_13491,N_13455);
nand U13588 (N_13588,N_13375,N_13389);
or U13589 (N_13589,N_13449,N_13454);
nand U13590 (N_13590,N_13423,N_13484);
xor U13591 (N_13591,N_13467,N_13490);
nand U13592 (N_13592,N_13450,N_13465);
and U13593 (N_13593,N_13413,N_13466);
or U13594 (N_13594,N_13393,N_13494);
or U13595 (N_13595,N_13407,N_13426);
nand U13596 (N_13596,N_13407,N_13455);
nor U13597 (N_13597,N_13491,N_13475);
and U13598 (N_13598,N_13420,N_13407);
xor U13599 (N_13599,N_13470,N_13432);
xnor U13600 (N_13600,N_13435,N_13412);
nor U13601 (N_13601,N_13430,N_13400);
or U13602 (N_13602,N_13468,N_13425);
xnor U13603 (N_13603,N_13483,N_13495);
nand U13604 (N_13604,N_13459,N_13456);
nand U13605 (N_13605,N_13485,N_13474);
nor U13606 (N_13606,N_13479,N_13408);
xnor U13607 (N_13607,N_13381,N_13449);
nand U13608 (N_13608,N_13385,N_13413);
and U13609 (N_13609,N_13425,N_13460);
xor U13610 (N_13610,N_13388,N_13464);
or U13611 (N_13611,N_13425,N_13442);
and U13612 (N_13612,N_13404,N_13473);
nand U13613 (N_13613,N_13442,N_13393);
nor U13614 (N_13614,N_13415,N_13437);
and U13615 (N_13615,N_13378,N_13389);
or U13616 (N_13616,N_13411,N_13419);
and U13617 (N_13617,N_13477,N_13488);
nor U13618 (N_13618,N_13443,N_13477);
nand U13619 (N_13619,N_13377,N_13382);
nor U13620 (N_13620,N_13457,N_13390);
and U13621 (N_13621,N_13435,N_13440);
xor U13622 (N_13622,N_13376,N_13424);
xnor U13623 (N_13623,N_13435,N_13375);
or U13624 (N_13624,N_13485,N_13486);
or U13625 (N_13625,N_13526,N_13518);
nor U13626 (N_13626,N_13568,N_13549);
nor U13627 (N_13627,N_13555,N_13573);
xor U13628 (N_13628,N_13514,N_13624);
or U13629 (N_13629,N_13543,N_13547);
xor U13630 (N_13630,N_13561,N_13579);
nand U13631 (N_13631,N_13591,N_13502);
nor U13632 (N_13632,N_13595,N_13509);
xnor U13633 (N_13633,N_13607,N_13545);
nand U13634 (N_13634,N_13531,N_13505);
nand U13635 (N_13635,N_13539,N_13521);
nand U13636 (N_13636,N_13524,N_13522);
nor U13637 (N_13637,N_13558,N_13528);
or U13638 (N_13638,N_13551,N_13608);
or U13639 (N_13639,N_13620,N_13615);
or U13640 (N_13640,N_13546,N_13616);
and U13641 (N_13641,N_13604,N_13541);
nor U13642 (N_13642,N_13556,N_13504);
nor U13643 (N_13643,N_13581,N_13576);
and U13644 (N_13644,N_13596,N_13592);
nor U13645 (N_13645,N_13507,N_13577);
or U13646 (N_13646,N_13605,N_13602);
or U13647 (N_13647,N_13584,N_13618);
and U13648 (N_13648,N_13617,N_13571);
and U13649 (N_13649,N_13588,N_13530);
nand U13650 (N_13650,N_13525,N_13613);
xnor U13651 (N_13651,N_13523,N_13560);
nor U13652 (N_13652,N_13550,N_13567);
nor U13653 (N_13653,N_13508,N_13621);
or U13654 (N_13654,N_13601,N_13544);
or U13655 (N_13655,N_13597,N_13611);
and U13656 (N_13656,N_13610,N_13506);
and U13657 (N_13657,N_13553,N_13619);
xor U13658 (N_13658,N_13540,N_13519);
nand U13659 (N_13659,N_13520,N_13580);
nor U13660 (N_13660,N_13554,N_13578);
nand U13661 (N_13661,N_13532,N_13527);
nand U13662 (N_13662,N_13537,N_13623);
nor U13663 (N_13663,N_13622,N_13538);
nor U13664 (N_13664,N_13582,N_13515);
nor U13665 (N_13665,N_13565,N_13587);
nand U13666 (N_13666,N_13594,N_13563);
nor U13667 (N_13667,N_13533,N_13590);
nand U13668 (N_13668,N_13542,N_13535);
nand U13669 (N_13669,N_13599,N_13572);
or U13670 (N_13670,N_13552,N_13516);
nor U13671 (N_13671,N_13562,N_13570);
nand U13672 (N_13672,N_13585,N_13557);
or U13673 (N_13673,N_13598,N_13501);
nor U13674 (N_13674,N_13600,N_13574);
nand U13675 (N_13675,N_13583,N_13529);
or U13676 (N_13676,N_13512,N_13536);
nand U13677 (N_13677,N_13559,N_13534);
xnor U13678 (N_13678,N_13564,N_13603);
nand U13679 (N_13679,N_13548,N_13609);
and U13680 (N_13680,N_13569,N_13614);
xnor U13681 (N_13681,N_13500,N_13606);
or U13682 (N_13682,N_13517,N_13513);
xnor U13683 (N_13683,N_13510,N_13503);
nand U13684 (N_13684,N_13612,N_13589);
or U13685 (N_13685,N_13575,N_13586);
xnor U13686 (N_13686,N_13511,N_13566);
or U13687 (N_13687,N_13593,N_13597);
xnor U13688 (N_13688,N_13577,N_13530);
nand U13689 (N_13689,N_13550,N_13616);
nand U13690 (N_13690,N_13534,N_13518);
nor U13691 (N_13691,N_13616,N_13620);
nand U13692 (N_13692,N_13581,N_13574);
nor U13693 (N_13693,N_13519,N_13501);
nor U13694 (N_13694,N_13542,N_13528);
or U13695 (N_13695,N_13547,N_13562);
and U13696 (N_13696,N_13600,N_13597);
xor U13697 (N_13697,N_13565,N_13622);
or U13698 (N_13698,N_13594,N_13551);
nand U13699 (N_13699,N_13599,N_13541);
nand U13700 (N_13700,N_13524,N_13601);
or U13701 (N_13701,N_13542,N_13579);
xor U13702 (N_13702,N_13526,N_13536);
nand U13703 (N_13703,N_13621,N_13525);
nand U13704 (N_13704,N_13549,N_13620);
or U13705 (N_13705,N_13537,N_13566);
nand U13706 (N_13706,N_13513,N_13567);
nand U13707 (N_13707,N_13526,N_13562);
and U13708 (N_13708,N_13597,N_13621);
xor U13709 (N_13709,N_13557,N_13526);
nor U13710 (N_13710,N_13602,N_13623);
nor U13711 (N_13711,N_13519,N_13570);
nand U13712 (N_13712,N_13614,N_13537);
nor U13713 (N_13713,N_13617,N_13619);
xor U13714 (N_13714,N_13611,N_13563);
nor U13715 (N_13715,N_13623,N_13544);
xnor U13716 (N_13716,N_13595,N_13608);
nor U13717 (N_13717,N_13530,N_13595);
nand U13718 (N_13718,N_13562,N_13587);
xnor U13719 (N_13719,N_13602,N_13622);
nand U13720 (N_13720,N_13527,N_13559);
nor U13721 (N_13721,N_13571,N_13594);
and U13722 (N_13722,N_13514,N_13566);
nand U13723 (N_13723,N_13546,N_13561);
or U13724 (N_13724,N_13533,N_13624);
xor U13725 (N_13725,N_13565,N_13522);
nand U13726 (N_13726,N_13504,N_13533);
xor U13727 (N_13727,N_13557,N_13618);
and U13728 (N_13728,N_13513,N_13518);
or U13729 (N_13729,N_13507,N_13553);
and U13730 (N_13730,N_13559,N_13513);
nor U13731 (N_13731,N_13521,N_13616);
and U13732 (N_13732,N_13526,N_13560);
nand U13733 (N_13733,N_13556,N_13536);
nand U13734 (N_13734,N_13540,N_13612);
or U13735 (N_13735,N_13591,N_13603);
nand U13736 (N_13736,N_13611,N_13512);
xnor U13737 (N_13737,N_13502,N_13603);
nand U13738 (N_13738,N_13555,N_13543);
nor U13739 (N_13739,N_13561,N_13611);
or U13740 (N_13740,N_13563,N_13613);
xor U13741 (N_13741,N_13515,N_13616);
and U13742 (N_13742,N_13542,N_13530);
or U13743 (N_13743,N_13526,N_13524);
or U13744 (N_13744,N_13508,N_13588);
nor U13745 (N_13745,N_13548,N_13558);
and U13746 (N_13746,N_13535,N_13579);
nor U13747 (N_13747,N_13550,N_13613);
and U13748 (N_13748,N_13521,N_13514);
or U13749 (N_13749,N_13504,N_13550);
nor U13750 (N_13750,N_13657,N_13655);
and U13751 (N_13751,N_13737,N_13629);
xnor U13752 (N_13752,N_13656,N_13627);
or U13753 (N_13753,N_13680,N_13700);
and U13754 (N_13754,N_13745,N_13689);
xor U13755 (N_13755,N_13631,N_13742);
nor U13756 (N_13756,N_13632,N_13638);
or U13757 (N_13757,N_13626,N_13625);
nand U13758 (N_13758,N_13723,N_13714);
nor U13759 (N_13759,N_13715,N_13729);
and U13760 (N_13760,N_13706,N_13674);
and U13761 (N_13761,N_13675,N_13672);
nor U13762 (N_13762,N_13707,N_13720);
or U13763 (N_13763,N_13712,N_13730);
or U13764 (N_13764,N_13662,N_13660);
nor U13765 (N_13765,N_13630,N_13667);
nand U13766 (N_13766,N_13713,N_13710);
nand U13767 (N_13767,N_13646,N_13684);
nand U13768 (N_13768,N_13643,N_13698);
or U13769 (N_13769,N_13702,N_13735);
xor U13770 (N_13770,N_13708,N_13651);
nand U13771 (N_13771,N_13695,N_13633);
xor U13772 (N_13772,N_13724,N_13733);
nor U13773 (N_13773,N_13736,N_13716);
nand U13774 (N_13774,N_13658,N_13652);
and U13775 (N_13775,N_13699,N_13678);
or U13776 (N_13776,N_13640,N_13649);
or U13777 (N_13777,N_13683,N_13670);
and U13778 (N_13778,N_13725,N_13746);
and U13779 (N_13779,N_13642,N_13682);
and U13780 (N_13780,N_13749,N_13728);
nand U13781 (N_13781,N_13653,N_13732);
xnor U13782 (N_13782,N_13691,N_13721);
or U13783 (N_13783,N_13748,N_13692);
and U13784 (N_13784,N_13666,N_13644);
or U13785 (N_13785,N_13654,N_13681);
and U13786 (N_13786,N_13696,N_13731);
nor U13787 (N_13787,N_13687,N_13726);
xor U13788 (N_13788,N_13701,N_13694);
and U13789 (N_13789,N_13676,N_13739);
and U13790 (N_13790,N_13717,N_13677);
and U13791 (N_13791,N_13645,N_13690);
nand U13792 (N_13792,N_13711,N_13740);
nand U13793 (N_13793,N_13636,N_13668);
xnor U13794 (N_13794,N_13704,N_13635);
nor U13795 (N_13795,N_13628,N_13639);
or U13796 (N_13796,N_13705,N_13718);
nor U13797 (N_13797,N_13673,N_13741);
nor U13798 (N_13798,N_13679,N_13719);
and U13799 (N_13799,N_13663,N_13669);
and U13800 (N_13800,N_13665,N_13685);
and U13801 (N_13801,N_13709,N_13661);
nor U13802 (N_13802,N_13650,N_13722);
xnor U13803 (N_13803,N_13738,N_13734);
nor U13804 (N_13804,N_13671,N_13641);
xnor U13805 (N_13805,N_13659,N_13703);
nor U13806 (N_13806,N_13743,N_13697);
nor U13807 (N_13807,N_13637,N_13686);
xor U13808 (N_13808,N_13647,N_13727);
nor U13809 (N_13809,N_13747,N_13744);
and U13810 (N_13810,N_13664,N_13688);
and U13811 (N_13811,N_13648,N_13693);
nand U13812 (N_13812,N_13634,N_13739);
nand U13813 (N_13813,N_13650,N_13645);
xor U13814 (N_13814,N_13662,N_13627);
and U13815 (N_13815,N_13640,N_13667);
nand U13816 (N_13816,N_13627,N_13658);
xnor U13817 (N_13817,N_13697,N_13656);
and U13818 (N_13818,N_13737,N_13736);
or U13819 (N_13819,N_13689,N_13733);
or U13820 (N_13820,N_13735,N_13627);
nor U13821 (N_13821,N_13709,N_13676);
and U13822 (N_13822,N_13633,N_13641);
xor U13823 (N_13823,N_13707,N_13695);
xor U13824 (N_13824,N_13649,N_13705);
nor U13825 (N_13825,N_13655,N_13642);
and U13826 (N_13826,N_13702,N_13717);
nor U13827 (N_13827,N_13657,N_13682);
or U13828 (N_13828,N_13718,N_13723);
nor U13829 (N_13829,N_13638,N_13658);
nor U13830 (N_13830,N_13634,N_13745);
or U13831 (N_13831,N_13627,N_13638);
xnor U13832 (N_13832,N_13741,N_13732);
nand U13833 (N_13833,N_13680,N_13657);
xor U13834 (N_13834,N_13644,N_13686);
xnor U13835 (N_13835,N_13659,N_13725);
nor U13836 (N_13836,N_13688,N_13685);
nor U13837 (N_13837,N_13630,N_13745);
or U13838 (N_13838,N_13685,N_13638);
nand U13839 (N_13839,N_13719,N_13746);
nand U13840 (N_13840,N_13642,N_13720);
nand U13841 (N_13841,N_13732,N_13711);
nor U13842 (N_13842,N_13649,N_13716);
or U13843 (N_13843,N_13625,N_13686);
and U13844 (N_13844,N_13719,N_13744);
nand U13845 (N_13845,N_13691,N_13742);
nand U13846 (N_13846,N_13723,N_13686);
or U13847 (N_13847,N_13636,N_13731);
xnor U13848 (N_13848,N_13704,N_13689);
nor U13849 (N_13849,N_13741,N_13716);
and U13850 (N_13850,N_13724,N_13662);
nor U13851 (N_13851,N_13641,N_13730);
nand U13852 (N_13852,N_13633,N_13652);
xnor U13853 (N_13853,N_13690,N_13633);
nand U13854 (N_13854,N_13648,N_13681);
or U13855 (N_13855,N_13712,N_13685);
nand U13856 (N_13856,N_13662,N_13705);
xor U13857 (N_13857,N_13745,N_13695);
and U13858 (N_13858,N_13721,N_13660);
nor U13859 (N_13859,N_13720,N_13659);
nand U13860 (N_13860,N_13718,N_13714);
or U13861 (N_13861,N_13682,N_13629);
or U13862 (N_13862,N_13744,N_13656);
xor U13863 (N_13863,N_13680,N_13654);
nand U13864 (N_13864,N_13657,N_13689);
or U13865 (N_13865,N_13697,N_13667);
xor U13866 (N_13866,N_13638,N_13635);
and U13867 (N_13867,N_13699,N_13649);
xor U13868 (N_13868,N_13678,N_13740);
and U13869 (N_13869,N_13647,N_13639);
xor U13870 (N_13870,N_13710,N_13734);
nor U13871 (N_13871,N_13746,N_13633);
or U13872 (N_13872,N_13712,N_13656);
nand U13873 (N_13873,N_13719,N_13637);
nor U13874 (N_13874,N_13661,N_13649);
nand U13875 (N_13875,N_13755,N_13826);
nand U13876 (N_13876,N_13822,N_13770);
or U13877 (N_13877,N_13771,N_13868);
nand U13878 (N_13878,N_13779,N_13758);
and U13879 (N_13879,N_13842,N_13843);
nor U13880 (N_13880,N_13812,N_13848);
nor U13881 (N_13881,N_13844,N_13780);
and U13882 (N_13882,N_13807,N_13814);
or U13883 (N_13883,N_13782,N_13831);
nor U13884 (N_13884,N_13870,N_13792);
nor U13885 (N_13885,N_13841,N_13793);
nand U13886 (N_13886,N_13796,N_13799);
xor U13887 (N_13887,N_13804,N_13836);
or U13888 (N_13888,N_13762,N_13845);
and U13889 (N_13889,N_13830,N_13821);
and U13890 (N_13890,N_13819,N_13853);
nand U13891 (N_13891,N_13835,N_13858);
nor U13892 (N_13892,N_13787,N_13874);
nand U13893 (N_13893,N_13851,N_13873);
nor U13894 (N_13894,N_13774,N_13777);
nor U13895 (N_13895,N_13808,N_13862);
nand U13896 (N_13896,N_13863,N_13794);
nand U13897 (N_13897,N_13817,N_13764);
and U13898 (N_13898,N_13806,N_13856);
and U13899 (N_13899,N_13776,N_13813);
and U13900 (N_13900,N_13761,N_13784);
or U13901 (N_13901,N_13781,N_13800);
xor U13902 (N_13902,N_13810,N_13785);
xor U13903 (N_13903,N_13765,N_13865);
nor U13904 (N_13904,N_13798,N_13839);
and U13905 (N_13905,N_13791,N_13789);
nor U13906 (N_13906,N_13786,N_13820);
xnor U13907 (N_13907,N_13852,N_13763);
or U13908 (N_13908,N_13759,N_13827);
or U13909 (N_13909,N_13861,N_13802);
nand U13910 (N_13910,N_13754,N_13767);
nand U13911 (N_13911,N_13867,N_13797);
nand U13912 (N_13912,N_13773,N_13816);
or U13913 (N_13913,N_13859,N_13857);
xnor U13914 (N_13914,N_13869,N_13772);
nand U13915 (N_13915,N_13757,N_13750);
nor U13916 (N_13916,N_13871,N_13854);
and U13917 (N_13917,N_13850,N_13849);
nor U13918 (N_13918,N_13795,N_13855);
nor U13919 (N_13919,N_13756,N_13809);
xor U13920 (N_13920,N_13824,N_13846);
xor U13921 (N_13921,N_13790,N_13752);
or U13922 (N_13922,N_13837,N_13828);
nor U13923 (N_13923,N_13825,N_13753);
nand U13924 (N_13924,N_13872,N_13788);
xnor U13925 (N_13925,N_13803,N_13864);
xnor U13926 (N_13926,N_13818,N_13829);
or U13927 (N_13927,N_13834,N_13805);
nand U13928 (N_13928,N_13833,N_13838);
nand U13929 (N_13929,N_13801,N_13847);
or U13930 (N_13930,N_13760,N_13823);
xor U13931 (N_13931,N_13811,N_13840);
xnor U13932 (N_13932,N_13815,N_13768);
nand U13933 (N_13933,N_13769,N_13775);
xnor U13934 (N_13934,N_13766,N_13866);
or U13935 (N_13935,N_13860,N_13751);
nand U13936 (N_13936,N_13783,N_13778);
or U13937 (N_13937,N_13832,N_13822);
and U13938 (N_13938,N_13858,N_13869);
nand U13939 (N_13939,N_13840,N_13820);
xnor U13940 (N_13940,N_13823,N_13839);
nand U13941 (N_13941,N_13799,N_13765);
nor U13942 (N_13942,N_13845,N_13763);
nor U13943 (N_13943,N_13768,N_13769);
nor U13944 (N_13944,N_13862,N_13822);
or U13945 (N_13945,N_13845,N_13829);
nand U13946 (N_13946,N_13804,N_13798);
and U13947 (N_13947,N_13811,N_13750);
or U13948 (N_13948,N_13816,N_13775);
or U13949 (N_13949,N_13804,N_13753);
or U13950 (N_13950,N_13818,N_13824);
nor U13951 (N_13951,N_13824,N_13814);
nor U13952 (N_13952,N_13803,N_13872);
and U13953 (N_13953,N_13843,N_13795);
nand U13954 (N_13954,N_13859,N_13754);
xnor U13955 (N_13955,N_13768,N_13868);
and U13956 (N_13956,N_13827,N_13780);
or U13957 (N_13957,N_13783,N_13864);
or U13958 (N_13958,N_13771,N_13801);
nor U13959 (N_13959,N_13765,N_13863);
and U13960 (N_13960,N_13839,N_13830);
and U13961 (N_13961,N_13765,N_13869);
and U13962 (N_13962,N_13794,N_13781);
nand U13963 (N_13963,N_13830,N_13808);
and U13964 (N_13964,N_13826,N_13775);
nor U13965 (N_13965,N_13837,N_13846);
or U13966 (N_13966,N_13815,N_13764);
xnor U13967 (N_13967,N_13827,N_13870);
or U13968 (N_13968,N_13792,N_13763);
and U13969 (N_13969,N_13827,N_13812);
or U13970 (N_13970,N_13859,N_13871);
nand U13971 (N_13971,N_13765,N_13809);
nor U13972 (N_13972,N_13812,N_13757);
xor U13973 (N_13973,N_13863,N_13807);
or U13974 (N_13974,N_13804,N_13873);
nor U13975 (N_13975,N_13760,N_13836);
nor U13976 (N_13976,N_13760,N_13831);
or U13977 (N_13977,N_13778,N_13857);
nor U13978 (N_13978,N_13818,N_13845);
nor U13979 (N_13979,N_13820,N_13808);
nand U13980 (N_13980,N_13828,N_13812);
nor U13981 (N_13981,N_13836,N_13861);
and U13982 (N_13982,N_13848,N_13754);
nor U13983 (N_13983,N_13781,N_13817);
nand U13984 (N_13984,N_13868,N_13804);
or U13985 (N_13985,N_13853,N_13755);
and U13986 (N_13986,N_13842,N_13765);
xnor U13987 (N_13987,N_13775,N_13864);
and U13988 (N_13988,N_13819,N_13866);
or U13989 (N_13989,N_13840,N_13823);
xnor U13990 (N_13990,N_13783,N_13832);
or U13991 (N_13991,N_13794,N_13864);
xnor U13992 (N_13992,N_13864,N_13840);
xnor U13993 (N_13993,N_13817,N_13793);
nand U13994 (N_13994,N_13775,N_13807);
nand U13995 (N_13995,N_13818,N_13756);
nor U13996 (N_13996,N_13780,N_13812);
or U13997 (N_13997,N_13787,N_13785);
and U13998 (N_13998,N_13826,N_13821);
or U13999 (N_13999,N_13820,N_13799);
nor U14000 (N_14000,N_13919,N_13996);
nor U14001 (N_14001,N_13988,N_13924);
xor U14002 (N_14002,N_13977,N_13952);
xnor U14003 (N_14003,N_13997,N_13940);
or U14004 (N_14004,N_13968,N_13958);
nand U14005 (N_14005,N_13884,N_13910);
xnor U14006 (N_14006,N_13932,N_13999);
nand U14007 (N_14007,N_13975,N_13893);
nor U14008 (N_14008,N_13913,N_13907);
nor U14009 (N_14009,N_13939,N_13905);
nand U14010 (N_14010,N_13938,N_13898);
and U14011 (N_14011,N_13935,N_13887);
nand U14012 (N_14012,N_13894,N_13993);
and U14013 (N_14013,N_13895,N_13899);
nand U14014 (N_14014,N_13920,N_13953);
and U14015 (N_14015,N_13954,N_13971);
nand U14016 (N_14016,N_13908,N_13880);
nand U14017 (N_14017,N_13959,N_13950);
or U14018 (N_14018,N_13883,N_13890);
and U14019 (N_14019,N_13973,N_13921);
nand U14020 (N_14020,N_13897,N_13981);
xor U14021 (N_14021,N_13942,N_13900);
or U14022 (N_14022,N_13889,N_13989);
nor U14023 (N_14023,N_13927,N_13955);
xnor U14024 (N_14024,N_13946,N_13928);
and U14025 (N_14025,N_13960,N_13912);
nand U14026 (N_14026,N_13964,N_13943);
nor U14027 (N_14027,N_13976,N_13987);
nand U14028 (N_14028,N_13965,N_13985);
nor U14029 (N_14029,N_13998,N_13882);
nor U14030 (N_14030,N_13923,N_13881);
nand U14031 (N_14031,N_13949,N_13945);
and U14032 (N_14032,N_13896,N_13931);
nand U14033 (N_14033,N_13937,N_13947);
xor U14034 (N_14034,N_13994,N_13948);
and U14035 (N_14035,N_13962,N_13915);
and U14036 (N_14036,N_13929,N_13986);
xor U14037 (N_14037,N_13925,N_13875);
xnor U14038 (N_14038,N_13877,N_13970);
xor U14039 (N_14039,N_13992,N_13933);
nand U14040 (N_14040,N_13982,N_13990);
and U14041 (N_14041,N_13906,N_13979);
xor U14042 (N_14042,N_13885,N_13984);
or U14043 (N_14043,N_13914,N_13878);
and U14044 (N_14044,N_13876,N_13926);
nor U14045 (N_14045,N_13903,N_13918);
xnor U14046 (N_14046,N_13922,N_13995);
or U14047 (N_14047,N_13916,N_13961);
and U14048 (N_14048,N_13963,N_13892);
nand U14049 (N_14049,N_13966,N_13974);
xor U14050 (N_14050,N_13941,N_13891);
or U14051 (N_14051,N_13991,N_13909);
or U14052 (N_14052,N_13930,N_13944);
or U14053 (N_14053,N_13978,N_13901);
or U14054 (N_14054,N_13917,N_13956);
or U14055 (N_14055,N_13934,N_13972);
nor U14056 (N_14056,N_13967,N_13904);
xnor U14057 (N_14057,N_13911,N_13888);
and U14058 (N_14058,N_13957,N_13969);
xnor U14059 (N_14059,N_13902,N_13980);
and U14060 (N_14060,N_13951,N_13879);
nor U14061 (N_14061,N_13983,N_13936);
xnor U14062 (N_14062,N_13886,N_13999);
nor U14063 (N_14063,N_13899,N_13902);
and U14064 (N_14064,N_13910,N_13886);
nor U14065 (N_14065,N_13921,N_13966);
nand U14066 (N_14066,N_13973,N_13954);
nand U14067 (N_14067,N_13987,N_13905);
xnor U14068 (N_14068,N_13971,N_13921);
nand U14069 (N_14069,N_13938,N_13942);
or U14070 (N_14070,N_13897,N_13979);
xnor U14071 (N_14071,N_13977,N_13877);
xnor U14072 (N_14072,N_13970,N_13963);
xnor U14073 (N_14073,N_13889,N_13956);
nand U14074 (N_14074,N_13889,N_13916);
xnor U14075 (N_14075,N_13981,N_13903);
or U14076 (N_14076,N_13907,N_13934);
and U14077 (N_14077,N_13964,N_13961);
xnor U14078 (N_14078,N_13899,N_13877);
nor U14079 (N_14079,N_13908,N_13952);
nor U14080 (N_14080,N_13902,N_13884);
nand U14081 (N_14081,N_13898,N_13960);
xor U14082 (N_14082,N_13945,N_13921);
nor U14083 (N_14083,N_13915,N_13875);
and U14084 (N_14084,N_13997,N_13974);
xor U14085 (N_14085,N_13937,N_13889);
or U14086 (N_14086,N_13996,N_13889);
nor U14087 (N_14087,N_13943,N_13892);
or U14088 (N_14088,N_13900,N_13945);
and U14089 (N_14089,N_13973,N_13995);
nand U14090 (N_14090,N_13949,N_13958);
and U14091 (N_14091,N_13906,N_13974);
nand U14092 (N_14092,N_13953,N_13952);
and U14093 (N_14093,N_13984,N_13894);
nor U14094 (N_14094,N_13962,N_13918);
and U14095 (N_14095,N_13936,N_13935);
nand U14096 (N_14096,N_13998,N_13884);
or U14097 (N_14097,N_13968,N_13988);
or U14098 (N_14098,N_13900,N_13968);
nor U14099 (N_14099,N_13913,N_13887);
nand U14100 (N_14100,N_13902,N_13985);
xnor U14101 (N_14101,N_13894,N_13968);
or U14102 (N_14102,N_13898,N_13964);
or U14103 (N_14103,N_13968,N_13972);
and U14104 (N_14104,N_13908,N_13895);
nand U14105 (N_14105,N_13892,N_13971);
or U14106 (N_14106,N_13893,N_13966);
or U14107 (N_14107,N_13888,N_13922);
or U14108 (N_14108,N_13886,N_13951);
and U14109 (N_14109,N_13892,N_13913);
or U14110 (N_14110,N_13891,N_13998);
or U14111 (N_14111,N_13920,N_13917);
or U14112 (N_14112,N_13983,N_13998);
xor U14113 (N_14113,N_13909,N_13906);
and U14114 (N_14114,N_13927,N_13922);
nor U14115 (N_14115,N_13976,N_13902);
nand U14116 (N_14116,N_13991,N_13977);
nand U14117 (N_14117,N_13909,N_13914);
nand U14118 (N_14118,N_13941,N_13933);
nor U14119 (N_14119,N_13880,N_13975);
nand U14120 (N_14120,N_13970,N_13954);
nor U14121 (N_14121,N_13911,N_13997);
xnor U14122 (N_14122,N_13981,N_13933);
nor U14123 (N_14123,N_13950,N_13977);
or U14124 (N_14124,N_13887,N_13910);
or U14125 (N_14125,N_14073,N_14051);
or U14126 (N_14126,N_14064,N_14087);
xnor U14127 (N_14127,N_14111,N_14017);
xnor U14128 (N_14128,N_14098,N_14068);
nand U14129 (N_14129,N_14008,N_14114);
nor U14130 (N_14130,N_14034,N_14022);
or U14131 (N_14131,N_14023,N_14103);
and U14132 (N_14132,N_14077,N_14007);
nor U14133 (N_14133,N_14019,N_14108);
nand U14134 (N_14134,N_14083,N_14124);
and U14135 (N_14135,N_14041,N_14076);
nor U14136 (N_14136,N_14096,N_14009);
xnor U14137 (N_14137,N_14115,N_14052);
and U14138 (N_14138,N_14030,N_14021);
and U14139 (N_14139,N_14113,N_14048);
nor U14140 (N_14140,N_14045,N_14059);
nor U14141 (N_14141,N_14097,N_14006);
or U14142 (N_14142,N_14027,N_14122);
nor U14143 (N_14143,N_14025,N_14075);
nand U14144 (N_14144,N_14112,N_14013);
or U14145 (N_14145,N_14080,N_14101);
nand U14146 (N_14146,N_14010,N_14116);
and U14147 (N_14147,N_14053,N_14109);
nor U14148 (N_14148,N_14002,N_14038);
and U14149 (N_14149,N_14031,N_14082);
nor U14150 (N_14150,N_14047,N_14012);
or U14151 (N_14151,N_14079,N_14037);
or U14152 (N_14152,N_14090,N_14093);
xnor U14153 (N_14153,N_14107,N_14094);
nor U14154 (N_14154,N_14057,N_14042);
xor U14155 (N_14155,N_14065,N_14060);
nor U14156 (N_14156,N_14084,N_14049);
xnor U14157 (N_14157,N_14000,N_14016);
and U14158 (N_14158,N_14028,N_14100);
and U14159 (N_14159,N_14063,N_14001);
or U14160 (N_14160,N_14102,N_14099);
xor U14161 (N_14161,N_14061,N_14091);
nand U14162 (N_14162,N_14029,N_14043);
and U14163 (N_14163,N_14092,N_14072);
nor U14164 (N_14164,N_14069,N_14024);
nor U14165 (N_14165,N_14046,N_14056);
and U14166 (N_14166,N_14110,N_14011);
nand U14167 (N_14167,N_14074,N_14070);
or U14168 (N_14168,N_14085,N_14088);
nor U14169 (N_14169,N_14020,N_14005);
or U14170 (N_14170,N_14106,N_14036);
xor U14171 (N_14171,N_14123,N_14062);
or U14172 (N_14172,N_14033,N_14015);
and U14173 (N_14173,N_14120,N_14066);
xnor U14174 (N_14174,N_14119,N_14032);
xnor U14175 (N_14175,N_14078,N_14081);
xor U14176 (N_14176,N_14014,N_14071);
nand U14177 (N_14177,N_14117,N_14003);
xnor U14178 (N_14178,N_14104,N_14044);
nor U14179 (N_14179,N_14089,N_14105);
nor U14180 (N_14180,N_14121,N_14067);
or U14181 (N_14181,N_14004,N_14054);
or U14182 (N_14182,N_14118,N_14055);
nor U14183 (N_14183,N_14026,N_14058);
or U14184 (N_14184,N_14040,N_14018);
xnor U14185 (N_14185,N_14035,N_14039);
xnor U14186 (N_14186,N_14095,N_14050);
nand U14187 (N_14187,N_14086,N_14082);
or U14188 (N_14188,N_14010,N_14038);
or U14189 (N_14189,N_14092,N_14062);
nand U14190 (N_14190,N_14017,N_14120);
nor U14191 (N_14191,N_14012,N_14031);
or U14192 (N_14192,N_14086,N_14027);
xnor U14193 (N_14193,N_14097,N_14106);
or U14194 (N_14194,N_14120,N_14024);
or U14195 (N_14195,N_14044,N_14087);
nand U14196 (N_14196,N_14101,N_14096);
nor U14197 (N_14197,N_14097,N_14010);
or U14198 (N_14198,N_14092,N_14096);
nor U14199 (N_14199,N_14050,N_14037);
nor U14200 (N_14200,N_14086,N_14043);
nor U14201 (N_14201,N_14054,N_14103);
or U14202 (N_14202,N_14085,N_14062);
nor U14203 (N_14203,N_14009,N_14018);
xnor U14204 (N_14204,N_14086,N_14079);
and U14205 (N_14205,N_14087,N_14121);
nor U14206 (N_14206,N_14067,N_14063);
xor U14207 (N_14207,N_14105,N_14008);
xor U14208 (N_14208,N_14083,N_14060);
and U14209 (N_14209,N_14040,N_14033);
nand U14210 (N_14210,N_14021,N_14120);
nand U14211 (N_14211,N_14076,N_14111);
or U14212 (N_14212,N_14053,N_14011);
and U14213 (N_14213,N_14064,N_14107);
and U14214 (N_14214,N_14058,N_14120);
and U14215 (N_14215,N_14113,N_14052);
and U14216 (N_14216,N_14039,N_14100);
nor U14217 (N_14217,N_14011,N_14068);
xnor U14218 (N_14218,N_14031,N_14117);
and U14219 (N_14219,N_14023,N_14028);
nor U14220 (N_14220,N_14051,N_14094);
or U14221 (N_14221,N_14004,N_14049);
or U14222 (N_14222,N_14000,N_14059);
and U14223 (N_14223,N_14024,N_14084);
or U14224 (N_14224,N_14050,N_14015);
nor U14225 (N_14225,N_14062,N_14124);
nand U14226 (N_14226,N_14094,N_14124);
nand U14227 (N_14227,N_14062,N_14089);
or U14228 (N_14228,N_14119,N_14074);
nand U14229 (N_14229,N_14079,N_14031);
xor U14230 (N_14230,N_14040,N_14119);
nand U14231 (N_14231,N_14013,N_14038);
and U14232 (N_14232,N_14058,N_14105);
nor U14233 (N_14233,N_14047,N_14081);
and U14234 (N_14234,N_14124,N_14090);
or U14235 (N_14235,N_14083,N_14014);
nor U14236 (N_14236,N_14088,N_14056);
nand U14237 (N_14237,N_14013,N_14086);
xor U14238 (N_14238,N_14024,N_14010);
nand U14239 (N_14239,N_14090,N_14029);
nor U14240 (N_14240,N_14029,N_14042);
and U14241 (N_14241,N_14012,N_14037);
or U14242 (N_14242,N_14083,N_14028);
and U14243 (N_14243,N_14055,N_14006);
nor U14244 (N_14244,N_14109,N_14111);
nand U14245 (N_14245,N_14083,N_14054);
or U14246 (N_14246,N_14060,N_14042);
nand U14247 (N_14247,N_14056,N_14111);
and U14248 (N_14248,N_14073,N_14084);
and U14249 (N_14249,N_14101,N_14084);
and U14250 (N_14250,N_14152,N_14158);
nand U14251 (N_14251,N_14243,N_14185);
or U14252 (N_14252,N_14178,N_14220);
and U14253 (N_14253,N_14127,N_14193);
nand U14254 (N_14254,N_14165,N_14176);
nor U14255 (N_14255,N_14169,N_14140);
nand U14256 (N_14256,N_14190,N_14159);
or U14257 (N_14257,N_14160,N_14177);
or U14258 (N_14258,N_14211,N_14167);
xnor U14259 (N_14259,N_14137,N_14173);
nor U14260 (N_14260,N_14182,N_14210);
nor U14261 (N_14261,N_14235,N_14223);
nand U14262 (N_14262,N_14228,N_14163);
nor U14263 (N_14263,N_14237,N_14241);
or U14264 (N_14264,N_14191,N_14180);
xnor U14265 (N_14265,N_14156,N_14164);
and U14266 (N_14266,N_14227,N_14148);
nand U14267 (N_14267,N_14144,N_14179);
or U14268 (N_14268,N_14172,N_14147);
nor U14269 (N_14269,N_14206,N_14198);
xnor U14270 (N_14270,N_14189,N_14155);
or U14271 (N_14271,N_14192,N_14209);
and U14272 (N_14272,N_14151,N_14161);
xnor U14273 (N_14273,N_14232,N_14183);
and U14274 (N_14274,N_14146,N_14203);
nand U14275 (N_14275,N_14130,N_14226);
xnor U14276 (N_14276,N_14150,N_14145);
nand U14277 (N_14277,N_14157,N_14230);
or U14278 (N_14278,N_14149,N_14132);
xnor U14279 (N_14279,N_14187,N_14212);
xnor U14280 (N_14280,N_14143,N_14129);
xnor U14281 (N_14281,N_14205,N_14236);
nor U14282 (N_14282,N_14231,N_14171);
or U14283 (N_14283,N_14136,N_14181);
nor U14284 (N_14284,N_14201,N_14135);
nor U14285 (N_14285,N_14168,N_14217);
nand U14286 (N_14286,N_14204,N_14248);
nand U14287 (N_14287,N_14229,N_14186);
or U14288 (N_14288,N_14138,N_14128);
nor U14289 (N_14289,N_14166,N_14238);
nand U14290 (N_14290,N_14224,N_14188);
xnor U14291 (N_14291,N_14249,N_14125);
xor U14292 (N_14292,N_14214,N_14153);
nand U14293 (N_14293,N_14194,N_14246);
xnor U14294 (N_14294,N_14216,N_14233);
nor U14295 (N_14295,N_14134,N_14141);
nand U14296 (N_14296,N_14247,N_14170);
xor U14297 (N_14297,N_14126,N_14213);
xor U14298 (N_14298,N_14221,N_14218);
or U14299 (N_14299,N_14234,N_14154);
or U14300 (N_14300,N_14175,N_14142);
and U14301 (N_14301,N_14242,N_14208);
nor U14302 (N_14302,N_14195,N_14199);
xor U14303 (N_14303,N_14174,N_14244);
nand U14304 (N_14304,N_14197,N_14207);
nor U14305 (N_14305,N_14196,N_14184);
nand U14306 (N_14306,N_14131,N_14200);
and U14307 (N_14307,N_14215,N_14162);
or U14308 (N_14308,N_14219,N_14139);
and U14309 (N_14309,N_14202,N_14225);
or U14310 (N_14310,N_14245,N_14222);
and U14311 (N_14311,N_14133,N_14240);
nand U14312 (N_14312,N_14239,N_14159);
nand U14313 (N_14313,N_14154,N_14171);
or U14314 (N_14314,N_14140,N_14147);
nor U14315 (N_14315,N_14162,N_14198);
xor U14316 (N_14316,N_14168,N_14172);
nor U14317 (N_14317,N_14125,N_14187);
nor U14318 (N_14318,N_14190,N_14217);
or U14319 (N_14319,N_14137,N_14154);
and U14320 (N_14320,N_14205,N_14224);
and U14321 (N_14321,N_14176,N_14129);
and U14322 (N_14322,N_14132,N_14161);
nor U14323 (N_14323,N_14204,N_14247);
nand U14324 (N_14324,N_14136,N_14140);
nor U14325 (N_14325,N_14156,N_14172);
nand U14326 (N_14326,N_14243,N_14232);
or U14327 (N_14327,N_14152,N_14199);
and U14328 (N_14328,N_14235,N_14125);
xor U14329 (N_14329,N_14130,N_14230);
xor U14330 (N_14330,N_14139,N_14177);
nand U14331 (N_14331,N_14223,N_14193);
and U14332 (N_14332,N_14228,N_14213);
xnor U14333 (N_14333,N_14135,N_14213);
xor U14334 (N_14334,N_14246,N_14197);
xor U14335 (N_14335,N_14203,N_14194);
or U14336 (N_14336,N_14196,N_14202);
nand U14337 (N_14337,N_14246,N_14222);
or U14338 (N_14338,N_14166,N_14141);
nand U14339 (N_14339,N_14220,N_14138);
xnor U14340 (N_14340,N_14175,N_14168);
xnor U14341 (N_14341,N_14205,N_14193);
xnor U14342 (N_14342,N_14238,N_14135);
or U14343 (N_14343,N_14145,N_14191);
xor U14344 (N_14344,N_14150,N_14139);
or U14345 (N_14345,N_14158,N_14247);
or U14346 (N_14346,N_14217,N_14179);
or U14347 (N_14347,N_14158,N_14188);
and U14348 (N_14348,N_14132,N_14211);
and U14349 (N_14349,N_14249,N_14181);
nor U14350 (N_14350,N_14130,N_14214);
and U14351 (N_14351,N_14194,N_14154);
nor U14352 (N_14352,N_14192,N_14153);
xor U14353 (N_14353,N_14225,N_14245);
xor U14354 (N_14354,N_14214,N_14212);
or U14355 (N_14355,N_14214,N_14188);
or U14356 (N_14356,N_14136,N_14212);
nand U14357 (N_14357,N_14192,N_14201);
nor U14358 (N_14358,N_14204,N_14152);
nand U14359 (N_14359,N_14217,N_14218);
and U14360 (N_14360,N_14245,N_14138);
xor U14361 (N_14361,N_14141,N_14232);
xnor U14362 (N_14362,N_14198,N_14179);
xor U14363 (N_14363,N_14169,N_14128);
xor U14364 (N_14364,N_14241,N_14224);
nand U14365 (N_14365,N_14214,N_14135);
nor U14366 (N_14366,N_14172,N_14177);
or U14367 (N_14367,N_14153,N_14236);
nor U14368 (N_14368,N_14171,N_14135);
or U14369 (N_14369,N_14140,N_14154);
nor U14370 (N_14370,N_14242,N_14203);
xor U14371 (N_14371,N_14199,N_14217);
or U14372 (N_14372,N_14225,N_14215);
xor U14373 (N_14373,N_14155,N_14136);
nand U14374 (N_14374,N_14185,N_14248);
nand U14375 (N_14375,N_14307,N_14325);
xor U14376 (N_14376,N_14314,N_14258);
nand U14377 (N_14377,N_14322,N_14369);
xnor U14378 (N_14378,N_14294,N_14275);
or U14379 (N_14379,N_14335,N_14374);
xor U14380 (N_14380,N_14306,N_14256);
and U14381 (N_14381,N_14330,N_14336);
nor U14382 (N_14382,N_14349,N_14362);
nor U14383 (N_14383,N_14341,N_14360);
or U14384 (N_14384,N_14264,N_14346);
or U14385 (N_14385,N_14357,N_14365);
and U14386 (N_14386,N_14254,N_14354);
nand U14387 (N_14387,N_14276,N_14350);
or U14388 (N_14388,N_14323,N_14293);
nand U14389 (N_14389,N_14372,N_14267);
or U14390 (N_14390,N_14319,N_14257);
nor U14391 (N_14391,N_14344,N_14290);
nand U14392 (N_14392,N_14270,N_14315);
xor U14393 (N_14393,N_14373,N_14329);
nand U14394 (N_14394,N_14255,N_14281);
nand U14395 (N_14395,N_14269,N_14340);
xor U14396 (N_14396,N_14310,N_14288);
xnor U14397 (N_14397,N_14320,N_14298);
xor U14398 (N_14398,N_14282,N_14287);
nor U14399 (N_14399,N_14368,N_14345);
xnor U14400 (N_14400,N_14356,N_14263);
nor U14401 (N_14401,N_14291,N_14366);
nor U14402 (N_14402,N_14347,N_14250);
nand U14403 (N_14403,N_14266,N_14338);
xor U14404 (N_14404,N_14337,N_14268);
nand U14405 (N_14405,N_14280,N_14311);
nor U14406 (N_14406,N_14284,N_14262);
and U14407 (N_14407,N_14334,N_14261);
or U14408 (N_14408,N_14265,N_14318);
nand U14409 (N_14409,N_14364,N_14363);
nand U14410 (N_14410,N_14292,N_14332);
and U14411 (N_14411,N_14260,N_14299);
nor U14412 (N_14412,N_14339,N_14342);
and U14413 (N_14413,N_14316,N_14326);
and U14414 (N_14414,N_14273,N_14277);
nor U14415 (N_14415,N_14328,N_14321);
or U14416 (N_14416,N_14300,N_14353);
xor U14417 (N_14417,N_14271,N_14355);
nand U14418 (N_14418,N_14252,N_14305);
and U14419 (N_14419,N_14274,N_14303);
xor U14420 (N_14420,N_14331,N_14309);
or U14421 (N_14421,N_14333,N_14352);
and U14422 (N_14422,N_14317,N_14253);
nand U14423 (N_14423,N_14278,N_14324);
and U14424 (N_14424,N_14259,N_14297);
and U14425 (N_14425,N_14286,N_14367);
xor U14426 (N_14426,N_14295,N_14313);
or U14427 (N_14427,N_14343,N_14285);
nand U14428 (N_14428,N_14296,N_14272);
or U14429 (N_14429,N_14348,N_14361);
and U14430 (N_14430,N_14359,N_14251);
nand U14431 (N_14431,N_14301,N_14283);
xor U14432 (N_14432,N_14308,N_14312);
xnor U14433 (N_14433,N_14304,N_14351);
nor U14434 (N_14434,N_14371,N_14327);
nor U14435 (N_14435,N_14289,N_14279);
nand U14436 (N_14436,N_14358,N_14302);
nand U14437 (N_14437,N_14370,N_14305);
or U14438 (N_14438,N_14288,N_14324);
and U14439 (N_14439,N_14351,N_14328);
xnor U14440 (N_14440,N_14267,N_14273);
nand U14441 (N_14441,N_14278,N_14294);
nor U14442 (N_14442,N_14258,N_14327);
xor U14443 (N_14443,N_14358,N_14296);
and U14444 (N_14444,N_14282,N_14315);
nand U14445 (N_14445,N_14259,N_14334);
or U14446 (N_14446,N_14343,N_14365);
nor U14447 (N_14447,N_14333,N_14366);
or U14448 (N_14448,N_14372,N_14273);
nand U14449 (N_14449,N_14256,N_14339);
nor U14450 (N_14450,N_14351,N_14330);
nand U14451 (N_14451,N_14304,N_14318);
and U14452 (N_14452,N_14272,N_14255);
xor U14453 (N_14453,N_14261,N_14336);
xnor U14454 (N_14454,N_14324,N_14254);
and U14455 (N_14455,N_14292,N_14353);
nor U14456 (N_14456,N_14267,N_14298);
or U14457 (N_14457,N_14265,N_14300);
xnor U14458 (N_14458,N_14256,N_14278);
and U14459 (N_14459,N_14326,N_14252);
xor U14460 (N_14460,N_14316,N_14335);
or U14461 (N_14461,N_14324,N_14302);
xor U14462 (N_14462,N_14349,N_14263);
nand U14463 (N_14463,N_14293,N_14332);
xor U14464 (N_14464,N_14347,N_14308);
and U14465 (N_14465,N_14366,N_14252);
nand U14466 (N_14466,N_14258,N_14328);
nor U14467 (N_14467,N_14282,N_14279);
nor U14468 (N_14468,N_14288,N_14335);
and U14469 (N_14469,N_14360,N_14372);
nor U14470 (N_14470,N_14294,N_14263);
nand U14471 (N_14471,N_14331,N_14261);
nand U14472 (N_14472,N_14334,N_14293);
nor U14473 (N_14473,N_14349,N_14294);
or U14474 (N_14474,N_14273,N_14374);
xnor U14475 (N_14475,N_14267,N_14300);
xnor U14476 (N_14476,N_14320,N_14282);
xor U14477 (N_14477,N_14347,N_14283);
and U14478 (N_14478,N_14332,N_14259);
xor U14479 (N_14479,N_14287,N_14362);
or U14480 (N_14480,N_14356,N_14333);
nor U14481 (N_14481,N_14359,N_14317);
and U14482 (N_14482,N_14277,N_14339);
xnor U14483 (N_14483,N_14373,N_14348);
or U14484 (N_14484,N_14256,N_14298);
and U14485 (N_14485,N_14319,N_14298);
and U14486 (N_14486,N_14325,N_14345);
or U14487 (N_14487,N_14261,N_14341);
nand U14488 (N_14488,N_14334,N_14260);
and U14489 (N_14489,N_14354,N_14323);
or U14490 (N_14490,N_14302,N_14357);
and U14491 (N_14491,N_14319,N_14367);
xnor U14492 (N_14492,N_14330,N_14345);
or U14493 (N_14493,N_14281,N_14356);
and U14494 (N_14494,N_14325,N_14373);
or U14495 (N_14495,N_14258,N_14277);
nand U14496 (N_14496,N_14283,N_14350);
or U14497 (N_14497,N_14275,N_14273);
nor U14498 (N_14498,N_14367,N_14296);
xnor U14499 (N_14499,N_14322,N_14263);
and U14500 (N_14500,N_14375,N_14434);
nor U14501 (N_14501,N_14465,N_14497);
nand U14502 (N_14502,N_14445,N_14407);
and U14503 (N_14503,N_14397,N_14444);
and U14504 (N_14504,N_14457,N_14386);
nor U14505 (N_14505,N_14414,N_14449);
nor U14506 (N_14506,N_14395,N_14472);
or U14507 (N_14507,N_14468,N_14381);
xor U14508 (N_14508,N_14470,N_14393);
nand U14509 (N_14509,N_14463,N_14428);
nor U14510 (N_14510,N_14438,N_14439);
nor U14511 (N_14511,N_14394,N_14420);
nor U14512 (N_14512,N_14402,N_14419);
and U14513 (N_14513,N_14400,N_14443);
or U14514 (N_14514,N_14454,N_14426);
xor U14515 (N_14515,N_14433,N_14416);
and U14516 (N_14516,N_14485,N_14398);
nand U14517 (N_14517,N_14489,N_14427);
xnor U14518 (N_14518,N_14496,N_14459);
and U14519 (N_14519,N_14392,N_14480);
nand U14520 (N_14520,N_14477,N_14490);
or U14521 (N_14521,N_14475,N_14474);
nor U14522 (N_14522,N_14429,N_14435);
nand U14523 (N_14523,N_14483,N_14430);
or U14524 (N_14524,N_14462,N_14432);
xnor U14525 (N_14525,N_14442,N_14441);
nor U14526 (N_14526,N_14379,N_14384);
nand U14527 (N_14527,N_14380,N_14401);
and U14528 (N_14528,N_14437,N_14415);
nand U14529 (N_14529,N_14486,N_14455);
and U14530 (N_14530,N_14447,N_14425);
or U14531 (N_14531,N_14493,N_14453);
nor U14532 (N_14532,N_14417,N_14450);
and U14533 (N_14533,N_14484,N_14421);
and U14534 (N_14534,N_14498,N_14409);
nand U14535 (N_14535,N_14405,N_14469);
nand U14536 (N_14536,N_14488,N_14388);
nand U14537 (N_14537,N_14451,N_14391);
xnor U14538 (N_14538,N_14385,N_14390);
nor U14539 (N_14539,N_14431,N_14436);
xnor U14540 (N_14540,N_14456,N_14424);
nor U14541 (N_14541,N_14458,N_14478);
nor U14542 (N_14542,N_14422,N_14413);
or U14543 (N_14543,N_14452,N_14448);
and U14544 (N_14544,N_14404,N_14499);
nor U14545 (N_14545,N_14403,N_14411);
nand U14546 (N_14546,N_14377,N_14382);
nand U14547 (N_14547,N_14464,N_14473);
xor U14548 (N_14548,N_14410,N_14461);
nand U14549 (N_14549,N_14383,N_14479);
or U14550 (N_14550,N_14467,N_14399);
nand U14551 (N_14551,N_14412,N_14389);
nor U14552 (N_14552,N_14471,N_14440);
xnor U14553 (N_14553,N_14466,N_14495);
or U14554 (N_14554,N_14446,N_14481);
xnor U14555 (N_14555,N_14494,N_14491);
nand U14556 (N_14556,N_14492,N_14408);
nand U14557 (N_14557,N_14482,N_14423);
nor U14558 (N_14558,N_14378,N_14476);
xor U14559 (N_14559,N_14487,N_14418);
or U14560 (N_14560,N_14376,N_14460);
nor U14561 (N_14561,N_14396,N_14406);
xnor U14562 (N_14562,N_14387,N_14402);
or U14563 (N_14563,N_14424,N_14388);
or U14564 (N_14564,N_14412,N_14456);
xnor U14565 (N_14565,N_14466,N_14490);
and U14566 (N_14566,N_14461,N_14482);
nand U14567 (N_14567,N_14398,N_14409);
nor U14568 (N_14568,N_14411,N_14455);
and U14569 (N_14569,N_14417,N_14480);
nand U14570 (N_14570,N_14451,N_14439);
nor U14571 (N_14571,N_14472,N_14437);
and U14572 (N_14572,N_14464,N_14469);
xor U14573 (N_14573,N_14443,N_14421);
nor U14574 (N_14574,N_14450,N_14494);
nor U14575 (N_14575,N_14463,N_14484);
nand U14576 (N_14576,N_14433,N_14387);
xnor U14577 (N_14577,N_14472,N_14418);
nor U14578 (N_14578,N_14406,N_14469);
or U14579 (N_14579,N_14458,N_14399);
nand U14580 (N_14580,N_14396,N_14486);
and U14581 (N_14581,N_14412,N_14454);
xor U14582 (N_14582,N_14486,N_14376);
nor U14583 (N_14583,N_14487,N_14401);
nand U14584 (N_14584,N_14395,N_14452);
nor U14585 (N_14585,N_14393,N_14490);
and U14586 (N_14586,N_14488,N_14485);
or U14587 (N_14587,N_14489,N_14449);
xor U14588 (N_14588,N_14486,N_14398);
xor U14589 (N_14589,N_14492,N_14435);
and U14590 (N_14590,N_14440,N_14499);
and U14591 (N_14591,N_14394,N_14453);
xnor U14592 (N_14592,N_14419,N_14479);
nand U14593 (N_14593,N_14408,N_14473);
and U14594 (N_14594,N_14436,N_14473);
nand U14595 (N_14595,N_14406,N_14431);
nand U14596 (N_14596,N_14391,N_14406);
or U14597 (N_14597,N_14417,N_14379);
nor U14598 (N_14598,N_14497,N_14470);
and U14599 (N_14599,N_14419,N_14388);
or U14600 (N_14600,N_14490,N_14445);
nor U14601 (N_14601,N_14499,N_14395);
nand U14602 (N_14602,N_14482,N_14391);
nand U14603 (N_14603,N_14415,N_14416);
nor U14604 (N_14604,N_14390,N_14447);
xnor U14605 (N_14605,N_14392,N_14394);
nand U14606 (N_14606,N_14391,N_14398);
and U14607 (N_14607,N_14375,N_14446);
nor U14608 (N_14608,N_14422,N_14417);
or U14609 (N_14609,N_14422,N_14489);
xor U14610 (N_14610,N_14468,N_14375);
and U14611 (N_14611,N_14447,N_14405);
xnor U14612 (N_14612,N_14446,N_14387);
xnor U14613 (N_14613,N_14457,N_14409);
xnor U14614 (N_14614,N_14438,N_14486);
xor U14615 (N_14615,N_14379,N_14479);
xor U14616 (N_14616,N_14452,N_14387);
xnor U14617 (N_14617,N_14480,N_14439);
and U14618 (N_14618,N_14406,N_14446);
nor U14619 (N_14619,N_14440,N_14389);
nand U14620 (N_14620,N_14459,N_14422);
nor U14621 (N_14621,N_14443,N_14464);
or U14622 (N_14622,N_14417,N_14388);
xnor U14623 (N_14623,N_14379,N_14408);
nor U14624 (N_14624,N_14414,N_14411);
and U14625 (N_14625,N_14524,N_14521);
nor U14626 (N_14626,N_14512,N_14598);
or U14627 (N_14627,N_14567,N_14518);
xor U14628 (N_14628,N_14551,N_14547);
nand U14629 (N_14629,N_14624,N_14592);
xnor U14630 (N_14630,N_14613,N_14610);
or U14631 (N_14631,N_14515,N_14594);
or U14632 (N_14632,N_14591,N_14590);
xnor U14633 (N_14633,N_14579,N_14607);
and U14634 (N_14634,N_14614,N_14585);
nand U14635 (N_14635,N_14573,N_14501);
xnor U14636 (N_14636,N_14576,N_14578);
or U14637 (N_14637,N_14517,N_14570);
nor U14638 (N_14638,N_14522,N_14619);
or U14639 (N_14639,N_14623,N_14596);
or U14640 (N_14640,N_14548,N_14603);
and U14641 (N_14641,N_14510,N_14565);
nor U14642 (N_14642,N_14611,N_14526);
or U14643 (N_14643,N_14597,N_14513);
nand U14644 (N_14644,N_14507,N_14555);
nand U14645 (N_14645,N_14519,N_14534);
nor U14646 (N_14646,N_14580,N_14504);
and U14647 (N_14647,N_14581,N_14599);
or U14648 (N_14648,N_14538,N_14574);
nand U14649 (N_14649,N_14546,N_14533);
or U14650 (N_14650,N_14568,N_14500);
xor U14651 (N_14651,N_14604,N_14560);
nor U14652 (N_14652,N_14527,N_14605);
nor U14653 (N_14653,N_14525,N_14539);
or U14654 (N_14654,N_14587,N_14564);
nor U14655 (N_14655,N_14621,N_14561);
nand U14656 (N_14656,N_14584,N_14540);
nor U14657 (N_14657,N_14528,N_14503);
nor U14658 (N_14658,N_14549,N_14558);
xor U14659 (N_14659,N_14616,N_14536);
xnor U14660 (N_14660,N_14618,N_14520);
xnor U14661 (N_14661,N_14617,N_14532);
nand U14662 (N_14662,N_14552,N_14535);
and U14663 (N_14663,N_14550,N_14569);
nand U14664 (N_14664,N_14529,N_14505);
nor U14665 (N_14665,N_14553,N_14506);
nand U14666 (N_14666,N_14582,N_14543);
and U14667 (N_14667,N_14537,N_14523);
nand U14668 (N_14668,N_14559,N_14609);
nor U14669 (N_14669,N_14541,N_14588);
nor U14670 (N_14670,N_14571,N_14562);
xor U14671 (N_14671,N_14586,N_14595);
nor U14672 (N_14672,N_14554,N_14602);
or U14673 (N_14673,N_14572,N_14589);
nor U14674 (N_14674,N_14622,N_14600);
or U14675 (N_14675,N_14601,N_14583);
and U14676 (N_14676,N_14531,N_14516);
nand U14677 (N_14677,N_14514,N_14575);
nand U14678 (N_14678,N_14563,N_14556);
nor U14679 (N_14679,N_14542,N_14530);
nand U14680 (N_14680,N_14545,N_14508);
xor U14681 (N_14681,N_14612,N_14511);
or U14682 (N_14682,N_14608,N_14593);
nor U14683 (N_14683,N_14502,N_14509);
nor U14684 (N_14684,N_14557,N_14620);
nor U14685 (N_14685,N_14615,N_14544);
xor U14686 (N_14686,N_14577,N_14566);
nor U14687 (N_14687,N_14606,N_14522);
nand U14688 (N_14688,N_14591,N_14564);
and U14689 (N_14689,N_14607,N_14515);
or U14690 (N_14690,N_14512,N_14526);
or U14691 (N_14691,N_14597,N_14580);
and U14692 (N_14692,N_14620,N_14537);
xor U14693 (N_14693,N_14541,N_14514);
or U14694 (N_14694,N_14577,N_14580);
xnor U14695 (N_14695,N_14605,N_14532);
or U14696 (N_14696,N_14574,N_14604);
xnor U14697 (N_14697,N_14614,N_14583);
and U14698 (N_14698,N_14576,N_14513);
and U14699 (N_14699,N_14505,N_14603);
and U14700 (N_14700,N_14572,N_14575);
xor U14701 (N_14701,N_14575,N_14536);
xnor U14702 (N_14702,N_14555,N_14577);
nand U14703 (N_14703,N_14570,N_14617);
or U14704 (N_14704,N_14586,N_14605);
and U14705 (N_14705,N_14523,N_14557);
xnor U14706 (N_14706,N_14603,N_14518);
nor U14707 (N_14707,N_14609,N_14590);
nand U14708 (N_14708,N_14558,N_14577);
and U14709 (N_14709,N_14540,N_14516);
xor U14710 (N_14710,N_14560,N_14516);
xor U14711 (N_14711,N_14570,N_14600);
or U14712 (N_14712,N_14613,N_14558);
xnor U14713 (N_14713,N_14525,N_14516);
and U14714 (N_14714,N_14508,N_14568);
xor U14715 (N_14715,N_14561,N_14500);
nor U14716 (N_14716,N_14533,N_14583);
nand U14717 (N_14717,N_14617,N_14511);
nor U14718 (N_14718,N_14615,N_14532);
or U14719 (N_14719,N_14554,N_14528);
and U14720 (N_14720,N_14501,N_14524);
nor U14721 (N_14721,N_14504,N_14543);
xor U14722 (N_14722,N_14561,N_14603);
nor U14723 (N_14723,N_14601,N_14514);
or U14724 (N_14724,N_14616,N_14587);
nor U14725 (N_14725,N_14531,N_14600);
xnor U14726 (N_14726,N_14582,N_14606);
nand U14727 (N_14727,N_14605,N_14608);
nor U14728 (N_14728,N_14615,N_14579);
xor U14729 (N_14729,N_14584,N_14530);
or U14730 (N_14730,N_14530,N_14515);
xnor U14731 (N_14731,N_14562,N_14523);
nor U14732 (N_14732,N_14533,N_14586);
nand U14733 (N_14733,N_14546,N_14521);
nor U14734 (N_14734,N_14516,N_14521);
or U14735 (N_14735,N_14538,N_14514);
nand U14736 (N_14736,N_14582,N_14563);
nand U14737 (N_14737,N_14543,N_14595);
xor U14738 (N_14738,N_14606,N_14590);
and U14739 (N_14739,N_14517,N_14504);
nand U14740 (N_14740,N_14552,N_14536);
nor U14741 (N_14741,N_14622,N_14580);
nor U14742 (N_14742,N_14525,N_14562);
nand U14743 (N_14743,N_14590,N_14525);
nand U14744 (N_14744,N_14539,N_14616);
nor U14745 (N_14745,N_14589,N_14518);
xnor U14746 (N_14746,N_14596,N_14609);
or U14747 (N_14747,N_14619,N_14590);
xnor U14748 (N_14748,N_14623,N_14609);
or U14749 (N_14749,N_14598,N_14544);
nand U14750 (N_14750,N_14731,N_14638);
and U14751 (N_14751,N_14675,N_14739);
xor U14752 (N_14752,N_14634,N_14656);
xor U14753 (N_14753,N_14691,N_14724);
xor U14754 (N_14754,N_14690,N_14736);
and U14755 (N_14755,N_14685,N_14651);
or U14756 (N_14756,N_14672,N_14734);
nor U14757 (N_14757,N_14646,N_14700);
nand U14758 (N_14758,N_14657,N_14729);
xnor U14759 (N_14759,N_14655,N_14706);
xnor U14760 (N_14760,N_14716,N_14707);
nor U14761 (N_14761,N_14689,N_14713);
or U14762 (N_14762,N_14649,N_14653);
and U14763 (N_14763,N_14682,N_14712);
nor U14764 (N_14764,N_14666,N_14635);
nand U14765 (N_14765,N_14696,N_14714);
xnor U14766 (N_14766,N_14630,N_14715);
nand U14767 (N_14767,N_14744,N_14628);
nor U14768 (N_14768,N_14721,N_14665);
xnor U14769 (N_14769,N_14722,N_14702);
and U14770 (N_14770,N_14699,N_14667);
nor U14771 (N_14771,N_14726,N_14684);
or U14772 (N_14772,N_14677,N_14629);
and U14773 (N_14773,N_14743,N_14633);
nand U14774 (N_14774,N_14660,N_14661);
or U14775 (N_14775,N_14710,N_14676);
nor U14776 (N_14776,N_14705,N_14674);
nor U14777 (N_14777,N_14701,N_14748);
nand U14778 (N_14778,N_14732,N_14664);
xor U14779 (N_14779,N_14745,N_14703);
nand U14780 (N_14780,N_14718,N_14632);
and U14781 (N_14781,N_14730,N_14727);
and U14782 (N_14782,N_14687,N_14668);
nor U14783 (N_14783,N_14637,N_14695);
nor U14784 (N_14784,N_14709,N_14673);
xnor U14785 (N_14785,N_14738,N_14642);
nand U14786 (N_14786,N_14688,N_14693);
xnor U14787 (N_14787,N_14670,N_14742);
or U14788 (N_14788,N_14694,N_14711);
and U14789 (N_14789,N_14717,N_14650);
nand U14790 (N_14790,N_14678,N_14704);
nor U14791 (N_14791,N_14698,N_14733);
nand U14792 (N_14792,N_14680,N_14708);
xor U14793 (N_14793,N_14627,N_14692);
nor U14794 (N_14794,N_14643,N_14697);
and U14795 (N_14795,N_14639,N_14679);
or U14796 (N_14796,N_14654,N_14648);
and U14797 (N_14797,N_14652,N_14681);
and U14798 (N_14798,N_14662,N_14625);
xnor U14799 (N_14799,N_14645,N_14647);
nor U14800 (N_14800,N_14659,N_14746);
and U14801 (N_14801,N_14658,N_14741);
nand U14802 (N_14802,N_14669,N_14720);
nand U14803 (N_14803,N_14747,N_14686);
nor U14804 (N_14804,N_14640,N_14626);
or U14805 (N_14805,N_14636,N_14671);
and U14806 (N_14806,N_14644,N_14723);
nand U14807 (N_14807,N_14728,N_14737);
and U14808 (N_14808,N_14725,N_14735);
and U14809 (N_14809,N_14663,N_14631);
nand U14810 (N_14810,N_14749,N_14719);
xor U14811 (N_14811,N_14740,N_14683);
nor U14812 (N_14812,N_14641,N_14625);
or U14813 (N_14813,N_14655,N_14708);
xnor U14814 (N_14814,N_14682,N_14726);
nand U14815 (N_14815,N_14740,N_14659);
nand U14816 (N_14816,N_14649,N_14725);
nand U14817 (N_14817,N_14710,N_14696);
and U14818 (N_14818,N_14668,N_14729);
xnor U14819 (N_14819,N_14650,N_14676);
or U14820 (N_14820,N_14721,N_14711);
nand U14821 (N_14821,N_14667,N_14689);
or U14822 (N_14822,N_14688,N_14709);
xor U14823 (N_14823,N_14639,N_14671);
nand U14824 (N_14824,N_14651,N_14716);
nor U14825 (N_14825,N_14708,N_14748);
or U14826 (N_14826,N_14630,N_14675);
nor U14827 (N_14827,N_14634,N_14666);
nor U14828 (N_14828,N_14645,N_14700);
nor U14829 (N_14829,N_14711,N_14661);
nand U14830 (N_14830,N_14625,N_14699);
nor U14831 (N_14831,N_14625,N_14647);
or U14832 (N_14832,N_14731,N_14729);
nand U14833 (N_14833,N_14674,N_14670);
nor U14834 (N_14834,N_14634,N_14628);
nor U14835 (N_14835,N_14707,N_14741);
xnor U14836 (N_14836,N_14726,N_14713);
nand U14837 (N_14837,N_14625,N_14702);
nor U14838 (N_14838,N_14626,N_14699);
xnor U14839 (N_14839,N_14683,N_14671);
and U14840 (N_14840,N_14701,N_14731);
xnor U14841 (N_14841,N_14661,N_14739);
nor U14842 (N_14842,N_14712,N_14711);
or U14843 (N_14843,N_14712,N_14630);
or U14844 (N_14844,N_14678,N_14663);
nand U14845 (N_14845,N_14690,N_14705);
xor U14846 (N_14846,N_14660,N_14689);
and U14847 (N_14847,N_14626,N_14740);
nand U14848 (N_14848,N_14702,N_14738);
nor U14849 (N_14849,N_14740,N_14640);
nand U14850 (N_14850,N_14734,N_14650);
and U14851 (N_14851,N_14687,N_14667);
nand U14852 (N_14852,N_14626,N_14694);
xnor U14853 (N_14853,N_14692,N_14735);
xnor U14854 (N_14854,N_14651,N_14640);
xnor U14855 (N_14855,N_14713,N_14670);
xor U14856 (N_14856,N_14638,N_14694);
or U14857 (N_14857,N_14643,N_14666);
xnor U14858 (N_14858,N_14709,N_14738);
nor U14859 (N_14859,N_14689,N_14642);
or U14860 (N_14860,N_14662,N_14697);
or U14861 (N_14861,N_14711,N_14710);
nor U14862 (N_14862,N_14625,N_14697);
or U14863 (N_14863,N_14629,N_14634);
or U14864 (N_14864,N_14744,N_14666);
nor U14865 (N_14865,N_14717,N_14636);
or U14866 (N_14866,N_14653,N_14678);
nand U14867 (N_14867,N_14728,N_14677);
xnor U14868 (N_14868,N_14672,N_14694);
xnor U14869 (N_14869,N_14690,N_14647);
and U14870 (N_14870,N_14749,N_14693);
xnor U14871 (N_14871,N_14717,N_14632);
xor U14872 (N_14872,N_14710,N_14627);
nor U14873 (N_14873,N_14744,N_14678);
or U14874 (N_14874,N_14713,N_14696);
and U14875 (N_14875,N_14843,N_14790);
nor U14876 (N_14876,N_14776,N_14831);
nor U14877 (N_14877,N_14772,N_14841);
nor U14878 (N_14878,N_14784,N_14751);
or U14879 (N_14879,N_14823,N_14762);
and U14880 (N_14880,N_14811,N_14805);
nor U14881 (N_14881,N_14809,N_14803);
or U14882 (N_14882,N_14781,N_14782);
and U14883 (N_14883,N_14807,N_14839);
nand U14884 (N_14884,N_14791,N_14793);
xnor U14885 (N_14885,N_14800,N_14820);
or U14886 (N_14886,N_14761,N_14840);
and U14887 (N_14887,N_14774,N_14851);
xnor U14888 (N_14888,N_14765,N_14810);
or U14889 (N_14889,N_14873,N_14788);
and U14890 (N_14890,N_14799,N_14853);
nand U14891 (N_14891,N_14814,N_14794);
and U14892 (N_14892,N_14834,N_14802);
xor U14893 (N_14893,N_14871,N_14767);
nand U14894 (N_14894,N_14849,N_14816);
nand U14895 (N_14895,N_14847,N_14861);
xor U14896 (N_14896,N_14797,N_14842);
nand U14897 (N_14897,N_14779,N_14862);
xor U14898 (N_14898,N_14815,N_14818);
and U14899 (N_14899,N_14753,N_14783);
nor U14900 (N_14900,N_14764,N_14826);
or U14901 (N_14901,N_14758,N_14798);
or U14902 (N_14902,N_14827,N_14837);
or U14903 (N_14903,N_14756,N_14838);
xnor U14904 (N_14904,N_14845,N_14770);
nor U14905 (N_14905,N_14795,N_14808);
nand U14906 (N_14906,N_14866,N_14868);
xor U14907 (N_14907,N_14848,N_14759);
nor U14908 (N_14908,N_14817,N_14771);
nand U14909 (N_14909,N_14796,N_14863);
nand U14910 (N_14910,N_14760,N_14768);
nand U14911 (N_14911,N_14850,N_14828);
xor U14912 (N_14912,N_14836,N_14824);
nand U14913 (N_14913,N_14773,N_14789);
nor U14914 (N_14914,N_14801,N_14830);
or U14915 (N_14915,N_14869,N_14752);
nor U14916 (N_14916,N_14785,N_14835);
nor U14917 (N_14917,N_14872,N_14860);
nand U14918 (N_14918,N_14786,N_14775);
or U14919 (N_14919,N_14874,N_14819);
nand U14920 (N_14920,N_14792,N_14754);
and U14921 (N_14921,N_14855,N_14858);
and U14922 (N_14922,N_14804,N_14778);
xnor U14923 (N_14923,N_14854,N_14755);
and U14924 (N_14924,N_14859,N_14812);
nand U14925 (N_14925,N_14750,N_14832);
nand U14926 (N_14926,N_14766,N_14829);
xnor U14927 (N_14927,N_14856,N_14865);
nand U14928 (N_14928,N_14757,N_14825);
or U14929 (N_14929,N_14870,N_14769);
nor U14930 (N_14930,N_14846,N_14864);
or U14931 (N_14931,N_14813,N_14852);
nor U14932 (N_14932,N_14763,N_14833);
or U14933 (N_14933,N_14787,N_14821);
xnor U14934 (N_14934,N_14857,N_14822);
and U14935 (N_14935,N_14806,N_14844);
and U14936 (N_14936,N_14780,N_14867);
nand U14937 (N_14937,N_14777,N_14847);
nor U14938 (N_14938,N_14786,N_14761);
nor U14939 (N_14939,N_14823,N_14870);
and U14940 (N_14940,N_14786,N_14839);
xnor U14941 (N_14941,N_14831,N_14830);
and U14942 (N_14942,N_14856,N_14827);
xnor U14943 (N_14943,N_14781,N_14777);
nand U14944 (N_14944,N_14843,N_14755);
xnor U14945 (N_14945,N_14840,N_14784);
xnor U14946 (N_14946,N_14845,N_14862);
nor U14947 (N_14947,N_14857,N_14869);
or U14948 (N_14948,N_14792,N_14854);
nand U14949 (N_14949,N_14775,N_14857);
or U14950 (N_14950,N_14840,N_14801);
or U14951 (N_14951,N_14782,N_14851);
xnor U14952 (N_14952,N_14800,N_14798);
or U14953 (N_14953,N_14853,N_14773);
nand U14954 (N_14954,N_14849,N_14819);
xnor U14955 (N_14955,N_14814,N_14870);
and U14956 (N_14956,N_14768,N_14773);
or U14957 (N_14957,N_14829,N_14804);
nor U14958 (N_14958,N_14827,N_14795);
nor U14959 (N_14959,N_14817,N_14869);
xnor U14960 (N_14960,N_14802,N_14779);
nand U14961 (N_14961,N_14799,N_14842);
nor U14962 (N_14962,N_14793,N_14844);
xor U14963 (N_14963,N_14771,N_14872);
and U14964 (N_14964,N_14868,N_14793);
nor U14965 (N_14965,N_14800,N_14815);
or U14966 (N_14966,N_14847,N_14868);
and U14967 (N_14967,N_14850,N_14782);
and U14968 (N_14968,N_14760,N_14823);
xnor U14969 (N_14969,N_14750,N_14812);
xnor U14970 (N_14970,N_14853,N_14761);
xnor U14971 (N_14971,N_14837,N_14843);
nand U14972 (N_14972,N_14818,N_14870);
or U14973 (N_14973,N_14823,N_14776);
or U14974 (N_14974,N_14752,N_14780);
nand U14975 (N_14975,N_14783,N_14838);
and U14976 (N_14976,N_14867,N_14830);
or U14977 (N_14977,N_14853,N_14753);
nand U14978 (N_14978,N_14829,N_14816);
and U14979 (N_14979,N_14842,N_14753);
nor U14980 (N_14980,N_14845,N_14841);
and U14981 (N_14981,N_14849,N_14813);
nand U14982 (N_14982,N_14811,N_14832);
or U14983 (N_14983,N_14827,N_14838);
xor U14984 (N_14984,N_14762,N_14825);
nand U14985 (N_14985,N_14870,N_14848);
nand U14986 (N_14986,N_14767,N_14783);
nand U14987 (N_14987,N_14775,N_14805);
nand U14988 (N_14988,N_14831,N_14783);
and U14989 (N_14989,N_14872,N_14841);
nor U14990 (N_14990,N_14750,N_14840);
or U14991 (N_14991,N_14869,N_14797);
or U14992 (N_14992,N_14833,N_14794);
and U14993 (N_14993,N_14833,N_14807);
or U14994 (N_14994,N_14752,N_14776);
nand U14995 (N_14995,N_14789,N_14809);
nor U14996 (N_14996,N_14801,N_14854);
and U14997 (N_14997,N_14809,N_14815);
and U14998 (N_14998,N_14849,N_14851);
xnor U14999 (N_14999,N_14829,N_14776);
xor UO_0 (O_0,N_14931,N_14988);
nand UO_1 (O_1,N_14944,N_14939);
xnor UO_2 (O_2,N_14932,N_14911);
nor UO_3 (O_3,N_14930,N_14902);
and UO_4 (O_4,N_14928,N_14904);
and UO_5 (O_5,N_14876,N_14885);
or UO_6 (O_6,N_14884,N_14877);
or UO_7 (O_7,N_14887,N_14990);
or UO_8 (O_8,N_14976,N_14969);
nor UO_9 (O_9,N_14978,N_14905);
or UO_10 (O_10,N_14963,N_14949);
nand UO_11 (O_11,N_14907,N_14878);
xnor UO_12 (O_12,N_14958,N_14897);
or UO_13 (O_13,N_14924,N_14901);
nor UO_14 (O_14,N_14881,N_14968);
or UO_15 (O_15,N_14956,N_14940);
or UO_16 (O_16,N_14955,N_14889);
or UO_17 (O_17,N_14879,N_14964);
xor UO_18 (O_18,N_14993,N_14972);
xor UO_19 (O_19,N_14914,N_14975);
or UO_20 (O_20,N_14883,N_14926);
and UO_21 (O_21,N_14951,N_14945);
nor UO_22 (O_22,N_14893,N_14937);
nor UO_23 (O_23,N_14917,N_14910);
nand UO_24 (O_24,N_14938,N_14986);
and UO_25 (O_25,N_14959,N_14967);
nand UO_26 (O_26,N_14915,N_14891);
xnor UO_27 (O_27,N_14933,N_14935);
nand UO_28 (O_28,N_14906,N_14985);
xor UO_29 (O_29,N_14980,N_14965);
xor UO_30 (O_30,N_14903,N_14983);
nand UO_31 (O_31,N_14888,N_14982);
nand UO_32 (O_32,N_14996,N_14999);
and UO_33 (O_33,N_14941,N_14921);
nor UO_34 (O_34,N_14979,N_14961);
or UO_35 (O_35,N_14957,N_14966);
and UO_36 (O_36,N_14886,N_14908);
nand UO_37 (O_37,N_14991,N_14875);
nor UO_38 (O_38,N_14936,N_14971);
or UO_39 (O_39,N_14987,N_14913);
xnor UO_40 (O_40,N_14948,N_14880);
or UO_41 (O_41,N_14954,N_14890);
and UO_42 (O_42,N_14923,N_14989);
and UO_43 (O_43,N_14953,N_14947);
nor UO_44 (O_44,N_14998,N_14943);
nor UO_45 (O_45,N_14984,N_14920);
nand UO_46 (O_46,N_14919,N_14900);
or UO_47 (O_47,N_14962,N_14973);
xnor UO_48 (O_48,N_14942,N_14981);
nor UO_49 (O_49,N_14896,N_14922);
or UO_50 (O_50,N_14892,N_14970);
or UO_51 (O_51,N_14977,N_14895);
and UO_52 (O_52,N_14918,N_14894);
nor UO_53 (O_53,N_14925,N_14909);
nor UO_54 (O_54,N_14929,N_14952);
nand UO_55 (O_55,N_14912,N_14960);
and UO_56 (O_56,N_14898,N_14899);
or UO_57 (O_57,N_14934,N_14995);
or UO_58 (O_58,N_14992,N_14946);
nand UO_59 (O_59,N_14882,N_14997);
and UO_60 (O_60,N_14916,N_14927);
and UO_61 (O_61,N_14974,N_14994);
or UO_62 (O_62,N_14950,N_14938);
and UO_63 (O_63,N_14967,N_14878);
or UO_64 (O_64,N_14912,N_14916);
or UO_65 (O_65,N_14880,N_14957);
and UO_66 (O_66,N_14942,N_14890);
nand UO_67 (O_67,N_14887,N_14983);
xnor UO_68 (O_68,N_14945,N_14974);
nand UO_69 (O_69,N_14912,N_14931);
or UO_70 (O_70,N_14902,N_14979);
xor UO_71 (O_71,N_14897,N_14887);
nand UO_72 (O_72,N_14993,N_14960);
and UO_73 (O_73,N_14885,N_14899);
and UO_74 (O_74,N_14977,N_14997);
xnor UO_75 (O_75,N_14922,N_14882);
or UO_76 (O_76,N_14894,N_14959);
xor UO_77 (O_77,N_14997,N_14883);
xnor UO_78 (O_78,N_14971,N_14981);
or UO_79 (O_79,N_14983,N_14910);
nand UO_80 (O_80,N_14883,N_14974);
and UO_81 (O_81,N_14932,N_14984);
nand UO_82 (O_82,N_14899,N_14927);
and UO_83 (O_83,N_14920,N_14887);
nand UO_84 (O_84,N_14949,N_14915);
nor UO_85 (O_85,N_14935,N_14938);
xnor UO_86 (O_86,N_14969,N_14965);
and UO_87 (O_87,N_14981,N_14884);
xnor UO_88 (O_88,N_14922,N_14934);
or UO_89 (O_89,N_14896,N_14951);
xor UO_90 (O_90,N_14894,N_14998);
and UO_91 (O_91,N_14896,N_14910);
and UO_92 (O_92,N_14955,N_14877);
nand UO_93 (O_93,N_14894,N_14972);
nor UO_94 (O_94,N_14928,N_14923);
and UO_95 (O_95,N_14987,N_14966);
xor UO_96 (O_96,N_14990,N_14992);
and UO_97 (O_97,N_14944,N_14915);
xor UO_98 (O_98,N_14979,N_14929);
xor UO_99 (O_99,N_14984,N_14909);
and UO_100 (O_100,N_14984,N_14941);
or UO_101 (O_101,N_14933,N_14945);
nand UO_102 (O_102,N_14889,N_14887);
nor UO_103 (O_103,N_14886,N_14884);
xor UO_104 (O_104,N_14891,N_14984);
and UO_105 (O_105,N_14949,N_14988);
xnor UO_106 (O_106,N_14937,N_14878);
and UO_107 (O_107,N_14993,N_14875);
xor UO_108 (O_108,N_14905,N_14926);
xnor UO_109 (O_109,N_14889,N_14964);
nand UO_110 (O_110,N_14886,N_14921);
nand UO_111 (O_111,N_14936,N_14973);
or UO_112 (O_112,N_14878,N_14888);
xor UO_113 (O_113,N_14950,N_14915);
nand UO_114 (O_114,N_14892,N_14879);
nand UO_115 (O_115,N_14993,N_14937);
or UO_116 (O_116,N_14969,N_14893);
or UO_117 (O_117,N_14913,N_14956);
xor UO_118 (O_118,N_14926,N_14936);
xnor UO_119 (O_119,N_14919,N_14878);
xor UO_120 (O_120,N_14992,N_14924);
nand UO_121 (O_121,N_14901,N_14885);
nand UO_122 (O_122,N_14918,N_14932);
nor UO_123 (O_123,N_14936,N_14993);
nor UO_124 (O_124,N_14909,N_14924);
nor UO_125 (O_125,N_14904,N_14921);
or UO_126 (O_126,N_14914,N_14973);
and UO_127 (O_127,N_14883,N_14897);
nand UO_128 (O_128,N_14904,N_14877);
nand UO_129 (O_129,N_14892,N_14933);
or UO_130 (O_130,N_14997,N_14903);
nand UO_131 (O_131,N_14968,N_14892);
or UO_132 (O_132,N_14936,N_14891);
nor UO_133 (O_133,N_14977,N_14920);
nand UO_134 (O_134,N_14976,N_14883);
and UO_135 (O_135,N_14942,N_14886);
xnor UO_136 (O_136,N_14913,N_14877);
nor UO_137 (O_137,N_14894,N_14913);
nor UO_138 (O_138,N_14887,N_14914);
nand UO_139 (O_139,N_14875,N_14881);
nand UO_140 (O_140,N_14971,N_14944);
nor UO_141 (O_141,N_14924,N_14995);
xnor UO_142 (O_142,N_14960,N_14896);
or UO_143 (O_143,N_14907,N_14996);
and UO_144 (O_144,N_14885,N_14987);
or UO_145 (O_145,N_14895,N_14938);
nor UO_146 (O_146,N_14956,N_14925);
or UO_147 (O_147,N_14935,N_14878);
and UO_148 (O_148,N_14906,N_14898);
and UO_149 (O_149,N_14882,N_14949);
nand UO_150 (O_150,N_14943,N_14988);
nand UO_151 (O_151,N_14938,N_14982);
xor UO_152 (O_152,N_14922,N_14926);
nor UO_153 (O_153,N_14941,N_14944);
xnor UO_154 (O_154,N_14891,N_14919);
nor UO_155 (O_155,N_14940,N_14979);
and UO_156 (O_156,N_14898,N_14918);
nor UO_157 (O_157,N_14940,N_14876);
nand UO_158 (O_158,N_14966,N_14971);
or UO_159 (O_159,N_14916,N_14933);
xor UO_160 (O_160,N_14971,N_14876);
nand UO_161 (O_161,N_14939,N_14989);
nand UO_162 (O_162,N_14985,N_14919);
or UO_163 (O_163,N_14949,N_14984);
and UO_164 (O_164,N_14982,N_14964);
nand UO_165 (O_165,N_14979,N_14965);
xnor UO_166 (O_166,N_14911,N_14991);
xor UO_167 (O_167,N_14907,N_14979);
xor UO_168 (O_168,N_14943,N_14877);
xor UO_169 (O_169,N_14927,N_14909);
nor UO_170 (O_170,N_14952,N_14993);
xor UO_171 (O_171,N_14938,N_14975);
or UO_172 (O_172,N_14964,N_14929);
and UO_173 (O_173,N_14920,N_14949);
and UO_174 (O_174,N_14960,N_14976);
nand UO_175 (O_175,N_14990,N_14989);
xnor UO_176 (O_176,N_14916,N_14997);
xnor UO_177 (O_177,N_14875,N_14912);
or UO_178 (O_178,N_14880,N_14951);
nor UO_179 (O_179,N_14994,N_14956);
nor UO_180 (O_180,N_14946,N_14901);
nor UO_181 (O_181,N_14907,N_14985);
and UO_182 (O_182,N_14957,N_14962);
xor UO_183 (O_183,N_14876,N_14942);
xnor UO_184 (O_184,N_14888,N_14939);
or UO_185 (O_185,N_14954,N_14977);
and UO_186 (O_186,N_14989,N_14987);
nor UO_187 (O_187,N_14906,N_14934);
nor UO_188 (O_188,N_14928,N_14877);
or UO_189 (O_189,N_14972,N_14911);
or UO_190 (O_190,N_14942,N_14884);
or UO_191 (O_191,N_14922,N_14951);
nand UO_192 (O_192,N_14949,N_14905);
xor UO_193 (O_193,N_14976,N_14988);
or UO_194 (O_194,N_14980,N_14918);
and UO_195 (O_195,N_14966,N_14907);
nand UO_196 (O_196,N_14938,N_14984);
and UO_197 (O_197,N_14900,N_14941);
nand UO_198 (O_198,N_14980,N_14937);
xnor UO_199 (O_199,N_14914,N_14909);
and UO_200 (O_200,N_14949,N_14892);
nand UO_201 (O_201,N_14949,N_14911);
and UO_202 (O_202,N_14904,N_14981);
nand UO_203 (O_203,N_14998,N_14983);
nor UO_204 (O_204,N_14968,N_14988);
nor UO_205 (O_205,N_14967,N_14902);
and UO_206 (O_206,N_14879,N_14899);
xor UO_207 (O_207,N_14973,N_14924);
or UO_208 (O_208,N_14963,N_14959);
xnor UO_209 (O_209,N_14923,N_14880);
nor UO_210 (O_210,N_14930,N_14932);
nor UO_211 (O_211,N_14986,N_14907);
xnor UO_212 (O_212,N_14983,N_14971);
and UO_213 (O_213,N_14907,N_14905);
xnor UO_214 (O_214,N_14981,N_14954);
or UO_215 (O_215,N_14948,N_14910);
and UO_216 (O_216,N_14939,N_14955);
xor UO_217 (O_217,N_14909,N_14944);
and UO_218 (O_218,N_14946,N_14985);
xnor UO_219 (O_219,N_14989,N_14880);
or UO_220 (O_220,N_14954,N_14998);
and UO_221 (O_221,N_14890,N_14983);
nand UO_222 (O_222,N_14932,N_14993);
or UO_223 (O_223,N_14903,N_14976);
xor UO_224 (O_224,N_14982,N_14948);
nand UO_225 (O_225,N_14940,N_14937);
and UO_226 (O_226,N_14884,N_14919);
xnor UO_227 (O_227,N_14927,N_14968);
and UO_228 (O_228,N_14878,N_14987);
nor UO_229 (O_229,N_14944,N_14884);
or UO_230 (O_230,N_14889,N_14900);
and UO_231 (O_231,N_14946,N_14911);
or UO_232 (O_232,N_14944,N_14947);
nand UO_233 (O_233,N_14914,N_14956);
nand UO_234 (O_234,N_14936,N_14945);
nor UO_235 (O_235,N_14983,N_14957);
and UO_236 (O_236,N_14975,N_14949);
or UO_237 (O_237,N_14897,N_14921);
nor UO_238 (O_238,N_14885,N_14954);
nor UO_239 (O_239,N_14911,N_14994);
or UO_240 (O_240,N_14901,N_14984);
or UO_241 (O_241,N_14918,N_14976);
and UO_242 (O_242,N_14910,N_14920);
xor UO_243 (O_243,N_14932,N_14890);
and UO_244 (O_244,N_14982,N_14942);
and UO_245 (O_245,N_14989,N_14977);
and UO_246 (O_246,N_14895,N_14909);
or UO_247 (O_247,N_14895,N_14970);
or UO_248 (O_248,N_14887,N_14976);
and UO_249 (O_249,N_14977,N_14902);
and UO_250 (O_250,N_14964,N_14959);
xor UO_251 (O_251,N_14979,N_14969);
nand UO_252 (O_252,N_14980,N_14878);
nand UO_253 (O_253,N_14896,N_14921);
nand UO_254 (O_254,N_14930,N_14922);
nand UO_255 (O_255,N_14924,N_14972);
xor UO_256 (O_256,N_14970,N_14952);
and UO_257 (O_257,N_14912,N_14970);
and UO_258 (O_258,N_14969,N_14978);
xnor UO_259 (O_259,N_14982,N_14978);
nand UO_260 (O_260,N_14886,N_14986);
and UO_261 (O_261,N_14945,N_14931);
nand UO_262 (O_262,N_14890,N_14949);
xnor UO_263 (O_263,N_14907,N_14977);
nor UO_264 (O_264,N_14947,N_14913);
and UO_265 (O_265,N_14903,N_14896);
nor UO_266 (O_266,N_14876,N_14910);
and UO_267 (O_267,N_14964,N_14958);
and UO_268 (O_268,N_14901,N_14876);
nor UO_269 (O_269,N_14936,N_14907);
or UO_270 (O_270,N_14902,N_14953);
xor UO_271 (O_271,N_14936,N_14898);
xnor UO_272 (O_272,N_14918,N_14933);
nand UO_273 (O_273,N_14989,N_14944);
or UO_274 (O_274,N_14950,N_14972);
xor UO_275 (O_275,N_14949,N_14933);
nand UO_276 (O_276,N_14983,N_14939);
or UO_277 (O_277,N_14946,N_14934);
nor UO_278 (O_278,N_14978,N_14914);
or UO_279 (O_279,N_14937,N_14939);
nand UO_280 (O_280,N_14955,N_14966);
nor UO_281 (O_281,N_14946,N_14893);
nand UO_282 (O_282,N_14910,N_14930);
and UO_283 (O_283,N_14968,N_14930);
nor UO_284 (O_284,N_14951,N_14985);
and UO_285 (O_285,N_14880,N_14907);
xnor UO_286 (O_286,N_14942,N_14987);
or UO_287 (O_287,N_14876,N_14884);
and UO_288 (O_288,N_14967,N_14957);
or UO_289 (O_289,N_14901,N_14992);
nand UO_290 (O_290,N_14875,N_14946);
nor UO_291 (O_291,N_14893,N_14895);
xnor UO_292 (O_292,N_14892,N_14998);
xnor UO_293 (O_293,N_14923,N_14919);
or UO_294 (O_294,N_14975,N_14925);
nand UO_295 (O_295,N_14892,N_14952);
and UO_296 (O_296,N_14999,N_14892);
nand UO_297 (O_297,N_14985,N_14999);
and UO_298 (O_298,N_14925,N_14883);
and UO_299 (O_299,N_14957,N_14931);
or UO_300 (O_300,N_14904,N_14930);
xnor UO_301 (O_301,N_14879,N_14955);
xnor UO_302 (O_302,N_14929,N_14890);
nor UO_303 (O_303,N_14972,N_14962);
nor UO_304 (O_304,N_14971,N_14999);
xor UO_305 (O_305,N_14888,N_14976);
nor UO_306 (O_306,N_14965,N_14877);
and UO_307 (O_307,N_14967,N_14903);
nor UO_308 (O_308,N_14938,N_14909);
xor UO_309 (O_309,N_14983,N_14927);
xor UO_310 (O_310,N_14917,N_14909);
xor UO_311 (O_311,N_14985,N_14898);
nor UO_312 (O_312,N_14880,N_14914);
and UO_313 (O_313,N_14974,N_14980);
nand UO_314 (O_314,N_14881,N_14990);
nand UO_315 (O_315,N_14956,N_14999);
nor UO_316 (O_316,N_14962,N_14965);
xnor UO_317 (O_317,N_14949,N_14893);
xor UO_318 (O_318,N_14948,N_14897);
xnor UO_319 (O_319,N_14919,N_14876);
xnor UO_320 (O_320,N_14950,N_14924);
or UO_321 (O_321,N_14963,N_14947);
nand UO_322 (O_322,N_14938,N_14981);
and UO_323 (O_323,N_14987,N_14917);
xor UO_324 (O_324,N_14959,N_14896);
nor UO_325 (O_325,N_14949,N_14924);
nor UO_326 (O_326,N_14933,N_14898);
or UO_327 (O_327,N_14943,N_14933);
nor UO_328 (O_328,N_14975,N_14984);
or UO_329 (O_329,N_14987,N_14965);
or UO_330 (O_330,N_14943,N_14997);
xor UO_331 (O_331,N_14899,N_14991);
or UO_332 (O_332,N_14876,N_14987);
nor UO_333 (O_333,N_14930,N_14980);
nand UO_334 (O_334,N_14986,N_14898);
nor UO_335 (O_335,N_14958,N_14911);
nor UO_336 (O_336,N_14949,N_14921);
nor UO_337 (O_337,N_14887,N_14918);
or UO_338 (O_338,N_14979,N_14941);
and UO_339 (O_339,N_14961,N_14958);
xor UO_340 (O_340,N_14891,N_14928);
nor UO_341 (O_341,N_14936,N_14910);
nor UO_342 (O_342,N_14888,N_14943);
xor UO_343 (O_343,N_14967,N_14950);
nand UO_344 (O_344,N_14877,N_14997);
nand UO_345 (O_345,N_14940,N_14913);
or UO_346 (O_346,N_14929,N_14920);
nand UO_347 (O_347,N_14946,N_14919);
or UO_348 (O_348,N_14895,N_14898);
nor UO_349 (O_349,N_14920,N_14958);
or UO_350 (O_350,N_14885,N_14897);
or UO_351 (O_351,N_14928,N_14998);
and UO_352 (O_352,N_14943,N_14940);
nor UO_353 (O_353,N_14892,N_14943);
and UO_354 (O_354,N_14917,N_14883);
nand UO_355 (O_355,N_14970,N_14984);
nor UO_356 (O_356,N_14916,N_14985);
nand UO_357 (O_357,N_14965,N_14941);
nand UO_358 (O_358,N_14922,N_14944);
nor UO_359 (O_359,N_14986,N_14965);
or UO_360 (O_360,N_14952,N_14878);
nand UO_361 (O_361,N_14934,N_14939);
nand UO_362 (O_362,N_14911,N_14891);
or UO_363 (O_363,N_14959,N_14919);
or UO_364 (O_364,N_14886,N_14997);
nor UO_365 (O_365,N_14905,N_14919);
and UO_366 (O_366,N_14891,N_14893);
or UO_367 (O_367,N_14985,N_14933);
xor UO_368 (O_368,N_14930,N_14885);
or UO_369 (O_369,N_14916,N_14891);
nand UO_370 (O_370,N_14901,N_14920);
nor UO_371 (O_371,N_14926,N_14928);
or UO_372 (O_372,N_14998,N_14976);
xor UO_373 (O_373,N_14922,N_14995);
and UO_374 (O_374,N_14994,N_14941);
nor UO_375 (O_375,N_14943,N_14878);
nor UO_376 (O_376,N_14903,N_14913);
nor UO_377 (O_377,N_14968,N_14891);
nor UO_378 (O_378,N_14908,N_14881);
or UO_379 (O_379,N_14936,N_14897);
or UO_380 (O_380,N_14925,N_14966);
nor UO_381 (O_381,N_14977,N_14952);
or UO_382 (O_382,N_14875,N_14894);
nor UO_383 (O_383,N_14988,N_14891);
xnor UO_384 (O_384,N_14910,N_14976);
nor UO_385 (O_385,N_14905,N_14957);
and UO_386 (O_386,N_14924,N_14964);
nor UO_387 (O_387,N_14946,N_14999);
xor UO_388 (O_388,N_14987,N_14936);
nor UO_389 (O_389,N_14983,N_14940);
and UO_390 (O_390,N_14964,N_14947);
xor UO_391 (O_391,N_14891,N_14997);
and UO_392 (O_392,N_14886,N_14982);
nand UO_393 (O_393,N_14878,N_14940);
or UO_394 (O_394,N_14965,N_14985);
xnor UO_395 (O_395,N_14882,N_14906);
nand UO_396 (O_396,N_14986,N_14884);
nor UO_397 (O_397,N_14914,N_14924);
nor UO_398 (O_398,N_14985,N_14905);
and UO_399 (O_399,N_14970,N_14882);
and UO_400 (O_400,N_14914,N_14995);
or UO_401 (O_401,N_14998,N_14951);
xnor UO_402 (O_402,N_14884,N_14915);
and UO_403 (O_403,N_14947,N_14907);
and UO_404 (O_404,N_14916,N_14911);
xor UO_405 (O_405,N_14979,N_14919);
nor UO_406 (O_406,N_14922,N_14939);
or UO_407 (O_407,N_14968,N_14902);
or UO_408 (O_408,N_14993,N_14997);
and UO_409 (O_409,N_14921,N_14917);
nand UO_410 (O_410,N_14893,N_14901);
nand UO_411 (O_411,N_14992,N_14899);
nand UO_412 (O_412,N_14932,N_14968);
and UO_413 (O_413,N_14887,N_14924);
nor UO_414 (O_414,N_14976,N_14902);
nand UO_415 (O_415,N_14939,N_14974);
nor UO_416 (O_416,N_14879,N_14940);
xnor UO_417 (O_417,N_14980,N_14912);
nor UO_418 (O_418,N_14949,N_14909);
nand UO_419 (O_419,N_14944,N_14943);
nand UO_420 (O_420,N_14910,N_14921);
xor UO_421 (O_421,N_14950,N_14885);
xor UO_422 (O_422,N_14955,N_14881);
nand UO_423 (O_423,N_14910,N_14927);
xor UO_424 (O_424,N_14883,N_14963);
nand UO_425 (O_425,N_14912,N_14983);
and UO_426 (O_426,N_14898,N_14915);
and UO_427 (O_427,N_14949,N_14961);
nor UO_428 (O_428,N_14890,N_14934);
nand UO_429 (O_429,N_14890,N_14948);
xnor UO_430 (O_430,N_14951,N_14965);
and UO_431 (O_431,N_14949,N_14925);
or UO_432 (O_432,N_14932,N_14958);
nand UO_433 (O_433,N_14882,N_14886);
xor UO_434 (O_434,N_14945,N_14995);
or UO_435 (O_435,N_14931,N_14977);
nand UO_436 (O_436,N_14929,N_14981);
nor UO_437 (O_437,N_14915,N_14880);
and UO_438 (O_438,N_14888,N_14914);
nor UO_439 (O_439,N_14893,N_14923);
nor UO_440 (O_440,N_14884,N_14909);
xnor UO_441 (O_441,N_14919,N_14913);
and UO_442 (O_442,N_14938,N_14928);
xnor UO_443 (O_443,N_14950,N_14991);
or UO_444 (O_444,N_14944,N_14906);
or UO_445 (O_445,N_14933,N_14896);
or UO_446 (O_446,N_14963,N_14933);
xor UO_447 (O_447,N_14892,N_14953);
or UO_448 (O_448,N_14892,N_14947);
and UO_449 (O_449,N_14987,N_14902);
nor UO_450 (O_450,N_14947,N_14926);
and UO_451 (O_451,N_14992,N_14890);
nor UO_452 (O_452,N_14949,N_14897);
nor UO_453 (O_453,N_14902,N_14934);
or UO_454 (O_454,N_14887,N_14946);
nor UO_455 (O_455,N_14970,N_14953);
or UO_456 (O_456,N_14982,N_14979);
or UO_457 (O_457,N_14882,N_14895);
and UO_458 (O_458,N_14989,N_14960);
or UO_459 (O_459,N_14964,N_14940);
nand UO_460 (O_460,N_14923,N_14969);
or UO_461 (O_461,N_14991,N_14993);
nand UO_462 (O_462,N_14932,N_14902);
and UO_463 (O_463,N_14972,N_14932);
or UO_464 (O_464,N_14985,N_14924);
and UO_465 (O_465,N_14907,N_14937);
or UO_466 (O_466,N_14929,N_14957);
and UO_467 (O_467,N_14891,N_14940);
and UO_468 (O_468,N_14926,N_14975);
xnor UO_469 (O_469,N_14933,N_14965);
xor UO_470 (O_470,N_14966,N_14964);
or UO_471 (O_471,N_14898,N_14926);
nor UO_472 (O_472,N_14972,N_14970);
nor UO_473 (O_473,N_14908,N_14981);
nor UO_474 (O_474,N_14986,N_14990);
nand UO_475 (O_475,N_14900,N_14938);
xor UO_476 (O_476,N_14991,N_14923);
nor UO_477 (O_477,N_14993,N_14929);
xor UO_478 (O_478,N_14947,N_14895);
nor UO_479 (O_479,N_14916,N_14878);
or UO_480 (O_480,N_14939,N_14948);
and UO_481 (O_481,N_14981,N_14902);
nand UO_482 (O_482,N_14961,N_14929);
nor UO_483 (O_483,N_14942,N_14948);
or UO_484 (O_484,N_14941,N_14940);
xor UO_485 (O_485,N_14923,N_14929);
and UO_486 (O_486,N_14985,N_14925);
nand UO_487 (O_487,N_14990,N_14941);
nor UO_488 (O_488,N_14928,N_14956);
nor UO_489 (O_489,N_14897,N_14924);
or UO_490 (O_490,N_14978,N_14998);
nand UO_491 (O_491,N_14940,N_14890);
nor UO_492 (O_492,N_14969,N_14990);
nand UO_493 (O_493,N_14891,N_14939);
and UO_494 (O_494,N_14877,N_14951);
nand UO_495 (O_495,N_14948,N_14972);
or UO_496 (O_496,N_14953,N_14950);
nand UO_497 (O_497,N_14891,N_14932);
xor UO_498 (O_498,N_14882,N_14950);
or UO_499 (O_499,N_14968,N_14877);
nor UO_500 (O_500,N_14990,N_14915);
and UO_501 (O_501,N_14933,N_14957);
nor UO_502 (O_502,N_14968,N_14964);
and UO_503 (O_503,N_14959,N_14907);
xor UO_504 (O_504,N_14935,N_14916);
and UO_505 (O_505,N_14939,N_14981);
xor UO_506 (O_506,N_14981,N_14926);
nor UO_507 (O_507,N_14981,N_14878);
nand UO_508 (O_508,N_14987,N_14945);
and UO_509 (O_509,N_14875,N_14919);
or UO_510 (O_510,N_14939,N_14882);
and UO_511 (O_511,N_14971,N_14925);
xnor UO_512 (O_512,N_14934,N_14915);
and UO_513 (O_513,N_14875,N_14898);
and UO_514 (O_514,N_14959,N_14893);
nor UO_515 (O_515,N_14941,N_14951);
or UO_516 (O_516,N_14970,N_14909);
xnor UO_517 (O_517,N_14876,N_14887);
and UO_518 (O_518,N_14962,N_14922);
nor UO_519 (O_519,N_14910,N_14986);
xor UO_520 (O_520,N_14930,N_14979);
or UO_521 (O_521,N_14999,N_14994);
nand UO_522 (O_522,N_14993,N_14894);
and UO_523 (O_523,N_14900,N_14975);
xnor UO_524 (O_524,N_14992,N_14972);
and UO_525 (O_525,N_14937,N_14899);
nand UO_526 (O_526,N_14925,N_14939);
or UO_527 (O_527,N_14879,N_14990);
and UO_528 (O_528,N_14950,N_14946);
and UO_529 (O_529,N_14939,N_14912);
xor UO_530 (O_530,N_14896,N_14887);
or UO_531 (O_531,N_14921,N_14912);
or UO_532 (O_532,N_14947,N_14966);
and UO_533 (O_533,N_14970,N_14990);
nand UO_534 (O_534,N_14993,N_14968);
nand UO_535 (O_535,N_14884,N_14890);
and UO_536 (O_536,N_14974,N_14940);
xor UO_537 (O_537,N_14891,N_14938);
xnor UO_538 (O_538,N_14905,N_14943);
and UO_539 (O_539,N_14975,N_14959);
nor UO_540 (O_540,N_14975,N_14896);
or UO_541 (O_541,N_14977,N_14933);
xor UO_542 (O_542,N_14890,N_14938);
nand UO_543 (O_543,N_14886,N_14878);
or UO_544 (O_544,N_14980,N_14968);
xor UO_545 (O_545,N_14902,N_14890);
and UO_546 (O_546,N_14969,N_14891);
xnor UO_547 (O_547,N_14925,N_14897);
nand UO_548 (O_548,N_14922,N_14971);
and UO_549 (O_549,N_14930,N_14997);
nand UO_550 (O_550,N_14968,N_14958);
xnor UO_551 (O_551,N_14933,N_14953);
or UO_552 (O_552,N_14902,N_14978);
and UO_553 (O_553,N_14892,N_14979);
xnor UO_554 (O_554,N_14975,N_14972);
or UO_555 (O_555,N_14949,N_14877);
nor UO_556 (O_556,N_14898,N_14949);
or UO_557 (O_557,N_14918,N_14975);
nand UO_558 (O_558,N_14996,N_14963);
xnor UO_559 (O_559,N_14934,N_14971);
xnor UO_560 (O_560,N_14916,N_14977);
nand UO_561 (O_561,N_14975,N_14936);
xnor UO_562 (O_562,N_14926,N_14937);
nor UO_563 (O_563,N_14876,N_14896);
or UO_564 (O_564,N_14980,N_14907);
nand UO_565 (O_565,N_14909,N_14977);
and UO_566 (O_566,N_14944,N_14928);
and UO_567 (O_567,N_14944,N_14991);
or UO_568 (O_568,N_14878,N_14958);
nor UO_569 (O_569,N_14988,N_14898);
nor UO_570 (O_570,N_14915,N_14982);
xor UO_571 (O_571,N_14940,N_14985);
nand UO_572 (O_572,N_14975,N_14960);
nand UO_573 (O_573,N_14895,N_14897);
nand UO_574 (O_574,N_14969,N_14994);
nor UO_575 (O_575,N_14906,N_14891);
nand UO_576 (O_576,N_14936,N_14948);
and UO_577 (O_577,N_14943,N_14966);
nand UO_578 (O_578,N_14878,N_14914);
or UO_579 (O_579,N_14942,N_14901);
and UO_580 (O_580,N_14965,N_14913);
and UO_581 (O_581,N_14979,N_14908);
nand UO_582 (O_582,N_14970,N_14926);
xor UO_583 (O_583,N_14981,N_14915);
xnor UO_584 (O_584,N_14985,N_14984);
xor UO_585 (O_585,N_14900,N_14907);
nor UO_586 (O_586,N_14966,N_14900);
nand UO_587 (O_587,N_14920,N_14952);
nand UO_588 (O_588,N_14995,N_14889);
or UO_589 (O_589,N_14908,N_14980);
nand UO_590 (O_590,N_14920,N_14911);
or UO_591 (O_591,N_14910,N_14912);
nand UO_592 (O_592,N_14985,N_14892);
nand UO_593 (O_593,N_14955,N_14876);
xor UO_594 (O_594,N_14998,N_14988);
nand UO_595 (O_595,N_14995,N_14908);
xnor UO_596 (O_596,N_14952,N_14985);
or UO_597 (O_597,N_14880,N_14947);
or UO_598 (O_598,N_14880,N_14889);
nor UO_599 (O_599,N_14991,N_14942);
and UO_600 (O_600,N_14967,N_14921);
or UO_601 (O_601,N_14976,N_14917);
and UO_602 (O_602,N_14887,N_14948);
and UO_603 (O_603,N_14988,N_14951);
nand UO_604 (O_604,N_14897,N_14899);
nor UO_605 (O_605,N_14924,N_14989);
nand UO_606 (O_606,N_14971,N_14905);
or UO_607 (O_607,N_14919,N_14972);
xnor UO_608 (O_608,N_14981,N_14941);
nor UO_609 (O_609,N_14928,N_14913);
and UO_610 (O_610,N_14927,N_14991);
nand UO_611 (O_611,N_14936,N_14912);
nor UO_612 (O_612,N_14964,N_14960);
nand UO_613 (O_613,N_14890,N_14878);
and UO_614 (O_614,N_14933,N_14962);
or UO_615 (O_615,N_14939,N_14901);
and UO_616 (O_616,N_14974,N_14912);
nand UO_617 (O_617,N_14970,N_14876);
and UO_618 (O_618,N_14881,N_14947);
nand UO_619 (O_619,N_14888,N_14945);
or UO_620 (O_620,N_14953,N_14881);
nand UO_621 (O_621,N_14969,N_14943);
nor UO_622 (O_622,N_14889,N_14890);
xor UO_623 (O_623,N_14928,N_14884);
or UO_624 (O_624,N_14966,N_14915);
xnor UO_625 (O_625,N_14877,N_14977);
and UO_626 (O_626,N_14962,N_14980);
or UO_627 (O_627,N_14890,N_14930);
or UO_628 (O_628,N_14965,N_14880);
or UO_629 (O_629,N_14962,N_14943);
nor UO_630 (O_630,N_14916,N_14950);
nor UO_631 (O_631,N_14987,N_14998);
xnor UO_632 (O_632,N_14945,N_14906);
and UO_633 (O_633,N_14928,N_14901);
and UO_634 (O_634,N_14963,N_14920);
and UO_635 (O_635,N_14888,N_14884);
and UO_636 (O_636,N_14950,N_14904);
or UO_637 (O_637,N_14997,N_14946);
nand UO_638 (O_638,N_14911,N_14963);
nor UO_639 (O_639,N_14931,N_14955);
nor UO_640 (O_640,N_14918,N_14889);
or UO_641 (O_641,N_14984,N_14990);
nor UO_642 (O_642,N_14893,N_14882);
nor UO_643 (O_643,N_14930,N_14878);
nand UO_644 (O_644,N_14956,N_14887);
nor UO_645 (O_645,N_14998,N_14910);
or UO_646 (O_646,N_14919,N_14971);
and UO_647 (O_647,N_14993,N_14916);
or UO_648 (O_648,N_14963,N_14971);
xnor UO_649 (O_649,N_14892,N_14930);
and UO_650 (O_650,N_14959,N_14962);
xor UO_651 (O_651,N_14905,N_14955);
nor UO_652 (O_652,N_14894,N_14876);
and UO_653 (O_653,N_14880,N_14924);
and UO_654 (O_654,N_14906,N_14939);
or UO_655 (O_655,N_14987,N_14927);
nand UO_656 (O_656,N_14983,N_14967);
and UO_657 (O_657,N_14902,N_14997);
nor UO_658 (O_658,N_14933,N_14921);
or UO_659 (O_659,N_14960,N_14898);
xnor UO_660 (O_660,N_14903,N_14939);
xor UO_661 (O_661,N_14910,N_14947);
or UO_662 (O_662,N_14877,N_14969);
or UO_663 (O_663,N_14974,N_14922);
xor UO_664 (O_664,N_14974,N_14917);
or UO_665 (O_665,N_14973,N_14904);
nand UO_666 (O_666,N_14899,N_14930);
nand UO_667 (O_667,N_14995,N_14962);
xor UO_668 (O_668,N_14977,N_14922);
or UO_669 (O_669,N_14961,N_14886);
and UO_670 (O_670,N_14915,N_14883);
nor UO_671 (O_671,N_14950,N_14952);
or UO_672 (O_672,N_14955,N_14998);
xnor UO_673 (O_673,N_14905,N_14963);
nand UO_674 (O_674,N_14996,N_14959);
and UO_675 (O_675,N_14881,N_14978);
xnor UO_676 (O_676,N_14947,N_14942);
xnor UO_677 (O_677,N_14886,N_14934);
nand UO_678 (O_678,N_14899,N_14967);
and UO_679 (O_679,N_14909,N_14883);
xnor UO_680 (O_680,N_14953,N_14993);
and UO_681 (O_681,N_14926,N_14920);
and UO_682 (O_682,N_14942,N_14983);
nor UO_683 (O_683,N_14970,N_14996);
or UO_684 (O_684,N_14979,N_14955);
or UO_685 (O_685,N_14941,N_14958);
or UO_686 (O_686,N_14974,N_14942);
xnor UO_687 (O_687,N_14903,N_14917);
xnor UO_688 (O_688,N_14972,N_14900);
xnor UO_689 (O_689,N_14944,N_14885);
or UO_690 (O_690,N_14899,N_14888);
xnor UO_691 (O_691,N_14964,N_14895);
xnor UO_692 (O_692,N_14926,N_14915);
nor UO_693 (O_693,N_14939,N_14914);
or UO_694 (O_694,N_14968,N_14975);
nand UO_695 (O_695,N_14994,N_14899);
xnor UO_696 (O_696,N_14883,N_14986);
and UO_697 (O_697,N_14881,N_14963);
nor UO_698 (O_698,N_14938,N_14998);
and UO_699 (O_699,N_14964,N_14957);
nor UO_700 (O_700,N_14875,N_14968);
nand UO_701 (O_701,N_14934,N_14879);
or UO_702 (O_702,N_14884,N_14933);
nor UO_703 (O_703,N_14951,N_14924);
nor UO_704 (O_704,N_14983,N_14978);
xnor UO_705 (O_705,N_14909,N_14894);
nor UO_706 (O_706,N_14982,N_14893);
or UO_707 (O_707,N_14996,N_14943);
and UO_708 (O_708,N_14893,N_14935);
nand UO_709 (O_709,N_14917,N_14882);
and UO_710 (O_710,N_14969,N_14916);
or UO_711 (O_711,N_14891,N_14907);
nor UO_712 (O_712,N_14969,N_14934);
and UO_713 (O_713,N_14908,N_14907);
and UO_714 (O_714,N_14975,N_14964);
nand UO_715 (O_715,N_14892,N_14951);
nand UO_716 (O_716,N_14934,N_14897);
xor UO_717 (O_717,N_14878,N_14997);
nor UO_718 (O_718,N_14920,N_14938);
nand UO_719 (O_719,N_14897,N_14915);
xnor UO_720 (O_720,N_14894,N_14945);
nor UO_721 (O_721,N_14930,N_14938);
nand UO_722 (O_722,N_14977,N_14927);
nand UO_723 (O_723,N_14983,N_14953);
xnor UO_724 (O_724,N_14929,N_14968);
or UO_725 (O_725,N_14895,N_14971);
nand UO_726 (O_726,N_14875,N_14981);
or UO_727 (O_727,N_14889,N_14956);
nor UO_728 (O_728,N_14900,N_14933);
or UO_729 (O_729,N_14970,N_14983);
nand UO_730 (O_730,N_14957,N_14943);
xnor UO_731 (O_731,N_14938,N_14956);
or UO_732 (O_732,N_14965,N_14983);
nor UO_733 (O_733,N_14934,N_14996);
or UO_734 (O_734,N_14917,N_14955);
or UO_735 (O_735,N_14900,N_14947);
nand UO_736 (O_736,N_14922,N_14891);
nor UO_737 (O_737,N_14992,N_14940);
or UO_738 (O_738,N_14908,N_14917);
xor UO_739 (O_739,N_14963,N_14909);
and UO_740 (O_740,N_14928,N_14917);
nor UO_741 (O_741,N_14927,N_14947);
xor UO_742 (O_742,N_14944,N_14923);
nand UO_743 (O_743,N_14971,N_14910);
xor UO_744 (O_744,N_14896,N_14977);
and UO_745 (O_745,N_14930,N_14895);
xor UO_746 (O_746,N_14991,N_14907);
nand UO_747 (O_747,N_14895,N_14981);
nor UO_748 (O_748,N_14933,N_14928);
xnor UO_749 (O_749,N_14964,N_14994);
nand UO_750 (O_750,N_14983,N_14919);
nor UO_751 (O_751,N_14890,N_14901);
and UO_752 (O_752,N_14899,N_14877);
nand UO_753 (O_753,N_14911,N_14962);
xor UO_754 (O_754,N_14886,N_14965);
or UO_755 (O_755,N_14970,N_14889);
nor UO_756 (O_756,N_14881,N_14924);
or UO_757 (O_757,N_14936,N_14951);
or UO_758 (O_758,N_14998,N_14959);
and UO_759 (O_759,N_14978,N_14933);
nor UO_760 (O_760,N_14965,N_14888);
nor UO_761 (O_761,N_14891,N_14900);
nor UO_762 (O_762,N_14894,N_14919);
nor UO_763 (O_763,N_14992,N_14983);
nand UO_764 (O_764,N_14964,N_14987);
nor UO_765 (O_765,N_14883,N_14994);
or UO_766 (O_766,N_14988,N_14946);
nor UO_767 (O_767,N_14984,N_14880);
and UO_768 (O_768,N_14939,N_14960);
nor UO_769 (O_769,N_14936,N_14900);
or UO_770 (O_770,N_14949,N_14918);
nor UO_771 (O_771,N_14987,N_14944);
or UO_772 (O_772,N_14988,N_14942);
xnor UO_773 (O_773,N_14939,N_14953);
nand UO_774 (O_774,N_14995,N_14970);
and UO_775 (O_775,N_14902,N_14985);
xor UO_776 (O_776,N_14952,N_14995);
nand UO_777 (O_777,N_14895,N_14998);
or UO_778 (O_778,N_14924,N_14889);
xor UO_779 (O_779,N_14960,N_14900);
and UO_780 (O_780,N_14904,N_14905);
or UO_781 (O_781,N_14980,N_14894);
nand UO_782 (O_782,N_14948,N_14891);
and UO_783 (O_783,N_14978,N_14962);
nand UO_784 (O_784,N_14990,N_14979);
or UO_785 (O_785,N_14936,N_14917);
or UO_786 (O_786,N_14886,N_14918);
nor UO_787 (O_787,N_14883,N_14899);
xor UO_788 (O_788,N_14923,N_14892);
or UO_789 (O_789,N_14947,N_14879);
and UO_790 (O_790,N_14941,N_14931);
nor UO_791 (O_791,N_14928,N_14882);
nand UO_792 (O_792,N_14943,N_14954);
xnor UO_793 (O_793,N_14994,N_14918);
nor UO_794 (O_794,N_14931,N_14970);
nand UO_795 (O_795,N_14918,N_14948);
and UO_796 (O_796,N_14961,N_14953);
and UO_797 (O_797,N_14886,N_14920);
nand UO_798 (O_798,N_14879,N_14875);
nand UO_799 (O_799,N_14930,N_14911);
and UO_800 (O_800,N_14953,N_14932);
and UO_801 (O_801,N_14906,N_14917);
and UO_802 (O_802,N_14980,N_14994);
and UO_803 (O_803,N_14960,N_14970);
and UO_804 (O_804,N_14931,N_14949);
nand UO_805 (O_805,N_14991,N_14919);
nor UO_806 (O_806,N_14954,N_14973);
and UO_807 (O_807,N_14964,N_14884);
and UO_808 (O_808,N_14937,N_14987);
nand UO_809 (O_809,N_14917,N_14893);
or UO_810 (O_810,N_14892,N_14976);
or UO_811 (O_811,N_14878,N_14921);
nand UO_812 (O_812,N_14918,N_14967);
nand UO_813 (O_813,N_14981,N_14945);
nor UO_814 (O_814,N_14950,N_14910);
nor UO_815 (O_815,N_14878,N_14948);
xnor UO_816 (O_816,N_14991,N_14969);
xor UO_817 (O_817,N_14942,N_14915);
nand UO_818 (O_818,N_14964,N_14944);
nand UO_819 (O_819,N_14980,N_14938);
nor UO_820 (O_820,N_14876,N_14900);
xor UO_821 (O_821,N_14891,N_14899);
and UO_822 (O_822,N_14961,N_14916);
xor UO_823 (O_823,N_14940,N_14932);
nand UO_824 (O_824,N_14942,N_14892);
xnor UO_825 (O_825,N_14893,N_14881);
nor UO_826 (O_826,N_14878,N_14978);
or UO_827 (O_827,N_14913,N_14889);
nor UO_828 (O_828,N_14926,N_14958);
nand UO_829 (O_829,N_14943,N_14923);
xnor UO_830 (O_830,N_14959,N_14955);
nor UO_831 (O_831,N_14952,N_14905);
nand UO_832 (O_832,N_14987,N_14957);
or UO_833 (O_833,N_14980,N_14877);
or UO_834 (O_834,N_14972,N_14979);
and UO_835 (O_835,N_14975,N_14889);
xor UO_836 (O_836,N_14922,N_14979);
xor UO_837 (O_837,N_14893,N_14936);
or UO_838 (O_838,N_14980,N_14951);
or UO_839 (O_839,N_14930,N_14985);
and UO_840 (O_840,N_14915,N_14890);
and UO_841 (O_841,N_14982,N_14980);
nand UO_842 (O_842,N_14886,N_14932);
or UO_843 (O_843,N_14966,N_14965);
or UO_844 (O_844,N_14920,N_14925);
and UO_845 (O_845,N_14981,N_14994);
or UO_846 (O_846,N_14887,N_14969);
and UO_847 (O_847,N_14930,N_14970);
nor UO_848 (O_848,N_14880,N_14893);
xor UO_849 (O_849,N_14995,N_14918);
nand UO_850 (O_850,N_14945,N_14940);
or UO_851 (O_851,N_14940,N_14971);
nand UO_852 (O_852,N_14927,N_14904);
or UO_853 (O_853,N_14922,N_14960);
nand UO_854 (O_854,N_14971,N_14962);
nor UO_855 (O_855,N_14917,N_14996);
nand UO_856 (O_856,N_14963,N_14977);
xnor UO_857 (O_857,N_14894,N_14987);
or UO_858 (O_858,N_14939,N_14886);
or UO_859 (O_859,N_14983,N_14948);
or UO_860 (O_860,N_14878,N_14965);
and UO_861 (O_861,N_14939,N_14916);
and UO_862 (O_862,N_14900,N_14934);
nor UO_863 (O_863,N_14989,N_14890);
nor UO_864 (O_864,N_14981,N_14997);
xnor UO_865 (O_865,N_14923,N_14971);
and UO_866 (O_866,N_14931,N_14890);
nand UO_867 (O_867,N_14939,N_14993);
or UO_868 (O_868,N_14971,N_14918);
nand UO_869 (O_869,N_14913,N_14931);
nor UO_870 (O_870,N_14920,N_14968);
and UO_871 (O_871,N_14931,N_14876);
nand UO_872 (O_872,N_14910,N_14908);
xor UO_873 (O_873,N_14886,N_14979);
nor UO_874 (O_874,N_14904,N_14971);
nor UO_875 (O_875,N_14952,N_14953);
nand UO_876 (O_876,N_14990,N_14939);
nand UO_877 (O_877,N_14886,N_14970);
xor UO_878 (O_878,N_14968,N_14977);
xor UO_879 (O_879,N_14990,N_14943);
xor UO_880 (O_880,N_14984,N_14937);
and UO_881 (O_881,N_14910,N_14981);
nand UO_882 (O_882,N_14902,N_14940);
nor UO_883 (O_883,N_14950,N_14926);
or UO_884 (O_884,N_14954,N_14886);
or UO_885 (O_885,N_14902,N_14926);
and UO_886 (O_886,N_14877,N_14902);
nand UO_887 (O_887,N_14920,N_14943);
nand UO_888 (O_888,N_14895,N_14992);
or UO_889 (O_889,N_14964,N_14963);
nor UO_890 (O_890,N_14905,N_14931);
nor UO_891 (O_891,N_14949,N_14966);
nand UO_892 (O_892,N_14972,N_14891);
nor UO_893 (O_893,N_14984,N_14930);
or UO_894 (O_894,N_14980,N_14986);
nand UO_895 (O_895,N_14876,N_14996);
xor UO_896 (O_896,N_14957,N_14896);
and UO_897 (O_897,N_14875,N_14967);
or UO_898 (O_898,N_14955,N_14980);
or UO_899 (O_899,N_14991,N_14966);
and UO_900 (O_900,N_14998,N_14929);
nor UO_901 (O_901,N_14903,N_14909);
nand UO_902 (O_902,N_14977,N_14994);
xor UO_903 (O_903,N_14928,N_14962);
nand UO_904 (O_904,N_14911,N_14913);
and UO_905 (O_905,N_14892,N_14978);
nand UO_906 (O_906,N_14920,N_14992);
nand UO_907 (O_907,N_14965,N_14908);
or UO_908 (O_908,N_14882,N_14907);
xor UO_909 (O_909,N_14946,N_14994);
nand UO_910 (O_910,N_14895,N_14925);
nor UO_911 (O_911,N_14958,N_14992);
and UO_912 (O_912,N_14928,N_14968);
and UO_913 (O_913,N_14962,N_14936);
nor UO_914 (O_914,N_14894,N_14902);
xor UO_915 (O_915,N_14991,N_14901);
nand UO_916 (O_916,N_14929,N_14958);
or UO_917 (O_917,N_14993,N_14892);
or UO_918 (O_918,N_14922,N_14893);
nand UO_919 (O_919,N_14993,N_14887);
or UO_920 (O_920,N_14895,N_14903);
or UO_921 (O_921,N_14976,N_14875);
nor UO_922 (O_922,N_14977,N_14898);
or UO_923 (O_923,N_14995,N_14993);
or UO_924 (O_924,N_14954,N_14947);
xnor UO_925 (O_925,N_14942,N_14912);
nand UO_926 (O_926,N_14890,N_14916);
nand UO_927 (O_927,N_14903,N_14998);
nand UO_928 (O_928,N_14930,N_14978);
and UO_929 (O_929,N_14964,N_14890);
and UO_930 (O_930,N_14907,N_14999);
or UO_931 (O_931,N_14920,N_14922);
and UO_932 (O_932,N_14998,N_14939);
nor UO_933 (O_933,N_14917,N_14958);
nand UO_934 (O_934,N_14906,N_14948);
or UO_935 (O_935,N_14899,N_14908);
xnor UO_936 (O_936,N_14888,N_14959);
and UO_937 (O_937,N_14960,N_14895);
nand UO_938 (O_938,N_14939,N_14887);
xor UO_939 (O_939,N_14945,N_14914);
nand UO_940 (O_940,N_14996,N_14891);
or UO_941 (O_941,N_14905,N_14944);
xnor UO_942 (O_942,N_14929,N_14944);
and UO_943 (O_943,N_14947,N_14923);
nor UO_944 (O_944,N_14912,N_14962);
xnor UO_945 (O_945,N_14901,N_14985);
nor UO_946 (O_946,N_14907,N_14976);
nand UO_947 (O_947,N_14885,N_14974);
xnor UO_948 (O_948,N_14885,N_14917);
xnor UO_949 (O_949,N_14946,N_14981);
xnor UO_950 (O_950,N_14926,N_14998);
xor UO_951 (O_951,N_14986,N_14956);
or UO_952 (O_952,N_14907,N_14950);
nor UO_953 (O_953,N_14933,N_14903);
and UO_954 (O_954,N_14898,N_14943);
nor UO_955 (O_955,N_14918,N_14907);
nand UO_956 (O_956,N_14893,N_14988);
or UO_957 (O_957,N_14951,N_14876);
or UO_958 (O_958,N_14961,N_14980);
nor UO_959 (O_959,N_14937,N_14986);
nor UO_960 (O_960,N_14963,N_14940);
xor UO_961 (O_961,N_14888,N_14912);
nor UO_962 (O_962,N_14881,N_14901);
and UO_963 (O_963,N_14964,N_14914);
xnor UO_964 (O_964,N_14998,N_14896);
xnor UO_965 (O_965,N_14927,N_14903);
or UO_966 (O_966,N_14890,N_14961);
and UO_967 (O_967,N_14933,N_14885);
nand UO_968 (O_968,N_14948,N_14886);
or UO_969 (O_969,N_14900,N_14929);
nand UO_970 (O_970,N_14903,N_14961);
nor UO_971 (O_971,N_14988,N_14989);
nand UO_972 (O_972,N_14883,N_14930);
and UO_973 (O_973,N_14888,N_14967);
xnor UO_974 (O_974,N_14941,N_14896);
nand UO_975 (O_975,N_14911,N_14908);
xnor UO_976 (O_976,N_14893,N_14900);
xor UO_977 (O_977,N_14925,N_14906);
nor UO_978 (O_978,N_14970,N_14901);
nor UO_979 (O_979,N_14985,N_14945);
xnor UO_980 (O_980,N_14976,N_14964);
nand UO_981 (O_981,N_14987,N_14971);
nand UO_982 (O_982,N_14878,N_14900);
nor UO_983 (O_983,N_14990,N_14891);
and UO_984 (O_984,N_14936,N_14941);
or UO_985 (O_985,N_14940,N_14931);
nand UO_986 (O_986,N_14963,N_14930);
nor UO_987 (O_987,N_14881,N_14915);
and UO_988 (O_988,N_14928,N_14941);
nand UO_989 (O_989,N_14950,N_14917);
nor UO_990 (O_990,N_14900,N_14928);
xnor UO_991 (O_991,N_14998,N_14931);
and UO_992 (O_992,N_14944,N_14974);
nor UO_993 (O_993,N_14920,N_14923);
and UO_994 (O_994,N_14957,N_14988);
xor UO_995 (O_995,N_14905,N_14920);
nand UO_996 (O_996,N_14897,N_14995);
nand UO_997 (O_997,N_14953,N_14915);
xnor UO_998 (O_998,N_14966,N_14974);
nor UO_999 (O_999,N_14973,N_14999);
nor UO_1000 (O_1000,N_14997,N_14905);
xor UO_1001 (O_1001,N_14914,N_14913);
and UO_1002 (O_1002,N_14950,N_14921);
nand UO_1003 (O_1003,N_14996,N_14899);
nor UO_1004 (O_1004,N_14990,N_14960);
and UO_1005 (O_1005,N_14915,N_14999);
xnor UO_1006 (O_1006,N_14955,N_14985);
and UO_1007 (O_1007,N_14926,N_14890);
and UO_1008 (O_1008,N_14887,N_14943);
nor UO_1009 (O_1009,N_14933,N_14999);
xnor UO_1010 (O_1010,N_14985,N_14911);
nor UO_1011 (O_1011,N_14996,N_14944);
nand UO_1012 (O_1012,N_14884,N_14900);
or UO_1013 (O_1013,N_14985,N_14983);
xnor UO_1014 (O_1014,N_14966,N_14959);
xnor UO_1015 (O_1015,N_14936,N_14918);
and UO_1016 (O_1016,N_14992,N_14928);
xor UO_1017 (O_1017,N_14928,N_14879);
nor UO_1018 (O_1018,N_14890,N_14956);
nor UO_1019 (O_1019,N_14925,N_14952);
xnor UO_1020 (O_1020,N_14899,N_14954);
nor UO_1021 (O_1021,N_14904,N_14964);
nand UO_1022 (O_1022,N_14881,N_14958);
or UO_1023 (O_1023,N_14969,N_14926);
and UO_1024 (O_1024,N_14965,N_14974);
and UO_1025 (O_1025,N_14889,N_14974);
nand UO_1026 (O_1026,N_14965,N_14943);
nor UO_1027 (O_1027,N_14954,N_14962);
xor UO_1028 (O_1028,N_14902,N_14944);
or UO_1029 (O_1029,N_14875,N_14921);
nor UO_1030 (O_1030,N_14940,N_14923);
or UO_1031 (O_1031,N_14902,N_14975);
nand UO_1032 (O_1032,N_14986,N_14923);
and UO_1033 (O_1033,N_14924,N_14908);
xnor UO_1034 (O_1034,N_14917,N_14962);
nand UO_1035 (O_1035,N_14966,N_14914);
or UO_1036 (O_1036,N_14940,N_14885);
nand UO_1037 (O_1037,N_14944,N_14882);
nor UO_1038 (O_1038,N_14884,N_14927);
nor UO_1039 (O_1039,N_14999,N_14919);
xor UO_1040 (O_1040,N_14893,N_14887);
or UO_1041 (O_1041,N_14984,N_14923);
and UO_1042 (O_1042,N_14929,N_14935);
xnor UO_1043 (O_1043,N_14911,N_14926);
or UO_1044 (O_1044,N_14983,N_14896);
and UO_1045 (O_1045,N_14987,N_14982);
or UO_1046 (O_1046,N_14976,N_14953);
nor UO_1047 (O_1047,N_14974,N_14995);
or UO_1048 (O_1048,N_14886,N_14931);
xor UO_1049 (O_1049,N_14915,N_14920);
xor UO_1050 (O_1050,N_14934,N_14977);
nor UO_1051 (O_1051,N_14927,N_14926);
xnor UO_1052 (O_1052,N_14968,N_14959);
nor UO_1053 (O_1053,N_14994,N_14892);
nand UO_1054 (O_1054,N_14909,N_14990);
nand UO_1055 (O_1055,N_14908,N_14937);
xnor UO_1056 (O_1056,N_14878,N_14995);
and UO_1057 (O_1057,N_14930,N_14897);
or UO_1058 (O_1058,N_14990,N_14922);
nand UO_1059 (O_1059,N_14989,N_14915);
xnor UO_1060 (O_1060,N_14943,N_14999);
nand UO_1061 (O_1061,N_14929,N_14914);
and UO_1062 (O_1062,N_14877,N_14982);
and UO_1063 (O_1063,N_14878,N_14969);
xnor UO_1064 (O_1064,N_14949,N_14888);
xnor UO_1065 (O_1065,N_14889,N_14881);
xnor UO_1066 (O_1066,N_14906,N_14935);
and UO_1067 (O_1067,N_14941,N_14963);
nand UO_1068 (O_1068,N_14937,N_14988);
or UO_1069 (O_1069,N_14977,N_14881);
nor UO_1070 (O_1070,N_14906,N_14955);
and UO_1071 (O_1071,N_14992,N_14960);
xnor UO_1072 (O_1072,N_14890,N_14945);
xnor UO_1073 (O_1073,N_14944,N_14975);
or UO_1074 (O_1074,N_14968,N_14990);
nor UO_1075 (O_1075,N_14888,N_14926);
xor UO_1076 (O_1076,N_14882,N_14909);
and UO_1077 (O_1077,N_14902,N_14912);
xor UO_1078 (O_1078,N_14876,N_14995);
xnor UO_1079 (O_1079,N_14887,N_14932);
nand UO_1080 (O_1080,N_14972,N_14988);
xnor UO_1081 (O_1081,N_14922,N_14887);
xnor UO_1082 (O_1082,N_14985,N_14934);
xor UO_1083 (O_1083,N_14903,N_14922);
nand UO_1084 (O_1084,N_14985,N_14990);
or UO_1085 (O_1085,N_14898,N_14950);
and UO_1086 (O_1086,N_14912,N_14961);
and UO_1087 (O_1087,N_14940,N_14927);
xor UO_1088 (O_1088,N_14955,N_14911);
xor UO_1089 (O_1089,N_14900,N_14917);
or UO_1090 (O_1090,N_14898,N_14953);
or UO_1091 (O_1091,N_14964,N_14880);
or UO_1092 (O_1092,N_14944,N_14875);
or UO_1093 (O_1093,N_14900,N_14961);
nand UO_1094 (O_1094,N_14979,N_14909);
and UO_1095 (O_1095,N_14929,N_14980);
and UO_1096 (O_1096,N_14958,N_14905);
and UO_1097 (O_1097,N_14907,N_14916);
or UO_1098 (O_1098,N_14993,N_14947);
nand UO_1099 (O_1099,N_14917,N_14929);
or UO_1100 (O_1100,N_14920,N_14913);
and UO_1101 (O_1101,N_14907,N_14974);
xnor UO_1102 (O_1102,N_14884,N_14960);
nand UO_1103 (O_1103,N_14904,N_14977);
xnor UO_1104 (O_1104,N_14898,N_14974);
or UO_1105 (O_1105,N_14897,N_14959);
nand UO_1106 (O_1106,N_14947,N_14955);
nand UO_1107 (O_1107,N_14901,N_14904);
or UO_1108 (O_1108,N_14954,N_14894);
nor UO_1109 (O_1109,N_14895,N_14916);
xnor UO_1110 (O_1110,N_14953,N_14912);
nand UO_1111 (O_1111,N_14875,N_14907);
and UO_1112 (O_1112,N_14979,N_14936);
nor UO_1113 (O_1113,N_14982,N_14901);
nor UO_1114 (O_1114,N_14918,N_14888);
or UO_1115 (O_1115,N_14970,N_14894);
or UO_1116 (O_1116,N_14965,N_14991);
or UO_1117 (O_1117,N_14976,N_14882);
nor UO_1118 (O_1118,N_14952,N_14879);
or UO_1119 (O_1119,N_14886,N_14969);
nand UO_1120 (O_1120,N_14973,N_14911);
nor UO_1121 (O_1121,N_14883,N_14895);
xnor UO_1122 (O_1122,N_14908,N_14920);
xnor UO_1123 (O_1123,N_14929,N_14919);
or UO_1124 (O_1124,N_14995,N_14916);
nand UO_1125 (O_1125,N_14923,N_14961);
xnor UO_1126 (O_1126,N_14892,N_14967);
xor UO_1127 (O_1127,N_14876,N_14915);
xor UO_1128 (O_1128,N_14934,N_14931);
or UO_1129 (O_1129,N_14941,N_14998);
and UO_1130 (O_1130,N_14905,N_14889);
or UO_1131 (O_1131,N_14989,N_14945);
nand UO_1132 (O_1132,N_14961,N_14906);
xnor UO_1133 (O_1133,N_14976,N_14948);
and UO_1134 (O_1134,N_14977,N_14924);
nor UO_1135 (O_1135,N_14992,N_14981);
nor UO_1136 (O_1136,N_14892,N_14902);
or UO_1137 (O_1137,N_14955,N_14897);
nor UO_1138 (O_1138,N_14943,N_14885);
nand UO_1139 (O_1139,N_14932,N_14973);
and UO_1140 (O_1140,N_14906,N_14991);
nor UO_1141 (O_1141,N_14978,N_14896);
and UO_1142 (O_1142,N_14878,N_14902);
and UO_1143 (O_1143,N_14958,N_14978);
nand UO_1144 (O_1144,N_14938,N_14918);
and UO_1145 (O_1145,N_14964,N_14928);
xor UO_1146 (O_1146,N_14877,N_14978);
and UO_1147 (O_1147,N_14997,N_14901);
and UO_1148 (O_1148,N_14948,N_14907);
or UO_1149 (O_1149,N_14945,N_14946);
nand UO_1150 (O_1150,N_14978,N_14951);
nor UO_1151 (O_1151,N_14918,N_14953);
nand UO_1152 (O_1152,N_14916,N_14906);
nor UO_1153 (O_1153,N_14945,N_14882);
xnor UO_1154 (O_1154,N_14963,N_14969);
nand UO_1155 (O_1155,N_14877,N_14945);
xnor UO_1156 (O_1156,N_14984,N_14987);
and UO_1157 (O_1157,N_14911,N_14894);
xnor UO_1158 (O_1158,N_14916,N_14919);
or UO_1159 (O_1159,N_14943,N_14925);
nor UO_1160 (O_1160,N_14915,N_14962);
and UO_1161 (O_1161,N_14911,N_14921);
or UO_1162 (O_1162,N_14924,N_14938);
xnor UO_1163 (O_1163,N_14884,N_14977);
or UO_1164 (O_1164,N_14953,N_14928);
nand UO_1165 (O_1165,N_14920,N_14888);
xnor UO_1166 (O_1166,N_14925,N_14891);
or UO_1167 (O_1167,N_14994,N_14982);
xor UO_1168 (O_1168,N_14980,N_14886);
and UO_1169 (O_1169,N_14961,N_14996);
nor UO_1170 (O_1170,N_14916,N_14897);
nor UO_1171 (O_1171,N_14955,N_14935);
or UO_1172 (O_1172,N_14981,N_14940);
nor UO_1173 (O_1173,N_14943,N_14936);
or UO_1174 (O_1174,N_14889,N_14904);
nor UO_1175 (O_1175,N_14889,N_14991);
and UO_1176 (O_1176,N_14958,N_14918);
nand UO_1177 (O_1177,N_14936,N_14942);
or UO_1178 (O_1178,N_14891,N_14902);
xor UO_1179 (O_1179,N_14927,N_14986);
nand UO_1180 (O_1180,N_14982,N_14966);
nand UO_1181 (O_1181,N_14998,N_14883);
or UO_1182 (O_1182,N_14920,N_14959);
or UO_1183 (O_1183,N_14932,N_14979);
nand UO_1184 (O_1184,N_14990,N_14997);
nor UO_1185 (O_1185,N_14971,N_14986);
xnor UO_1186 (O_1186,N_14877,N_14909);
nand UO_1187 (O_1187,N_14995,N_14986);
xnor UO_1188 (O_1188,N_14923,N_14957);
or UO_1189 (O_1189,N_14889,N_14911);
nand UO_1190 (O_1190,N_14970,N_14935);
or UO_1191 (O_1191,N_14944,N_14955);
nand UO_1192 (O_1192,N_14926,N_14979);
xor UO_1193 (O_1193,N_14900,N_14890);
nand UO_1194 (O_1194,N_14901,N_14994);
or UO_1195 (O_1195,N_14889,N_14935);
or UO_1196 (O_1196,N_14918,N_14943);
nor UO_1197 (O_1197,N_14993,N_14979);
nor UO_1198 (O_1198,N_14994,N_14996);
or UO_1199 (O_1199,N_14919,N_14892);
xnor UO_1200 (O_1200,N_14992,N_14883);
or UO_1201 (O_1201,N_14987,N_14941);
or UO_1202 (O_1202,N_14969,N_14875);
and UO_1203 (O_1203,N_14932,N_14908);
nor UO_1204 (O_1204,N_14980,N_14934);
xor UO_1205 (O_1205,N_14938,N_14929);
and UO_1206 (O_1206,N_14920,N_14991);
xor UO_1207 (O_1207,N_14905,N_14938);
xor UO_1208 (O_1208,N_14928,N_14885);
nand UO_1209 (O_1209,N_14948,N_14920);
nand UO_1210 (O_1210,N_14988,N_14996);
or UO_1211 (O_1211,N_14958,N_14990);
nor UO_1212 (O_1212,N_14991,N_14985);
nand UO_1213 (O_1213,N_14922,N_14992);
nand UO_1214 (O_1214,N_14982,N_14917);
nand UO_1215 (O_1215,N_14926,N_14962);
xnor UO_1216 (O_1216,N_14979,N_14885);
and UO_1217 (O_1217,N_14889,N_14949);
nand UO_1218 (O_1218,N_14961,N_14971);
and UO_1219 (O_1219,N_14948,N_14934);
nand UO_1220 (O_1220,N_14905,N_14946);
and UO_1221 (O_1221,N_14943,N_14948);
nor UO_1222 (O_1222,N_14929,N_14995);
or UO_1223 (O_1223,N_14879,N_14995);
nor UO_1224 (O_1224,N_14955,N_14958);
nor UO_1225 (O_1225,N_14933,N_14912);
or UO_1226 (O_1226,N_14956,N_14894);
or UO_1227 (O_1227,N_14963,N_14956);
and UO_1228 (O_1228,N_14952,N_14882);
nor UO_1229 (O_1229,N_14875,N_14995);
and UO_1230 (O_1230,N_14986,N_14981);
nor UO_1231 (O_1231,N_14925,N_14923);
and UO_1232 (O_1232,N_14892,N_14887);
nand UO_1233 (O_1233,N_14917,N_14990);
nand UO_1234 (O_1234,N_14958,N_14895);
xnor UO_1235 (O_1235,N_14875,N_14996);
nor UO_1236 (O_1236,N_14928,N_14993);
or UO_1237 (O_1237,N_14924,N_14961);
xor UO_1238 (O_1238,N_14925,N_14988);
or UO_1239 (O_1239,N_14884,N_14994);
nor UO_1240 (O_1240,N_14914,N_14957);
nand UO_1241 (O_1241,N_14917,N_14890);
nand UO_1242 (O_1242,N_14882,N_14921);
xor UO_1243 (O_1243,N_14996,N_14960);
or UO_1244 (O_1244,N_14908,N_14902);
and UO_1245 (O_1245,N_14890,N_14879);
or UO_1246 (O_1246,N_14881,N_14995);
and UO_1247 (O_1247,N_14914,N_14991);
and UO_1248 (O_1248,N_14963,N_14937);
or UO_1249 (O_1249,N_14983,N_14951);
nor UO_1250 (O_1250,N_14950,N_14876);
nand UO_1251 (O_1251,N_14989,N_14922);
nand UO_1252 (O_1252,N_14878,N_14982);
or UO_1253 (O_1253,N_14888,N_14952);
nand UO_1254 (O_1254,N_14925,N_14915);
or UO_1255 (O_1255,N_14900,N_14994);
or UO_1256 (O_1256,N_14940,N_14944);
nor UO_1257 (O_1257,N_14975,N_14991);
xnor UO_1258 (O_1258,N_14991,N_14979);
nand UO_1259 (O_1259,N_14937,N_14960);
nor UO_1260 (O_1260,N_14987,N_14999);
nand UO_1261 (O_1261,N_14899,N_14962);
xnor UO_1262 (O_1262,N_14929,N_14911);
and UO_1263 (O_1263,N_14888,N_14951);
nor UO_1264 (O_1264,N_14971,N_14892);
xor UO_1265 (O_1265,N_14875,N_14883);
or UO_1266 (O_1266,N_14961,N_14891);
nor UO_1267 (O_1267,N_14989,N_14975);
and UO_1268 (O_1268,N_14925,N_14877);
nor UO_1269 (O_1269,N_14981,N_14907);
xnor UO_1270 (O_1270,N_14954,N_14918);
and UO_1271 (O_1271,N_14919,N_14997);
or UO_1272 (O_1272,N_14942,N_14959);
or UO_1273 (O_1273,N_14954,N_14909);
nor UO_1274 (O_1274,N_14956,N_14897);
and UO_1275 (O_1275,N_14988,N_14900);
nor UO_1276 (O_1276,N_14912,N_14956);
and UO_1277 (O_1277,N_14960,N_14935);
xnor UO_1278 (O_1278,N_14941,N_14886);
or UO_1279 (O_1279,N_14892,N_14891);
or UO_1280 (O_1280,N_14905,N_14979);
or UO_1281 (O_1281,N_14998,N_14912);
xnor UO_1282 (O_1282,N_14998,N_14904);
nor UO_1283 (O_1283,N_14930,N_14880);
nand UO_1284 (O_1284,N_14912,N_14966);
nor UO_1285 (O_1285,N_14974,N_14905);
xnor UO_1286 (O_1286,N_14922,N_14949);
nand UO_1287 (O_1287,N_14945,N_14964);
or UO_1288 (O_1288,N_14989,N_14929);
nand UO_1289 (O_1289,N_14937,N_14903);
or UO_1290 (O_1290,N_14942,N_14997);
nor UO_1291 (O_1291,N_14905,N_14968);
xnor UO_1292 (O_1292,N_14962,N_14996);
xnor UO_1293 (O_1293,N_14886,N_14978);
nor UO_1294 (O_1294,N_14985,N_14897);
nor UO_1295 (O_1295,N_14981,N_14923);
nand UO_1296 (O_1296,N_14909,N_14940);
nor UO_1297 (O_1297,N_14983,N_14964);
and UO_1298 (O_1298,N_14922,N_14899);
xor UO_1299 (O_1299,N_14897,N_14939);
and UO_1300 (O_1300,N_14994,N_14972);
or UO_1301 (O_1301,N_14896,N_14958);
and UO_1302 (O_1302,N_14983,N_14893);
nand UO_1303 (O_1303,N_14967,N_14987);
nor UO_1304 (O_1304,N_14909,N_14986);
xnor UO_1305 (O_1305,N_14980,N_14890);
and UO_1306 (O_1306,N_14933,N_14942);
nand UO_1307 (O_1307,N_14988,N_14909);
nand UO_1308 (O_1308,N_14985,N_14986);
nor UO_1309 (O_1309,N_14936,N_14885);
and UO_1310 (O_1310,N_14881,N_14982);
nor UO_1311 (O_1311,N_14931,N_14909);
nand UO_1312 (O_1312,N_14941,N_14902);
xnor UO_1313 (O_1313,N_14999,N_14990);
or UO_1314 (O_1314,N_14959,N_14979);
nand UO_1315 (O_1315,N_14918,N_14923);
nor UO_1316 (O_1316,N_14945,N_14892);
nor UO_1317 (O_1317,N_14899,N_14999);
nor UO_1318 (O_1318,N_14935,N_14967);
or UO_1319 (O_1319,N_14880,N_14882);
and UO_1320 (O_1320,N_14923,N_14876);
nor UO_1321 (O_1321,N_14988,N_14987);
and UO_1322 (O_1322,N_14958,N_14885);
nor UO_1323 (O_1323,N_14930,N_14967);
nor UO_1324 (O_1324,N_14892,N_14932);
xnor UO_1325 (O_1325,N_14906,N_14926);
or UO_1326 (O_1326,N_14983,N_14977);
xor UO_1327 (O_1327,N_14940,N_14935);
xor UO_1328 (O_1328,N_14972,N_14969);
and UO_1329 (O_1329,N_14900,N_14964);
or UO_1330 (O_1330,N_14950,N_14888);
and UO_1331 (O_1331,N_14886,N_14938);
and UO_1332 (O_1332,N_14905,N_14984);
and UO_1333 (O_1333,N_14892,N_14885);
xor UO_1334 (O_1334,N_14877,N_14935);
or UO_1335 (O_1335,N_14914,N_14950);
or UO_1336 (O_1336,N_14977,N_14975);
nand UO_1337 (O_1337,N_14990,N_14962);
nand UO_1338 (O_1338,N_14987,N_14955);
or UO_1339 (O_1339,N_14950,N_14936);
xor UO_1340 (O_1340,N_14973,N_14922);
or UO_1341 (O_1341,N_14966,N_14975);
or UO_1342 (O_1342,N_14977,N_14899);
nand UO_1343 (O_1343,N_14911,N_14936);
nor UO_1344 (O_1344,N_14949,N_14916);
nand UO_1345 (O_1345,N_14937,N_14979);
and UO_1346 (O_1346,N_14921,N_14937);
xnor UO_1347 (O_1347,N_14925,N_14947);
nor UO_1348 (O_1348,N_14969,N_14971);
and UO_1349 (O_1349,N_14914,N_14892);
and UO_1350 (O_1350,N_14895,N_14936);
nor UO_1351 (O_1351,N_14947,N_14875);
nand UO_1352 (O_1352,N_14983,N_14922);
and UO_1353 (O_1353,N_14998,N_14967);
xor UO_1354 (O_1354,N_14909,N_14980);
or UO_1355 (O_1355,N_14916,N_14965);
nand UO_1356 (O_1356,N_14910,N_14909);
xnor UO_1357 (O_1357,N_14908,N_14982);
xor UO_1358 (O_1358,N_14979,N_14899);
or UO_1359 (O_1359,N_14908,N_14875);
nand UO_1360 (O_1360,N_14902,N_14961);
xnor UO_1361 (O_1361,N_14936,N_14956);
nor UO_1362 (O_1362,N_14894,N_14897);
xor UO_1363 (O_1363,N_14935,N_14875);
xnor UO_1364 (O_1364,N_14995,N_14992);
and UO_1365 (O_1365,N_14933,N_14915);
or UO_1366 (O_1366,N_14923,N_14890);
or UO_1367 (O_1367,N_14992,N_14906);
and UO_1368 (O_1368,N_14999,N_14898);
or UO_1369 (O_1369,N_14999,N_14928);
nand UO_1370 (O_1370,N_14964,N_14912);
or UO_1371 (O_1371,N_14947,N_14890);
and UO_1372 (O_1372,N_14903,N_14884);
and UO_1373 (O_1373,N_14964,N_14962);
and UO_1374 (O_1374,N_14933,N_14950);
and UO_1375 (O_1375,N_14994,N_14925);
xnor UO_1376 (O_1376,N_14936,N_14976);
and UO_1377 (O_1377,N_14876,N_14920);
and UO_1378 (O_1378,N_14934,N_14938);
and UO_1379 (O_1379,N_14903,N_14991);
or UO_1380 (O_1380,N_14901,N_14926);
nand UO_1381 (O_1381,N_14897,N_14943);
or UO_1382 (O_1382,N_14938,N_14879);
and UO_1383 (O_1383,N_14895,N_14880);
nand UO_1384 (O_1384,N_14995,N_14880);
or UO_1385 (O_1385,N_14880,N_14931);
nand UO_1386 (O_1386,N_14970,N_14922);
or UO_1387 (O_1387,N_14914,N_14883);
nor UO_1388 (O_1388,N_14965,N_14900);
xnor UO_1389 (O_1389,N_14946,N_14882);
xnor UO_1390 (O_1390,N_14879,N_14908);
nor UO_1391 (O_1391,N_14972,N_14877);
or UO_1392 (O_1392,N_14998,N_14986);
and UO_1393 (O_1393,N_14981,N_14963);
nand UO_1394 (O_1394,N_14931,N_14887);
and UO_1395 (O_1395,N_14882,N_14988);
nor UO_1396 (O_1396,N_14882,N_14974);
nand UO_1397 (O_1397,N_14915,N_14998);
nor UO_1398 (O_1398,N_14888,N_14885);
nand UO_1399 (O_1399,N_14979,N_14914);
nor UO_1400 (O_1400,N_14880,N_14906);
xnor UO_1401 (O_1401,N_14983,N_14909);
or UO_1402 (O_1402,N_14917,N_14997);
nand UO_1403 (O_1403,N_14906,N_14973);
and UO_1404 (O_1404,N_14921,N_14881);
nor UO_1405 (O_1405,N_14917,N_14984);
or UO_1406 (O_1406,N_14878,N_14882);
nor UO_1407 (O_1407,N_14984,N_14889);
nand UO_1408 (O_1408,N_14894,N_14988);
nor UO_1409 (O_1409,N_14999,N_14926);
and UO_1410 (O_1410,N_14930,N_14995);
and UO_1411 (O_1411,N_14912,N_14940);
xor UO_1412 (O_1412,N_14891,N_14905);
or UO_1413 (O_1413,N_14913,N_14893);
nand UO_1414 (O_1414,N_14927,N_14965);
nor UO_1415 (O_1415,N_14979,N_14978);
nor UO_1416 (O_1416,N_14973,N_14902);
nand UO_1417 (O_1417,N_14946,N_14894);
and UO_1418 (O_1418,N_14935,N_14931);
or UO_1419 (O_1419,N_14948,N_14879);
and UO_1420 (O_1420,N_14896,N_14891);
xor UO_1421 (O_1421,N_14875,N_14977);
nor UO_1422 (O_1422,N_14879,N_14997);
and UO_1423 (O_1423,N_14979,N_14967);
nand UO_1424 (O_1424,N_14905,N_14972);
nor UO_1425 (O_1425,N_14878,N_14999);
and UO_1426 (O_1426,N_14952,N_14895);
nor UO_1427 (O_1427,N_14934,N_14908);
and UO_1428 (O_1428,N_14905,N_14897);
nor UO_1429 (O_1429,N_14995,N_14991);
nand UO_1430 (O_1430,N_14949,N_14875);
xnor UO_1431 (O_1431,N_14905,N_14892);
nor UO_1432 (O_1432,N_14879,N_14929);
nand UO_1433 (O_1433,N_14952,N_14877);
and UO_1434 (O_1434,N_14991,N_14938);
nand UO_1435 (O_1435,N_14984,N_14894);
xnor UO_1436 (O_1436,N_14933,N_14955);
nor UO_1437 (O_1437,N_14905,N_14973);
or UO_1438 (O_1438,N_14994,N_14890);
xnor UO_1439 (O_1439,N_14928,N_14966);
and UO_1440 (O_1440,N_14892,N_14980);
and UO_1441 (O_1441,N_14971,N_14890);
and UO_1442 (O_1442,N_14987,N_14962);
and UO_1443 (O_1443,N_14993,N_14907);
xnor UO_1444 (O_1444,N_14952,N_14998);
nor UO_1445 (O_1445,N_14900,N_14921);
xnor UO_1446 (O_1446,N_14876,N_14882);
or UO_1447 (O_1447,N_14988,N_14981);
xnor UO_1448 (O_1448,N_14988,N_14929);
or UO_1449 (O_1449,N_14946,N_14927);
xnor UO_1450 (O_1450,N_14899,N_14928);
and UO_1451 (O_1451,N_14916,N_14968);
nand UO_1452 (O_1452,N_14890,N_14960);
nor UO_1453 (O_1453,N_14917,N_14934);
xor UO_1454 (O_1454,N_14966,N_14882);
nor UO_1455 (O_1455,N_14942,N_14909);
or UO_1456 (O_1456,N_14995,N_14926);
and UO_1457 (O_1457,N_14898,N_14991);
or UO_1458 (O_1458,N_14985,N_14917);
or UO_1459 (O_1459,N_14922,N_14876);
xor UO_1460 (O_1460,N_14958,N_14949);
xor UO_1461 (O_1461,N_14877,N_14985);
and UO_1462 (O_1462,N_14906,N_14981);
xnor UO_1463 (O_1463,N_14939,N_14904);
or UO_1464 (O_1464,N_14885,N_14951);
or UO_1465 (O_1465,N_14971,N_14960);
or UO_1466 (O_1466,N_14900,N_14959);
nand UO_1467 (O_1467,N_14892,N_14941);
or UO_1468 (O_1468,N_14977,N_14949);
or UO_1469 (O_1469,N_14921,N_14909);
xnor UO_1470 (O_1470,N_14938,N_14955);
nand UO_1471 (O_1471,N_14877,N_14961);
nor UO_1472 (O_1472,N_14953,N_14954);
or UO_1473 (O_1473,N_14913,N_14902);
or UO_1474 (O_1474,N_14911,N_14931);
or UO_1475 (O_1475,N_14988,N_14969);
or UO_1476 (O_1476,N_14905,N_14900);
xor UO_1477 (O_1477,N_14947,N_14914);
xor UO_1478 (O_1478,N_14970,N_14993);
and UO_1479 (O_1479,N_14968,N_14996);
nor UO_1480 (O_1480,N_14924,N_14900);
xor UO_1481 (O_1481,N_14877,N_14887);
xnor UO_1482 (O_1482,N_14928,N_14883);
nand UO_1483 (O_1483,N_14882,N_14956);
xnor UO_1484 (O_1484,N_14949,N_14910);
nand UO_1485 (O_1485,N_14959,N_14944);
or UO_1486 (O_1486,N_14935,N_14969);
nor UO_1487 (O_1487,N_14921,N_14954);
or UO_1488 (O_1488,N_14904,N_14913);
xnor UO_1489 (O_1489,N_14897,N_14997);
xnor UO_1490 (O_1490,N_14981,N_14961);
or UO_1491 (O_1491,N_14901,N_14999);
nor UO_1492 (O_1492,N_14952,N_14885);
nand UO_1493 (O_1493,N_14896,N_14997);
and UO_1494 (O_1494,N_14951,N_14993);
nand UO_1495 (O_1495,N_14925,N_14905);
or UO_1496 (O_1496,N_14902,N_14938);
nor UO_1497 (O_1497,N_14910,N_14902);
nand UO_1498 (O_1498,N_14897,N_14891);
nand UO_1499 (O_1499,N_14932,N_14941);
and UO_1500 (O_1500,N_14891,N_14986);
xor UO_1501 (O_1501,N_14960,N_14875);
xnor UO_1502 (O_1502,N_14913,N_14955);
xor UO_1503 (O_1503,N_14895,N_14989);
or UO_1504 (O_1504,N_14981,N_14965);
and UO_1505 (O_1505,N_14959,N_14909);
or UO_1506 (O_1506,N_14943,N_14950);
and UO_1507 (O_1507,N_14973,N_14916);
or UO_1508 (O_1508,N_14978,N_14965);
or UO_1509 (O_1509,N_14891,N_14944);
or UO_1510 (O_1510,N_14973,N_14965);
and UO_1511 (O_1511,N_14980,N_14953);
xor UO_1512 (O_1512,N_14974,N_14969);
or UO_1513 (O_1513,N_14884,N_14912);
and UO_1514 (O_1514,N_14929,N_14886);
nor UO_1515 (O_1515,N_14901,N_14967);
or UO_1516 (O_1516,N_14973,N_14899);
or UO_1517 (O_1517,N_14973,N_14913);
nand UO_1518 (O_1518,N_14961,N_14897);
and UO_1519 (O_1519,N_14947,N_14893);
or UO_1520 (O_1520,N_14963,N_14973);
nand UO_1521 (O_1521,N_14989,N_14956);
and UO_1522 (O_1522,N_14929,N_14983);
or UO_1523 (O_1523,N_14996,N_14995);
nand UO_1524 (O_1524,N_14981,N_14931);
nor UO_1525 (O_1525,N_14889,N_14939);
xor UO_1526 (O_1526,N_14977,N_14914);
and UO_1527 (O_1527,N_14928,N_14929);
or UO_1528 (O_1528,N_14943,N_14896);
and UO_1529 (O_1529,N_14912,N_14969);
or UO_1530 (O_1530,N_14879,N_14935);
xor UO_1531 (O_1531,N_14946,N_14902);
nand UO_1532 (O_1532,N_14888,N_14924);
or UO_1533 (O_1533,N_14913,N_14961);
and UO_1534 (O_1534,N_14985,N_14918);
nor UO_1535 (O_1535,N_14878,N_14910);
xnor UO_1536 (O_1536,N_14938,N_14994);
or UO_1537 (O_1537,N_14994,N_14910);
nand UO_1538 (O_1538,N_14995,N_14886);
nor UO_1539 (O_1539,N_14946,N_14890);
nor UO_1540 (O_1540,N_14961,N_14901);
or UO_1541 (O_1541,N_14931,N_14976);
nor UO_1542 (O_1542,N_14881,N_14904);
and UO_1543 (O_1543,N_14976,N_14920);
nor UO_1544 (O_1544,N_14981,N_14948);
xnor UO_1545 (O_1545,N_14958,N_14959);
nand UO_1546 (O_1546,N_14938,N_14999);
nor UO_1547 (O_1547,N_14942,N_14907);
xor UO_1548 (O_1548,N_14941,N_14945);
or UO_1549 (O_1549,N_14944,N_14934);
or UO_1550 (O_1550,N_14919,N_14879);
nand UO_1551 (O_1551,N_14956,N_14990);
nor UO_1552 (O_1552,N_14985,N_14941);
nor UO_1553 (O_1553,N_14991,N_14894);
nand UO_1554 (O_1554,N_14985,N_14921);
or UO_1555 (O_1555,N_14996,N_14915);
and UO_1556 (O_1556,N_14948,N_14965);
or UO_1557 (O_1557,N_14965,N_14894);
nor UO_1558 (O_1558,N_14910,N_14978);
nor UO_1559 (O_1559,N_14881,N_14957);
and UO_1560 (O_1560,N_14955,N_14996);
nand UO_1561 (O_1561,N_14991,N_14963);
xnor UO_1562 (O_1562,N_14883,N_14879);
and UO_1563 (O_1563,N_14918,N_14917);
nor UO_1564 (O_1564,N_14952,N_14907);
nand UO_1565 (O_1565,N_14900,N_14984);
xnor UO_1566 (O_1566,N_14944,N_14877);
nand UO_1567 (O_1567,N_14948,N_14978);
nor UO_1568 (O_1568,N_14928,N_14915);
or UO_1569 (O_1569,N_14886,N_14915);
or UO_1570 (O_1570,N_14894,N_14887);
and UO_1571 (O_1571,N_14924,N_14991);
or UO_1572 (O_1572,N_14926,N_14895);
xnor UO_1573 (O_1573,N_14912,N_14897);
or UO_1574 (O_1574,N_14945,N_14969);
nand UO_1575 (O_1575,N_14985,N_14959);
or UO_1576 (O_1576,N_14954,N_14936);
or UO_1577 (O_1577,N_14912,N_14905);
nor UO_1578 (O_1578,N_14960,N_14930);
or UO_1579 (O_1579,N_14995,N_14950);
or UO_1580 (O_1580,N_14930,N_14921);
xor UO_1581 (O_1581,N_14983,N_14880);
and UO_1582 (O_1582,N_14938,N_14945);
or UO_1583 (O_1583,N_14973,N_14944);
or UO_1584 (O_1584,N_14953,N_14922);
and UO_1585 (O_1585,N_14921,N_14946);
nor UO_1586 (O_1586,N_14898,N_14979);
xor UO_1587 (O_1587,N_14935,N_14985);
and UO_1588 (O_1588,N_14953,N_14958);
nand UO_1589 (O_1589,N_14948,N_14969);
nor UO_1590 (O_1590,N_14902,N_14989);
and UO_1591 (O_1591,N_14895,N_14988);
nor UO_1592 (O_1592,N_14993,N_14878);
nand UO_1593 (O_1593,N_14979,N_14964);
or UO_1594 (O_1594,N_14957,N_14928);
nand UO_1595 (O_1595,N_14884,N_14946);
xor UO_1596 (O_1596,N_14881,N_14997);
or UO_1597 (O_1597,N_14929,N_14884);
nor UO_1598 (O_1598,N_14931,N_14978);
and UO_1599 (O_1599,N_14904,N_14876);
or UO_1600 (O_1600,N_14974,N_14960);
nor UO_1601 (O_1601,N_14911,N_14879);
xor UO_1602 (O_1602,N_14899,N_14982);
nand UO_1603 (O_1603,N_14966,N_14995);
xor UO_1604 (O_1604,N_14996,N_14964);
nor UO_1605 (O_1605,N_14888,N_14921);
nor UO_1606 (O_1606,N_14913,N_14980);
nor UO_1607 (O_1607,N_14880,N_14980);
xnor UO_1608 (O_1608,N_14908,N_14913);
or UO_1609 (O_1609,N_14930,N_14961);
xor UO_1610 (O_1610,N_14953,N_14988);
or UO_1611 (O_1611,N_14966,N_14913);
or UO_1612 (O_1612,N_14957,N_14917);
nand UO_1613 (O_1613,N_14977,N_14890);
nor UO_1614 (O_1614,N_14982,N_14924);
nor UO_1615 (O_1615,N_14980,N_14947);
and UO_1616 (O_1616,N_14942,N_14941);
nand UO_1617 (O_1617,N_14992,N_14903);
and UO_1618 (O_1618,N_14905,N_14977);
nor UO_1619 (O_1619,N_14945,N_14918);
and UO_1620 (O_1620,N_14974,N_14987);
and UO_1621 (O_1621,N_14966,N_14942);
or UO_1622 (O_1622,N_14994,N_14927);
or UO_1623 (O_1623,N_14892,N_14986);
or UO_1624 (O_1624,N_14885,N_14910);
nand UO_1625 (O_1625,N_14954,N_14888);
or UO_1626 (O_1626,N_14890,N_14898);
nand UO_1627 (O_1627,N_14987,N_14922);
nor UO_1628 (O_1628,N_14886,N_14943);
nor UO_1629 (O_1629,N_14976,N_14919);
or UO_1630 (O_1630,N_14926,N_14976);
nand UO_1631 (O_1631,N_14979,N_14958);
and UO_1632 (O_1632,N_14875,N_14957);
and UO_1633 (O_1633,N_14999,N_14981);
xor UO_1634 (O_1634,N_14972,N_14896);
xnor UO_1635 (O_1635,N_14881,N_14992);
xnor UO_1636 (O_1636,N_14888,N_14955);
or UO_1637 (O_1637,N_14885,N_14984);
nor UO_1638 (O_1638,N_14876,N_14966);
nand UO_1639 (O_1639,N_14945,N_14880);
nand UO_1640 (O_1640,N_14967,N_14958);
nand UO_1641 (O_1641,N_14937,N_14909);
and UO_1642 (O_1642,N_14962,N_14935);
nand UO_1643 (O_1643,N_14939,N_14977);
or UO_1644 (O_1644,N_14898,N_14993);
nor UO_1645 (O_1645,N_14943,N_14981);
or UO_1646 (O_1646,N_14878,N_14979);
or UO_1647 (O_1647,N_14965,N_14902);
xnor UO_1648 (O_1648,N_14972,N_14958);
or UO_1649 (O_1649,N_14942,N_14903);
nor UO_1650 (O_1650,N_14879,N_14902);
or UO_1651 (O_1651,N_14944,N_14954);
nand UO_1652 (O_1652,N_14889,N_14978);
nand UO_1653 (O_1653,N_14904,N_14906);
nor UO_1654 (O_1654,N_14991,N_14972);
xor UO_1655 (O_1655,N_14941,N_14929);
nand UO_1656 (O_1656,N_14998,N_14985);
nand UO_1657 (O_1657,N_14931,N_14926);
nor UO_1658 (O_1658,N_14931,N_14983);
nor UO_1659 (O_1659,N_14882,N_14993);
and UO_1660 (O_1660,N_14962,N_14904);
and UO_1661 (O_1661,N_14884,N_14993);
xnor UO_1662 (O_1662,N_14888,N_14925);
nor UO_1663 (O_1663,N_14980,N_14875);
nand UO_1664 (O_1664,N_14973,N_14985);
nand UO_1665 (O_1665,N_14989,N_14912);
nor UO_1666 (O_1666,N_14891,N_14934);
or UO_1667 (O_1667,N_14911,N_14919);
and UO_1668 (O_1668,N_14991,N_14978);
xor UO_1669 (O_1669,N_14998,N_14921);
or UO_1670 (O_1670,N_14932,N_14962);
nor UO_1671 (O_1671,N_14948,N_14962);
xor UO_1672 (O_1672,N_14954,N_14925);
and UO_1673 (O_1673,N_14976,N_14930);
nand UO_1674 (O_1674,N_14896,N_14877);
xor UO_1675 (O_1675,N_14933,N_14902);
and UO_1676 (O_1676,N_14937,N_14977);
and UO_1677 (O_1677,N_14977,N_14888);
and UO_1678 (O_1678,N_14933,N_14888);
and UO_1679 (O_1679,N_14996,N_14958);
xor UO_1680 (O_1680,N_14985,N_14994);
and UO_1681 (O_1681,N_14927,N_14993);
nand UO_1682 (O_1682,N_14938,N_14983);
nand UO_1683 (O_1683,N_14961,N_14931);
nand UO_1684 (O_1684,N_14950,N_14989);
xor UO_1685 (O_1685,N_14997,N_14935);
or UO_1686 (O_1686,N_14980,N_14887);
xor UO_1687 (O_1687,N_14888,N_14983);
or UO_1688 (O_1688,N_14931,N_14906);
or UO_1689 (O_1689,N_14999,N_14923);
xnor UO_1690 (O_1690,N_14950,N_14899);
nand UO_1691 (O_1691,N_14913,N_14998);
and UO_1692 (O_1692,N_14923,N_14915);
or UO_1693 (O_1693,N_14888,N_14957);
nand UO_1694 (O_1694,N_14991,N_14895);
xnor UO_1695 (O_1695,N_14877,N_14959);
xor UO_1696 (O_1696,N_14931,N_14884);
nor UO_1697 (O_1697,N_14955,N_14950);
xor UO_1698 (O_1698,N_14893,N_14989);
xnor UO_1699 (O_1699,N_14921,N_14997);
nand UO_1700 (O_1700,N_14974,N_14935);
nand UO_1701 (O_1701,N_14891,N_14973);
nor UO_1702 (O_1702,N_14875,N_14910);
nand UO_1703 (O_1703,N_14909,N_14876);
nand UO_1704 (O_1704,N_14966,N_14963);
nand UO_1705 (O_1705,N_14903,N_14902);
and UO_1706 (O_1706,N_14924,N_14986);
nand UO_1707 (O_1707,N_14970,N_14981);
xnor UO_1708 (O_1708,N_14964,N_14991);
and UO_1709 (O_1709,N_14960,N_14899);
or UO_1710 (O_1710,N_14979,N_14888);
or UO_1711 (O_1711,N_14891,N_14987);
nand UO_1712 (O_1712,N_14972,N_14929);
and UO_1713 (O_1713,N_14978,N_14936);
nand UO_1714 (O_1714,N_14968,N_14938);
and UO_1715 (O_1715,N_14947,N_14888);
nand UO_1716 (O_1716,N_14941,N_14953);
nand UO_1717 (O_1717,N_14973,N_14907);
nor UO_1718 (O_1718,N_14993,N_14911);
and UO_1719 (O_1719,N_14923,N_14924);
nand UO_1720 (O_1720,N_14897,N_14957);
xor UO_1721 (O_1721,N_14989,N_14921);
and UO_1722 (O_1722,N_14914,N_14993);
or UO_1723 (O_1723,N_14967,N_14961);
xnor UO_1724 (O_1724,N_14904,N_14938);
or UO_1725 (O_1725,N_14973,N_14900);
nand UO_1726 (O_1726,N_14981,N_14897);
and UO_1727 (O_1727,N_14963,N_14922);
xor UO_1728 (O_1728,N_14895,N_14887);
xnor UO_1729 (O_1729,N_14982,N_14974);
and UO_1730 (O_1730,N_14997,N_14972);
nor UO_1731 (O_1731,N_14929,N_14976);
nand UO_1732 (O_1732,N_14920,N_14895);
xnor UO_1733 (O_1733,N_14914,N_14896);
nor UO_1734 (O_1734,N_14924,N_14922);
nand UO_1735 (O_1735,N_14902,N_14914);
nand UO_1736 (O_1736,N_14920,N_14892);
and UO_1737 (O_1737,N_14881,N_14964);
nand UO_1738 (O_1738,N_14881,N_14922);
xnor UO_1739 (O_1739,N_14999,N_14929);
nor UO_1740 (O_1740,N_14992,N_14913);
nor UO_1741 (O_1741,N_14892,N_14884);
xor UO_1742 (O_1742,N_14983,N_14930);
or UO_1743 (O_1743,N_14898,N_14881);
xnor UO_1744 (O_1744,N_14966,N_14934);
or UO_1745 (O_1745,N_14914,N_14916);
nor UO_1746 (O_1746,N_14951,N_14890);
nand UO_1747 (O_1747,N_14879,N_14878);
and UO_1748 (O_1748,N_14926,N_14956);
nor UO_1749 (O_1749,N_14995,N_14994);
nor UO_1750 (O_1750,N_14967,N_14925);
or UO_1751 (O_1751,N_14948,N_14971);
nand UO_1752 (O_1752,N_14987,N_14990);
or UO_1753 (O_1753,N_14909,N_14908);
nand UO_1754 (O_1754,N_14999,N_14949);
or UO_1755 (O_1755,N_14969,N_14910);
and UO_1756 (O_1756,N_14968,N_14912);
nand UO_1757 (O_1757,N_14949,N_14880);
nor UO_1758 (O_1758,N_14976,N_14962);
and UO_1759 (O_1759,N_14946,N_14928);
nor UO_1760 (O_1760,N_14972,N_14981);
nand UO_1761 (O_1761,N_14946,N_14932);
nor UO_1762 (O_1762,N_14931,N_14936);
xnor UO_1763 (O_1763,N_14992,N_14978);
or UO_1764 (O_1764,N_14887,N_14883);
and UO_1765 (O_1765,N_14881,N_14989);
and UO_1766 (O_1766,N_14898,N_14878);
nand UO_1767 (O_1767,N_14965,N_14938);
nor UO_1768 (O_1768,N_14998,N_14878);
or UO_1769 (O_1769,N_14959,N_14905);
nor UO_1770 (O_1770,N_14963,N_14995);
and UO_1771 (O_1771,N_14970,N_14920);
and UO_1772 (O_1772,N_14892,N_14961);
and UO_1773 (O_1773,N_14959,N_14982);
and UO_1774 (O_1774,N_14941,N_14903);
xor UO_1775 (O_1775,N_14990,N_14920);
and UO_1776 (O_1776,N_14907,N_14928);
xor UO_1777 (O_1777,N_14985,N_14982);
or UO_1778 (O_1778,N_14906,N_14893);
nor UO_1779 (O_1779,N_14878,N_14889);
xor UO_1780 (O_1780,N_14929,N_14908);
and UO_1781 (O_1781,N_14970,N_14924);
nor UO_1782 (O_1782,N_14944,N_14984);
or UO_1783 (O_1783,N_14879,N_14885);
xnor UO_1784 (O_1784,N_14971,N_14975);
nor UO_1785 (O_1785,N_14991,N_14936);
nand UO_1786 (O_1786,N_14993,N_14996);
nand UO_1787 (O_1787,N_14883,N_14900);
nor UO_1788 (O_1788,N_14958,N_14946);
xor UO_1789 (O_1789,N_14919,N_14963);
nand UO_1790 (O_1790,N_14885,N_14883);
xor UO_1791 (O_1791,N_14891,N_14880);
nand UO_1792 (O_1792,N_14939,N_14931);
and UO_1793 (O_1793,N_14936,N_14977);
nand UO_1794 (O_1794,N_14913,N_14936);
nand UO_1795 (O_1795,N_14970,N_14910);
or UO_1796 (O_1796,N_14916,N_14970);
nor UO_1797 (O_1797,N_14971,N_14945);
or UO_1798 (O_1798,N_14907,N_14895);
and UO_1799 (O_1799,N_14976,N_14955);
nand UO_1800 (O_1800,N_14893,N_14897);
xor UO_1801 (O_1801,N_14945,N_14925);
nor UO_1802 (O_1802,N_14917,N_14931);
xor UO_1803 (O_1803,N_14931,N_14877);
or UO_1804 (O_1804,N_14940,N_14918);
nand UO_1805 (O_1805,N_14948,N_14919);
xnor UO_1806 (O_1806,N_14909,N_14987);
or UO_1807 (O_1807,N_14895,N_14975);
or UO_1808 (O_1808,N_14933,N_14989);
nor UO_1809 (O_1809,N_14927,N_14939);
and UO_1810 (O_1810,N_14994,N_14903);
xnor UO_1811 (O_1811,N_14979,N_14903);
xnor UO_1812 (O_1812,N_14890,N_14895);
nor UO_1813 (O_1813,N_14963,N_14917);
and UO_1814 (O_1814,N_14927,N_14997);
nor UO_1815 (O_1815,N_14931,N_14937);
nor UO_1816 (O_1816,N_14978,N_14875);
xnor UO_1817 (O_1817,N_14995,N_14969);
and UO_1818 (O_1818,N_14961,N_14995);
xnor UO_1819 (O_1819,N_14902,N_14960);
or UO_1820 (O_1820,N_14878,N_14966);
and UO_1821 (O_1821,N_14885,N_14896);
nand UO_1822 (O_1822,N_14986,N_14875);
and UO_1823 (O_1823,N_14889,N_14907);
or UO_1824 (O_1824,N_14897,N_14986);
xnor UO_1825 (O_1825,N_14926,N_14941);
or UO_1826 (O_1826,N_14923,N_14941);
nor UO_1827 (O_1827,N_14995,N_14883);
and UO_1828 (O_1828,N_14969,N_14954);
or UO_1829 (O_1829,N_14881,N_14962);
xor UO_1830 (O_1830,N_14879,N_14980);
or UO_1831 (O_1831,N_14985,N_14967);
and UO_1832 (O_1832,N_14994,N_14983);
nand UO_1833 (O_1833,N_14924,N_14910);
and UO_1834 (O_1834,N_14963,N_14955);
nor UO_1835 (O_1835,N_14930,N_14950);
and UO_1836 (O_1836,N_14918,N_14979);
nor UO_1837 (O_1837,N_14923,N_14896);
nand UO_1838 (O_1838,N_14995,N_14887);
xor UO_1839 (O_1839,N_14892,N_14982);
and UO_1840 (O_1840,N_14883,N_14977);
xor UO_1841 (O_1841,N_14935,N_14897);
nand UO_1842 (O_1842,N_14895,N_14901);
nor UO_1843 (O_1843,N_14998,N_14948);
or UO_1844 (O_1844,N_14913,N_14883);
and UO_1845 (O_1845,N_14961,N_14941);
nand UO_1846 (O_1846,N_14884,N_14945);
and UO_1847 (O_1847,N_14878,N_14892);
or UO_1848 (O_1848,N_14982,N_14904);
nor UO_1849 (O_1849,N_14954,N_14999);
nor UO_1850 (O_1850,N_14960,N_14962);
or UO_1851 (O_1851,N_14981,N_14901);
xnor UO_1852 (O_1852,N_14967,N_14896);
and UO_1853 (O_1853,N_14993,N_14962);
nor UO_1854 (O_1854,N_14976,N_14991);
xnor UO_1855 (O_1855,N_14914,N_14998);
nand UO_1856 (O_1856,N_14875,N_14911);
nand UO_1857 (O_1857,N_14922,N_14904);
and UO_1858 (O_1858,N_14904,N_14900);
xnor UO_1859 (O_1859,N_14988,N_14986);
nor UO_1860 (O_1860,N_14886,N_14922);
xor UO_1861 (O_1861,N_14884,N_14924);
nand UO_1862 (O_1862,N_14948,N_14992);
xor UO_1863 (O_1863,N_14938,N_14885);
or UO_1864 (O_1864,N_14883,N_14904);
nor UO_1865 (O_1865,N_14893,N_14892);
nor UO_1866 (O_1866,N_14910,N_14926);
xor UO_1867 (O_1867,N_14935,N_14911);
nand UO_1868 (O_1868,N_14994,N_14882);
nand UO_1869 (O_1869,N_14919,N_14993);
nand UO_1870 (O_1870,N_14946,N_14935);
or UO_1871 (O_1871,N_14890,N_14882);
and UO_1872 (O_1872,N_14875,N_14945);
nand UO_1873 (O_1873,N_14887,N_14965);
or UO_1874 (O_1874,N_14902,N_14880);
nor UO_1875 (O_1875,N_14884,N_14956);
nor UO_1876 (O_1876,N_14902,N_14896);
xnor UO_1877 (O_1877,N_14943,N_14912);
xnor UO_1878 (O_1878,N_14900,N_14978);
xnor UO_1879 (O_1879,N_14958,N_14921);
nand UO_1880 (O_1880,N_14934,N_14893);
nand UO_1881 (O_1881,N_14917,N_14907);
xor UO_1882 (O_1882,N_14965,N_14882);
and UO_1883 (O_1883,N_14877,N_14900);
nand UO_1884 (O_1884,N_14937,N_14911);
and UO_1885 (O_1885,N_14904,N_14931);
or UO_1886 (O_1886,N_14975,N_14917);
and UO_1887 (O_1887,N_14939,N_14958);
or UO_1888 (O_1888,N_14938,N_14915);
and UO_1889 (O_1889,N_14993,N_14905);
nand UO_1890 (O_1890,N_14936,N_14996);
xnor UO_1891 (O_1891,N_14974,N_14981);
or UO_1892 (O_1892,N_14937,N_14898);
nand UO_1893 (O_1893,N_14988,N_14877);
or UO_1894 (O_1894,N_14910,N_14899);
nand UO_1895 (O_1895,N_14875,N_14975);
nand UO_1896 (O_1896,N_14962,N_14969);
and UO_1897 (O_1897,N_14966,N_14916);
nand UO_1898 (O_1898,N_14903,N_14885);
xor UO_1899 (O_1899,N_14905,N_14885);
nand UO_1900 (O_1900,N_14930,N_14974);
or UO_1901 (O_1901,N_14979,N_14997);
nand UO_1902 (O_1902,N_14908,N_14975);
nor UO_1903 (O_1903,N_14985,N_14987);
or UO_1904 (O_1904,N_14986,N_14885);
nand UO_1905 (O_1905,N_14947,N_14957);
or UO_1906 (O_1906,N_14921,N_14940);
nand UO_1907 (O_1907,N_14936,N_14927);
and UO_1908 (O_1908,N_14951,N_14925);
or UO_1909 (O_1909,N_14978,N_14989);
nor UO_1910 (O_1910,N_14883,N_14931);
nand UO_1911 (O_1911,N_14928,N_14954);
nor UO_1912 (O_1912,N_14905,N_14924);
and UO_1913 (O_1913,N_14978,N_14913);
xor UO_1914 (O_1914,N_14914,N_14932);
xnor UO_1915 (O_1915,N_14925,N_14978);
xor UO_1916 (O_1916,N_14895,N_14892);
xor UO_1917 (O_1917,N_14941,N_14989);
or UO_1918 (O_1918,N_14910,N_14894);
xnor UO_1919 (O_1919,N_14943,N_14994);
or UO_1920 (O_1920,N_14912,N_14903);
nor UO_1921 (O_1921,N_14906,N_14959);
nand UO_1922 (O_1922,N_14885,N_14932);
nor UO_1923 (O_1923,N_14932,N_14915);
xor UO_1924 (O_1924,N_14900,N_14970);
xnor UO_1925 (O_1925,N_14933,N_14987);
or UO_1926 (O_1926,N_14990,N_14964);
or UO_1927 (O_1927,N_14939,N_14976);
and UO_1928 (O_1928,N_14912,N_14963);
or UO_1929 (O_1929,N_14897,N_14974);
or UO_1930 (O_1930,N_14915,N_14968);
nand UO_1931 (O_1931,N_14935,N_14990);
nor UO_1932 (O_1932,N_14992,N_14917);
nor UO_1933 (O_1933,N_14971,N_14933);
and UO_1934 (O_1934,N_14991,N_14960);
and UO_1935 (O_1935,N_14998,N_14889);
nand UO_1936 (O_1936,N_14921,N_14943);
xor UO_1937 (O_1937,N_14884,N_14875);
or UO_1938 (O_1938,N_14954,N_14996);
or UO_1939 (O_1939,N_14906,N_14982);
and UO_1940 (O_1940,N_14910,N_14961);
nor UO_1941 (O_1941,N_14963,N_14900);
nor UO_1942 (O_1942,N_14941,N_14920);
or UO_1943 (O_1943,N_14971,N_14998);
nor UO_1944 (O_1944,N_14905,N_14875);
and UO_1945 (O_1945,N_14986,N_14968);
nand UO_1946 (O_1946,N_14936,N_14990);
xnor UO_1947 (O_1947,N_14876,N_14893);
or UO_1948 (O_1948,N_14897,N_14967);
xor UO_1949 (O_1949,N_14952,N_14875);
and UO_1950 (O_1950,N_14894,N_14967);
xor UO_1951 (O_1951,N_14939,N_14994);
or UO_1952 (O_1952,N_14908,N_14974);
and UO_1953 (O_1953,N_14962,N_14889);
nand UO_1954 (O_1954,N_14898,N_14934);
or UO_1955 (O_1955,N_14942,N_14975);
xnor UO_1956 (O_1956,N_14926,N_14886);
xnor UO_1957 (O_1957,N_14989,N_14891);
nor UO_1958 (O_1958,N_14908,N_14954);
xnor UO_1959 (O_1959,N_14880,N_14890);
and UO_1960 (O_1960,N_14961,N_14947);
xor UO_1961 (O_1961,N_14958,N_14947);
or UO_1962 (O_1962,N_14904,N_14985);
and UO_1963 (O_1963,N_14896,N_14929);
or UO_1964 (O_1964,N_14884,N_14937);
or UO_1965 (O_1965,N_14880,N_14985);
nand UO_1966 (O_1966,N_14964,N_14984);
and UO_1967 (O_1967,N_14958,N_14980);
xnor UO_1968 (O_1968,N_14932,N_14994);
or UO_1969 (O_1969,N_14918,N_14941);
and UO_1970 (O_1970,N_14929,N_14955);
xnor UO_1971 (O_1971,N_14920,N_14935);
and UO_1972 (O_1972,N_14919,N_14947);
nand UO_1973 (O_1973,N_14883,N_14936);
and UO_1974 (O_1974,N_14891,N_14962);
and UO_1975 (O_1975,N_14908,N_14914);
nand UO_1976 (O_1976,N_14900,N_14945);
nor UO_1977 (O_1977,N_14916,N_14955);
xnor UO_1978 (O_1978,N_14991,N_14937);
xor UO_1979 (O_1979,N_14928,N_14950);
or UO_1980 (O_1980,N_14901,N_14948);
nand UO_1981 (O_1981,N_14877,N_14979);
nand UO_1982 (O_1982,N_14944,N_14880);
and UO_1983 (O_1983,N_14885,N_14956);
or UO_1984 (O_1984,N_14875,N_14954);
nand UO_1985 (O_1985,N_14926,N_14893);
nand UO_1986 (O_1986,N_14948,N_14904);
nor UO_1987 (O_1987,N_14944,N_14917);
nor UO_1988 (O_1988,N_14953,N_14964);
and UO_1989 (O_1989,N_14967,N_14923);
nand UO_1990 (O_1990,N_14925,N_14896);
nor UO_1991 (O_1991,N_14893,N_14933);
nand UO_1992 (O_1992,N_14897,N_14903);
xor UO_1993 (O_1993,N_14981,N_14996);
xnor UO_1994 (O_1994,N_14901,N_14963);
nor UO_1995 (O_1995,N_14899,N_14975);
and UO_1996 (O_1996,N_14918,N_14879);
nand UO_1997 (O_1997,N_14965,N_14891);
and UO_1998 (O_1998,N_14928,N_14897);
nor UO_1999 (O_1999,N_14880,N_14941);
endmodule