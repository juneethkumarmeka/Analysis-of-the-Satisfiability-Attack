module basic_500_3000_500_5_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_69,In_291);
and U1 (N_1,In_251,In_482);
or U2 (N_2,In_422,In_155);
or U3 (N_3,In_46,In_295);
nand U4 (N_4,In_309,In_3);
nand U5 (N_5,In_273,In_97);
nand U6 (N_6,In_488,In_497);
or U7 (N_7,In_186,In_411);
and U8 (N_8,In_459,In_337);
nand U9 (N_9,In_384,In_51);
nand U10 (N_10,In_329,In_179);
and U11 (N_11,In_481,In_63);
and U12 (N_12,In_70,In_91);
nand U13 (N_13,In_107,In_338);
nor U14 (N_14,In_156,In_446);
or U15 (N_15,In_55,In_294);
or U16 (N_16,In_456,In_450);
or U17 (N_17,In_374,In_5);
nor U18 (N_18,In_138,In_435);
and U19 (N_19,In_408,In_188);
or U20 (N_20,In_114,In_81);
nand U21 (N_21,In_310,In_150);
or U22 (N_22,In_451,In_161);
and U23 (N_23,In_135,In_204);
nand U24 (N_24,In_230,In_244);
xor U25 (N_25,In_176,In_255);
xor U26 (N_26,In_163,In_203);
nand U27 (N_27,In_217,In_42);
nor U28 (N_28,In_101,In_257);
nand U29 (N_29,In_151,In_166);
nor U30 (N_30,In_202,In_480);
nor U31 (N_31,In_145,In_494);
nand U32 (N_32,In_349,In_298);
nand U33 (N_33,In_22,In_376);
and U34 (N_34,In_245,In_276);
xor U35 (N_35,In_287,In_493);
nand U36 (N_36,In_26,In_261);
xor U37 (N_37,In_127,In_192);
or U38 (N_38,In_316,In_403);
nand U39 (N_39,In_423,In_100);
xor U40 (N_40,In_409,In_312);
nor U41 (N_41,In_79,In_73);
nand U42 (N_42,In_381,In_264);
nor U43 (N_43,In_371,In_102);
nand U44 (N_44,In_327,In_357);
and U45 (N_45,In_36,In_277);
nor U46 (N_46,In_170,In_428);
and U47 (N_47,In_306,In_468);
or U48 (N_48,In_317,In_144);
or U49 (N_49,In_66,In_282);
nor U50 (N_50,In_86,In_486);
and U51 (N_51,In_490,In_333);
nor U52 (N_52,In_142,In_275);
nand U53 (N_53,In_246,In_231);
and U54 (N_54,In_483,In_242);
nor U55 (N_55,In_87,In_302);
nor U56 (N_56,In_475,In_64);
nor U57 (N_57,In_279,In_352);
nor U58 (N_58,In_99,In_15);
or U59 (N_59,In_126,In_199);
and U60 (N_60,In_159,In_14);
nand U61 (N_61,In_44,In_339);
xnor U62 (N_62,In_139,In_375);
xor U63 (N_63,In_28,In_267);
or U64 (N_64,In_141,In_223);
or U65 (N_65,In_94,In_311);
or U66 (N_66,In_346,In_443);
or U67 (N_67,In_303,In_414);
and U68 (N_68,In_72,In_367);
and U69 (N_69,In_247,In_249);
and U70 (N_70,In_62,In_61);
nor U71 (N_71,In_149,In_290);
nor U72 (N_72,In_17,In_189);
or U73 (N_73,In_361,In_53);
nor U74 (N_74,In_196,In_154);
nor U75 (N_75,In_354,In_307);
nand U76 (N_76,In_108,In_413);
or U77 (N_77,In_415,In_392);
nand U78 (N_78,In_129,In_296);
nor U79 (N_79,In_12,In_300);
nor U80 (N_80,In_110,In_308);
and U81 (N_81,In_183,In_104);
nand U82 (N_82,In_85,In_187);
nand U83 (N_83,In_390,In_9);
nand U84 (N_84,In_229,In_165);
and U85 (N_85,In_225,In_118);
or U86 (N_86,In_74,In_334);
nor U87 (N_87,In_436,In_498);
and U88 (N_88,In_11,In_353);
nand U89 (N_89,In_75,In_485);
or U90 (N_90,In_0,In_119);
nand U91 (N_91,In_227,In_132);
or U92 (N_92,In_113,In_343);
and U93 (N_93,In_116,In_226);
nor U94 (N_94,In_274,In_134);
nor U95 (N_95,In_252,In_174);
or U96 (N_96,In_146,In_140);
and U97 (N_97,In_470,In_258);
or U98 (N_98,In_404,In_476);
nor U99 (N_99,In_347,In_454);
nor U100 (N_100,In_467,In_92);
nor U101 (N_101,In_248,In_340);
or U102 (N_102,In_355,In_167);
nor U103 (N_103,In_315,In_40);
and U104 (N_104,In_124,In_181);
nor U105 (N_105,In_350,In_19);
nor U106 (N_106,In_469,In_152);
nor U107 (N_107,In_313,In_172);
nor U108 (N_108,In_211,In_109);
and U109 (N_109,In_331,In_289);
and U110 (N_110,In_236,In_65);
and U111 (N_111,In_373,In_464);
or U112 (N_112,In_366,In_106);
or U113 (N_113,In_499,In_364);
nor U114 (N_114,In_418,In_360);
nand U115 (N_115,In_380,In_173);
and U116 (N_116,In_115,In_128);
nor U117 (N_117,In_356,In_447);
nand U118 (N_118,In_377,In_424);
and U119 (N_119,In_440,In_383);
nand U120 (N_120,In_452,In_38);
and U121 (N_121,In_431,In_35);
nand U122 (N_122,In_260,In_318);
nand U123 (N_123,In_330,In_487);
or U124 (N_124,In_112,In_250);
nand U125 (N_125,In_484,In_175);
nand U126 (N_126,In_228,In_105);
nand U127 (N_127,In_320,In_402);
and U128 (N_128,In_362,In_238);
nand U129 (N_129,In_259,In_365);
and U130 (N_130,In_123,In_269);
and U131 (N_131,In_336,In_299);
and U132 (N_132,In_58,In_263);
and U133 (N_133,In_24,In_213);
nand U134 (N_134,In_496,In_222);
nor U135 (N_135,In_478,In_345);
and U136 (N_136,In_45,In_281);
and U137 (N_137,In_399,In_130);
or U138 (N_138,In_98,In_6);
nor U139 (N_139,In_358,In_253);
and U140 (N_140,In_393,In_344);
or U141 (N_141,In_398,In_368);
or U142 (N_142,In_283,In_216);
or U143 (N_143,In_219,In_412);
and U144 (N_144,In_83,In_180);
or U145 (N_145,In_7,In_2);
and U146 (N_146,In_293,In_406);
nand U147 (N_147,In_465,In_385);
and U148 (N_148,In_18,In_215);
xnor U149 (N_149,In_191,In_492);
nand U150 (N_150,In_270,In_442);
nor U151 (N_151,In_59,In_31);
nor U152 (N_152,In_437,In_444);
nor U153 (N_153,In_438,In_93);
nand U154 (N_154,In_201,In_68);
and U155 (N_155,In_448,In_212);
nor U156 (N_156,In_397,In_241);
and U157 (N_157,In_67,In_471);
or U158 (N_158,In_389,In_265);
nor U159 (N_159,In_474,In_477);
and U160 (N_160,In_41,In_426);
nor U161 (N_161,In_49,In_433);
and U162 (N_162,In_445,In_305);
nand U163 (N_163,In_420,In_158);
and U164 (N_164,In_185,In_271);
nor U165 (N_165,In_164,In_10);
and U166 (N_166,In_221,In_455);
nor U167 (N_167,In_190,In_314);
nor U168 (N_168,In_78,In_495);
xor U169 (N_169,In_233,In_168);
nand U170 (N_170,In_157,In_4);
and U171 (N_171,In_297,In_160);
and U172 (N_172,In_472,In_195);
and U173 (N_173,In_432,In_378);
and U174 (N_174,In_489,In_71);
or U175 (N_175,In_370,In_268);
nor U176 (N_176,In_461,In_326);
xnor U177 (N_177,In_439,In_286);
nand U178 (N_178,In_117,In_30);
nand U179 (N_179,In_218,In_325);
and U180 (N_180,In_278,In_348);
nand U181 (N_181,In_209,In_20);
or U182 (N_182,In_88,In_388);
and U183 (N_183,In_205,In_200);
nand U184 (N_184,In_429,In_272);
nor U185 (N_185,In_232,In_405);
and U186 (N_186,In_194,In_60);
and U187 (N_187,In_491,In_33);
and U188 (N_188,In_453,In_80);
nand U189 (N_189,In_319,In_162);
or U190 (N_190,In_103,In_23);
or U191 (N_191,In_43,In_285);
nand U192 (N_192,In_147,In_198);
or U193 (N_193,In_284,In_396);
xnor U194 (N_194,In_430,In_54);
and U195 (N_195,In_256,In_13);
or U196 (N_196,In_214,In_341);
nand U197 (N_197,In_449,In_137);
or U198 (N_198,In_280,In_29);
nand U199 (N_199,In_458,In_56);
or U200 (N_200,In_16,In_133);
nand U201 (N_201,In_125,In_419);
xor U202 (N_202,In_153,In_359);
nand U203 (N_203,In_34,In_441);
and U204 (N_204,In_235,In_21);
nor U205 (N_205,In_410,In_466);
or U206 (N_206,In_328,In_322);
or U207 (N_207,In_8,In_425);
and U208 (N_208,In_131,In_351);
and U209 (N_209,In_76,In_234);
or U210 (N_210,In_479,In_394);
nand U211 (N_211,In_84,In_395);
nor U212 (N_212,In_120,In_473);
nor U213 (N_213,In_266,In_89);
or U214 (N_214,In_1,In_90);
or U215 (N_215,In_169,In_324);
nor U216 (N_216,In_121,In_143);
or U217 (N_217,In_210,In_47);
nor U218 (N_218,In_184,In_37);
and U219 (N_219,In_292,In_379);
and U220 (N_220,In_382,In_335);
nor U221 (N_221,In_27,In_421);
nor U222 (N_222,In_240,In_206);
or U223 (N_223,In_52,In_457);
nor U224 (N_224,In_178,In_288);
or U225 (N_225,In_369,In_363);
nor U226 (N_226,In_323,In_224);
or U227 (N_227,In_460,In_342);
and U228 (N_228,In_182,In_332);
nand U229 (N_229,In_462,In_401);
and U230 (N_230,In_136,In_197);
and U231 (N_231,In_463,In_148);
nor U232 (N_232,In_386,In_177);
or U233 (N_233,In_207,In_262);
or U234 (N_234,In_96,In_48);
or U235 (N_235,In_32,In_82);
nand U236 (N_236,In_77,In_321);
or U237 (N_237,In_193,In_301);
or U238 (N_238,In_400,In_372);
or U239 (N_239,In_171,In_254);
and U240 (N_240,In_427,In_111);
nor U241 (N_241,In_208,In_417);
or U242 (N_242,In_407,In_122);
nand U243 (N_243,In_239,In_57);
and U244 (N_244,In_39,In_50);
nand U245 (N_245,In_95,In_416);
or U246 (N_246,In_304,In_243);
nand U247 (N_247,In_434,In_387);
nand U248 (N_248,In_391,In_25);
nand U249 (N_249,In_237,In_220);
and U250 (N_250,In_172,In_38);
nor U251 (N_251,In_70,In_459);
or U252 (N_252,In_348,In_359);
or U253 (N_253,In_351,In_354);
or U254 (N_254,In_460,In_11);
nand U255 (N_255,In_36,In_232);
nor U256 (N_256,In_315,In_234);
nand U257 (N_257,In_195,In_92);
and U258 (N_258,In_206,In_65);
nor U259 (N_259,In_240,In_441);
nor U260 (N_260,In_192,In_349);
nand U261 (N_261,In_450,In_127);
nor U262 (N_262,In_56,In_372);
or U263 (N_263,In_145,In_89);
or U264 (N_264,In_95,In_97);
or U265 (N_265,In_452,In_439);
or U266 (N_266,In_274,In_424);
nand U267 (N_267,In_38,In_183);
nor U268 (N_268,In_398,In_371);
nand U269 (N_269,In_274,In_61);
or U270 (N_270,In_405,In_213);
and U271 (N_271,In_221,In_492);
and U272 (N_272,In_193,In_317);
and U273 (N_273,In_490,In_314);
nor U274 (N_274,In_246,In_355);
nor U275 (N_275,In_356,In_358);
or U276 (N_276,In_496,In_54);
or U277 (N_277,In_38,In_345);
nand U278 (N_278,In_238,In_460);
nor U279 (N_279,In_426,In_431);
nand U280 (N_280,In_390,In_273);
nor U281 (N_281,In_69,In_385);
or U282 (N_282,In_204,In_106);
nor U283 (N_283,In_392,In_383);
and U284 (N_284,In_339,In_145);
nor U285 (N_285,In_87,In_216);
nand U286 (N_286,In_7,In_201);
nor U287 (N_287,In_228,In_418);
or U288 (N_288,In_132,In_428);
xor U289 (N_289,In_52,In_23);
nand U290 (N_290,In_373,In_30);
or U291 (N_291,In_403,In_199);
nor U292 (N_292,In_180,In_171);
xor U293 (N_293,In_155,In_363);
nor U294 (N_294,In_62,In_79);
or U295 (N_295,In_62,In_446);
and U296 (N_296,In_391,In_2);
and U297 (N_297,In_164,In_234);
nand U298 (N_298,In_477,In_48);
and U299 (N_299,In_386,In_461);
or U300 (N_300,In_357,In_370);
and U301 (N_301,In_405,In_289);
nand U302 (N_302,In_116,In_86);
or U303 (N_303,In_297,In_74);
and U304 (N_304,In_57,In_353);
and U305 (N_305,In_214,In_457);
and U306 (N_306,In_314,In_404);
and U307 (N_307,In_268,In_226);
nor U308 (N_308,In_48,In_173);
or U309 (N_309,In_216,In_245);
nand U310 (N_310,In_322,In_301);
nor U311 (N_311,In_7,In_17);
nand U312 (N_312,In_278,In_100);
and U313 (N_313,In_93,In_164);
and U314 (N_314,In_485,In_441);
nor U315 (N_315,In_174,In_380);
or U316 (N_316,In_307,In_352);
nor U317 (N_317,In_393,In_279);
nor U318 (N_318,In_325,In_492);
nor U319 (N_319,In_41,In_98);
nand U320 (N_320,In_185,In_487);
xnor U321 (N_321,In_261,In_28);
nor U322 (N_322,In_295,In_452);
nand U323 (N_323,In_456,In_43);
and U324 (N_324,In_69,In_441);
or U325 (N_325,In_365,In_230);
nand U326 (N_326,In_222,In_378);
nand U327 (N_327,In_309,In_278);
or U328 (N_328,In_289,In_272);
and U329 (N_329,In_422,In_89);
and U330 (N_330,In_475,In_345);
nor U331 (N_331,In_346,In_404);
and U332 (N_332,In_143,In_32);
nand U333 (N_333,In_273,In_299);
nor U334 (N_334,In_291,In_475);
and U335 (N_335,In_170,In_266);
nor U336 (N_336,In_240,In_487);
or U337 (N_337,In_197,In_248);
nand U338 (N_338,In_341,In_442);
or U339 (N_339,In_102,In_453);
or U340 (N_340,In_106,In_193);
and U341 (N_341,In_161,In_194);
nand U342 (N_342,In_21,In_341);
or U343 (N_343,In_101,In_31);
or U344 (N_344,In_477,In_181);
nand U345 (N_345,In_383,In_174);
nor U346 (N_346,In_43,In_365);
nand U347 (N_347,In_35,In_331);
nand U348 (N_348,In_338,In_41);
nand U349 (N_349,In_132,In_221);
xnor U350 (N_350,In_203,In_310);
and U351 (N_351,In_207,In_205);
or U352 (N_352,In_344,In_384);
xnor U353 (N_353,In_165,In_248);
or U354 (N_354,In_258,In_375);
and U355 (N_355,In_252,In_345);
or U356 (N_356,In_385,In_420);
and U357 (N_357,In_336,In_322);
nand U358 (N_358,In_480,In_145);
nand U359 (N_359,In_161,In_22);
nor U360 (N_360,In_373,In_429);
xor U361 (N_361,In_474,In_442);
and U362 (N_362,In_46,In_71);
nor U363 (N_363,In_72,In_45);
nor U364 (N_364,In_162,In_155);
and U365 (N_365,In_173,In_441);
nand U366 (N_366,In_152,In_311);
and U367 (N_367,In_264,In_329);
nand U368 (N_368,In_173,In_298);
nand U369 (N_369,In_351,In_300);
or U370 (N_370,In_98,In_84);
nor U371 (N_371,In_333,In_23);
and U372 (N_372,In_264,In_219);
nand U373 (N_373,In_286,In_60);
nand U374 (N_374,In_36,In_126);
or U375 (N_375,In_311,In_163);
and U376 (N_376,In_439,In_132);
nor U377 (N_377,In_371,In_173);
nor U378 (N_378,In_41,In_184);
and U379 (N_379,In_440,In_303);
and U380 (N_380,In_251,In_408);
and U381 (N_381,In_57,In_414);
and U382 (N_382,In_479,In_313);
or U383 (N_383,In_142,In_8);
or U384 (N_384,In_95,In_105);
nand U385 (N_385,In_426,In_60);
and U386 (N_386,In_408,In_497);
nand U387 (N_387,In_232,In_463);
xor U388 (N_388,In_160,In_405);
nand U389 (N_389,In_450,In_305);
nand U390 (N_390,In_3,In_380);
and U391 (N_391,In_15,In_132);
nor U392 (N_392,In_434,In_285);
and U393 (N_393,In_16,In_420);
nor U394 (N_394,In_36,In_86);
nor U395 (N_395,In_439,In_334);
or U396 (N_396,In_474,In_466);
and U397 (N_397,In_155,In_330);
and U398 (N_398,In_221,In_495);
nand U399 (N_399,In_111,In_72);
nand U400 (N_400,In_419,In_378);
or U401 (N_401,In_134,In_229);
xor U402 (N_402,In_234,In_290);
and U403 (N_403,In_213,In_1);
or U404 (N_404,In_280,In_458);
and U405 (N_405,In_188,In_68);
and U406 (N_406,In_396,In_450);
or U407 (N_407,In_18,In_220);
or U408 (N_408,In_220,In_460);
or U409 (N_409,In_50,In_135);
nand U410 (N_410,In_287,In_238);
nand U411 (N_411,In_189,In_144);
nand U412 (N_412,In_209,In_313);
nor U413 (N_413,In_170,In_150);
xor U414 (N_414,In_254,In_196);
nor U415 (N_415,In_12,In_143);
or U416 (N_416,In_183,In_145);
and U417 (N_417,In_65,In_286);
nor U418 (N_418,In_270,In_348);
nor U419 (N_419,In_335,In_47);
nor U420 (N_420,In_414,In_167);
nor U421 (N_421,In_356,In_279);
and U422 (N_422,In_199,In_129);
nor U423 (N_423,In_302,In_296);
xor U424 (N_424,In_414,In_93);
or U425 (N_425,In_155,In_59);
nor U426 (N_426,In_359,In_398);
or U427 (N_427,In_173,In_190);
or U428 (N_428,In_272,In_228);
nand U429 (N_429,In_225,In_423);
or U430 (N_430,In_281,In_472);
xor U431 (N_431,In_92,In_368);
and U432 (N_432,In_91,In_426);
nand U433 (N_433,In_87,In_53);
nand U434 (N_434,In_312,In_402);
or U435 (N_435,In_408,In_212);
and U436 (N_436,In_155,In_451);
nand U437 (N_437,In_27,In_0);
xor U438 (N_438,In_219,In_91);
nor U439 (N_439,In_106,In_477);
nor U440 (N_440,In_348,In_211);
nor U441 (N_441,In_57,In_113);
or U442 (N_442,In_390,In_144);
or U443 (N_443,In_207,In_386);
and U444 (N_444,In_71,In_441);
and U445 (N_445,In_403,In_432);
xnor U446 (N_446,In_103,In_259);
nor U447 (N_447,In_123,In_317);
or U448 (N_448,In_209,In_9);
and U449 (N_449,In_331,In_338);
or U450 (N_450,In_37,In_170);
and U451 (N_451,In_16,In_135);
nor U452 (N_452,In_251,In_388);
and U453 (N_453,In_420,In_182);
and U454 (N_454,In_390,In_355);
nor U455 (N_455,In_381,In_290);
or U456 (N_456,In_39,In_86);
and U457 (N_457,In_42,In_416);
or U458 (N_458,In_252,In_320);
nor U459 (N_459,In_45,In_74);
and U460 (N_460,In_460,In_428);
or U461 (N_461,In_198,In_410);
or U462 (N_462,In_56,In_382);
nor U463 (N_463,In_19,In_442);
and U464 (N_464,In_300,In_327);
and U465 (N_465,In_12,In_442);
nand U466 (N_466,In_345,In_268);
nand U467 (N_467,In_89,In_498);
nor U468 (N_468,In_294,In_138);
xor U469 (N_469,In_289,In_330);
or U470 (N_470,In_60,In_332);
or U471 (N_471,In_324,In_327);
or U472 (N_472,In_7,In_112);
and U473 (N_473,In_93,In_281);
and U474 (N_474,In_20,In_107);
and U475 (N_475,In_40,In_55);
or U476 (N_476,In_27,In_335);
nor U477 (N_477,In_421,In_124);
nand U478 (N_478,In_117,In_253);
nand U479 (N_479,In_480,In_221);
xnor U480 (N_480,In_88,In_228);
nand U481 (N_481,In_272,In_73);
or U482 (N_482,In_33,In_441);
and U483 (N_483,In_450,In_275);
and U484 (N_484,In_238,In_139);
or U485 (N_485,In_68,In_80);
and U486 (N_486,In_287,In_170);
nor U487 (N_487,In_409,In_51);
nand U488 (N_488,In_338,In_234);
or U489 (N_489,In_46,In_370);
and U490 (N_490,In_31,In_385);
nand U491 (N_491,In_134,In_222);
nand U492 (N_492,In_46,In_134);
and U493 (N_493,In_392,In_423);
nor U494 (N_494,In_450,In_118);
or U495 (N_495,In_427,In_117);
and U496 (N_496,In_460,In_472);
nand U497 (N_497,In_362,In_52);
and U498 (N_498,In_81,In_332);
or U499 (N_499,In_243,In_492);
nor U500 (N_500,In_325,In_421);
or U501 (N_501,In_464,In_7);
nand U502 (N_502,In_5,In_210);
nor U503 (N_503,In_283,In_18);
and U504 (N_504,In_55,In_107);
xnor U505 (N_505,In_196,In_204);
and U506 (N_506,In_93,In_4);
or U507 (N_507,In_189,In_245);
nand U508 (N_508,In_59,In_176);
nand U509 (N_509,In_322,In_305);
or U510 (N_510,In_475,In_376);
and U511 (N_511,In_11,In_303);
nor U512 (N_512,In_308,In_257);
nand U513 (N_513,In_387,In_104);
nand U514 (N_514,In_418,In_23);
and U515 (N_515,In_236,In_374);
nor U516 (N_516,In_342,In_185);
nor U517 (N_517,In_364,In_241);
and U518 (N_518,In_38,In_308);
and U519 (N_519,In_385,In_261);
nor U520 (N_520,In_280,In_305);
or U521 (N_521,In_332,In_355);
nand U522 (N_522,In_443,In_427);
nor U523 (N_523,In_140,In_105);
nand U524 (N_524,In_126,In_10);
nor U525 (N_525,In_468,In_193);
nand U526 (N_526,In_192,In_324);
nand U527 (N_527,In_323,In_32);
nor U528 (N_528,In_229,In_278);
or U529 (N_529,In_265,In_195);
or U530 (N_530,In_463,In_196);
nand U531 (N_531,In_361,In_130);
or U532 (N_532,In_89,In_251);
nor U533 (N_533,In_42,In_496);
nand U534 (N_534,In_319,In_173);
or U535 (N_535,In_392,In_335);
and U536 (N_536,In_68,In_171);
or U537 (N_537,In_300,In_238);
and U538 (N_538,In_237,In_365);
or U539 (N_539,In_460,In_252);
or U540 (N_540,In_239,In_23);
nor U541 (N_541,In_145,In_338);
and U542 (N_542,In_9,In_203);
nand U543 (N_543,In_249,In_265);
nand U544 (N_544,In_161,In_368);
nand U545 (N_545,In_473,In_371);
or U546 (N_546,In_486,In_36);
or U547 (N_547,In_450,In_115);
or U548 (N_548,In_284,In_34);
or U549 (N_549,In_48,In_29);
nor U550 (N_550,In_72,In_113);
nor U551 (N_551,In_215,In_323);
nand U552 (N_552,In_142,In_174);
or U553 (N_553,In_48,In_231);
nor U554 (N_554,In_348,In_454);
and U555 (N_555,In_488,In_96);
nor U556 (N_556,In_452,In_50);
and U557 (N_557,In_149,In_105);
xor U558 (N_558,In_99,In_495);
nand U559 (N_559,In_127,In_260);
and U560 (N_560,In_410,In_189);
nor U561 (N_561,In_398,In_222);
xor U562 (N_562,In_319,In_158);
and U563 (N_563,In_143,In_139);
or U564 (N_564,In_236,In_316);
nand U565 (N_565,In_107,In_202);
and U566 (N_566,In_347,In_111);
nand U567 (N_567,In_54,In_3);
nand U568 (N_568,In_76,In_417);
and U569 (N_569,In_387,In_21);
and U570 (N_570,In_59,In_274);
nor U571 (N_571,In_316,In_119);
nand U572 (N_572,In_290,In_76);
or U573 (N_573,In_84,In_303);
and U574 (N_574,In_285,In_238);
or U575 (N_575,In_440,In_496);
nand U576 (N_576,In_7,In_296);
and U577 (N_577,In_279,In_1);
and U578 (N_578,In_17,In_237);
nand U579 (N_579,In_51,In_325);
nand U580 (N_580,In_78,In_215);
nand U581 (N_581,In_472,In_187);
and U582 (N_582,In_32,In_215);
nand U583 (N_583,In_356,In_138);
or U584 (N_584,In_267,In_246);
nand U585 (N_585,In_168,In_98);
and U586 (N_586,In_468,In_362);
and U587 (N_587,In_445,In_492);
nand U588 (N_588,In_186,In_164);
nand U589 (N_589,In_376,In_367);
nor U590 (N_590,In_88,In_456);
nand U591 (N_591,In_486,In_143);
or U592 (N_592,In_478,In_448);
and U593 (N_593,In_357,In_140);
and U594 (N_594,In_447,In_440);
and U595 (N_595,In_183,In_420);
or U596 (N_596,In_463,In_362);
nand U597 (N_597,In_178,In_63);
nand U598 (N_598,In_127,In_279);
nand U599 (N_599,In_381,In_240);
and U600 (N_600,N_54,N_527);
nor U601 (N_601,N_298,N_550);
nand U602 (N_602,N_237,N_377);
nor U603 (N_603,N_347,N_161);
or U604 (N_604,N_22,N_339);
nand U605 (N_605,N_313,N_129);
nor U606 (N_606,N_352,N_62);
nand U607 (N_607,N_366,N_429);
and U608 (N_608,N_506,N_461);
and U609 (N_609,N_346,N_335);
nand U610 (N_610,N_547,N_189);
and U611 (N_611,N_583,N_584);
nand U612 (N_612,N_540,N_331);
nand U613 (N_613,N_78,N_211);
or U614 (N_614,N_172,N_100);
and U615 (N_615,N_576,N_254);
nor U616 (N_616,N_76,N_350);
or U617 (N_617,N_525,N_230);
nor U618 (N_618,N_521,N_68);
nand U619 (N_619,N_316,N_480);
nor U620 (N_620,N_288,N_191);
nand U621 (N_621,N_504,N_198);
or U622 (N_622,N_408,N_369);
or U623 (N_623,N_397,N_260);
nand U624 (N_624,N_505,N_487);
nand U625 (N_625,N_12,N_194);
nand U626 (N_626,N_243,N_577);
nand U627 (N_627,N_107,N_588);
nand U628 (N_628,N_482,N_184);
nand U629 (N_629,N_122,N_102);
nor U630 (N_630,N_465,N_249);
nand U631 (N_631,N_187,N_97);
or U632 (N_632,N_595,N_53);
nand U633 (N_633,N_45,N_72);
nor U634 (N_634,N_61,N_182);
xor U635 (N_635,N_312,N_579);
nand U636 (N_636,N_493,N_291);
nand U637 (N_637,N_455,N_532);
xor U638 (N_638,N_570,N_209);
nand U639 (N_639,N_150,N_565);
nor U640 (N_640,N_267,N_474);
and U641 (N_641,N_227,N_178);
nand U642 (N_642,N_195,N_158);
and U643 (N_643,N_40,N_420);
or U644 (N_644,N_58,N_30);
or U645 (N_645,N_293,N_35);
nor U646 (N_646,N_370,N_274);
xnor U647 (N_647,N_485,N_520);
nand U648 (N_648,N_250,N_19);
nand U649 (N_649,N_305,N_326);
and U650 (N_650,N_446,N_435);
nand U651 (N_651,N_507,N_134);
and U652 (N_652,N_73,N_476);
nand U653 (N_653,N_546,N_411);
and U654 (N_654,N_387,N_327);
and U655 (N_655,N_549,N_558);
or U656 (N_656,N_89,N_221);
or U657 (N_657,N_426,N_509);
nor U658 (N_658,N_141,N_497);
or U659 (N_659,N_29,N_373);
nand U660 (N_660,N_591,N_333);
nand U661 (N_661,N_475,N_283);
nand U662 (N_662,N_578,N_124);
and U663 (N_663,N_399,N_304);
nor U664 (N_664,N_155,N_207);
nor U665 (N_665,N_186,N_568);
nor U666 (N_666,N_265,N_382);
nor U667 (N_667,N_270,N_77);
and U668 (N_668,N_431,N_121);
nand U669 (N_669,N_197,N_167);
or U670 (N_670,N_92,N_323);
xor U671 (N_671,N_324,N_38);
or U672 (N_672,N_93,N_136);
nand U673 (N_673,N_33,N_552);
nor U674 (N_674,N_39,N_363);
nand U675 (N_675,N_244,N_164);
nand U676 (N_676,N_587,N_71);
nor U677 (N_677,N_135,N_553);
nand U678 (N_678,N_179,N_496);
nand U679 (N_679,N_137,N_126);
xnor U680 (N_680,N_433,N_18);
and U681 (N_681,N_364,N_534);
and U682 (N_682,N_241,N_372);
nor U683 (N_683,N_147,N_300);
nand U684 (N_684,N_282,N_251);
or U685 (N_685,N_87,N_59);
nand U686 (N_686,N_310,N_36);
and U687 (N_687,N_359,N_543);
and U688 (N_688,N_545,N_398);
nand U689 (N_689,N_539,N_119);
nor U690 (N_690,N_127,N_320);
and U691 (N_691,N_206,N_556);
or U692 (N_692,N_166,N_13);
and U693 (N_693,N_392,N_538);
and U694 (N_694,N_290,N_60);
nor U695 (N_695,N_342,N_81);
nand U696 (N_696,N_371,N_6);
or U697 (N_697,N_245,N_569);
or U698 (N_698,N_64,N_152);
or U699 (N_699,N_586,N_319);
and U700 (N_700,N_139,N_389);
and U701 (N_701,N_456,N_385);
nor U702 (N_702,N_1,N_308);
nor U703 (N_703,N_303,N_463);
nand U704 (N_704,N_458,N_99);
xor U705 (N_705,N_355,N_44);
nand U706 (N_706,N_55,N_390);
nand U707 (N_707,N_101,N_512);
and U708 (N_708,N_357,N_31);
nor U709 (N_709,N_272,N_516);
nand U710 (N_710,N_526,N_544);
nand U711 (N_711,N_515,N_354);
nor U712 (N_712,N_548,N_380);
nand U713 (N_713,N_154,N_306);
nor U714 (N_714,N_378,N_572);
or U715 (N_715,N_502,N_199);
and U716 (N_716,N_278,N_74);
and U717 (N_717,N_598,N_103);
nand U718 (N_718,N_48,N_84);
xnor U719 (N_719,N_314,N_560);
nor U720 (N_720,N_315,N_405);
nor U721 (N_721,N_273,N_330);
and U722 (N_722,N_110,N_460);
nor U723 (N_723,N_34,N_451);
and U724 (N_724,N_383,N_177);
and U725 (N_725,N_535,N_70);
and U726 (N_726,N_384,N_518);
xnor U727 (N_727,N_555,N_296);
or U728 (N_728,N_400,N_201);
and U729 (N_729,N_340,N_428);
nor U730 (N_730,N_111,N_138);
xnor U731 (N_731,N_449,N_542);
xor U732 (N_732,N_285,N_275);
nand U733 (N_733,N_489,N_156);
or U734 (N_734,N_286,N_90);
or U735 (N_735,N_256,N_259);
nand U736 (N_736,N_318,N_7);
nor U737 (N_737,N_344,N_453);
nor U738 (N_738,N_188,N_334);
nor U739 (N_739,N_143,N_203);
nor U740 (N_740,N_240,N_566);
nand U741 (N_741,N_128,N_541);
xor U742 (N_742,N_348,N_168);
nor U743 (N_743,N_503,N_105);
nand U744 (N_744,N_358,N_551);
nor U745 (N_745,N_14,N_50);
nor U746 (N_746,N_477,N_528);
or U747 (N_747,N_263,N_287);
xnor U748 (N_748,N_403,N_567);
and U749 (N_749,N_442,N_153);
or U750 (N_750,N_356,N_115);
nand U751 (N_751,N_94,N_24);
and U752 (N_752,N_106,N_581);
nor U753 (N_753,N_501,N_401);
or U754 (N_754,N_322,N_266);
or U755 (N_755,N_220,N_479);
or U756 (N_756,N_471,N_88);
or U757 (N_757,N_95,N_261);
or U758 (N_758,N_216,N_145);
or U759 (N_759,N_83,N_554);
nor U760 (N_760,N_268,N_590);
and U761 (N_761,N_255,N_146);
nor U762 (N_762,N_91,N_599);
or U763 (N_763,N_589,N_452);
and U764 (N_764,N_75,N_473);
nor U765 (N_765,N_557,N_430);
nand U766 (N_766,N_478,N_297);
nor U767 (N_767,N_65,N_580);
and U768 (N_768,N_46,N_404);
nor U769 (N_769,N_171,N_522);
nand U770 (N_770,N_8,N_269);
nor U771 (N_771,N_441,N_204);
nand U772 (N_772,N_537,N_183);
nand U773 (N_773,N_294,N_160);
nand U774 (N_774,N_32,N_112);
nand U775 (N_775,N_360,N_459);
and U776 (N_776,N_375,N_181);
or U777 (N_777,N_381,N_5);
and U778 (N_778,N_3,N_10);
nor U779 (N_779,N_328,N_500);
and U780 (N_780,N_511,N_226);
nor U781 (N_781,N_394,N_151);
nor U782 (N_782,N_190,N_142);
nand U783 (N_783,N_409,N_585);
or U784 (N_784,N_117,N_130);
nand U785 (N_785,N_510,N_529);
xor U786 (N_786,N_531,N_422);
or U787 (N_787,N_486,N_213);
nor U788 (N_788,N_440,N_281);
nand U789 (N_789,N_174,N_321);
and U790 (N_790,N_574,N_225);
or U791 (N_791,N_133,N_448);
and U792 (N_792,N_594,N_63);
or U793 (N_793,N_214,N_0);
or U794 (N_794,N_462,N_436);
nor U795 (N_795,N_262,N_11);
nor U796 (N_796,N_447,N_593);
nand U797 (N_797,N_271,N_341);
or U798 (N_798,N_193,N_242);
and U799 (N_799,N_118,N_402);
nand U800 (N_800,N_393,N_337);
or U801 (N_801,N_301,N_86);
nor U802 (N_802,N_571,N_311);
nor U803 (N_803,N_116,N_407);
or U804 (N_804,N_210,N_562);
nand U805 (N_805,N_332,N_239);
or U806 (N_806,N_80,N_376);
or U807 (N_807,N_252,N_98);
or U808 (N_808,N_247,N_425);
nand U809 (N_809,N_434,N_231);
nor U810 (N_810,N_472,N_597);
and U811 (N_811,N_57,N_484);
nor U812 (N_812,N_162,N_343);
nand U813 (N_813,N_492,N_236);
or U814 (N_814,N_196,N_564);
nand U815 (N_815,N_148,N_444);
xor U816 (N_816,N_66,N_217);
nor U817 (N_817,N_445,N_176);
and U818 (N_818,N_144,N_533);
and U819 (N_819,N_365,N_212);
nor U820 (N_820,N_253,N_28);
and U821 (N_821,N_386,N_9);
nand U822 (N_822,N_495,N_395);
or U823 (N_823,N_284,N_41);
nand U824 (N_824,N_16,N_43);
or U825 (N_825,N_424,N_416);
or U826 (N_826,N_292,N_450);
and U827 (N_827,N_185,N_51);
nor U828 (N_828,N_222,N_325);
nand U829 (N_829,N_257,N_170);
nor U830 (N_830,N_192,N_163);
nand U831 (N_831,N_361,N_519);
nand U832 (N_832,N_469,N_396);
nor U833 (N_833,N_439,N_559);
nor U834 (N_834,N_517,N_498);
or U835 (N_835,N_349,N_468);
nor U836 (N_836,N_466,N_362);
and U837 (N_837,N_218,N_582);
or U838 (N_838,N_229,N_317);
and U839 (N_839,N_248,N_596);
and U840 (N_840,N_47,N_427);
or U841 (N_841,N_488,N_329);
or U842 (N_842,N_17,N_125);
nand U843 (N_843,N_494,N_219);
or U844 (N_844,N_406,N_20);
or U845 (N_845,N_418,N_2);
or U846 (N_846,N_454,N_26);
or U847 (N_847,N_21,N_96);
nor U848 (N_848,N_464,N_23);
or U849 (N_849,N_52,N_419);
and U850 (N_850,N_367,N_309);
xor U851 (N_851,N_200,N_25);
and U852 (N_852,N_467,N_490);
nor U853 (N_853,N_246,N_353);
or U854 (N_854,N_85,N_432);
nand U855 (N_855,N_421,N_514);
nor U856 (N_856,N_561,N_276);
nand U857 (N_857,N_295,N_491);
nand U858 (N_858,N_499,N_113);
nor U859 (N_859,N_338,N_345);
or U860 (N_860,N_412,N_223);
nand U861 (N_861,N_523,N_592);
nor U862 (N_862,N_279,N_299);
and U863 (N_863,N_289,N_205);
nor U864 (N_864,N_109,N_438);
nor U865 (N_865,N_280,N_208);
xnor U866 (N_866,N_202,N_49);
nor U867 (N_867,N_513,N_258);
nor U868 (N_868,N_224,N_368);
or U869 (N_869,N_481,N_413);
nor U870 (N_870,N_120,N_108);
nor U871 (N_871,N_42,N_336);
nand U872 (N_872,N_159,N_4);
nor U873 (N_873,N_573,N_157);
nor U874 (N_874,N_232,N_234);
nand U875 (N_875,N_173,N_379);
nor U876 (N_876,N_82,N_391);
or U877 (N_877,N_351,N_417);
nand U878 (N_878,N_123,N_410);
nor U879 (N_879,N_423,N_56);
or U880 (N_880,N_508,N_175);
or U881 (N_881,N_536,N_215);
nand U882 (N_882,N_563,N_414);
or U883 (N_883,N_15,N_470);
nor U884 (N_884,N_374,N_69);
or U885 (N_885,N_437,N_238);
nand U886 (N_886,N_483,N_277);
or U887 (N_887,N_530,N_67);
nand U888 (N_888,N_37,N_235);
nand U889 (N_889,N_307,N_131);
and U890 (N_890,N_264,N_104);
or U891 (N_891,N_149,N_169);
nor U892 (N_892,N_114,N_524);
and U893 (N_893,N_233,N_27);
nand U894 (N_894,N_457,N_79);
and U895 (N_895,N_165,N_415);
or U896 (N_896,N_180,N_575);
nand U897 (N_897,N_228,N_140);
nand U898 (N_898,N_388,N_132);
and U899 (N_899,N_302,N_443);
and U900 (N_900,N_109,N_577);
nand U901 (N_901,N_162,N_145);
or U902 (N_902,N_276,N_162);
and U903 (N_903,N_155,N_11);
nand U904 (N_904,N_207,N_414);
and U905 (N_905,N_60,N_398);
and U906 (N_906,N_251,N_549);
xnor U907 (N_907,N_268,N_177);
or U908 (N_908,N_528,N_54);
and U909 (N_909,N_514,N_117);
or U910 (N_910,N_5,N_481);
nand U911 (N_911,N_422,N_436);
or U912 (N_912,N_159,N_527);
and U913 (N_913,N_399,N_427);
and U914 (N_914,N_126,N_152);
or U915 (N_915,N_122,N_51);
and U916 (N_916,N_560,N_296);
nand U917 (N_917,N_330,N_58);
and U918 (N_918,N_250,N_424);
and U919 (N_919,N_40,N_589);
nand U920 (N_920,N_466,N_152);
and U921 (N_921,N_216,N_565);
nor U922 (N_922,N_428,N_98);
nor U923 (N_923,N_569,N_142);
nor U924 (N_924,N_373,N_354);
and U925 (N_925,N_356,N_308);
nand U926 (N_926,N_218,N_392);
or U927 (N_927,N_267,N_597);
nor U928 (N_928,N_447,N_125);
nor U929 (N_929,N_238,N_337);
or U930 (N_930,N_526,N_179);
nand U931 (N_931,N_154,N_360);
nand U932 (N_932,N_343,N_426);
nand U933 (N_933,N_128,N_129);
nor U934 (N_934,N_302,N_534);
or U935 (N_935,N_425,N_1);
nand U936 (N_936,N_229,N_487);
nor U937 (N_937,N_482,N_430);
nand U938 (N_938,N_70,N_116);
nor U939 (N_939,N_121,N_98);
or U940 (N_940,N_266,N_320);
and U941 (N_941,N_111,N_295);
xor U942 (N_942,N_134,N_572);
or U943 (N_943,N_379,N_52);
nor U944 (N_944,N_163,N_482);
nor U945 (N_945,N_308,N_376);
and U946 (N_946,N_76,N_327);
and U947 (N_947,N_496,N_412);
and U948 (N_948,N_445,N_223);
nor U949 (N_949,N_499,N_79);
or U950 (N_950,N_23,N_394);
nor U951 (N_951,N_553,N_346);
nand U952 (N_952,N_480,N_134);
nand U953 (N_953,N_320,N_573);
nor U954 (N_954,N_469,N_231);
nand U955 (N_955,N_34,N_560);
or U956 (N_956,N_123,N_112);
or U957 (N_957,N_230,N_384);
or U958 (N_958,N_463,N_71);
nand U959 (N_959,N_242,N_570);
or U960 (N_960,N_204,N_71);
nand U961 (N_961,N_521,N_421);
nor U962 (N_962,N_328,N_64);
or U963 (N_963,N_431,N_332);
or U964 (N_964,N_104,N_252);
nor U965 (N_965,N_192,N_414);
and U966 (N_966,N_130,N_125);
nand U967 (N_967,N_129,N_386);
and U968 (N_968,N_138,N_576);
nor U969 (N_969,N_472,N_393);
and U970 (N_970,N_345,N_313);
nand U971 (N_971,N_588,N_131);
and U972 (N_972,N_261,N_519);
or U973 (N_973,N_278,N_176);
nand U974 (N_974,N_166,N_238);
or U975 (N_975,N_142,N_90);
or U976 (N_976,N_274,N_343);
or U977 (N_977,N_143,N_225);
nor U978 (N_978,N_331,N_72);
or U979 (N_979,N_523,N_79);
nor U980 (N_980,N_559,N_435);
and U981 (N_981,N_264,N_455);
nand U982 (N_982,N_39,N_20);
nand U983 (N_983,N_76,N_309);
nand U984 (N_984,N_347,N_222);
or U985 (N_985,N_526,N_259);
nor U986 (N_986,N_109,N_47);
and U987 (N_987,N_346,N_440);
nand U988 (N_988,N_77,N_1);
and U989 (N_989,N_387,N_508);
nor U990 (N_990,N_120,N_586);
nand U991 (N_991,N_292,N_519);
or U992 (N_992,N_356,N_243);
and U993 (N_993,N_270,N_109);
and U994 (N_994,N_61,N_121);
nand U995 (N_995,N_375,N_161);
nor U996 (N_996,N_436,N_15);
nand U997 (N_997,N_76,N_104);
nor U998 (N_998,N_277,N_519);
nand U999 (N_999,N_186,N_294);
nand U1000 (N_1000,N_151,N_547);
nand U1001 (N_1001,N_320,N_342);
and U1002 (N_1002,N_70,N_72);
and U1003 (N_1003,N_193,N_309);
and U1004 (N_1004,N_8,N_18);
or U1005 (N_1005,N_278,N_556);
nand U1006 (N_1006,N_300,N_203);
or U1007 (N_1007,N_152,N_409);
and U1008 (N_1008,N_46,N_517);
or U1009 (N_1009,N_139,N_303);
and U1010 (N_1010,N_372,N_30);
and U1011 (N_1011,N_193,N_148);
and U1012 (N_1012,N_403,N_60);
nand U1013 (N_1013,N_109,N_291);
nand U1014 (N_1014,N_344,N_560);
or U1015 (N_1015,N_286,N_82);
and U1016 (N_1016,N_542,N_9);
or U1017 (N_1017,N_551,N_66);
nand U1018 (N_1018,N_225,N_575);
nand U1019 (N_1019,N_255,N_152);
or U1020 (N_1020,N_340,N_48);
nand U1021 (N_1021,N_138,N_34);
nor U1022 (N_1022,N_46,N_429);
and U1023 (N_1023,N_272,N_251);
and U1024 (N_1024,N_354,N_307);
or U1025 (N_1025,N_579,N_241);
nor U1026 (N_1026,N_325,N_19);
and U1027 (N_1027,N_159,N_189);
xnor U1028 (N_1028,N_241,N_244);
and U1029 (N_1029,N_479,N_470);
nand U1030 (N_1030,N_532,N_234);
or U1031 (N_1031,N_210,N_551);
or U1032 (N_1032,N_499,N_102);
nor U1033 (N_1033,N_106,N_188);
nor U1034 (N_1034,N_205,N_138);
or U1035 (N_1035,N_241,N_411);
nand U1036 (N_1036,N_111,N_54);
and U1037 (N_1037,N_270,N_274);
and U1038 (N_1038,N_358,N_59);
nor U1039 (N_1039,N_323,N_229);
nor U1040 (N_1040,N_214,N_593);
and U1041 (N_1041,N_9,N_58);
nand U1042 (N_1042,N_580,N_517);
xnor U1043 (N_1043,N_533,N_179);
nor U1044 (N_1044,N_265,N_21);
nor U1045 (N_1045,N_511,N_20);
and U1046 (N_1046,N_408,N_420);
or U1047 (N_1047,N_25,N_32);
nor U1048 (N_1048,N_481,N_499);
nor U1049 (N_1049,N_142,N_253);
or U1050 (N_1050,N_490,N_46);
or U1051 (N_1051,N_428,N_399);
or U1052 (N_1052,N_561,N_103);
or U1053 (N_1053,N_377,N_452);
or U1054 (N_1054,N_300,N_475);
nor U1055 (N_1055,N_167,N_165);
nor U1056 (N_1056,N_159,N_55);
nor U1057 (N_1057,N_147,N_461);
xor U1058 (N_1058,N_10,N_510);
or U1059 (N_1059,N_216,N_275);
or U1060 (N_1060,N_430,N_66);
nor U1061 (N_1061,N_151,N_197);
and U1062 (N_1062,N_87,N_291);
or U1063 (N_1063,N_389,N_256);
nor U1064 (N_1064,N_549,N_492);
nor U1065 (N_1065,N_424,N_542);
and U1066 (N_1066,N_324,N_555);
nor U1067 (N_1067,N_135,N_548);
or U1068 (N_1068,N_19,N_6);
nand U1069 (N_1069,N_70,N_103);
nor U1070 (N_1070,N_504,N_160);
nand U1071 (N_1071,N_520,N_154);
and U1072 (N_1072,N_573,N_416);
nand U1073 (N_1073,N_135,N_358);
and U1074 (N_1074,N_73,N_1);
and U1075 (N_1075,N_381,N_533);
nand U1076 (N_1076,N_536,N_450);
nor U1077 (N_1077,N_327,N_210);
nand U1078 (N_1078,N_362,N_201);
and U1079 (N_1079,N_271,N_546);
nor U1080 (N_1080,N_28,N_313);
or U1081 (N_1081,N_311,N_275);
and U1082 (N_1082,N_231,N_499);
or U1083 (N_1083,N_79,N_513);
and U1084 (N_1084,N_63,N_313);
nand U1085 (N_1085,N_162,N_172);
nand U1086 (N_1086,N_8,N_388);
and U1087 (N_1087,N_540,N_507);
or U1088 (N_1088,N_29,N_118);
and U1089 (N_1089,N_344,N_508);
nand U1090 (N_1090,N_0,N_588);
nor U1091 (N_1091,N_49,N_88);
and U1092 (N_1092,N_410,N_455);
nand U1093 (N_1093,N_88,N_556);
and U1094 (N_1094,N_36,N_43);
and U1095 (N_1095,N_243,N_282);
and U1096 (N_1096,N_255,N_453);
or U1097 (N_1097,N_321,N_409);
and U1098 (N_1098,N_2,N_284);
nand U1099 (N_1099,N_345,N_414);
nor U1100 (N_1100,N_395,N_191);
nor U1101 (N_1101,N_361,N_81);
nand U1102 (N_1102,N_250,N_257);
nor U1103 (N_1103,N_144,N_476);
and U1104 (N_1104,N_302,N_361);
or U1105 (N_1105,N_485,N_231);
nor U1106 (N_1106,N_26,N_19);
and U1107 (N_1107,N_99,N_243);
nor U1108 (N_1108,N_416,N_231);
or U1109 (N_1109,N_376,N_597);
and U1110 (N_1110,N_369,N_561);
nand U1111 (N_1111,N_212,N_409);
nand U1112 (N_1112,N_455,N_131);
nand U1113 (N_1113,N_585,N_23);
nand U1114 (N_1114,N_322,N_60);
nor U1115 (N_1115,N_244,N_19);
and U1116 (N_1116,N_466,N_7);
or U1117 (N_1117,N_254,N_338);
nor U1118 (N_1118,N_336,N_478);
and U1119 (N_1119,N_98,N_419);
and U1120 (N_1120,N_171,N_598);
and U1121 (N_1121,N_175,N_580);
and U1122 (N_1122,N_67,N_294);
and U1123 (N_1123,N_424,N_484);
nor U1124 (N_1124,N_373,N_146);
nor U1125 (N_1125,N_527,N_463);
and U1126 (N_1126,N_343,N_134);
and U1127 (N_1127,N_112,N_481);
and U1128 (N_1128,N_401,N_384);
and U1129 (N_1129,N_216,N_194);
nand U1130 (N_1130,N_105,N_405);
nand U1131 (N_1131,N_397,N_434);
or U1132 (N_1132,N_64,N_68);
nor U1133 (N_1133,N_430,N_406);
or U1134 (N_1134,N_329,N_326);
or U1135 (N_1135,N_71,N_110);
or U1136 (N_1136,N_108,N_253);
nand U1137 (N_1137,N_186,N_201);
nor U1138 (N_1138,N_508,N_390);
nor U1139 (N_1139,N_21,N_212);
nand U1140 (N_1140,N_553,N_29);
nand U1141 (N_1141,N_550,N_125);
or U1142 (N_1142,N_155,N_4);
and U1143 (N_1143,N_468,N_368);
and U1144 (N_1144,N_435,N_344);
nor U1145 (N_1145,N_399,N_390);
and U1146 (N_1146,N_84,N_95);
or U1147 (N_1147,N_279,N_129);
and U1148 (N_1148,N_79,N_303);
nor U1149 (N_1149,N_443,N_8);
nor U1150 (N_1150,N_450,N_111);
or U1151 (N_1151,N_489,N_531);
or U1152 (N_1152,N_550,N_587);
nor U1153 (N_1153,N_257,N_524);
or U1154 (N_1154,N_95,N_488);
xnor U1155 (N_1155,N_385,N_590);
nor U1156 (N_1156,N_305,N_303);
and U1157 (N_1157,N_161,N_326);
nor U1158 (N_1158,N_11,N_137);
nor U1159 (N_1159,N_382,N_97);
nand U1160 (N_1160,N_369,N_509);
or U1161 (N_1161,N_451,N_397);
nand U1162 (N_1162,N_223,N_566);
and U1163 (N_1163,N_456,N_130);
nor U1164 (N_1164,N_461,N_134);
or U1165 (N_1165,N_234,N_589);
or U1166 (N_1166,N_98,N_137);
nand U1167 (N_1167,N_466,N_381);
and U1168 (N_1168,N_575,N_257);
or U1169 (N_1169,N_438,N_67);
nand U1170 (N_1170,N_375,N_434);
nor U1171 (N_1171,N_92,N_302);
nand U1172 (N_1172,N_548,N_505);
or U1173 (N_1173,N_423,N_19);
or U1174 (N_1174,N_561,N_22);
or U1175 (N_1175,N_382,N_221);
nand U1176 (N_1176,N_287,N_516);
nor U1177 (N_1177,N_83,N_513);
or U1178 (N_1178,N_118,N_345);
and U1179 (N_1179,N_236,N_470);
nand U1180 (N_1180,N_404,N_323);
and U1181 (N_1181,N_476,N_228);
nor U1182 (N_1182,N_33,N_131);
nand U1183 (N_1183,N_6,N_283);
nor U1184 (N_1184,N_429,N_170);
nor U1185 (N_1185,N_147,N_524);
and U1186 (N_1186,N_431,N_336);
and U1187 (N_1187,N_226,N_289);
nand U1188 (N_1188,N_322,N_93);
nor U1189 (N_1189,N_470,N_550);
nand U1190 (N_1190,N_397,N_30);
or U1191 (N_1191,N_153,N_203);
or U1192 (N_1192,N_58,N_105);
and U1193 (N_1193,N_543,N_401);
nor U1194 (N_1194,N_365,N_249);
nand U1195 (N_1195,N_487,N_135);
or U1196 (N_1196,N_0,N_209);
or U1197 (N_1197,N_368,N_463);
and U1198 (N_1198,N_465,N_435);
or U1199 (N_1199,N_210,N_354);
or U1200 (N_1200,N_936,N_1100);
and U1201 (N_1201,N_906,N_603);
and U1202 (N_1202,N_1195,N_646);
or U1203 (N_1203,N_1016,N_782);
and U1204 (N_1204,N_1183,N_992);
and U1205 (N_1205,N_602,N_799);
nor U1206 (N_1206,N_970,N_801);
nand U1207 (N_1207,N_1174,N_761);
nand U1208 (N_1208,N_697,N_737);
nor U1209 (N_1209,N_889,N_600);
nand U1210 (N_1210,N_978,N_932);
nor U1211 (N_1211,N_708,N_1182);
nor U1212 (N_1212,N_1076,N_1090);
xor U1213 (N_1213,N_712,N_900);
nand U1214 (N_1214,N_1055,N_996);
or U1215 (N_1215,N_776,N_676);
nor U1216 (N_1216,N_771,N_633);
and U1217 (N_1217,N_947,N_909);
nand U1218 (N_1218,N_791,N_722);
nor U1219 (N_1219,N_1026,N_952);
nand U1220 (N_1220,N_832,N_640);
nor U1221 (N_1221,N_988,N_756);
nor U1222 (N_1222,N_916,N_1192);
nor U1223 (N_1223,N_891,N_1010);
and U1224 (N_1224,N_652,N_1101);
nand U1225 (N_1225,N_768,N_882);
nand U1226 (N_1226,N_885,N_1021);
or U1227 (N_1227,N_1000,N_655);
nand U1228 (N_1228,N_977,N_1027);
nor U1229 (N_1229,N_699,N_620);
nor U1230 (N_1230,N_1070,N_839);
nand U1231 (N_1231,N_1075,N_798);
or U1232 (N_1232,N_993,N_738);
or U1233 (N_1233,N_815,N_675);
nand U1234 (N_1234,N_758,N_661);
nand U1235 (N_1235,N_1030,N_783);
and U1236 (N_1236,N_868,N_824);
nand U1237 (N_1237,N_905,N_964);
and U1238 (N_1238,N_1050,N_904);
and U1239 (N_1239,N_1022,N_1179);
or U1240 (N_1240,N_1103,N_984);
and U1241 (N_1241,N_747,N_678);
and U1242 (N_1242,N_1163,N_662);
nor U1243 (N_1243,N_1032,N_898);
nor U1244 (N_1244,N_1116,N_751);
or U1245 (N_1245,N_744,N_1173);
nor U1246 (N_1246,N_704,N_615);
xor U1247 (N_1247,N_674,N_670);
and U1248 (N_1248,N_908,N_1064);
nand U1249 (N_1249,N_755,N_667);
or U1250 (N_1250,N_834,N_1108);
or U1251 (N_1251,N_1142,N_718);
nand U1252 (N_1252,N_1132,N_870);
and U1253 (N_1253,N_1031,N_843);
and U1254 (N_1254,N_1171,N_682);
nand U1255 (N_1255,N_881,N_770);
nand U1256 (N_1256,N_660,N_1036);
or U1257 (N_1257,N_767,N_1034);
nor U1258 (N_1258,N_1164,N_703);
and U1259 (N_1259,N_1001,N_1196);
or U1260 (N_1260,N_796,N_1046);
nand U1261 (N_1261,N_1194,N_1045);
nand U1262 (N_1262,N_622,N_884);
or U1263 (N_1263,N_1069,N_866);
xor U1264 (N_1264,N_1198,N_810);
nor U1265 (N_1265,N_873,N_800);
xnor U1266 (N_1266,N_1009,N_855);
or U1267 (N_1267,N_806,N_1135);
nor U1268 (N_1268,N_899,N_949);
nor U1269 (N_1269,N_642,N_886);
or U1270 (N_1270,N_903,N_943);
and U1271 (N_1271,N_1176,N_663);
nand U1272 (N_1272,N_1148,N_883);
nor U1273 (N_1273,N_1123,N_1134);
nor U1274 (N_1274,N_981,N_897);
nand U1275 (N_1275,N_894,N_994);
and U1276 (N_1276,N_705,N_725);
or U1277 (N_1277,N_926,N_1098);
nand U1278 (N_1278,N_957,N_789);
and U1279 (N_1279,N_1039,N_878);
nand U1280 (N_1280,N_630,N_690);
xnor U1281 (N_1281,N_757,N_1087);
nor U1282 (N_1282,N_962,N_609);
nand U1283 (N_1283,N_653,N_982);
nand U1284 (N_1284,N_1131,N_1102);
nand U1285 (N_1285,N_769,N_794);
nor U1286 (N_1286,N_845,N_1035);
and U1287 (N_1287,N_658,N_743);
nand U1288 (N_1288,N_1104,N_811);
and U1289 (N_1289,N_740,N_920);
nor U1290 (N_1290,N_1175,N_792);
and U1291 (N_1291,N_1130,N_1188);
and U1292 (N_1292,N_1165,N_732);
nor U1293 (N_1293,N_1144,N_805);
nand U1294 (N_1294,N_1153,N_1199);
nor U1295 (N_1295,N_1154,N_635);
or U1296 (N_1296,N_1184,N_989);
nor U1297 (N_1297,N_605,N_752);
or U1298 (N_1298,N_765,N_1178);
and U1299 (N_1299,N_679,N_973);
nand U1300 (N_1300,N_611,N_668);
nor U1301 (N_1301,N_736,N_1141);
and U1302 (N_1302,N_1172,N_692);
nor U1303 (N_1303,N_945,N_863);
nand U1304 (N_1304,N_976,N_1110);
xnor U1305 (N_1305,N_1043,N_601);
or U1306 (N_1306,N_681,N_944);
xor U1307 (N_1307,N_1189,N_913);
and U1308 (N_1308,N_968,N_731);
or U1309 (N_1309,N_876,N_1020);
xor U1310 (N_1310,N_733,N_840);
or U1311 (N_1311,N_745,N_1073);
xor U1312 (N_1312,N_616,N_1105);
and U1313 (N_1313,N_841,N_665);
or U1314 (N_1314,N_717,N_1119);
or U1315 (N_1315,N_750,N_707);
or U1316 (N_1316,N_1003,N_803);
or U1317 (N_1317,N_1006,N_1125);
nand U1318 (N_1318,N_948,N_809);
and U1319 (N_1319,N_639,N_659);
nand U1320 (N_1320,N_934,N_1107);
and U1321 (N_1321,N_685,N_930);
and U1322 (N_1322,N_688,N_941);
and U1323 (N_1323,N_1155,N_1028);
nand U1324 (N_1324,N_995,N_632);
and U1325 (N_1325,N_623,N_730);
nor U1326 (N_1326,N_1139,N_787);
nor U1327 (N_1327,N_1150,N_649);
xnor U1328 (N_1328,N_713,N_1080);
nor U1329 (N_1329,N_619,N_951);
and U1330 (N_1330,N_1088,N_825);
or U1331 (N_1331,N_1044,N_813);
nor U1332 (N_1332,N_818,N_1067);
and U1333 (N_1333,N_1061,N_777);
and U1334 (N_1334,N_1057,N_1099);
nand U1335 (N_1335,N_1047,N_775);
nor U1336 (N_1336,N_902,N_860);
and U1337 (N_1337,N_935,N_1082);
and U1338 (N_1338,N_650,N_946);
and U1339 (N_1339,N_647,N_654);
nand U1340 (N_1340,N_759,N_966);
or U1341 (N_1341,N_861,N_929);
nor U1342 (N_1342,N_1112,N_1012);
or U1343 (N_1343,N_854,N_910);
or U1344 (N_1344,N_680,N_980);
nand U1345 (N_1345,N_624,N_762);
nor U1346 (N_1346,N_1096,N_1152);
or U1347 (N_1347,N_786,N_1126);
and U1348 (N_1348,N_1072,N_735);
or U1349 (N_1349,N_698,N_1011);
nand U1350 (N_1350,N_1180,N_638);
or U1351 (N_1351,N_967,N_802);
nand U1352 (N_1352,N_833,N_1078);
or U1353 (N_1353,N_911,N_748);
and U1354 (N_1354,N_626,N_835);
and U1355 (N_1355,N_636,N_1138);
or U1356 (N_1356,N_779,N_817);
or U1357 (N_1357,N_629,N_634);
or U1358 (N_1358,N_875,N_846);
nand U1359 (N_1359,N_925,N_795);
nor U1360 (N_1360,N_1086,N_890);
or U1361 (N_1361,N_742,N_956);
nand U1362 (N_1362,N_1186,N_1193);
nand U1363 (N_1363,N_656,N_1007);
nand U1364 (N_1364,N_971,N_871);
and U1365 (N_1365,N_669,N_1106);
nor U1366 (N_1366,N_686,N_921);
or U1367 (N_1367,N_727,N_888);
or U1368 (N_1368,N_960,N_856);
and U1369 (N_1369,N_961,N_1002);
nand U1370 (N_1370,N_1143,N_726);
and U1371 (N_1371,N_772,N_612);
or U1372 (N_1372,N_1068,N_1084);
or U1373 (N_1373,N_784,N_694);
nand U1374 (N_1374,N_922,N_892);
nand U1375 (N_1375,N_1097,N_1118);
or U1376 (N_1376,N_1159,N_1127);
or U1377 (N_1377,N_901,N_1091);
or U1378 (N_1378,N_1053,N_729);
and U1379 (N_1379,N_604,N_711);
nor U1380 (N_1380,N_1197,N_672);
or U1381 (N_1381,N_1089,N_723);
or U1382 (N_1382,N_931,N_1017);
nor U1383 (N_1383,N_938,N_827);
nand U1384 (N_1384,N_780,N_1162);
nand U1385 (N_1385,N_621,N_1121);
nand U1386 (N_1386,N_618,N_1117);
nand U1387 (N_1387,N_928,N_702);
and U1388 (N_1388,N_1156,N_608);
or U1389 (N_1389,N_706,N_693);
or U1390 (N_1390,N_1093,N_1120);
nor U1391 (N_1391,N_797,N_847);
nor U1392 (N_1392,N_859,N_1052);
nor U1393 (N_1393,N_1074,N_979);
or U1394 (N_1394,N_969,N_822);
and U1395 (N_1395,N_1095,N_773);
and U1396 (N_1396,N_919,N_1040);
and U1397 (N_1397,N_657,N_923);
or U1398 (N_1398,N_651,N_983);
and U1399 (N_1399,N_1048,N_1013);
or U1400 (N_1400,N_1167,N_1015);
nand U1401 (N_1401,N_720,N_637);
nand U1402 (N_1402,N_1018,N_1124);
or U1403 (N_1403,N_1008,N_953);
and U1404 (N_1404,N_754,N_1071);
nand U1405 (N_1405,N_721,N_927);
and U1406 (N_1406,N_781,N_763);
nor U1407 (N_1407,N_1014,N_924);
and U1408 (N_1408,N_1114,N_857);
nor U1409 (N_1409,N_648,N_912);
or U1410 (N_1410,N_1170,N_987);
and U1411 (N_1411,N_1185,N_684);
and U1412 (N_1412,N_1160,N_741);
nor U1413 (N_1413,N_851,N_820);
and U1414 (N_1414,N_1133,N_790);
and U1415 (N_1415,N_1151,N_778);
nand U1416 (N_1416,N_848,N_997);
and U1417 (N_1417,N_1169,N_643);
and U1418 (N_1418,N_606,N_628);
and U1419 (N_1419,N_895,N_631);
and U1420 (N_1420,N_614,N_942);
or U1421 (N_1421,N_625,N_918);
or U1422 (N_1422,N_974,N_807);
nor U1423 (N_1423,N_965,N_1166);
nor U1424 (N_1424,N_1059,N_893);
nor U1425 (N_1425,N_724,N_950);
or U1426 (N_1426,N_1092,N_607);
or U1427 (N_1427,N_814,N_739);
or U1428 (N_1428,N_880,N_788);
nor U1429 (N_1429,N_879,N_641);
or U1430 (N_1430,N_937,N_1063);
nand U1431 (N_1431,N_998,N_1049);
and U1432 (N_1432,N_831,N_749);
and U1433 (N_1433,N_939,N_785);
xnor U1434 (N_1434,N_933,N_867);
or U1435 (N_1435,N_1122,N_1136);
or U1436 (N_1436,N_1129,N_842);
or U1437 (N_1437,N_990,N_849);
or U1438 (N_1438,N_677,N_714);
and U1439 (N_1439,N_746,N_700);
nand U1440 (N_1440,N_972,N_793);
and U1441 (N_1441,N_1023,N_1060);
or U1442 (N_1442,N_963,N_1094);
or U1443 (N_1443,N_838,N_1024);
and U1444 (N_1444,N_955,N_760);
or U1445 (N_1445,N_1177,N_940);
or U1446 (N_1446,N_954,N_695);
and U1447 (N_1447,N_1161,N_716);
and U1448 (N_1448,N_819,N_986);
and U1449 (N_1449,N_1038,N_715);
nand U1450 (N_1450,N_1042,N_1033);
or U1451 (N_1451,N_1187,N_613);
nand U1452 (N_1452,N_671,N_734);
or U1453 (N_1453,N_1058,N_1149);
nand U1454 (N_1454,N_877,N_1145);
or U1455 (N_1455,N_645,N_830);
nand U1456 (N_1456,N_959,N_1065);
nand U1457 (N_1457,N_673,N_975);
nand U1458 (N_1458,N_864,N_627);
or U1459 (N_1459,N_689,N_852);
and U1460 (N_1460,N_1191,N_1051);
or U1461 (N_1461,N_766,N_719);
or U1462 (N_1462,N_1109,N_1168);
and U1463 (N_1463,N_1111,N_1005);
nor U1464 (N_1464,N_829,N_1054);
nand U1465 (N_1465,N_753,N_823);
nand U1466 (N_1466,N_1137,N_808);
or U1467 (N_1467,N_844,N_644);
or U1468 (N_1468,N_1037,N_858);
and U1469 (N_1469,N_816,N_999);
xor U1470 (N_1470,N_812,N_764);
nand U1471 (N_1471,N_1146,N_687);
or U1472 (N_1472,N_837,N_991);
and U1473 (N_1473,N_1004,N_1062);
or U1474 (N_1474,N_610,N_1041);
and U1475 (N_1475,N_701,N_1083);
and U1476 (N_1476,N_710,N_683);
and U1477 (N_1477,N_1081,N_862);
nor U1478 (N_1478,N_666,N_1079);
nor U1479 (N_1479,N_664,N_896);
or U1480 (N_1480,N_836,N_958);
nand U1481 (N_1481,N_853,N_826);
nand U1482 (N_1482,N_1181,N_828);
and U1483 (N_1483,N_1157,N_850);
or U1484 (N_1484,N_874,N_617);
or U1485 (N_1485,N_869,N_1077);
or U1486 (N_1486,N_1085,N_917);
and U1487 (N_1487,N_1140,N_691);
and U1488 (N_1488,N_1190,N_1019);
or U1489 (N_1489,N_1029,N_872);
nor U1490 (N_1490,N_1025,N_865);
nand U1491 (N_1491,N_774,N_821);
and U1492 (N_1492,N_1115,N_1147);
nor U1493 (N_1493,N_1128,N_887);
nor U1494 (N_1494,N_1113,N_804);
and U1495 (N_1495,N_907,N_728);
nand U1496 (N_1496,N_1158,N_1056);
nor U1497 (N_1497,N_985,N_915);
and U1498 (N_1498,N_709,N_914);
and U1499 (N_1499,N_1066,N_696);
and U1500 (N_1500,N_1067,N_805);
and U1501 (N_1501,N_1155,N_997);
and U1502 (N_1502,N_857,N_836);
and U1503 (N_1503,N_1053,N_608);
nand U1504 (N_1504,N_731,N_646);
nand U1505 (N_1505,N_1113,N_740);
or U1506 (N_1506,N_988,N_1154);
nor U1507 (N_1507,N_1199,N_912);
xnor U1508 (N_1508,N_721,N_961);
nor U1509 (N_1509,N_1023,N_667);
or U1510 (N_1510,N_919,N_1090);
or U1511 (N_1511,N_737,N_927);
nand U1512 (N_1512,N_1078,N_1006);
nand U1513 (N_1513,N_1183,N_663);
nor U1514 (N_1514,N_1186,N_721);
nor U1515 (N_1515,N_1010,N_602);
nand U1516 (N_1516,N_915,N_878);
or U1517 (N_1517,N_896,N_883);
or U1518 (N_1518,N_811,N_1119);
nor U1519 (N_1519,N_822,N_967);
xnor U1520 (N_1520,N_656,N_607);
and U1521 (N_1521,N_668,N_1107);
nor U1522 (N_1522,N_674,N_1100);
and U1523 (N_1523,N_1004,N_928);
and U1524 (N_1524,N_1120,N_714);
nand U1525 (N_1525,N_854,N_747);
nand U1526 (N_1526,N_1010,N_1078);
or U1527 (N_1527,N_1189,N_1096);
or U1528 (N_1528,N_737,N_720);
or U1529 (N_1529,N_606,N_748);
and U1530 (N_1530,N_604,N_1144);
xor U1531 (N_1531,N_877,N_1051);
nor U1532 (N_1532,N_1158,N_617);
xor U1533 (N_1533,N_749,N_798);
or U1534 (N_1534,N_782,N_703);
nand U1535 (N_1535,N_638,N_971);
or U1536 (N_1536,N_874,N_799);
nor U1537 (N_1537,N_833,N_936);
nand U1538 (N_1538,N_871,N_906);
nor U1539 (N_1539,N_1022,N_653);
nor U1540 (N_1540,N_1182,N_1187);
or U1541 (N_1541,N_690,N_711);
nand U1542 (N_1542,N_896,N_889);
and U1543 (N_1543,N_868,N_1034);
nor U1544 (N_1544,N_771,N_622);
nor U1545 (N_1545,N_852,N_771);
nand U1546 (N_1546,N_895,N_874);
and U1547 (N_1547,N_1182,N_810);
or U1548 (N_1548,N_1196,N_1156);
nor U1549 (N_1549,N_773,N_643);
or U1550 (N_1550,N_1131,N_824);
and U1551 (N_1551,N_663,N_1008);
or U1552 (N_1552,N_1160,N_1151);
or U1553 (N_1553,N_641,N_660);
nand U1554 (N_1554,N_988,N_1031);
nor U1555 (N_1555,N_616,N_1093);
nand U1556 (N_1556,N_739,N_663);
nand U1557 (N_1557,N_737,N_803);
nand U1558 (N_1558,N_1016,N_785);
nor U1559 (N_1559,N_1087,N_802);
nand U1560 (N_1560,N_857,N_1128);
nor U1561 (N_1561,N_703,N_747);
xnor U1562 (N_1562,N_626,N_1019);
or U1563 (N_1563,N_926,N_745);
and U1564 (N_1564,N_1194,N_762);
nor U1565 (N_1565,N_1083,N_1097);
or U1566 (N_1566,N_631,N_786);
and U1567 (N_1567,N_1108,N_931);
or U1568 (N_1568,N_677,N_1020);
nor U1569 (N_1569,N_1033,N_1032);
and U1570 (N_1570,N_1068,N_1066);
or U1571 (N_1571,N_1046,N_798);
and U1572 (N_1572,N_973,N_776);
or U1573 (N_1573,N_858,N_805);
or U1574 (N_1574,N_935,N_1023);
nor U1575 (N_1575,N_940,N_733);
nand U1576 (N_1576,N_881,N_627);
nor U1577 (N_1577,N_714,N_756);
nand U1578 (N_1578,N_946,N_1186);
nand U1579 (N_1579,N_1188,N_1108);
xnor U1580 (N_1580,N_642,N_758);
or U1581 (N_1581,N_1136,N_820);
and U1582 (N_1582,N_1107,N_647);
nor U1583 (N_1583,N_957,N_834);
nand U1584 (N_1584,N_739,N_698);
and U1585 (N_1585,N_919,N_839);
nor U1586 (N_1586,N_606,N_919);
or U1587 (N_1587,N_738,N_690);
or U1588 (N_1588,N_1161,N_675);
nand U1589 (N_1589,N_1090,N_760);
nor U1590 (N_1590,N_629,N_876);
or U1591 (N_1591,N_1098,N_989);
nor U1592 (N_1592,N_1127,N_636);
nand U1593 (N_1593,N_608,N_1101);
nor U1594 (N_1594,N_1117,N_997);
nand U1595 (N_1595,N_1093,N_1044);
nor U1596 (N_1596,N_795,N_840);
nand U1597 (N_1597,N_682,N_631);
xnor U1598 (N_1598,N_786,N_686);
nor U1599 (N_1599,N_1150,N_1186);
nor U1600 (N_1600,N_739,N_856);
and U1601 (N_1601,N_1003,N_1136);
and U1602 (N_1602,N_661,N_644);
or U1603 (N_1603,N_661,N_1065);
nand U1604 (N_1604,N_849,N_1080);
nor U1605 (N_1605,N_844,N_645);
or U1606 (N_1606,N_1161,N_801);
and U1607 (N_1607,N_618,N_943);
nand U1608 (N_1608,N_1139,N_903);
and U1609 (N_1609,N_656,N_925);
or U1610 (N_1610,N_713,N_705);
nor U1611 (N_1611,N_797,N_1142);
nor U1612 (N_1612,N_1136,N_819);
nand U1613 (N_1613,N_652,N_616);
nor U1614 (N_1614,N_1031,N_708);
nand U1615 (N_1615,N_1158,N_644);
or U1616 (N_1616,N_911,N_1061);
or U1617 (N_1617,N_873,N_657);
or U1618 (N_1618,N_771,N_1068);
nand U1619 (N_1619,N_987,N_1140);
and U1620 (N_1620,N_626,N_664);
or U1621 (N_1621,N_764,N_1144);
and U1622 (N_1622,N_983,N_915);
nor U1623 (N_1623,N_604,N_1054);
nand U1624 (N_1624,N_862,N_994);
nor U1625 (N_1625,N_805,N_704);
and U1626 (N_1626,N_1182,N_1006);
nand U1627 (N_1627,N_757,N_783);
or U1628 (N_1628,N_1084,N_974);
or U1629 (N_1629,N_1155,N_894);
nand U1630 (N_1630,N_963,N_718);
and U1631 (N_1631,N_1042,N_1152);
and U1632 (N_1632,N_817,N_898);
nor U1633 (N_1633,N_1029,N_846);
nand U1634 (N_1634,N_976,N_889);
and U1635 (N_1635,N_1072,N_788);
nor U1636 (N_1636,N_1053,N_1007);
nand U1637 (N_1637,N_1113,N_1044);
nand U1638 (N_1638,N_1084,N_1089);
and U1639 (N_1639,N_723,N_778);
or U1640 (N_1640,N_957,N_910);
nor U1641 (N_1641,N_1082,N_764);
nor U1642 (N_1642,N_1197,N_1096);
nor U1643 (N_1643,N_1012,N_829);
or U1644 (N_1644,N_788,N_1082);
nand U1645 (N_1645,N_937,N_698);
and U1646 (N_1646,N_897,N_919);
and U1647 (N_1647,N_1073,N_863);
xnor U1648 (N_1648,N_1007,N_813);
and U1649 (N_1649,N_977,N_996);
and U1650 (N_1650,N_1184,N_1139);
and U1651 (N_1651,N_613,N_717);
and U1652 (N_1652,N_603,N_778);
and U1653 (N_1653,N_788,N_925);
xnor U1654 (N_1654,N_705,N_803);
and U1655 (N_1655,N_772,N_729);
nand U1656 (N_1656,N_796,N_1006);
nor U1657 (N_1657,N_676,N_603);
nand U1658 (N_1658,N_727,N_1091);
xor U1659 (N_1659,N_1142,N_725);
or U1660 (N_1660,N_877,N_1170);
nor U1661 (N_1661,N_798,N_1131);
nand U1662 (N_1662,N_1030,N_786);
and U1663 (N_1663,N_1057,N_866);
or U1664 (N_1664,N_797,N_980);
nor U1665 (N_1665,N_920,N_971);
nor U1666 (N_1666,N_968,N_1107);
or U1667 (N_1667,N_1063,N_730);
nand U1668 (N_1668,N_744,N_800);
nor U1669 (N_1669,N_780,N_1085);
nor U1670 (N_1670,N_916,N_627);
nor U1671 (N_1671,N_728,N_736);
and U1672 (N_1672,N_610,N_1066);
xnor U1673 (N_1673,N_727,N_1109);
or U1674 (N_1674,N_821,N_883);
or U1675 (N_1675,N_1172,N_762);
or U1676 (N_1676,N_792,N_1077);
nand U1677 (N_1677,N_618,N_791);
or U1678 (N_1678,N_778,N_1067);
or U1679 (N_1679,N_991,N_630);
or U1680 (N_1680,N_932,N_683);
nor U1681 (N_1681,N_666,N_635);
nand U1682 (N_1682,N_785,N_786);
nor U1683 (N_1683,N_1134,N_1136);
nand U1684 (N_1684,N_1114,N_730);
nor U1685 (N_1685,N_613,N_747);
and U1686 (N_1686,N_681,N_1023);
nand U1687 (N_1687,N_680,N_778);
or U1688 (N_1688,N_637,N_651);
nor U1689 (N_1689,N_824,N_839);
xnor U1690 (N_1690,N_1021,N_752);
or U1691 (N_1691,N_760,N_951);
nand U1692 (N_1692,N_912,N_862);
or U1693 (N_1693,N_891,N_735);
nor U1694 (N_1694,N_866,N_1093);
and U1695 (N_1695,N_837,N_771);
nor U1696 (N_1696,N_1097,N_1019);
and U1697 (N_1697,N_885,N_940);
nand U1698 (N_1698,N_925,N_751);
nor U1699 (N_1699,N_921,N_809);
and U1700 (N_1700,N_650,N_694);
or U1701 (N_1701,N_642,N_1155);
or U1702 (N_1702,N_995,N_1151);
or U1703 (N_1703,N_744,N_717);
or U1704 (N_1704,N_808,N_1190);
xor U1705 (N_1705,N_784,N_1085);
and U1706 (N_1706,N_764,N_1198);
and U1707 (N_1707,N_1015,N_1090);
or U1708 (N_1708,N_787,N_732);
nor U1709 (N_1709,N_1080,N_957);
or U1710 (N_1710,N_1021,N_967);
and U1711 (N_1711,N_661,N_665);
nand U1712 (N_1712,N_1088,N_1174);
nor U1713 (N_1713,N_680,N_1063);
and U1714 (N_1714,N_649,N_1117);
nand U1715 (N_1715,N_1141,N_621);
nor U1716 (N_1716,N_1194,N_702);
nor U1717 (N_1717,N_789,N_1036);
nor U1718 (N_1718,N_886,N_654);
nor U1719 (N_1719,N_942,N_908);
and U1720 (N_1720,N_944,N_617);
nor U1721 (N_1721,N_967,N_863);
nor U1722 (N_1722,N_1093,N_1165);
nor U1723 (N_1723,N_1122,N_737);
nor U1724 (N_1724,N_1164,N_1121);
nor U1725 (N_1725,N_994,N_976);
nor U1726 (N_1726,N_1117,N_931);
nand U1727 (N_1727,N_834,N_1037);
nor U1728 (N_1728,N_902,N_636);
or U1729 (N_1729,N_700,N_1101);
or U1730 (N_1730,N_819,N_774);
nand U1731 (N_1731,N_1103,N_921);
nor U1732 (N_1732,N_916,N_855);
or U1733 (N_1733,N_996,N_876);
nand U1734 (N_1734,N_1016,N_728);
nor U1735 (N_1735,N_811,N_816);
or U1736 (N_1736,N_861,N_952);
nor U1737 (N_1737,N_1139,N_1109);
and U1738 (N_1738,N_941,N_610);
nor U1739 (N_1739,N_713,N_756);
and U1740 (N_1740,N_715,N_1118);
and U1741 (N_1741,N_970,N_1175);
or U1742 (N_1742,N_945,N_683);
nand U1743 (N_1743,N_800,N_827);
xnor U1744 (N_1744,N_822,N_1092);
or U1745 (N_1745,N_1101,N_924);
nand U1746 (N_1746,N_600,N_634);
nand U1747 (N_1747,N_970,N_1043);
nor U1748 (N_1748,N_818,N_1180);
nand U1749 (N_1749,N_740,N_1052);
and U1750 (N_1750,N_1094,N_804);
nor U1751 (N_1751,N_974,N_1177);
nand U1752 (N_1752,N_881,N_1012);
nor U1753 (N_1753,N_901,N_950);
nor U1754 (N_1754,N_1048,N_756);
nor U1755 (N_1755,N_822,N_1038);
nor U1756 (N_1756,N_891,N_656);
nor U1757 (N_1757,N_686,N_1197);
nand U1758 (N_1758,N_978,N_1056);
nand U1759 (N_1759,N_676,N_963);
and U1760 (N_1760,N_813,N_818);
or U1761 (N_1761,N_884,N_604);
nand U1762 (N_1762,N_1017,N_1115);
nor U1763 (N_1763,N_932,N_610);
nand U1764 (N_1764,N_931,N_1032);
or U1765 (N_1765,N_602,N_800);
or U1766 (N_1766,N_855,N_917);
nand U1767 (N_1767,N_697,N_790);
or U1768 (N_1768,N_738,N_900);
nand U1769 (N_1769,N_1046,N_1068);
nand U1770 (N_1770,N_683,N_1059);
nand U1771 (N_1771,N_1095,N_830);
nand U1772 (N_1772,N_623,N_774);
or U1773 (N_1773,N_888,N_621);
nand U1774 (N_1774,N_1124,N_1104);
or U1775 (N_1775,N_998,N_1081);
nand U1776 (N_1776,N_608,N_687);
nand U1777 (N_1777,N_699,N_638);
nor U1778 (N_1778,N_985,N_674);
and U1779 (N_1779,N_930,N_977);
and U1780 (N_1780,N_1075,N_802);
xor U1781 (N_1781,N_786,N_1015);
nand U1782 (N_1782,N_1071,N_1184);
and U1783 (N_1783,N_916,N_949);
nor U1784 (N_1784,N_632,N_1152);
and U1785 (N_1785,N_1025,N_1135);
nor U1786 (N_1786,N_1110,N_729);
nor U1787 (N_1787,N_693,N_983);
and U1788 (N_1788,N_822,N_790);
nor U1789 (N_1789,N_1074,N_1159);
and U1790 (N_1790,N_1157,N_936);
and U1791 (N_1791,N_610,N_980);
nand U1792 (N_1792,N_942,N_827);
and U1793 (N_1793,N_663,N_680);
and U1794 (N_1794,N_1089,N_897);
and U1795 (N_1795,N_782,N_812);
nor U1796 (N_1796,N_706,N_765);
nand U1797 (N_1797,N_695,N_994);
nand U1798 (N_1798,N_1168,N_1010);
and U1799 (N_1799,N_692,N_752);
nand U1800 (N_1800,N_1397,N_1770);
nor U1801 (N_1801,N_1422,N_1798);
and U1802 (N_1802,N_1539,N_1760);
nand U1803 (N_1803,N_1266,N_1726);
nor U1804 (N_1804,N_1558,N_1700);
and U1805 (N_1805,N_1547,N_1553);
nand U1806 (N_1806,N_1343,N_1781);
nor U1807 (N_1807,N_1716,N_1666);
nor U1808 (N_1808,N_1670,N_1404);
and U1809 (N_1809,N_1660,N_1645);
or U1810 (N_1810,N_1505,N_1483);
or U1811 (N_1811,N_1329,N_1571);
or U1812 (N_1812,N_1545,N_1290);
or U1813 (N_1813,N_1515,N_1574);
nand U1814 (N_1814,N_1210,N_1302);
or U1815 (N_1815,N_1467,N_1363);
or U1816 (N_1816,N_1465,N_1695);
and U1817 (N_1817,N_1650,N_1447);
nand U1818 (N_1818,N_1618,N_1629);
or U1819 (N_1819,N_1484,N_1261);
or U1820 (N_1820,N_1573,N_1622);
nor U1821 (N_1821,N_1487,N_1643);
and U1822 (N_1822,N_1354,N_1698);
nand U1823 (N_1823,N_1448,N_1240);
nand U1824 (N_1824,N_1632,N_1534);
nor U1825 (N_1825,N_1427,N_1358);
nand U1826 (N_1826,N_1682,N_1379);
or U1827 (N_1827,N_1294,N_1353);
and U1828 (N_1828,N_1771,N_1405);
nand U1829 (N_1829,N_1456,N_1491);
or U1830 (N_1830,N_1316,N_1480);
nand U1831 (N_1831,N_1348,N_1355);
nor U1832 (N_1832,N_1678,N_1287);
or U1833 (N_1833,N_1518,N_1351);
nor U1834 (N_1834,N_1417,N_1498);
nand U1835 (N_1835,N_1520,N_1267);
and U1836 (N_1836,N_1318,N_1502);
nand U1837 (N_1837,N_1367,N_1658);
and U1838 (N_1838,N_1299,N_1663);
and U1839 (N_1839,N_1739,N_1537);
nand U1840 (N_1840,N_1708,N_1309);
nor U1841 (N_1841,N_1228,N_1747);
nand U1842 (N_1842,N_1426,N_1400);
nor U1843 (N_1843,N_1461,N_1260);
nor U1844 (N_1844,N_1754,N_1550);
or U1845 (N_1845,N_1703,N_1369);
nor U1846 (N_1846,N_1300,N_1415);
or U1847 (N_1847,N_1576,N_1514);
or U1848 (N_1848,N_1625,N_1671);
and U1849 (N_1849,N_1375,N_1635);
nand U1850 (N_1850,N_1603,N_1773);
and U1851 (N_1851,N_1508,N_1540);
nor U1852 (N_1852,N_1307,N_1684);
or U1853 (N_1853,N_1614,N_1373);
nor U1854 (N_1854,N_1292,N_1735);
nand U1855 (N_1855,N_1499,N_1697);
xnor U1856 (N_1856,N_1651,N_1399);
nand U1857 (N_1857,N_1460,N_1445);
and U1858 (N_1858,N_1580,N_1243);
nor U1859 (N_1859,N_1203,N_1255);
and U1860 (N_1860,N_1497,N_1291);
and U1861 (N_1861,N_1257,N_1711);
or U1862 (N_1862,N_1564,N_1283);
or U1863 (N_1863,N_1420,N_1689);
or U1864 (N_1864,N_1278,N_1477);
nand U1865 (N_1865,N_1282,N_1259);
and U1866 (N_1866,N_1264,N_1271);
or U1867 (N_1867,N_1249,N_1724);
xnor U1868 (N_1868,N_1552,N_1423);
and U1869 (N_1869,N_1721,N_1297);
nand U1870 (N_1870,N_1601,N_1357);
nor U1871 (N_1871,N_1503,N_1738);
nand U1872 (N_1872,N_1234,N_1380);
and U1873 (N_1873,N_1659,N_1269);
nor U1874 (N_1874,N_1667,N_1389);
nand U1875 (N_1875,N_1285,N_1270);
nor U1876 (N_1876,N_1326,N_1216);
and U1877 (N_1877,N_1332,N_1599);
nor U1878 (N_1878,N_1330,N_1471);
and U1879 (N_1879,N_1317,N_1741);
nand U1880 (N_1880,N_1296,N_1687);
and U1881 (N_1881,N_1606,N_1313);
or U1882 (N_1882,N_1734,N_1541);
or U1883 (N_1883,N_1474,N_1769);
nand U1884 (N_1884,N_1247,N_1311);
nand U1885 (N_1885,N_1275,N_1672);
nand U1886 (N_1886,N_1429,N_1665);
nor U1887 (N_1887,N_1374,N_1376);
or U1888 (N_1888,N_1386,N_1489);
and U1889 (N_1889,N_1683,N_1458);
nor U1890 (N_1890,N_1623,N_1214);
nor U1891 (N_1891,N_1293,N_1594);
nand U1892 (N_1892,N_1680,N_1425);
or U1893 (N_1893,N_1649,N_1706);
xor U1894 (N_1894,N_1767,N_1281);
nor U1895 (N_1895,N_1496,N_1325);
or U1896 (N_1896,N_1277,N_1604);
nor U1897 (N_1897,N_1419,N_1349);
and U1898 (N_1898,N_1555,N_1786);
and U1899 (N_1899,N_1432,N_1339);
xor U1900 (N_1900,N_1361,N_1661);
or U1901 (N_1901,N_1251,N_1522);
nand U1902 (N_1902,N_1342,N_1410);
or U1903 (N_1903,N_1433,N_1794);
nor U1904 (N_1904,N_1200,N_1208);
nor U1905 (N_1905,N_1345,N_1506);
or U1906 (N_1906,N_1476,N_1755);
or U1907 (N_1907,N_1602,N_1364);
and U1908 (N_1908,N_1322,N_1372);
or U1909 (N_1909,N_1621,N_1414);
or U1910 (N_1910,N_1685,N_1679);
nand U1911 (N_1911,N_1637,N_1779);
xnor U1912 (N_1912,N_1615,N_1352);
nand U1913 (N_1913,N_1745,N_1761);
or U1914 (N_1914,N_1593,N_1305);
and U1915 (N_1915,N_1793,N_1220);
nor U1916 (N_1916,N_1308,N_1718);
or U1917 (N_1917,N_1455,N_1273);
nand U1918 (N_1918,N_1385,N_1715);
or U1919 (N_1919,N_1640,N_1705);
or U1920 (N_1920,N_1336,N_1219);
and U1921 (N_1921,N_1639,N_1790);
and U1922 (N_1922,N_1562,N_1335);
and U1923 (N_1923,N_1230,N_1608);
or U1924 (N_1924,N_1535,N_1301);
and U1925 (N_1925,N_1206,N_1624);
and U1926 (N_1926,N_1519,N_1548);
nor U1927 (N_1927,N_1704,N_1398);
nor U1928 (N_1928,N_1304,N_1766);
nor U1929 (N_1929,N_1331,N_1396);
nor U1930 (N_1930,N_1482,N_1713);
and U1931 (N_1931,N_1529,N_1543);
and U1932 (N_1932,N_1512,N_1213);
nor U1933 (N_1933,N_1556,N_1551);
or U1934 (N_1934,N_1407,N_1241);
nand U1935 (N_1935,N_1488,N_1383);
nand U1936 (N_1936,N_1204,N_1239);
nor U1937 (N_1937,N_1648,N_1218);
and U1938 (N_1938,N_1561,N_1626);
nand U1939 (N_1939,N_1590,N_1674);
and U1940 (N_1940,N_1238,N_1406);
or U1941 (N_1941,N_1589,N_1584);
nor U1942 (N_1942,N_1653,N_1746);
and U1943 (N_1943,N_1436,N_1408);
nor U1944 (N_1944,N_1725,N_1748);
nor U1945 (N_1945,N_1466,N_1306);
nand U1946 (N_1946,N_1559,N_1457);
nor U1947 (N_1947,N_1394,N_1450);
or U1948 (N_1948,N_1217,N_1475);
or U1949 (N_1949,N_1530,N_1759);
or U1950 (N_1950,N_1628,N_1523);
or U1951 (N_1951,N_1310,N_1609);
nor U1952 (N_1952,N_1500,N_1231);
nor U1953 (N_1953,N_1638,N_1538);
or U1954 (N_1954,N_1526,N_1597);
nand U1955 (N_1955,N_1542,N_1350);
nor U1956 (N_1956,N_1586,N_1756);
nand U1957 (N_1957,N_1409,N_1472);
nand U1958 (N_1958,N_1333,N_1613);
xor U1959 (N_1959,N_1712,N_1578);
nor U1960 (N_1960,N_1315,N_1280);
or U1961 (N_1961,N_1510,N_1323);
nor U1962 (N_1962,N_1588,N_1531);
xor U1963 (N_1963,N_1642,N_1740);
or U1964 (N_1964,N_1356,N_1463);
nor U1965 (N_1965,N_1235,N_1710);
and U1966 (N_1966,N_1596,N_1494);
nand U1967 (N_1967,N_1565,N_1776);
xor U1968 (N_1968,N_1693,N_1513);
and U1969 (N_1969,N_1486,N_1692);
nor U1970 (N_1970,N_1749,N_1451);
or U1971 (N_1971,N_1733,N_1620);
nor U1972 (N_1972,N_1532,N_1647);
nor U1973 (N_1973,N_1441,N_1676);
and U1974 (N_1974,N_1401,N_1569);
nor U1975 (N_1975,N_1378,N_1709);
nor U1976 (N_1976,N_1464,N_1566);
nand U1977 (N_1977,N_1751,N_1320);
nand U1978 (N_1978,N_1485,N_1469);
nand U1979 (N_1979,N_1223,N_1493);
or U1980 (N_1980,N_1575,N_1567);
and U1981 (N_1981,N_1424,N_1262);
nor U1982 (N_1982,N_1656,N_1511);
and U1983 (N_1983,N_1341,N_1359);
and U1984 (N_1984,N_1382,N_1611);
nand U1985 (N_1985,N_1205,N_1517);
or U1986 (N_1986,N_1347,N_1371);
or U1987 (N_1987,N_1459,N_1254);
and U1988 (N_1988,N_1321,N_1797);
and U1989 (N_1989,N_1757,N_1224);
nand U1990 (N_1990,N_1612,N_1616);
nand U1991 (N_1991,N_1211,N_1582);
or U1992 (N_1992,N_1446,N_1274);
or U1993 (N_1993,N_1634,N_1473);
nand U1994 (N_1994,N_1595,N_1652);
nor U1995 (N_1995,N_1750,N_1438);
and U1996 (N_1996,N_1434,N_1744);
and U1997 (N_1997,N_1258,N_1758);
nand U1998 (N_1998,N_1403,N_1344);
or U1999 (N_1999,N_1365,N_1610);
nor U2000 (N_2000,N_1252,N_1752);
nand U2001 (N_2001,N_1334,N_1314);
nand U2002 (N_2002,N_1319,N_1490);
and U2003 (N_2003,N_1443,N_1557);
nand U2004 (N_2004,N_1242,N_1468);
and U2005 (N_2005,N_1362,N_1546);
xor U2006 (N_2006,N_1544,N_1720);
nor U2007 (N_2007,N_1699,N_1619);
or U2008 (N_2008,N_1250,N_1742);
nand U2009 (N_2009,N_1504,N_1799);
and U2010 (N_2010,N_1780,N_1675);
nor U2011 (N_2011,N_1743,N_1536);
and U2012 (N_2012,N_1337,N_1572);
nand U2013 (N_2013,N_1501,N_1694);
or U2014 (N_2014,N_1591,N_1783);
nor U2015 (N_2015,N_1636,N_1662);
nand U2016 (N_2016,N_1737,N_1585);
and U2017 (N_2017,N_1245,N_1600);
or U2018 (N_2018,N_1728,N_1253);
nor U2019 (N_2019,N_1527,N_1598);
nor U2020 (N_2020,N_1340,N_1392);
and U2021 (N_2021,N_1338,N_1212);
and U2022 (N_2022,N_1690,N_1444);
nand U2023 (N_2023,N_1732,N_1237);
nand U2024 (N_2024,N_1495,N_1644);
and U2025 (N_2025,N_1681,N_1554);
and U2026 (N_2026,N_1244,N_1246);
nand U2027 (N_2027,N_1366,N_1630);
nor U2028 (N_2028,N_1655,N_1528);
or U2029 (N_2029,N_1657,N_1226);
and U2030 (N_2030,N_1627,N_1201);
or U2031 (N_2031,N_1452,N_1525);
nor U2032 (N_2032,N_1722,N_1775);
and U2033 (N_2033,N_1763,N_1787);
and U2034 (N_2034,N_1507,N_1449);
or U2035 (N_2035,N_1388,N_1232);
nor U2036 (N_2036,N_1411,N_1723);
nor U2037 (N_2037,N_1222,N_1717);
nor U2038 (N_2038,N_1284,N_1286);
nand U2039 (N_2039,N_1288,N_1453);
nor U2040 (N_2040,N_1521,N_1577);
and U2041 (N_2041,N_1202,N_1646);
and U2042 (N_2042,N_1324,N_1289);
or U2043 (N_2043,N_1298,N_1265);
nand U2044 (N_2044,N_1207,N_1524);
nor U2045 (N_2045,N_1509,N_1607);
and U2046 (N_2046,N_1796,N_1479);
and U2047 (N_2047,N_1568,N_1753);
nand U2048 (N_2048,N_1765,N_1669);
and U2049 (N_2049,N_1516,N_1440);
nor U2050 (N_2050,N_1581,N_1360);
or U2051 (N_2051,N_1442,N_1256);
and U2052 (N_2052,N_1784,N_1328);
nor U2053 (N_2053,N_1549,N_1402);
and U2054 (N_2054,N_1416,N_1370);
nand U2055 (N_2055,N_1393,N_1470);
nor U2056 (N_2056,N_1719,N_1731);
nor U2057 (N_2057,N_1772,N_1686);
nor U2058 (N_2058,N_1563,N_1673);
nand U2059 (N_2059,N_1268,N_1688);
or U2060 (N_2060,N_1462,N_1791);
nor U2061 (N_2061,N_1789,N_1762);
nor U2062 (N_2062,N_1418,N_1579);
nor U2063 (N_2063,N_1327,N_1592);
nor U2064 (N_2064,N_1492,N_1439);
nand U2065 (N_2065,N_1714,N_1225);
and U2066 (N_2066,N_1390,N_1664);
nand U2067 (N_2067,N_1263,N_1785);
nand U2068 (N_2068,N_1533,N_1788);
or U2069 (N_2069,N_1413,N_1736);
and U2070 (N_2070,N_1387,N_1381);
or U2071 (N_2071,N_1428,N_1641);
nor U2072 (N_2072,N_1764,N_1215);
and U2073 (N_2073,N_1454,N_1227);
and U2074 (N_2074,N_1412,N_1587);
and U2075 (N_2075,N_1368,N_1696);
and U2076 (N_2076,N_1481,N_1229);
nor U2077 (N_2077,N_1276,N_1295);
and U2078 (N_2078,N_1209,N_1236);
nor U2079 (N_2079,N_1377,N_1570);
nand U2080 (N_2080,N_1437,N_1792);
or U2081 (N_2081,N_1768,N_1395);
or U2082 (N_2082,N_1312,N_1435);
and U2083 (N_2083,N_1478,N_1702);
or U2084 (N_2084,N_1617,N_1346);
and U2085 (N_2085,N_1248,N_1691);
nor U2086 (N_2086,N_1774,N_1430);
and U2087 (N_2087,N_1633,N_1701);
or U2088 (N_2088,N_1668,N_1654);
nor U2089 (N_2089,N_1421,N_1560);
or U2090 (N_2090,N_1605,N_1795);
nand U2091 (N_2091,N_1729,N_1631);
or U2092 (N_2092,N_1391,N_1677);
nand U2093 (N_2093,N_1730,N_1727);
or U2094 (N_2094,N_1583,N_1233);
nor U2095 (N_2095,N_1279,N_1778);
or U2096 (N_2096,N_1431,N_1384);
or U2097 (N_2097,N_1303,N_1782);
nand U2098 (N_2098,N_1221,N_1272);
and U2099 (N_2099,N_1707,N_1777);
nand U2100 (N_2100,N_1710,N_1232);
nand U2101 (N_2101,N_1547,N_1466);
or U2102 (N_2102,N_1612,N_1551);
nor U2103 (N_2103,N_1639,N_1268);
nand U2104 (N_2104,N_1579,N_1294);
and U2105 (N_2105,N_1606,N_1245);
and U2106 (N_2106,N_1479,N_1428);
nand U2107 (N_2107,N_1247,N_1558);
nor U2108 (N_2108,N_1614,N_1669);
or U2109 (N_2109,N_1354,N_1215);
and U2110 (N_2110,N_1689,N_1322);
xnor U2111 (N_2111,N_1579,N_1233);
and U2112 (N_2112,N_1771,N_1331);
nand U2113 (N_2113,N_1503,N_1473);
or U2114 (N_2114,N_1744,N_1221);
or U2115 (N_2115,N_1282,N_1680);
xnor U2116 (N_2116,N_1205,N_1274);
nor U2117 (N_2117,N_1720,N_1209);
or U2118 (N_2118,N_1621,N_1241);
nand U2119 (N_2119,N_1726,N_1444);
or U2120 (N_2120,N_1472,N_1439);
and U2121 (N_2121,N_1233,N_1456);
nand U2122 (N_2122,N_1253,N_1357);
or U2123 (N_2123,N_1692,N_1715);
and U2124 (N_2124,N_1600,N_1471);
and U2125 (N_2125,N_1672,N_1735);
nand U2126 (N_2126,N_1419,N_1354);
nand U2127 (N_2127,N_1705,N_1750);
nand U2128 (N_2128,N_1412,N_1440);
and U2129 (N_2129,N_1455,N_1301);
or U2130 (N_2130,N_1611,N_1645);
and U2131 (N_2131,N_1464,N_1696);
or U2132 (N_2132,N_1679,N_1373);
or U2133 (N_2133,N_1720,N_1348);
nor U2134 (N_2134,N_1338,N_1754);
and U2135 (N_2135,N_1773,N_1286);
or U2136 (N_2136,N_1389,N_1714);
or U2137 (N_2137,N_1487,N_1334);
and U2138 (N_2138,N_1778,N_1325);
nor U2139 (N_2139,N_1207,N_1756);
nand U2140 (N_2140,N_1620,N_1386);
or U2141 (N_2141,N_1451,N_1347);
or U2142 (N_2142,N_1362,N_1622);
and U2143 (N_2143,N_1748,N_1687);
nand U2144 (N_2144,N_1262,N_1227);
nand U2145 (N_2145,N_1260,N_1695);
and U2146 (N_2146,N_1307,N_1617);
and U2147 (N_2147,N_1666,N_1288);
or U2148 (N_2148,N_1396,N_1337);
nand U2149 (N_2149,N_1320,N_1459);
nor U2150 (N_2150,N_1339,N_1315);
nand U2151 (N_2151,N_1412,N_1503);
nor U2152 (N_2152,N_1300,N_1734);
nand U2153 (N_2153,N_1495,N_1655);
nor U2154 (N_2154,N_1201,N_1740);
nand U2155 (N_2155,N_1581,N_1784);
and U2156 (N_2156,N_1510,N_1280);
and U2157 (N_2157,N_1552,N_1360);
and U2158 (N_2158,N_1787,N_1513);
nand U2159 (N_2159,N_1627,N_1360);
nor U2160 (N_2160,N_1500,N_1301);
nor U2161 (N_2161,N_1572,N_1472);
nand U2162 (N_2162,N_1210,N_1490);
nand U2163 (N_2163,N_1734,N_1573);
or U2164 (N_2164,N_1663,N_1430);
or U2165 (N_2165,N_1409,N_1488);
nand U2166 (N_2166,N_1653,N_1499);
nand U2167 (N_2167,N_1643,N_1370);
or U2168 (N_2168,N_1759,N_1405);
or U2169 (N_2169,N_1421,N_1797);
or U2170 (N_2170,N_1644,N_1524);
and U2171 (N_2171,N_1527,N_1313);
and U2172 (N_2172,N_1744,N_1757);
and U2173 (N_2173,N_1343,N_1574);
and U2174 (N_2174,N_1302,N_1666);
and U2175 (N_2175,N_1352,N_1228);
nand U2176 (N_2176,N_1388,N_1667);
nor U2177 (N_2177,N_1668,N_1552);
and U2178 (N_2178,N_1352,N_1728);
and U2179 (N_2179,N_1313,N_1724);
or U2180 (N_2180,N_1734,N_1342);
nand U2181 (N_2181,N_1597,N_1443);
nor U2182 (N_2182,N_1327,N_1345);
nand U2183 (N_2183,N_1542,N_1698);
xor U2184 (N_2184,N_1443,N_1366);
nand U2185 (N_2185,N_1398,N_1443);
and U2186 (N_2186,N_1201,N_1454);
or U2187 (N_2187,N_1358,N_1219);
and U2188 (N_2188,N_1646,N_1343);
nand U2189 (N_2189,N_1748,N_1499);
nand U2190 (N_2190,N_1532,N_1334);
and U2191 (N_2191,N_1321,N_1759);
or U2192 (N_2192,N_1587,N_1670);
or U2193 (N_2193,N_1328,N_1764);
nand U2194 (N_2194,N_1422,N_1579);
and U2195 (N_2195,N_1673,N_1534);
nand U2196 (N_2196,N_1542,N_1745);
nor U2197 (N_2197,N_1443,N_1494);
or U2198 (N_2198,N_1639,N_1219);
xnor U2199 (N_2199,N_1644,N_1636);
nand U2200 (N_2200,N_1569,N_1403);
nor U2201 (N_2201,N_1280,N_1745);
and U2202 (N_2202,N_1400,N_1722);
nor U2203 (N_2203,N_1565,N_1223);
nand U2204 (N_2204,N_1534,N_1303);
and U2205 (N_2205,N_1312,N_1289);
xnor U2206 (N_2206,N_1444,N_1650);
nand U2207 (N_2207,N_1492,N_1229);
or U2208 (N_2208,N_1546,N_1502);
and U2209 (N_2209,N_1703,N_1661);
nor U2210 (N_2210,N_1596,N_1358);
or U2211 (N_2211,N_1734,N_1587);
xor U2212 (N_2212,N_1604,N_1306);
or U2213 (N_2213,N_1203,N_1607);
or U2214 (N_2214,N_1514,N_1602);
and U2215 (N_2215,N_1367,N_1449);
and U2216 (N_2216,N_1599,N_1543);
nand U2217 (N_2217,N_1555,N_1771);
or U2218 (N_2218,N_1519,N_1413);
or U2219 (N_2219,N_1240,N_1773);
nand U2220 (N_2220,N_1368,N_1301);
nand U2221 (N_2221,N_1327,N_1322);
nor U2222 (N_2222,N_1408,N_1792);
nand U2223 (N_2223,N_1583,N_1260);
nor U2224 (N_2224,N_1263,N_1253);
nand U2225 (N_2225,N_1541,N_1357);
and U2226 (N_2226,N_1607,N_1658);
or U2227 (N_2227,N_1341,N_1521);
nor U2228 (N_2228,N_1487,N_1213);
and U2229 (N_2229,N_1519,N_1398);
nand U2230 (N_2230,N_1500,N_1425);
nand U2231 (N_2231,N_1722,N_1547);
or U2232 (N_2232,N_1248,N_1383);
and U2233 (N_2233,N_1787,N_1764);
and U2234 (N_2234,N_1487,N_1457);
and U2235 (N_2235,N_1604,N_1430);
nand U2236 (N_2236,N_1261,N_1737);
and U2237 (N_2237,N_1661,N_1613);
nand U2238 (N_2238,N_1710,N_1280);
and U2239 (N_2239,N_1379,N_1658);
nor U2240 (N_2240,N_1274,N_1309);
nor U2241 (N_2241,N_1271,N_1411);
or U2242 (N_2242,N_1333,N_1747);
or U2243 (N_2243,N_1558,N_1691);
or U2244 (N_2244,N_1232,N_1497);
or U2245 (N_2245,N_1758,N_1272);
nand U2246 (N_2246,N_1303,N_1579);
nor U2247 (N_2247,N_1222,N_1688);
nand U2248 (N_2248,N_1250,N_1666);
nand U2249 (N_2249,N_1702,N_1226);
and U2250 (N_2250,N_1676,N_1691);
or U2251 (N_2251,N_1664,N_1753);
nand U2252 (N_2252,N_1629,N_1401);
and U2253 (N_2253,N_1325,N_1763);
nand U2254 (N_2254,N_1632,N_1541);
and U2255 (N_2255,N_1212,N_1303);
and U2256 (N_2256,N_1701,N_1462);
nor U2257 (N_2257,N_1308,N_1574);
nand U2258 (N_2258,N_1552,N_1458);
nand U2259 (N_2259,N_1707,N_1704);
and U2260 (N_2260,N_1471,N_1232);
and U2261 (N_2261,N_1216,N_1679);
nand U2262 (N_2262,N_1370,N_1606);
nor U2263 (N_2263,N_1741,N_1733);
and U2264 (N_2264,N_1464,N_1206);
and U2265 (N_2265,N_1572,N_1214);
nor U2266 (N_2266,N_1625,N_1699);
nand U2267 (N_2267,N_1570,N_1255);
and U2268 (N_2268,N_1294,N_1255);
and U2269 (N_2269,N_1696,N_1348);
nand U2270 (N_2270,N_1313,N_1427);
nor U2271 (N_2271,N_1314,N_1522);
nand U2272 (N_2272,N_1580,N_1583);
nand U2273 (N_2273,N_1619,N_1397);
and U2274 (N_2274,N_1498,N_1526);
or U2275 (N_2275,N_1683,N_1799);
nor U2276 (N_2276,N_1257,N_1275);
and U2277 (N_2277,N_1443,N_1635);
nand U2278 (N_2278,N_1706,N_1684);
and U2279 (N_2279,N_1294,N_1226);
nor U2280 (N_2280,N_1426,N_1781);
and U2281 (N_2281,N_1281,N_1237);
nor U2282 (N_2282,N_1531,N_1352);
nor U2283 (N_2283,N_1700,N_1267);
and U2284 (N_2284,N_1249,N_1564);
nor U2285 (N_2285,N_1331,N_1760);
nor U2286 (N_2286,N_1526,N_1310);
nand U2287 (N_2287,N_1454,N_1331);
nor U2288 (N_2288,N_1293,N_1552);
nand U2289 (N_2289,N_1479,N_1327);
nor U2290 (N_2290,N_1475,N_1248);
nor U2291 (N_2291,N_1486,N_1490);
or U2292 (N_2292,N_1772,N_1604);
nand U2293 (N_2293,N_1700,N_1796);
or U2294 (N_2294,N_1585,N_1268);
nor U2295 (N_2295,N_1559,N_1665);
or U2296 (N_2296,N_1707,N_1261);
nor U2297 (N_2297,N_1211,N_1678);
nand U2298 (N_2298,N_1679,N_1474);
or U2299 (N_2299,N_1219,N_1786);
or U2300 (N_2300,N_1479,N_1633);
nor U2301 (N_2301,N_1538,N_1328);
and U2302 (N_2302,N_1560,N_1673);
and U2303 (N_2303,N_1618,N_1649);
and U2304 (N_2304,N_1278,N_1425);
and U2305 (N_2305,N_1538,N_1473);
and U2306 (N_2306,N_1535,N_1608);
nor U2307 (N_2307,N_1262,N_1243);
and U2308 (N_2308,N_1372,N_1324);
or U2309 (N_2309,N_1210,N_1786);
nand U2310 (N_2310,N_1230,N_1601);
and U2311 (N_2311,N_1520,N_1613);
nor U2312 (N_2312,N_1211,N_1722);
or U2313 (N_2313,N_1480,N_1563);
nand U2314 (N_2314,N_1402,N_1525);
nor U2315 (N_2315,N_1436,N_1291);
nand U2316 (N_2316,N_1342,N_1641);
and U2317 (N_2317,N_1536,N_1399);
or U2318 (N_2318,N_1650,N_1389);
and U2319 (N_2319,N_1742,N_1416);
and U2320 (N_2320,N_1339,N_1441);
nand U2321 (N_2321,N_1326,N_1335);
nand U2322 (N_2322,N_1377,N_1411);
nand U2323 (N_2323,N_1468,N_1416);
or U2324 (N_2324,N_1213,N_1373);
nand U2325 (N_2325,N_1332,N_1286);
and U2326 (N_2326,N_1337,N_1320);
and U2327 (N_2327,N_1347,N_1780);
nor U2328 (N_2328,N_1412,N_1231);
nand U2329 (N_2329,N_1346,N_1724);
and U2330 (N_2330,N_1417,N_1723);
and U2331 (N_2331,N_1335,N_1448);
nand U2332 (N_2332,N_1543,N_1208);
or U2333 (N_2333,N_1745,N_1794);
nor U2334 (N_2334,N_1560,N_1644);
or U2335 (N_2335,N_1727,N_1655);
and U2336 (N_2336,N_1424,N_1465);
nand U2337 (N_2337,N_1380,N_1552);
nor U2338 (N_2338,N_1251,N_1315);
nor U2339 (N_2339,N_1456,N_1745);
nor U2340 (N_2340,N_1326,N_1428);
nor U2341 (N_2341,N_1330,N_1628);
or U2342 (N_2342,N_1603,N_1506);
and U2343 (N_2343,N_1752,N_1596);
or U2344 (N_2344,N_1453,N_1517);
or U2345 (N_2345,N_1715,N_1242);
nand U2346 (N_2346,N_1684,N_1686);
or U2347 (N_2347,N_1752,N_1254);
or U2348 (N_2348,N_1292,N_1514);
nand U2349 (N_2349,N_1436,N_1325);
nor U2350 (N_2350,N_1686,N_1703);
or U2351 (N_2351,N_1691,N_1665);
or U2352 (N_2352,N_1596,N_1794);
and U2353 (N_2353,N_1395,N_1689);
or U2354 (N_2354,N_1614,N_1477);
nor U2355 (N_2355,N_1594,N_1353);
and U2356 (N_2356,N_1241,N_1415);
nand U2357 (N_2357,N_1745,N_1277);
or U2358 (N_2358,N_1365,N_1230);
and U2359 (N_2359,N_1202,N_1647);
nor U2360 (N_2360,N_1751,N_1738);
xnor U2361 (N_2361,N_1616,N_1707);
nor U2362 (N_2362,N_1722,N_1589);
and U2363 (N_2363,N_1465,N_1257);
or U2364 (N_2364,N_1671,N_1561);
and U2365 (N_2365,N_1405,N_1249);
nand U2366 (N_2366,N_1538,N_1722);
nor U2367 (N_2367,N_1469,N_1466);
nor U2368 (N_2368,N_1673,N_1747);
or U2369 (N_2369,N_1387,N_1562);
nand U2370 (N_2370,N_1383,N_1793);
or U2371 (N_2371,N_1338,N_1782);
nand U2372 (N_2372,N_1537,N_1782);
or U2373 (N_2373,N_1224,N_1730);
nand U2374 (N_2374,N_1551,N_1779);
nand U2375 (N_2375,N_1614,N_1327);
nand U2376 (N_2376,N_1695,N_1449);
nor U2377 (N_2377,N_1249,N_1354);
nor U2378 (N_2378,N_1278,N_1420);
nand U2379 (N_2379,N_1684,N_1242);
xnor U2380 (N_2380,N_1221,N_1726);
or U2381 (N_2381,N_1398,N_1421);
or U2382 (N_2382,N_1660,N_1692);
nor U2383 (N_2383,N_1727,N_1420);
nor U2384 (N_2384,N_1240,N_1425);
and U2385 (N_2385,N_1415,N_1437);
or U2386 (N_2386,N_1668,N_1537);
or U2387 (N_2387,N_1776,N_1375);
nor U2388 (N_2388,N_1769,N_1391);
nor U2389 (N_2389,N_1230,N_1208);
nor U2390 (N_2390,N_1791,N_1588);
nor U2391 (N_2391,N_1576,N_1533);
or U2392 (N_2392,N_1450,N_1315);
nand U2393 (N_2393,N_1495,N_1731);
or U2394 (N_2394,N_1722,N_1671);
nor U2395 (N_2395,N_1382,N_1629);
nand U2396 (N_2396,N_1227,N_1516);
or U2397 (N_2397,N_1219,N_1338);
nand U2398 (N_2398,N_1426,N_1790);
or U2399 (N_2399,N_1551,N_1314);
or U2400 (N_2400,N_1969,N_2196);
or U2401 (N_2401,N_2323,N_1986);
or U2402 (N_2402,N_1822,N_2173);
nor U2403 (N_2403,N_2243,N_2129);
nor U2404 (N_2404,N_2127,N_2358);
and U2405 (N_2405,N_2334,N_2302);
or U2406 (N_2406,N_2044,N_2037);
nand U2407 (N_2407,N_1965,N_2264);
nand U2408 (N_2408,N_2342,N_2031);
nand U2409 (N_2409,N_2242,N_2078);
nor U2410 (N_2410,N_1935,N_1896);
nand U2411 (N_2411,N_1962,N_1800);
or U2412 (N_2412,N_2319,N_2343);
and U2413 (N_2413,N_2199,N_2133);
and U2414 (N_2414,N_1842,N_2113);
nand U2415 (N_2415,N_2318,N_2105);
nor U2416 (N_2416,N_1874,N_2390);
or U2417 (N_2417,N_2035,N_1967);
and U2418 (N_2418,N_1988,N_1817);
nor U2419 (N_2419,N_2398,N_2089);
and U2420 (N_2420,N_1899,N_2200);
or U2421 (N_2421,N_1903,N_1846);
or U2422 (N_2422,N_2259,N_1886);
or U2423 (N_2423,N_2189,N_2174);
xor U2424 (N_2424,N_2191,N_2224);
or U2425 (N_2425,N_2081,N_2206);
or U2426 (N_2426,N_2304,N_2294);
and U2427 (N_2427,N_2040,N_2145);
nor U2428 (N_2428,N_1914,N_2177);
or U2429 (N_2429,N_2024,N_2307);
nor U2430 (N_2430,N_2399,N_2141);
nand U2431 (N_2431,N_2114,N_1921);
or U2432 (N_2432,N_1824,N_2027);
nand U2433 (N_2433,N_1918,N_2159);
nor U2434 (N_2434,N_2063,N_1989);
nor U2435 (N_2435,N_2134,N_1825);
nand U2436 (N_2436,N_2384,N_2231);
or U2437 (N_2437,N_1995,N_1902);
nor U2438 (N_2438,N_1900,N_2085);
and U2439 (N_2439,N_2363,N_2303);
and U2440 (N_2440,N_2279,N_2204);
xor U2441 (N_2441,N_1898,N_2347);
and U2442 (N_2442,N_2023,N_2149);
nor U2443 (N_2443,N_2290,N_2077);
nor U2444 (N_2444,N_2253,N_1930);
nand U2445 (N_2445,N_2160,N_2122);
nor U2446 (N_2446,N_2360,N_1904);
or U2447 (N_2447,N_2104,N_2041);
or U2448 (N_2448,N_1907,N_2103);
or U2449 (N_2449,N_2060,N_1819);
and U2450 (N_2450,N_1980,N_1922);
nand U2451 (N_2451,N_2240,N_2192);
nor U2452 (N_2452,N_1805,N_2119);
or U2453 (N_2453,N_2282,N_1857);
or U2454 (N_2454,N_2088,N_2255);
nor U2455 (N_2455,N_2228,N_1939);
and U2456 (N_2456,N_2135,N_2272);
or U2457 (N_2457,N_1868,N_1936);
or U2458 (N_2458,N_1873,N_2115);
nor U2459 (N_2459,N_2066,N_1864);
nand U2460 (N_2460,N_2260,N_2324);
nand U2461 (N_2461,N_1820,N_1806);
or U2462 (N_2462,N_2297,N_2288);
or U2463 (N_2463,N_2393,N_1855);
nand U2464 (N_2464,N_2274,N_1870);
nor U2465 (N_2465,N_1883,N_1998);
nand U2466 (N_2466,N_1830,N_2169);
nor U2467 (N_2467,N_2366,N_2331);
xor U2468 (N_2468,N_2090,N_1976);
or U2469 (N_2469,N_1933,N_2335);
nand U2470 (N_2470,N_1837,N_2352);
or U2471 (N_2471,N_1829,N_2170);
and U2472 (N_2472,N_2202,N_2117);
and U2473 (N_2473,N_2179,N_2010);
xnor U2474 (N_2474,N_2018,N_1926);
nand U2475 (N_2475,N_2107,N_2396);
and U2476 (N_2476,N_2292,N_2190);
nor U2477 (N_2477,N_1890,N_1880);
and U2478 (N_2478,N_2147,N_1894);
nand U2479 (N_2479,N_2344,N_1836);
and U2480 (N_2480,N_2234,N_2161);
nor U2481 (N_2481,N_2152,N_2211);
nand U2482 (N_2482,N_1951,N_1821);
nand U2483 (N_2483,N_2167,N_1885);
or U2484 (N_2484,N_1938,N_1801);
or U2485 (N_2485,N_2101,N_2053);
nor U2486 (N_2486,N_2079,N_2021);
nor U2487 (N_2487,N_1952,N_1985);
and U2488 (N_2488,N_2182,N_2245);
nand U2489 (N_2489,N_1917,N_1959);
nand U2490 (N_2490,N_1839,N_2042);
or U2491 (N_2491,N_1966,N_2164);
nand U2492 (N_2492,N_1809,N_2359);
nand U2493 (N_2493,N_1960,N_1889);
or U2494 (N_2494,N_2267,N_1961);
and U2495 (N_2495,N_1975,N_1942);
nor U2496 (N_2496,N_2136,N_2386);
or U2497 (N_2497,N_1990,N_1957);
nand U2498 (N_2498,N_2373,N_2311);
xor U2499 (N_2499,N_2312,N_2100);
or U2500 (N_2500,N_2310,N_1972);
nor U2501 (N_2501,N_2193,N_2020);
nand U2502 (N_2502,N_1982,N_1901);
and U2503 (N_2503,N_1863,N_2009);
nor U2504 (N_2504,N_1915,N_2383);
or U2505 (N_2505,N_2388,N_1848);
nand U2506 (N_2506,N_1808,N_2356);
and U2507 (N_2507,N_2256,N_2295);
nand U2508 (N_2508,N_2087,N_2291);
or U2509 (N_2509,N_2249,N_2284);
nor U2510 (N_2510,N_2299,N_2368);
or U2511 (N_2511,N_2011,N_2171);
nand U2512 (N_2512,N_1861,N_1944);
or U2513 (N_2513,N_1844,N_2380);
nand U2514 (N_2514,N_2265,N_1826);
nand U2515 (N_2515,N_2203,N_2034);
and U2516 (N_2516,N_2013,N_1947);
nor U2517 (N_2517,N_2233,N_1828);
nor U2518 (N_2518,N_2301,N_2340);
xnor U2519 (N_2519,N_1879,N_1888);
nor U2520 (N_2520,N_2032,N_1812);
nand U2521 (N_2521,N_1875,N_2188);
or U2522 (N_2522,N_1994,N_1992);
xor U2523 (N_2523,N_2139,N_2391);
or U2524 (N_2524,N_1814,N_1971);
nand U2525 (N_2525,N_2002,N_1866);
and U2526 (N_2526,N_1831,N_2225);
nand U2527 (N_2527,N_1973,N_1813);
or U2528 (N_2528,N_2055,N_2350);
nor U2529 (N_2529,N_2073,N_1862);
or U2530 (N_2530,N_1802,N_2165);
or U2531 (N_2531,N_1923,N_2070);
and U2532 (N_2532,N_1934,N_2019);
or U2533 (N_2533,N_2154,N_1878);
nand U2534 (N_2534,N_1849,N_2280);
or U2535 (N_2535,N_1832,N_2287);
xor U2536 (N_2536,N_2195,N_2395);
nand U2537 (N_2537,N_1943,N_2314);
nand U2538 (N_2538,N_2376,N_2345);
nand U2539 (N_2539,N_1996,N_2208);
and U2540 (N_2540,N_2254,N_2125);
and U2541 (N_2541,N_2364,N_1893);
and U2542 (N_2542,N_2030,N_2250);
and U2543 (N_2543,N_2246,N_2095);
nor U2544 (N_2544,N_2248,N_1940);
and U2545 (N_2545,N_1948,N_2099);
or U2546 (N_2546,N_2207,N_2048);
and U2547 (N_2547,N_2194,N_2258);
nand U2548 (N_2548,N_2014,N_2144);
nand U2549 (N_2549,N_1835,N_1911);
nand U2550 (N_2550,N_2049,N_2330);
or U2551 (N_2551,N_1924,N_2283);
or U2552 (N_2552,N_2385,N_2325);
nor U2553 (N_2553,N_2198,N_2074);
nor U2554 (N_2554,N_1997,N_2351);
or U2555 (N_2555,N_1981,N_1946);
xnor U2556 (N_2556,N_2241,N_1860);
or U2557 (N_2557,N_2271,N_2375);
and U2558 (N_2558,N_2273,N_2362);
or U2559 (N_2559,N_1810,N_2006);
nand U2560 (N_2560,N_2069,N_1823);
and U2561 (N_2561,N_2214,N_2217);
and U2562 (N_2562,N_2051,N_2332);
nand U2563 (N_2563,N_2232,N_2112);
nor U2564 (N_2564,N_2337,N_2238);
and U2565 (N_2565,N_2308,N_2205);
and U2566 (N_2566,N_2150,N_1937);
or U2567 (N_2567,N_2372,N_2381);
and U2568 (N_2568,N_2336,N_2065);
nor U2569 (N_2569,N_1963,N_2361);
or U2570 (N_2570,N_1983,N_2237);
and U2571 (N_2571,N_2007,N_2353);
and U2572 (N_2572,N_2275,N_2175);
nand U2573 (N_2573,N_1818,N_2235);
or U2574 (N_2574,N_1887,N_1927);
nand U2575 (N_2575,N_1931,N_2339);
or U2576 (N_2576,N_2181,N_2052);
and U2577 (N_2577,N_2116,N_2118);
or U2578 (N_2578,N_2168,N_2015);
and U2579 (N_2579,N_2091,N_2028);
or U2580 (N_2580,N_1859,N_2215);
or U2581 (N_2581,N_1984,N_2183);
xnor U2582 (N_2582,N_1858,N_2220);
and U2583 (N_2583,N_2397,N_2096);
or U2584 (N_2584,N_1932,N_2016);
or U2585 (N_2585,N_2132,N_1925);
or U2586 (N_2586,N_2148,N_2140);
or U2587 (N_2587,N_2157,N_1847);
nor U2588 (N_2588,N_1803,N_2050);
and U2589 (N_2589,N_1977,N_2263);
or U2590 (N_2590,N_1991,N_2075);
xor U2591 (N_2591,N_2138,N_1851);
nand U2592 (N_2592,N_2338,N_1958);
nor U2593 (N_2593,N_1891,N_2045);
nand U2594 (N_2594,N_2370,N_2309);
and U2595 (N_2595,N_2185,N_1941);
xnor U2596 (N_2596,N_1852,N_2076);
or U2597 (N_2597,N_2084,N_2367);
nand U2598 (N_2598,N_1811,N_2278);
and U2599 (N_2599,N_2223,N_2180);
nor U2600 (N_2600,N_2389,N_1970);
nand U2601 (N_2601,N_1838,N_1905);
and U2602 (N_2602,N_1850,N_2313);
nor U2603 (N_2603,N_2382,N_2124);
nor U2604 (N_2604,N_2093,N_2355);
and U2605 (N_2605,N_2329,N_1871);
nand U2606 (N_2606,N_2058,N_1913);
nand U2607 (N_2607,N_1954,N_2276);
and U2608 (N_2608,N_2008,N_2285);
xor U2609 (N_2609,N_2328,N_2394);
or U2610 (N_2610,N_2251,N_2266);
and U2611 (N_2611,N_2158,N_2155);
nand U2612 (N_2612,N_1949,N_2247);
nand U2613 (N_2613,N_2082,N_2106);
nor U2614 (N_2614,N_2239,N_2109);
and U2615 (N_2615,N_2341,N_1816);
or U2616 (N_2616,N_2377,N_2004);
or U2617 (N_2617,N_2346,N_2333);
nand U2618 (N_2618,N_1950,N_1945);
nand U2619 (N_2619,N_2320,N_2257);
nand U2620 (N_2620,N_2162,N_2221);
or U2621 (N_2621,N_2316,N_2230);
nor U2622 (N_2622,N_2186,N_2387);
or U2623 (N_2623,N_2327,N_2046);
nor U2624 (N_2624,N_1897,N_2210);
and U2625 (N_2625,N_1841,N_2003);
and U2626 (N_2626,N_2296,N_1993);
xor U2627 (N_2627,N_2317,N_2005);
nand U2628 (N_2628,N_1929,N_2163);
or U2629 (N_2629,N_2094,N_2268);
or U2630 (N_2630,N_2137,N_2038);
or U2631 (N_2631,N_2068,N_2121);
and U2632 (N_2632,N_1978,N_2128);
or U2633 (N_2633,N_1906,N_2348);
nand U2634 (N_2634,N_2000,N_2123);
and U2635 (N_2635,N_2143,N_2057);
nor U2636 (N_2636,N_2354,N_2286);
or U2637 (N_2637,N_2305,N_2083);
nor U2638 (N_2638,N_2212,N_2166);
and U2639 (N_2639,N_2054,N_2244);
nand U2640 (N_2640,N_2097,N_2120);
or U2641 (N_2641,N_2126,N_2374);
nand U2642 (N_2642,N_2306,N_1840);
nand U2643 (N_2643,N_2064,N_2321);
nor U2644 (N_2644,N_1834,N_1895);
or U2645 (N_2645,N_2326,N_1953);
nand U2646 (N_2646,N_2289,N_2378);
nor U2647 (N_2647,N_2086,N_2236);
or U2648 (N_2648,N_2261,N_1876);
or U2649 (N_2649,N_1979,N_1987);
nand U2650 (N_2650,N_2379,N_1892);
or U2651 (N_2651,N_2156,N_1845);
xor U2652 (N_2652,N_2218,N_2098);
nand U2653 (N_2653,N_2036,N_2209);
nor U2654 (N_2654,N_2300,N_2056);
nand U2655 (N_2655,N_2102,N_2262);
and U2656 (N_2656,N_1807,N_1910);
xor U2657 (N_2657,N_2033,N_2187);
and U2658 (N_2658,N_2365,N_2146);
nand U2659 (N_2659,N_1908,N_1919);
nand U2660 (N_2660,N_2047,N_1865);
nor U2661 (N_2661,N_2322,N_1867);
nor U2662 (N_2662,N_2178,N_1869);
and U2663 (N_2663,N_2022,N_2067);
and U2664 (N_2664,N_2061,N_2281);
nand U2665 (N_2665,N_1974,N_1956);
nand U2666 (N_2666,N_2357,N_2270);
and U2667 (N_2667,N_2092,N_2012);
nor U2668 (N_2668,N_2111,N_1920);
nand U2669 (N_2669,N_2216,N_2213);
nor U2670 (N_2670,N_1999,N_2153);
nor U2671 (N_2671,N_2197,N_2226);
and U2672 (N_2672,N_2298,N_2071);
nand U2673 (N_2673,N_2222,N_1928);
nor U2674 (N_2674,N_1872,N_1964);
nor U2675 (N_2675,N_2043,N_2072);
and U2676 (N_2676,N_2142,N_1912);
or U2677 (N_2677,N_2269,N_2371);
or U2678 (N_2678,N_1827,N_2184);
or U2679 (N_2679,N_1815,N_2029);
and U2680 (N_2680,N_2252,N_1881);
or U2681 (N_2681,N_2392,N_2151);
or U2682 (N_2682,N_1804,N_1882);
and U2683 (N_2683,N_1916,N_2131);
nor U2684 (N_2684,N_2026,N_2172);
nand U2685 (N_2685,N_1854,N_2017);
nand U2686 (N_2686,N_1833,N_2130);
and U2687 (N_2687,N_2108,N_2227);
nand U2688 (N_2688,N_1968,N_2059);
nor U2689 (N_2689,N_2039,N_2349);
or U2690 (N_2690,N_2293,N_1877);
or U2691 (N_2691,N_2025,N_1955);
nand U2692 (N_2692,N_2315,N_2001);
and U2693 (N_2693,N_2277,N_1843);
nor U2694 (N_2694,N_2229,N_2219);
nor U2695 (N_2695,N_2110,N_2369);
or U2696 (N_2696,N_1884,N_2080);
nand U2697 (N_2697,N_1853,N_2176);
or U2698 (N_2698,N_1909,N_1856);
nor U2699 (N_2699,N_2062,N_2201);
nand U2700 (N_2700,N_1843,N_1976);
nand U2701 (N_2701,N_2104,N_1984);
and U2702 (N_2702,N_1904,N_2363);
or U2703 (N_2703,N_1874,N_2273);
nand U2704 (N_2704,N_2016,N_1935);
and U2705 (N_2705,N_2240,N_2354);
and U2706 (N_2706,N_1957,N_2383);
or U2707 (N_2707,N_1959,N_2292);
nor U2708 (N_2708,N_1878,N_2390);
nor U2709 (N_2709,N_2139,N_1963);
nor U2710 (N_2710,N_2262,N_2094);
nand U2711 (N_2711,N_2013,N_2265);
nor U2712 (N_2712,N_1806,N_2299);
nand U2713 (N_2713,N_2366,N_2249);
or U2714 (N_2714,N_1958,N_1967);
nor U2715 (N_2715,N_2145,N_1887);
nand U2716 (N_2716,N_1978,N_1939);
or U2717 (N_2717,N_2181,N_2303);
or U2718 (N_2718,N_1806,N_2001);
or U2719 (N_2719,N_2221,N_1879);
and U2720 (N_2720,N_2140,N_2153);
or U2721 (N_2721,N_2152,N_1872);
or U2722 (N_2722,N_1813,N_2020);
or U2723 (N_2723,N_2315,N_2289);
nand U2724 (N_2724,N_2158,N_2159);
and U2725 (N_2725,N_2375,N_2282);
nor U2726 (N_2726,N_2337,N_1919);
nor U2727 (N_2727,N_2106,N_2286);
and U2728 (N_2728,N_2387,N_2360);
nand U2729 (N_2729,N_2037,N_2190);
nor U2730 (N_2730,N_2134,N_2211);
nand U2731 (N_2731,N_1907,N_2004);
nand U2732 (N_2732,N_2287,N_2132);
or U2733 (N_2733,N_2109,N_1825);
and U2734 (N_2734,N_2004,N_2108);
nand U2735 (N_2735,N_2090,N_2136);
nor U2736 (N_2736,N_1885,N_2268);
and U2737 (N_2737,N_2046,N_2278);
or U2738 (N_2738,N_2361,N_1935);
or U2739 (N_2739,N_2112,N_1837);
nor U2740 (N_2740,N_2161,N_1801);
or U2741 (N_2741,N_1925,N_2138);
nand U2742 (N_2742,N_2067,N_1930);
nand U2743 (N_2743,N_2308,N_1889);
nand U2744 (N_2744,N_2236,N_2107);
and U2745 (N_2745,N_2066,N_2091);
and U2746 (N_2746,N_2141,N_2051);
and U2747 (N_2747,N_1895,N_2071);
or U2748 (N_2748,N_1842,N_1948);
nand U2749 (N_2749,N_2159,N_1979);
nand U2750 (N_2750,N_2333,N_2174);
and U2751 (N_2751,N_2252,N_2330);
or U2752 (N_2752,N_2197,N_1837);
nand U2753 (N_2753,N_1854,N_2257);
nand U2754 (N_2754,N_2121,N_2042);
and U2755 (N_2755,N_2096,N_2260);
or U2756 (N_2756,N_2015,N_2293);
and U2757 (N_2757,N_2030,N_2358);
nand U2758 (N_2758,N_2229,N_1822);
nand U2759 (N_2759,N_1916,N_2311);
and U2760 (N_2760,N_2223,N_2276);
or U2761 (N_2761,N_2335,N_2200);
nor U2762 (N_2762,N_1896,N_1932);
nor U2763 (N_2763,N_2309,N_1988);
and U2764 (N_2764,N_1877,N_1929);
nor U2765 (N_2765,N_1910,N_2278);
nand U2766 (N_2766,N_2359,N_2157);
and U2767 (N_2767,N_2152,N_1807);
or U2768 (N_2768,N_2062,N_2189);
and U2769 (N_2769,N_2132,N_2019);
xor U2770 (N_2770,N_2170,N_1993);
nor U2771 (N_2771,N_1889,N_2055);
nand U2772 (N_2772,N_2213,N_2125);
nor U2773 (N_2773,N_1961,N_1822);
and U2774 (N_2774,N_1866,N_2232);
nor U2775 (N_2775,N_2223,N_2102);
nand U2776 (N_2776,N_2030,N_2208);
and U2777 (N_2777,N_1950,N_2144);
or U2778 (N_2778,N_2023,N_2358);
nand U2779 (N_2779,N_1803,N_1855);
and U2780 (N_2780,N_2253,N_2211);
or U2781 (N_2781,N_2138,N_2050);
nand U2782 (N_2782,N_2379,N_2118);
nor U2783 (N_2783,N_1848,N_1997);
or U2784 (N_2784,N_2063,N_2135);
or U2785 (N_2785,N_2371,N_1825);
and U2786 (N_2786,N_1928,N_1823);
nor U2787 (N_2787,N_2240,N_2137);
nor U2788 (N_2788,N_2359,N_2107);
nor U2789 (N_2789,N_2318,N_1982);
or U2790 (N_2790,N_2375,N_1996);
or U2791 (N_2791,N_1958,N_1947);
or U2792 (N_2792,N_2024,N_1971);
and U2793 (N_2793,N_2297,N_2161);
nand U2794 (N_2794,N_2081,N_1804);
nor U2795 (N_2795,N_2022,N_2081);
or U2796 (N_2796,N_2121,N_2270);
or U2797 (N_2797,N_2214,N_2316);
or U2798 (N_2798,N_1928,N_2387);
nor U2799 (N_2799,N_1813,N_2023);
nand U2800 (N_2800,N_2186,N_2002);
nor U2801 (N_2801,N_1810,N_1949);
nor U2802 (N_2802,N_1941,N_2026);
nand U2803 (N_2803,N_2237,N_2252);
nand U2804 (N_2804,N_2316,N_2330);
and U2805 (N_2805,N_1816,N_2113);
and U2806 (N_2806,N_2276,N_1827);
nand U2807 (N_2807,N_2369,N_1928);
or U2808 (N_2808,N_2116,N_1975);
or U2809 (N_2809,N_2032,N_1809);
nor U2810 (N_2810,N_1878,N_1818);
nand U2811 (N_2811,N_2324,N_2116);
and U2812 (N_2812,N_2314,N_2191);
and U2813 (N_2813,N_1940,N_2272);
nand U2814 (N_2814,N_2249,N_1888);
nor U2815 (N_2815,N_1907,N_2066);
nand U2816 (N_2816,N_2096,N_2234);
and U2817 (N_2817,N_2221,N_2012);
nand U2818 (N_2818,N_2006,N_2184);
and U2819 (N_2819,N_2069,N_2025);
xnor U2820 (N_2820,N_1995,N_1897);
nor U2821 (N_2821,N_2030,N_1818);
nor U2822 (N_2822,N_1817,N_2277);
nand U2823 (N_2823,N_2048,N_2040);
nand U2824 (N_2824,N_2095,N_1989);
nand U2825 (N_2825,N_2081,N_2211);
nor U2826 (N_2826,N_2135,N_2311);
and U2827 (N_2827,N_2238,N_2338);
and U2828 (N_2828,N_1830,N_2120);
nand U2829 (N_2829,N_2361,N_2319);
nand U2830 (N_2830,N_1820,N_2045);
or U2831 (N_2831,N_1908,N_1917);
or U2832 (N_2832,N_1925,N_2305);
or U2833 (N_2833,N_2253,N_2348);
nor U2834 (N_2834,N_1918,N_1897);
and U2835 (N_2835,N_2059,N_1800);
and U2836 (N_2836,N_1967,N_2184);
nor U2837 (N_2837,N_2008,N_2094);
nor U2838 (N_2838,N_2222,N_1828);
and U2839 (N_2839,N_1990,N_2139);
and U2840 (N_2840,N_2132,N_2336);
nor U2841 (N_2841,N_2222,N_2230);
and U2842 (N_2842,N_2107,N_2341);
nand U2843 (N_2843,N_2196,N_2297);
or U2844 (N_2844,N_2241,N_2344);
nor U2845 (N_2845,N_2338,N_1860);
nor U2846 (N_2846,N_1857,N_1860);
nor U2847 (N_2847,N_2177,N_1806);
and U2848 (N_2848,N_2258,N_2337);
or U2849 (N_2849,N_2179,N_2187);
or U2850 (N_2850,N_2149,N_2220);
or U2851 (N_2851,N_2090,N_2333);
and U2852 (N_2852,N_2380,N_2255);
nor U2853 (N_2853,N_1825,N_2159);
nor U2854 (N_2854,N_2202,N_1978);
or U2855 (N_2855,N_2353,N_1938);
nor U2856 (N_2856,N_1864,N_1888);
nor U2857 (N_2857,N_1926,N_2145);
nand U2858 (N_2858,N_2328,N_1889);
nand U2859 (N_2859,N_2001,N_2005);
and U2860 (N_2860,N_2131,N_2316);
nor U2861 (N_2861,N_2046,N_2072);
or U2862 (N_2862,N_2112,N_2290);
or U2863 (N_2863,N_2074,N_2030);
xor U2864 (N_2864,N_2015,N_2298);
and U2865 (N_2865,N_2181,N_1838);
nor U2866 (N_2866,N_2330,N_1990);
or U2867 (N_2867,N_2308,N_1927);
nand U2868 (N_2868,N_2264,N_1813);
and U2869 (N_2869,N_1913,N_2099);
or U2870 (N_2870,N_2260,N_1892);
nand U2871 (N_2871,N_2305,N_2136);
nor U2872 (N_2872,N_2049,N_2396);
or U2873 (N_2873,N_2328,N_2060);
or U2874 (N_2874,N_1916,N_1991);
nor U2875 (N_2875,N_2031,N_2112);
or U2876 (N_2876,N_1968,N_2396);
or U2877 (N_2877,N_2310,N_1993);
nand U2878 (N_2878,N_1819,N_2119);
nor U2879 (N_2879,N_2240,N_2251);
or U2880 (N_2880,N_2262,N_2160);
and U2881 (N_2881,N_2025,N_1835);
nor U2882 (N_2882,N_2033,N_1956);
nor U2883 (N_2883,N_2059,N_1852);
nor U2884 (N_2884,N_2145,N_2193);
nand U2885 (N_2885,N_1864,N_2004);
and U2886 (N_2886,N_2189,N_2114);
nand U2887 (N_2887,N_2096,N_1909);
and U2888 (N_2888,N_1927,N_2346);
nor U2889 (N_2889,N_2285,N_2334);
and U2890 (N_2890,N_2239,N_2146);
nand U2891 (N_2891,N_2077,N_2093);
or U2892 (N_2892,N_2153,N_1831);
and U2893 (N_2893,N_2355,N_2235);
nand U2894 (N_2894,N_1858,N_2268);
nor U2895 (N_2895,N_1805,N_1857);
or U2896 (N_2896,N_2228,N_2131);
and U2897 (N_2897,N_1952,N_2336);
nor U2898 (N_2898,N_1922,N_2042);
nand U2899 (N_2899,N_1807,N_1888);
and U2900 (N_2900,N_2334,N_1900);
nor U2901 (N_2901,N_2294,N_2218);
nor U2902 (N_2902,N_2051,N_2227);
nand U2903 (N_2903,N_2391,N_2143);
nand U2904 (N_2904,N_1867,N_2197);
or U2905 (N_2905,N_2021,N_1911);
nor U2906 (N_2906,N_2074,N_2206);
nand U2907 (N_2907,N_2326,N_1834);
nor U2908 (N_2908,N_1860,N_2123);
or U2909 (N_2909,N_2384,N_2240);
and U2910 (N_2910,N_2228,N_2000);
nor U2911 (N_2911,N_2037,N_2382);
or U2912 (N_2912,N_2317,N_1899);
or U2913 (N_2913,N_2113,N_1820);
nor U2914 (N_2914,N_2072,N_1885);
nor U2915 (N_2915,N_2395,N_1895);
or U2916 (N_2916,N_2211,N_1964);
and U2917 (N_2917,N_1828,N_2238);
nor U2918 (N_2918,N_1951,N_1871);
nand U2919 (N_2919,N_2264,N_2143);
and U2920 (N_2920,N_2079,N_2220);
nor U2921 (N_2921,N_2353,N_2347);
and U2922 (N_2922,N_1878,N_2149);
nand U2923 (N_2923,N_2249,N_2352);
or U2924 (N_2924,N_2174,N_2037);
nor U2925 (N_2925,N_1955,N_2014);
or U2926 (N_2926,N_2376,N_2006);
nor U2927 (N_2927,N_2360,N_2386);
and U2928 (N_2928,N_2197,N_2270);
or U2929 (N_2929,N_1877,N_2358);
nand U2930 (N_2930,N_2301,N_2190);
nand U2931 (N_2931,N_2294,N_1801);
nor U2932 (N_2932,N_1922,N_2175);
or U2933 (N_2933,N_1972,N_2205);
nand U2934 (N_2934,N_2132,N_1894);
and U2935 (N_2935,N_2010,N_2240);
or U2936 (N_2936,N_2336,N_2216);
and U2937 (N_2937,N_1965,N_2350);
or U2938 (N_2938,N_2077,N_1840);
and U2939 (N_2939,N_1803,N_1869);
and U2940 (N_2940,N_2173,N_2291);
nand U2941 (N_2941,N_2052,N_1942);
and U2942 (N_2942,N_2105,N_2031);
and U2943 (N_2943,N_1851,N_1943);
nand U2944 (N_2944,N_2243,N_2373);
xor U2945 (N_2945,N_1888,N_2389);
nand U2946 (N_2946,N_2106,N_1942);
or U2947 (N_2947,N_2258,N_2118);
or U2948 (N_2948,N_2195,N_2302);
and U2949 (N_2949,N_1957,N_2048);
nand U2950 (N_2950,N_2257,N_1804);
nand U2951 (N_2951,N_1824,N_2184);
nand U2952 (N_2952,N_2232,N_2379);
nand U2953 (N_2953,N_2272,N_2277);
xor U2954 (N_2954,N_2184,N_2399);
nand U2955 (N_2955,N_1892,N_2329);
nor U2956 (N_2956,N_2394,N_2179);
nor U2957 (N_2957,N_2170,N_1905);
and U2958 (N_2958,N_1944,N_2117);
or U2959 (N_2959,N_2075,N_2299);
xnor U2960 (N_2960,N_2023,N_2269);
and U2961 (N_2961,N_2378,N_2329);
nor U2962 (N_2962,N_2080,N_1839);
or U2963 (N_2963,N_1952,N_2192);
nand U2964 (N_2964,N_2391,N_1912);
or U2965 (N_2965,N_1809,N_2097);
or U2966 (N_2966,N_2026,N_2330);
or U2967 (N_2967,N_2005,N_2181);
or U2968 (N_2968,N_1963,N_2217);
or U2969 (N_2969,N_2378,N_2139);
and U2970 (N_2970,N_2195,N_2043);
or U2971 (N_2971,N_1975,N_2158);
and U2972 (N_2972,N_1842,N_2262);
and U2973 (N_2973,N_1928,N_2064);
or U2974 (N_2974,N_2242,N_1817);
and U2975 (N_2975,N_2020,N_2292);
and U2976 (N_2976,N_2079,N_1902);
nand U2977 (N_2977,N_1897,N_2011);
or U2978 (N_2978,N_1819,N_1821);
nand U2979 (N_2979,N_2339,N_2335);
and U2980 (N_2980,N_2143,N_2048);
xor U2981 (N_2981,N_1979,N_1810);
nor U2982 (N_2982,N_1846,N_2281);
nor U2983 (N_2983,N_1899,N_2053);
nand U2984 (N_2984,N_2055,N_2075);
nand U2985 (N_2985,N_2347,N_1850);
and U2986 (N_2986,N_2195,N_1982);
or U2987 (N_2987,N_1800,N_2373);
and U2988 (N_2988,N_2064,N_2046);
and U2989 (N_2989,N_2277,N_2149);
nand U2990 (N_2990,N_2085,N_1933);
and U2991 (N_2991,N_1877,N_1999);
nor U2992 (N_2992,N_2347,N_2051);
or U2993 (N_2993,N_2336,N_1909);
nand U2994 (N_2994,N_2095,N_2391);
and U2995 (N_2995,N_2297,N_2220);
nor U2996 (N_2996,N_2084,N_2318);
nand U2997 (N_2997,N_2113,N_1924);
and U2998 (N_2998,N_2309,N_1904);
nor U2999 (N_2999,N_1841,N_2116);
and UO_0 (O_0,N_2533,N_2596);
and UO_1 (O_1,N_2659,N_2783);
nand UO_2 (O_2,N_2446,N_2492);
xor UO_3 (O_3,N_2511,N_2697);
nand UO_4 (O_4,N_2407,N_2848);
or UO_5 (O_5,N_2491,N_2456);
xor UO_6 (O_6,N_2925,N_2543);
nor UO_7 (O_7,N_2732,N_2776);
nand UO_8 (O_8,N_2426,N_2453);
nand UO_9 (O_9,N_2849,N_2865);
nand UO_10 (O_10,N_2610,N_2569);
nand UO_11 (O_11,N_2406,N_2825);
and UO_12 (O_12,N_2701,N_2904);
or UO_13 (O_13,N_2837,N_2753);
and UO_14 (O_14,N_2708,N_2726);
and UO_15 (O_15,N_2998,N_2463);
and UO_16 (O_16,N_2704,N_2728);
nor UO_17 (O_17,N_2601,N_2551);
nand UO_18 (O_18,N_2907,N_2950);
nand UO_19 (O_19,N_2789,N_2804);
or UO_20 (O_20,N_2748,N_2488);
and UO_21 (O_21,N_2476,N_2421);
nand UO_22 (O_22,N_2498,N_2740);
nor UO_23 (O_23,N_2892,N_2626);
nand UO_24 (O_24,N_2887,N_2960);
nand UO_25 (O_25,N_2823,N_2768);
nor UO_26 (O_26,N_2425,N_2644);
nor UO_27 (O_27,N_2983,N_2988);
or UO_28 (O_28,N_2869,N_2747);
or UO_29 (O_29,N_2790,N_2878);
and UO_30 (O_30,N_2750,N_2941);
or UO_31 (O_31,N_2741,N_2599);
and UO_32 (O_32,N_2861,N_2400);
nand UO_33 (O_33,N_2975,N_2974);
and UO_34 (O_34,N_2875,N_2549);
or UO_35 (O_35,N_2444,N_2935);
nand UO_36 (O_36,N_2588,N_2594);
nand UO_37 (O_37,N_2884,N_2852);
nor UO_38 (O_38,N_2509,N_2508);
nor UO_39 (O_39,N_2623,N_2868);
and UO_40 (O_40,N_2836,N_2835);
nor UO_41 (O_41,N_2627,N_2537);
and UO_42 (O_42,N_2535,N_2756);
nor UO_43 (O_43,N_2416,N_2777);
or UO_44 (O_44,N_2656,N_2553);
and UO_45 (O_45,N_2763,N_2724);
or UO_46 (O_46,N_2822,N_2710);
or UO_47 (O_47,N_2513,N_2672);
nand UO_48 (O_48,N_2688,N_2735);
or UO_49 (O_49,N_2885,N_2477);
nor UO_50 (O_50,N_2938,N_2413);
and UO_51 (O_51,N_2987,N_2515);
or UO_52 (O_52,N_2678,N_2702);
nor UO_53 (O_53,N_2432,N_2972);
or UO_54 (O_54,N_2690,N_2670);
nand UO_55 (O_55,N_2826,N_2489);
nand UO_56 (O_56,N_2992,N_2954);
xnor UO_57 (O_57,N_2872,N_2854);
nand UO_58 (O_58,N_2454,N_2891);
nor UO_59 (O_59,N_2721,N_2937);
and UO_60 (O_60,N_2745,N_2900);
nand UO_61 (O_61,N_2990,N_2662);
or UO_62 (O_62,N_2729,N_2405);
nor UO_63 (O_63,N_2703,N_2597);
nand UO_64 (O_64,N_2786,N_2720);
nand UO_65 (O_65,N_2566,N_2953);
nand UO_66 (O_66,N_2984,N_2738);
and UO_67 (O_67,N_2445,N_2700);
nor UO_68 (O_68,N_2994,N_2927);
nand UO_69 (O_69,N_2449,N_2734);
nor UO_70 (O_70,N_2810,N_2482);
and UO_71 (O_71,N_2842,N_2814);
or UO_72 (O_72,N_2618,N_2539);
xnor UO_73 (O_73,N_2602,N_2780);
and UO_74 (O_74,N_2465,N_2434);
or UO_75 (O_75,N_2773,N_2595);
nor UO_76 (O_76,N_2430,N_2442);
nand UO_77 (O_77,N_2800,N_2930);
nand UO_78 (O_78,N_2859,N_2796);
or UO_79 (O_79,N_2536,N_2815);
nor UO_80 (O_80,N_2813,N_2468);
or UO_81 (O_81,N_2530,N_2752);
nand UO_82 (O_82,N_2910,N_2547);
nand UO_83 (O_83,N_2824,N_2903);
nor UO_84 (O_84,N_2723,N_2495);
and UO_85 (O_85,N_2467,N_2527);
or UO_86 (O_86,N_2788,N_2794);
or UO_87 (O_87,N_2666,N_2902);
or UO_88 (O_88,N_2531,N_2895);
and UO_89 (O_89,N_2541,N_2685);
or UO_90 (O_90,N_2557,N_2447);
nand UO_91 (O_91,N_2478,N_2739);
and UO_92 (O_92,N_2905,N_2933);
or UO_93 (O_93,N_2830,N_2590);
nor UO_94 (O_94,N_2846,N_2554);
nor UO_95 (O_95,N_2718,N_2612);
or UO_96 (O_96,N_2643,N_2414);
nand UO_97 (O_97,N_2576,N_2562);
and UO_98 (O_98,N_2665,N_2845);
and UO_99 (O_99,N_2673,N_2585);
and UO_100 (O_100,N_2401,N_2567);
nor UO_101 (O_101,N_2521,N_2897);
nor UO_102 (O_102,N_2909,N_2829);
and UO_103 (O_103,N_2419,N_2692);
nor UO_104 (O_104,N_2448,N_2968);
or UO_105 (O_105,N_2879,N_2816);
nand UO_106 (O_106,N_2986,N_2956);
nor UO_107 (O_107,N_2844,N_2713);
nand UO_108 (O_108,N_2642,N_2450);
nor UO_109 (O_109,N_2481,N_2991);
nand UO_110 (O_110,N_2649,N_2969);
and UO_111 (O_111,N_2727,N_2894);
nand UO_112 (O_112,N_2451,N_2742);
nor UO_113 (O_113,N_2962,N_2435);
nor UO_114 (O_114,N_2877,N_2838);
and UO_115 (O_115,N_2946,N_2831);
or UO_116 (O_116,N_2613,N_2751);
and UO_117 (O_117,N_2779,N_2607);
or UO_118 (O_118,N_2422,N_2577);
nand UO_119 (O_119,N_2538,N_2605);
or UO_120 (O_120,N_2841,N_2733);
or UO_121 (O_121,N_2676,N_2973);
nor UO_122 (O_122,N_2943,N_2757);
and UO_123 (O_123,N_2827,N_2646);
nand UO_124 (O_124,N_2514,N_2880);
nor UO_125 (O_125,N_2647,N_2412);
and UO_126 (O_126,N_2455,N_2944);
and UO_127 (O_127,N_2461,N_2918);
or UO_128 (O_128,N_2853,N_2806);
and UO_129 (O_129,N_2486,N_2572);
nor UO_130 (O_130,N_2764,N_2970);
and UO_131 (O_131,N_2696,N_2614);
nor UO_132 (O_132,N_2712,N_2522);
or UO_133 (O_133,N_2843,N_2559);
nand UO_134 (O_134,N_2939,N_2801);
xor UO_135 (O_135,N_2948,N_2929);
nor UO_136 (O_136,N_2743,N_2667);
nor UO_137 (O_137,N_2487,N_2862);
nor UO_138 (O_138,N_2893,N_2867);
and UO_139 (O_139,N_2581,N_2999);
or UO_140 (O_140,N_2663,N_2469);
nor UO_141 (O_141,N_2997,N_2638);
or UO_142 (O_142,N_2617,N_2503);
nor UO_143 (O_143,N_2424,N_2512);
nand UO_144 (O_144,N_2959,N_2494);
nand UO_145 (O_145,N_2771,N_2571);
nor UO_146 (O_146,N_2466,N_2808);
or UO_147 (O_147,N_2803,N_2631);
or UO_148 (O_148,N_2716,N_2528);
nand UO_149 (O_149,N_2410,N_2525);
and UO_150 (O_150,N_2499,N_2565);
or UO_151 (O_151,N_2811,N_2587);
or UO_152 (O_152,N_2493,N_2709);
nor UO_153 (O_153,N_2978,N_2661);
or UO_154 (O_154,N_2655,N_2749);
or UO_155 (O_155,N_2504,N_2886);
and UO_156 (O_156,N_2603,N_2479);
and UO_157 (O_157,N_2573,N_2687);
nor UO_158 (O_158,N_2650,N_2634);
and UO_159 (O_159,N_2715,N_2855);
xnor UO_160 (O_160,N_2438,N_2622);
or UO_161 (O_161,N_2961,N_2473);
and UO_162 (O_162,N_2611,N_2427);
or UO_163 (O_163,N_2758,N_2985);
nand UO_164 (O_164,N_2653,N_2964);
nand UO_165 (O_165,N_2575,N_2589);
or UO_166 (O_166,N_2660,N_2963);
nand UO_167 (O_167,N_2934,N_2586);
or UO_168 (O_168,N_2440,N_2698);
or UO_169 (O_169,N_2420,N_2408);
nor UO_170 (O_170,N_2564,N_2923);
nand UO_171 (O_171,N_2847,N_2669);
xnor UO_172 (O_172,N_2922,N_2532);
xor UO_173 (O_173,N_2664,N_2797);
nor UO_174 (O_174,N_2980,N_2402);
nand UO_175 (O_175,N_2439,N_2632);
or UO_176 (O_176,N_2556,N_2819);
nor UO_177 (O_177,N_2470,N_2785);
and UO_178 (O_178,N_2529,N_2926);
nor UO_179 (O_179,N_2637,N_2496);
and UO_180 (O_180,N_2686,N_2545);
nor UO_181 (O_181,N_2462,N_2876);
nand UO_182 (O_182,N_2707,N_2863);
xnor UO_183 (O_183,N_2722,N_2888);
nor UO_184 (O_184,N_2472,N_2982);
nand UO_185 (O_185,N_2931,N_2693);
and UO_186 (O_186,N_2592,N_2570);
nand UO_187 (O_187,N_2681,N_2654);
and UO_188 (O_188,N_2608,N_2787);
nand UO_189 (O_189,N_2736,N_2624);
nand UO_190 (O_190,N_2677,N_2730);
nor UO_191 (O_191,N_2593,N_2609);
nor UO_192 (O_192,N_2981,N_2744);
nor UO_193 (O_193,N_2898,N_2520);
nand UO_194 (O_194,N_2917,N_2807);
nand UO_195 (O_195,N_2967,N_2415);
and UO_196 (O_196,N_2851,N_2431);
nor UO_197 (O_197,N_2640,N_2755);
nand UO_198 (O_198,N_2404,N_2674);
nand UO_199 (O_199,N_2578,N_2552);
or UO_200 (O_200,N_2652,N_2574);
nor UO_201 (O_201,N_2915,N_2809);
or UO_202 (O_202,N_2436,N_2714);
nor UO_203 (O_203,N_2598,N_2616);
or UO_204 (O_204,N_2546,N_2857);
nor UO_205 (O_205,N_2770,N_2784);
and UO_206 (O_206,N_2914,N_2782);
nand UO_207 (O_207,N_2719,N_2890);
nand UO_208 (O_208,N_2497,N_2550);
or UO_209 (O_209,N_2615,N_2899);
or UO_210 (O_210,N_2940,N_2474);
nand UO_211 (O_211,N_2629,N_2500);
nor UO_212 (O_212,N_2641,N_2924);
xnor UO_213 (O_213,N_2799,N_2684);
or UO_214 (O_214,N_2584,N_2619);
or UO_215 (O_215,N_2418,N_2699);
nand UO_216 (O_216,N_2871,N_2883);
nor UO_217 (O_217,N_2912,N_2945);
nor UO_218 (O_218,N_2630,N_2490);
and UO_219 (O_219,N_2977,N_2775);
nor UO_220 (O_220,N_2458,N_2766);
nand UO_221 (O_221,N_2913,N_2437);
or UO_222 (O_222,N_2942,N_2648);
nor UO_223 (O_223,N_2821,N_2475);
or UO_224 (O_224,N_2772,N_2639);
or UO_225 (O_225,N_2901,N_2731);
and UO_226 (O_226,N_2561,N_2621);
nand UO_227 (O_227,N_2812,N_2761);
and UO_228 (O_228,N_2460,N_2548);
nand UO_229 (O_229,N_2781,N_2441);
nor UO_230 (O_230,N_2778,N_2896);
and UO_231 (O_231,N_2563,N_2881);
or UO_232 (O_232,N_2671,N_2820);
nor UO_233 (O_233,N_2517,N_2452);
nand UO_234 (O_234,N_2502,N_2409);
or UO_235 (O_235,N_2464,N_2657);
and UO_236 (O_236,N_2429,N_2568);
and UO_237 (O_237,N_2911,N_2580);
nor UO_238 (O_238,N_2759,N_2765);
or UO_239 (O_239,N_2832,N_2484);
xor UO_240 (O_240,N_2874,N_2866);
nand UO_241 (O_241,N_2762,N_2850);
or UO_242 (O_242,N_2633,N_2966);
nor UO_243 (O_243,N_2403,N_2417);
or UO_244 (O_244,N_2480,N_2620);
or UO_245 (O_245,N_2889,N_2955);
or UO_246 (O_246,N_2754,N_2995);
and UO_247 (O_247,N_2428,N_2706);
and UO_248 (O_248,N_2864,N_2993);
nand UO_249 (O_249,N_2635,N_2711);
nand UO_250 (O_250,N_2658,N_2856);
nand UO_251 (O_251,N_2947,N_2604);
nor UO_252 (O_252,N_2979,N_2834);
nor UO_253 (O_253,N_2774,N_2510);
nor UO_254 (O_254,N_2443,N_2996);
nor UO_255 (O_255,N_2818,N_2833);
or UO_256 (O_256,N_2989,N_2952);
or UO_257 (O_257,N_2628,N_2555);
and UO_258 (O_258,N_2506,N_2583);
or UO_259 (O_259,N_2957,N_2936);
and UO_260 (O_260,N_2518,N_2958);
and UO_261 (O_261,N_2858,N_2683);
nand UO_262 (O_262,N_2651,N_2524);
or UO_263 (O_263,N_2908,N_2919);
and UO_264 (O_264,N_2680,N_2507);
and UO_265 (O_265,N_2802,N_2725);
nand UO_266 (O_266,N_2600,N_2873);
or UO_267 (O_267,N_2928,N_2691);
nand UO_268 (O_268,N_2793,N_2526);
nor UO_269 (O_269,N_2860,N_2951);
xor UO_270 (O_270,N_2689,N_2679);
or UO_271 (O_271,N_2817,N_2457);
xor UO_272 (O_272,N_2976,N_2916);
nor UO_273 (O_273,N_2839,N_2949);
and UO_274 (O_274,N_2636,N_2920);
and UO_275 (O_275,N_2798,N_2540);
and UO_276 (O_276,N_2519,N_2791);
nor UO_277 (O_277,N_2523,N_2737);
nand UO_278 (O_278,N_2717,N_2932);
or UO_279 (O_279,N_2534,N_2483);
and UO_280 (O_280,N_2805,N_2870);
nand UO_281 (O_281,N_2767,N_2544);
or UO_282 (O_282,N_2471,N_2501);
nand UO_283 (O_283,N_2423,N_2705);
or UO_284 (O_284,N_2882,N_2582);
or UO_285 (O_285,N_2625,N_2459);
nor UO_286 (O_286,N_2485,N_2695);
and UO_287 (O_287,N_2746,N_2675);
nor UO_288 (O_288,N_2591,N_2921);
and UO_289 (O_289,N_2505,N_2694);
or UO_290 (O_290,N_2542,N_2795);
nand UO_291 (O_291,N_2645,N_2769);
nor UO_292 (O_292,N_2606,N_2516);
and UO_293 (O_293,N_2840,N_2828);
and UO_294 (O_294,N_2433,N_2971);
nand UO_295 (O_295,N_2668,N_2965);
nor UO_296 (O_296,N_2792,N_2579);
nand UO_297 (O_297,N_2682,N_2558);
or UO_298 (O_298,N_2411,N_2906);
nand UO_299 (O_299,N_2760,N_2560);
nand UO_300 (O_300,N_2835,N_2471);
or UO_301 (O_301,N_2554,N_2849);
nand UO_302 (O_302,N_2893,N_2546);
nor UO_303 (O_303,N_2846,N_2789);
xnor UO_304 (O_304,N_2885,N_2956);
nand UO_305 (O_305,N_2721,N_2499);
or UO_306 (O_306,N_2520,N_2996);
nand UO_307 (O_307,N_2411,N_2806);
xor UO_308 (O_308,N_2508,N_2410);
nand UO_309 (O_309,N_2491,N_2455);
nor UO_310 (O_310,N_2695,N_2633);
nand UO_311 (O_311,N_2954,N_2505);
nand UO_312 (O_312,N_2446,N_2501);
and UO_313 (O_313,N_2623,N_2911);
or UO_314 (O_314,N_2801,N_2947);
nand UO_315 (O_315,N_2510,N_2690);
and UO_316 (O_316,N_2869,N_2622);
and UO_317 (O_317,N_2593,N_2565);
or UO_318 (O_318,N_2699,N_2742);
and UO_319 (O_319,N_2696,N_2581);
nand UO_320 (O_320,N_2900,N_2523);
and UO_321 (O_321,N_2896,N_2464);
nor UO_322 (O_322,N_2989,N_2878);
nand UO_323 (O_323,N_2709,N_2896);
or UO_324 (O_324,N_2497,N_2983);
or UO_325 (O_325,N_2948,N_2972);
nor UO_326 (O_326,N_2993,N_2771);
and UO_327 (O_327,N_2501,N_2472);
or UO_328 (O_328,N_2892,N_2569);
and UO_329 (O_329,N_2529,N_2989);
and UO_330 (O_330,N_2435,N_2849);
nand UO_331 (O_331,N_2731,N_2544);
or UO_332 (O_332,N_2491,N_2830);
and UO_333 (O_333,N_2753,N_2917);
nand UO_334 (O_334,N_2937,N_2779);
and UO_335 (O_335,N_2640,N_2822);
and UO_336 (O_336,N_2741,N_2519);
and UO_337 (O_337,N_2460,N_2811);
nor UO_338 (O_338,N_2807,N_2929);
nand UO_339 (O_339,N_2980,N_2743);
or UO_340 (O_340,N_2884,N_2879);
nor UO_341 (O_341,N_2758,N_2639);
and UO_342 (O_342,N_2753,N_2956);
and UO_343 (O_343,N_2585,N_2633);
or UO_344 (O_344,N_2623,N_2563);
or UO_345 (O_345,N_2618,N_2658);
and UO_346 (O_346,N_2492,N_2510);
nor UO_347 (O_347,N_2477,N_2807);
nand UO_348 (O_348,N_2813,N_2429);
or UO_349 (O_349,N_2822,N_2648);
or UO_350 (O_350,N_2663,N_2953);
nand UO_351 (O_351,N_2511,N_2585);
nor UO_352 (O_352,N_2788,N_2740);
or UO_353 (O_353,N_2979,N_2719);
or UO_354 (O_354,N_2519,N_2607);
nor UO_355 (O_355,N_2479,N_2616);
and UO_356 (O_356,N_2558,N_2552);
or UO_357 (O_357,N_2727,N_2838);
nand UO_358 (O_358,N_2849,N_2907);
nand UO_359 (O_359,N_2504,N_2490);
and UO_360 (O_360,N_2573,N_2420);
and UO_361 (O_361,N_2780,N_2427);
nor UO_362 (O_362,N_2853,N_2773);
and UO_363 (O_363,N_2615,N_2850);
and UO_364 (O_364,N_2698,N_2822);
and UO_365 (O_365,N_2832,N_2767);
nand UO_366 (O_366,N_2633,N_2638);
or UO_367 (O_367,N_2963,N_2857);
and UO_368 (O_368,N_2439,N_2850);
nand UO_369 (O_369,N_2668,N_2549);
nor UO_370 (O_370,N_2963,N_2914);
nand UO_371 (O_371,N_2645,N_2690);
or UO_372 (O_372,N_2663,N_2666);
nor UO_373 (O_373,N_2948,N_2677);
nand UO_374 (O_374,N_2482,N_2459);
and UO_375 (O_375,N_2736,N_2909);
and UO_376 (O_376,N_2794,N_2935);
nand UO_377 (O_377,N_2513,N_2914);
and UO_378 (O_378,N_2698,N_2997);
nand UO_379 (O_379,N_2841,N_2783);
nor UO_380 (O_380,N_2854,N_2618);
nor UO_381 (O_381,N_2414,N_2881);
and UO_382 (O_382,N_2606,N_2779);
nand UO_383 (O_383,N_2968,N_2667);
or UO_384 (O_384,N_2500,N_2984);
and UO_385 (O_385,N_2522,N_2588);
nor UO_386 (O_386,N_2420,N_2658);
nand UO_387 (O_387,N_2459,N_2914);
nor UO_388 (O_388,N_2905,N_2827);
and UO_389 (O_389,N_2744,N_2613);
or UO_390 (O_390,N_2839,N_2488);
or UO_391 (O_391,N_2708,N_2830);
nand UO_392 (O_392,N_2952,N_2597);
nand UO_393 (O_393,N_2964,N_2823);
nand UO_394 (O_394,N_2439,N_2946);
nand UO_395 (O_395,N_2689,N_2528);
or UO_396 (O_396,N_2726,N_2627);
nor UO_397 (O_397,N_2888,N_2511);
nand UO_398 (O_398,N_2535,N_2547);
or UO_399 (O_399,N_2859,N_2968);
or UO_400 (O_400,N_2678,N_2810);
nor UO_401 (O_401,N_2862,N_2550);
nand UO_402 (O_402,N_2946,N_2633);
or UO_403 (O_403,N_2572,N_2813);
and UO_404 (O_404,N_2946,N_2485);
or UO_405 (O_405,N_2879,N_2525);
and UO_406 (O_406,N_2489,N_2745);
or UO_407 (O_407,N_2756,N_2430);
or UO_408 (O_408,N_2548,N_2586);
and UO_409 (O_409,N_2796,N_2645);
and UO_410 (O_410,N_2901,N_2565);
and UO_411 (O_411,N_2465,N_2892);
and UO_412 (O_412,N_2983,N_2476);
nor UO_413 (O_413,N_2596,N_2802);
nor UO_414 (O_414,N_2989,N_2400);
or UO_415 (O_415,N_2631,N_2640);
nor UO_416 (O_416,N_2827,N_2752);
and UO_417 (O_417,N_2576,N_2784);
or UO_418 (O_418,N_2612,N_2457);
nand UO_419 (O_419,N_2872,N_2622);
or UO_420 (O_420,N_2475,N_2930);
and UO_421 (O_421,N_2539,N_2589);
or UO_422 (O_422,N_2581,N_2708);
nor UO_423 (O_423,N_2837,N_2483);
or UO_424 (O_424,N_2955,N_2992);
nand UO_425 (O_425,N_2988,N_2405);
nor UO_426 (O_426,N_2780,N_2420);
nor UO_427 (O_427,N_2720,N_2963);
and UO_428 (O_428,N_2967,N_2733);
and UO_429 (O_429,N_2510,N_2948);
nand UO_430 (O_430,N_2780,N_2804);
nor UO_431 (O_431,N_2634,N_2663);
nand UO_432 (O_432,N_2762,N_2407);
nand UO_433 (O_433,N_2477,N_2431);
nand UO_434 (O_434,N_2725,N_2718);
nand UO_435 (O_435,N_2487,N_2613);
or UO_436 (O_436,N_2711,N_2626);
and UO_437 (O_437,N_2572,N_2617);
nor UO_438 (O_438,N_2411,N_2703);
and UO_439 (O_439,N_2457,N_2619);
or UO_440 (O_440,N_2717,N_2593);
or UO_441 (O_441,N_2698,N_2844);
or UO_442 (O_442,N_2983,N_2460);
nand UO_443 (O_443,N_2760,N_2495);
nor UO_444 (O_444,N_2748,N_2719);
nand UO_445 (O_445,N_2988,N_2637);
and UO_446 (O_446,N_2526,N_2494);
nand UO_447 (O_447,N_2772,N_2746);
or UO_448 (O_448,N_2727,N_2499);
and UO_449 (O_449,N_2925,N_2534);
and UO_450 (O_450,N_2818,N_2663);
nand UO_451 (O_451,N_2978,N_2893);
nand UO_452 (O_452,N_2909,N_2800);
nand UO_453 (O_453,N_2645,N_2838);
nand UO_454 (O_454,N_2982,N_2830);
or UO_455 (O_455,N_2407,N_2481);
or UO_456 (O_456,N_2565,N_2573);
nor UO_457 (O_457,N_2930,N_2982);
nor UO_458 (O_458,N_2850,N_2642);
or UO_459 (O_459,N_2999,N_2961);
or UO_460 (O_460,N_2727,N_2658);
or UO_461 (O_461,N_2977,N_2720);
and UO_462 (O_462,N_2629,N_2950);
or UO_463 (O_463,N_2421,N_2798);
and UO_464 (O_464,N_2671,N_2621);
nor UO_465 (O_465,N_2481,N_2885);
and UO_466 (O_466,N_2546,N_2793);
nand UO_467 (O_467,N_2565,N_2594);
nor UO_468 (O_468,N_2959,N_2762);
nand UO_469 (O_469,N_2892,N_2417);
nand UO_470 (O_470,N_2563,N_2843);
or UO_471 (O_471,N_2914,N_2558);
nand UO_472 (O_472,N_2538,N_2483);
or UO_473 (O_473,N_2477,N_2766);
and UO_474 (O_474,N_2769,N_2780);
or UO_475 (O_475,N_2878,N_2507);
and UO_476 (O_476,N_2646,N_2825);
and UO_477 (O_477,N_2900,N_2787);
nor UO_478 (O_478,N_2586,N_2539);
nand UO_479 (O_479,N_2964,N_2462);
nor UO_480 (O_480,N_2795,N_2966);
or UO_481 (O_481,N_2566,N_2502);
nand UO_482 (O_482,N_2833,N_2587);
or UO_483 (O_483,N_2743,N_2424);
and UO_484 (O_484,N_2858,N_2446);
nand UO_485 (O_485,N_2477,N_2724);
nor UO_486 (O_486,N_2707,N_2745);
and UO_487 (O_487,N_2464,N_2835);
nand UO_488 (O_488,N_2813,N_2683);
or UO_489 (O_489,N_2448,N_2839);
nor UO_490 (O_490,N_2757,N_2736);
or UO_491 (O_491,N_2505,N_2929);
or UO_492 (O_492,N_2445,N_2405);
or UO_493 (O_493,N_2546,N_2526);
nor UO_494 (O_494,N_2796,N_2814);
or UO_495 (O_495,N_2443,N_2737);
or UO_496 (O_496,N_2677,N_2822);
and UO_497 (O_497,N_2619,N_2595);
nand UO_498 (O_498,N_2776,N_2648);
nand UO_499 (O_499,N_2503,N_2925);
endmodule