module basic_500_3000_500_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_405,In_7);
and U1 (N_1,In_442,In_498);
or U2 (N_2,In_11,In_398);
xnor U3 (N_3,In_157,In_55);
nand U4 (N_4,In_263,In_258);
xor U5 (N_5,In_423,In_485);
nor U6 (N_6,In_205,In_23);
nor U7 (N_7,In_289,In_220);
nand U8 (N_8,In_381,In_100);
nand U9 (N_9,In_51,In_169);
and U10 (N_10,In_76,In_265);
or U11 (N_11,In_111,In_363);
xor U12 (N_12,In_62,In_217);
nor U13 (N_13,In_12,In_104);
xnor U14 (N_14,In_449,In_224);
nor U15 (N_15,In_88,In_207);
xor U16 (N_16,In_186,In_252);
and U17 (N_17,In_251,In_378);
nand U18 (N_18,In_313,In_479);
or U19 (N_19,In_216,In_57);
or U20 (N_20,In_326,In_61);
or U21 (N_21,In_191,In_60);
nor U22 (N_22,In_358,In_180);
and U23 (N_23,In_310,In_283);
nand U24 (N_24,In_330,In_231);
nand U25 (N_25,In_379,In_236);
and U26 (N_26,In_126,In_245);
nand U27 (N_27,In_412,In_271);
or U28 (N_28,In_113,In_455);
nor U29 (N_29,In_377,In_78);
nand U30 (N_30,In_346,In_254);
nand U31 (N_31,In_425,In_345);
nor U32 (N_32,In_431,In_153);
or U33 (N_33,In_452,In_305);
and U34 (N_34,In_144,In_44);
or U35 (N_35,In_360,In_471);
or U36 (N_36,In_351,In_323);
or U37 (N_37,In_47,In_404);
or U38 (N_38,In_63,In_112);
or U39 (N_39,In_80,In_376);
nand U40 (N_40,In_204,In_141);
nor U41 (N_41,In_149,In_364);
nor U42 (N_42,In_30,In_71);
nand U43 (N_43,In_403,In_460);
or U44 (N_44,In_188,In_136);
xnor U45 (N_45,In_170,In_147);
nor U46 (N_46,In_84,In_318);
nand U47 (N_47,In_53,In_439);
or U48 (N_48,In_337,In_266);
and U49 (N_49,In_120,In_371);
and U50 (N_50,In_117,In_419);
nor U51 (N_51,In_276,In_480);
and U52 (N_52,In_122,In_331);
nand U53 (N_53,In_50,In_278);
nor U54 (N_54,In_168,In_394);
nand U55 (N_55,In_262,In_66);
and U56 (N_56,In_464,In_357);
and U57 (N_57,In_13,In_83);
and U58 (N_58,In_70,In_467);
nand U59 (N_59,In_465,In_154);
nor U60 (N_60,In_417,In_230);
or U61 (N_61,In_274,N_34);
nand U62 (N_62,In_185,In_174);
and U63 (N_63,In_332,In_20);
nand U64 (N_64,N_19,In_253);
or U65 (N_65,In_118,In_409);
xnor U66 (N_66,In_21,In_34);
or U67 (N_67,In_290,In_334);
nand U68 (N_68,In_56,In_416);
or U69 (N_69,In_82,In_375);
and U70 (N_70,In_396,In_336);
xnor U71 (N_71,N_22,In_324);
or U72 (N_72,In_384,In_408);
xor U73 (N_73,In_355,In_247);
and U74 (N_74,N_26,In_68);
and U75 (N_75,In_94,In_132);
nand U76 (N_76,In_31,In_99);
nand U77 (N_77,In_308,In_478);
nand U78 (N_78,In_158,In_294);
and U79 (N_79,In_52,In_472);
xnor U80 (N_80,In_487,In_194);
xor U81 (N_81,N_36,In_382);
and U82 (N_82,N_4,N_25);
nor U83 (N_83,In_429,In_182);
and U84 (N_84,In_391,In_219);
or U85 (N_85,In_352,In_228);
nand U86 (N_86,In_361,N_0);
nand U87 (N_87,N_10,In_192);
or U88 (N_88,In_437,In_415);
and U89 (N_89,In_243,N_32);
nor U90 (N_90,In_295,In_125);
nor U91 (N_91,In_495,In_386);
or U92 (N_92,In_493,In_162);
or U93 (N_93,In_299,N_48);
xor U94 (N_94,In_264,In_356);
xnor U95 (N_95,N_42,In_282);
or U96 (N_96,In_447,In_223);
or U97 (N_97,In_444,In_476);
nor U98 (N_98,In_209,In_221);
or U99 (N_99,In_333,In_427);
xnor U100 (N_100,In_463,In_5);
nand U101 (N_101,In_275,In_183);
nand U102 (N_102,In_319,In_212);
nor U103 (N_103,In_89,In_67);
nand U104 (N_104,In_4,N_18);
xor U105 (N_105,In_206,In_75);
and U106 (N_106,In_309,In_387);
and U107 (N_107,In_281,In_6);
nand U108 (N_108,In_291,In_414);
nand U109 (N_109,In_106,In_389);
nor U110 (N_110,In_422,In_448);
and U111 (N_111,N_8,In_321);
nor U112 (N_112,In_108,N_13);
and U113 (N_113,In_250,In_229);
and U114 (N_114,In_232,In_369);
and U115 (N_115,In_46,In_8);
nor U116 (N_116,In_164,In_41);
or U117 (N_117,In_165,In_33);
or U118 (N_118,N_35,N_59);
and U119 (N_119,In_139,In_298);
nor U120 (N_120,N_54,In_246);
xor U121 (N_121,N_45,In_202);
and U122 (N_122,In_443,N_23);
nor U123 (N_123,N_57,In_240);
xor U124 (N_124,In_436,In_344);
xor U125 (N_125,In_15,N_65);
nor U126 (N_126,In_311,In_244);
nor U127 (N_127,N_61,In_114);
or U128 (N_128,In_433,N_82);
nor U129 (N_129,In_26,In_441);
and U130 (N_130,In_201,In_198);
nand U131 (N_131,In_137,In_187);
or U132 (N_132,In_193,N_12);
nor U133 (N_133,In_374,In_285);
nand U134 (N_134,N_79,In_435);
and U135 (N_135,In_167,In_257);
xor U136 (N_136,In_72,In_348);
xor U137 (N_137,N_94,In_163);
xor U138 (N_138,In_1,In_73);
nand U139 (N_139,In_37,N_92);
or U140 (N_140,In_36,N_89);
or U141 (N_141,In_411,N_110);
and U142 (N_142,In_45,In_401);
or U143 (N_143,In_0,In_155);
nand U144 (N_144,In_359,In_19);
nor U145 (N_145,In_256,N_97);
or U146 (N_146,In_372,N_91);
nand U147 (N_147,In_316,In_325);
nor U148 (N_148,N_17,In_119);
and U149 (N_149,N_114,In_85);
nor U150 (N_150,In_430,In_179);
nor U151 (N_151,In_453,In_488);
nor U152 (N_152,In_211,N_15);
and U153 (N_153,In_134,In_123);
or U154 (N_154,In_484,In_197);
xor U155 (N_155,In_64,In_91);
or U156 (N_156,In_96,N_77);
and U157 (N_157,N_95,In_184);
xor U158 (N_158,In_312,In_335);
or U159 (N_159,N_58,In_367);
xnor U160 (N_160,In_454,N_30);
nand U161 (N_161,N_86,N_87);
nand U162 (N_162,N_60,N_1);
nand U163 (N_163,In_473,In_392);
or U164 (N_164,In_420,In_16);
nor U165 (N_165,N_49,N_50);
and U166 (N_166,In_90,In_29);
or U167 (N_167,In_74,In_199);
xnor U168 (N_168,N_3,In_65);
nand U169 (N_169,N_111,N_100);
and U170 (N_170,In_426,In_272);
and U171 (N_171,N_103,In_397);
and U172 (N_172,In_116,In_434);
or U173 (N_173,In_424,In_77);
xor U174 (N_174,In_421,In_286);
and U175 (N_175,In_215,In_292);
or U176 (N_176,N_51,N_62);
or U177 (N_177,In_69,In_457);
and U178 (N_178,N_72,In_92);
nand U179 (N_179,In_297,In_59);
and U180 (N_180,In_368,In_400);
xor U181 (N_181,In_273,N_159);
xnor U182 (N_182,N_123,In_79);
nand U183 (N_183,In_418,In_482);
xor U184 (N_184,In_135,In_131);
xor U185 (N_185,N_172,In_402);
xnor U186 (N_186,In_172,N_29);
nor U187 (N_187,In_343,In_269);
xnor U188 (N_188,In_38,In_115);
nor U189 (N_189,N_129,In_87);
xnor U190 (N_190,N_7,In_238);
and U191 (N_191,In_200,N_43);
and U192 (N_192,In_239,In_210);
nor U193 (N_193,In_48,In_49);
or U194 (N_194,In_314,In_339);
or U195 (N_195,N_132,N_24);
nor U196 (N_196,In_268,In_341);
xnor U197 (N_197,N_76,N_38);
nand U198 (N_198,N_83,In_196);
nor U199 (N_199,N_153,N_127);
nand U200 (N_200,N_63,In_35);
xnor U201 (N_201,In_181,In_171);
or U202 (N_202,In_303,N_39);
and U203 (N_203,In_327,N_64);
nor U204 (N_204,In_320,In_474);
xnor U205 (N_205,In_161,In_296);
xnor U206 (N_206,N_71,N_78);
xor U207 (N_207,In_17,In_300);
and U208 (N_208,In_176,N_108);
xor U209 (N_209,N_116,In_160);
nand U210 (N_210,N_68,In_304);
or U211 (N_211,In_28,In_128);
nand U212 (N_212,In_148,In_248);
and U213 (N_213,In_225,N_47);
nor U214 (N_214,In_97,N_93);
and U215 (N_215,N_117,N_109);
xor U216 (N_216,In_481,N_148);
and U217 (N_217,N_141,In_350);
xnor U218 (N_218,In_383,In_25);
xnor U219 (N_219,In_302,In_173);
or U220 (N_220,N_113,In_143);
nand U221 (N_221,In_407,In_390);
nor U222 (N_222,N_81,In_178);
and U223 (N_223,N_178,In_151);
nor U224 (N_224,In_475,N_143);
and U225 (N_225,N_53,In_9);
or U226 (N_226,N_27,In_105);
and U227 (N_227,In_489,In_190);
nand U228 (N_228,In_456,In_491);
and U229 (N_229,In_293,In_365);
nor U230 (N_230,In_329,N_69);
nand U231 (N_231,In_301,In_459);
xor U232 (N_232,In_203,N_121);
or U233 (N_233,In_121,In_146);
or U234 (N_234,In_42,In_152);
xor U235 (N_235,N_73,N_90);
and U236 (N_236,N_174,In_462);
and U237 (N_237,N_162,In_445);
nor U238 (N_238,In_10,N_101);
nor U239 (N_239,N_28,N_144);
xnor U240 (N_240,In_140,N_183);
or U241 (N_241,N_186,In_24);
nand U242 (N_242,In_142,N_158);
or U243 (N_243,N_119,N_215);
nor U244 (N_244,N_176,In_342);
and U245 (N_245,In_393,N_31);
or U246 (N_246,N_197,N_37);
nand U247 (N_247,N_160,N_140);
or U248 (N_248,N_96,In_410);
nor U249 (N_249,N_207,N_212);
or U250 (N_250,In_492,N_181);
nand U251 (N_251,N_238,N_224);
xnor U252 (N_252,In_226,In_54);
xor U253 (N_253,N_193,In_288);
nor U254 (N_254,In_241,N_175);
xnor U255 (N_255,N_122,N_164);
or U256 (N_256,N_201,N_66);
nand U257 (N_257,In_438,In_189);
or U258 (N_258,N_232,N_152);
xnor U259 (N_259,In_446,N_217);
nor U260 (N_260,In_340,N_102);
xor U261 (N_261,In_237,In_499);
or U262 (N_262,N_84,N_112);
nand U263 (N_263,N_204,N_105);
or U264 (N_264,N_157,In_129);
nor U265 (N_265,In_103,In_477);
and U266 (N_266,N_115,N_211);
and U267 (N_267,In_496,N_40);
or U268 (N_268,In_267,N_55);
nand U269 (N_269,N_206,In_322);
nor U270 (N_270,In_40,In_195);
nor U271 (N_271,N_169,N_52);
xor U272 (N_272,In_440,N_184);
and U273 (N_273,In_385,N_104);
or U274 (N_274,N_220,N_214);
and U275 (N_275,N_191,In_451);
xor U276 (N_276,N_21,N_227);
nor U277 (N_277,In_406,N_170);
nor U278 (N_278,N_223,N_219);
and U279 (N_279,N_5,N_146);
nand U280 (N_280,In_107,N_145);
or U281 (N_281,In_27,In_338);
nor U282 (N_282,N_185,N_130);
nand U283 (N_283,N_156,In_156);
and U284 (N_284,N_75,N_222);
xor U285 (N_285,N_177,N_189);
xnor U286 (N_286,In_175,In_287);
or U287 (N_287,In_213,N_221);
xnor U288 (N_288,In_413,N_188);
and U289 (N_289,N_88,In_255);
nand U290 (N_290,N_203,In_124);
xor U291 (N_291,In_222,N_182);
or U292 (N_292,In_110,In_306);
nor U293 (N_293,In_469,N_142);
xnor U294 (N_294,In_208,In_249);
nand U295 (N_295,In_43,N_139);
or U296 (N_296,N_234,N_237);
and U297 (N_297,N_161,N_155);
nor U298 (N_298,In_483,N_14);
or U299 (N_299,N_41,N_179);
nor U300 (N_300,N_70,N_6);
and U301 (N_301,N_126,N_180);
and U302 (N_302,In_349,N_163);
xor U303 (N_303,N_165,N_279);
xor U304 (N_304,N_297,In_14);
or U305 (N_305,In_395,In_22);
xor U306 (N_306,N_283,N_290);
nand U307 (N_307,In_497,N_216);
nand U308 (N_308,In_315,In_18);
and U309 (N_309,In_461,N_299);
xor U310 (N_310,In_138,In_58);
nand U311 (N_311,In_159,In_234);
nor U312 (N_312,N_138,In_32);
or U313 (N_313,N_276,In_277);
and U314 (N_314,N_128,In_145);
nor U315 (N_315,In_166,N_125);
xnor U316 (N_316,N_289,In_307);
and U317 (N_317,N_257,In_95);
and U318 (N_318,N_173,In_259);
and U319 (N_319,N_229,N_2);
or U320 (N_320,N_275,N_284);
and U321 (N_321,N_209,In_260);
xnor U322 (N_322,In_458,N_208);
nor U323 (N_323,N_171,N_67);
or U324 (N_324,N_98,N_274);
xor U325 (N_325,In_366,In_347);
xnor U326 (N_326,N_271,N_259);
nand U327 (N_327,N_198,N_251);
or U328 (N_328,N_277,N_147);
nor U329 (N_329,N_267,In_450);
nor U330 (N_330,In_353,In_280);
or U331 (N_331,In_399,N_151);
xor U332 (N_332,In_177,N_252);
or U333 (N_333,In_233,N_33);
nand U334 (N_334,N_137,N_44);
or U335 (N_335,N_241,N_133);
xor U336 (N_336,N_244,N_268);
xnor U337 (N_337,N_194,N_260);
nand U338 (N_338,N_281,N_205);
xnor U339 (N_339,N_233,In_486);
and U340 (N_340,N_256,N_239);
nand U341 (N_341,N_135,N_150);
and U342 (N_342,In_127,N_190);
nand U343 (N_343,N_202,N_231);
nand U344 (N_344,N_187,In_373);
and U345 (N_345,N_107,N_262);
or U346 (N_346,In_370,N_131);
and U347 (N_347,N_287,In_227);
nor U348 (N_348,In_468,In_130);
and U349 (N_349,In_354,N_240);
or U350 (N_350,N_288,N_248);
and U351 (N_351,N_85,N_99);
and U352 (N_352,N_266,N_258);
or U353 (N_353,N_235,In_98);
or U354 (N_354,N_295,N_16);
nor U355 (N_355,In_235,N_282);
nand U356 (N_356,N_9,N_154);
nor U357 (N_357,In_261,N_254);
or U358 (N_358,N_120,N_149);
and U359 (N_359,N_298,N_296);
nand U360 (N_360,N_332,N_321);
xor U361 (N_361,N_356,N_192);
and U362 (N_362,N_166,N_355);
nand U363 (N_363,N_247,N_342);
and U364 (N_364,In_328,N_199);
and U365 (N_365,In_270,N_74);
and U366 (N_366,N_323,N_293);
xor U367 (N_367,N_269,N_350);
or U368 (N_368,N_280,N_308);
xor U369 (N_369,N_46,N_56);
and U370 (N_370,N_118,In_432);
or U371 (N_371,In_102,N_230);
or U372 (N_372,In_93,N_359);
or U373 (N_373,N_309,N_272);
xnor U374 (N_374,N_213,N_168);
and U375 (N_375,N_236,In_2);
or U376 (N_376,N_318,In_284);
nor U377 (N_377,N_320,N_346);
nor U378 (N_378,N_80,N_311);
and U379 (N_379,In_109,N_264);
xnor U380 (N_380,In_279,N_273);
nor U381 (N_381,N_226,N_249);
and U382 (N_382,N_124,N_243);
and U383 (N_383,In_466,N_345);
nor U384 (N_384,N_261,N_200);
and U385 (N_385,N_306,N_210);
xor U386 (N_386,N_314,N_316);
or U387 (N_387,In_86,N_330);
nor U388 (N_388,N_134,N_343);
and U389 (N_389,N_225,N_270);
xnor U390 (N_390,In_470,N_319);
nand U391 (N_391,N_344,N_358);
xnor U392 (N_392,N_250,N_305);
xor U393 (N_393,In_218,N_352);
nor U394 (N_394,N_255,N_246);
or U395 (N_395,N_245,N_348);
or U396 (N_396,N_106,N_195);
xor U397 (N_397,N_329,N_335);
nand U398 (N_398,N_196,N_253);
or U399 (N_399,N_337,N_136);
nand U400 (N_400,In_242,N_294);
or U401 (N_401,N_242,N_292);
and U402 (N_402,N_341,N_347);
nand U403 (N_403,N_336,N_310);
or U404 (N_404,N_303,In_150);
and U405 (N_405,In_380,N_339);
nand U406 (N_406,N_326,N_340);
nor U407 (N_407,N_315,N_218);
xnor U408 (N_408,N_301,N_333);
nor U409 (N_409,In_317,N_338);
nand U410 (N_410,N_286,N_322);
nand U411 (N_411,N_312,In_388);
xor U412 (N_412,N_334,N_357);
nand U413 (N_413,N_263,N_285);
and U414 (N_414,In_490,N_354);
nor U415 (N_415,In_3,N_331);
nor U416 (N_416,N_265,N_278);
and U417 (N_417,In_362,N_291);
or U418 (N_418,In_81,N_351);
or U419 (N_419,N_324,N_300);
nand U420 (N_420,N_307,N_376);
nor U421 (N_421,N_228,N_418);
nor U422 (N_422,N_412,N_407);
or U423 (N_423,N_397,N_374);
and U424 (N_424,N_385,N_406);
nor U425 (N_425,N_313,N_390);
and U426 (N_426,N_373,N_362);
nand U427 (N_427,N_393,N_403);
nand U428 (N_428,N_409,In_214);
or U429 (N_429,In_101,N_405);
or U430 (N_430,N_372,N_380);
xor U431 (N_431,N_167,N_349);
nand U432 (N_432,N_384,N_398);
and U433 (N_433,N_416,N_365);
or U434 (N_434,N_382,In_133);
or U435 (N_435,N_387,N_410);
nor U436 (N_436,N_400,N_402);
or U437 (N_437,N_394,N_399);
nor U438 (N_438,N_395,N_20);
nor U439 (N_439,N_377,N_325);
nor U440 (N_440,N_11,N_367);
xnor U441 (N_441,N_396,In_39);
or U442 (N_442,N_361,N_383);
nand U443 (N_443,N_353,N_391);
nor U444 (N_444,N_419,N_328);
nor U445 (N_445,N_369,N_414);
nor U446 (N_446,N_413,In_494);
or U447 (N_447,N_415,N_388);
nor U448 (N_448,N_389,N_392);
xor U449 (N_449,In_428,N_381);
nand U450 (N_450,N_302,N_404);
nand U451 (N_451,N_379,N_368);
xnor U452 (N_452,N_327,N_408);
or U453 (N_453,N_366,N_417);
nor U454 (N_454,N_375,N_370);
or U455 (N_455,N_360,N_411);
xnor U456 (N_456,N_364,N_401);
xor U457 (N_457,N_317,N_386);
or U458 (N_458,N_378,N_363);
xnor U459 (N_459,N_371,N_304);
nor U460 (N_460,N_371,N_392);
xnor U461 (N_461,N_20,N_349);
or U462 (N_462,N_372,N_407);
nor U463 (N_463,N_361,N_409);
nand U464 (N_464,N_228,In_494);
or U465 (N_465,N_381,N_375);
nor U466 (N_466,In_214,N_361);
xnor U467 (N_467,N_361,In_39);
nand U468 (N_468,N_377,N_328);
and U469 (N_469,N_391,N_384);
or U470 (N_470,N_417,N_397);
xnor U471 (N_471,N_386,N_20);
and U472 (N_472,N_369,In_214);
or U473 (N_473,N_402,In_214);
nor U474 (N_474,In_101,N_394);
xnor U475 (N_475,N_362,N_366);
and U476 (N_476,N_307,N_378);
and U477 (N_477,N_391,N_393);
nand U478 (N_478,N_410,N_377);
or U479 (N_479,N_384,N_390);
nand U480 (N_480,N_442,N_458);
and U481 (N_481,N_479,N_463);
and U482 (N_482,N_468,N_466);
xor U483 (N_483,N_447,N_453);
xor U484 (N_484,N_434,N_435);
xor U485 (N_485,N_450,N_448);
nor U486 (N_486,N_444,N_427);
nor U487 (N_487,N_432,N_440);
nor U488 (N_488,N_433,N_422);
nor U489 (N_489,N_428,N_424);
nor U490 (N_490,N_426,N_451);
or U491 (N_491,N_438,N_460);
or U492 (N_492,N_471,N_470);
or U493 (N_493,N_475,N_446);
or U494 (N_494,N_477,N_445);
or U495 (N_495,N_461,N_472);
or U496 (N_496,N_430,N_457);
and U497 (N_497,N_443,N_449);
or U498 (N_498,N_465,N_421);
nand U499 (N_499,N_452,N_476);
or U500 (N_500,N_467,N_420);
nor U501 (N_501,N_423,N_436);
or U502 (N_502,N_459,N_437);
xnor U503 (N_503,N_456,N_441);
or U504 (N_504,N_474,N_478);
nor U505 (N_505,N_431,N_473);
nor U506 (N_506,N_425,N_454);
or U507 (N_507,N_464,N_469);
nor U508 (N_508,N_455,N_439);
nand U509 (N_509,N_462,N_429);
nor U510 (N_510,N_464,N_450);
nor U511 (N_511,N_458,N_456);
or U512 (N_512,N_451,N_469);
or U513 (N_513,N_440,N_471);
or U514 (N_514,N_429,N_473);
nor U515 (N_515,N_478,N_422);
and U516 (N_516,N_478,N_433);
nor U517 (N_517,N_435,N_472);
and U518 (N_518,N_423,N_472);
nand U519 (N_519,N_444,N_467);
or U520 (N_520,N_454,N_444);
nor U521 (N_521,N_474,N_447);
nand U522 (N_522,N_458,N_427);
xnor U523 (N_523,N_433,N_477);
xor U524 (N_524,N_453,N_444);
nand U525 (N_525,N_426,N_456);
or U526 (N_526,N_456,N_445);
nor U527 (N_527,N_446,N_439);
or U528 (N_528,N_433,N_479);
or U529 (N_529,N_423,N_469);
nor U530 (N_530,N_451,N_475);
nand U531 (N_531,N_472,N_449);
nor U532 (N_532,N_429,N_445);
xor U533 (N_533,N_453,N_458);
or U534 (N_534,N_451,N_478);
and U535 (N_535,N_435,N_466);
xor U536 (N_536,N_460,N_463);
and U537 (N_537,N_431,N_468);
nor U538 (N_538,N_440,N_468);
or U539 (N_539,N_446,N_472);
and U540 (N_540,N_535,N_512);
nor U541 (N_541,N_536,N_518);
or U542 (N_542,N_525,N_523);
or U543 (N_543,N_527,N_514);
and U544 (N_544,N_485,N_533);
xnor U545 (N_545,N_494,N_504);
or U546 (N_546,N_537,N_489);
xnor U547 (N_547,N_502,N_531);
nand U548 (N_548,N_491,N_532);
xor U549 (N_549,N_515,N_520);
nand U550 (N_550,N_530,N_522);
and U551 (N_551,N_526,N_480);
nor U552 (N_552,N_488,N_511);
or U553 (N_553,N_509,N_510);
xnor U554 (N_554,N_519,N_507);
and U555 (N_555,N_506,N_539);
nor U556 (N_556,N_490,N_534);
nor U557 (N_557,N_498,N_484);
and U558 (N_558,N_538,N_524);
xnor U559 (N_559,N_501,N_513);
or U560 (N_560,N_517,N_482);
nor U561 (N_561,N_521,N_500);
and U562 (N_562,N_499,N_528);
nor U563 (N_563,N_508,N_496);
nor U564 (N_564,N_497,N_486);
xor U565 (N_565,N_516,N_495);
nor U566 (N_566,N_492,N_529);
xor U567 (N_567,N_493,N_503);
xnor U568 (N_568,N_481,N_505);
nor U569 (N_569,N_487,N_483);
nand U570 (N_570,N_531,N_529);
nor U571 (N_571,N_485,N_483);
xor U572 (N_572,N_523,N_504);
or U573 (N_573,N_520,N_500);
nor U574 (N_574,N_521,N_523);
nor U575 (N_575,N_532,N_507);
xor U576 (N_576,N_481,N_524);
xnor U577 (N_577,N_536,N_528);
or U578 (N_578,N_523,N_508);
nand U579 (N_579,N_502,N_524);
or U580 (N_580,N_510,N_514);
nor U581 (N_581,N_506,N_501);
or U582 (N_582,N_493,N_527);
or U583 (N_583,N_486,N_496);
and U584 (N_584,N_489,N_501);
and U585 (N_585,N_496,N_503);
nand U586 (N_586,N_523,N_481);
xnor U587 (N_587,N_535,N_497);
xor U588 (N_588,N_508,N_491);
or U589 (N_589,N_522,N_520);
xnor U590 (N_590,N_498,N_492);
or U591 (N_591,N_508,N_513);
nor U592 (N_592,N_526,N_524);
xor U593 (N_593,N_526,N_536);
or U594 (N_594,N_522,N_491);
xor U595 (N_595,N_517,N_515);
or U596 (N_596,N_496,N_515);
nand U597 (N_597,N_537,N_505);
and U598 (N_598,N_521,N_522);
nor U599 (N_599,N_480,N_529);
xor U600 (N_600,N_574,N_543);
and U601 (N_601,N_561,N_576);
xnor U602 (N_602,N_579,N_597);
xor U603 (N_603,N_572,N_583);
and U604 (N_604,N_541,N_542);
xnor U605 (N_605,N_556,N_594);
nor U606 (N_606,N_565,N_564);
and U607 (N_607,N_558,N_562);
nand U608 (N_608,N_546,N_550);
nand U609 (N_609,N_578,N_545);
nand U610 (N_610,N_596,N_573);
nor U611 (N_611,N_560,N_595);
or U612 (N_612,N_570,N_575);
nand U613 (N_613,N_587,N_590);
nor U614 (N_614,N_586,N_554);
nand U615 (N_615,N_549,N_568);
and U616 (N_616,N_567,N_592);
xor U617 (N_617,N_577,N_580);
xor U618 (N_618,N_591,N_555);
or U619 (N_619,N_589,N_593);
xnor U620 (N_620,N_566,N_557);
and U621 (N_621,N_548,N_571);
nor U622 (N_622,N_569,N_581);
xor U623 (N_623,N_588,N_552);
and U624 (N_624,N_599,N_584);
xor U625 (N_625,N_585,N_547);
and U626 (N_626,N_598,N_544);
or U627 (N_627,N_551,N_582);
nand U628 (N_628,N_540,N_563);
and U629 (N_629,N_559,N_553);
nor U630 (N_630,N_563,N_570);
nor U631 (N_631,N_559,N_555);
nand U632 (N_632,N_565,N_546);
xnor U633 (N_633,N_590,N_586);
xnor U634 (N_634,N_553,N_572);
nand U635 (N_635,N_580,N_561);
xnor U636 (N_636,N_569,N_566);
xor U637 (N_637,N_593,N_586);
and U638 (N_638,N_553,N_561);
nor U639 (N_639,N_569,N_578);
nand U640 (N_640,N_598,N_561);
nor U641 (N_641,N_542,N_552);
nor U642 (N_642,N_564,N_599);
or U643 (N_643,N_576,N_591);
nand U644 (N_644,N_578,N_567);
and U645 (N_645,N_596,N_545);
or U646 (N_646,N_562,N_589);
or U647 (N_647,N_548,N_567);
xnor U648 (N_648,N_579,N_560);
or U649 (N_649,N_586,N_552);
or U650 (N_650,N_562,N_584);
nor U651 (N_651,N_548,N_590);
and U652 (N_652,N_585,N_573);
xor U653 (N_653,N_541,N_565);
or U654 (N_654,N_599,N_595);
nor U655 (N_655,N_597,N_560);
or U656 (N_656,N_540,N_549);
and U657 (N_657,N_552,N_596);
and U658 (N_658,N_552,N_583);
xor U659 (N_659,N_544,N_572);
or U660 (N_660,N_608,N_656);
and U661 (N_661,N_645,N_640);
nor U662 (N_662,N_639,N_617);
nand U663 (N_663,N_609,N_624);
nand U664 (N_664,N_649,N_653);
nor U665 (N_665,N_657,N_627);
and U666 (N_666,N_619,N_641);
nor U667 (N_667,N_626,N_613);
or U668 (N_668,N_646,N_614);
xor U669 (N_669,N_605,N_632);
nand U670 (N_670,N_637,N_650);
nand U671 (N_671,N_620,N_644);
nor U672 (N_672,N_630,N_603);
or U673 (N_673,N_612,N_621);
or U674 (N_674,N_633,N_602);
nor U675 (N_675,N_607,N_643);
nand U676 (N_676,N_623,N_610);
or U677 (N_677,N_634,N_652);
and U678 (N_678,N_655,N_642);
and U679 (N_679,N_625,N_651);
and U680 (N_680,N_636,N_635);
and U681 (N_681,N_622,N_629);
nor U682 (N_682,N_601,N_647);
and U683 (N_683,N_615,N_631);
nor U684 (N_684,N_638,N_606);
or U685 (N_685,N_600,N_618);
or U686 (N_686,N_616,N_604);
and U687 (N_687,N_628,N_648);
and U688 (N_688,N_658,N_611);
xor U689 (N_689,N_659,N_654);
xnor U690 (N_690,N_649,N_603);
xnor U691 (N_691,N_647,N_605);
nor U692 (N_692,N_653,N_635);
nand U693 (N_693,N_635,N_658);
nand U694 (N_694,N_648,N_618);
nand U695 (N_695,N_608,N_633);
xnor U696 (N_696,N_631,N_659);
or U697 (N_697,N_603,N_652);
xor U698 (N_698,N_638,N_618);
nand U699 (N_699,N_648,N_658);
nor U700 (N_700,N_651,N_623);
xor U701 (N_701,N_636,N_644);
nand U702 (N_702,N_643,N_639);
nor U703 (N_703,N_613,N_642);
or U704 (N_704,N_638,N_614);
xnor U705 (N_705,N_629,N_612);
or U706 (N_706,N_639,N_627);
or U707 (N_707,N_655,N_635);
xor U708 (N_708,N_626,N_611);
nor U709 (N_709,N_641,N_644);
xnor U710 (N_710,N_600,N_616);
or U711 (N_711,N_626,N_620);
nor U712 (N_712,N_612,N_619);
nor U713 (N_713,N_610,N_635);
nor U714 (N_714,N_643,N_653);
and U715 (N_715,N_629,N_624);
and U716 (N_716,N_609,N_641);
or U717 (N_717,N_630,N_600);
and U718 (N_718,N_611,N_642);
or U719 (N_719,N_640,N_650);
nand U720 (N_720,N_691,N_700);
nand U721 (N_721,N_667,N_669);
nand U722 (N_722,N_704,N_676);
xor U723 (N_723,N_692,N_705);
xnor U724 (N_724,N_661,N_680);
nand U725 (N_725,N_682,N_679);
or U726 (N_726,N_703,N_701);
nand U727 (N_727,N_670,N_715);
nand U728 (N_728,N_668,N_697);
and U729 (N_729,N_698,N_674);
and U730 (N_730,N_714,N_689);
and U731 (N_731,N_685,N_686);
and U732 (N_732,N_666,N_681);
nand U733 (N_733,N_707,N_711);
and U734 (N_734,N_665,N_696);
nor U735 (N_735,N_709,N_713);
xnor U736 (N_736,N_675,N_664);
or U737 (N_737,N_719,N_718);
nor U738 (N_738,N_678,N_662);
nor U739 (N_739,N_694,N_710);
and U740 (N_740,N_716,N_673);
nand U741 (N_741,N_663,N_688);
xnor U742 (N_742,N_690,N_706);
xnor U743 (N_743,N_708,N_660);
xnor U744 (N_744,N_702,N_672);
and U745 (N_745,N_693,N_695);
nand U746 (N_746,N_712,N_683);
or U747 (N_747,N_684,N_699);
or U748 (N_748,N_671,N_717);
xnor U749 (N_749,N_687,N_677);
or U750 (N_750,N_664,N_693);
nand U751 (N_751,N_698,N_699);
nand U752 (N_752,N_714,N_705);
or U753 (N_753,N_679,N_688);
and U754 (N_754,N_717,N_714);
and U755 (N_755,N_716,N_669);
and U756 (N_756,N_718,N_682);
nor U757 (N_757,N_670,N_676);
nor U758 (N_758,N_665,N_671);
and U759 (N_759,N_675,N_718);
and U760 (N_760,N_672,N_676);
or U761 (N_761,N_695,N_661);
nor U762 (N_762,N_663,N_682);
and U763 (N_763,N_712,N_711);
nand U764 (N_764,N_690,N_682);
nor U765 (N_765,N_689,N_671);
nor U766 (N_766,N_719,N_705);
nor U767 (N_767,N_708,N_691);
nand U768 (N_768,N_678,N_693);
xnor U769 (N_769,N_679,N_699);
or U770 (N_770,N_663,N_685);
xnor U771 (N_771,N_662,N_692);
nand U772 (N_772,N_661,N_691);
or U773 (N_773,N_713,N_675);
nand U774 (N_774,N_676,N_673);
nand U775 (N_775,N_708,N_664);
or U776 (N_776,N_707,N_687);
or U777 (N_777,N_673,N_712);
and U778 (N_778,N_682,N_660);
and U779 (N_779,N_698,N_671);
xor U780 (N_780,N_724,N_776);
or U781 (N_781,N_768,N_727);
or U782 (N_782,N_754,N_767);
or U783 (N_783,N_752,N_730);
nand U784 (N_784,N_778,N_739);
and U785 (N_785,N_731,N_770);
nor U786 (N_786,N_760,N_745);
or U787 (N_787,N_774,N_726);
nor U788 (N_788,N_775,N_750);
xnor U789 (N_789,N_720,N_741);
and U790 (N_790,N_734,N_744);
or U791 (N_791,N_772,N_766);
nand U792 (N_792,N_757,N_742);
or U793 (N_793,N_723,N_763);
xor U794 (N_794,N_747,N_771);
and U795 (N_795,N_736,N_769);
nor U796 (N_796,N_728,N_761);
and U797 (N_797,N_737,N_779);
nor U798 (N_798,N_722,N_756);
or U799 (N_799,N_733,N_740);
nor U800 (N_800,N_748,N_759);
and U801 (N_801,N_773,N_729);
xnor U802 (N_802,N_721,N_746);
or U803 (N_803,N_735,N_732);
nor U804 (N_804,N_753,N_738);
nor U805 (N_805,N_777,N_762);
or U806 (N_806,N_743,N_725);
or U807 (N_807,N_765,N_749);
or U808 (N_808,N_758,N_751);
and U809 (N_809,N_764,N_755);
xor U810 (N_810,N_776,N_725);
and U811 (N_811,N_767,N_735);
or U812 (N_812,N_769,N_729);
xnor U813 (N_813,N_773,N_768);
or U814 (N_814,N_724,N_763);
xnor U815 (N_815,N_778,N_722);
nor U816 (N_816,N_734,N_743);
nor U817 (N_817,N_776,N_743);
xnor U818 (N_818,N_720,N_776);
nor U819 (N_819,N_723,N_776);
and U820 (N_820,N_738,N_749);
xnor U821 (N_821,N_729,N_744);
xor U822 (N_822,N_724,N_723);
or U823 (N_823,N_720,N_763);
xor U824 (N_824,N_748,N_752);
nor U825 (N_825,N_751,N_768);
nand U826 (N_826,N_741,N_730);
and U827 (N_827,N_750,N_746);
nor U828 (N_828,N_778,N_724);
and U829 (N_829,N_755,N_762);
or U830 (N_830,N_770,N_762);
nand U831 (N_831,N_755,N_730);
xor U832 (N_832,N_746,N_753);
xnor U833 (N_833,N_762,N_764);
nand U834 (N_834,N_726,N_733);
xor U835 (N_835,N_721,N_730);
or U836 (N_836,N_774,N_760);
nand U837 (N_837,N_771,N_745);
nor U838 (N_838,N_750,N_766);
nor U839 (N_839,N_748,N_724);
nand U840 (N_840,N_832,N_809);
nand U841 (N_841,N_839,N_802);
nand U842 (N_842,N_795,N_784);
and U843 (N_843,N_787,N_817);
nand U844 (N_844,N_781,N_805);
xor U845 (N_845,N_797,N_819);
nand U846 (N_846,N_807,N_803);
nor U847 (N_847,N_790,N_782);
nand U848 (N_848,N_792,N_829);
or U849 (N_849,N_831,N_833);
and U850 (N_850,N_806,N_825);
nor U851 (N_851,N_793,N_828);
and U852 (N_852,N_836,N_813);
or U853 (N_853,N_788,N_799);
xor U854 (N_854,N_794,N_835);
xor U855 (N_855,N_834,N_786);
or U856 (N_856,N_811,N_785);
nand U857 (N_857,N_827,N_815);
and U858 (N_858,N_822,N_789);
nand U859 (N_859,N_814,N_821);
and U860 (N_860,N_796,N_816);
and U861 (N_861,N_810,N_798);
nor U862 (N_862,N_830,N_826);
or U863 (N_863,N_823,N_838);
nand U864 (N_864,N_820,N_780);
nor U865 (N_865,N_818,N_800);
xnor U866 (N_866,N_791,N_804);
nor U867 (N_867,N_837,N_783);
and U868 (N_868,N_824,N_812);
nand U869 (N_869,N_808,N_801);
xor U870 (N_870,N_782,N_787);
or U871 (N_871,N_799,N_837);
or U872 (N_872,N_834,N_805);
xnor U873 (N_873,N_790,N_820);
nand U874 (N_874,N_784,N_813);
or U875 (N_875,N_834,N_800);
nand U876 (N_876,N_834,N_814);
nor U877 (N_877,N_831,N_808);
xor U878 (N_878,N_830,N_823);
or U879 (N_879,N_831,N_799);
nor U880 (N_880,N_825,N_805);
or U881 (N_881,N_780,N_810);
nand U882 (N_882,N_835,N_781);
nand U883 (N_883,N_795,N_827);
nand U884 (N_884,N_827,N_787);
nand U885 (N_885,N_838,N_839);
and U886 (N_886,N_815,N_817);
xor U887 (N_887,N_834,N_781);
xor U888 (N_888,N_813,N_823);
and U889 (N_889,N_801,N_832);
xnor U890 (N_890,N_810,N_791);
nand U891 (N_891,N_822,N_812);
xnor U892 (N_892,N_801,N_797);
nor U893 (N_893,N_838,N_828);
and U894 (N_894,N_794,N_837);
nand U895 (N_895,N_812,N_819);
and U896 (N_896,N_823,N_810);
nand U897 (N_897,N_802,N_825);
nand U898 (N_898,N_822,N_830);
or U899 (N_899,N_833,N_784);
xnor U900 (N_900,N_892,N_847);
and U901 (N_901,N_859,N_861);
nand U902 (N_902,N_889,N_856);
and U903 (N_903,N_897,N_884);
nand U904 (N_904,N_875,N_850);
and U905 (N_905,N_868,N_881);
nor U906 (N_906,N_873,N_852);
and U907 (N_907,N_854,N_853);
nor U908 (N_908,N_894,N_891);
and U909 (N_909,N_893,N_872);
nand U910 (N_910,N_883,N_858);
and U911 (N_911,N_899,N_878);
and U912 (N_912,N_879,N_867);
xor U913 (N_913,N_896,N_885);
nor U914 (N_914,N_877,N_874);
nor U915 (N_915,N_841,N_886);
and U916 (N_916,N_876,N_844);
and U917 (N_917,N_869,N_880);
nor U918 (N_918,N_845,N_864);
nand U919 (N_919,N_857,N_851);
nand U920 (N_920,N_860,N_842);
xnor U921 (N_921,N_862,N_840);
and U922 (N_922,N_870,N_849);
or U923 (N_923,N_846,N_843);
or U924 (N_924,N_871,N_848);
nor U925 (N_925,N_866,N_855);
or U926 (N_926,N_887,N_882);
nand U927 (N_927,N_890,N_865);
xnor U928 (N_928,N_898,N_895);
xnor U929 (N_929,N_888,N_863);
nor U930 (N_930,N_878,N_867);
and U931 (N_931,N_843,N_895);
and U932 (N_932,N_899,N_880);
nand U933 (N_933,N_865,N_847);
and U934 (N_934,N_874,N_896);
xnor U935 (N_935,N_849,N_883);
or U936 (N_936,N_845,N_879);
nor U937 (N_937,N_846,N_883);
nor U938 (N_938,N_865,N_889);
and U939 (N_939,N_870,N_888);
xor U940 (N_940,N_880,N_860);
xor U941 (N_941,N_845,N_856);
and U942 (N_942,N_884,N_895);
and U943 (N_943,N_843,N_870);
or U944 (N_944,N_845,N_849);
or U945 (N_945,N_878,N_879);
xor U946 (N_946,N_857,N_864);
xnor U947 (N_947,N_857,N_888);
and U948 (N_948,N_885,N_871);
xor U949 (N_949,N_860,N_894);
and U950 (N_950,N_845,N_893);
or U951 (N_951,N_849,N_858);
and U952 (N_952,N_845,N_866);
xnor U953 (N_953,N_843,N_865);
nand U954 (N_954,N_876,N_888);
and U955 (N_955,N_890,N_891);
xnor U956 (N_956,N_854,N_843);
or U957 (N_957,N_899,N_854);
nor U958 (N_958,N_843,N_879);
or U959 (N_959,N_848,N_887);
or U960 (N_960,N_947,N_946);
nand U961 (N_961,N_911,N_937);
nor U962 (N_962,N_933,N_901);
and U963 (N_963,N_950,N_922);
and U964 (N_964,N_913,N_917);
and U965 (N_965,N_919,N_957);
nor U966 (N_966,N_909,N_932);
nor U967 (N_967,N_959,N_910);
xor U968 (N_968,N_943,N_948);
xnor U969 (N_969,N_921,N_914);
nor U970 (N_970,N_927,N_925);
and U971 (N_971,N_928,N_916);
nand U972 (N_972,N_938,N_958);
and U973 (N_973,N_915,N_912);
xnor U974 (N_974,N_952,N_942);
nand U975 (N_975,N_934,N_904);
xor U976 (N_976,N_931,N_944);
or U977 (N_977,N_926,N_918);
and U978 (N_978,N_955,N_953);
xor U979 (N_979,N_908,N_907);
xnor U980 (N_980,N_940,N_949);
xnor U981 (N_981,N_951,N_936);
or U982 (N_982,N_903,N_935);
and U983 (N_983,N_906,N_902);
xnor U984 (N_984,N_954,N_920);
xnor U985 (N_985,N_923,N_939);
or U986 (N_986,N_900,N_905);
nand U987 (N_987,N_930,N_941);
xnor U988 (N_988,N_929,N_924);
and U989 (N_989,N_956,N_945);
nand U990 (N_990,N_906,N_912);
nand U991 (N_991,N_930,N_937);
or U992 (N_992,N_957,N_955);
and U993 (N_993,N_911,N_913);
xnor U994 (N_994,N_907,N_953);
xnor U995 (N_995,N_958,N_953);
xor U996 (N_996,N_909,N_902);
nor U997 (N_997,N_905,N_947);
nor U998 (N_998,N_913,N_954);
and U999 (N_999,N_925,N_922);
or U1000 (N_1000,N_909,N_937);
or U1001 (N_1001,N_931,N_920);
nor U1002 (N_1002,N_940,N_921);
nand U1003 (N_1003,N_905,N_913);
nand U1004 (N_1004,N_948,N_910);
nor U1005 (N_1005,N_907,N_943);
nor U1006 (N_1006,N_923,N_903);
and U1007 (N_1007,N_923,N_906);
nand U1008 (N_1008,N_941,N_955);
and U1009 (N_1009,N_902,N_914);
and U1010 (N_1010,N_914,N_918);
or U1011 (N_1011,N_939,N_953);
nand U1012 (N_1012,N_956,N_926);
or U1013 (N_1013,N_945,N_921);
nor U1014 (N_1014,N_905,N_929);
nor U1015 (N_1015,N_924,N_936);
or U1016 (N_1016,N_903,N_910);
nand U1017 (N_1017,N_917,N_951);
or U1018 (N_1018,N_918,N_959);
or U1019 (N_1019,N_956,N_930);
nor U1020 (N_1020,N_1009,N_990);
nand U1021 (N_1021,N_998,N_960);
or U1022 (N_1022,N_1008,N_965);
nor U1023 (N_1023,N_974,N_961);
nand U1024 (N_1024,N_1000,N_999);
and U1025 (N_1025,N_1004,N_1006);
nand U1026 (N_1026,N_968,N_979);
xnor U1027 (N_1027,N_972,N_1002);
or U1028 (N_1028,N_982,N_1014);
nor U1029 (N_1029,N_975,N_1010);
or U1030 (N_1030,N_973,N_976);
nand U1031 (N_1031,N_1019,N_1005);
nand U1032 (N_1032,N_1012,N_1015);
nor U1033 (N_1033,N_971,N_970);
nor U1034 (N_1034,N_1001,N_994);
and U1035 (N_1035,N_997,N_986);
and U1036 (N_1036,N_993,N_964);
nand U1037 (N_1037,N_969,N_995);
and U1038 (N_1038,N_1003,N_988);
nand U1039 (N_1039,N_1016,N_991);
and U1040 (N_1040,N_987,N_1018);
or U1041 (N_1041,N_985,N_1017);
or U1042 (N_1042,N_983,N_992);
nand U1043 (N_1043,N_984,N_977);
nand U1044 (N_1044,N_1013,N_996);
nor U1045 (N_1045,N_981,N_967);
nor U1046 (N_1046,N_1007,N_962);
nand U1047 (N_1047,N_989,N_966);
and U1048 (N_1048,N_963,N_978);
nor U1049 (N_1049,N_980,N_1011);
nand U1050 (N_1050,N_964,N_1009);
nand U1051 (N_1051,N_973,N_972);
nand U1052 (N_1052,N_1011,N_1010);
nor U1053 (N_1053,N_1005,N_972);
nor U1054 (N_1054,N_996,N_963);
nor U1055 (N_1055,N_1013,N_972);
and U1056 (N_1056,N_994,N_1007);
nand U1057 (N_1057,N_997,N_1009);
nor U1058 (N_1058,N_980,N_1006);
nand U1059 (N_1059,N_1005,N_995);
and U1060 (N_1060,N_1003,N_1013);
xnor U1061 (N_1061,N_984,N_980);
or U1062 (N_1062,N_972,N_967);
xor U1063 (N_1063,N_969,N_962);
nand U1064 (N_1064,N_1002,N_998);
xor U1065 (N_1065,N_983,N_991);
nor U1066 (N_1066,N_965,N_963);
and U1067 (N_1067,N_997,N_1007);
and U1068 (N_1068,N_1000,N_994);
xor U1069 (N_1069,N_963,N_987);
nor U1070 (N_1070,N_988,N_1005);
nor U1071 (N_1071,N_987,N_1008);
nand U1072 (N_1072,N_1016,N_967);
nand U1073 (N_1073,N_963,N_974);
nand U1074 (N_1074,N_969,N_986);
xnor U1075 (N_1075,N_965,N_973);
nand U1076 (N_1076,N_995,N_984);
or U1077 (N_1077,N_994,N_969);
and U1078 (N_1078,N_1013,N_1000);
or U1079 (N_1079,N_998,N_966);
xor U1080 (N_1080,N_1027,N_1020);
and U1081 (N_1081,N_1034,N_1025);
xnor U1082 (N_1082,N_1058,N_1066);
or U1083 (N_1083,N_1026,N_1077);
nor U1084 (N_1084,N_1071,N_1022);
and U1085 (N_1085,N_1048,N_1035);
or U1086 (N_1086,N_1021,N_1042);
or U1087 (N_1087,N_1040,N_1045);
nand U1088 (N_1088,N_1049,N_1073);
and U1089 (N_1089,N_1052,N_1078);
and U1090 (N_1090,N_1051,N_1050);
xnor U1091 (N_1091,N_1068,N_1028);
nand U1092 (N_1092,N_1039,N_1074);
nand U1093 (N_1093,N_1079,N_1056);
or U1094 (N_1094,N_1044,N_1057);
nand U1095 (N_1095,N_1043,N_1053);
nand U1096 (N_1096,N_1064,N_1070);
and U1097 (N_1097,N_1067,N_1024);
xor U1098 (N_1098,N_1030,N_1075);
and U1099 (N_1099,N_1072,N_1038);
nor U1100 (N_1100,N_1059,N_1055);
or U1101 (N_1101,N_1046,N_1032);
nand U1102 (N_1102,N_1033,N_1069);
nand U1103 (N_1103,N_1076,N_1061);
nor U1104 (N_1104,N_1047,N_1063);
xnor U1105 (N_1105,N_1054,N_1037);
nand U1106 (N_1106,N_1065,N_1031);
nor U1107 (N_1107,N_1023,N_1036);
nand U1108 (N_1108,N_1062,N_1029);
or U1109 (N_1109,N_1041,N_1060);
or U1110 (N_1110,N_1049,N_1041);
and U1111 (N_1111,N_1049,N_1062);
or U1112 (N_1112,N_1068,N_1064);
and U1113 (N_1113,N_1070,N_1078);
nand U1114 (N_1114,N_1055,N_1038);
nand U1115 (N_1115,N_1065,N_1073);
and U1116 (N_1116,N_1021,N_1030);
xor U1117 (N_1117,N_1023,N_1031);
or U1118 (N_1118,N_1078,N_1028);
and U1119 (N_1119,N_1022,N_1044);
xor U1120 (N_1120,N_1064,N_1020);
nor U1121 (N_1121,N_1078,N_1056);
or U1122 (N_1122,N_1042,N_1074);
nand U1123 (N_1123,N_1040,N_1033);
or U1124 (N_1124,N_1056,N_1031);
or U1125 (N_1125,N_1057,N_1067);
nor U1126 (N_1126,N_1045,N_1069);
and U1127 (N_1127,N_1039,N_1027);
nor U1128 (N_1128,N_1030,N_1036);
xor U1129 (N_1129,N_1028,N_1020);
xor U1130 (N_1130,N_1059,N_1021);
nor U1131 (N_1131,N_1053,N_1036);
and U1132 (N_1132,N_1042,N_1071);
nor U1133 (N_1133,N_1046,N_1066);
xnor U1134 (N_1134,N_1029,N_1021);
or U1135 (N_1135,N_1075,N_1057);
nor U1136 (N_1136,N_1078,N_1059);
nand U1137 (N_1137,N_1022,N_1068);
nor U1138 (N_1138,N_1053,N_1078);
and U1139 (N_1139,N_1068,N_1034);
nand U1140 (N_1140,N_1088,N_1100);
nor U1141 (N_1141,N_1082,N_1136);
xor U1142 (N_1142,N_1095,N_1133);
nor U1143 (N_1143,N_1125,N_1121);
nand U1144 (N_1144,N_1104,N_1092);
xor U1145 (N_1145,N_1090,N_1138);
nor U1146 (N_1146,N_1120,N_1084);
or U1147 (N_1147,N_1099,N_1106);
xor U1148 (N_1148,N_1123,N_1114);
or U1149 (N_1149,N_1127,N_1096);
nand U1150 (N_1150,N_1081,N_1134);
or U1151 (N_1151,N_1112,N_1139);
xnor U1152 (N_1152,N_1102,N_1137);
and U1153 (N_1153,N_1115,N_1131);
and U1154 (N_1154,N_1091,N_1108);
nor U1155 (N_1155,N_1124,N_1094);
nand U1156 (N_1156,N_1126,N_1111);
nor U1157 (N_1157,N_1101,N_1097);
or U1158 (N_1158,N_1083,N_1122);
xor U1159 (N_1159,N_1098,N_1110);
or U1160 (N_1160,N_1080,N_1103);
xor U1161 (N_1161,N_1105,N_1107);
or U1162 (N_1162,N_1118,N_1086);
or U1163 (N_1163,N_1085,N_1089);
or U1164 (N_1164,N_1087,N_1119);
or U1165 (N_1165,N_1116,N_1093);
nand U1166 (N_1166,N_1130,N_1128);
xor U1167 (N_1167,N_1132,N_1113);
and U1168 (N_1168,N_1109,N_1129);
xnor U1169 (N_1169,N_1117,N_1135);
nand U1170 (N_1170,N_1114,N_1091);
nand U1171 (N_1171,N_1112,N_1130);
xor U1172 (N_1172,N_1124,N_1110);
nor U1173 (N_1173,N_1101,N_1083);
or U1174 (N_1174,N_1101,N_1117);
nand U1175 (N_1175,N_1085,N_1086);
and U1176 (N_1176,N_1131,N_1092);
nor U1177 (N_1177,N_1132,N_1099);
and U1178 (N_1178,N_1123,N_1118);
or U1179 (N_1179,N_1100,N_1105);
nor U1180 (N_1180,N_1117,N_1136);
nand U1181 (N_1181,N_1139,N_1095);
nor U1182 (N_1182,N_1109,N_1104);
nor U1183 (N_1183,N_1124,N_1129);
nand U1184 (N_1184,N_1096,N_1103);
nor U1185 (N_1185,N_1139,N_1108);
nand U1186 (N_1186,N_1129,N_1107);
or U1187 (N_1187,N_1124,N_1125);
or U1188 (N_1188,N_1122,N_1134);
nor U1189 (N_1189,N_1106,N_1110);
nand U1190 (N_1190,N_1127,N_1113);
and U1191 (N_1191,N_1131,N_1139);
nor U1192 (N_1192,N_1081,N_1082);
or U1193 (N_1193,N_1134,N_1111);
or U1194 (N_1194,N_1103,N_1118);
xnor U1195 (N_1195,N_1122,N_1136);
xor U1196 (N_1196,N_1119,N_1109);
or U1197 (N_1197,N_1120,N_1093);
xnor U1198 (N_1198,N_1087,N_1129);
or U1199 (N_1199,N_1084,N_1128);
xor U1200 (N_1200,N_1164,N_1178);
or U1201 (N_1201,N_1186,N_1155);
xnor U1202 (N_1202,N_1190,N_1191);
nand U1203 (N_1203,N_1159,N_1193);
xor U1204 (N_1204,N_1167,N_1196);
xnor U1205 (N_1205,N_1189,N_1199);
xor U1206 (N_1206,N_1175,N_1162);
nor U1207 (N_1207,N_1185,N_1140);
nand U1208 (N_1208,N_1165,N_1147);
xnor U1209 (N_1209,N_1195,N_1176);
nand U1210 (N_1210,N_1143,N_1157);
xor U1211 (N_1211,N_1156,N_1198);
nand U1212 (N_1212,N_1197,N_1188);
or U1213 (N_1213,N_1182,N_1171);
nor U1214 (N_1214,N_1174,N_1181);
nand U1215 (N_1215,N_1149,N_1154);
nand U1216 (N_1216,N_1179,N_1184);
nor U1217 (N_1217,N_1144,N_1148);
xor U1218 (N_1218,N_1180,N_1151);
xor U1219 (N_1219,N_1192,N_1153);
xnor U1220 (N_1220,N_1141,N_1194);
or U1221 (N_1221,N_1160,N_1173);
nand U1222 (N_1222,N_1169,N_1142);
and U1223 (N_1223,N_1168,N_1177);
and U1224 (N_1224,N_1187,N_1170);
and U1225 (N_1225,N_1163,N_1150);
and U1226 (N_1226,N_1158,N_1161);
xnor U1227 (N_1227,N_1183,N_1172);
nand U1228 (N_1228,N_1152,N_1146);
xnor U1229 (N_1229,N_1166,N_1145);
and U1230 (N_1230,N_1183,N_1194);
nor U1231 (N_1231,N_1164,N_1149);
xor U1232 (N_1232,N_1166,N_1156);
nor U1233 (N_1233,N_1181,N_1180);
or U1234 (N_1234,N_1167,N_1157);
xor U1235 (N_1235,N_1198,N_1166);
xnor U1236 (N_1236,N_1184,N_1166);
nor U1237 (N_1237,N_1176,N_1197);
xor U1238 (N_1238,N_1195,N_1144);
or U1239 (N_1239,N_1145,N_1154);
nor U1240 (N_1240,N_1197,N_1141);
nand U1241 (N_1241,N_1185,N_1156);
nor U1242 (N_1242,N_1194,N_1145);
nor U1243 (N_1243,N_1197,N_1191);
and U1244 (N_1244,N_1191,N_1170);
nand U1245 (N_1245,N_1150,N_1187);
or U1246 (N_1246,N_1140,N_1153);
and U1247 (N_1247,N_1147,N_1194);
and U1248 (N_1248,N_1149,N_1170);
xor U1249 (N_1249,N_1161,N_1195);
and U1250 (N_1250,N_1189,N_1190);
or U1251 (N_1251,N_1176,N_1163);
xnor U1252 (N_1252,N_1188,N_1171);
nor U1253 (N_1253,N_1168,N_1141);
and U1254 (N_1254,N_1144,N_1153);
and U1255 (N_1255,N_1149,N_1193);
nor U1256 (N_1256,N_1183,N_1179);
nor U1257 (N_1257,N_1155,N_1187);
nand U1258 (N_1258,N_1144,N_1178);
and U1259 (N_1259,N_1180,N_1185);
or U1260 (N_1260,N_1203,N_1230);
and U1261 (N_1261,N_1257,N_1224);
or U1262 (N_1262,N_1207,N_1214);
xor U1263 (N_1263,N_1204,N_1200);
nor U1264 (N_1264,N_1222,N_1237);
xnor U1265 (N_1265,N_1223,N_1227);
and U1266 (N_1266,N_1259,N_1221);
and U1267 (N_1267,N_1218,N_1246);
xor U1268 (N_1268,N_1220,N_1210);
or U1269 (N_1269,N_1256,N_1209);
or U1270 (N_1270,N_1253,N_1229);
or U1271 (N_1271,N_1235,N_1211);
nor U1272 (N_1272,N_1250,N_1201);
and U1273 (N_1273,N_1244,N_1239);
xor U1274 (N_1274,N_1242,N_1258);
nor U1275 (N_1275,N_1254,N_1251);
nor U1276 (N_1276,N_1238,N_1217);
or U1277 (N_1277,N_1213,N_1245);
and U1278 (N_1278,N_1219,N_1255);
nand U1279 (N_1279,N_1248,N_1247);
nand U1280 (N_1280,N_1212,N_1252);
and U1281 (N_1281,N_1240,N_1231);
and U1282 (N_1282,N_1243,N_1233);
nor U1283 (N_1283,N_1228,N_1208);
nand U1284 (N_1284,N_1215,N_1234);
xor U1285 (N_1285,N_1202,N_1241);
nor U1286 (N_1286,N_1216,N_1225);
nand U1287 (N_1287,N_1206,N_1226);
or U1288 (N_1288,N_1249,N_1232);
xor U1289 (N_1289,N_1236,N_1205);
xnor U1290 (N_1290,N_1248,N_1246);
xor U1291 (N_1291,N_1226,N_1208);
or U1292 (N_1292,N_1200,N_1246);
or U1293 (N_1293,N_1233,N_1216);
nand U1294 (N_1294,N_1211,N_1250);
and U1295 (N_1295,N_1224,N_1250);
or U1296 (N_1296,N_1249,N_1211);
or U1297 (N_1297,N_1219,N_1237);
nand U1298 (N_1298,N_1253,N_1242);
nand U1299 (N_1299,N_1209,N_1217);
or U1300 (N_1300,N_1202,N_1256);
or U1301 (N_1301,N_1257,N_1245);
nor U1302 (N_1302,N_1225,N_1228);
xor U1303 (N_1303,N_1256,N_1253);
or U1304 (N_1304,N_1242,N_1244);
or U1305 (N_1305,N_1248,N_1237);
xor U1306 (N_1306,N_1214,N_1256);
xnor U1307 (N_1307,N_1256,N_1245);
nand U1308 (N_1308,N_1231,N_1224);
or U1309 (N_1309,N_1206,N_1253);
and U1310 (N_1310,N_1222,N_1258);
xnor U1311 (N_1311,N_1216,N_1220);
nor U1312 (N_1312,N_1251,N_1225);
or U1313 (N_1313,N_1259,N_1230);
and U1314 (N_1314,N_1232,N_1256);
or U1315 (N_1315,N_1246,N_1237);
or U1316 (N_1316,N_1225,N_1204);
nor U1317 (N_1317,N_1227,N_1234);
nand U1318 (N_1318,N_1250,N_1244);
xnor U1319 (N_1319,N_1216,N_1244);
nor U1320 (N_1320,N_1307,N_1312);
nand U1321 (N_1321,N_1265,N_1303);
nor U1322 (N_1322,N_1272,N_1314);
and U1323 (N_1323,N_1295,N_1308);
nor U1324 (N_1324,N_1285,N_1302);
nor U1325 (N_1325,N_1317,N_1266);
xnor U1326 (N_1326,N_1305,N_1309);
and U1327 (N_1327,N_1316,N_1279);
xor U1328 (N_1328,N_1293,N_1304);
and U1329 (N_1329,N_1289,N_1275);
and U1330 (N_1330,N_1297,N_1271);
xnor U1331 (N_1331,N_1313,N_1260);
xnor U1332 (N_1332,N_1310,N_1263);
nand U1333 (N_1333,N_1291,N_1276);
xnor U1334 (N_1334,N_1286,N_1283);
and U1335 (N_1335,N_1315,N_1298);
or U1336 (N_1336,N_1287,N_1290);
xor U1337 (N_1337,N_1301,N_1268);
xnor U1338 (N_1338,N_1306,N_1296);
xor U1339 (N_1339,N_1288,N_1278);
nor U1340 (N_1340,N_1294,N_1282);
and U1341 (N_1341,N_1270,N_1318);
and U1342 (N_1342,N_1267,N_1299);
nand U1343 (N_1343,N_1273,N_1319);
nand U1344 (N_1344,N_1264,N_1274);
nor U1345 (N_1345,N_1261,N_1281);
or U1346 (N_1346,N_1280,N_1269);
nor U1347 (N_1347,N_1300,N_1284);
xnor U1348 (N_1348,N_1311,N_1277);
and U1349 (N_1349,N_1262,N_1292);
and U1350 (N_1350,N_1278,N_1267);
and U1351 (N_1351,N_1286,N_1305);
or U1352 (N_1352,N_1304,N_1270);
and U1353 (N_1353,N_1300,N_1261);
or U1354 (N_1354,N_1307,N_1281);
xor U1355 (N_1355,N_1289,N_1311);
xnor U1356 (N_1356,N_1294,N_1291);
xnor U1357 (N_1357,N_1309,N_1292);
and U1358 (N_1358,N_1286,N_1268);
xor U1359 (N_1359,N_1314,N_1303);
or U1360 (N_1360,N_1303,N_1264);
xor U1361 (N_1361,N_1273,N_1260);
xnor U1362 (N_1362,N_1299,N_1280);
nor U1363 (N_1363,N_1313,N_1312);
xnor U1364 (N_1364,N_1268,N_1264);
nor U1365 (N_1365,N_1272,N_1276);
or U1366 (N_1366,N_1262,N_1269);
and U1367 (N_1367,N_1305,N_1260);
xnor U1368 (N_1368,N_1264,N_1301);
nand U1369 (N_1369,N_1269,N_1292);
or U1370 (N_1370,N_1306,N_1267);
or U1371 (N_1371,N_1271,N_1314);
nor U1372 (N_1372,N_1280,N_1297);
and U1373 (N_1373,N_1277,N_1271);
xnor U1374 (N_1374,N_1292,N_1277);
xnor U1375 (N_1375,N_1310,N_1268);
and U1376 (N_1376,N_1262,N_1313);
and U1377 (N_1377,N_1293,N_1294);
and U1378 (N_1378,N_1260,N_1280);
nor U1379 (N_1379,N_1300,N_1305);
xnor U1380 (N_1380,N_1370,N_1371);
or U1381 (N_1381,N_1375,N_1352);
xnor U1382 (N_1382,N_1368,N_1341);
or U1383 (N_1383,N_1351,N_1323);
nand U1384 (N_1384,N_1337,N_1364);
or U1385 (N_1385,N_1344,N_1355);
nand U1386 (N_1386,N_1357,N_1354);
or U1387 (N_1387,N_1353,N_1378);
or U1388 (N_1388,N_1333,N_1359);
or U1389 (N_1389,N_1324,N_1374);
nand U1390 (N_1390,N_1346,N_1342);
or U1391 (N_1391,N_1369,N_1325);
or U1392 (N_1392,N_1328,N_1360);
nand U1393 (N_1393,N_1358,N_1361);
nand U1394 (N_1394,N_1347,N_1321);
xnor U1395 (N_1395,N_1334,N_1362);
and U1396 (N_1396,N_1356,N_1339);
or U1397 (N_1397,N_1329,N_1326);
and U1398 (N_1398,N_1373,N_1336);
or U1399 (N_1399,N_1332,N_1330);
nor U1400 (N_1400,N_1322,N_1379);
and U1401 (N_1401,N_1320,N_1350);
or U1402 (N_1402,N_1376,N_1348);
nand U1403 (N_1403,N_1349,N_1377);
and U1404 (N_1404,N_1345,N_1343);
nor U1405 (N_1405,N_1365,N_1335);
or U1406 (N_1406,N_1327,N_1340);
nor U1407 (N_1407,N_1363,N_1331);
or U1408 (N_1408,N_1338,N_1366);
xor U1409 (N_1409,N_1372,N_1367);
nand U1410 (N_1410,N_1333,N_1371);
nand U1411 (N_1411,N_1344,N_1336);
nor U1412 (N_1412,N_1322,N_1324);
xor U1413 (N_1413,N_1366,N_1369);
or U1414 (N_1414,N_1374,N_1356);
xnor U1415 (N_1415,N_1324,N_1363);
nand U1416 (N_1416,N_1366,N_1339);
or U1417 (N_1417,N_1375,N_1350);
or U1418 (N_1418,N_1339,N_1350);
nor U1419 (N_1419,N_1325,N_1375);
nor U1420 (N_1420,N_1342,N_1323);
or U1421 (N_1421,N_1320,N_1349);
nor U1422 (N_1422,N_1340,N_1366);
nor U1423 (N_1423,N_1359,N_1379);
and U1424 (N_1424,N_1328,N_1359);
nor U1425 (N_1425,N_1327,N_1349);
xor U1426 (N_1426,N_1365,N_1353);
nor U1427 (N_1427,N_1347,N_1371);
xnor U1428 (N_1428,N_1343,N_1373);
xnor U1429 (N_1429,N_1356,N_1366);
and U1430 (N_1430,N_1370,N_1335);
nand U1431 (N_1431,N_1344,N_1364);
nand U1432 (N_1432,N_1351,N_1335);
xor U1433 (N_1433,N_1372,N_1359);
or U1434 (N_1434,N_1335,N_1356);
and U1435 (N_1435,N_1331,N_1346);
nand U1436 (N_1436,N_1341,N_1365);
nor U1437 (N_1437,N_1355,N_1341);
xor U1438 (N_1438,N_1341,N_1346);
nor U1439 (N_1439,N_1326,N_1337);
xor U1440 (N_1440,N_1396,N_1434);
xor U1441 (N_1441,N_1404,N_1432);
or U1442 (N_1442,N_1394,N_1390);
or U1443 (N_1443,N_1438,N_1393);
nor U1444 (N_1444,N_1397,N_1387);
nand U1445 (N_1445,N_1423,N_1392);
xnor U1446 (N_1446,N_1398,N_1403);
and U1447 (N_1447,N_1406,N_1410);
xor U1448 (N_1448,N_1413,N_1388);
nor U1449 (N_1449,N_1384,N_1389);
or U1450 (N_1450,N_1437,N_1382);
nor U1451 (N_1451,N_1391,N_1422);
and U1452 (N_1452,N_1431,N_1418);
xor U1453 (N_1453,N_1417,N_1420);
or U1454 (N_1454,N_1428,N_1405);
nand U1455 (N_1455,N_1429,N_1385);
nor U1456 (N_1456,N_1407,N_1430);
or U1457 (N_1457,N_1425,N_1419);
nor U1458 (N_1458,N_1383,N_1415);
nor U1459 (N_1459,N_1409,N_1439);
xnor U1460 (N_1460,N_1400,N_1426);
nand U1461 (N_1461,N_1435,N_1411);
nor U1462 (N_1462,N_1433,N_1380);
or U1463 (N_1463,N_1395,N_1386);
xnor U1464 (N_1464,N_1427,N_1421);
and U1465 (N_1465,N_1402,N_1414);
or U1466 (N_1466,N_1412,N_1424);
or U1467 (N_1467,N_1436,N_1381);
xnor U1468 (N_1468,N_1408,N_1399);
and U1469 (N_1469,N_1401,N_1416);
nand U1470 (N_1470,N_1394,N_1399);
or U1471 (N_1471,N_1432,N_1394);
nor U1472 (N_1472,N_1411,N_1384);
or U1473 (N_1473,N_1395,N_1431);
nand U1474 (N_1474,N_1382,N_1414);
nand U1475 (N_1475,N_1417,N_1387);
or U1476 (N_1476,N_1435,N_1422);
nand U1477 (N_1477,N_1410,N_1400);
xnor U1478 (N_1478,N_1408,N_1423);
or U1479 (N_1479,N_1406,N_1396);
xnor U1480 (N_1480,N_1399,N_1406);
nor U1481 (N_1481,N_1428,N_1382);
and U1482 (N_1482,N_1431,N_1405);
nand U1483 (N_1483,N_1418,N_1386);
xnor U1484 (N_1484,N_1417,N_1424);
or U1485 (N_1485,N_1437,N_1399);
nor U1486 (N_1486,N_1404,N_1394);
nand U1487 (N_1487,N_1416,N_1437);
xor U1488 (N_1488,N_1414,N_1394);
and U1489 (N_1489,N_1384,N_1406);
xnor U1490 (N_1490,N_1429,N_1436);
and U1491 (N_1491,N_1406,N_1402);
or U1492 (N_1492,N_1410,N_1384);
xnor U1493 (N_1493,N_1406,N_1411);
or U1494 (N_1494,N_1405,N_1435);
xnor U1495 (N_1495,N_1409,N_1398);
xnor U1496 (N_1496,N_1385,N_1383);
and U1497 (N_1497,N_1402,N_1391);
nor U1498 (N_1498,N_1404,N_1417);
nor U1499 (N_1499,N_1387,N_1433);
nor U1500 (N_1500,N_1470,N_1457);
nor U1501 (N_1501,N_1496,N_1450);
nand U1502 (N_1502,N_1488,N_1494);
nand U1503 (N_1503,N_1448,N_1486);
nand U1504 (N_1504,N_1487,N_1499);
xnor U1505 (N_1505,N_1485,N_1445);
xor U1506 (N_1506,N_1493,N_1472);
xnor U1507 (N_1507,N_1443,N_1462);
nor U1508 (N_1508,N_1464,N_1449);
or U1509 (N_1509,N_1495,N_1492);
nor U1510 (N_1510,N_1453,N_1482);
nand U1511 (N_1511,N_1459,N_1468);
and U1512 (N_1512,N_1478,N_1491);
nor U1513 (N_1513,N_1498,N_1483);
or U1514 (N_1514,N_1460,N_1471);
xnor U1515 (N_1515,N_1466,N_1440);
nand U1516 (N_1516,N_1481,N_1469);
and U1517 (N_1517,N_1444,N_1484);
xor U1518 (N_1518,N_1458,N_1473);
nand U1519 (N_1519,N_1476,N_1451);
or U1520 (N_1520,N_1497,N_1467);
nor U1521 (N_1521,N_1465,N_1463);
or U1522 (N_1522,N_1480,N_1490);
nand U1523 (N_1523,N_1442,N_1479);
nor U1524 (N_1524,N_1441,N_1455);
nand U1525 (N_1525,N_1475,N_1456);
nor U1526 (N_1526,N_1446,N_1489);
nand U1527 (N_1527,N_1461,N_1477);
nor U1528 (N_1528,N_1474,N_1452);
nand U1529 (N_1529,N_1447,N_1454);
or U1530 (N_1530,N_1441,N_1442);
and U1531 (N_1531,N_1462,N_1473);
nor U1532 (N_1532,N_1497,N_1493);
xnor U1533 (N_1533,N_1456,N_1487);
and U1534 (N_1534,N_1493,N_1484);
nor U1535 (N_1535,N_1466,N_1446);
nor U1536 (N_1536,N_1443,N_1498);
nand U1537 (N_1537,N_1498,N_1470);
xor U1538 (N_1538,N_1452,N_1449);
nor U1539 (N_1539,N_1482,N_1457);
nand U1540 (N_1540,N_1454,N_1459);
xnor U1541 (N_1541,N_1495,N_1463);
nand U1542 (N_1542,N_1454,N_1464);
xor U1543 (N_1543,N_1463,N_1492);
or U1544 (N_1544,N_1475,N_1477);
nor U1545 (N_1545,N_1440,N_1492);
or U1546 (N_1546,N_1454,N_1469);
or U1547 (N_1547,N_1496,N_1474);
and U1548 (N_1548,N_1463,N_1443);
nor U1549 (N_1549,N_1457,N_1481);
and U1550 (N_1550,N_1497,N_1465);
nor U1551 (N_1551,N_1482,N_1462);
nand U1552 (N_1552,N_1461,N_1465);
nor U1553 (N_1553,N_1486,N_1492);
xnor U1554 (N_1554,N_1467,N_1482);
nand U1555 (N_1555,N_1463,N_1464);
or U1556 (N_1556,N_1484,N_1454);
or U1557 (N_1557,N_1465,N_1472);
or U1558 (N_1558,N_1474,N_1490);
and U1559 (N_1559,N_1460,N_1496);
xnor U1560 (N_1560,N_1553,N_1513);
nand U1561 (N_1561,N_1539,N_1543);
or U1562 (N_1562,N_1506,N_1503);
or U1563 (N_1563,N_1549,N_1557);
xnor U1564 (N_1564,N_1534,N_1530);
and U1565 (N_1565,N_1516,N_1542);
or U1566 (N_1566,N_1515,N_1538);
nand U1567 (N_1567,N_1502,N_1508);
nor U1568 (N_1568,N_1558,N_1509);
nor U1569 (N_1569,N_1531,N_1517);
and U1570 (N_1570,N_1537,N_1545);
or U1571 (N_1571,N_1512,N_1511);
or U1572 (N_1572,N_1533,N_1554);
or U1573 (N_1573,N_1521,N_1550);
or U1574 (N_1574,N_1546,N_1519);
nand U1575 (N_1575,N_1541,N_1535);
nor U1576 (N_1576,N_1536,N_1525);
xnor U1577 (N_1577,N_1529,N_1555);
and U1578 (N_1578,N_1544,N_1552);
nand U1579 (N_1579,N_1520,N_1528);
or U1580 (N_1580,N_1510,N_1559);
and U1581 (N_1581,N_1524,N_1504);
nand U1582 (N_1582,N_1500,N_1527);
nor U1583 (N_1583,N_1501,N_1514);
nor U1584 (N_1584,N_1526,N_1548);
and U1585 (N_1585,N_1556,N_1540);
xor U1586 (N_1586,N_1547,N_1551);
or U1587 (N_1587,N_1523,N_1522);
xnor U1588 (N_1588,N_1505,N_1518);
nor U1589 (N_1589,N_1532,N_1507);
nor U1590 (N_1590,N_1552,N_1554);
nor U1591 (N_1591,N_1548,N_1528);
and U1592 (N_1592,N_1539,N_1547);
nor U1593 (N_1593,N_1515,N_1541);
xor U1594 (N_1594,N_1525,N_1547);
xor U1595 (N_1595,N_1512,N_1540);
or U1596 (N_1596,N_1542,N_1504);
and U1597 (N_1597,N_1547,N_1557);
or U1598 (N_1598,N_1540,N_1542);
nor U1599 (N_1599,N_1511,N_1528);
or U1600 (N_1600,N_1540,N_1541);
xnor U1601 (N_1601,N_1557,N_1506);
xor U1602 (N_1602,N_1505,N_1537);
nor U1603 (N_1603,N_1514,N_1545);
nor U1604 (N_1604,N_1521,N_1532);
and U1605 (N_1605,N_1540,N_1554);
xor U1606 (N_1606,N_1515,N_1522);
nand U1607 (N_1607,N_1522,N_1554);
and U1608 (N_1608,N_1523,N_1547);
and U1609 (N_1609,N_1513,N_1531);
and U1610 (N_1610,N_1528,N_1523);
nor U1611 (N_1611,N_1549,N_1522);
nor U1612 (N_1612,N_1510,N_1519);
or U1613 (N_1613,N_1550,N_1520);
nand U1614 (N_1614,N_1509,N_1512);
nor U1615 (N_1615,N_1528,N_1536);
and U1616 (N_1616,N_1523,N_1559);
and U1617 (N_1617,N_1530,N_1531);
or U1618 (N_1618,N_1532,N_1519);
and U1619 (N_1619,N_1538,N_1524);
or U1620 (N_1620,N_1588,N_1562);
nor U1621 (N_1621,N_1607,N_1563);
nand U1622 (N_1622,N_1606,N_1603);
nand U1623 (N_1623,N_1590,N_1613);
nand U1624 (N_1624,N_1598,N_1584);
and U1625 (N_1625,N_1570,N_1571);
nand U1626 (N_1626,N_1594,N_1569);
and U1627 (N_1627,N_1566,N_1612);
and U1628 (N_1628,N_1580,N_1591);
nor U1629 (N_1629,N_1572,N_1595);
xor U1630 (N_1630,N_1610,N_1611);
nor U1631 (N_1631,N_1589,N_1592);
nor U1632 (N_1632,N_1585,N_1561);
xor U1633 (N_1633,N_1600,N_1575);
nor U1634 (N_1634,N_1615,N_1599);
and U1635 (N_1635,N_1583,N_1596);
or U1636 (N_1636,N_1565,N_1581);
nor U1637 (N_1637,N_1574,N_1573);
or U1638 (N_1638,N_1618,N_1608);
xor U1639 (N_1639,N_1586,N_1597);
nand U1640 (N_1640,N_1619,N_1602);
and U1641 (N_1641,N_1567,N_1564);
xor U1642 (N_1642,N_1604,N_1616);
or U1643 (N_1643,N_1605,N_1601);
and U1644 (N_1644,N_1576,N_1568);
and U1645 (N_1645,N_1617,N_1582);
and U1646 (N_1646,N_1614,N_1577);
xor U1647 (N_1647,N_1587,N_1579);
and U1648 (N_1648,N_1593,N_1560);
nor U1649 (N_1649,N_1578,N_1609);
nand U1650 (N_1650,N_1591,N_1604);
nor U1651 (N_1651,N_1569,N_1582);
nor U1652 (N_1652,N_1593,N_1606);
xnor U1653 (N_1653,N_1599,N_1582);
nor U1654 (N_1654,N_1605,N_1588);
nor U1655 (N_1655,N_1610,N_1583);
or U1656 (N_1656,N_1615,N_1607);
or U1657 (N_1657,N_1596,N_1574);
xnor U1658 (N_1658,N_1594,N_1589);
nand U1659 (N_1659,N_1600,N_1594);
nand U1660 (N_1660,N_1593,N_1582);
xnor U1661 (N_1661,N_1615,N_1570);
nand U1662 (N_1662,N_1617,N_1608);
nand U1663 (N_1663,N_1591,N_1607);
and U1664 (N_1664,N_1611,N_1598);
xor U1665 (N_1665,N_1581,N_1618);
xor U1666 (N_1666,N_1611,N_1600);
or U1667 (N_1667,N_1616,N_1605);
nor U1668 (N_1668,N_1601,N_1610);
nand U1669 (N_1669,N_1587,N_1612);
xnor U1670 (N_1670,N_1605,N_1589);
or U1671 (N_1671,N_1603,N_1592);
xor U1672 (N_1672,N_1570,N_1604);
nand U1673 (N_1673,N_1613,N_1560);
or U1674 (N_1674,N_1614,N_1581);
nand U1675 (N_1675,N_1577,N_1608);
or U1676 (N_1676,N_1615,N_1585);
and U1677 (N_1677,N_1613,N_1577);
xor U1678 (N_1678,N_1570,N_1603);
or U1679 (N_1679,N_1603,N_1594);
nand U1680 (N_1680,N_1671,N_1655);
nor U1681 (N_1681,N_1664,N_1661);
xor U1682 (N_1682,N_1624,N_1623);
or U1683 (N_1683,N_1649,N_1669);
nand U1684 (N_1684,N_1628,N_1676);
nor U1685 (N_1685,N_1657,N_1633);
nand U1686 (N_1686,N_1630,N_1662);
xnor U1687 (N_1687,N_1634,N_1621);
or U1688 (N_1688,N_1620,N_1658);
and U1689 (N_1689,N_1636,N_1635);
xnor U1690 (N_1690,N_1677,N_1679);
nand U1691 (N_1691,N_1643,N_1625);
xor U1692 (N_1692,N_1647,N_1644);
or U1693 (N_1693,N_1639,N_1663);
or U1694 (N_1694,N_1629,N_1654);
xor U1695 (N_1695,N_1656,N_1660);
nand U1696 (N_1696,N_1666,N_1652);
xnor U1697 (N_1697,N_1627,N_1674);
and U1698 (N_1698,N_1641,N_1626);
xnor U1699 (N_1699,N_1653,N_1665);
nor U1700 (N_1700,N_1670,N_1672);
or U1701 (N_1701,N_1632,N_1631);
xnor U1702 (N_1702,N_1646,N_1668);
nor U1703 (N_1703,N_1638,N_1622);
or U1704 (N_1704,N_1667,N_1642);
nor U1705 (N_1705,N_1640,N_1675);
nor U1706 (N_1706,N_1650,N_1659);
xor U1707 (N_1707,N_1637,N_1678);
xor U1708 (N_1708,N_1645,N_1651);
nand U1709 (N_1709,N_1673,N_1648);
and U1710 (N_1710,N_1669,N_1642);
xnor U1711 (N_1711,N_1654,N_1664);
and U1712 (N_1712,N_1624,N_1670);
nor U1713 (N_1713,N_1620,N_1637);
xnor U1714 (N_1714,N_1627,N_1678);
and U1715 (N_1715,N_1671,N_1621);
and U1716 (N_1716,N_1622,N_1673);
and U1717 (N_1717,N_1665,N_1647);
nor U1718 (N_1718,N_1645,N_1673);
or U1719 (N_1719,N_1622,N_1672);
and U1720 (N_1720,N_1640,N_1628);
xnor U1721 (N_1721,N_1657,N_1667);
or U1722 (N_1722,N_1667,N_1661);
xor U1723 (N_1723,N_1675,N_1676);
and U1724 (N_1724,N_1628,N_1677);
xor U1725 (N_1725,N_1620,N_1633);
and U1726 (N_1726,N_1671,N_1678);
nand U1727 (N_1727,N_1640,N_1635);
nor U1728 (N_1728,N_1630,N_1624);
xnor U1729 (N_1729,N_1639,N_1679);
and U1730 (N_1730,N_1640,N_1674);
and U1731 (N_1731,N_1679,N_1622);
xnor U1732 (N_1732,N_1676,N_1641);
xor U1733 (N_1733,N_1624,N_1658);
and U1734 (N_1734,N_1647,N_1626);
nand U1735 (N_1735,N_1635,N_1630);
nor U1736 (N_1736,N_1626,N_1640);
nand U1737 (N_1737,N_1675,N_1663);
nand U1738 (N_1738,N_1667,N_1634);
nor U1739 (N_1739,N_1668,N_1633);
and U1740 (N_1740,N_1727,N_1732);
nor U1741 (N_1741,N_1696,N_1688);
nor U1742 (N_1742,N_1726,N_1703);
nor U1743 (N_1743,N_1736,N_1691);
and U1744 (N_1744,N_1733,N_1693);
and U1745 (N_1745,N_1718,N_1720);
and U1746 (N_1746,N_1735,N_1692);
or U1747 (N_1747,N_1707,N_1687);
and U1748 (N_1748,N_1738,N_1708);
xnor U1749 (N_1749,N_1716,N_1680);
and U1750 (N_1750,N_1694,N_1719);
xnor U1751 (N_1751,N_1689,N_1700);
and U1752 (N_1752,N_1712,N_1690);
nand U1753 (N_1753,N_1717,N_1695);
nor U1754 (N_1754,N_1684,N_1701);
and U1755 (N_1755,N_1724,N_1714);
nor U1756 (N_1756,N_1705,N_1722);
nor U1757 (N_1757,N_1704,N_1706);
xor U1758 (N_1758,N_1713,N_1739);
or U1759 (N_1759,N_1731,N_1737);
nand U1760 (N_1760,N_1728,N_1697);
nor U1761 (N_1761,N_1682,N_1685);
nand U1762 (N_1762,N_1734,N_1711);
xnor U1763 (N_1763,N_1681,N_1699);
and U1764 (N_1764,N_1702,N_1723);
nand U1765 (N_1765,N_1686,N_1683);
xor U1766 (N_1766,N_1725,N_1730);
and U1767 (N_1767,N_1721,N_1709);
xnor U1768 (N_1768,N_1710,N_1729);
nand U1769 (N_1769,N_1715,N_1698);
xnor U1770 (N_1770,N_1726,N_1724);
nand U1771 (N_1771,N_1694,N_1731);
and U1772 (N_1772,N_1701,N_1736);
nand U1773 (N_1773,N_1723,N_1729);
nor U1774 (N_1774,N_1728,N_1707);
or U1775 (N_1775,N_1712,N_1699);
xor U1776 (N_1776,N_1714,N_1689);
nor U1777 (N_1777,N_1734,N_1682);
nor U1778 (N_1778,N_1711,N_1680);
nand U1779 (N_1779,N_1694,N_1722);
and U1780 (N_1780,N_1690,N_1735);
nor U1781 (N_1781,N_1723,N_1720);
xor U1782 (N_1782,N_1730,N_1694);
nand U1783 (N_1783,N_1726,N_1706);
nand U1784 (N_1784,N_1702,N_1738);
and U1785 (N_1785,N_1728,N_1708);
and U1786 (N_1786,N_1681,N_1682);
and U1787 (N_1787,N_1693,N_1729);
or U1788 (N_1788,N_1727,N_1725);
or U1789 (N_1789,N_1688,N_1704);
xnor U1790 (N_1790,N_1708,N_1727);
nor U1791 (N_1791,N_1733,N_1723);
nand U1792 (N_1792,N_1687,N_1699);
or U1793 (N_1793,N_1697,N_1714);
nand U1794 (N_1794,N_1723,N_1708);
or U1795 (N_1795,N_1713,N_1693);
nor U1796 (N_1796,N_1709,N_1729);
nand U1797 (N_1797,N_1691,N_1699);
and U1798 (N_1798,N_1692,N_1720);
or U1799 (N_1799,N_1737,N_1713);
xor U1800 (N_1800,N_1743,N_1755);
xnor U1801 (N_1801,N_1788,N_1741);
or U1802 (N_1802,N_1794,N_1779);
or U1803 (N_1803,N_1762,N_1759);
xor U1804 (N_1804,N_1761,N_1764);
nand U1805 (N_1805,N_1746,N_1772);
xor U1806 (N_1806,N_1750,N_1742);
or U1807 (N_1807,N_1752,N_1773);
xor U1808 (N_1808,N_1757,N_1781);
or U1809 (N_1809,N_1778,N_1753);
and U1810 (N_1810,N_1744,N_1776);
xor U1811 (N_1811,N_1748,N_1767);
nand U1812 (N_1812,N_1769,N_1754);
and U1813 (N_1813,N_1798,N_1774);
or U1814 (N_1814,N_1787,N_1784);
and U1815 (N_1815,N_1796,N_1747);
nor U1816 (N_1816,N_1740,N_1770);
xnor U1817 (N_1817,N_1777,N_1760);
or U1818 (N_1818,N_1789,N_1780);
xnor U1819 (N_1819,N_1751,N_1745);
or U1820 (N_1820,N_1771,N_1766);
xnor U1821 (N_1821,N_1795,N_1790);
xnor U1822 (N_1822,N_1785,N_1782);
nor U1823 (N_1823,N_1749,N_1775);
nand U1824 (N_1824,N_1793,N_1765);
or U1825 (N_1825,N_1768,N_1797);
and U1826 (N_1826,N_1799,N_1758);
nor U1827 (N_1827,N_1783,N_1763);
nand U1828 (N_1828,N_1756,N_1786);
or U1829 (N_1829,N_1792,N_1791);
nor U1830 (N_1830,N_1746,N_1748);
nand U1831 (N_1831,N_1798,N_1763);
nand U1832 (N_1832,N_1796,N_1772);
or U1833 (N_1833,N_1745,N_1788);
nand U1834 (N_1834,N_1766,N_1743);
nand U1835 (N_1835,N_1754,N_1766);
xor U1836 (N_1836,N_1796,N_1757);
xor U1837 (N_1837,N_1741,N_1757);
nand U1838 (N_1838,N_1783,N_1745);
nand U1839 (N_1839,N_1785,N_1781);
nor U1840 (N_1840,N_1763,N_1746);
nand U1841 (N_1841,N_1771,N_1741);
or U1842 (N_1842,N_1782,N_1747);
nand U1843 (N_1843,N_1778,N_1790);
and U1844 (N_1844,N_1787,N_1770);
nand U1845 (N_1845,N_1777,N_1787);
nor U1846 (N_1846,N_1781,N_1764);
or U1847 (N_1847,N_1773,N_1794);
nor U1848 (N_1848,N_1744,N_1775);
and U1849 (N_1849,N_1775,N_1752);
and U1850 (N_1850,N_1794,N_1750);
and U1851 (N_1851,N_1759,N_1792);
xor U1852 (N_1852,N_1740,N_1774);
nor U1853 (N_1853,N_1770,N_1751);
or U1854 (N_1854,N_1799,N_1790);
xnor U1855 (N_1855,N_1799,N_1750);
or U1856 (N_1856,N_1752,N_1751);
or U1857 (N_1857,N_1753,N_1782);
or U1858 (N_1858,N_1774,N_1796);
nor U1859 (N_1859,N_1797,N_1777);
or U1860 (N_1860,N_1857,N_1814);
xnor U1861 (N_1861,N_1809,N_1819);
and U1862 (N_1862,N_1813,N_1833);
nor U1863 (N_1863,N_1802,N_1811);
and U1864 (N_1864,N_1817,N_1847);
or U1865 (N_1865,N_1842,N_1841);
xor U1866 (N_1866,N_1827,N_1822);
or U1867 (N_1867,N_1821,N_1828);
nor U1868 (N_1868,N_1806,N_1855);
xnor U1869 (N_1869,N_1848,N_1820);
xor U1870 (N_1870,N_1812,N_1826);
nand U1871 (N_1871,N_1803,N_1840);
nand U1872 (N_1872,N_1844,N_1851);
or U1873 (N_1873,N_1832,N_1843);
or U1874 (N_1874,N_1853,N_1830);
xor U1875 (N_1875,N_1856,N_1849);
and U1876 (N_1876,N_1859,N_1831);
xnor U1877 (N_1877,N_1823,N_1845);
nand U1878 (N_1878,N_1854,N_1837);
or U1879 (N_1879,N_1829,N_1858);
or U1880 (N_1880,N_1835,N_1836);
xnor U1881 (N_1881,N_1815,N_1839);
and U1882 (N_1882,N_1810,N_1838);
nand U1883 (N_1883,N_1852,N_1805);
and U1884 (N_1884,N_1846,N_1834);
nand U1885 (N_1885,N_1808,N_1824);
or U1886 (N_1886,N_1801,N_1850);
nor U1887 (N_1887,N_1807,N_1816);
xor U1888 (N_1888,N_1818,N_1800);
and U1889 (N_1889,N_1825,N_1804);
xor U1890 (N_1890,N_1804,N_1836);
and U1891 (N_1891,N_1823,N_1857);
xor U1892 (N_1892,N_1842,N_1820);
and U1893 (N_1893,N_1841,N_1808);
and U1894 (N_1894,N_1806,N_1841);
and U1895 (N_1895,N_1821,N_1837);
and U1896 (N_1896,N_1803,N_1835);
nand U1897 (N_1897,N_1855,N_1848);
xnor U1898 (N_1898,N_1833,N_1804);
nor U1899 (N_1899,N_1852,N_1827);
nand U1900 (N_1900,N_1852,N_1804);
nand U1901 (N_1901,N_1835,N_1817);
xor U1902 (N_1902,N_1820,N_1854);
nor U1903 (N_1903,N_1829,N_1857);
xnor U1904 (N_1904,N_1839,N_1824);
nand U1905 (N_1905,N_1837,N_1835);
xor U1906 (N_1906,N_1827,N_1853);
or U1907 (N_1907,N_1810,N_1832);
nor U1908 (N_1908,N_1813,N_1821);
and U1909 (N_1909,N_1810,N_1857);
nor U1910 (N_1910,N_1816,N_1812);
and U1911 (N_1911,N_1814,N_1810);
or U1912 (N_1912,N_1824,N_1854);
xnor U1913 (N_1913,N_1835,N_1832);
and U1914 (N_1914,N_1800,N_1846);
or U1915 (N_1915,N_1858,N_1825);
nor U1916 (N_1916,N_1801,N_1824);
and U1917 (N_1917,N_1837,N_1809);
and U1918 (N_1918,N_1830,N_1858);
nor U1919 (N_1919,N_1830,N_1854);
or U1920 (N_1920,N_1860,N_1875);
nand U1921 (N_1921,N_1919,N_1866);
xor U1922 (N_1922,N_1887,N_1904);
and U1923 (N_1923,N_1890,N_1883);
nand U1924 (N_1924,N_1898,N_1865);
xor U1925 (N_1925,N_1906,N_1910);
nor U1926 (N_1926,N_1902,N_1889);
nor U1927 (N_1927,N_1907,N_1894);
nor U1928 (N_1928,N_1897,N_1908);
and U1929 (N_1929,N_1879,N_1899);
and U1930 (N_1930,N_1881,N_1909);
nand U1931 (N_1931,N_1882,N_1903);
xnor U1932 (N_1932,N_1916,N_1874);
or U1933 (N_1933,N_1884,N_1869);
and U1934 (N_1934,N_1867,N_1873);
nor U1935 (N_1935,N_1868,N_1870);
or U1936 (N_1936,N_1915,N_1862);
xor U1937 (N_1937,N_1905,N_1878);
nand U1938 (N_1938,N_1871,N_1888);
nand U1939 (N_1939,N_1917,N_1896);
and U1940 (N_1940,N_1913,N_1893);
and U1941 (N_1941,N_1885,N_1912);
or U1942 (N_1942,N_1914,N_1872);
nand U1943 (N_1943,N_1880,N_1863);
and U1944 (N_1944,N_1891,N_1901);
xor U1945 (N_1945,N_1900,N_1895);
nor U1946 (N_1946,N_1876,N_1886);
xor U1947 (N_1947,N_1864,N_1892);
nand U1948 (N_1948,N_1911,N_1877);
nand U1949 (N_1949,N_1861,N_1918);
xnor U1950 (N_1950,N_1899,N_1886);
nor U1951 (N_1951,N_1903,N_1885);
xor U1952 (N_1952,N_1863,N_1865);
and U1953 (N_1953,N_1897,N_1910);
xnor U1954 (N_1954,N_1914,N_1907);
nand U1955 (N_1955,N_1869,N_1910);
xor U1956 (N_1956,N_1905,N_1883);
or U1957 (N_1957,N_1861,N_1885);
xor U1958 (N_1958,N_1897,N_1887);
or U1959 (N_1959,N_1864,N_1869);
or U1960 (N_1960,N_1872,N_1896);
and U1961 (N_1961,N_1891,N_1914);
nor U1962 (N_1962,N_1912,N_1915);
nor U1963 (N_1963,N_1896,N_1904);
and U1964 (N_1964,N_1900,N_1917);
xor U1965 (N_1965,N_1867,N_1864);
or U1966 (N_1966,N_1879,N_1891);
or U1967 (N_1967,N_1898,N_1913);
xnor U1968 (N_1968,N_1867,N_1878);
or U1969 (N_1969,N_1900,N_1889);
xor U1970 (N_1970,N_1895,N_1916);
and U1971 (N_1971,N_1919,N_1869);
xnor U1972 (N_1972,N_1911,N_1891);
nand U1973 (N_1973,N_1909,N_1868);
nand U1974 (N_1974,N_1864,N_1907);
or U1975 (N_1975,N_1865,N_1877);
or U1976 (N_1976,N_1874,N_1894);
nand U1977 (N_1977,N_1875,N_1869);
or U1978 (N_1978,N_1906,N_1880);
or U1979 (N_1979,N_1914,N_1885);
nor U1980 (N_1980,N_1935,N_1955);
nand U1981 (N_1981,N_1952,N_1928);
and U1982 (N_1982,N_1929,N_1964);
or U1983 (N_1983,N_1930,N_1946);
and U1984 (N_1984,N_1934,N_1961);
xor U1985 (N_1985,N_1933,N_1979);
nor U1986 (N_1986,N_1939,N_1957);
nor U1987 (N_1987,N_1976,N_1925);
xnor U1988 (N_1988,N_1927,N_1954);
nor U1989 (N_1989,N_1958,N_1953);
xnor U1990 (N_1990,N_1969,N_1973);
xnor U1991 (N_1991,N_1975,N_1970);
and U1992 (N_1992,N_1950,N_1966);
xnor U1993 (N_1993,N_1949,N_1947);
nor U1994 (N_1994,N_1924,N_1972);
and U1995 (N_1995,N_1920,N_1959);
xor U1996 (N_1996,N_1974,N_1923);
or U1997 (N_1997,N_1956,N_1962);
and U1998 (N_1998,N_1941,N_1922);
or U1999 (N_1999,N_1932,N_1968);
or U2000 (N_2000,N_1971,N_1965);
nor U2001 (N_2001,N_1943,N_1945);
or U2002 (N_2002,N_1978,N_1942);
xor U2003 (N_2003,N_1948,N_1921);
nor U2004 (N_2004,N_1960,N_1940);
and U2005 (N_2005,N_1937,N_1977);
nor U2006 (N_2006,N_1944,N_1963);
xnor U2007 (N_2007,N_1931,N_1936);
or U2008 (N_2008,N_1926,N_1967);
nor U2009 (N_2009,N_1951,N_1938);
xor U2010 (N_2010,N_1948,N_1949);
and U2011 (N_2011,N_1971,N_1931);
or U2012 (N_2012,N_1969,N_1961);
nor U2013 (N_2013,N_1961,N_1922);
nor U2014 (N_2014,N_1967,N_1963);
or U2015 (N_2015,N_1975,N_1939);
nor U2016 (N_2016,N_1963,N_1951);
xnor U2017 (N_2017,N_1977,N_1974);
nand U2018 (N_2018,N_1920,N_1942);
or U2019 (N_2019,N_1979,N_1961);
nand U2020 (N_2020,N_1979,N_1978);
or U2021 (N_2021,N_1978,N_1931);
or U2022 (N_2022,N_1940,N_1938);
nor U2023 (N_2023,N_1949,N_1937);
nand U2024 (N_2024,N_1943,N_1964);
or U2025 (N_2025,N_1978,N_1923);
nor U2026 (N_2026,N_1968,N_1920);
or U2027 (N_2027,N_1922,N_1946);
nor U2028 (N_2028,N_1936,N_1959);
nor U2029 (N_2029,N_1967,N_1969);
xnor U2030 (N_2030,N_1938,N_1964);
and U2031 (N_2031,N_1941,N_1961);
or U2032 (N_2032,N_1951,N_1961);
or U2033 (N_2033,N_1976,N_1952);
nand U2034 (N_2034,N_1963,N_1923);
xnor U2035 (N_2035,N_1924,N_1929);
xor U2036 (N_2036,N_1958,N_1928);
xnor U2037 (N_2037,N_1952,N_1949);
or U2038 (N_2038,N_1935,N_1965);
or U2039 (N_2039,N_1979,N_1960);
or U2040 (N_2040,N_2012,N_2000);
nor U2041 (N_2041,N_2038,N_2031);
nor U2042 (N_2042,N_2032,N_1981);
and U2043 (N_2043,N_1998,N_1992);
xnor U2044 (N_2044,N_2035,N_1997);
nand U2045 (N_2045,N_2018,N_1983);
xnor U2046 (N_2046,N_2036,N_1988);
xnor U2047 (N_2047,N_2013,N_1982);
or U2048 (N_2048,N_2024,N_2007);
and U2049 (N_2049,N_2015,N_2004);
xor U2050 (N_2050,N_2028,N_2005);
nand U2051 (N_2051,N_2001,N_1994);
xnor U2052 (N_2052,N_1989,N_2016);
and U2053 (N_2053,N_2008,N_1987);
nor U2054 (N_2054,N_2039,N_1996);
nor U2055 (N_2055,N_2029,N_2026);
and U2056 (N_2056,N_2037,N_2003);
nor U2057 (N_2057,N_2021,N_1984);
nor U2058 (N_2058,N_2002,N_2017);
and U2059 (N_2059,N_2022,N_1995);
nand U2060 (N_2060,N_2011,N_1990);
nand U2061 (N_2061,N_2027,N_2023);
nor U2062 (N_2062,N_2034,N_2030);
nor U2063 (N_2063,N_1999,N_2009);
nand U2064 (N_2064,N_1993,N_2006);
nor U2065 (N_2065,N_2014,N_1980);
and U2066 (N_2066,N_1991,N_2020);
xor U2067 (N_2067,N_1986,N_1985);
nor U2068 (N_2068,N_2019,N_2010);
nand U2069 (N_2069,N_2033,N_2025);
nor U2070 (N_2070,N_2016,N_2034);
xnor U2071 (N_2071,N_2014,N_2037);
or U2072 (N_2072,N_1995,N_2005);
xnor U2073 (N_2073,N_1988,N_1998);
and U2074 (N_2074,N_2018,N_2010);
or U2075 (N_2075,N_2016,N_2013);
nor U2076 (N_2076,N_1993,N_1987);
or U2077 (N_2077,N_2023,N_2013);
nand U2078 (N_2078,N_2033,N_2024);
or U2079 (N_2079,N_2037,N_2018);
and U2080 (N_2080,N_1991,N_2033);
xor U2081 (N_2081,N_2013,N_2021);
nand U2082 (N_2082,N_2027,N_1997);
or U2083 (N_2083,N_1981,N_1996);
or U2084 (N_2084,N_2002,N_2022);
xnor U2085 (N_2085,N_2009,N_2021);
xnor U2086 (N_2086,N_2022,N_2017);
or U2087 (N_2087,N_1986,N_2033);
and U2088 (N_2088,N_2016,N_2000);
nand U2089 (N_2089,N_1981,N_2025);
or U2090 (N_2090,N_2036,N_2019);
nand U2091 (N_2091,N_2036,N_1990);
nand U2092 (N_2092,N_1998,N_2009);
and U2093 (N_2093,N_2005,N_1983);
and U2094 (N_2094,N_2008,N_2033);
or U2095 (N_2095,N_1983,N_1998);
or U2096 (N_2096,N_2029,N_2037);
nand U2097 (N_2097,N_2022,N_1985);
xor U2098 (N_2098,N_2005,N_2027);
or U2099 (N_2099,N_1995,N_2028);
nor U2100 (N_2100,N_2088,N_2077);
nand U2101 (N_2101,N_2067,N_2086);
nor U2102 (N_2102,N_2081,N_2092);
nor U2103 (N_2103,N_2089,N_2048);
nand U2104 (N_2104,N_2068,N_2076);
nor U2105 (N_2105,N_2073,N_2065);
xor U2106 (N_2106,N_2043,N_2083);
and U2107 (N_2107,N_2079,N_2060);
nand U2108 (N_2108,N_2069,N_2064);
nor U2109 (N_2109,N_2087,N_2082);
nand U2110 (N_2110,N_2097,N_2053);
or U2111 (N_2111,N_2090,N_2072);
xor U2112 (N_2112,N_2084,N_2061);
nor U2113 (N_2113,N_2044,N_2091);
xnor U2114 (N_2114,N_2098,N_2099);
nand U2115 (N_2115,N_2071,N_2045);
and U2116 (N_2116,N_2057,N_2050);
nor U2117 (N_2117,N_2049,N_2059);
nor U2118 (N_2118,N_2074,N_2047);
xor U2119 (N_2119,N_2056,N_2080);
nor U2120 (N_2120,N_2041,N_2046);
or U2121 (N_2121,N_2075,N_2042);
nor U2122 (N_2122,N_2063,N_2052);
and U2123 (N_2123,N_2066,N_2070);
or U2124 (N_2124,N_2062,N_2058);
xnor U2125 (N_2125,N_2055,N_2094);
or U2126 (N_2126,N_2078,N_2085);
nor U2127 (N_2127,N_2095,N_2096);
and U2128 (N_2128,N_2093,N_2054);
xor U2129 (N_2129,N_2051,N_2040);
xor U2130 (N_2130,N_2048,N_2069);
and U2131 (N_2131,N_2083,N_2089);
nand U2132 (N_2132,N_2058,N_2045);
or U2133 (N_2133,N_2088,N_2091);
and U2134 (N_2134,N_2076,N_2050);
nand U2135 (N_2135,N_2087,N_2043);
xor U2136 (N_2136,N_2053,N_2058);
xor U2137 (N_2137,N_2084,N_2093);
nor U2138 (N_2138,N_2089,N_2071);
nor U2139 (N_2139,N_2094,N_2056);
xnor U2140 (N_2140,N_2089,N_2082);
nand U2141 (N_2141,N_2051,N_2095);
or U2142 (N_2142,N_2048,N_2076);
nand U2143 (N_2143,N_2062,N_2073);
and U2144 (N_2144,N_2071,N_2070);
or U2145 (N_2145,N_2087,N_2057);
and U2146 (N_2146,N_2066,N_2072);
xnor U2147 (N_2147,N_2084,N_2076);
xnor U2148 (N_2148,N_2050,N_2051);
or U2149 (N_2149,N_2054,N_2091);
or U2150 (N_2150,N_2064,N_2047);
xnor U2151 (N_2151,N_2082,N_2076);
and U2152 (N_2152,N_2046,N_2053);
and U2153 (N_2153,N_2058,N_2047);
or U2154 (N_2154,N_2046,N_2073);
xnor U2155 (N_2155,N_2083,N_2064);
xor U2156 (N_2156,N_2065,N_2043);
nor U2157 (N_2157,N_2072,N_2095);
nor U2158 (N_2158,N_2080,N_2076);
xnor U2159 (N_2159,N_2071,N_2090);
or U2160 (N_2160,N_2153,N_2136);
nor U2161 (N_2161,N_2110,N_2150);
nor U2162 (N_2162,N_2147,N_2130);
nor U2163 (N_2163,N_2106,N_2133);
or U2164 (N_2164,N_2132,N_2125);
nor U2165 (N_2165,N_2141,N_2154);
nand U2166 (N_2166,N_2121,N_2142);
xnor U2167 (N_2167,N_2139,N_2155);
or U2168 (N_2168,N_2135,N_2137);
nand U2169 (N_2169,N_2124,N_2118);
nor U2170 (N_2170,N_2152,N_2128);
or U2171 (N_2171,N_2158,N_2129);
or U2172 (N_2172,N_2145,N_2157);
nor U2173 (N_2173,N_2159,N_2107);
xnor U2174 (N_2174,N_2149,N_2127);
nand U2175 (N_2175,N_2119,N_2120);
and U2176 (N_2176,N_2100,N_2151);
and U2177 (N_2177,N_2111,N_2156);
or U2178 (N_2178,N_2122,N_2138);
nand U2179 (N_2179,N_2104,N_2105);
xor U2180 (N_2180,N_2101,N_2126);
and U2181 (N_2181,N_2146,N_2123);
nand U2182 (N_2182,N_2117,N_2114);
and U2183 (N_2183,N_2113,N_2115);
xor U2184 (N_2184,N_2144,N_2109);
or U2185 (N_2185,N_2108,N_2134);
xnor U2186 (N_2186,N_2112,N_2116);
xnor U2187 (N_2187,N_2131,N_2140);
nor U2188 (N_2188,N_2143,N_2102);
or U2189 (N_2189,N_2103,N_2148);
nand U2190 (N_2190,N_2132,N_2111);
nor U2191 (N_2191,N_2115,N_2120);
and U2192 (N_2192,N_2100,N_2122);
nor U2193 (N_2193,N_2149,N_2135);
nand U2194 (N_2194,N_2129,N_2136);
nand U2195 (N_2195,N_2125,N_2114);
nand U2196 (N_2196,N_2107,N_2153);
or U2197 (N_2197,N_2128,N_2140);
nor U2198 (N_2198,N_2139,N_2153);
nand U2199 (N_2199,N_2128,N_2144);
nor U2200 (N_2200,N_2116,N_2108);
or U2201 (N_2201,N_2128,N_2116);
xnor U2202 (N_2202,N_2151,N_2144);
xor U2203 (N_2203,N_2112,N_2151);
and U2204 (N_2204,N_2112,N_2126);
and U2205 (N_2205,N_2100,N_2148);
or U2206 (N_2206,N_2124,N_2112);
nor U2207 (N_2207,N_2127,N_2151);
or U2208 (N_2208,N_2130,N_2141);
xor U2209 (N_2209,N_2138,N_2127);
xor U2210 (N_2210,N_2153,N_2115);
xor U2211 (N_2211,N_2148,N_2117);
xnor U2212 (N_2212,N_2150,N_2118);
nor U2213 (N_2213,N_2103,N_2145);
xnor U2214 (N_2214,N_2104,N_2111);
and U2215 (N_2215,N_2121,N_2101);
xor U2216 (N_2216,N_2116,N_2114);
and U2217 (N_2217,N_2123,N_2132);
nand U2218 (N_2218,N_2124,N_2146);
or U2219 (N_2219,N_2126,N_2134);
nand U2220 (N_2220,N_2191,N_2212);
nand U2221 (N_2221,N_2170,N_2199);
and U2222 (N_2222,N_2219,N_2171);
nor U2223 (N_2223,N_2196,N_2164);
or U2224 (N_2224,N_2218,N_2189);
and U2225 (N_2225,N_2175,N_2167);
and U2226 (N_2226,N_2190,N_2188);
nor U2227 (N_2227,N_2216,N_2177);
nor U2228 (N_2228,N_2179,N_2180);
and U2229 (N_2229,N_2206,N_2161);
and U2230 (N_2230,N_2181,N_2176);
nand U2231 (N_2231,N_2204,N_2178);
and U2232 (N_2232,N_2165,N_2202);
or U2233 (N_2233,N_2186,N_2185);
xnor U2234 (N_2234,N_2208,N_2211);
or U2235 (N_2235,N_2210,N_2166);
and U2236 (N_2236,N_2183,N_2197);
xor U2237 (N_2237,N_2184,N_2214);
nand U2238 (N_2238,N_2194,N_2160);
and U2239 (N_2239,N_2201,N_2172);
or U2240 (N_2240,N_2192,N_2195);
xor U2241 (N_2241,N_2193,N_2174);
nand U2242 (N_2242,N_2215,N_2182);
nor U2243 (N_2243,N_2173,N_2162);
nor U2244 (N_2244,N_2169,N_2198);
nand U2245 (N_2245,N_2168,N_2200);
nor U2246 (N_2246,N_2207,N_2213);
nor U2247 (N_2247,N_2163,N_2205);
nand U2248 (N_2248,N_2187,N_2209);
nand U2249 (N_2249,N_2203,N_2217);
nand U2250 (N_2250,N_2193,N_2197);
xnor U2251 (N_2251,N_2209,N_2210);
nand U2252 (N_2252,N_2208,N_2177);
nor U2253 (N_2253,N_2205,N_2177);
nor U2254 (N_2254,N_2209,N_2202);
or U2255 (N_2255,N_2219,N_2185);
nor U2256 (N_2256,N_2205,N_2197);
or U2257 (N_2257,N_2209,N_2190);
and U2258 (N_2258,N_2163,N_2213);
and U2259 (N_2259,N_2197,N_2194);
and U2260 (N_2260,N_2189,N_2179);
or U2261 (N_2261,N_2210,N_2208);
and U2262 (N_2262,N_2214,N_2173);
nor U2263 (N_2263,N_2190,N_2196);
xnor U2264 (N_2264,N_2185,N_2160);
nand U2265 (N_2265,N_2177,N_2168);
nor U2266 (N_2266,N_2175,N_2186);
nand U2267 (N_2267,N_2169,N_2185);
nand U2268 (N_2268,N_2190,N_2219);
and U2269 (N_2269,N_2185,N_2207);
xor U2270 (N_2270,N_2160,N_2179);
or U2271 (N_2271,N_2179,N_2204);
or U2272 (N_2272,N_2168,N_2212);
nor U2273 (N_2273,N_2200,N_2207);
nand U2274 (N_2274,N_2204,N_2195);
and U2275 (N_2275,N_2212,N_2195);
nand U2276 (N_2276,N_2195,N_2215);
nand U2277 (N_2277,N_2178,N_2209);
or U2278 (N_2278,N_2178,N_2184);
and U2279 (N_2279,N_2213,N_2198);
and U2280 (N_2280,N_2229,N_2237);
nand U2281 (N_2281,N_2233,N_2279);
xor U2282 (N_2282,N_2223,N_2245);
or U2283 (N_2283,N_2228,N_2267);
xor U2284 (N_2284,N_2240,N_2260);
xnor U2285 (N_2285,N_2221,N_2269);
xor U2286 (N_2286,N_2275,N_2261);
nor U2287 (N_2287,N_2255,N_2254);
nand U2288 (N_2288,N_2250,N_2263);
nor U2289 (N_2289,N_2244,N_2256);
or U2290 (N_2290,N_2276,N_2270);
and U2291 (N_2291,N_2220,N_2234);
xor U2292 (N_2292,N_2265,N_2273);
nand U2293 (N_2293,N_2238,N_2262);
and U2294 (N_2294,N_2231,N_2251);
or U2295 (N_2295,N_2246,N_2259);
or U2296 (N_2296,N_2257,N_2230);
and U2297 (N_2297,N_2271,N_2268);
or U2298 (N_2298,N_2222,N_2278);
or U2299 (N_2299,N_2243,N_2227);
and U2300 (N_2300,N_2266,N_2252);
xor U2301 (N_2301,N_2224,N_2277);
nand U2302 (N_2302,N_2249,N_2236);
nor U2303 (N_2303,N_2242,N_2226);
nand U2304 (N_2304,N_2232,N_2247);
xnor U2305 (N_2305,N_2272,N_2264);
nor U2306 (N_2306,N_2258,N_2274);
nor U2307 (N_2307,N_2253,N_2239);
nor U2308 (N_2308,N_2241,N_2225);
nor U2309 (N_2309,N_2235,N_2248);
xor U2310 (N_2310,N_2263,N_2239);
xor U2311 (N_2311,N_2236,N_2238);
nand U2312 (N_2312,N_2265,N_2254);
nand U2313 (N_2313,N_2243,N_2245);
xor U2314 (N_2314,N_2257,N_2238);
and U2315 (N_2315,N_2246,N_2233);
or U2316 (N_2316,N_2279,N_2270);
nor U2317 (N_2317,N_2276,N_2227);
nor U2318 (N_2318,N_2235,N_2236);
and U2319 (N_2319,N_2249,N_2257);
nand U2320 (N_2320,N_2232,N_2269);
xnor U2321 (N_2321,N_2272,N_2238);
nor U2322 (N_2322,N_2264,N_2251);
nor U2323 (N_2323,N_2247,N_2234);
nor U2324 (N_2324,N_2266,N_2253);
nand U2325 (N_2325,N_2226,N_2264);
nand U2326 (N_2326,N_2270,N_2254);
or U2327 (N_2327,N_2250,N_2257);
and U2328 (N_2328,N_2275,N_2237);
and U2329 (N_2329,N_2231,N_2259);
nand U2330 (N_2330,N_2235,N_2240);
nor U2331 (N_2331,N_2254,N_2245);
and U2332 (N_2332,N_2229,N_2235);
nand U2333 (N_2333,N_2245,N_2231);
nand U2334 (N_2334,N_2262,N_2223);
or U2335 (N_2335,N_2236,N_2262);
xor U2336 (N_2336,N_2232,N_2271);
nand U2337 (N_2337,N_2239,N_2244);
or U2338 (N_2338,N_2251,N_2272);
or U2339 (N_2339,N_2232,N_2224);
nand U2340 (N_2340,N_2331,N_2329);
and U2341 (N_2341,N_2307,N_2322);
nand U2342 (N_2342,N_2287,N_2300);
nor U2343 (N_2343,N_2317,N_2292);
nand U2344 (N_2344,N_2304,N_2321);
nand U2345 (N_2345,N_2325,N_2294);
nor U2346 (N_2346,N_2282,N_2326);
and U2347 (N_2347,N_2296,N_2323);
nor U2348 (N_2348,N_2285,N_2299);
and U2349 (N_2349,N_2291,N_2303);
nand U2350 (N_2350,N_2314,N_2332);
nand U2351 (N_2351,N_2335,N_2301);
nor U2352 (N_2352,N_2284,N_2308);
or U2353 (N_2353,N_2283,N_2336);
xnor U2354 (N_2354,N_2313,N_2315);
xor U2355 (N_2355,N_2298,N_2286);
and U2356 (N_2356,N_2310,N_2328);
nor U2357 (N_2357,N_2320,N_2318);
nand U2358 (N_2358,N_2338,N_2330);
or U2359 (N_2359,N_2319,N_2281);
and U2360 (N_2360,N_2302,N_2337);
nand U2361 (N_2361,N_2293,N_2290);
or U2362 (N_2362,N_2295,N_2312);
or U2363 (N_2363,N_2297,N_2333);
nor U2364 (N_2364,N_2316,N_2309);
and U2365 (N_2365,N_2311,N_2324);
and U2366 (N_2366,N_2306,N_2327);
xor U2367 (N_2367,N_2280,N_2288);
and U2368 (N_2368,N_2305,N_2334);
nand U2369 (N_2369,N_2289,N_2339);
or U2370 (N_2370,N_2291,N_2280);
nand U2371 (N_2371,N_2338,N_2299);
or U2372 (N_2372,N_2315,N_2324);
nand U2373 (N_2373,N_2309,N_2294);
nor U2374 (N_2374,N_2307,N_2309);
and U2375 (N_2375,N_2288,N_2292);
and U2376 (N_2376,N_2311,N_2286);
nand U2377 (N_2377,N_2307,N_2311);
xor U2378 (N_2378,N_2313,N_2317);
or U2379 (N_2379,N_2325,N_2313);
or U2380 (N_2380,N_2320,N_2304);
nand U2381 (N_2381,N_2297,N_2307);
nand U2382 (N_2382,N_2316,N_2293);
or U2383 (N_2383,N_2338,N_2339);
or U2384 (N_2384,N_2306,N_2331);
nand U2385 (N_2385,N_2336,N_2314);
nor U2386 (N_2386,N_2320,N_2305);
xnor U2387 (N_2387,N_2312,N_2322);
xnor U2388 (N_2388,N_2336,N_2317);
nand U2389 (N_2389,N_2288,N_2286);
nor U2390 (N_2390,N_2302,N_2303);
or U2391 (N_2391,N_2330,N_2300);
or U2392 (N_2392,N_2293,N_2285);
nor U2393 (N_2393,N_2288,N_2312);
nor U2394 (N_2394,N_2326,N_2324);
or U2395 (N_2395,N_2303,N_2329);
or U2396 (N_2396,N_2333,N_2323);
and U2397 (N_2397,N_2296,N_2334);
or U2398 (N_2398,N_2301,N_2309);
nand U2399 (N_2399,N_2293,N_2283);
xnor U2400 (N_2400,N_2399,N_2374);
nand U2401 (N_2401,N_2384,N_2358);
nand U2402 (N_2402,N_2343,N_2379);
xnor U2403 (N_2403,N_2372,N_2357);
xnor U2404 (N_2404,N_2363,N_2392);
or U2405 (N_2405,N_2345,N_2395);
or U2406 (N_2406,N_2370,N_2362);
nor U2407 (N_2407,N_2366,N_2356);
and U2408 (N_2408,N_2382,N_2368);
or U2409 (N_2409,N_2386,N_2398);
nand U2410 (N_2410,N_2355,N_2342);
or U2411 (N_2411,N_2394,N_2364);
and U2412 (N_2412,N_2361,N_2348);
nor U2413 (N_2413,N_2391,N_2371);
nor U2414 (N_2414,N_2350,N_2365);
nand U2415 (N_2415,N_2377,N_2346);
nand U2416 (N_2416,N_2385,N_2351);
nand U2417 (N_2417,N_2359,N_2390);
nor U2418 (N_2418,N_2344,N_2378);
nor U2419 (N_2419,N_2341,N_2360);
nand U2420 (N_2420,N_2375,N_2352);
nand U2421 (N_2421,N_2349,N_2340);
or U2422 (N_2422,N_2367,N_2369);
or U2423 (N_2423,N_2396,N_2381);
and U2424 (N_2424,N_2387,N_2354);
nor U2425 (N_2425,N_2393,N_2397);
xnor U2426 (N_2426,N_2373,N_2389);
or U2427 (N_2427,N_2380,N_2376);
nor U2428 (N_2428,N_2388,N_2383);
nand U2429 (N_2429,N_2353,N_2347);
nand U2430 (N_2430,N_2370,N_2384);
nor U2431 (N_2431,N_2360,N_2347);
nand U2432 (N_2432,N_2364,N_2366);
xnor U2433 (N_2433,N_2363,N_2384);
and U2434 (N_2434,N_2362,N_2353);
or U2435 (N_2435,N_2347,N_2396);
nand U2436 (N_2436,N_2343,N_2373);
nand U2437 (N_2437,N_2353,N_2396);
or U2438 (N_2438,N_2346,N_2380);
and U2439 (N_2439,N_2378,N_2355);
and U2440 (N_2440,N_2382,N_2359);
nor U2441 (N_2441,N_2391,N_2372);
xor U2442 (N_2442,N_2391,N_2383);
nand U2443 (N_2443,N_2351,N_2353);
and U2444 (N_2444,N_2350,N_2358);
and U2445 (N_2445,N_2385,N_2387);
or U2446 (N_2446,N_2354,N_2344);
nand U2447 (N_2447,N_2386,N_2341);
nand U2448 (N_2448,N_2380,N_2352);
nor U2449 (N_2449,N_2354,N_2348);
nor U2450 (N_2450,N_2388,N_2360);
xnor U2451 (N_2451,N_2375,N_2351);
and U2452 (N_2452,N_2356,N_2353);
xor U2453 (N_2453,N_2364,N_2350);
xor U2454 (N_2454,N_2392,N_2395);
nor U2455 (N_2455,N_2343,N_2345);
nand U2456 (N_2456,N_2378,N_2356);
and U2457 (N_2457,N_2352,N_2384);
nand U2458 (N_2458,N_2368,N_2349);
xnor U2459 (N_2459,N_2398,N_2362);
and U2460 (N_2460,N_2402,N_2413);
xnor U2461 (N_2461,N_2440,N_2442);
xor U2462 (N_2462,N_2453,N_2456);
xnor U2463 (N_2463,N_2437,N_2421);
nand U2464 (N_2464,N_2430,N_2435);
xnor U2465 (N_2465,N_2408,N_2427);
nand U2466 (N_2466,N_2415,N_2443);
nand U2467 (N_2467,N_2410,N_2401);
xnor U2468 (N_2468,N_2425,N_2436);
nor U2469 (N_2469,N_2438,N_2448);
nand U2470 (N_2470,N_2444,N_2400);
nor U2471 (N_2471,N_2459,N_2452);
or U2472 (N_2472,N_2420,N_2439);
xor U2473 (N_2473,N_2423,N_2451);
nand U2474 (N_2474,N_2446,N_2416);
nor U2475 (N_2475,N_2414,N_2412);
and U2476 (N_2476,N_2445,N_2411);
xor U2477 (N_2477,N_2405,N_2450);
nand U2478 (N_2478,N_2422,N_2426);
or U2479 (N_2479,N_2418,N_2424);
nor U2480 (N_2480,N_2417,N_2447);
xnor U2481 (N_2481,N_2441,N_2403);
nor U2482 (N_2482,N_2429,N_2406);
or U2483 (N_2483,N_2458,N_2428);
nor U2484 (N_2484,N_2434,N_2404);
and U2485 (N_2485,N_2455,N_2407);
xnor U2486 (N_2486,N_2432,N_2409);
and U2487 (N_2487,N_2454,N_2419);
nand U2488 (N_2488,N_2457,N_2433);
nor U2489 (N_2489,N_2449,N_2431);
or U2490 (N_2490,N_2443,N_2410);
or U2491 (N_2491,N_2404,N_2423);
or U2492 (N_2492,N_2440,N_2437);
or U2493 (N_2493,N_2426,N_2403);
or U2494 (N_2494,N_2440,N_2438);
or U2495 (N_2495,N_2406,N_2448);
nor U2496 (N_2496,N_2402,N_2411);
xnor U2497 (N_2497,N_2450,N_2430);
or U2498 (N_2498,N_2419,N_2427);
and U2499 (N_2499,N_2457,N_2446);
and U2500 (N_2500,N_2446,N_2443);
nand U2501 (N_2501,N_2449,N_2410);
nand U2502 (N_2502,N_2457,N_2431);
nor U2503 (N_2503,N_2448,N_2400);
xnor U2504 (N_2504,N_2403,N_2457);
or U2505 (N_2505,N_2421,N_2418);
nand U2506 (N_2506,N_2422,N_2436);
xor U2507 (N_2507,N_2408,N_2444);
or U2508 (N_2508,N_2454,N_2437);
nor U2509 (N_2509,N_2449,N_2424);
xor U2510 (N_2510,N_2412,N_2434);
nand U2511 (N_2511,N_2416,N_2430);
or U2512 (N_2512,N_2410,N_2441);
nand U2513 (N_2513,N_2425,N_2432);
and U2514 (N_2514,N_2403,N_2453);
and U2515 (N_2515,N_2413,N_2426);
nand U2516 (N_2516,N_2459,N_2427);
and U2517 (N_2517,N_2437,N_2459);
and U2518 (N_2518,N_2458,N_2424);
nand U2519 (N_2519,N_2429,N_2432);
and U2520 (N_2520,N_2495,N_2501);
nand U2521 (N_2521,N_2510,N_2514);
nand U2522 (N_2522,N_2487,N_2498);
nand U2523 (N_2523,N_2463,N_2468);
and U2524 (N_2524,N_2462,N_2517);
or U2525 (N_2525,N_2465,N_2482);
xnor U2526 (N_2526,N_2489,N_2467);
nor U2527 (N_2527,N_2483,N_2488);
nand U2528 (N_2528,N_2479,N_2506);
or U2529 (N_2529,N_2518,N_2478);
nand U2530 (N_2530,N_2466,N_2475);
xnor U2531 (N_2531,N_2471,N_2490);
or U2532 (N_2532,N_2507,N_2473);
xor U2533 (N_2533,N_2516,N_2491);
and U2534 (N_2534,N_2484,N_2509);
and U2535 (N_2535,N_2499,N_2476);
or U2536 (N_2536,N_2515,N_2481);
or U2537 (N_2537,N_2461,N_2474);
xor U2538 (N_2538,N_2519,N_2511);
and U2539 (N_2539,N_2500,N_2494);
nand U2540 (N_2540,N_2464,N_2503);
and U2541 (N_2541,N_2460,N_2486);
xor U2542 (N_2542,N_2480,N_2477);
and U2543 (N_2543,N_2502,N_2497);
nand U2544 (N_2544,N_2485,N_2512);
xnor U2545 (N_2545,N_2504,N_2469);
nor U2546 (N_2546,N_2493,N_2472);
or U2547 (N_2547,N_2505,N_2508);
and U2548 (N_2548,N_2513,N_2470);
nor U2549 (N_2549,N_2496,N_2492);
nor U2550 (N_2550,N_2518,N_2471);
nor U2551 (N_2551,N_2463,N_2489);
and U2552 (N_2552,N_2487,N_2510);
and U2553 (N_2553,N_2510,N_2493);
nand U2554 (N_2554,N_2471,N_2467);
and U2555 (N_2555,N_2487,N_2464);
nor U2556 (N_2556,N_2472,N_2510);
nor U2557 (N_2557,N_2480,N_2501);
and U2558 (N_2558,N_2517,N_2496);
nor U2559 (N_2559,N_2471,N_2460);
xor U2560 (N_2560,N_2508,N_2517);
nor U2561 (N_2561,N_2487,N_2476);
nand U2562 (N_2562,N_2493,N_2501);
and U2563 (N_2563,N_2465,N_2509);
nand U2564 (N_2564,N_2497,N_2493);
nor U2565 (N_2565,N_2502,N_2461);
nor U2566 (N_2566,N_2503,N_2519);
and U2567 (N_2567,N_2492,N_2464);
or U2568 (N_2568,N_2468,N_2510);
or U2569 (N_2569,N_2500,N_2478);
xor U2570 (N_2570,N_2480,N_2464);
or U2571 (N_2571,N_2510,N_2494);
and U2572 (N_2572,N_2499,N_2484);
nor U2573 (N_2573,N_2472,N_2463);
and U2574 (N_2574,N_2476,N_2473);
nand U2575 (N_2575,N_2490,N_2511);
nor U2576 (N_2576,N_2482,N_2490);
and U2577 (N_2577,N_2462,N_2496);
nor U2578 (N_2578,N_2482,N_2473);
nand U2579 (N_2579,N_2478,N_2490);
and U2580 (N_2580,N_2565,N_2568);
xor U2581 (N_2581,N_2544,N_2556);
and U2582 (N_2582,N_2551,N_2554);
nor U2583 (N_2583,N_2530,N_2569);
or U2584 (N_2584,N_2559,N_2537);
xor U2585 (N_2585,N_2553,N_2532);
and U2586 (N_2586,N_2521,N_2577);
xor U2587 (N_2587,N_2538,N_2555);
or U2588 (N_2588,N_2541,N_2535);
nand U2589 (N_2589,N_2528,N_2549);
or U2590 (N_2590,N_2520,N_2552);
xnor U2591 (N_2591,N_2562,N_2546);
xnor U2592 (N_2592,N_2540,N_2523);
nand U2593 (N_2593,N_2579,N_2527);
xnor U2594 (N_2594,N_2533,N_2566);
nand U2595 (N_2595,N_2567,N_2563);
xor U2596 (N_2596,N_2531,N_2560);
or U2597 (N_2597,N_2574,N_2561);
or U2598 (N_2598,N_2529,N_2570);
and U2599 (N_2599,N_2526,N_2543);
and U2600 (N_2600,N_2542,N_2547);
nand U2601 (N_2601,N_2572,N_2522);
nand U2602 (N_2602,N_2578,N_2545);
nor U2603 (N_2603,N_2524,N_2557);
xnor U2604 (N_2604,N_2573,N_2575);
xnor U2605 (N_2605,N_2548,N_2571);
nor U2606 (N_2606,N_2536,N_2525);
nor U2607 (N_2607,N_2576,N_2534);
nor U2608 (N_2608,N_2558,N_2564);
or U2609 (N_2609,N_2550,N_2539);
and U2610 (N_2610,N_2544,N_2549);
and U2611 (N_2611,N_2556,N_2558);
nor U2612 (N_2612,N_2564,N_2528);
and U2613 (N_2613,N_2545,N_2543);
nor U2614 (N_2614,N_2575,N_2546);
and U2615 (N_2615,N_2544,N_2560);
nor U2616 (N_2616,N_2543,N_2555);
and U2617 (N_2617,N_2553,N_2566);
and U2618 (N_2618,N_2520,N_2575);
nand U2619 (N_2619,N_2526,N_2560);
nor U2620 (N_2620,N_2534,N_2538);
or U2621 (N_2621,N_2554,N_2542);
xor U2622 (N_2622,N_2566,N_2540);
or U2623 (N_2623,N_2570,N_2560);
nor U2624 (N_2624,N_2562,N_2539);
and U2625 (N_2625,N_2576,N_2578);
xor U2626 (N_2626,N_2559,N_2536);
xnor U2627 (N_2627,N_2540,N_2538);
or U2628 (N_2628,N_2579,N_2525);
and U2629 (N_2629,N_2549,N_2556);
and U2630 (N_2630,N_2558,N_2541);
and U2631 (N_2631,N_2520,N_2565);
or U2632 (N_2632,N_2526,N_2545);
or U2633 (N_2633,N_2532,N_2577);
nor U2634 (N_2634,N_2569,N_2556);
nor U2635 (N_2635,N_2561,N_2526);
nor U2636 (N_2636,N_2543,N_2567);
xor U2637 (N_2637,N_2527,N_2564);
and U2638 (N_2638,N_2569,N_2561);
nor U2639 (N_2639,N_2572,N_2576);
nand U2640 (N_2640,N_2634,N_2590);
nor U2641 (N_2641,N_2622,N_2591);
or U2642 (N_2642,N_2633,N_2615);
and U2643 (N_2643,N_2620,N_2621);
nand U2644 (N_2644,N_2580,N_2635);
xor U2645 (N_2645,N_2587,N_2585);
xor U2646 (N_2646,N_2628,N_2589);
and U2647 (N_2647,N_2626,N_2627);
or U2648 (N_2648,N_2602,N_2632);
nor U2649 (N_2649,N_2618,N_2593);
and U2650 (N_2650,N_2639,N_2614);
nor U2651 (N_2651,N_2595,N_2583);
and U2652 (N_2652,N_2631,N_2599);
nor U2653 (N_2653,N_2616,N_2596);
xor U2654 (N_2654,N_2609,N_2598);
or U2655 (N_2655,N_2588,N_2610);
nor U2656 (N_2656,N_2581,N_2600);
nor U2657 (N_2657,N_2636,N_2617);
or U2658 (N_2658,N_2605,N_2612);
xor U2659 (N_2659,N_2584,N_2629);
and U2660 (N_2660,N_2638,N_2586);
nor U2661 (N_2661,N_2604,N_2619);
nor U2662 (N_2662,N_2594,N_2597);
nand U2663 (N_2663,N_2601,N_2624);
and U2664 (N_2664,N_2630,N_2608);
or U2665 (N_2665,N_2625,N_2606);
and U2666 (N_2666,N_2582,N_2623);
xnor U2667 (N_2667,N_2603,N_2637);
nor U2668 (N_2668,N_2613,N_2611);
or U2669 (N_2669,N_2592,N_2607);
or U2670 (N_2670,N_2608,N_2635);
nand U2671 (N_2671,N_2598,N_2610);
and U2672 (N_2672,N_2609,N_2608);
xnor U2673 (N_2673,N_2633,N_2621);
nor U2674 (N_2674,N_2589,N_2622);
and U2675 (N_2675,N_2586,N_2603);
nor U2676 (N_2676,N_2613,N_2634);
nor U2677 (N_2677,N_2610,N_2602);
nor U2678 (N_2678,N_2632,N_2621);
nand U2679 (N_2679,N_2636,N_2600);
or U2680 (N_2680,N_2611,N_2584);
xor U2681 (N_2681,N_2581,N_2617);
or U2682 (N_2682,N_2635,N_2588);
nor U2683 (N_2683,N_2619,N_2614);
or U2684 (N_2684,N_2612,N_2582);
nor U2685 (N_2685,N_2585,N_2626);
xor U2686 (N_2686,N_2639,N_2594);
and U2687 (N_2687,N_2603,N_2613);
nand U2688 (N_2688,N_2622,N_2613);
xor U2689 (N_2689,N_2588,N_2626);
or U2690 (N_2690,N_2601,N_2607);
xnor U2691 (N_2691,N_2588,N_2591);
nand U2692 (N_2692,N_2617,N_2612);
xor U2693 (N_2693,N_2613,N_2638);
xnor U2694 (N_2694,N_2612,N_2631);
nor U2695 (N_2695,N_2619,N_2596);
and U2696 (N_2696,N_2587,N_2604);
nor U2697 (N_2697,N_2605,N_2582);
or U2698 (N_2698,N_2616,N_2604);
nand U2699 (N_2699,N_2629,N_2594);
xor U2700 (N_2700,N_2642,N_2669);
and U2701 (N_2701,N_2663,N_2681);
xnor U2702 (N_2702,N_2696,N_2684);
and U2703 (N_2703,N_2689,N_2646);
xor U2704 (N_2704,N_2697,N_2673);
or U2705 (N_2705,N_2698,N_2658);
xnor U2706 (N_2706,N_2693,N_2676);
nand U2707 (N_2707,N_2644,N_2692);
nor U2708 (N_2708,N_2665,N_2672);
nand U2709 (N_2709,N_2662,N_2666);
nand U2710 (N_2710,N_2647,N_2641);
or U2711 (N_2711,N_2640,N_2649);
or U2712 (N_2712,N_2683,N_2687);
nand U2713 (N_2713,N_2685,N_2680);
nand U2714 (N_2714,N_2699,N_2654);
xnor U2715 (N_2715,N_2688,N_2650);
nand U2716 (N_2716,N_2670,N_2668);
or U2717 (N_2717,N_2677,N_2682);
or U2718 (N_2718,N_2694,N_2659);
xor U2719 (N_2719,N_2674,N_2657);
and U2720 (N_2720,N_2691,N_2660);
nor U2721 (N_2721,N_2679,N_2675);
and U2722 (N_2722,N_2655,N_2667);
nor U2723 (N_2723,N_2643,N_2648);
nor U2724 (N_2724,N_2664,N_2686);
or U2725 (N_2725,N_2653,N_2656);
nand U2726 (N_2726,N_2661,N_2651);
or U2727 (N_2727,N_2678,N_2671);
xnor U2728 (N_2728,N_2695,N_2652);
or U2729 (N_2729,N_2645,N_2690);
nand U2730 (N_2730,N_2643,N_2641);
and U2731 (N_2731,N_2647,N_2655);
and U2732 (N_2732,N_2662,N_2663);
nor U2733 (N_2733,N_2672,N_2689);
and U2734 (N_2734,N_2684,N_2669);
xnor U2735 (N_2735,N_2696,N_2691);
xor U2736 (N_2736,N_2666,N_2654);
xor U2737 (N_2737,N_2684,N_2643);
and U2738 (N_2738,N_2650,N_2652);
nor U2739 (N_2739,N_2659,N_2670);
xnor U2740 (N_2740,N_2682,N_2679);
and U2741 (N_2741,N_2674,N_2663);
or U2742 (N_2742,N_2662,N_2683);
xor U2743 (N_2743,N_2671,N_2690);
nand U2744 (N_2744,N_2671,N_2660);
xnor U2745 (N_2745,N_2654,N_2690);
nand U2746 (N_2746,N_2684,N_2665);
or U2747 (N_2747,N_2640,N_2683);
and U2748 (N_2748,N_2660,N_2695);
xor U2749 (N_2749,N_2642,N_2695);
xor U2750 (N_2750,N_2682,N_2643);
nand U2751 (N_2751,N_2696,N_2690);
xor U2752 (N_2752,N_2684,N_2648);
nor U2753 (N_2753,N_2693,N_2643);
nand U2754 (N_2754,N_2699,N_2696);
or U2755 (N_2755,N_2652,N_2653);
nand U2756 (N_2756,N_2655,N_2699);
xnor U2757 (N_2757,N_2682,N_2657);
xor U2758 (N_2758,N_2670,N_2677);
and U2759 (N_2759,N_2660,N_2659);
nand U2760 (N_2760,N_2703,N_2705);
nand U2761 (N_2761,N_2718,N_2729);
and U2762 (N_2762,N_2734,N_2717);
xnor U2763 (N_2763,N_2730,N_2736);
nor U2764 (N_2764,N_2709,N_2723);
xnor U2765 (N_2765,N_2716,N_2724);
xor U2766 (N_2766,N_2750,N_2733);
or U2767 (N_2767,N_2756,N_2713);
nand U2768 (N_2768,N_2735,N_2728);
nand U2769 (N_2769,N_2720,N_2753);
or U2770 (N_2770,N_2749,N_2702);
nand U2771 (N_2771,N_2711,N_2712);
xor U2772 (N_2772,N_2743,N_2751);
and U2773 (N_2773,N_2744,N_2731);
and U2774 (N_2774,N_2722,N_2701);
and U2775 (N_2775,N_2745,N_2732);
nor U2776 (N_2776,N_2738,N_2739);
or U2777 (N_2777,N_2727,N_2748);
nand U2778 (N_2778,N_2746,N_2742);
xnor U2779 (N_2779,N_2747,N_2707);
nand U2780 (N_2780,N_2726,N_2752);
xor U2781 (N_2781,N_2715,N_2719);
xor U2782 (N_2782,N_2754,N_2700);
or U2783 (N_2783,N_2725,N_2741);
and U2784 (N_2784,N_2714,N_2708);
and U2785 (N_2785,N_2721,N_2759);
and U2786 (N_2786,N_2757,N_2704);
nor U2787 (N_2787,N_2740,N_2737);
xor U2788 (N_2788,N_2758,N_2710);
and U2789 (N_2789,N_2755,N_2706);
and U2790 (N_2790,N_2742,N_2757);
nand U2791 (N_2791,N_2750,N_2713);
xor U2792 (N_2792,N_2700,N_2725);
and U2793 (N_2793,N_2759,N_2718);
and U2794 (N_2794,N_2758,N_2744);
nand U2795 (N_2795,N_2743,N_2740);
or U2796 (N_2796,N_2752,N_2744);
or U2797 (N_2797,N_2724,N_2730);
nand U2798 (N_2798,N_2725,N_2720);
and U2799 (N_2799,N_2742,N_2758);
nand U2800 (N_2800,N_2726,N_2715);
xnor U2801 (N_2801,N_2706,N_2742);
nor U2802 (N_2802,N_2759,N_2728);
nor U2803 (N_2803,N_2721,N_2700);
or U2804 (N_2804,N_2712,N_2730);
nor U2805 (N_2805,N_2713,N_2748);
or U2806 (N_2806,N_2740,N_2727);
xnor U2807 (N_2807,N_2737,N_2703);
nor U2808 (N_2808,N_2711,N_2729);
or U2809 (N_2809,N_2701,N_2721);
nor U2810 (N_2810,N_2717,N_2720);
nand U2811 (N_2811,N_2734,N_2722);
or U2812 (N_2812,N_2746,N_2721);
and U2813 (N_2813,N_2754,N_2737);
xnor U2814 (N_2814,N_2751,N_2727);
nand U2815 (N_2815,N_2702,N_2733);
or U2816 (N_2816,N_2736,N_2740);
xor U2817 (N_2817,N_2722,N_2752);
and U2818 (N_2818,N_2738,N_2708);
xnor U2819 (N_2819,N_2737,N_2719);
nand U2820 (N_2820,N_2796,N_2799);
xnor U2821 (N_2821,N_2781,N_2818);
xnor U2822 (N_2822,N_2786,N_2813);
nand U2823 (N_2823,N_2762,N_2817);
nand U2824 (N_2824,N_2780,N_2794);
nor U2825 (N_2825,N_2815,N_2767);
and U2826 (N_2826,N_2782,N_2787);
and U2827 (N_2827,N_2788,N_2765);
or U2828 (N_2828,N_2777,N_2790);
or U2829 (N_2829,N_2811,N_2795);
nand U2830 (N_2830,N_2792,N_2806);
or U2831 (N_2831,N_2771,N_2760);
nand U2832 (N_2832,N_2785,N_2778);
xor U2833 (N_2833,N_2791,N_2779);
and U2834 (N_2834,N_2766,N_2768);
nand U2835 (N_2835,N_2772,N_2804);
nor U2836 (N_2836,N_2763,N_2801);
xnor U2837 (N_2837,N_2784,N_2800);
xor U2838 (N_2838,N_2814,N_2802);
and U2839 (N_2839,N_2776,N_2808);
nor U2840 (N_2840,N_2809,N_2810);
nand U2841 (N_2841,N_2774,N_2803);
nor U2842 (N_2842,N_2773,N_2797);
xor U2843 (N_2843,N_2812,N_2793);
nor U2844 (N_2844,N_2816,N_2789);
and U2845 (N_2845,N_2819,N_2807);
nand U2846 (N_2846,N_2761,N_2783);
xnor U2847 (N_2847,N_2805,N_2775);
and U2848 (N_2848,N_2798,N_2769);
nand U2849 (N_2849,N_2770,N_2764);
xnor U2850 (N_2850,N_2776,N_2777);
nand U2851 (N_2851,N_2778,N_2792);
nor U2852 (N_2852,N_2766,N_2772);
xor U2853 (N_2853,N_2810,N_2798);
or U2854 (N_2854,N_2795,N_2766);
xor U2855 (N_2855,N_2803,N_2782);
or U2856 (N_2856,N_2786,N_2799);
nor U2857 (N_2857,N_2811,N_2819);
or U2858 (N_2858,N_2782,N_2814);
nor U2859 (N_2859,N_2786,N_2776);
and U2860 (N_2860,N_2818,N_2786);
or U2861 (N_2861,N_2782,N_2796);
xor U2862 (N_2862,N_2810,N_2812);
nand U2863 (N_2863,N_2796,N_2792);
xnor U2864 (N_2864,N_2761,N_2816);
and U2865 (N_2865,N_2819,N_2813);
xor U2866 (N_2866,N_2772,N_2813);
xnor U2867 (N_2867,N_2787,N_2780);
nor U2868 (N_2868,N_2808,N_2793);
or U2869 (N_2869,N_2763,N_2767);
nand U2870 (N_2870,N_2760,N_2786);
nand U2871 (N_2871,N_2764,N_2808);
nor U2872 (N_2872,N_2766,N_2792);
nor U2873 (N_2873,N_2814,N_2768);
xor U2874 (N_2874,N_2790,N_2817);
nand U2875 (N_2875,N_2763,N_2819);
nor U2876 (N_2876,N_2814,N_2769);
nand U2877 (N_2877,N_2779,N_2771);
and U2878 (N_2878,N_2793,N_2784);
and U2879 (N_2879,N_2802,N_2764);
and U2880 (N_2880,N_2824,N_2869);
xnor U2881 (N_2881,N_2845,N_2835);
xnor U2882 (N_2882,N_2828,N_2820);
or U2883 (N_2883,N_2844,N_2847);
and U2884 (N_2884,N_2878,N_2857);
nand U2885 (N_2885,N_2825,N_2849);
xnor U2886 (N_2886,N_2863,N_2826);
or U2887 (N_2887,N_2842,N_2850);
or U2888 (N_2888,N_2822,N_2831);
or U2889 (N_2889,N_2823,N_2859);
and U2890 (N_2890,N_2853,N_2837);
and U2891 (N_2891,N_2855,N_2868);
or U2892 (N_2892,N_2867,N_2866);
and U2893 (N_2893,N_2838,N_2846);
or U2894 (N_2894,N_2854,N_2860);
or U2895 (N_2895,N_2875,N_2843);
nand U2896 (N_2896,N_2879,N_2832);
or U2897 (N_2897,N_2852,N_2877);
nand U2898 (N_2898,N_2851,N_2861);
nand U2899 (N_2899,N_2873,N_2862);
xnor U2900 (N_2900,N_2865,N_2830);
and U2901 (N_2901,N_2856,N_2827);
nand U2902 (N_2902,N_2858,N_2872);
or U2903 (N_2903,N_2829,N_2870);
and U2904 (N_2904,N_2836,N_2833);
or U2905 (N_2905,N_2821,N_2848);
xnor U2906 (N_2906,N_2840,N_2864);
and U2907 (N_2907,N_2876,N_2834);
nand U2908 (N_2908,N_2841,N_2839);
and U2909 (N_2909,N_2871,N_2874);
and U2910 (N_2910,N_2842,N_2861);
nand U2911 (N_2911,N_2842,N_2823);
or U2912 (N_2912,N_2820,N_2864);
xor U2913 (N_2913,N_2858,N_2874);
xnor U2914 (N_2914,N_2854,N_2874);
and U2915 (N_2915,N_2829,N_2871);
nor U2916 (N_2916,N_2827,N_2821);
nand U2917 (N_2917,N_2825,N_2875);
nor U2918 (N_2918,N_2823,N_2824);
nand U2919 (N_2919,N_2877,N_2875);
nor U2920 (N_2920,N_2837,N_2830);
and U2921 (N_2921,N_2846,N_2857);
or U2922 (N_2922,N_2876,N_2841);
xor U2923 (N_2923,N_2862,N_2840);
or U2924 (N_2924,N_2845,N_2873);
or U2925 (N_2925,N_2877,N_2839);
nor U2926 (N_2926,N_2838,N_2859);
nand U2927 (N_2927,N_2871,N_2832);
or U2928 (N_2928,N_2866,N_2859);
and U2929 (N_2929,N_2878,N_2845);
xor U2930 (N_2930,N_2844,N_2871);
nor U2931 (N_2931,N_2831,N_2859);
xor U2932 (N_2932,N_2875,N_2855);
nand U2933 (N_2933,N_2874,N_2872);
or U2934 (N_2934,N_2876,N_2857);
or U2935 (N_2935,N_2829,N_2856);
and U2936 (N_2936,N_2850,N_2863);
and U2937 (N_2937,N_2872,N_2846);
nor U2938 (N_2938,N_2844,N_2865);
nor U2939 (N_2939,N_2851,N_2843);
xor U2940 (N_2940,N_2895,N_2886);
and U2941 (N_2941,N_2891,N_2901);
nand U2942 (N_2942,N_2912,N_2904);
nand U2943 (N_2943,N_2897,N_2902);
and U2944 (N_2944,N_2924,N_2898);
xnor U2945 (N_2945,N_2884,N_2919);
nor U2946 (N_2946,N_2909,N_2908);
or U2947 (N_2947,N_2893,N_2910);
and U2948 (N_2948,N_2915,N_2922);
or U2949 (N_2949,N_2934,N_2885);
nand U2950 (N_2950,N_2892,N_2889);
or U2951 (N_2951,N_2929,N_2887);
and U2952 (N_2952,N_2916,N_2894);
or U2953 (N_2953,N_2931,N_2907);
xnor U2954 (N_2954,N_2882,N_2930);
or U2955 (N_2955,N_2938,N_2900);
nor U2956 (N_2956,N_2936,N_2903);
and U2957 (N_2957,N_2896,N_2928);
or U2958 (N_2958,N_2935,N_2906);
nor U2959 (N_2959,N_2888,N_2905);
or U2960 (N_2960,N_2939,N_2925);
nor U2961 (N_2961,N_2881,N_2890);
xor U2962 (N_2962,N_2927,N_2880);
xnor U2963 (N_2963,N_2923,N_2883);
nand U2964 (N_2964,N_2932,N_2914);
xnor U2965 (N_2965,N_2920,N_2933);
nor U2966 (N_2966,N_2899,N_2911);
and U2967 (N_2967,N_2921,N_2926);
xor U2968 (N_2968,N_2917,N_2937);
and U2969 (N_2969,N_2918,N_2913);
and U2970 (N_2970,N_2915,N_2930);
nor U2971 (N_2971,N_2932,N_2880);
nor U2972 (N_2972,N_2892,N_2922);
xnor U2973 (N_2973,N_2888,N_2936);
or U2974 (N_2974,N_2906,N_2898);
xor U2975 (N_2975,N_2893,N_2909);
or U2976 (N_2976,N_2933,N_2932);
and U2977 (N_2977,N_2930,N_2904);
nand U2978 (N_2978,N_2931,N_2906);
and U2979 (N_2979,N_2930,N_2896);
xor U2980 (N_2980,N_2883,N_2936);
and U2981 (N_2981,N_2913,N_2892);
and U2982 (N_2982,N_2913,N_2925);
xor U2983 (N_2983,N_2937,N_2885);
nor U2984 (N_2984,N_2930,N_2912);
and U2985 (N_2985,N_2899,N_2935);
nand U2986 (N_2986,N_2899,N_2898);
xor U2987 (N_2987,N_2911,N_2908);
nand U2988 (N_2988,N_2906,N_2907);
nor U2989 (N_2989,N_2928,N_2914);
and U2990 (N_2990,N_2883,N_2916);
xnor U2991 (N_2991,N_2886,N_2925);
nand U2992 (N_2992,N_2903,N_2901);
nand U2993 (N_2993,N_2896,N_2918);
nor U2994 (N_2994,N_2927,N_2909);
and U2995 (N_2995,N_2931,N_2939);
xor U2996 (N_2996,N_2937,N_2933);
and U2997 (N_2997,N_2895,N_2907);
and U2998 (N_2998,N_2885,N_2939);
nor U2999 (N_2999,N_2935,N_2894);
and UO_0 (O_0,N_2956,N_2976);
nand UO_1 (O_1,N_2969,N_2985);
xor UO_2 (O_2,N_2981,N_2957);
nand UO_3 (O_3,N_2973,N_2979);
or UO_4 (O_4,N_2994,N_2941);
nor UO_5 (O_5,N_2967,N_2991);
nand UO_6 (O_6,N_2945,N_2983);
xnor UO_7 (O_7,N_2955,N_2963);
and UO_8 (O_8,N_2964,N_2996);
nand UO_9 (O_9,N_2975,N_2950);
xnor UO_10 (O_10,N_2947,N_2953);
or UO_11 (O_11,N_2988,N_2968);
and UO_12 (O_12,N_2962,N_2949);
nor UO_13 (O_13,N_2954,N_2970);
nor UO_14 (O_14,N_2997,N_2952);
or UO_15 (O_15,N_2974,N_2986);
nand UO_16 (O_16,N_2984,N_2971);
nand UO_17 (O_17,N_2999,N_2965);
nor UO_18 (O_18,N_2982,N_2992);
xnor UO_19 (O_19,N_2972,N_2959);
xnor UO_20 (O_20,N_2977,N_2995);
nand UO_21 (O_21,N_2944,N_2966);
xor UO_22 (O_22,N_2989,N_2948);
xnor UO_23 (O_23,N_2958,N_2961);
nor UO_24 (O_24,N_2951,N_2998);
and UO_25 (O_25,N_2987,N_2978);
and UO_26 (O_26,N_2946,N_2980);
nand UO_27 (O_27,N_2990,N_2960);
nor UO_28 (O_28,N_2993,N_2943);
or UO_29 (O_29,N_2940,N_2942);
and UO_30 (O_30,N_2982,N_2946);
and UO_31 (O_31,N_2976,N_2952);
nand UO_32 (O_32,N_2943,N_2991);
xnor UO_33 (O_33,N_2995,N_2978);
and UO_34 (O_34,N_2957,N_2990);
nand UO_35 (O_35,N_2978,N_2991);
and UO_36 (O_36,N_2949,N_2990);
nand UO_37 (O_37,N_2954,N_2992);
and UO_38 (O_38,N_2953,N_2968);
nor UO_39 (O_39,N_2982,N_2958);
nand UO_40 (O_40,N_2977,N_2960);
and UO_41 (O_41,N_2952,N_2995);
xor UO_42 (O_42,N_2941,N_2971);
or UO_43 (O_43,N_2971,N_2956);
and UO_44 (O_44,N_2960,N_2953);
xor UO_45 (O_45,N_2948,N_2967);
and UO_46 (O_46,N_2984,N_2988);
nor UO_47 (O_47,N_2951,N_2973);
or UO_48 (O_48,N_2945,N_2973);
xnor UO_49 (O_49,N_2987,N_2942);
xnor UO_50 (O_50,N_2963,N_2978);
and UO_51 (O_51,N_2945,N_2976);
nor UO_52 (O_52,N_2944,N_2958);
nand UO_53 (O_53,N_2959,N_2973);
nand UO_54 (O_54,N_2981,N_2973);
nor UO_55 (O_55,N_2976,N_2948);
nand UO_56 (O_56,N_2991,N_2949);
xnor UO_57 (O_57,N_2994,N_2988);
nand UO_58 (O_58,N_2998,N_2941);
or UO_59 (O_59,N_2949,N_2964);
and UO_60 (O_60,N_2990,N_2955);
xnor UO_61 (O_61,N_2957,N_2962);
nand UO_62 (O_62,N_2998,N_2961);
and UO_63 (O_63,N_2955,N_2998);
nand UO_64 (O_64,N_2970,N_2996);
xor UO_65 (O_65,N_2953,N_2977);
nand UO_66 (O_66,N_2974,N_2961);
and UO_67 (O_67,N_2979,N_2950);
and UO_68 (O_68,N_2951,N_2964);
nor UO_69 (O_69,N_2981,N_2968);
or UO_70 (O_70,N_2950,N_2942);
nor UO_71 (O_71,N_2960,N_2958);
nor UO_72 (O_72,N_2993,N_2944);
nor UO_73 (O_73,N_2953,N_2993);
xor UO_74 (O_74,N_2972,N_2996);
or UO_75 (O_75,N_2946,N_2979);
xnor UO_76 (O_76,N_2973,N_2946);
xnor UO_77 (O_77,N_2952,N_2980);
and UO_78 (O_78,N_2944,N_2996);
and UO_79 (O_79,N_2967,N_2946);
nand UO_80 (O_80,N_2977,N_2988);
nor UO_81 (O_81,N_2984,N_2975);
and UO_82 (O_82,N_2989,N_2997);
nor UO_83 (O_83,N_2972,N_2998);
and UO_84 (O_84,N_2986,N_2941);
nand UO_85 (O_85,N_2986,N_2981);
xnor UO_86 (O_86,N_2946,N_2985);
xnor UO_87 (O_87,N_2946,N_2959);
and UO_88 (O_88,N_2994,N_2997);
nor UO_89 (O_89,N_2993,N_2987);
nand UO_90 (O_90,N_2984,N_2995);
xnor UO_91 (O_91,N_2999,N_2958);
and UO_92 (O_92,N_2978,N_2976);
xnor UO_93 (O_93,N_2972,N_2982);
xor UO_94 (O_94,N_2951,N_2953);
nand UO_95 (O_95,N_2969,N_2959);
nand UO_96 (O_96,N_2987,N_2983);
and UO_97 (O_97,N_2949,N_2980);
or UO_98 (O_98,N_2986,N_2963);
xor UO_99 (O_99,N_2990,N_2956);
nand UO_100 (O_100,N_2959,N_2960);
nor UO_101 (O_101,N_2969,N_2965);
nor UO_102 (O_102,N_2957,N_2995);
or UO_103 (O_103,N_2977,N_2974);
or UO_104 (O_104,N_2980,N_2996);
or UO_105 (O_105,N_2954,N_2989);
and UO_106 (O_106,N_2979,N_2954);
and UO_107 (O_107,N_2950,N_2981);
nand UO_108 (O_108,N_2980,N_2991);
nand UO_109 (O_109,N_2990,N_2971);
nand UO_110 (O_110,N_2944,N_2986);
xor UO_111 (O_111,N_2962,N_2987);
nor UO_112 (O_112,N_2994,N_2978);
and UO_113 (O_113,N_2956,N_2970);
or UO_114 (O_114,N_2967,N_2945);
nand UO_115 (O_115,N_2976,N_2941);
xor UO_116 (O_116,N_2950,N_2962);
xnor UO_117 (O_117,N_2976,N_2967);
and UO_118 (O_118,N_2953,N_2990);
nand UO_119 (O_119,N_2993,N_2998);
nor UO_120 (O_120,N_2970,N_2983);
and UO_121 (O_121,N_2967,N_2972);
and UO_122 (O_122,N_2944,N_2973);
xnor UO_123 (O_123,N_2964,N_2981);
nand UO_124 (O_124,N_2966,N_2985);
nand UO_125 (O_125,N_2996,N_2990);
xor UO_126 (O_126,N_2964,N_2973);
or UO_127 (O_127,N_2970,N_2999);
and UO_128 (O_128,N_2998,N_2964);
nand UO_129 (O_129,N_2951,N_2999);
xnor UO_130 (O_130,N_2947,N_2988);
xor UO_131 (O_131,N_2970,N_2959);
nand UO_132 (O_132,N_2949,N_2944);
or UO_133 (O_133,N_2943,N_2990);
and UO_134 (O_134,N_2979,N_2956);
xnor UO_135 (O_135,N_2952,N_2949);
and UO_136 (O_136,N_2956,N_2987);
or UO_137 (O_137,N_2976,N_2975);
and UO_138 (O_138,N_2956,N_2951);
or UO_139 (O_139,N_2952,N_2974);
and UO_140 (O_140,N_2955,N_2943);
or UO_141 (O_141,N_2940,N_2987);
xnor UO_142 (O_142,N_2949,N_2950);
nor UO_143 (O_143,N_2947,N_2971);
nor UO_144 (O_144,N_2999,N_2973);
or UO_145 (O_145,N_2956,N_2978);
xnor UO_146 (O_146,N_2973,N_2984);
or UO_147 (O_147,N_2982,N_2948);
or UO_148 (O_148,N_2978,N_2960);
xor UO_149 (O_149,N_2991,N_2965);
and UO_150 (O_150,N_2980,N_2966);
xor UO_151 (O_151,N_2943,N_2994);
nand UO_152 (O_152,N_2941,N_2982);
and UO_153 (O_153,N_2986,N_2984);
or UO_154 (O_154,N_2956,N_2949);
nor UO_155 (O_155,N_2962,N_2947);
nor UO_156 (O_156,N_2947,N_2984);
xnor UO_157 (O_157,N_2949,N_2968);
or UO_158 (O_158,N_2945,N_2943);
xnor UO_159 (O_159,N_2989,N_2996);
or UO_160 (O_160,N_2966,N_2982);
nand UO_161 (O_161,N_2980,N_2957);
and UO_162 (O_162,N_2986,N_2989);
or UO_163 (O_163,N_2972,N_2957);
and UO_164 (O_164,N_2977,N_2964);
and UO_165 (O_165,N_2974,N_2992);
xor UO_166 (O_166,N_2988,N_2948);
or UO_167 (O_167,N_2996,N_2954);
or UO_168 (O_168,N_2944,N_2972);
nor UO_169 (O_169,N_2971,N_2986);
and UO_170 (O_170,N_2949,N_2977);
and UO_171 (O_171,N_2953,N_2992);
and UO_172 (O_172,N_2987,N_2990);
and UO_173 (O_173,N_2984,N_2965);
xor UO_174 (O_174,N_2991,N_2945);
or UO_175 (O_175,N_2996,N_2950);
or UO_176 (O_176,N_2947,N_2957);
nor UO_177 (O_177,N_2996,N_2985);
nor UO_178 (O_178,N_2951,N_2995);
xor UO_179 (O_179,N_2976,N_2982);
nor UO_180 (O_180,N_2980,N_2959);
xor UO_181 (O_181,N_2960,N_2993);
and UO_182 (O_182,N_2947,N_2961);
nand UO_183 (O_183,N_2984,N_2962);
nand UO_184 (O_184,N_2991,N_2969);
and UO_185 (O_185,N_2955,N_2956);
xnor UO_186 (O_186,N_2965,N_2985);
and UO_187 (O_187,N_2973,N_2960);
and UO_188 (O_188,N_2956,N_2944);
nor UO_189 (O_189,N_2944,N_2990);
nand UO_190 (O_190,N_2994,N_2986);
nand UO_191 (O_191,N_2978,N_2997);
xnor UO_192 (O_192,N_2992,N_2969);
or UO_193 (O_193,N_2952,N_2964);
xnor UO_194 (O_194,N_2961,N_2976);
nand UO_195 (O_195,N_2950,N_2945);
and UO_196 (O_196,N_2961,N_2960);
or UO_197 (O_197,N_2940,N_2941);
xor UO_198 (O_198,N_2959,N_2977);
nor UO_199 (O_199,N_2958,N_2974);
nor UO_200 (O_200,N_2995,N_2993);
and UO_201 (O_201,N_2996,N_2981);
nor UO_202 (O_202,N_2983,N_2971);
nand UO_203 (O_203,N_2956,N_2965);
or UO_204 (O_204,N_2946,N_2995);
or UO_205 (O_205,N_2940,N_2956);
nand UO_206 (O_206,N_2949,N_2943);
nor UO_207 (O_207,N_2966,N_2952);
nand UO_208 (O_208,N_2946,N_2950);
nor UO_209 (O_209,N_2958,N_2946);
or UO_210 (O_210,N_2952,N_2999);
nor UO_211 (O_211,N_2978,N_2967);
nor UO_212 (O_212,N_2954,N_2949);
and UO_213 (O_213,N_2994,N_2968);
or UO_214 (O_214,N_2991,N_2995);
nor UO_215 (O_215,N_2995,N_2981);
and UO_216 (O_216,N_2988,N_2964);
or UO_217 (O_217,N_2943,N_2971);
xor UO_218 (O_218,N_2943,N_2941);
xor UO_219 (O_219,N_2948,N_2996);
and UO_220 (O_220,N_2974,N_2940);
nor UO_221 (O_221,N_2976,N_2993);
or UO_222 (O_222,N_2979,N_2983);
or UO_223 (O_223,N_2971,N_2961);
nand UO_224 (O_224,N_2997,N_2960);
and UO_225 (O_225,N_2966,N_2977);
xor UO_226 (O_226,N_2969,N_2996);
xor UO_227 (O_227,N_2940,N_2965);
xnor UO_228 (O_228,N_2972,N_2992);
or UO_229 (O_229,N_2965,N_2967);
xnor UO_230 (O_230,N_2994,N_2980);
nor UO_231 (O_231,N_2986,N_2943);
nor UO_232 (O_232,N_2974,N_2979);
and UO_233 (O_233,N_2980,N_2940);
nand UO_234 (O_234,N_2987,N_2953);
or UO_235 (O_235,N_2975,N_2983);
xor UO_236 (O_236,N_2947,N_2996);
xnor UO_237 (O_237,N_2991,N_2956);
or UO_238 (O_238,N_2953,N_2964);
or UO_239 (O_239,N_2982,N_2953);
nand UO_240 (O_240,N_2981,N_2959);
nand UO_241 (O_241,N_2954,N_2985);
nand UO_242 (O_242,N_2996,N_2956);
and UO_243 (O_243,N_2975,N_2996);
and UO_244 (O_244,N_2988,N_2981);
and UO_245 (O_245,N_2968,N_2962);
and UO_246 (O_246,N_2972,N_2979);
and UO_247 (O_247,N_2998,N_2947);
nor UO_248 (O_248,N_2975,N_2944);
nand UO_249 (O_249,N_2957,N_2965);
and UO_250 (O_250,N_2975,N_2993);
nand UO_251 (O_251,N_2986,N_2993);
nand UO_252 (O_252,N_2973,N_2942);
nand UO_253 (O_253,N_2989,N_2994);
nand UO_254 (O_254,N_2941,N_2967);
and UO_255 (O_255,N_2975,N_2999);
and UO_256 (O_256,N_2944,N_2967);
nor UO_257 (O_257,N_2965,N_2971);
and UO_258 (O_258,N_2963,N_2960);
and UO_259 (O_259,N_2985,N_2944);
xor UO_260 (O_260,N_2951,N_2942);
nor UO_261 (O_261,N_2986,N_2996);
xor UO_262 (O_262,N_2949,N_2974);
nand UO_263 (O_263,N_2940,N_2983);
nand UO_264 (O_264,N_2953,N_2999);
or UO_265 (O_265,N_2996,N_2999);
or UO_266 (O_266,N_2981,N_2991);
nor UO_267 (O_267,N_2973,N_2985);
nor UO_268 (O_268,N_2942,N_2972);
nand UO_269 (O_269,N_2991,N_2996);
and UO_270 (O_270,N_2989,N_2987);
xor UO_271 (O_271,N_2994,N_2987);
and UO_272 (O_272,N_2946,N_2968);
xor UO_273 (O_273,N_2947,N_2978);
nor UO_274 (O_274,N_2944,N_2978);
nor UO_275 (O_275,N_2975,N_2987);
and UO_276 (O_276,N_2995,N_2998);
xor UO_277 (O_277,N_2952,N_2958);
nor UO_278 (O_278,N_2966,N_2948);
nor UO_279 (O_279,N_2996,N_2951);
and UO_280 (O_280,N_2962,N_2983);
xor UO_281 (O_281,N_2960,N_2972);
and UO_282 (O_282,N_2940,N_2954);
and UO_283 (O_283,N_2971,N_2985);
nand UO_284 (O_284,N_2941,N_2970);
xor UO_285 (O_285,N_2988,N_2999);
xor UO_286 (O_286,N_2975,N_2953);
xnor UO_287 (O_287,N_2959,N_2958);
nand UO_288 (O_288,N_2962,N_2956);
or UO_289 (O_289,N_2946,N_2947);
and UO_290 (O_290,N_2980,N_2945);
xor UO_291 (O_291,N_2976,N_2957);
and UO_292 (O_292,N_2970,N_2957);
nand UO_293 (O_293,N_2953,N_2971);
xnor UO_294 (O_294,N_2945,N_2946);
or UO_295 (O_295,N_2996,N_2940);
nor UO_296 (O_296,N_2960,N_2983);
nand UO_297 (O_297,N_2964,N_2987);
and UO_298 (O_298,N_2978,N_2942);
nand UO_299 (O_299,N_2981,N_2961);
xor UO_300 (O_300,N_2985,N_2955);
and UO_301 (O_301,N_2955,N_2992);
nand UO_302 (O_302,N_2943,N_2980);
nand UO_303 (O_303,N_2940,N_2972);
or UO_304 (O_304,N_2982,N_2995);
nand UO_305 (O_305,N_2982,N_2981);
or UO_306 (O_306,N_2983,N_2995);
nand UO_307 (O_307,N_2984,N_2983);
or UO_308 (O_308,N_2996,N_2945);
nor UO_309 (O_309,N_2991,N_2984);
and UO_310 (O_310,N_2987,N_2958);
and UO_311 (O_311,N_2981,N_2969);
nand UO_312 (O_312,N_2992,N_2948);
nor UO_313 (O_313,N_2960,N_2951);
xor UO_314 (O_314,N_2981,N_2954);
nor UO_315 (O_315,N_2979,N_2998);
xor UO_316 (O_316,N_2983,N_2956);
xor UO_317 (O_317,N_2971,N_2989);
xor UO_318 (O_318,N_2981,N_2994);
nand UO_319 (O_319,N_2965,N_2989);
or UO_320 (O_320,N_2982,N_2994);
nand UO_321 (O_321,N_2970,N_2987);
nor UO_322 (O_322,N_2947,N_2990);
xor UO_323 (O_323,N_2956,N_2986);
nand UO_324 (O_324,N_2978,N_2962);
nand UO_325 (O_325,N_2977,N_2963);
or UO_326 (O_326,N_2994,N_2985);
or UO_327 (O_327,N_2970,N_2953);
xor UO_328 (O_328,N_2982,N_2985);
nand UO_329 (O_329,N_2957,N_2983);
or UO_330 (O_330,N_2999,N_2986);
or UO_331 (O_331,N_2992,N_2946);
xor UO_332 (O_332,N_2989,N_2993);
nand UO_333 (O_333,N_2944,N_2948);
nand UO_334 (O_334,N_2945,N_2940);
nand UO_335 (O_335,N_2946,N_2942);
xor UO_336 (O_336,N_2956,N_2959);
and UO_337 (O_337,N_2993,N_2961);
and UO_338 (O_338,N_2990,N_2963);
and UO_339 (O_339,N_2968,N_2975);
nand UO_340 (O_340,N_2961,N_2952);
xor UO_341 (O_341,N_2974,N_2959);
nand UO_342 (O_342,N_2990,N_2970);
xor UO_343 (O_343,N_2985,N_2989);
nor UO_344 (O_344,N_2949,N_2967);
nand UO_345 (O_345,N_2997,N_2962);
nand UO_346 (O_346,N_2989,N_2990);
and UO_347 (O_347,N_2978,N_2966);
or UO_348 (O_348,N_2957,N_2953);
nand UO_349 (O_349,N_2945,N_2969);
nor UO_350 (O_350,N_2946,N_2989);
xnor UO_351 (O_351,N_2950,N_2951);
nand UO_352 (O_352,N_2946,N_2970);
nor UO_353 (O_353,N_2955,N_2995);
xor UO_354 (O_354,N_2950,N_2957);
or UO_355 (O_355,N_2974,N_2960);
or UO_356 (O_356,N_2981,N_2958);
or UO_357 (O_357,N_2943,N_2967);
or UO_358 (O_358,N_2969,N_2966);
or UO_359 (O_359,N_2982,N_2989);
nor UO_360 (O_360,N_2960,N_2956);
or UO_361 (O_361,N_2990,N_2945);
nor UO_362 (O_362,N_2947,N_2963);
nand UO_363 (O_363,N_2984,N_2974);
nand UO_364 (O_364,N_2987,N_2972);
nand UO_365 (O_365,N_2977,N_2986);
xor UO_366 (O_366,N_2966,N_2983);
nand UO_367 (O_367,N_2973,N_2961);
nand UO_368 (O_368,N_2982,N_2956);
xnor UO_369 (O_369,N_2964,N_2947);
nand UO_370 (O_370,N_2940,N_2943);
and UO_371 (O_371,N_2959,N_2995);
xor UO_372 (O_372,N_2983,N_2988);
and UO_373 (O_373,N_2945,N_2994);
and UO_374 (O_374,N_2982,N_2965);
or UO_375 (O_375,N_2968,N_2963);
and UO_376 (O_376,N_2959,N_2985);
or UO_377 (O_377,N_2974,N_2976);
and UO_378 (O_378,N_2989,N_2964);
and UO_379 (O_379,N_2957,N_2987);
xnor UO_380 (O_380,N_2959,N_2957);
or UO_381 (O_381,N_2974,N_2983);
or UO_382 (O_382,N_2962,N_2988);
xnor UO_383 (O_383,N_2959,N_2983);
xnor UO_384 (O_384,N_2954,N_2967);
xnor UO_385 (O_385,N_2981,N_2944);
nand UO_386 (O_386,N_2965,N_2980);
xor UO_387 (O_387,N_2963,N_2984);
nand UO_388 (O_388,N_2966,N_2960);
nand UO_389 (O_389,N_2965,N_2994);
and UO_390 (O_390,N_2956,N_2950);
xor UO_391 (O_391,N_2986,N_2946);
or UO_392 (O_392,N_2979,N_2971);
or UO_393 (O_393,N_2945,N_2998);
or UO_394 (O_394,N_2984,N_2946);
and UO_395 (O_395,N_2998,N_2952);
nand UO_396 (O_396,N_2991,N_2941);
or UO_397 (O_397,N_2946,N_2957);
nand UO_398 (O_398,N_2975,N_2997);
nand UO_399 (O_399,N_2990,N_2975);
and UO_400 (O_400,N_2962,N_2959);
and UO_401 (O_401,N_2967,N_2950);
nand UO_402 (O_402,N_2980,N_2941);
or UO_403 (O_403,N_2973,N_2987);
xor UO_404 (O_404,N_2979,N_2945);
or UO_405 (O_405,N_2971,N_2958);
and UO_406 (O_406,N_2963,N_2953);
nand UO_407 (O_407,N_2979,N_2992);
or UO_408 (O_408,N_2942,N_2957);
nand UO_409 (O_409,N_2970,N_2966);
or UO_410 (O_410,N_2954,N_2982);
nand UO_411 (O_411,N_2979,N_2989);
or UO_412 (O_412,N_2959,N_2988);
or UO_413 (O_413,N_2978,N_2961);
nor UO_414 (O_414,N_2949,N_2963);
xnor UO_415 (O_415,N_2967,N_2969);
nor UO_416 (O_416,N_2968,N_2955);
xor UO_417 (O_417,N_2965,N_2978);
and UO_418 (O_418,N_2956,N_2953);
xnor UO_419 (O_419,N_2998,N_2984);
xor UO_420 (O_420,N_2980,N_2988);
nand UO_421 (O_421,N_2984,N_2944);
or UO_422 (O_422,N_2987,N_2965);
or UO_423 (O_423,N_2982,N_2942);
xor UO_424 (O_424,N_2989,N_2991);
nand UO_425 (O_425,N_2965,N_2992);
nand UO_426 (O_426,N_2969,N_2980);
or UO_427 (O_427,N_2974,N_2945);
and UO_428 (O_428,N_2971,N_2975);
or UO_429 (O_429,N_2966,N_2946);
nand UO_430 (O_430,N_2995,N_2980);
xnor UO_431 (O_431,N_2955,N_2961);
nand UO_432 (O_432,N_2984,N_2968);
nand UO_433 (O_433,N_2947,N_2969);
and UO_434 (O_434,N_2942,N_2947);
or UO_435 (O_435,N_2988,N_2966);
or UO_436 (O_436,N_2943,N_2962);
or UO_437 (O_437,N_2977,N_2947);
or UO_438 (O_438,N_2956,N_2985);
or UO_439 (O_439,N_2945,N_2968);
xnor UO_440 (O_440,N_2985,N_2948);
or UO_441 (O_441,N_2993,N_2996);
or UO_442 (O_442,N_2969,N_2955);
and UO_443 (O_443,N_2974,N_2982);
xor UO_444 (O_444,N_2949,N_2948);
nand UO_445 (O_445,N_2950,N_2987);
and UO_446 (O_446,N_2988,N_2954);
nor UO_447 (O_447,N_2970,N_2944);
or UO_448 (O_448,N_2985,N_2988);
or UO_449 (O_449,N_2994,N_2952);
and UO_450 (O_450,N_2984,N_2964);
xnor UO_451 (O_451,N_2958,N_2984);
and UO_452 (O_452,N_2959,N_2949);
nor UO_453 (O_453,N_2999,N_2947);
nand UO_454 (O_454,N_2977,N_2978);
and UO_455 (O_455,N_2983,N_2942);
and UO_456 (O_456,N_2973,N_2991);
nor UO_457 (O_457,N_2950,N_2966);
xor UO_458 (O_458,N_2993,N_2972);
nor UO_459 (O_459,N_2968,N_2961);
and UO_460 (O_460,N_2968,N_2974);
and UO_461 (O_461,N_2973,N_2983);
nand UO_462 (O_462,N_2983,N_2949);
and UO_463 (O_463,N_2987,N_2963);
or UO_464 (O_464,N_2961,N_2950);
nor UO_465 (O_465,N_2965,N_2947);
nand UO_466 (O_466,N_2997,N_2948);
xnor UO_467 (O_467,N_2986,N_2955);
xor UO_468 (O_468,N_2981,N_2985);
nor UO_469 (O_469,N_2955,N_2979);
nand UO_470 (O_470,N_2976,N_2947);
and UO_471 (O_471,N_2959,N_2971);
and UO_472 (O_472,N_2983,N_2997);
nor UO_473 (O_473,N_2974,N_2999);
xor UO_474 (O_474,N_2945,N_2966);
or UO_475 (O_475,N_2985,N_2972);
xor UO_476 (O_476,N_2978,N_2986);
nand UO_477 (O_477,N_2946,N_2991);
or UO_478 (O_478,N_2989,N_2983);
and UO_479 (O_479,N_2942,N_2964);
nand UO_480 (O_480,N_2981,N_2971);
nand UO_481 (O_481,N_2940,N_2960);
nor UO_482 (O_482,N_2987,N_2967);
nor UO_483 (O_483,N_2997,N_2977);
xor UO_484 (O_484,N_2996,N_2955);
or UO_485 (O_485,N_2949,N_2996);
xor UO_486 (O_486,N_2998,N_2942);
or UO_487 (O_487,N_2994,N_2942);
or UO_488 (O_488,N_2984,N_2942);
xor UO_489 (O_489,N_2975,N_2946);
and UO_490 (O_490,N_2980,N_2958);
xnor UO_491 (O_491,N_2967,N_2985);
or UO_492 (O_492,N_2990,N_2942);
and UO_493 (O_493,N_2942,N_2970);
nor UO_494 (O_494,N_2983,N_2994);
or UO_495 (O_495,N_2982,N_2979);
and UO_496 (O_496,N_2942,N_2955);
nor UO_497 (O_497,N_2989,N_2955);
or UO_498 (O_498,N_2951,N_2982);
nor UO_499 (O_499,N_2997,N_2947);
endmodule