module basic_750_5000_1000_50_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_633,In_720);
or U1 (N_1,In_351,In_176);
and U2 (N_2,In_583,In_380);
nor U3 (N_3,In_449,In_644);
and U4 (N_4,In_672,In_111);
or U5 (N_5,In_262,In_737);
or U6 (N_6,In_463,In_649);
nor U7 (N_7,In_427,In_187);
and U8 (N_8,In_130,In_31);
nor U9 (N_9,In_25,In_586);
nor U10 (N_10,In_406,In_582);
or U11 (N_11,In_159,In_437);
xor U12 (N_12,In_614,In_482);
or U13 (N_13,In_599,In_597);
xnor U14 (N_14,In_496,In_106);
nand U15 (N_15,In_151,In_578);
nor U16 (N_16,In_363,In_180);
and U17 (N_17,In_626,In_569);
and U18 (N_18,In_472,In_272);
nand U19 (N_19,In_192,In_728);
nand U20 (N_20,In_28,In_348);
nor U21 (N_21,In_331,In_654);
nand U22 (N_22,In_598,In_345);
nor U23 (N_23,In_89,In_369);
or U24 (N_24,In_319,In_148);
and U25 (N_25,In_109,In_228);
or U26 (N_26,In_710,In_600);
and U27 (N_27,In_123,In_204);
and U28 (N_28,In_212,In_142);
nor U29 (N_29,In_201,In_709);
or U30 (N_30,In_0,In_383);
and U31 (N_31,In_155,In_152);
and U32 (N_32,In_459,In_513);
nand U33 (N_33,In_703,In_305);
nor U34 (N_34,In_622,In_743);
nand U35 (N_35,In_617,In_244);
or U36 (N_36,In_211,In_362);
xnor U37 (N_37,In_516,In_475);
nand U38 (N_38,In_556,In_81);
nand U39 (N_39,In_120,In_446);
and U40 (N_40,In_367,In_13);
nand U41 (N_41,In_515,In_317);
or U42 (N_42,In_718,In_87);
and U43 (N_43,In_386,In_181);
nand U44 (N_44,In_267,In_371);
nand U45 (N_45,In_542,In_687);
nand U46 (N_46,In_342,In_392);
nand U47 (N_47,In_609,In_659);
or U48 (N_48,In_602,In_154);
or U49 (N_49,In_717,In_424);
nor U50 (N_50,In_539,In_567);
nand U51 (N_51,In_107,In_389);
xnor U52 (N_52,In_396,In_403);
xor U53 (N_53,In_686,In_511);
nor U54 (N_54,In_671,In_388);
or U55 (N_55,In_603,In_354);
or U56 (N_56,In_101,In_283);
nand U57 (N_57,In_105,In_382);
nor U58 (N_58,In_534,In_564);
or U59 (N_59,In_69,In_713);
or U60 (N_60,In_210,In_410);
nor U61 (N_61,In_52,In_575);
or U62 (N_62,In_476,In_714);
and U63 (N_63,In_337,In_208);
xnor U64 (N_64,In_218,In_316);
and U65 (N_65,In_263,In_335);
and U66 (N_66,In_332,In_420);
xnor U67 (N_67,In_546,In_184);
and U68 (N_68,In_118,In_224);
nand U69 (N_69,In_127,In_502);
or U70 (N_70,In_697,In_333);
nand U71 (N_71,In_77,In_115);
nand U72 (N_72,In_174,In_349);
nor U73 (N_73,In_40,In_723);
or U74 (N_74,In_615,In_78);
nor U75 (N_75,In_565,In_97);
or U76 (N_76,In_494,In_477);
nor U77 (N_77,In_233,In_311);
xor U78 (N_78,In_601,In_65);
and U79 (N_79,In_230,In_408);
nand U80 (N_80,In_533,In_458);
nor U81 (N_81,In_580,In_480);
xor U82 (N_82,In_676,In_685);
and U83 (N_83,In_699,In_253);
xnor U84 (N_84,In_315,In_327);
or U85 (N_85,In_499,In_295);
nand U86 (N_86,In_229,In_72);
and U87 (N_87,In_219,In_287);
nor U88 (N_88,In_606,In_145);
and U89 (N_89,In_167,In_632);
or U90 (N_90,In_468,In_535);
nand U91 (N_91,In_103,In_241);
nor U92 (N_92,In_140,In_59);
nor U93 (N_93,In_278,In_226);
and U94 (N_94,In_456,In_221);
nor U95 (N_95,In_455,In_510);
and U96 (N_96,In_498,In_225);
or U97 (N_97,In_265,In_397);
nor U98 (N_98,In_18,In_621);
nand U99 (N_99,In_435,In_312);
or U100 (N_100,In_175,In_726);
xor U101 (N_101,N_49,In_135);
or U102 (N_102,N_31,In_343);
or U103 (N_103,In_310,In_273);
nor U104 (N_104,In_462,In_339);
and U105 (N_105,In_85,In_189);
nand U106 (N_106,In_661,In_722);
nor U107 (N_107,In_506,In_402);
or U108 (N_108,N_8,N_24);
xnor U109 (N_109,In_745,In_683);
nand U110 (N_110,In_270,In_238);
nand U111 (N_111,N_26,In_326);
nand U112 (N_112,In_252,In_490);
nor U113 (N_113,In_747,In_652);
xor U114 (N_114,In_55,N_18);
nor U115 (N_115,In_23,In_520);
or U116 (N_116,In_119,In_635);
nand U117 (N_117,In_356,In_27);
nor U118 (N_118,In_376,In_607);
or U119 (N_119,In_156,In_716);
xor U120 (N_120,N_63,In_725);
and U121 (N_121,N_2,In_215);
nand U122 (N_122,In_46,In_261);
nand U123 (N_123,In_596,In_438);
nor U124 (N_124,In_730,N_4);
nor U125 (N_125,In_604,In_338);
nor U126 (N_126,In_347,In_536);
and U127 (N_127,In_129,In_553);
and U128 (N_128,In_418,In_688);
nor U129 (N_129,N_73,In_409);
nand U130 (N_130,In_405,In_99);
nor U131 (N_131,In_60,In_74);
nand U132 (N_132,In_577,In_594);
nor U133 (N_133,In_613,In_377);
and U134 (N_134,In_680,In_417);
nor U135 (N_135,In_630,N_16);
or U136 (N_136,In_138,In_150);
nor U137 (N_137,In_341,In_558);
xnor U138 (N_138,In_746,In_724);
or U139 (N_139,N_32,In_268);
or U140 (N_140,In_442,In_441);
and U141 (N_141,N_3,In_595);
nand U142 (N_142,In_641,In_731);
nor U143 (N_143,In_705,In_6);
and U144 (N_144,In_443,In_572);
nand U145 (N_145,In_374,In_400);
or U146 (N_146,N_91,In_675);
and U147 (N_147,In_308,In_281);
nand U148 (N_148,N_19,In_368);
nand U149 (N_149,In_271,In_209);
or U150 (N_150,N_79,In_289);
and U151 (N_151,In_484,N_20);
nand U152 (N_152,In_514,In_309);
or U153 (N_153,In_610,In_372);
nand U154 (N_154,In_668,In_82);
xor U155 (N_155,In_29,In_474);
nand U156 (N_156,In_67,N_13);
nor U157 (N_157,N_28,In_413);
and U158 (N_158,In_693,In_620);
nand U159 (N_159,In_530,In_227);
and U160 (N_160,N_87,N_6);
nand U161 (N_161,In_447,In_203);
or U162 (N_162,In_508,In_44);
nor U163 (N_163,In_398,In_117);
nand U164 (N_164,In_94,In_220);
nand U165 (N_165,In_414,N_83);
nand U166 (N_166,In_179,In_76);
or U167 (N_167,In_346,In_658);
nand U168 (N_168,In_395,In_86);
and U169 (N_169,In_170,In_231);
nor U170 (N_170,N_7,In_681);
nand U171 (N_171,In_216,In_526);
nor U172 (N_172,In_290,In_197);
and U173 (N_173,In_532,In_370);
or U174 (N_174,In_200,In_584);
nor U175 (N_175,In_576,In_605);
or U176 (N_176,In_637,In_670);
xor U177 (N_177,N_56,In_242);
nand U178 (N_178,In_519,In_75);
nand U179 (N_179,In_297,In_149);
and U180 (N_180,In_591,In_694);
and U181 (N_181,In_571,In_436);
nor U182 (N_182,In_139,In_550);
or U183 (N_183,In_450,In_399);
or U184 (N_184,In_39,In_375);
nor U185 (N_185,In_232,In_1);
and U186 (N_186,N_78,In_300);
and U187 (N_187,N_84,In_104);
or U188 (N_188,N_64,In_143);
or U189 (N_189,In_291,In_512);
and U190 (N_190,N_11,In_147);
xor U191 (N_191,N_40,In_34);
nand U192 (N_192,In_581,In_660);
xnor U193 (N_193,In_173,In_298);
nor U194 (N_194,In_266,In_222);
nor U195 (N_195,In_320,In_7);
and U196 (N_196,In_733,In_568);
and U197 (N_197,In_715,In_691);
nand U198 (N_198,In_529,In_381);
nand U199 (N_199,In_285,In_545);
and U200 (N_200,In_49,In_68);
or U201 (N_201,N_146,In_689);
and U202 (N_202,In_740,In_698);
and U203 (N_203,In_169,N_191);
nand U204 (N_204,N_170,N_45);
or U205 (N_205,In_634,In_695);
or U206 (N_206,N_173,N_159);
xnor U207 (N_207,N_152,N_5);
or U208 (N_208,In_523,N_154);
nor U209 (N_209,In_561,In_525);
xor U210 (N_210,In_656,In_58);
nor U211 (N_211,N_96,N_76);
xnor U212 (N_212,N_115,In_531);
and U213 (N_213,N_179,In_144);
nor U214 (N_214,In_61,In_554);
nand U215 (N_215,In_639,In_128);
nand U216 (N_216,N_143,In_264);
nor U217 (N_217,In_647,In_505);
or U218 (N_218,N_109,In_547);
nand U219 (N_219,N_134,In_276);
or U220 (N_220,In_719,In_419);
or U221 (N_221,In_440,In_422);
nand U222 (N_222,In_153,N_141);
nor U223 (N_223,In_146,In_416);
nand U224 (N_224,In_157,In_122);
and U225 (N_225,In_282,N_55);
nor U226 (N_226,N_137,In_359);
and U227 (N_227,In_178,N_22);
nand U228 (N_228,In_537,N_132);
nor U229 (N_229,In_251,In_579);
nor U230 (N_230,In_318,N_25);
or U231 (N_231,In_432,In_528);
and U232 (N_232,In_84,In_629);
xor U233 (N_233,In_702,In_552);
xor U234 (N_234,In_36,In_744);
or U235 (N_235,In_454,N_94);
nand U236 (N_236,In_729,N_195);
nand U237 (N_237,In_663,In_678);
xnor U238 (N_238,In_682,N_147);
nand U239 (N_239,In_205,In_83);
and U240 (N_240,In_95,In_88);
nand U241 (N_241,In_33,In_194);
nor U242 (N_242,In_121,N_44);
nor U243 (N_243,N_165,In_471);
nand U244 (N_244,In_302,In_162);
xor U245 (N_245,N_99,N_95);
or U246 (N_246,N_161,In_551);
nand U247 (N_247,In_373,In_428);
nand U248 (N_248,N_62,N_53);
xor U249 (N_249,In_674,In_464);
nand U250 (N_250,In_650,N_140);
and U251 (N_251,In_645,In_361);
or U252 (N_252,In_217,In_141);
or U253 (N_253,In_466,In_71);
or U254 (N_254,In_288,N_21);
and U255 (N_255,N_133,In_679);
xor U256 (N_256,In_448,In_469);
or U257 (N_257,In_182,In_379);
nand U258 (N_258,In_589,In_735);
nand U259 (N_259,In_636,In_473);
nor U260 (N_260,N_93,In_704);
nand U261 (N_261,In_50,In_616);
or U262 (N_262,N_122,N_85);
xnor U263 (N_263,In_538,N_184);
and U264 (N_264,In_240,N_144);
and U265 (N_265,In_711,In_131);
xor U266 (N_266,N_51,N_97);
nand U267 (N_267,N_166,N_172);
and U268 (N_268,In_648,In_223);
or U269 (N_269,In_191,N_42);
or U270 (N_270,In_465,In_543);
and U271 (N_271,In_415,In_236);
nand U272 (N_272,In_116,N_75);
nor U273 (N_273,In_387,In_665);
xor U274 (N_274,In_549,N_194);
nand U275 (N_275,In_133,N_9);
and U276 (N_276,In_412,In_451);
nor U277 (N_277,In_5,In_485);
nand U278 (N_278,In_559,N_118);
nand U279 (N_279,In_366,In_736);
nand U280 (N_280,In_12,N_102);
nand U281 (N_281,In_334,In_38);
and U282 (N_282,N_125,In_113);
nor U283 (N_283,In_165,In_394);
nand U284 (N_284,N_60,In_353);
and U285 (N_285,In_669,N_46);
xnor U286 (N_286,In_108,N_66);
or U287 (N_287,In_560,In_196);
or U288 (N_288,In_453,N_104);
or U289 (N_289,In_80,In_56);
or U290 (N_290,In_277,N_103);
nor U291 (N_291,N_164,N_54);
nor U292 (N_292,In_344,In_235);
nand U293 (N_293,N_61,In_37);
nand U294 (N_294,In_62,N_10);
nor U295 (N_295,In_623,In_4);
or U296 (N_296,N_182,N_82);
xnor U297 (N_297,In_246,In_279);
nand U298 (N_298,N_70,In_357);
and U299 (N_299,In_306,In_585);
and U300 (N_300,In_137,N_177);
or U301 (N_301,In_612,In_213);
nand U302 (N_302,N_47,In_425);
and U303 (N_303,N_175,N_289);
and U304 (N_304,In_488,N_174);
nor U305 (N_305,N_252,In_202);
xor U306 (N_306,N_167,N_180);
and U307 (N_307,N_72,In_314);
nor U308 (N_308,In_17,N_43);
xnor U309 (N_309,In_41,N_185);
xor U310 (N_310,In_664,In_254);
nand U311 (N_311,In_673,In_110);
or U312 (N_312,N_124,N_261);
nand U313 (N_313,In_43,In_470);
and U314 (N_314,In_256,In_26);
or U315 (N_315,In_54,In_350);
and U316 (N_316,In_696,In_98);
xor U317 (N_317,N_230,In_352);
nor U318 (N_318,N_92,In_323);
nand U319 (N_319,In_324,N_292);
or U320 (N_320,N_258,In_421);
and U321 (N_321,In_21,In_284);
nor U322 (N_322,N_59,In_708);
nor U323 (N_323,In_24,In_8);
nand U324 (N_324,In_748,In_20);
or U325 (N_325,N_206,N_98);
nor U326 (N_326,In_631,In_573);
or U327 (N_327,N_1,In_646);
nand U328 (N_328,N_114,In_30);
nor U329 (N_329,N_218,N_226);
nor U330 (N_330,N_37,N_169);
nand U331 (N_331,N_110,N_284);
nand U332 (N_332,In_677,N_150);
nor U333 (N_333,In_299,In_732);
or U334 (N_334,In_293,N_278);
and U335 (N_335,In_330,N_36);
nor U336 (N_336,In_364,N_120);
nor U337 (N_337,N_39,In_439);
and U338 (N_338,N_293,N_71);
nor U339 (N_339,N_101,N_211);
nor U340 (N_340,N_156,In_183);
nand U341 (N_341,In_325,In_63);
and U342 (N_342,In_426,N_223);
nor U343 (N_343,N_129,In_79);
nand U344 (N_344,N_222,N_162);
and U345 (N_345,In_642,In_358);
nor U346 (N_346,In_625,In_294);
and U347 (N_347,In_42,N_214);
and U348 (N_348,In_391,In_507);
and U349 (N_349,N_272,In_501);
nand U350 (N_350,In_574,N_247);
nand U351 (N_351,N_112,N_149);
or U352 (N_352,In_478,In_237);
and U353 (N_353,In_11,In_22);
nor U354 (N_354,In_292,In_190);
or U355 (N_355,In_247,In_739);
and U356 (N_356,N_113,In_35);
and U357 (N_357,N_227,In_521);
nor U358 (N_358,N_263,N_192);
nand U359 (N_359,In_692,N_245);
and U360 (N_360,N_229,In_667);
nand U361 (N_361,In_548,In_164);
and U362 (N_362,N_208,N_186);
nand U363 (N_363,In_322,N_216);
nand U364 (N_364,In_53,In_45);
nor U365 (N_365,In_274,In_245);
and U366 (N_366,In_163,In_177);
nand U367 (N_367,N_281,In_125);
or U368 (N_368,In_541,N_57);
nor U369 (N_369,In_2,In_503);
nand U370 (N_370,N_267,In_51);
nor U371 (N_371,In_185,In_378);
or U372 (N_372,In_234,In_214);
nor U373 (N_373,In_114,In_522);
nand U374 (N_374,In_701,N_205);
and U375 (N_375,In_64,N_196);
and U376 (N_376,N_273,N_197);
xnor U377 (N_377,N_232,In_102);
xor U378 (N_378,In_401,In_186);
and U379 (N_379,N_240,N_243);
xor U380 (N_380,In_168,In_92);
nor U381 (N_381,N_121,In_497);
or U382 (N_382,N_100,In_258);
and U383 (N_383,N_259,N_210);
and U384 (N_384,In_742,N_219);
or U385 (N_385,In_269,N_241);
nand U386 (N_386,N_264,N_52);
or U387 (N_387,N_119,N_295);
nand U388 (N_388,In_707,N_260);
nor U389 (N_389,In_198,In_562);
nor U390 (N_390,In_304,In_566);
or U391 (N_391,In_248,In_411);
or U392 (N_392,In_429,In_624);
and U393 (N_393,In_239,In_452);
and U394 (N_394,N_203,N_190);
and U395 (N_395,In_206,In_445);
nor U396 (N_396,N_127,N_131);
and U397 (N_397,In_741,N_33);
or U398 (N_398,N_198,In_544);
nor U399 (N_399,N_280,N_276);
nor U400 (N_400,N_354,N_130);
nand U401 (N_401,N_189,N_328);
and U402 (N_402,In_321,In_275);
or U403 (N_403,N_376,N_246);
xor U404 (N_404,In_619,In_608);
xnor U405 (N_405,N_116,N_212);
nor U406 (N_406,N_30,N_357);
or U407 (N_407,In_91,N_355);
nor U408 (N_408,In_15,N_88);
nor U409 (N_409,N_283,N_251);
nor U410 (N_410,N_364,N_142);
and U411 (N_411,In_518,N_326);
and U412 (N_412,In_188,N_145);
or U413 (N_413,N_366,In_495);
and U414 (N_414,N_309,N_389);
and U415 (N_415,N_23,In_486);
or U416 (N_416,In_627,N_231);
nor U417 (N_417,In_457,In_690);
and U418 (N_418,N_234,N_153);
xor U419 (N_419,In_307,N_373);
or U420 (N_420,N_136,In_136);
or U421 (N_421,In_250,N_123);
and U422 (N_422,N_349,N_378);
nand U423 (N_423,N_81,N_271);
and U424 (N_424,N_343,N_307);
nor U425 (N_425,N_244,N_80);
xnor U426 (N_426,N_320,In_260);
or U427 (N_427,N_238,N_316);
or U428 (N_428,In_161,N_67);
or U429 (N_429,In_100,N_265);
nand U430 (N_430,In_160,N_270);
nand U431 (N_431,N_90,In_3);
or U432 (N_432,N_331,N_237);
nor U433 (N_433,In_492,N_380);
nor U434 (N_434,In_509,N_358);
and U435 (N_435,N_399,In_195);
nor U436 (N_436,N_250,N_294);
nor U437 (N_437,N_207,In_280);
and U438 (N_438,N_287,N_356);
or U439 (N_439,N_363,In_489);
nor U440 (N_440,N_105,N_353);
nand U441 (N_441,N_350,In_517);
or U442 (N_442,N_369,In_727);
nand U443 (N_443,N_257,N_288);
and U444 (N_444,In_32,N_346);
or U445 (N_445,In_721,N_297);
nor U446 (N_446,N_303,N_318);
or U447 (N_447,N_248,N_74);
and U448 (N_448,In_700,In_14);
nor U449 (N_449,In_444,In_112);
nand U450 (N_450,N_298,N_155);
xor U451 (N_451,N_168,N_262);
and U452 (N_452,N_351,N_334);
nor U453 (N_453,N_342,In_592);
nor U454 (N_454,In_433,N_176);
xor U455 (N_455,N_388,N_128);
and U456 (N_456,N_213,N_340);
nor U457 (N_457,N_86,N_29);
or U458 (N_458,N_200,In_73);
nand U459 (N_459,N_126,N_317);
and U460 (N_460,N_217,N_117);
and U461 (N_461,N_359,N_148);
and U462 (N_462,N_345,N_305);
nand U463 (N_463,N_225,N_171);
nor U464 (N_464,N_239,N_193);
xor U465 (N_465,N_348,N_183);
nor U466 (N_466,N_301,N_188);
and U467 (N_467,N_352,N_325);
nand U468 (N_468,N_135,N_277);
or U469 (N_469,In_491,N_220);
nor U470 (N_470,N_201,N_181);
or U471 (N_471,In_93,N_361);
nand U472 (N_472,N_337,In_9);
nand U473 (N_473,N_204,In_481);
nand U474 (N_474,In_618,N_89);
and U475 (N_475,N_151,N_370);
nor U476 (N_476,In_66,In_407);
nand U477 (N_477,N_310,N_14);
nor U478 (N_478,In_540,In_611);
nor U479 (N_479,In_355,N_323);
and U480 (N_480,N_315,N_377);
or U481 (N_481,N_269,In_19);
or U482 (N_482,N_34,In_493);
nor U483 (N_483,In_749,N_398);
nand U484 (N_484,N_286,In_557);
or U485 (N_485,In_132,N_255);
nand U486 (N_486,In_257,In_460);
nand U487 (N_487,N_319,N_268);
and U488 (N_488,In_259,In_527);
and U489 (N_489,N_139,In_738);
nor U490 (N_490,N_215,In_487);
nor U491 (N_491,N_108,In_657);
nand U492 (N_492,N_209,In_158);
and U493 (N_493,N_344,In_385);
nand U494 (N_494,N_372,N_158);
nor U495 (N_495,N_336,N_157);
nor U496 (N_496,In_563,N_324);
and U497 (N_497,N_68,N_392);
and U498 (N_498,N_65,N_12);
nand U499 (N_499,In_134,In_479);
and U500 (N_500,N_432,N_418);
or U501 (N_501,N_467,N_457);
nand U502 (N_502,In_199,N_312);
and U503 (N_503,In_588,N_473);
nor U504 (N_504,In_16,N_327);
nor U505 (N_505,N_329,N_444);
or U506 (N_506,In_431,N_406);
nor U507 (N_507,N_368,N_417);
xor U508 (N_508,N_497,N_313);
or U509 (N_509,N_486,N_470);
or U510 (N_510,N_415,N_448);
nand U511 (N_511,In_328,In_336);
or U512 (N_512,N_106,N_381);
xnor U513 (N_513,N_423,N_479);
and U514 (N_514,N_362,N_256);
nor U515 (N_515,N_498,N_178);
or U516 (N_516,N_439,N_441);
or U517 (N_517,In_638,N_442);
nor U518 (N_518,N_274,N_476);
and U519 (N_519,N_333,N_367);
nor U520 (N_520,N_412,N_474);
nand U521 (N_521,N_224,N_38);
nand U522 (N_522,In_193,N_405);
nor U523 (N_523,In_593,N_304);
nand U524 (N_524,N_456,N_426);
nor U525 (N_525,In_734,In_171);
nor U526 (N_526,N_409,N_458);
nand U527 (N_527,In_587,In_666);
xnor U528 (N_528,N_379,In_47);
nor U529 (N_529,In_365,N_496);
nor U530 (N_530,N_382,N_430);
xnor U531 (N_531,N_464,N_77);
nor U532 (N_532,N_386,In_313);
and U533 (N_533,N_452,N_433);
nand U534 (N_534,In_655,N_481);
or U535 (N_535,N_17,N_468);
or U536 (N_536,N_111,N_35);
nor U537 (N_537,In_48,In_483);
nand U538 (N_538,N_254,N_275);
and U539 (N_539,In_70,In_90);
or U540 (N_540,N_332,N_487);
or U541 (N_541,N_495,N_494);
and U542 (N_542,N_438,N_347);
nor U543 (N_543,N_484,N_299);
and U544 (N_544,N_461,N_385);
or U545 (N_545,N_365,N_374);
or U546 (N_546,N_27,N_431);
nand U547 (N_547,N_330,N_472);
or U548 (N_548,N_463,N_475);
or U549 (N_549,N_401,N_58);
nor U550 (N_550,N_493,In_255);
or U551 (N_551,N_390,In_570);
and U552 (N_552,N_440,N_422);
nand U553 (N_553,N_459,N_436);
and U554 (N_554,In_662,N_454);
nand U555 (N_555,N_480,In_126);
nor U556 (N_556,N_477,In_286);
and U557 (N_557,N_163,N_428);
xor U558 (N_558,In_243,In_712);
and U559 (N_559,N_446,N_478);
or U560 (N_560,N_314,In_390);
and U561 (N_561,N_249,In_57);
or U562 (N_562,N_420,N_0);
or U563 (N_563,In_467,In_524);
nand U564 (N_564,N_300,N_202);
or U565 (N_565,N_445,N_306);
nand U566 (N_566,N_235,In_96);
and U567 (N_567,N_492,In_303);
xor U568 (N_568,N_279,In_10);
xor U569 (N_569,N_413,N_50);
or U570 (N_570,In_393,N_434);
nand U571 (N_571,In_706,N_471);
nand U572 (N_572,In_166,N_308);
or U573 (N_573,N_338,N_419);
and U574 (N_574,In_340,N_400);
and U575 (N_575,In_384,N_296);
or U576 (N_576,In_301,N_414);
and U577 (N_577,In_500,N_488);
and U578 (N_578,N_437,In_423);
nor U579 (N_579,N_499,N_285);
and U580 (N_580,N_408,N_321);
nor U581 (N_581,N_396,N_48);
and U582 (N_582,N_375,N_485);
or U583 (N_583,N_397,N_233);
or U584 (N_584,N_384,In_172);
nor U585 (N_585,N_435,N_483);
xnor U586 (N_586,N_466,N_469);
nand U587 (N_587,N_425,In_124);
nand U588 (N_588,N_290,N_395);
or U589 (N_589,In_434,N_443);
and U590 (N_590,N_427,N_460);
or U591 (N_591,In_651,N_302);
and U592 (N_592,N_455,N_429);
and U593 (N_593,N_138,N_311);
xor U594 (N_594,N_424,In_461);
and U595 (N_595,In_329,N_187);
nor U596 (N_596,N_482,N_387);
nand U597 (N_597,N_160,N_15);
and U598 (N_598,N_393,N_291);
and U599 (N_599,N_462,N_402);
nor U600 (N_600,N_339,N_519);
nand U601 (N_601,N_500,N_562);
nor U602 (N_602,N_391,N_543);
and U603 (N_603,In_643,N_199);
or U604 (N_604,N_553,N_410);
nor U605 (N_605,N_555,N_489);
and U606 (N_606,N_564,N_221);
nor U607 (N_607,N_574,N_563);
xor U608 (N_608,N_594,N_537);
xor U609 (N_609,In_504,N_575);
nor U610 (N_610,N_546,N_536);
nand U611 (N_611,N_411,N_341);
nor U612 (N_612,N_566,In_590);
and U613 (N_613,In_628,N_534);
and U614 (N_614,N_236,N_41);
nand U615 (N_615,In_555,N_588);
or U616 (N_616,N_421,N_590);
or U617 (N_617,N_451,N_540);
and U618 (N_618,N_512,N_514);
or U619 (N_619,N_541,N_450);
or U620 (N_620,N_583,N_554);
xnor U621 (N_621,N_580,N_525);
or U622 (N_622,N_503,N_577);
nand U623 (N_623,In_640,N_506);
nand U624 (N_624,N_599,N_228);
or U625 (N_625,N_491,N_570);
and U626 (N_626,N_490,N_515);
nor U627 (N_627,N_582,N_383);
and U628 (N_628,N_559,N_394);
nand U629 (N_629,N_360,N_522);
nand U630 (N_630,N_516,N_547);
nand U631 (N_631,N_579,In_207);
and U632 (N_632,N_510,N_545);
nor U633 (N_633,N_548,N_586);
or U634 (N_634,N_416,N_505);
or U635 (N_635,N_107,N_521);
or U636 (N_636,N_576,N_465);
or U637 (N_637,N_517,N_592);
or U638 (N_638,N_544,In_296);
or U639 (N_639,N_556,N_509);
nand U640 (N_640,N_266,N_453);
nor U641 (N_641,N_529,N_571);
nor U642 (N_642,N_561,In_249);
and U643 (N_643,N_523,N_242);
nand U644 (N_644,N_532,In_360);
and U645 (N_645,N_404,N_584);
xor U646 (N_646,N_585,N_502);
nand U647 (N_647,N_403,N_371);
nand U648 (N_648,N_542,N_597);
or U649 (N_649,In_404,N_504);
nand U650 (N_650,N_572,N_518);
nand U651 (N_651,N_593,N_551);
and U652 (N_652,N_568,N_560);
nor U653 (N_653,N_507,N_596);
nand U654 (N_654,In_430,N_520);
or U655 (N_655,N_449,N_526);
nand U656 (N_656,N_447,N_513);
xor U657 (N_657,N_531,N_282);
or U658 (N_658,N_527,N_595);
and U659 (N_659,N_569,N_550);
nor U660 (N_660,N_558,N_322);
and U661 (N_661,N_557,N_581);
or U662 (N_662,N_508,N_535);
nor U663 (N_663,N_549,N_567);
nand U664 (N_664,N_598,N_589);
nor U665 (N_665,N_539,N_407);
and U666 (N_666,N_591,N_552);
and U667 (N_667,N_530,N_253);
nor U668 (N_668,In_653,N_335);
nor U669 (N_669,N_511,N_538);
nand U670 (N_670,N_528,N_578);
and U671 (N_671,N_573,N_524);
nand U672 (N_672,In_684,N_69);
and U673 (N_673,N_501,N_587);
or U674 (N_674,N_565,N_533);
nor U675 (N_675,N_576,N_559);
xor U676 (N_676,N_545,N_515);
and U677 (N_677,N_504,N_552);
nand U678 (N_678,N_571,N_549);
nor U679 (N_679,N_590,N_507);
nor U680 (N_680,N_571,N_520);
nand U681 (N_681,N_407,N_556);
xor U682 (N_682,N_558,N_561);
or U683 (N_683,N_228,N_221);
and U684 (N_684,In_249,In_430);
or U685 (N_685,N_539,N_597);
and U686 (N_686,N_530,N_571);
or U687 (N_687,N_599,N_522);
nor U688 (N_688,N_341,N_544);
nand U689 (N_689,N_341,N_266);
nand U690 (N_690,N_531,N_595);
nand U691 (N_691,N_228,N_416);
nor U692 (N_692,N_371,In_404);
and U693 (N_693,N_199,N_548);
and U694 (N_694,N_595,N_549);
nand U695 (N_695,N_517,N_576);
or U696 (N_696,N_236,N_543);
and U697 (N_697,N_555,N_536);
nand U698 (N_698,N_586,N_532);
nor U699 (N_699,N_543,N_571);
nand U700 (N_700,N_675,N_611);
or U701 (N_701,N_676,N_682);
nor U702 (N_702,N_698,N_681);
nor U703 (N_703,N_692,N_651);
or U704 (N_704,N_694,N_663);
or U705 (N_705,N_680,N_635);
nand U706 (N_706,N_613,N_622);
or U707 (N_707,N_607,N_670);
and U708 (N_708,N_603,N_661);
nor U709 (N_709,N_628,N_688);
nand U710 (N_710,N_686,N_650);
or U711 (N_711,N_699,N_695);
and U712 (N_712,N_644,N_642);
or U713 (N_713,N_636,N_679);
and U714 (N_714,N_623,N_677);
and U715 (N_715,N_606,N_659);
xor U716 (N_716,N_652,N_647);
xor U717 (N_717,N_619,N_673);
or U718 (N_718,N_641,N_634);
nor U719 (N_719,N_610,N_625);
nand U720 (N_720,N_639,N_687);
and U721 (N_721,N_665,N_648);
nor U722 (N_722,N_616,N_666);
or U723 (N_723,N_660,N_685);
and U724 (N_724,N_646,N_600);
or U725 (N_725,N_671,N_618);
or U726 (N_726,N_620,N_684);
and U727 (N_727,N_658,N_662);
nand U728 (N_728,N_653,N_689);
nand U729 (N_729,N_637,N_668);
nand U730 (N_730,N_696,N_664);
nand U731 (N_731,N_657,N_631);
nor U732 (N_732,N_632,N_605);
or U733 (N_733,N_656,N_649);
nor U734 (N_734,N_629,N_627);
and U735 (N_735,N_697,N_633);
nor U736 (N_736,N_617,N_638);
and U737 (N_737,N_640,N_604);
and U738 (N_738,N_678,N_691);
nand U739 (N_739,N_690,N_602);
and U740 (N_740,N_615,N_630);
or U741 (N_741,N_612,N_609);
nand U742 (N_742,N_683,N_626);
and U743 (N_743,N_672,N_674);
nor U744 (N_744,N_645,N_643);
and U745 (N_745,N_654,N_614);
or U746 (N_746,N_621,N_655);
or U747 (N_747,N_693,N_667);
or U748 (N_748,N_669,N_608);
or U749 (N_749,N_624,N_601);
and U750 (N_750,N_657,N_671);
and U751 (N_751,N_668,N_676);
and U752 (N_752,N_644,N_693);
nand U753 (N_753,N_666,N_693);
nor U754 (N_754,N_696,N_609);
xnor U755 (N_755,N_617,N_618);
nand U756 (N_756,N_661,N_695);
xnor U757 (N_757,N_670,N_651);
or U758 (N_758,N_688,N_602);
nor U759 (N_759,N_668,N_677);
or U760 (N_760,N_602,N_614);
nand U761 (N_761,N_685,N_619);
nor U762 (N_762,N_604,N_644);
nand U763 (N_763,N_628,N_636);
xor U764 (N_764,N_639,N_682);
and U765 (N_765,N_612,N_608);
or U766 (N_766,N_694,N_661);
nor U767 (N_767,N_659,N_609);
and U768 (N_768,N_663,N_672);
or U769 (N_769,N_653,N_648);
nand U770 (N_770,N_673,N_677);
nand U771 (N_771,N_639,N_667);
nor U772 (N_772,N_619,N_664);
xor U773 (N_773,N_612,N_634);
xnor U774 (N_774,N_661,N_666);
and U775 (N_775,N_698,N_633);
xor U776 (N_776,N_623,N_683);
nor U777 (N_777,N_658,N_623);
nand U778 (N_778,N_674,N_673);
and U779 (N_779,N_671,N_629);
nor U780 (N_780,N_678,N_616);
or U781 (N_781,N_605,N_614);
xnor U782 (N_782,N_672,N_645);
or U783 (N_783,N_604,N_662);
nand U784 (N_784,N_686,N_687);
nand U785 (N_785,N_652,N_683);
or U786 (N_786,N_663,N_668);
nor U787 (N_787,N_663,N_632);
nor U788 (N_788,N_656,N_658);
or U789 (N_789,N_670,N_660);
and U790 (N_790,N_631,N_667);
and U791 (N_791,N_634,N_657);
nand U792 (N_792,N_664,N_672);
and U793 (N_793,N_662,N_679);
nand U794 (N_794,N_695,N_633);
and U795 (N_795,N_638,N_685);
or U796 (N_796,N_659,N_621);
nor U797 (N_797,N_668,N_651);
nand U798 (N_798,N_615,N_620);
and U799 (N_799,N_667,N_679);
and U800 (N_800,N_766,N_784);
nor U801 (N_801,N_758,N_710);
and U802 (N_802,N_755,N_760);
or U803 (N_803,N_721,N_748);
nand U804 (N_804,N_799,N_743);
nor U805 (N_805,N_734,N_708);
nor U806 (N_806,N_788,N_779);
and U807 (N_807,N_752,N_744);
or U808 (N_808,N_717,N_780);
or U809 (N_809,N_777,N_764);
or U810 (N_810,N_761,N_737);
nor U811 (N_811,N_733,N_776);
and U812 (N_812,N_749,N_709);
nor U813 (N_813,N_742,N_705);
nand U814 (N_814,N_785,N_723);
nor U815 (N_815,N_778,N_753);
or U816 (N_816,N_715,N_794);
and U817 (N_817,N_740,N_798);
and U818 (N_818,N_750,N_772);
or U819 (N_819,N_728,N_716);
nand U820 (N_820,N_738,N_725);
or U821 (N_821,N_797,N_735);
xnor U822 (N_822,N_703,N_775);
nand U823 (N_823,N_736,N_754);
and U824 (N_824,N_759,N_747);
nor U825 (N_825,N_792,N_793);
and U826 (N_826,N_768,N_751);
and U827 (N_827,N_790,N_701);
nand U828 (N_828,N_730,N_781);
nand U829 (N_829,N_763,N_746);
and U830 (N_830,N_718,N_713);
or U831 (N_831,N_770,N_739);
and U832 (N_832,N_722,N_773);
and U833 (N_833,N_714,N_783);
xnor U834 (N_834,N_767,N_757);
nand U835 (N_835,N_732,N_706);
and U836 (N_836,N_731,N_787);
nor U837 (N_837,N_712,N_726);
or U838 (N_838,N_762,N_707);
or U839 (N_839,N_720,N_700);
nand U840 (N_840,N_791,N_786);
nor U841 (N_841,N_727,N_729);
nor U842 (N_842,N_719,N_796);
or U843 (N_843,N_771,N_769);
nor U844 (N_844,N_724,N_765);
nor U845 (N_845,N_741,N_782);
and U846 (N_846,N_711,N_702);
xnor U847 (N_847,N_789,N_704);
nand U848 (N_848,N_774,N_745);
and U849 (N_849,N_756,N_795);
nor U850 (N_850,N_721,N_747);
or U851 (N_851,N_757,N_703);
nand U852 (N_852,N_740,N_796);
and U853 (N_853,N_790,N_756);
nand U854 (N_854,N_701,N_783);
or U855 (N_855,N_789,N_715);
nor U856 (N_856,N_743,N_725);
nor U857 (N_857,N_708,N_779);
and U858 (N_858,N_707,N_761);
nand U859 (N_859,N_795,N_728);
nand U860 (N_860,N_769,N_780);
nor U861 (N_861,N_761,N_702);
nand U862 (N_862,N_748,N_799);
or U863 (N_863,N_751,N_746);
and U864 (N_864,N_792,N_774);
or U865 (N_865,N_721,N_703);
nand U866 (N_866,N_722,N_784);
nand U867 (N_867,N_795,N_798);
and U868 (N_868,N_720,N_728);
and U869 (N_869,N_747,N_770);
and U870 (N_870,N_730,N_722);
and U871 (N_871,N_726,N_756);
or U872 (N_872,N_715,N_710);
nor U873 (N_873,N_794,N_746);
nand U874 (N_874,N_702,N_744);
or U875 (N_875,N_719,N_738);
nand U876 (N_876,N_721,N_769);
nor U877 (N_877,N_706,N_799);
xor U878 (N_878,N_713,N_724);
or U879 (N_879,N_783,N_755);
nand U880 (N_880,N_784,N_736);
nor U881 (N_881,N_721,N_735);
nand U882 (N_882,N_767,N_720);
and U883 (N_883,N_769,N_774);
nand U884 (N_884,N_753,N_726);
and U885 (N_885,N_710,N_787);
nand U886 (N_886,N_721,N_793);
or U887 (N_887,N_715,N_707);
and U888 (N_888,N_748,N_781);
nand U889 (N_889,N_748,N_795);
nor U890 (N_890,N_736,N_768);
nor U891 (N_891,N_719,N_785);
nor U892 (N_892,N_721,N_723);
xor U893 (N_893,N_735,N_736);
nor U894 (N_894,N_723,N_769);
nor U895 (N_895,N_709,N_702);
nor U896 (N_896,N_778,N_745);
nor U897 (N_897,N_786,N_759);
and U898 (N_898,N_776,N_732);
and U899 (N_899,N_749,N_776);
and U900 (N_900,N_836,N_870);
nor U901 (N_901,N_864,N_896);
nand U902 (N_902,N_822,N_898);
and U903 (N_903,N_832,N_812);
nor U904 (N_904,N_853,N_897);
and U905 (N_905,N_804,N_820);
nand U906 (N_906,N_841,N_878);
nor U907 (N_907,N_852,N_858);
or U908 (N_908,N_844,N_875);
or U909 (N_909,N_816,N_879);
and U910 (N_910,N_838,N_866);
and U911 (N_911,N_803,N_800);
and U912 (N_912,N_885,N_839);
nor U913 (N_913,N_846,N_842);
xor U914 (N_914,N_821,N_865);
nand U915 (N_915,N_880,N_833);
xnor U916 (N_916,N_881,N_891);
nand U917 (N_917,N_869,N_801);
and U918 (N_918,N_817,N_888);
or U919 (N_919,N_835,N_863);
or U920 (N_920,N_855,N_894);
and U921 (N_921,N_807,N_882);
nor U922 (N_922,N_868,N_819);
nand U923 (N_923,N_861,N_830);
or U924 (N_924,N_840,N_872);
and U925 (N_925,N_854,N_828);
nor U926 (N_926,N_808,N_825);
and U927 (N_927,N_890,N_826);
nand U928 (N_928,N_887,N_843);
or U929 (N_929,N_893,N_815);
or U930 (N_930,N_892,N_862);
or U931 (N_931,N_810,N_813);
nand U932 (N_932,N_829,N_823);
or U933 (N_933,N_857,N_895);
or U934 (N_934,N_876,N_851);
nand U935 (N_935,N_873,N_834);
or U936 (N_936,N_847,N_859);
nor U937 (N_937,N_871,N_856);
nor U938 (N_938,N_818,N_849);
nand U939 (N_939,N_831,N_824);
nor U940 (N_940,N_874,N_809);
nor U941 (N_941,N_848,N_805);
xor U942 (N_942,N_802,N_877);
and U943 (N_943,N_806,N_860);
nor U944 (N_944,N_883,N_845);
or U945 (N_945,N_867,N_814);
and U946 (N_946,N_886,N_837);
nor U947 (N_947,N_884,N_811);
or U948 (N_948,N_889,N_899);
nand U949 (N_949,N_827,N_850);
or U950 (N_950,N_874,N_819);
nand U951 (N_951,N_852,N_873);
and U952 (N_952,N_811,N_849);
or U953 (N_953,N_824,N_862);
nor U954 (N_954,N_895,N_891);
or U955 (N_955,N_858,N_881);
or U956 (N_956,N_830,N_839);
or U957 (N_957,N_889,N_878);
nand U958 (N_958,N_875,N_853);
nor U959 (N_959,N_870,N_888);
nand U960 (N_960,N_822,N_829);
xor U961 (N_961,N_824,N_871);
nand U962 (N_962,N_855,N_847);
xor U963 (N_963,N_851,N_883);
and U964 (N_964,N_821,N_846);
xnor U965 (N_965,N_886,N_810);
and U966 (N_966,N_822,N_834);
nand U967 (N_967,N_846,N_806);
nor U968 (N_968,N_803,N_869);
xor U969 (N_969,N_823,N_820);
nand U970 (N_970,N_856,N_833);
nor U971 (N_971,N_856,N_835);
or U972 (N_972,N_820,N_826);
and U973 (N_973,N_871,N_803);
nor U974 (N_974,N_869,N_812);
nand U975 (N_975,N_833,N_893);
nand U976 (N_976,N_878,N_853);
and U977 (N_977,N_816,N_839);
nor U978 (N_978,N_840,N_877);
nor U979 (N_979,N_823,N_874);
nand U980 (N_980,N_851,N_802);
and U981 (N_981,N_842,N_823);
nor U982 (N_982,N_806,N_878);
nor U983 (N_983,N_860,N_853);
nor U984 (N_984,N_845,N_822);
and U985 (N_985,N_823,N_839);
nor U986 (N_986,N_814,N_804);
xor U987 (N_987,N_886,N_876);
or U988 (N_988,N_885,N_834);
and U989 (N_989,N_848,N_808);
nor U990 (N_990,N_893,N_829);
or U991 (N_991,N_898,N_839);
nand U992 (N_992,N_848,N_815);
and U993 (N_993,N_845,N_852);
nor U994 (N_994,N_870,N_865);
xnor U995 (N_995,N_845,N_868);
or U996 (N_996,N_835,N_810);
and U997 (N_997,N_867,N_827);
or U998 (N_998,N_897,N_827);
nor U999 (N_999,N_877,N_831);
and U1000 (N_1000,N_985,N_923);
nor U1001 (N_1001,N_946,N_940);
xnor U1002 (N_1002,N_975,N_980);
and U1003 (N_1003,N_922,N_939);
nor U1004 (N_1004,N_915,N_996);
and U1005 (N_1005,N_929,N_974);
or U1006 (N_1006,N_943,N_932);
nor U1007 (N_1007,N_966,N_944);
and U1008 (N_1008,N_977,N_987);
and U1009 (N_1009,N_907,N_913);
or U1010 (N_1010,N_901,N_994);
and U1011 (N_1011,N_935,N_903);
nand U1012 (N_1012,N_937,N_954);
xor U1013 (N_1013,N_941,N_970);
or U1014 (N_1014,N_993,N_953);
nor U1015 (N_1015,N_908,N_938);
and U1016 (N_1016,N_917,N_955);
and U1017 (N_1017,N_968,N_900);
xnor U1018 (N_1018,N_918,N_927);
or U1019 (N_1019,N_902,N_995);
nand U1020 (N_1020,N_920,N_965);
nand U1021 (N_1021,N_919,N_961);
nor U1022 (N_1022,N_969,N_916);
nand U1023 (N_1023,N_924,N_958);
or U1024 (N_1024,N_982,N_992);
and U1025 (N_1025,N_959,N_921);
and U1026 (N_1026,N_971,N_952);
xor U1027 (N_1027,N_960,N_910);
and U1028 (N_1028,N_991,N_986);
xnor U1029 (N_1029,N_978,N_989);
and U1030 (N_1030,N_911,N_936);
or U1031 (N_1031,N_925,N_972);
or U1032 (N_1032,N_949,N_999);
xnor U1033 (N_1033,N_983,N_957);
xnor U1034 (N_1034,N_909,N_945);
or U1035 (N_1035,N_979,N_981);
and U1036 (N_1036,N_933,N_984);
xor U1037 (N_1037,N_964,N_904);
nand U1038 (N_1038,N_928,N_998);
and U1039 (N_1039,N_942,N_990);
or U1040 (N_1040,N_973,N_997);
and U1041 (N_1041,N_951,N_948);
nand U1042 (N_1042,N_947,N_930);
nor U1043 (N_1043,N_950,N_926);
nand U1044 (N_1044,N_976,N_906);
and U1045 (N_1045,N_967,N_963);
xor U1046 (N_1046,N_914,N_962);
and U1047 (N_1047,N_934,N_905);
or U1048 (N_1048,N_988,N_931);
nand U1049 (N_1049,N_956,N_912);
xnor U1050 (N_1050,N_996,N_959);
nand U1051 (N_1051,N_971,N_951);
and U1052 (N_1052,N_962,N_916);
xnor U1053 (N_1053,N_901,N_937);
or U1054 (N_1054,N_985,N_949);
nor U1055 (N_1055,N_915,N_962);
xor U1056 (N_1056,N_901,N_930);
and U1057 (N_1057,N_907,N_977);
nor U1058 (N_1058,N_984,N_904);
nor U1059 (N_1059,N_983,N_920);
nand U1060 (N_1060,N_904,N_973);
or U1061 (N_1061,N_948,N_977);
and U1062 (N_1062,N_993,N_931);
nand U1063 (N_1063,N_946,N_952);
xnor U1064 (N_1064,N_971,N_937);
nand U1065 (N_1065,N_921,N_925);
nor U1066 (N_1066,N_997,N_941);
and U1067 (N_1067,N_920,N_940);
nand U1068 (N_1068,N_990,N_998);
and U1069 (N_1069,N_928,N_952);
or U1070 (N_1070,N_948,N_979);
and U1071 (N_1071,N_974,N_991);
nor U1072 (N_1072,N_994,N_996);
xnor U1073 (N_1073,N_995,N_958);
nand U1074 (N_1074,N_920,N_988);
nand U1075 (N_1075,N_996,N_991);
xor U1076 (N_1076,N_908,N_963);
nand U1077 (N_1077,N_906,N_944);
nand U1078 (N_1078,N_967,N_975);
nand U1079 (N_1079,N_917,N_985);
and U1080 (N_1080,N_915,N_930);
nor U1081 (N_1081,N_919,N_900);
nand U1082 (N_1082,N_995,N_984);
nand U1083 (N_1083,N_929,N_985);
nor U1084 (N_1084,N_955,N_931);
or U1085 (N_1085,N_931,N_962);
or U1086 (N_1086,N_973,N_951);
xnor U1087 (N_1087,N_977,N_951);
or U1088 (N_1088,N_908,N_949);
nor U1089 (N_1089,N_915,N_916);
nand U1090 (N_1090,N_943,N_944);
and U1091 (N_1091,N_910,N_967);
nor U1092 (N_1092,N_939,N_927);
and U1093 (N_1093,N_948,N_935);
nand U1094 (N_1094,N_923,N_982);
nor U1095 (N_1095,N_917,N_967);
nand U1096 (N_1096,N_990,N_968);
or U1097 (N_1097,N_924,N_943);
nand U1098 (N_1098,N_976,N_991);
and U1099 (N_1099,N_938,N_946);
and U1100 (N_1100,N_1041,N_1001);
nor U1101 (N_1101,N_1062,N_1066);
nand U1102 (N_1102,N_1074,N_1000);
nand U1103 (N_1103,N_1077,N_1016);
nor U1104 (N_1104,N_1035,N_1009);
nand U1105 (N_1105,N_1068,N_1025);
nor U1106 (N_1106,N_1052,N_1048);
or U1107 (N_1107,N_1013,N_1055);
xnor U1108 (N_1108,N_1007,N_1004);
or U1109 (N_1109,N_1039,N_1020);
and U1110 (N_1110,N_1033,N_1056);
and U1111 (N_1111,N_1096,N_1046);
and U1112 (N_1112,N_1070,N_1085);
and U1113 (N_1113,N_1022,N_1099);
nand U1114 (N_1114,N_1042,N_1011);
nor U1115 (N_1115,N_1081,N_1019);
nor U1116 (N_1116,N_1026,N_1044);
or U1117 (N_1117,N_1092,N_1023);
xnor U1118 (N_1118,N_1031,N_1061);
or U1119 (N_1119,N_1008,N_1036);
nand U1120 (N_1120,N_1065,N_1053);
nor U1121 (N_1121,N_1021,N_1034);
or U1122 (N_1122,N_1091,N_1075);
or U1123 (N_1123,N_1029,N_1010);
or U1124 (N_1124,N_1082,N_1076);
nor U1125 (N_1125,N_1038,N_1006);
nand U1126 (N_1126,N_1086,N_1064);
or U1127 (N_1127,N_1043,N_1071);
nand U1128 (N_1128,N_1087,N_1017);
xnor U1129 (N_1129,N_1051,N_1024);
or U1130 (N_1130,N_1049,N_1067);
and U1131 (N_1131,N_1028,N_1037);
nand U1132 (N_1132,N_1059,N_1018);
nor U1133 (N_1133,N_1003,N_1083);
and U1134 (N_1134,N_1047,N_1088);
or U1135 (N_1135,N_1094,N_1045);
and U1136 (N_1136,N_1079,N_1090);
nand U1137 (N_1137,N_1095,N_1063);
and U1138 (N_1138,N_1073,N_1084);
or U1139 (N_1139,N_1015,N_1060);
xor U1140 (N_1140,N_1005,N_1014);
and U1141 (N_1141,N_1089,N_1097);
and U1142 (N_1142,N_1050,N_1093);
and U1143 (N_1143,N_1012,N_1002);
nand U1144 (N_1144,N_1072,N_1040);
and U1145 (N_1145,N_1098,N_1069);
nand U1146 (N_1146,N_1032,N_1027);
nand U1147 (N_1147,N_1078,N_1057);
or U1148 (N_1148,N_1080,N_1054);
nor U1149 (N_1149,N_1058,N_1030);
or U1150 (N_1150,N_1078,N_1071);
nor U1151 (N_1151,N_1001,N_1022);
nor U1152 (N_1152,N_1011,N_1080);
or U1153 (N_1153,N_1094,N_1011);
or U1154 (N_1154,N_1041,N_1040);
nor U1155 (N_1155,N_1070,N_1035);
nand U1156 (N_1156,N_1099,N_1045);
and U1157 (N_1157,N_1063,N_1085);
and U1158 (N_1158,N_1013,N_1004);
nor U1159 (N_1159,N_1056,N_1055);
or U1160 (N_1160,N_1070,N_1012);
nand U1161 (N_1161,N_1063,N_1091);
or U1162 (N_1162,N_1086,N_1080);
or U1163 (N_1163,N_1036,N_1034);
nor U1164 (N_1164,N_1072,N_1063);
and U1165 (N_1165,N_1001,N_1018);
and U1166 (N_1166,N_1005,N_1093);
and U1167 (N_1167,N_1051,N_1077);
nand U1168 (N_1168,N_1040,N_1026);
and U1169 (N_1169,N_1048,N_1077);
and U1170 (N_1170,N_1067,N_1066);
nand U1171 (N_1171,N_1032,N_1022);
nand U1172 (N_1172,N_1072,N_1042);
nand U1173 (N_1173,N_1081,N_1023);
and U1174 (N_1174,N_1097,N_1034);
and U1175 (N_1175,N_1060,N_1024);
and U1176 (N_1176,N_1057,N_1044);
xnor U1177 (N_1177,N_1059,N_1001);
or U1178 (N_1178,N_1032,N_1041);
xor U1179 (N_1179,N_1007,N_1091);
nor U1180 (N_1180,N_1047,N_1063);
nor U1181 (N_1181,N_1052,N_1082);
xor U1182 (N_1182,N_1074,N_1033);
nor U1183 (N_1183,N_1042,N_1057);
nor U1184 (N_1184,N_1050,N_1099);
and U1185 (N_1185,N_1024,N_1053);
xor U1186 (N_1186,N_1022,N_1080);
nand U1187 (N_1187,N_1063,N_1053);
or U1188 (N_1188,N_1020,N_1037);
or U1189 (N_1189,N_1091,N_1085);
and U1190 (N_1190,N_1002,N_1011);
and U1191 (N_1191,N_1074,N_1030);
or U1192 (N_1192,N_1052,N_1046);
nor U1193 (N_1193,N_1063,N_1070);
nand U1194 (N_1194,N_1028,N_1067);
nand U1195 (N_1195,N_1018,N_1037);
nor U1196 (N_1196,N_1056,N_1052);
nor U1197 (N_1197,N_1032,N_1037);
nor U1198 (N_1198,N_1063,N_1097);
and U1199 (N_1199,N_1018,N_1004);
and U1200 (N_1200,N_1126,N_1190);
or U1201 (N_1201,N_1121,N_1189);
xor U1202 (N_1202,N_1191,N_1157);
and U1203 (N_1203,N_1137,N_1101);
nand U1204 (N_1204,N_1106,N_1109);
xnor U1205 (N_1205,N_1135,N_1100);
nor U1206 (N_1206,N_1139,N_1177);
nor U1207 (N_1207,N_1174,N_1134);
nor U1208 (N_1208,N_1182,N_1130);
nand U1209 (N_1209,N_1199,N_1144);
nor U1210 (N_1210,N_1183,N_1119);
nor U1211 (N_1211,N_1112,N_1195);
and U1212 (N_1212,N_1103,N_1165);
or U1213 (N_1213,N_1151,N_1154);
and U1214 (N_1214,N_1133,N_1198);
nor U1215 (N_1215,N_1128,N_1170);
xnor U1216 (N_1216,N_1188,N_1107);
nor U1217 (N_1217,N_1132,N_1163);
nor U1218 (N_1218,N_1131,N_1152);
nor U1219 (N_1219,N_1113,N_1122);
xor U1220 (N_1220,N_1155,N_1184);
and U1221 (N_1221,N_1172,N_1197);
xor U1222 (N_1222,N_1173,N_1111);
xnor U1223 (N_1223,N_1160,N_1196);
and U1224 (N_1224,N_1114,N_1115);
or U1225 (N_1225,N_1176,N_1149);
or U1226 (N_1226,N_1166,N_1141);
nor U1227 (N_1227,N_1104,N_1178);
and U1228 (N_1228,N_1105,N_1142);
xnor U1229 (N_1229,N_1148,N_1120);
nor U1230 (N_1230,N_1118,N_1192);
and U1231 (N_1231,N_1169,N_1124);
or U1232 (N_1232,N_1167,N_1147);
and U1233 (N_1233,N_1168,N_1110);
nand U1234 (N_1234,N_1180,N_1145);
nand U1235 (N_1235,N_1164,N_1138);
nand U1236 (N_1236,N_1171,N_1146);
and U1237 (N_1237,N_1161,N_1158);
nor U1238 (N_1238,N_1116,N_1162);
xnor U1239 (N_1239,N_1175,N_1194);
or U1240 (N_1240,N_1117,N_1193);
and U1241 (N_1241,N_1159,N_1136);
nand U1242 (N_1242,N_1129,N_1140);
and U1243 (N_1243,N_1186,N_1123);
nand U1244 (N_1244,N_1181,N_1153);
nand U1245 (N_1245,N_1185,N_1127);
or U1246 (N_1246,N_1187,N_1150);
nand U1247 (N_1247,N_1108,N_1179);
nor U1248 (N_1248,N_1156,N_1143);
or U1249 (N_1249,N_1125,N_1102);
and U1250 (N_1250,N_1154,N_1117);
or U1251 (N_1251,N_1163,N_1126);
nor U1252 (N_1252,N_1161,N_1171);
or U1253 (N_1253,N_1199,N_1123);
nor U1254 (N_1254,N_1147,N_1199);
and U1255 (N_1255,N_1132,N_1175);
or U1256 (N_1256,N_1133,N_1125);
nor U1257 (N_1257,N_1139,N_1186);
or U1258 (N_1258,N_1165,N_1121);
nand U1259 (N_1259,N_1141,N_1179);
and U1260 (N_1260,N_1136,N_1161);
nor U1261 (N_1261,N_1181,N_1126);
or U1262 (N_1262,N_1141,N_1123);
or U1263 (N_1263,N_1105,N_1112);
nor U1264 (N_1264,N_1107,N_1129);
or U1265 (N_1265,N_1170,N_1134);
nand U1266 (N_1266,N_1109,N_1165);
or U1267 (N_1267,N_1149,N_1157);
and U1268 (N_1268,N_1190,N_1132);
nor U1269 (N_1269,N_1140,N_1175);
nand U1270 (N_1270,N_1147,N_1124);
nor U1271 (N_1271,N_1124,N_1144);
nand U1272 (N_1272,N_1194,N_1139);
and U1273 (N_1273,N_1153,N_1130);
nand U1274 (N_1274,N_1180,N_1164);
nand U1275 (N_1275,N_1197,N_1128);
xor U1276 (N_1276,N_1199,N_1143);
or U1277 (N_1277,N_1189,N_1126);
nand U1278 (N_1278,N_1189,N_1120);
nand U1279 (N_1279,N_1185,N_1180);
and U1280 (N_1280,N_1154,N_1145);
and U1281 (N_1281,N_1183,N_1180);
and U1282 (N_1282,N_1187,N_1112);
nand U1283 (N_1283,N_1151,N_1127);
or U1284 (N_1284,N_1163,N_1181);
nand U1285 (N_1285,N_1124,N_1159);
or U1286 (N_1286,N_1148,N_1160);
and U1287 (N_1287,N_1169,N_1111);
nor U1288 (N_1288,N_1100,N_1114);
nand U1289 (N_1289,N_1118,N_1125);
and U1290 (N_1290,N_1116,N_1121);
nor U1291 (N_1291,N_1136,N_1140);
xnor U1292 (N_1292,N_1192,N_1124);
or U1293 (N_1293,N_1183,N_1198);
nand U1294 (N_1294,N_1139,N_1126);
nor U1295 (N_1295,N_1166,N_1190);
nor U1296 (N_1296,N_1137,N_1125);
nand U1297 (N_1297,N_1100,N_1140);
and U1298 (N_1298,N_1158,N_1165);
and U1299 (N_1299,N_1148,N_1134);
or U1300 (N_1300,N_1209,N_1226);
and U1301 (N_1301,N_1208,N_1228);
or U1302 (N_1302,N_1269,N_1241);
or U1303 (N_1303,N_1256,N_1232);
xnor U1304 (N_1304,N_1267,N_1294);
or U1305 (N_1305,N_1246,N_1275);
nor U1306 (N_1306,N_1218,N_1274);
nand U1307 (N_1307,N_1252,N_1293);
or U1308 (N_1308,N_1236,N_1213);
and U1309 (N_1309,N_1263,N_1255);
nor U1310 (N_1310,N_1250,N_1235);
nand U1311 (N_1311,N_1272,N_1227);
xnor U1312 (N_1312,N_1262,N_1238);
or U1313 (N_1313,N_1230,N_1257);
xnor U1314 (N_1314,N_1289,N_1215);
or U1315 (N_1315,N_1265,N_1271);
or U1316 (N_1316,N_1247,N_1225);
nor U1317 (N_1317,N_1212,N_1281);
nand U1318 (N_1318,N_1251,N_1299);
or U1319 (N_1319,N_1268,N_1260);
xor U1320 (N_1320,N_1237,N_1243);
nor U1321 (N_1321,N_1234,N_1203);
and U1322 (N_1322,N_1277,N_1290);
or U1323 (N_1323,N_1282,N_1258);
nand U1324 (N_1324,N_1222,N_1292);
nand U1325 (N_1325,N_1286,N_1221);
or U1326 (N_1326,N_1204,N_1242);
or U1327 (N_1327,N_1210,N_1223);
and U1328 (N_1328,N_1291,N_1261);
nand U1329 (N_1329,N_1216,N_1280);
or U1330 (N_1330,N_1295,N_1287);
nand U1331 (N_1331,N_1244,N_1285);
nor U1332 (N_1332,N_1201,N_1219);
nor U1333 (N_1333,N_1284,N_1254);
or U1334 (N_1334,N_1239,N_1224);
nor U1335 (N_1335,N_1266,N_1214);
xnor U1336 (N_1336,N_1264,N_1200);
nor U1337 (N_1337,N_1276,N_1245);
xnor U1338 (N_1338,N_1253,N_1259);
and U1339 (N_1339,N_1270,N_1297);
nand U1340 (N_1340,N_1296,N_1220);
nor U1341 (N_1341,N_1217,N_1233);
nor U1342 (N_1342,N_1202,N_1279);
and U1343 (N_1343,N_1248,N_1207);
or U1344 (N_1344,N_1211,N_1288);
or U1345 (N_1345,N_1231,N_1273);
xnor U1346 (N_1346,N_1249,N_1278);
or U1347 (N_1347,N_1283,N_1206);
nor U1348 (N_1348,N_1298,N_1205);
xor U1349 (N_1349,N_1240,N_1229);
nand U1350 (N_1350,N_1265,N_1243);
nand U1351 (N_1351,N_1226,N_1288);
nor U1352 (N_1352,N_1291,N_1265);
and U1353 (N_1353,N_1265,N_1288);
and U1354 (N_1354,N_1223,N_1281);
nand U1355 (N_1355,N_1234,N_1245);
xnor U1356 (N_1356,N_1267,N_1247);
and U1357 (N_1357,N_1238,N_1288);
or U1358 (N_1358,N_1226,N_1214);
nand U1359 (N_1359,N_1236,N_1296);
or U1360 (N_1360,N_1260,N_1211);
and U1361 (N_1361,N_1200,N_1221);
or U1362 (N_1362,N_1293,N_1220);
nand U1363 (N_1363,N_1208,N_1276);
or U1364 (N_1364,N_1232,N_1274);
and U1365 (N_1365,N_1244,N_1265);
nor U1366 (N_1366,N_1290,N_1217);
nand U1367 (N_1367,N_1259,N_1257);
nor U1368 (N_1368,N_1261,N_1273);
and U1369 (N_1369,N_1276,N_1294);
or U1370 (N_1370,N_1247,N_1285);
or U1371 (N_1371,N_1291,N_1222);
xor U1372 (N_1372,N_1246,N_1201);
nor U1373 (N_1373,N_1204,N_1249);
nand U1374 (N_1374,N_1268,N_1275);
or U1375 (N_1375,N_1217,N_1207);
or U1376 (N_1376,N_1252,N_1297);
nand U1377 (N_1377,N_1224,N_1211);
and U1378 (N_1378,N_1210,N_1209);
nand U1379 (N_1379,N_1259,N_1268);
nand U1380 (N_1380,N_1204,N_1241);
nand U1381 (N_1381,N_1225,N_1270);
nand U1382 (N_1382,N_1278,N_1283);
nand U1383 (N_1383,N_1275,N_1224);
or U1384 (N_1384,N_1262,N_1212);
and U1385 (N_1385,N_1267,N_1244);
or U1386 (N_1386,N_1245,N_1289);
nand U1387 (N_1387,N_1233,N_1230);
nand U1388 (N_1388,N_1244,N_1251);
or U1389 (N_1389,N_1297,N_1267);
nor U1390 (N_1390,N_1219,N_1257);
or U1391 (N_1391,N_1266,N_1202);
or U1392 (N_1392,N_1240,N_1245);
or U1393 (N_1393,N_1227,N_1245);
nand U1394 (N_1394,N_1227,N_1208);
or U1395 (N_1395,N_1294,N_1284);
or U1396 (N_1396,N_1259,N_1229);
or U1397 (N_1397,N_1245,N_1201);
and U1398 (N_1398,N_1232,N_1205);
nor U1399 (N_1399,N_1218,N_1288);
nand U1400 (N_1400,N_1365,N_1395);
xnor U1401 (N_1401,N_1327,N_1332);
nor U1402 (N_1402,N_1324,N_1388);
nand U1403 (N_1403,N_1356,N_1335);
and U1404 (N_1404,N_1399,N_1330);
nand U1405 (N_1405,N_1345,N_1381);
or U1406 (N_1406,N_1385,N_1340);
nand U1407 (N_1407,N_1306,N_1316);
or U1408 (N_1408,N_1331,N_1361);
xor U1409 (N_1409,N_1338,N_1370);
or U1410 (N_1410,N_1337,N_1379);
xnor U1411 (N_1411,N_1367,N_1373);
or U1412 (N_1412,N_1344,N_1383);
or U1413 (N_1413,N_1359,N_1329);
and U1414 (N_1414,N_1378,N_1302);
nor U1415 (N_1415,N_1348,N_1339);
nand U1416 (N_1416,N_1328,N_1326);
or U1417 (N_1417,N_1387,N_1342);
or U1418 (N_1418,N_1375,N_1369);
xnor U1419 (N_1419,N_1374,N_1386);
nand U1420 (N_1420,N_1393,N_1310);
nand U1421 (N_1421,N_1300,N_1347);
nand U1422 (N_1422,N_1391,N_1308);
nand U1423 (N_1423,N_1355,N_1382);
and U1424 (N_1424,N_1318,N_1351);
nand U1425 (N_1425,N_1349,N_1320);
nand U1426 (N_1426,N_1305,N_1309);
nand U1427 (N_1427,N_1392,N_1363);
nand U1428 (N_1428,N_1353,N_1376);
or U1429 (N_1429,N_1372,N_1312);
or U1430 (N_1430,N_1319,N_1377);
or U1431 (N_1431,N_1390,N_1304);
nor U1432 (N_1432,N_1317,N_1389);
or U1433 (N_1433,N_1336,N_1314);
nand U1434 (N_1434,N_1311,N_1364);
or U1435 (N_1435,N_1357,N_1313);
and U1436 (N_1436,N_1301,N_1398);
and U1437 (N_1437,N_1384,N_1368);
or U1438 (N_1438,N_1371,N_1307);
nand U1439 (N_1439,N_1397,N_1396);
or U1440 (N_1440,N_1322,N_1360);
or U1441 (N_1441,N_1334,N_1354);
or U1442 (N_1442,N_1362,N_1315);
nand U1443 (N_1443,N_1323,N_1352);
or U1444 (N_1444,N_1333,N_1350);
xnor U1445 (N_1445,N_1341,N_1394);
nor U1446 (N_1446,N_1303,N_1343);
or U1447 (N_1447,N_1321,N_1366);
nand U1448 (N_1448,N_1358,N_1325);
and U1449 (N_1449,N_1380,N_1346);
or U1450 (N_1450,N_1329,N_1368);
nand U1451 (N_1451,N_1320,N_1343);
nand U1452 (N_1452,N_1359,N_1309);
xnor U1453 (N_1453,N_1356,N_1363);
and U1454 (N_1454,N_1337,N_1320);
nand U1455 (N_1455,N_1361,N_1347);
nand U1456 (N_1456,N_1364,N_1396);
nand U1457 (N_1457,N_1390,N_1364);
xnor U1458 (N_1458,N_1328,N_1378);
xor U1459 (N_1459,N_1378,N_1396);
nor U1460 (N_1460,N_1301,N_1372);
nand U1461 (N_1461,N_1375,N_1303);
and U1462 (N_1462,N_1351,N_1352);
nor U1463 (N_1463,N_1320,N_1367);
nor U1464 (N_1464,N_1317,N_1370);
or U1465 (N_1465,N_1342,N_1368);
or U1466 (N_1466,N_1398,N_1397);
and U1467 (N_1467,N_1311,N_1331);
nand U1468 (N_1468,N_1378,N_1352);
and U1469 (N_1469,N_1335,N_1353);
or U1470 (N_1470,N_1309,N_1321);
and U1471 (N_1471,N_1372,N_1371);
nor U1472 (N_1472,N_1378,N_1341);
or U1473 (N_1473,N_1346,N_1386);
and U1474 (N_1474,N_1394,N_1301);
nor U1475 (N_1475,N_1364,N_1332);
or U1476 (N_1476,N_1336,N_1338);
or U1477 (N_1477,N_1381,N_1315);
or U1478 (N_1478,N_1388,N_1326);
or U1479 (N_1479,N_1357,N_1366);
nand U1480 (N_1480,N_1300,N_1339);
or U1481 (N_1481,N_1325,N_1374);
and U1482 (N_1482,N_1398,N_1349);
nor U1483 (N_1483,N_1306,N_1374);
nand U1484 (N_1484,N_1305,N_1349);
nor U1485 (N_1485,N_1366,N_1331);
nor U1486 (N_1486,N_1398,N_1375);
or U1487 (N_1487,N_1379,N_1326);
or U1488 (N_1488,N_1373,N_1365);
or U1489 (N_1489,N_1314,N_1355);
or U1490 (N_1490,N_1318,N_1373);
and U1491 (N_1491,N_1359,N_1396);
and U1492 (N_1492,N_1307,N_1360);
nor U1493 (N_1493,N_1396,N_1384);
or U1494 (N_1494,N_1386,N_1370);
nor U1495 (N_1495,N_1383,N_1319);
nor U1496 (N_1496,N_1321,N_1316);
nand U1497 (N_1497,N_1386,N_1308);
nor U1498 (N_1498,N_1334,N_1350);
and U1499 (N_1499,N_1391,N_1327);
and U1500 (N_1500,N_1463,N_1407);
or U1501 (N_1501,N_1433,N_1471);
nand U1502 (N_1502,N_1414,N_1455);
or U1503 (N_1503,N_1495,N_1402);
or U1504 (N_1504,N_1469,N_1490);
nor U1505 (N_1505,N_1400,N_1410);
xor U1506 (N_1506,N_1441,N_1432);
nor U1507 (N_1507,N_1448,N_1484);
and U1508 (N_1508,N_1445,N_1419);
xnor U1509 (N_1509,N_1461,N_1435);
and U1510 (N_1510,N_1417,N_1440);
nand U1511 (N_1511,N_1439,N_1493);
nor U1512 (N_1512,N_1423,N_1498);
xnor U1513 (N_1513,N_1470,N_1497);
nor U1514 (N_1514,N_1427,N_1460);
xor U1515 (N_1515,N_1456,N_1476);
or U1516 (N_1516,N_1483,N_1450);
or U1517 (N_1517,N_1425,N_1466);
nor U1518 (N_1518,N_1465,N_1412);
xnor U1519 (N_1519,N_1447,N_1485);
nand U1520 (N_1520,N_1437,N_1473);
or U1521 (N_1521,N_1475,N_1442);
nor U1522 (N_1522,N_1472,N_1446);
and U1523 (N_1523,N_1426,N_1406);
nor U1524 (N_1524,N_1492,N_1494);
nand U1525 (N_1525,N_1457,N_1474);
xor U1526 (N_1526,N_1428,N_1487);
or U1527 (N_1527,N_1420,N_1413);
and U1528 (N_1528,N_1444,N_1449);
or U1529 (N_1529,N_1422,N_1409);
and U1530 (N_1530,N_1421,N_1411);
xnor U1531 (N_1531,N_1464,N_1452);
nor U1532 (N_1532,N_1479,N_1416);
nor U1533 (N_1533,N_1438,N_1401);
nor U1534 (N_1534,N_1415,N_1458);
nand U1535 (N_1535,N_1405,N_1403);
nor U1536 (N_1536,N_1467,N_1454);
nand U1537 (N_1537,N_1486,N_1404);
nand U1538 (N_1538,N_1443,N_1482);
nor U1539 (N_1539,N_1491,N_1434);
and U1540 (N_1540,N_1436,N_1489);
and U1541 (N_1541,N_1459,N_1480);
xor U1542 (N_1542,N_1424,N_1496);
or U1543 (N_1543,N_1431,N_1481);
xnor U1544 (N_1544,N_1430,N_1453);
and U1545 (N_1545,N_1478,N_1488);
or U1546 (N_1546,N_1451,N_1462);
nand U1547 (N_1547,N_1408,N_1418);
or U1548 (N_1548,N_1499,N_1429);
or U1549 (N_1549,N_1468,N_1477);
xnor U1550 (N_1550,N_1401,N_1493);
and U1551 (N_1551,N_1473,N_1494);
xor U1552 (N_1552,N_1463,N_1423);
or U1553 (N_1553,N_1445,N_1479);
nand U1554 (N_1554,N_1409,N_1425);
nor U1555 (N_1555,N_1416,N_1477);
or U1556 (N_1556,N_1488,N_1419);
nand U1557 (N_1557,N_1408,N_1480);
nand U1558 (N_1558,N_1414,N_1412);
nor U1559 (N_1559,N_1429,N_1447);
and U1560 (N_1560,N_1498,N_1418);
nor U1561 (N_1561,N_1469,N_1485);
nor U1562 (N_1562,N_1438,N_1410);
or U1563 (N_1563,N_1414,N_1460);
nor U1564 (N_1564,N_1493,N_1409);
or U1565 (N_1565,N_1424,N_1462);
or U1566 (N_1566,N_1421,N_1407);
or U1567 (N_1567,N_1423,N_1489);
xnor U1568 (N_1568,N_1407,N_1478);
or U1569 (N_1569,N_1422,N_1474);
nor U1570 (N_1570,N_1411,N_1486);
nor U1571 (N_1571,N_1458,N_1456);
nor U1572 (N_1572,N_1492,N_1496);
or U1573 (N_1573,N_1434,N_1413);
nor U1574 (N_1574,N_1434,N_1446);
nand U1575 (N_1575,N_1467,N_1433);
and U1576 (N_1576,N_1470,N_1420);
xnor U1577 (N_1577,N_1491,N_1415);
and U1578 (N_1578,N_1462,N_1404);
xor U1579 (N_1579,N_1498,N_1422);
and U1580 (N_1580,N_1416,N_1493);
nand U1581 (N_1581,N_1409,N_1437);
nand U1582 (N_1582,N_1430,N_1411);
xnor U1583 (N_1583,N_1437,N_1414);
nand U1584 (N_1584,N_1450,N_1472);
and U1585 (N_1585,N_1435,N_1470);
or U1586 (N_1586,N_1471,N_1487);
and U1587 (N_1587,N_1437,N_1404);
nor U1588 (N_1588,N_1428,N_1420);
nor U1589 (N_1589,N_1458,N_1485);
or U1590 (N_1590,N_1424,N_1448);
and U1591 (N_1591,N_1432,N_1413);
and U1592 (N_1592,N_1493,N_1488);
and U1593 (N_1593,N_1431,N_1440);
or U1594 (N_1594,N_1484,N_1441);
xnor U1595 (N_1595,N_1452,N_1419);
or U1596 (N_1596,N_1420,N_1435);
nor U1597 (N_1597,N_1406,N_1472);
nor U1598 (N_1598,N_1415,N_1406);
and U1599 (N_1599,N_1490,N_1441);
nor U1600 (N_1600,N_1561,N_1534);
or U1601 (N_1601,N_1595,N_1530);
nand U1602 (N_1602,N_1522,N_1528);
and U1603 (N_1603,N_1525,N_1501);
or U1604 (N_1604,N_1537,N_1564);
and U1605 (N_1605,N_1590,N_1541);
nand U1606 (N_1606,N_1588,N_1558);
and U1607 (N_1607,N_1524,N_1509);
nand U1608 (N_1608,N_1543,N_1547);
or U1609 (N_1609,N_1540,N_1569);
and U1610 (N_1610,N_1581,N_1553);
nand U1611 (N_1611,N_1503,N_1551);
nor U1612 (N_1612,N_1510,N_1531);
or U1613 (N_1613,N_1535,N_1532);
and U1614 (N_1614,N_1565,N_1527);
nor U1615 (N_1615,N_1533,N_1515);
xor U1616 (N_1616,N_1576,N_1512);
or U1617 (N_1617,N_1594,N_1545);
nand U1618 (N_1618,N_1566,N_1500);
nand U1619 (N_1619,N_1596,N_1507);
and U1620 (N_1620,N_1599,N_1587);
and U1621 (N_1621,N_1517,N_1560);
and U1622 (N_1622,N_1519,N_1578);
nand U1623 (N_1623,N_1567,N_1579);
or U1624 (N_1624,N_1518,N_1526);
nor U1625 (N_1625,N_1502,N_1570);
xnor U1626 (N_1626,N_1568,N_1555);
xor U1627 (N_1627,N_1556,N_1557);
nand U1628 (N_1628,N_1550,N_1506);
and U1629 (N_1629,N_1586,N_1589);
xor U1630 (N_1630,N_1574,N_1597);
or U1631 (N_1631,N_1592,N_1542);
or U1632 (N_1632,N_1571,N_1584);
and U1633 (N_1633,N_1577,N_1552);
nor U1634 (N_1634,N_1549,N_1554);
and U1635 (N_1635,N_1563,N_1582);
xnor U1636 (N_1636,N_1516,N_1575);
xnor U1637 (N_1637,N_1520,N_1513);
and U1638 (N_1638,N_1536,N_1539);
xnor U1639 (N_1639,N_1514,N_1544);
and U1640 (N_1640,N_1511,N_1559);
and U1641 (N_1641,N_1505,N_1591);
xnor U1642 (N_1642,N_1529,N_1508);
and U1643 (N_1643,N_1548,N_1593);
nor U1644 (N_1644,N_1504,N_1585);
nand U1645 (N_1645,N_1598,N_1562);
and U1646 (N_1646,N_1573,N_1523);
xor U1647 (N_1647,N_1546,N_1521);
and U1648 (N_1648,N_1538,N_1580);
and U1649 (N_1649,N_1572,N_1583);
nand U1650 (N_1650,N_1532,N_1543);
and U1651 (N_1651,N_1532,N_1588);
nor U1652 (N_1652,N_1570,N_1565);
or U1653 (N_1653,N_1529,N_1543);
or U1654 (N_1654,N_1505,N_1569);
nand U1655 (N_1655,N_1588,N_1534);
and U1656 (N_1656,N_1572,N_1593);
or U1657 (N_1657,N_1534,N_1579);
nand U1658 (N_1658,N_1507,N_1597);
or U1659 (N_1659,N_1596,N_1546);
and U1660 (N_1660,N_1570,N_1559);
nor U1661 (N_1661,N_1502,N_1521);
and U1662 (N_1662,N_1511,N_1567);
nand U1663 (N_1663,N_1513,N_1596);
and U1664 (N_1664,N_1573,N_1543);
xor U1665 (N_1665,N_1515,N_1508);
xnor U1666 (N_1666,N_1521,N_1506);
nor U1667 (N_1667,N_1572,N_1563);
or U1668 (N_1668,N_1596,N_1518);
and U1669 (N_1669,N_1580,N_1591);
or U1670 (N_1670,N_1513,N_1502);
nor U1671 (N_1671,N_1505,N_1577);
nand U1672 (N_1672,N_1512,N_1561);
nand U1673 (N_1673,N_1551,N_1526);
or U1674 (N_1674,N_1525,N_1549);
and U1675 (N_1675,N_1585,N_1541);
nand U1676 (N_1676,N_1570,N_1517);
and U1677 (N_1677,N_1532,N_1502);
or U1678 (N_1678,N_1592,N_1574);
and U1679 (N_1679,N_1504,N_1533);
nor U1680 (N_1680,N_1586,N_1529);
nor U1681 (N_1681,N_1522,N_1518);
or U1682 (N_1682,N_1565,N_1514);
nand U1683 (N_1683,N_1585,N_1574);
nand U1684 (N_1684,N_1584,N_1524);
and U1685 (N_1685,N_1506,N_1569);
and U1686 (N_1686,N_1547,N_1529);
nor U1687 (N_1687,N_1572,N_1592);
nand U1688 (N_1688,N_1542,N_1536);
xnor U1689 (N_1689,N_1577,N_1590);
nor U1690 (N_1690,N_1530,N_1552);
nor U1691 (N_1691,N_1580,N_1594);
or U1692 (N_1692,N_1596,N_1599);
nor U1693 (N_1693,N_1587,N_1557);
nor U1694 (N_1694,N_1500,N_1502);
and U1695 (N_1695,N_1506,N_1529);
and U1696 (N_1696,N_1560,N_1575);
nor U1697 (N_1697,N_1552,N_1554);
nor U1698 (N_1698,N_1551,N_1559);
and U1699 (N_1699,N_1583,N_1515);
and U1700 (N_1700,N_1696,N_1607);
nand U1701 (N_1701,N_1667,N_1650);
or U1702 (N_1702,N_1699,N_1602);
nand U1703 (N_1703,N_1606,N_1648);
nor U1704 (N_1704,N_1675,N_1661);
and U1705 (N_1705,N_1671,N_1639);
xor U1706 (N_1706,N_1621,N_1611);
and U1707 (N_1707,N_1681,N_1628);
and U1708 (N_1708,N_1614,N_1651);
or U1709 (N_1709,N_1687,N_1645);
nand U1710 (N_1710,N_1637,N_1672);
or U1711 (N_1711,N_1674,N_1643);
and U1712 (N_1712,N_1631,N_1619);
or U1713 (N_1713,N_1629,N_1601);
or U1714 (N_1714,N_1677,N_1657);
nand U1715 (N_1715,N_1647,N_1627);
or U1716 (N_1716,N_1689,N_1668);
nand U1717 (N_1717,N_1634,N_1633);
nor U1718 (N_1718,N_1603,N_1609);
nor U1719 (N_1719,N_1635,N_1623);
nand U1720 (N_1720,N_1698,N_1610);
nor U1721 (N_1721,N_1620,N_1659);
nand U1722 (N_1722,N_1605,N_1608);
and U1723 (N_1723,N_1646,N_1600);
nand U1724 (N_1724,N_1662,N_1697);
or U1725 (N_1725,N_1630,N_1618);
or U1726 (N_1726,N_1632,N_1694);
nor U1727 (N_1727,N_1652,N_1624);
xnor U1728 (N_1728,N_1679,N_1684);
nand U1729 (N_1729,N_1626,N_1612);
nand U1730 (N_1730,N_1693,N_1666);
or U1731 (N_1731,N_1655,N_1682);
and U1732 (N_1732,N_1670,N_1636);
and U1733 (N_1733,N_1641,N_1669);
nand U1734 (N_1734,N_1680,N_1663);
xnor U1735 (N_1735,N_1653,N_1683);
nand U1736 (N_1736,N_1695,N_1673);
nor U1737 (N_1737,N_1649,N_1678);
and U1738 (N_1738,N_1616,N_1686);
nor U1739 (N_1739,N_1656,N_1604);
xnor U1740 (N_1740,N_1615,N_1660);
nand U1741 (N_1741,N_1638,N_1622);
nor U1742 (N_1742,N_1685,N_1644);
and U1743 (N_1743,N_1617,N_1642);
and U1744 (N_1744,N_1690,N_1654);
nand U1745 (N_1745,N_1688,N_1676);
or U1746 (N_1746,N_1692,N_1658);
and U1747 (N_1747,N_1665,N_1613);
or U1748 (N_1748,N_1625,N_1664);
nand U1749 (N_1749,N_1691,N_1640);
or U1750 (N_1750,N_1664,N_1661);
xnor U1751 (N_1751,N_1617,N_1624);
nor U1752 (N_1752,N_1647,N_1602);
and U1753 (N_1753,N_1647,N_1621);
and U1754 (N_1754,N_1670,N_1682);
or U1755 (N_1755,N_1645,N_1682);
and U1756 (N_1756,N_1650,N_1624);
nand U1757 (N_1757,N_1618,N_1685);
nor U1758 (N_1758,N_1673,N_1610);
nand U1759 (N_1759,N_1691,N_1698);
or U1760 (N_1760,N_1655,N_1675);
nand U1761 (N_1761,N_1666,N_1626);
and U1762 (N_1762,N_1642,N_1629);
or U1763 (N_1763,N_1607,N_1637);
and U1764 (N_1764,N_1660,N_1637);
nor U1765 (N_1765,N_1664,N_1687);
nand U1766 (N_1766,N_1645,N_1658);
or U1767 (N_1767,N_1600,N_1636);
and U1768 (N_1768,N_1692,N_1646);
xnor U1769 (N_1769,N_1681,N_1630);
nor U1770 (N_1770,N_1675,N_1682);
and U1771 (N_1771,N_1645,N_1697);
or U1772 (N_1772,N_1629,N_1614);
nor U1773 (N_1773,N_1658,N_1653);
nand U1774 (N_1774,N_1687,N_1648);
nor U1775 (N_1775,N_1693,N_1600);
nor U1776 (N_1776,N_1623,N_1659);
nor U1777 (N_1777,N_1640,N_1626);
or U1778 (N_1778,N_1668,N_1623);
and U1779 (N_1779,N_1615,N_1664);
or U1780 (N_1780,N_1610,N_1669);
nand U1781 (N_1781,N_1627,N_1614);
and U1782 (N_1782,N_1607,N_1622);
and U1783 (N_1783,N_1629,N_1690);
or U1784 (N_1784,N_1640,N_1617);
xnor U1785 (N_1785,N_1630,N_1668);
and U1786 (N_1786,N_1676,N_1653);
nand U1787 (N_1787,N_1684,N_1658);
nor U1788 (N_1788,N_1602,N_1667);
xor U1789 (N_1789,N_1695,N_1622);
and U1790 (N_1790,N_1684,N_1681);
nor U1791 (N_1791,N_1649,N_1662);
xor U1792 (N_1792,N_1666,N_1617);
or U1793 (N_1793,N_1682,N_1668);
nor U1794 (N_1794,N_1666,N_1604);
and U1795 (N_1795,N_1603,N_1605);
and U1796 (N_1796,N_1647,N_1613);
xnor U1797 (N_1797,N_1655,N_1609);
nand U1798 (N_1798,N_1619,N_1614);
and U1799 (N_1799,N_1685,N_1651);
nor U1800 (N_1800,N_1790,N_1776);
nor U1801 (N_1801,N_1727,N_1763);
and U1802 (N_1802,N_1791,N_1712);
or U1803 (N_1803,N_1760,N_1725);
and U1804 (N_1804,N_1782,N_1795);
nor U1805 (N_1805,N_1785,N_1702);
nor U1806 (N_1806,N_1774,N_1718);
nor U1807 (N_1807,N_1743,N_1755);
or U1808 (N_1808,N_1740,N_1711);
nor U1809 (N_1809,N_1749,N_1723);
or U1810 (N_1810,N_1739,N_1713);
and U1811 (N_1811,N_1751,N_1741);
nand U1812 (N_1812,N_1704,N_1714);
xnor U1813 (N_1813,N_1750,N_1731);
nor U1814 (N_1814,N_1788,N_1744);
nand U1815 (N_1815,N_1767,N_1736);
or U1816 (N_1816,N_1730,N_1769);
nor U1817 (N_1817,N_1747,N_1762);
and U1818 (N_1818,N_1779,N_1783);
and U1819 (N_1819,N_1722,N_1734);
or U1820 (N_1820,N_1775,N_1721);
and U1821 (N_1821,N_1761,N_1748);
or U1822 (N_1822,N_1752,N_1710);
nor U1823 (N_1823,N_1746,N_1786);
or U1824 (N_1824,N_1715,N_1784);
xor U1825 (N_1825,N_1781,N_1799);
or U1826 (N_1826,N_1764,N_1737);
or U1827 (N_1827,N_1778,N_1735);
and U1828 (N_1828,N_1794,N_1770);
and U1829 (N_1829,N_1719,N_1745);
nand U1830 (N_1830,N_1773,N_1709);
nand U1831 (N_1831,N_1708,N_1758);
and U1832 (N_1832,N_1759,N_1724);
and U1833 (N_1833,N_1706,N_1797);
or U1834 (N_1834,N_1757,N_1768);
or U1835 (N_1835,N_1789,N_1798);
and U1836 (N_1836,N_1726,N_1753);
nor U1837 (N_1837,N_1796,N_1766);
nor U1838 (N_1838,N_1700,N_1738);
and U1839 (N_1839,N_1716,N_1705);
or U1840 (N_1840,N_1732,N_1754);
or U1841 (N_1841,N_1772,N_1787);
nand U1842 (N_1842,N_1703,N_1701);
or U1843 (N_1843,N_1729,N_1728);
nor U1844 (N_1844,N_1780,N_1720);
nand U1845 (N_1845,N_1707,N_1771);
nand U1846 (N_1846,N_1793,N_1717);
nor U1847 (N_1847,N_1742,N_1765);
xnor U1848 (N_1848,N_1756,N_1792);
xor U1849 (N_1849,N_1733,N_1777);
nand U1850 (N_1850,N_1765,N_1784);
and U1851 (N_1851,N_1767,N_1737);
and U1852 (N_1852,N_1709,N_1775);
or U1853 (N_1853,N_1792,N_1700);
and U1854 (N_1854,N_1777,N_1785);
xor U1855 (N_1855,N_1737,N_1798);
or U1856 (N_1856,N_1738,N_1737);
nand U1857 (N_1857,N_1799,N_1776);
and U1858 (N_1858,N_1703,N_1726);
or U1859 (N_1859,N_1733,N_1711);
nand U1860 (N_1860,N_1728,N_1797);
or U1861 (N_1861,N_1702,N_1717);
and U1862 (N_1862,N_1723,N_1772);
nand U1863 (N_1863,N_1768,N_1797);
nand U1864 (N_1864,N_1719,N_1795);
nor U1865 (N_1865,N_1736,N_1758);
nor U1866 (N_1866,N_1746,N_1794);
nor U1867 (N_1867,N_1784,N_1752);
nor U1868 (N_1868,N_1785,N_1723);
and U1869 (N_1869,N_1723,N_1702);
nor U1870 (N_1870,N_1753,N_1773);
and U1871 (N_1871,N_1758,N_1759);
and U1872 (N_1872,N_1745,N_1723);
or U1873 (N_1873,N_1748,N_1785);
or U1874 (N_1874,N_1767,N_1755);
nand U1875 (N_1875,N_1783,N_1712);
and U1876 (N_1876,N_1768,N_1784);
xor U1877 (N_1877,N_1703,N_1744);
nand U1878 (N_1878,N_1779,N_1729);
or U1879 (N_1879,N_1766,N_1707);
nor U1880 (N_1880,N_1763,N_1794);
nand U1881 (N_1881,N_1724,N_1754);
xor U1882 (N_1882,N_1746,N_1753);
nand U1883 (N_1883,N_1723,N_1779);
nor U1884 (N_1884,N_1723,N_1713);
or U1885 (N_1885,N_1726,N_1730);
nor U1886 (N_1886,N_1729,N_1785);
and U1887 (N_1887,N_1702,N_1798);
xor U1888 (N_1888,N_1776,N_1796);
and U1889 (N_1889,N_1746,N_1721);
nand U1890 (N_1890,N_1710,N_1747);
nor U1891 (N_1891,N_1738,N_1794);
nor U1892 (N_1892,N_1754,N_1751);
or U1893 (N_1893,N_1727,N_1744);
nand U1894 (N_1894,N_1749,N_1778);
nor U1895 (N_1895,N_1717,N_1720);
nand U1896 (N_1896,N_1791,N_1757);
and U1897 (N_1897,N_1780,N_1727);
nand U1898 (N_1898,N_1736,N_1770);
or U1899 (N_1899,N_1797,N_1741);
or U1900 (N_1900,N_1839,N_1838);
nor U1901 (N_1901,N_1814,N_1890);
xor U1902 (N_1902,N_1804,N_1848);
or U1903 (N_1903,N_1822,N_1823);
nand U1904 (N_1904,N_1871,N_1889);
nand U1905 (N_1905,N_1880,N_1835);
and U1906 (N_1906,N_1869,N_1851);
and U1907 (N_1907,N_1808,N_1861);
or U1908 (N_1908,N_1849,N_1827);
xor U1909 (N_1909,N_1874,N_1872);
nor U1910 (N_1910,N_1870,N_1896);
or U1911 (N_1911,N_1858,N_1883);
and U1912 (N_1912,N_1857,N_1886);
and U1913 (N_1913,N_1843,N_1862);
or U1914 (N_1914,N_1878,N_1842);
nor U1915 (N_1915,N_1806,N_1841);
nand U1916 (N_1916,N_1840,N_1859);
and U1917 (N_1917,N_1897,N_1819);
or U1918 (N_1918,N_1832,N_1833);
nand U1919 (N_1919,N_1854,N_1864);
or U1920 (N_1920,N_1898,N_1855);
nor U1921 (N_1921,N_1873,N_1847);
nor U1922 (N_1922,N_1893,N_1875);
nand U1923 (N_1923,N_1879,N_1811);
nand U1924 (N_1924,N_1830,N_1820);
or U1925 (N_1925,N_1846,N_1882);
or U1926 (N_1926,N_1845,N_1885);
or U1927 (N_1927,N_1834,N_1868);
nand U1928 (N_1928,N_1815,N_1828);
and U1929 (N_1929,N_1807,N_1829);
or U1930 (N_1930,N_1899,N_1802);
or U1931 (N_1931,N_1852,N_1853);
nor U1932 (N_1932,N_1831,N_1876);
nor U1933 (N_1933,N_1887,N_1801);
and U1934 (N_1934,N_1837,N_1865);
nand U1935 (N_1935,N_1821,N_1850);
or U1936 (N_1936,N_1884,N_1803);
nand U1937 (N_1937,N_1881,N_1816);
nand U1938 (N_1938,N_1891,N_1856);
and U1939 (N_1939,N_1844,N_1895);
nor U1940 (N_1940,N_1867,N_1894);
nor U1941 (N_1941,N_1825,N_1866);
nor U1942 (N_1942,N_1817,N_1800);
or U1943 (N_1943,N_1805,N_1877);
and U1944 (N_1944,N_1826,N_1824);
and U1945 (N_1945,N_1860,N_1809);
nand U1946 (N_1946,N_1813,N_1888);
nand U1947 (N_1947,N_1812,N_1818);
xor U1948 (N_1948,N_1836,N_1863);
and U1949 (N_1949,N_1892,N_1810);
or U1950 (N_1950,N_1874,N_1806);
nor U1951 (N_1951,N_1899,N_1882);
nand U1952 (N_1952,N_1830,N_1842);
nand U1953 (N_1953,N_1806,N_1833);
or U1954 (N_1954,N_1891,N_1834);
nand U1955 (N_1955,N_1861,N_1892);
nor U1956 (N_1956,N_1830,N_1804);
or U1957 (N_1957,N_1895,N_1824);
and U1958 (N_1958,N_1897,N_1832);
nand U1959 (N_1959,N_1845,N_1824);
or U1960 (N_1960,N_1831,N_1859);
nand U1961 (N_1961,N_1879,N_1858);
nor U1962 (N_1962,N_1854,N_1853);
or U1963 (N_1963,N_1814,N_1882);
nand U1964 (N_1964,N_1851,N_1866);
xnor U1965 (N_1965,N_1898,N_1884);
and U1966 (N_1966,N_1810,N_1877);
and U1967 (N_1967,N_1888,N_1866);
nor U1968 (N_1968,N_1844,N_1840);
and U1969 (N_1969,N_1852,N_1858);
nor U1970 (N_1970,N_1859,N_1874);
and U1971 (N_1971,N_1871,N_1826);
nand U1972 (N_1972,N_1894,N_1870);
or U1973 (N_1973,N_1815,N_1864);
and U1974 (N_1974,N_1872,N_1843);
or U1975 (N_1975,N_1853,N_1875);
nor U1976 (N_1976,N_1867,N_1866);
nor U1977 (N_1977,N_1822,N_1810);
nand U1978 (N_1978,N_1843,N_1855);
or U1979 (N_1979,N_1890,N_1801);
or U1980 (N_1980,N_1874,N_1884);
and U1981 (N_1981,N_1824,N_1836);
and U1982 (N_1982,N_1809,N_1802);
nand U1983 (N_1983,N_1802,N_1892);
nand U1984 (N_1984,N_1835,N_1889);
and U1985 (N_1985,N_1815,N_1839);
and U1986 (N_1986,N_1840,N_1897);
and U1987 (N_1987,N_1823,N_1866);
and U1988 (N_1988,N_1801,N_1862);
nor U1989 (N_1989,N_1802,N_1891);
xnor U1990 (N_1990,N_1832,N_1834);
xnor U1991 (N_1991,N_1846,N_1810);
or U1992 (N_1992,N_1885,N_1867);
nand U1993 (N_1993,N_1889,N_1880);
nor U1994 (N_1994,N_1890,N_1879);
and U1995 (N_1995,N_1806,N_1883);
and U1996 (N_1996,N_1834,N_1876);
nand U1997 (N_1997,N_1880,N_1884);
xor U1998 (N_1998,N_1814,N_1870);
nand U1999 (N_1999,N_1873,N_1885);
xor U2000 (N_2000,N_1914,N_1916);
and U2001 (N_2001,N_1977,N_1997);
or U2002 (N_2002,N_1992,N_1942);
nand U2003 (N_2003,N_1930,N_1989);
nor U2004 (N_2004,N_1981,N_1940);
and U2005 (N_2005,N_1978,N_1976);
nor U2006 (N_2006,N_1934,N_1904);
or U2007 (N_2007,N_1905,N_1929);
and U2008 (N_2008,N_1928,N_1944);
or U2009 (N_2009,N_1946,N_1907);
or U2010 (N_2010,N_1972,N_1964);
nor U2011 (N_2011,N_1911,N_1995);
and U2012 (N_2012,N_1952,N_1955);
xor U2013 (N_2013,N_1988,N_1980);
xnor U2014 (N_2014,N_1950,N_1908);
nand U2015 (N_2015,N_1913,N_1998);
nand U2016 (N_2016,N_1965,N_1951);
nor U2017 (N_2017,N_1948,N_1993);
nor U2018 (N_2018,N_1967,N_1984);
nor U2019 (N_2019,N_1917,N_1939);
nand U2020 (N_2020,N_1927,N_1902);
nand U2021 (N_2021,N_1994,N_1926);
nor U2022 (N_2022,N_1969,N_1931);
nand U2023 (N_2023,N_1910,N_1968);
nand U2024 (N_2024,N_1979,N_1937);
or U2025 (N_2025,N_1971,N_1933);
nor U2026 (N_2026,N_1919,N_1954);
nand U2027 (N_2027,N_1938,N_1959);
xor U2028 (N_2028,N_1903,N_1936);
and U2029 (N_2029,N_1945,N_1963);
and U2030 (N_2030,N_1990,N_1962);
and U2031 (N_2031,N_1923,N_1900);
and U2032 (N_2032,N_1953,N_1921);
xor U2033 (N_2033,N_1915,N_1941);
nand U2034 (N_2034,N_1956,N_1983);
or U2035 (N_2035,N_1912,N_1958);
nor U2036 (N_2036,N_1986,N_1922);
and U2037 (N_2037,N_1949,N_1966);
nor U2038 (N_2038,N_1901,N_1974);
or U2039 (N_2039,N_1991,N_1932);
nor U2040 (N_2040,N_1957,N_1975);
xnor U2041 (N_2041,N_1985,N_1925);
or U2042 (N_2042,N_1996,N_1947);
and U2043 (N_2043,N_1924,N_1906);
or U2044 (N_2044,N_1987,N_1909);
nand U2045 (N_2045,N_1970,N_1982);
or U2046 (N_2046,N_1918,N_1973);
nand U2047 (N_2047,N_1999,N_1943);
or U2048 (N_2048,N_1960,N_1920);
nor U2049 (N_2049,N_1961,N_1935);
and U2050 (N_2050,N_1904,N_1982);
and U2051 (N_2051,N_1931,N_1912);
nand U2052 (N_2052,N_1984,N_1961);
and U2053 (N_2053,N_1995,N_1910);
or U2054 (N_2054,N_1994,N_1928);
or U2055 (N_2055,N_1914,N_1924);
and U2056 (N_2056,N_1976,N_1975);
or U2057 (N_2057,N_1932,N_1935);
and U2058 (N_2058,N_1965,N_1958);
and U2059 (N_2059,N_1942,N_1989);
nand U2060 (N_2060,N_1974,N_1926);
nor U2061 (N_2061,N_1964,N_1990);
or U2062 (N_2062,N_1955,N_1983);
or U2063 (N_2063,N_1956,N_1989);
and U2064 (N_2064,N_1922,N_1931);
or U2065 (N_2065,N_1904,N_1989);
or U2066 (N_2066,N_1952,N_1901);
nand U2067 (N_2067,N_1971,N_1942);
and U2068 (N_2068,N_1953,N_1916);
and U2069 (N_2069,N_1940,N_1944);
nor U2070 (N_2070,N_1918,N_1910);
xnor U2071 (N_2071,N_1905,N_1950);
nand U2072 (N_2072,N_1902,N_1982);
nand U2073 (N_2073,N_1967,N_1937);
or U2074 (N_2074,N_1925,N_1962);
nor U2075 (N_2075,N_1942,N_1961);
and U2076 (N_2076,N_1994,N_1901);
xnor U2077 (N_2077,N_1967,N_1959);
nor U2078 (N_2078,N_1986,N_1923);
nor U2079 (N_2079,N_1948,N_1971);
and U2080 (N_2080,N_1956,N_1980);
nor U2081 (N_2081,N_1909,N_1906);
or U2082 (N_2082,N_1993,N_1919);
or U2083 (N_2083,N_1999,N_1968);
nand U2084 (N_2084,N_1938,N_1971);
and U2085 (N_2085,N_1991,N_1934);
or U2086 (N_2086,N_1965,N_1900);
or U2087 (N_2087,N_1905,N_1979);
nand U2088 (N_2088,N_1946,N_1949);
xnor U2089 (N_2089,N_1985,N_1977);
xnor U2090 (N_2090,N_1955,N_1925);
nand U2091 (N_2091,N_1938,N_1966);
and U2092 (N_2092,N_1996,N_1903);
xor U2093 (N_2093,N_1969,N_1913);
nand U2094 (N_2094,N_1933,N_1967);
and U2095 (N_2095,N_1996,N_1920);
nand U2096 (N_2096,N_1998,N_1939);
or U2097 (N_2097,N_1969,N_1907);
nor U2098 (N_2098,N_1939,N_1980);
and U2099 (N_2099,N_1951,N_1976);
and U2100 (N_2100,N_2080,N_2029);
nor U2101 (N_2101,N_2073,N_2022);
nand U2102 (N_2102,N_2066,N_2062);
nor U2103 (N_2103,N_2079,N_2097);
or U2104 (N_2104,N_2056,N_2060);
or U2105 (N_2105,N_2041,N_2094);
nor U2106 (N_2106,N_2082,N_2092);
and U2107 (N_2107,N_2004,N_2012);
xor U2108 (N_2108,N_2034,N_2040);
or U2109 (N_2109,N_2005,N_2074);
nand U2110 (N_2110,N_2055,N_2000);
and U2111 (N_2111,N_2076,N_2026);
or U2112 (N_2112,N_2027,N_2084);
nor U2113 (N_2113,N_2016,N_2039);
and U2114 (N_2114,N_2028,N_2023);
nor U2115 (N_2115,N_2037,N_2013);
nand U2116 (N_2116,N_2043,N_2024);
or U2117 (N_2117,N_2015,N_2058);
nor U2118 (N_2118,N_2048,N_2045);
nand U2119 (N_2119,N_2051,N_2030);
nand U2120 (N_2120,N_2007,N_2078);
nor U2121 (N_2121,N_2052,N_2087);
xnor U2122 (N_2122,N_2047,N_2008);
nand U2123 (N_2123,N_2020,N_2003);
nand U2124 (N_2124,N_2031,N_2001);
and U2125 (N_2125,N_2032,N_2017);
and U2126 (N_2126,N_2081,N_2014);
nor U2127 (N_2127,N_2083,N_2077);
nand U2128 (N_2128,N_2046,N_2088);
nor U2129 (N_2129,N_2099,N_2002);
or U2130 (N_2130,N_2063,N_2072);
and U2131 (N_2131,N_2068,N_2018);
and U2132 (N_2132,N_2070,N_2069);
or U2133 (N_2133,N_2067,N_2021);
or U2134 (N_2134,N_2093,N_2059);
or U2135 (N_2135,N_2061,N_2090);
nor U2136 (N_2136,N_2095,N_2044);
nor U2137 (N_2137,N_2019,N_2096);
nor U2138 (N_2138,N_2036,N_2085);
or U2139 (N_2139,N_2011,N_2064);
xor U2140 (N_2140,N_2006,N_2009);
and U2141 (N_2141,N_2038,N_2065);
or U2142 (N_2142,N_2089,N_2050);
nor U2143 (N_2143,N_2049,N_2042);
or U2144 (N_2144,N_2053,N_2057);
xnor U2145 (N_2145,N_2054,N_2075);
or U2146 (N_2146,N_2071,N_2091);
and U2147 (N_2147,N_2098,N_2025);
xor U2148 (N_2148,N_2010,N_2033);
xnor U2149 (N_2149,N_2086,N_2035);
nor U2150 (N_2150,N_2041,N_2000);
or U2151 (N_2151,N_2091,N_2060);
nor U2152 (N_2152,N_2070,N_2005);
and U2153 (N_2153,N_2003,N_2072);
nand U2154 (N_2154,N_2093,N_2092);
or U2155 (N_2155,N_2053,N_2083);
nor U2156 (N_2156,N_2064,N_2039);
nor U2157 (N_2157,N_2004,N_2001);
or U2158 (N_2158,N_2092,N_2083);
or U2159 (N_2159,N_2015,N_2092);
or U2160 (N_2160,N_2000,N_2019);
or U2161 (N_2161,N_2022,N_2059);
and U2162 (N_2162,N_2093,N_2025);
or U2163 (N_2163,N_2050,N_2087);
nor U2164 (N_2164,N_2061,N_2068);
xor U2165 (N_2165,N_2094,N_2096);
and U2166 (N_2166,N_2097,N_2013);
and U2167 (N_2167,N_2082,N_2095);
nor U2168 (N_2168,N_2076,N_2049);
or U2169 (N_2169,N_2079,N_2072);
and U2170 (N_2170,N_2057,N_2066);
nor U2171 (N_2171,N_2068,N_2042);
and U2172 (N_2172,N_2058,N_2086);
or U2173 (N_2173,N_2041,N_2079);
nand U2174 (N_2174,N_2042,N_2034);
and U2175 (N_2175,N_2061,N_2048);
and U2176 (N_2176,N_2096,N_2068);
or U2177 (N_2177,N_2032,N_2020);
or U2178 (N_2178,N_2021,N_2047);
nor U2179 (N_2179,N_2068,N_2053);
and U2180 (N_2180,N_2023,N_2031);
nand U2181 (N_2181,N_2061,N_2077);
and U2182 (N_2182,N_2062,N_2025);
or U2183 (N_2183,N_2080,N_2031);
and U2184 (N_2184,N_2027,N_2051);
nand U2185 (N_2185,N_2042,N_2069);
nand U2186 (N_2186,N_2069,N_2004);
or U2187 (N_2187,N_2033,N_2004);
nand U2188 (N_2188,N_2098,N_2040);
and U2189 (N_2189,N_2087,N_2008);
and U2190 (N_2190,N_2012,N_2068);
xnor U2191 (N_2191,N_2022,N_2027);
nor U2192 (N_2192,N_2083,N_2089);
nand U2193 (N_2193,N_2090,N_2042);
nand U2194 (N_2194,N_2057,N_2027);
and U2195 (N_2195,N_2089,N_2028);
nor U2196 (N_2196,N_2069,N_2064);
and U2197 (N_2197,N_2093,N_2068);
and U2198 (N_2198,N_2014,N_2088);
or U2199 (N_2199,N_2040,N_2039);
and U2200 (N_2200,N_2170,N_2187);
and U2201 (N_2201,N_2113,N_2143);
and U2202 (N_2202,N_2118,N_2181);
nand U2203 (N_2203,N_2107,N_2148);
nor U2204 (N_2204,N_2115,N_2108);
or U2205 (N_2205,N_2152,N_2126);
and U2206 (N_2206,N_2199,N_2186);
and U2207 (N_2207,N_2102,N_2153);
or U2208 (N_2208,N_2150,N_2184);
nand U2209 (N_2209,N_2111,N_2198);
nand U2210 (N_2210,N_2182,N_2154);
nand U2211 (N_2211,N_2120,N_2161);
nor U2212 (N_2212,N_2103,N_2142);
nand U2213 (N_2213,N_2159,N_2197);
nand U2214 (N_2214,N_2114,N_2109);
or U2215 (N_2215,N_2151,N_2155);
and U2216 (N_2216,N_2101,N_2172);
nor U2217 (N_2217,N_2123,N_2196);
xnor U2218 (N_2218,N_2136,N_2175);
and U2219 (N_2219,N_2192,N_2166);
nor U2220 (N_2220,N_2173,N_2171);
nor U2221 (N_2221,N_2139,N_2189);
and U2222 (N_2222,N_2156,N_2163);
nand U2223 (N_2223,N_2165,N_2149);
nand U2224 (N_2224,N_2183,N_2168);
and U2225 (N_2225,N_2140,N_2144);
or U2226 (N_2226,N_2169,N_2110);
nor U2227 (N_2227,N_2180,N_2116);
nand U2228 (N_2228,N_2177,N_2147);
nand U2229 (N_2229,N_2145,N_2138);
or U2230 (N_2230,N_2121,N_2117);
or U2231 (N_2231,N_2128,N_2106);
nor U2232 (N_2232,N_2130,N_2133);
and U2233 (N_2233,N_2176,N_2141);
and U2234 (N_2234,N_2137,N_2178);
nor U2235 (N_2235,N_2157,N_2132);
or U2236 (N_2236,N_2190,N_2195);
xor U2237 (N_2237,N_2134,N_2146);
nand U2238 (N_2238,N_2188,N_2191);
or U2239 (N_2239,N_2179,N_2124);
and U2240 (N_2240,N_2112,N_2105);
nand U2241 (N_2241,N_2125,N_2158);
nor U2242 (N_2242,N_2167,N_2162);
or U2243 (N_2243,N_2174,N_2185);
or U2244 (N_2244,N_2160,N_2131);
nor U2245 (N_2245,N_2104,N_2127);
and U2246 (N_2246,N_2100,N_2135);
nor U2247 (N_2247,N_2194,N_2129);
nor U2248 (N_2248,N_2193,N_2119);
or U2249 (N_2249,N_2122,N_2164);
or U2250 (N_2250,N_2148,N_2134);
nand U2251 (N_2251,N_2164,N_2165);
or U2252 (N_2252,N_2165,N_2124);
nor U2253 (N_2253,N_2102,N_2148);
xor U2254 (N_2254,N_2191,N_2101);
nor U2255 (N_2255,N_2178,N_2195);
and U2256 (N_2256,N_2127,N_2173);
or U2257 (N_2257,N_2157,N_2117);
or U2258 (N_2258,N_2190,N_2187);
or U2259 (N_2259,N_2129,N_2196);
or U2260 (N_2260,N_2154,N_2138);
nor U2261 (N_2261,N_2188,N_2132);
or U2262 (N_2262,N_2179,N_2150);
and U2263 (N_2263,N_2143,N_2157);
and U2264 (N_2264,N_2165,N_2194);
and U2265 (N_2265,N_2179,N_2186);
and U2266 (N_2266,N_2175,N_2158);
nor U2267 (N_2267,N_2130,N_2194);
or U2268 (N_2268,N_2120,N_2159);
or U2269 (N_2269,N_2145,N_2198);
nand U2270 (N_2270,N_2111,N_2169);
xnor U2271 (N_2271,N_2153,N_2124);
or U2272 (N_2272,N_2141,N_2130);
nand U2273 (N_2273,N_2110,N_2144);
and U2274 (N_2274,N_2112,N_2180);
or U2275 (N_2275,N_2188,N_2186);
nor U2276 (N_2276,N_2163,N_2143);
or U2277 (N_2277,N_2196,N_2118);
and U2278 (N_2278,N_2139,N_2137);
nor U2279 (N_2279,N_2135,N_2195);
or U2280 (N_2280,N_2145,N_2184);
or U2281 (N_2281,N_2175,N_2122);
nor U2282 (N_2282,N_2197,N_2166);
and U2283 (N_2283,N_2101,N_2147);
or U2284 (N_2284,N_2129,N_2171);
or U2285 (N_2285,N_2184,N_2163);
xor U2286 (N_2286,N_2106,N_2158);
or U2287 (N_2287,N_2127,N_2181);
and U2288 (N_2288,N_2192,N_2179);
or U2289 (N_2289,N_2138,N_2115);
nor U2290 (N_2290,N_2119,N_2165);
or U2291 (N_2291,N_2166,N_2151);
or U2292 (N_2292,N_2111,N_2157);
xor U2293 (N_2293,N_2141,N_2112);
or U2294 (N_2294,N_2165,N_2190);
nand U2295 (N_2295,N_2136,N_2149);
or U2296 (N_2296,N_2169,N_2166);
or U2297 (N_2297,N_2119,N_2167);
or U2298 (N_2298,N_2167,N_2143);
and U2299 (N_2299,N_2147,N_2143);
nor U2300 (N_2300,N_2249,N_2238);
xor U2301 (N_2301,N_2293,N_2252);
and U2302 (N_2302,N_2218,N_2245);
nor U2303 (N_2303,N_2210,N_2279);
nor U2304 (N_2304,N_2211,N_2267);
nand U2305 (N_2305,N_2294,N_2261);
nand U2306 (N_2306,N_2213,N_2228);
nand U2307 (N_2307,N_2223,N_2271);
and U2308 (N_2308,N_2226,N_2215);
and U2309 (N_2309,N_2285,N_2202);
or U2310 (N_2310,N_2295,N_2203);
and U2311 (N_2311,N_2236,N_2286);
or U2312 (N_2312,N_2263,N_2254);
nand U2313 (N_2313,N_2241,N_2214);
or U2314 (N_2314,N_2222,N_2250);
nor U2315 (N_2315,N_2278,N_2287);
nor U2316 (N_2316,N_2207,N_2298);
xor U2317 (N_2317,N_2262,N_2259);
and U2318 (N_2318,N_2231,N_2232);
and U2319 (N_2319,N_2219,N_2297);
nor U2320 (N_2320,N_2208,N_2273);
nor U2321 (N_2321,N_2264,N_2237);
or U2322 (N_2322,N_2200,N_2276);
or U2323 (N_2323,N_2227,N_2216);
nand U2324 (N_2324,N_2205,N_2234);
nand U2325 (N_2325,N_2248,N_2290);
or U2326 (N_2326,N_2220,N_2201);
nor U2327 (N_2327,N_2266,N_2224);
nor U2328 (N_2328,N_2281,N_2235);
nand U2329 (N_2329,N_2225,N_2246);
nor U2330 (N_2330,N_2277,N_2289);
nor U2331 (N_2331,N_2265,N_2291);
nor U2332 (N_2332,N_2258,N_2288);
nor U2333 (N_2333,N_2256,N_2251);
nand U2334 (N_2334,N_2270,N_2268);
nand U2335 (N_2335,N_2255,N_2269);
nor U2336 (N_2336,N_2260,N_2209);
nor U2337 (N_2337,N_2257,N_2239);
nor U2338 (N_2338,N_2283,N_2274);
nor U2339 (N_2339,N_2275,N_2253);
nand U2340 (N_2340,N_2244,N_2292);
and U2341 (N_2341,N_2206,N_2229);
nand U2342 (N_2342,N_2272,N_2282);
nand U2343 (N_2343,N_2296,N_2233);
nand U2344 (N_2344,N_2230,N_2280);
and U2345 (N_2345,N_2212,N_2299);
or U2346 (N_2346,N_2204,N_2242);
or U2347 (N_2347,N_2284,N_2221);
nor U2348 (N_2348,N_2240,N_2243);
nand U2349 (N_2349,N_2217,N_2247);
and U2350 (N_2350,N_2260,N_2219);
xnor U2351 (N_2351,N_2274,N_2252);
and U2352 (N_2352,N_2268,N_2216);
nor U2353 (N_2353,N_2206,N_2261);
nand U2354 (N_2354,N_2234,N_2247);
nor U2355 (N_2355,N_2291,N_2242);
and U2356 (N_2356,N_2220,N_2203);
or U2357 (N_2357,N_2228,N_2236);
and U2358 (N_2358,N_2253,N_2212);
and U2359 (N_2359,N_2213,N_2259);
nor U2360 (N_2360,N_2234,N_2291);
or U2361 (N_2361,N_2297,N_2222);
nand U2362 (N_2362,N_2263,N_2216);
nand U2363 (N_2363,N_2259,N_2205);
xor U2364 (N_2364,N_2290,N_2259);
nand U2365 (N_2365,N_2269,N_2253);
or U2366 (N_2366,N_2290,N_2227);
nor U2367 (N_2367,N_2216,N_2289);
xnor U2368 (N_2368,N_2229,N_2247);
nor U2369 (N_2369,N_2201,N_2245);
xnor U2370 (N_2370,N_2215,N_2265);
nor U2371 (N_2371,N_2260,N_2201);
nand U2372 (N_2372,N_2238,N_2223);
nor U2373 (N_2373,N_2213,N_2212);
nand U2374 (N_2374,N_2288,N_2299);
xnor U2375 (N_2375,N_2289,N_2295);
nor U2376 (N_2376,N_2226,N_2270);
nor U2377 (N_2377,N_2211,N_2260);
nor U2378 (N_2378,N_2257,N_2279);
or U2379 (N_2379,N_2258,N_2299);
xor U2380 (N_2380,N_2267,N_2279);
and U2381 (N_2381,N_2243,N_2234);
and U2382 (N_2382,N_2269,N_2260);
and U2383 (N_2383,N_2271,N_2250);
and U2384 (N_2384,N_2294,N_2258);
and U2385 (N_2385,N_2297,N_2262);
or U2386 (N_2386,N_2293,N_2262);
or U2387 (N_2387,N_2267,N_2209);
nand U2388 (N_2388,N_2253,N_2274);
nor U2389 (N_2389,N_2226,N_2246);
nand U2390 (N_2390,N_2241,N_2227);
or U2391 (N_2391,N_2262,N_2215);
nor U2392 (N_2392,N_2267,N_2252);
xor U2393 (N_2393,N_2205,N_2256);
xor U2394 (N_2394,N_2261,N_2280);
nand U2395 (N_2395,N_2277,N_2290);
xnor U2396 (N_2396,N_2259,N_2266);
or U2397 (N_2397,N_2279,N_2240);
xnor U2398 (N_2398,N_2288,N_2247);
nor U2399 (N_2399,N_2232,N_2221);
nor U2400 (N_2400,N_2358,N_2354);
and U2401 (N_2401,N_2375,N_2304);
nand U2402 (N_2402,N_2379,N_2352);
and U2403 (N_2403,N_2362,N_2320);
xnor U2404 (N_2404,N_2373,N_2335);
nand U2405 (N_2405,N_2328,N_2366);
and U2406 (N_2406,N_2302,N_2343);
or U2407 (N_2407,N_2365,N_2307);
nand U2408 (N_2408,N_2309,N_2312);
and U2409 (N_2409,N_2369,N_2303);
nand U2410 (N_2410,N_2367,N_2300);
or U2411 (N_2411,N_2322,N_2334);
nand U2412 (N_2412,N_2317,N_2372);
nand U2413 (N_2413,N_2361,N_2377);
nor U2414 (N_2414,N_2319,N_2313);
nand U2415 (N_2415,N_2323,N_2348);
and U2416 (N_2416,N_2314,N_2316);
or U2417 (N_2417,N_2376,N_2364);
nand U2418 (N_2418,N_2336,N_2349);
or U2419 (N_2419,N_2332,N_2310);
nor U2420 (N_2420,N_2350,N_2340);
or U2421 (N_2421,N_2357,N_2396);
or U2422 (N_2422,N_2351,N_2345);
or U2423 (N_2423,N_2383,N_2381);
or U2424 (N_2424,N_2398,N_2391);
nor U2425 (N_2425,N_2399,N_2392);
or U2426 (N_2426,N_2387,N_2311);
nor U2427 (N_2427,N_2327,N_2305);
and U2428 (N_2428,N_2363,N_2356);
nand U2429 (N_2429,N_2378,N_2318);
nor U2430 (N_2430,N_2338,N_2339);
xnor U2431 (N_2431,N_2359,N_2388);
or U2432 (N_2432,N_2389,N_2337);
nand U2433 (N_2433,N_2397,N_2385);
and U2434 (N_2434,N_2380,N_2394);
or U2435 (N_2435,N_2329,N_2321);
nand U2436 (N_2436,N_2330,N_2342);
or U2437 (N_2437,N_2306,N_2347);
nand U2438 (N_2438,N_2333,N_2390);
and U2439 (N_2439,N_2301,N_2315);
nor U2440 (N_2440,N_2360,N_2371);
and U2441 (N_2441,N_2395,N_2384);
xnor U2442 (N_2442,N_2374,N_2386);
or U2443 (N_2443,N_2326,N_2382);
nand U2444 (N_2444,N_2393,N_2344);
or U2445 (N_2445,N_2324,N_2331);
or U2446 (N_2446,N_2353,N_2355);
nand U2447 (N_2447,N_2370,N_2368);
nand U2448 (N_2448,N_2325,N_2308);
nand U2449 (N_2449,N_2341,N_2346);
xor U2450 (N_2450,N_2388,N_2328);
and U2451 (N_2451,N_2304,N_2394);
and U2452 (N_2452,N_2383,N_2311);
nand U2453 (N_2453,N_2307,N_2392);
and U2454 (N_2454,N_2396,N_2314);
nand U2455 (N_2455,N_2394,N_2329);
nand U2456 (N_2456,N_2348,N_2301);
or U2457 (N_2457,N_2369,N_2389);
nand U2458 (N_2458,N_2318,N_2338);
or U2459 (N_2459,N_2351,N_2376);
nand U2460 (N_2460,N_2318,N_2313);
nor U2461 (N_2461,N_2376,N_2383);
or U2462 (N_2462,N_2381,N_2347);
or U2463 (N_2463,N_2327,N_2315);
nor U2464 (N_2464,N_2309,N_2391);
nor U2465 (N_2465,N_2382,N_2330);
nand U2466 (N_2466,N_2346,N_2325);
nand U2467 (N_2467,N_2395,N_2349);
nand U2468 (N_2468,N_2393,N_2312);
and U2469 (N_2469,N_2350,N_2308);
or U2470 (N_2470,N_2387,N_2399);
or U2471 (N_2471,N_2381,N_2358);
or U2472 (N_2472,N_2306,N_2357);
and U2473 (N_2473,N_2396,N_2375);
or U2474 (N_2474,N_2324,N_2359);
nor U2475 (N_2475,N_2394,N_2347);
xor U2476 (N_2476,N_2318,N_2306);
xnor U2477 (N_2477,N_2389,N_2386);
nor U2478 (N_2478,N_2376,N_2357);
nand U2479 (N_2479,N_2330,N_2367);
and U2480 (N_2480,N_2338,N_2343);
nand U2481 (N_2481,N_2347,N_2396);
or U2482 (N_2482,N_2387,N_2359);
nand U2483 (N_2483,N_2381,N_2307);
nand U2484 (N_2484,N_2379,N_2341);
nor U2485 (N_2485,N_2322,N_2375);
and U2486 (N_2486,N_2342,N_2334);
nand U2487 (N_2487,N_2366,N_2369);
and U2488 (N_2488,N_2344,N_2322);
nand U2489 (N_2489,N_2310,N_2319);
or U2490 (N_2490,N_2321,N_2353);
nor U2491 (N_2491,N_2316,N_2342);
nand U2492 (N_2492,N_2367,N_2312);
and U2493 (N_2493,N_2301,N_2321);
nand U2494 (N_2494,N_2374,N_2335);
nand U2495 (N_2495,N_2391,N_2311);
nand U2496 (N_2496,N_2337,N_2324);
xnor U2497 (N_2497,N_2319,N_2387);
and U2498 (N_2498,N_2339,N_2375);
nor U2499 (N_2499,N_2354,N_2387);
nor U2500 (N_2500,N_2452,N_2493);
or U2501 (N_2501,N_2469,N_2456);
nand U2502 (N_2502,N_2450,N_2411);
nor U2503 (N_2503,N_2461,N_2409);
and U2504 (N_2504,N_2470,N_2481);
or U2505 (N_2505,N_2441,N_2467);
nor U2506 (N_2506,N_2476,N_2492);
nand U2507 (N_2507,N_2463,N_2413);
nand U2508 (N_2508,N_2430,N_2436);
or U2509 (N_2509,N_2419,N_2466);
or U2510 (N_2510,N_2485,N_2446);
and U2511 (N_2511,N_2400,N_2480);
and U2512 (N_2512,N_2421,N_2483);
or U2513 (N_2513,N_2479,N_2489);
nor U2514 (N_2514,N_2438,N_2462);
and U2515 (N_2515,N_2401,N_2488);
nor U2516 (N_2516,N_2459,N_2435);
xnor U2517 (N_2517,N_2460,N_2408);
or U2518 (N_2518,N_2407,N_2468);
or U2519 (N_2519,N_2418,N_2457);
or U2520 (N_2520,N_2471,N_2453);
nand U2521 (N_2521,N_2499,N_2443);
or U2522 (N_2522,N_2403,N_2472);
nor U2523 (N_2523,N_2412,N_2474);
nor U2524 (N_2524,N_2454,N_2426);
nand U2525 (N_2525,N_2473,N_2402);
nand U2526 (N_2526,N_2496,N_2424);
and U2527 (N_2527,N_2458,N_2464);
nand U2528 (N_2528,N_2410,N_2451);
and U2529 (N_2529,N_2455,N_2484);
nand U2530 (N_2530,N_2439,N_2429);
or U2531 (N_2531,N_2417,N_2448);
nor U2532 (N_2532,N_2465,N_2434);
nor U2533 (N_2533,N_2494,N_2420);
nand U2534 (N_2534,N_2475,N_2445);
or U2535 (N_2535,N_2437,N_2449);
nor U2536 (N_2536,N_2490,N_2487);
nor U2537 (N_2537,N_2497,N_2422);
or U2538 (N_2538,N_2444,N_2406);
xnor U2539 (N_2539,N_2423,N_2404);
xor U2540 (N_2540,N_2405,N_2440);
nor U2541 (N_2541,N_2415,N_2414);
xor U2542 (N_2542,N_2447,N_2432);
or U2543 (N_2543,N_2477,N_2431);
or U2544 (N_2544,N_2495,N_2433);
or U2545 (N_2545,N_2425,N_2491);
nor U2546 (N_2546,N_2486,N_2428);
nand U2547 (N_2547,N_2427,N_2478);
nor U2548 (N_2548,N_2442,N_2416);
nor U2549 (N_2549,N_2482,N_2498);
and U2550 (N_2550,N_2421,N_2439);
nand U2551 (N_2551,N_2484,N_2416);
and U2552 (N_2552,N_2411,N_2496);
and U2553 (N_2553,N_2484,N_2466);
nor U2554 (N_2554,N_2445,N_2450);
or U2555 (N_2555,N_2490,N_2438);
nor U2556 (N_2556,N_2442,N_2410);
or U2557 (N_2557,N_2489,N_2439);
and U2558 (N_2558,N_2474,N_2499);
and U2559 (N_2559,N_2450,N_2404);
xnor U2560 (N_2560,N_2467,N_2480);
nor U2561 (N_2561,N_2429,N_2418);
nor U2562 (N_2562,N_2490,N_2456);
and U2563 (N_2563,N_2415,N_2436);
nor U2564 (N_2564,N_2456,N_2479);
or U2565 (N_2565,N_2445,N_2433);
nor U2566 (N_2566,N_2460,N_2481);
nor U2567 (N_2567,N_2424,N_2452);
and U2568 (N_2568,N_2417,N_2423);
nor U2569 (N_2569,N_2411,N_2462);
or U2570 (N_2570,N_2411,N_2423);
and U2571 (N_2571,N_2414,N_2419);
nand U2572 (N_2572,N_2445,N_2481);
and U2573 (N_2573,N_2437,N_2482);
nand U2574 (N_2574,N_2489,N_2413);
and U2575 (N_2575,N_2418,N_2480);
nor U2576 (N_2576,N_2441,N_2490);
nand U2577 (N_2577,N_2413,N_2470);
nand U2578 (N_2578,N_2486,N_2457);
nor U2579 (N_2579,N_2466,N_2469);
or U2580 (N_2580,N_2450,N_2419);
nor U2581 (N_2581,N_2419,N_2475);
or U2582 (N_2582,N_2443,N_2435);
and U2583 (N_2583,N_2448,N_2426);
nand U2584 (N_2584,N_2460,N_2443);
and U2585 (N_2585,N_2499,N_2495);
or U2586 (N_2586,N_2446,N_2497);
and U2587 (N_2587,N_2498,N_2489);
and U2588 (N_2588,N_2400,N_2463);
and U2589 (N_2589,N_2480,N_2416);
nor U2590 (N_2590,N_2474,N_2443);
or U2591 (N_2591,N_2434,N_2453);
and U2592 (N_2592,N_2497,N_2489);
and U2593 (N_2593,N_2427,N_2482);
nand U2594 (N_2594,N_2498,N_2425);
and U2595 (N_2595,N_2470,N_2472);
nor U2596 (N_2596,N_2450,N_2479);
or U2597 (N_2597,N_2482,N_2477);
nand U2598 (N_2598,N_2460,N_2476);
nor U2599 (N_2599,N_2450,N_2455);
and U2600 (N_2600,N_2530,N_2511);
and U2601 (N_2601,N_2563,N_2583);
or U2602 (N_2602,N_2546,N_2596);
and U2603 (N_2603,N_2588,N_2595);
and U2604 (N_2604,N_2533,N_2585);
and U2605 (N_2605,N_2575,N_2535);
nand U2606 (N_2606,N_2528,N_2509);
nor U2607 (N_2607,N_2568,N_2569);
nand U2608 (N_2608,N_2566,N_2547);
and U2609 (N_2609,N_2518,N_2549);
nand U2610 (N_2610,N_2508,N_2539);
or U2611 (N_2611,N_2523,N_2597);
or U2612 (N_2612,N_2561,N_2504);
or U2613 (N_2613,N_2579,N_2513);
and U2614 (N_2614,N_2590,N_2537);
nor U2615 (N_2615,N_2525,N_2556);
and U2616 (N_2616,N_2515,N_2536);
and U2617 (N_2617,N_2514,N_2529);
nor U2618 (N_2618,N_2532,N_2582);
nand U2619 (N_2619,N_2543,N_2548);
nor U2620 (N_2620,N_2545,N_2519);
and U2621 (N_2621,N_2516,N_2540);
and U2622 (N_2622,N_2551,N_2506);
or U2623 (N_2623,N_2565,N_2507);
or U2624 (N_2624,N_2571,N_2538);
nor U2625 (N_2625,N_2584,N_2574);
or U2626 (N_2626,N_2503,N_2557);
or U2627 (N_2627,N_2589,N_2593);
xor U2628 (N_2628,N_2573,N_2520);
or U2629 (N_2629,N_2510,N_2581);
or U2630 (N_2630,N_2587,N_2558);
nand U2631 (N_2631,N_2592,N_2591);
nand U2632 (N_2632,N_2526,N_2521);
or U2633 (N_2633,N_2531,N_2550);
nand U2634 (N_2634,N_2580,N_2599);
or U2635 (N_2635,N_2554,N_2560);
nand U2636 (N_2636,N_2522,N_2517);
xor U2637 (N_2637,N_2505,N_2577);
or U2638 (N_2638,N_2544,N_2562);
nand U2639 (N_2639,N_2500,N_2570);
and U2640 (N_2640,N_2524,N_2576);
or U2641 (N_2641,N_2501,N_2512);
nand U2642 (N_2642,N_2564,N_2559);
or U2643 (N_2643,N_2572,N_2534);
xor U2644 (N_2644,N_2555,N_2567);
nor U2645 (N_2645,N_2594,N_2541);
and U2646 (N_2646,N_2586,N_2502);
nand U2647 (N_2647,N_2578,N_2553);
or U2648 (N_2648,N_2598,N_2552);
and U2649 (N_2649,N_2542,N_2527);
or U2650 (N_2650,N_2544,N_2580);
or U2651 (N_2651,N_2594,N_2519);
or U2652 (N_2652,N_2508,N_2574);
and U2653 (N_2653,N_2542,N_2537);
and U2654 (N_2654,N_2528,N_2571);
or U2655 (N_2655,N_2593,N_2592);
xnor U2656 (N_2656,N_2507,N_2562);
nand U2657 (N_2657,N_2514,N_2534);
nor U2658 (N_2658,N_2566,N_2505);
xor U2659 (N_2659,N_2586,N_2565);
xor U2660 (N_2660,N_2535,N_2552);
and U2661 (N_2661,N_2543,N_2581);
nor U2662 (N_2662,N_2513,N_2537);
xnor U2663 (N_2663,N_2521,N_2518);
nor U2664 (N_2664,N_2531,N_2590);
xor U2665 (N_2665,N_2505,N_2591);
or U2666 (N_2666,N_2589,N_2517);
or U2667 (N_2667,N_2527,N_2599);
and U2668 (N_2668,N_2546,N_2584);
nor U2669 (N_2669,N_2596,N_2507);
xor U2670 (N_2670,N_2517,N_2596);
nand U2671 (N_2671,N_2548,N_2572);
and U2672 (N_2672,N_2508,N_2533);
and U2673 (N_2673,N_2559,N_2583);
nand U2674 (N_2674,N_2570,N_2514);
nor U2675 (N_2675,N_2507,N_2543);
nor U2676 (N_2676,N_2523,N_2598);
xnor U2677 (N_2677,N_2515,N_2537);
and U2678 (N_2678,N_2515,N_2594);
nor U2679 (N_2679,N_2586,N_2594);
xnor U2680 (N_2680,N_2551,N_2514);
and U2681 (N_2681,N_2500,N_2540);
nor U2682 (N_2682,N_2579,N_2524);
or U2683 (N_2683,N_2547,N_2594);
nand U2684 (N_2684,N_2551,N_2597);
and U2685 (N_2685,N_2503,N_2588);
or U2686 (N_2686,N_2597,N_2576);
and U2687 (N_2687,N_2514,N_2515);
or U2688 (N_2688,N_2556,N_2517);
and U2689 (N_2689,N_2524,N_2585);
and U2690 (N_2690,N_2504,N_2565);
and U2691 (N_2691,N_2531,N_2528);
nor U2692 (N_2692,N_2538,N_2542);
nor U2693 (N_2693,N_2597,N_2574);
nand U2694 (N_2694,N_2560,N_2584);
xor U2695 (N_2695,N_2548,N_2535);
nor U2696 (N_2696,N_2543,N_2582);
or U2697 (N_2697,N_2591,N_2523);
and U2698 (N_2698,N_2512,N_2585);
nor U2699 (N_2699,N_2559,N_2549);
nand U2700 (N_2700,N_2673,N_2682);
or U2701 (N_2701,N_2634,N_2609);
nor U2702 (N_2702,N_2671,N_2657);
nor U2703 (N_2703,N_2604,N_2645);
and U2704 (N_2704,N_2662,N_2667);
or U2705 (N_2705,N_2636,N_2615);
nand U2706 (N_2706,N_2659,N_2686);
or U2707 (N_2707,N_2695,N_2640);
or U2708 (N_2708,N_2621,N_2696);
nand U2709 (N_2709,N_2653,N_2674);
and U2710 (N_2710,N_2633,N_2649);
or U2711 (N_2711,N_2614,N_2610);
or U2712 (N_2712,N_2687,N_2663);
and U2713 (N_2713,N_2675,N_2679);
and U2714 (N_2714,N_2643,N_2669);
xnor U2715 (N_2715,N_2651,N_2654);
xor U2716 (N_2716,N_2692,N_2638);
xor U2717 (N_2717,N_2631,N_2690);
nand U2718 (N_2718,N_2611,N_2664);
xor U2719 (N_2719,N_2666,N_2616);
and U2720 (N_2720,N_2655,N_2660);
nor U2721 (N_2721,N_2607,N_2697);
and U2722 (N_2722,N_2642,N_2632);
or U2723 (N_2723,N_2661,N_2647);
nand U2724 (N_2724,N_2698,N_2684);
nand U2725 (N_2725,N_2693,N_2691);
xnor U2726 (N_2726,N_2681,N_2622);
and U2727 (N_2727,N_2678,N_2618);
nor U2728 (N_2728,N_2656,N_2683);
or U2729 (N_2729,N_2648,N_2601);
nand U2730 (N_2730,N_2652,N_2677);
nor U2731 (N_2731,N_2699,N_2685);
or U2732 (N_2732,N_2646,N_2624);
nand U2733 (N_2733,N_2680,N_2619);
and U2734 (N_2734,N_2694,N_2635);
nor U2735 (N_2735,N_2600,N_2670);
nor U2736 (N_2736,N_2688,N_2620);
xor U2737 (N_2737,N_2627,N_2603);
nand U2738 (N_2738,N_2676,N_2606);
nor U2739 (N_2739,N_2625,N_2602);
nor U2740 (N_2740,N_2639,N_2665);
or U2741 (N_2741,N_2617,N_2644);
and U2742 (N_2742,N_2668,N_2637);
nand U2743 (N_2743,N_2672,N_2629);
nor U2744 (N_2744,N_2630,N_2650);
and U2745 (N_2745,N_2641,N_2628);
nor U2746 (N_2746,N_2608,N_2689);
or U2747 (N_2747,N_2612,N_2613);
nand U2748 (N_2748,N_2623,N_2626);
or U2749 (N_2749,N_2605,N_2658);
nor U2750 (N_2750,N_2606,N_2616);
nor U2751 (N_2751,N_2601,N_2600);
nand U2752 (N_2752,N_2690,N_2608);
xor U2753 (N_2753,N_2697,N_2666);
nor U2754 (N_2754,N_2699,N_2693);
or U2755 (N_2755,N_2623,N_2614);
and U2756 (N_2756,N_2689,N_2601);
or U2757 (N_2757,N_2666,N_2603);
and U2758 (N_2758,N_2613,N_2631);
and U2759 (N_2759,N_2663,N_2611);
nor U2760 (N_2760,N_2644,N_2606);
nand U2761 (N_2761,N_2699,N_2674);
and U2762 (N_2762,N_2605,N_2664);
nand U2763 (N_2763,N_2682,N_2605);
nand U2764 (N_2764,N_2694,N_2633);
nand U2765 (N_2765,N_2672,N_2694);
or U2766 (N_2766,N_2602,N_2612);
xnor U2767 (N_2767,N_2619,N_2641);
nor U2768 (N_2768,N_2688,N_2661);
nor U2769 (N_2769,N_2612,N_2631);
nor U2770 (N_2770,N_2687,N_2692);
or U2771 (N_2771,N_2608,N_2654);
or U2772 (N_2772,N_2691,N_2651);
and U2773 (N_2773,N_2692,N_2696);
nand U2774 (N_2774,N_2636,N_2673);
and U2775 (N_2775,N_2616,N_2621);
nor U2776 (N_2776,N_2680,N_2661);
and U2777 (N_2777,N_2695,N_2633);
xnor U2778 (N_2778,N_2664,N_2699);
and U2779 (N_2779,N_2641,N_2697);
nor U2780 (N_2780,N_2685,N_2659);
or U2781 (N_2781,N_2655,N_2642);
or U2782 (N_2782,N_2656,N_2689);
nand U2783 (N_2783,N_2603,N_2648);
or U2784 (N_2784,N_2698,N_2609);
xnor U2785 (N_2785,N_2620,N_2647);
nor U2786 (N_2786,N_2633,N_2670);
or U2787 (N_2787,N_2631,N_2663);
xnor U2788 (N_2788,N_2673,N_2612);
or U2789 (N_2789,N_2650,N_2672);
or U2790 (N_2790,N_2600,N_2672);
or U2791 (N_2791,N_2667,N_2624);
nor U2792 (N_2792,N_2615,N_2627);
or U2793 (N_2793,N_2637,N_2619);
and U2794 (N_2794,N_2646,N_2691);
xnor U2795 (N_2795,N_2637,N_2692);
or U2796 (N_2796,N_2697,N_2606);
or U2797 (N_2797,N_2603,N_2642);
nand U2798 (N_2798,N_2629,N_2692);
xor U2799 (N_2799,N_2606,N_2660);
nand U2800 (N_2800,N_2700,N_2752);
nand U2801 (N_2801,N_2736,N_2762);
or U2802 (N_2802,N_2714,N_2777);
nand U2803 (N_2803,N_2749,N_2760);
nand U2804 (N_2804,N_2742,N_2781);
or U2805 (N_2805,N_2765,N_2791);
or U2806 (N_2806,N_2730,N_2710);
nor U2807 (N_2807,N_2764,N_2773);
nand U2808 (N_2808,N_2741,N_2704);
nor U2809 (N_2809,N_2732,N_2794);
and U2810 (N_2810,N_2726,N_2783);
nor U2811 (N_2811,N_2718,N_2711);
nand U2812 (N_2812,N_2797,N_2793);
or U2813 (N_2813,N_2795,N_2701);
or U2814 (N_2814,N_2724,N_2747);
nor U2815 (N_2815,N_2739,N_2798);
nand U2816 (N_2816,N_2757,N_2750);
nand U2817 (N_2817,N_2720,N_2766);
nand U2818 (N_2818,N_2778,N_2790);
nor U2819 (N_2819,N_2788,N_2789);
nor U2820 (N_2820,N_2768,N_2774);
nor U2821 (N_2821,N_2782,N_2708);
or U2822 (N_2822,N_2713,N_2709);
xor U2823 (N_2823,N_2779,N_2784);
nor U2824 (N_2824,N_2716,N_2758);
and U2825 (N_2825,N_2706,N_2743);
nand U2826 (N_2826,N_2763,N_2703);
nand U2827 (N_2827,N_2796,N_2731);
and U2828 (N_2828,N_2722,N_2717);
xnor U2829 (N_2829,N_2767,N_2744);
nand U2830 (N_2830,N_2707,N_2771);
nand U2831 (N_2831,N_2754,N_2729);
nand U2832 (N_2832,N_2775,N_2740);
or U2833 (N_2833,N_2748,N_2737);
nor U2834 (N_2834,N_2770,N_2792);
nor U2835 (N_2835,N_2745,N_2776);
nand U2836 (N_2836,N_2787,N_2738);
or U2837 (N_2837,N_2780,N_2723);
nand U2838 (N_2838,N_2719,N_2761);
nand U2839 (N_2839,N_2734,N_2725);
nand U2840 (N_2840,N_2733,N_2753);
and U2841 (N_2841,N_2772,N_2702);
or U2842 (N_2842,N_2756,N_2705);
or U2843 (N_2843,N_2746,N_2712);
or U2844 (N_2844,N_2735,N_2715);
and U2845 (N_2845,N_2786,N_2785);
nand U2846 (N_2846,N_2759,N_2755);
and U2847 (N_2847,N_2721,N_2728);
and U2848 (N_2848,N_2799,N_2727);
nand U2849 (N_2849,N_2751,N_2769);
nor U2850 (N_2850,N_2794,N_2703);
nand U2851 (N_2851,N_2707,N_2746);
nor U2852 (N_2852,N_2792,N_2730);
or U2853 (N_2853,N_2727,N_2706);
and U2854 (N_2854,N_2721,N_2755);
nand U2855 (N_2855,N_2766,N_2761);
nand U2856 (N_2856,N_2776,N_2734);
nor U2857 (N_2857,N_2762,N_2700);
or U2858 (N_2858,N_2746,N_2711);
nor U2859 (N_2859,N_2794,N_2734);
nor U2860 (N_2860,N_2797,N_2752);
and U2861 (N_2861,N_2727,N_2772);
xnor U2862 (N_2862,N_2731,N_2706);
nand U2863 (N_2863,N_2786,N_2737);
nor U2864 (N_2864,N_2725,N_2791);
xor U2865 (N_2865,N_2792,N_2715);
nand U2866 (N_2866,N_2706,N_2772);
and U2867 (N_2867,N_2797,N_2701);
or U2868 (N_2868,N_2700,N_2721);
or U2869 (N_2869,N_2752,N_2788);
or U2870 (N_2870,N_2799,N_2733);
and U2871 (N_2871,N_2787,N_2756);
nand U2872 (N_2872,N_2730,N_2739);
and U2873 (N_2873,N_2736,N_2787);
or U2874 (N_2874,N_2797,N_2765);
nor U2875 (N_2875,N_2734,N_2732);
and U2876 (N_2876,N_2759,N_2773);
nand U2877 (N_2877,N_2765,N_2726);
or U2878 (N_2878,N_2733,N_2718);
xnor U2879 (N_2879,N_2753,N_2759);
nand U2880 (N_2880,N_2728,N_2741);
nor U2881 (N_2881,N_2787,N_2792);
or U2882 (N_2882,N_2796,N_2749);
nor U2883 (N_2883,N_2794,N_2756);
nor U2884 (N_2884,N_2710,N_2787);
xor U2885 (N_2885,N_2712,N_2701);
or U2886 (N_2886,N_2711,N_2753);
and U2887 (N_2887,N_2729,N_2705);
nand U2888 (N_2888,N_2714,N_2770);
and U2889 (N_2889,N_2715,N_2703);
and U2890 (N_2890,N_2755,N_2763);
or U2891 (N_2891,N_2739,N_2756);
nor U2892 (N_2892,N_2770,N_2743);
nor U2893 (N_2893,N_2785,N_2713);
or U2894 (N_2894,N_2781,N_2762);
and U2895 (N_2895,N_2773,N_2713);
nand U2896 (N_2896,N_2738,N_2711);
nand U2897 (N_2897,N_2765,N_2715);
nand U2898 (N_2898,N_2770,N_2793);
nor U2899 (N_2899,N_2766,N_2773);
nand U2900 (N_2900,N_2842,N_2849);
and U2901 (N_2901,N_2868,N_2888);
nand U2902 (N_2902,N_2884,N_2808);
nor U2903 (N_2903,N_2810,N_2855);
nand U2904 (N_2904,N_2850,N_2837);
nor U2905 (N_2905,N_2839,N_2805);
or U2906 (N_2906,N_2860,N_2800);
nor U2907 (N_2907,N_2823,N_2886);
or U2908 (N_2908,N_2829,N_2834);
or U2909 (N_2909,N_2831,N_2867);
and U2910 (N_2910,N_2802,N_2865);
nor U2911 (N_2911,N_2817,N_2896);
or U2912 (N_2912,N_2891,N_2811);
and U2913 (N_2913,N_2895,N_2876);
nand U2914 (N_2914,N_2846,N_2851);
nor U2915 (N_2915,N_2813,N_2852);
nand U2916 (N_2916,N_2821,N_2807);
or U2917 (N_2917,N_2801,N_2832);
and U2918 (N_2918,N_2824,N_2804);
nand U2919 (N_2919,N_2848,N_2883);
nor U2920 (N_2920,N_2841,N_2871);
nand U2921 (N_2921,N_2844,N_2815);
nand U2922 (N_2922,N_2872,N_2897);
nand U2923 (N_2923,N_2899,N_2887);
nor U2924 (N_2924,N_2892,N_2819);
nand U2925 (N_2925,N_2803,N_2882);
nand U2926 (N_2926,N_2854,N_2835);
and U2927 (N_2927,N_2863,N_2853);
xnor U2928 (N_2928,N_2893,N_2856);
nand U2929 (N_2929,N_2830,N_2869);
nor U2930 (N_2930,N_2875,N_2814);
nor U2931 (N_2931,N_2866,N_2827);
nor U2932 (N_2932,N_2845,N_2881);
nand U2933 (N_2933,N_2859,N_2877);
xor U2934 (N_2934,N_2879,N_2889);
nand U2935 (N_2935,N_2862,N_2885);
or U2936 (N_2936,N_2843,N_2858);
nand U2937 (N_2937,N_2878,N_2828);
and U2938 (N_2938,N_2864,N_2873);
nor U2939 (N_2939,N_2826,N_2820);
or U2940 (N_2940,N_2822,N_2833);
nand U2941 (N_2941,N_2812,N_2857);
nor U2942 (N_2942,N_2818,N_2806);
and U2943 (N_2943,N_2816,N_2840);
nor U2944 (N_2944,N_2836,N_2870);
or U2945 (N_2945,N_2825,N_2890);
or U2946 (N_2946,N_2880,N_2894);
nand U2947 (N_2947,N_2874,N_2847);
nor U2948 (N_2948,N_2898,N_2861);
or U2949 (N_2949,N_2838,N_2809);
or U2950 (N_2950,N_2816,N_2872);
nor U2951 (N_2951,N_2869,N_2820);
and U2952 (N_2952,N_2800,N_2865);
xnor U2953 (N_2953,N_2810,N_2846);
and U2954 (N_2954,N_2841,N_2880);
and U2955 (N_2955,N_2882,N_2873);
and U2956 (N_2956,N_2830,N_2876);
nor U2957 (N_2957,N_2812,N_2871);
nor U2958 (N_2958,N_2858,N_2839);
or U2959 (N_2959,N_2848,N_2825);
or U2960 (N_2960,N_2858,N_2878);
nor U2961 (N_2961,N_2872,N_2878);
and U2962 (N_2962,N_2874,N_2844);
nor U2963 (N_2963,N_2814,N_2802);
nor U2964 (N_2964,N_2845,N_2842);
nand U2965 (N_2965,N_2892,N_2862);
and U2966 (N_2966,N_2800,N_2833);
or U2967 (N_2967,N_2836,N_2874);
nor U2968 (N_2968,N_2833,N_2818);
and U2969 (N_2969,N_2880,N_2825);
or U2970 (N_2970,N_2885,N_2894);
nor U2971 (N_2971,N_2829,N_2815);
nand U2972 (N_2972,N_2867,N_2839);
nor U2973 (N_2973,N_2861,N_2832);
nor U2974 (N_2974,N_2809,N_2892);
nor U2975 (N_2975,N_2833,N_2841);
and U2976 (N_2976,N_2802,N_2896);
xnor U2977 (N_2977,N_2880,N_2813);
and U2978 (N_2978,N_2854,N_2853);
nor U2979 (N_2979,N_2804,N_2888);
nand U2980 (N_2980,N_2846,N_2830);
or U2981 (N_2981,N_2810,N_2803);
or U2982 (N_2982,N_2849,N_2882);
nor U2983 (N_2983,N_2854,N_2852);
and U2984 (N_2984,N_2828,N_2814);
nor U2985 (N_2985,N_2898,N_2849);
nand U2986 (N_2986,N_2862,N_2864);
and U2987 (N_2987,N_2879,N_2850);
nand U2988 (N_2988,N_2819,N_2845);
or U2989 (N_2989,N_2872,N_2823);
or U2990 (N_2990,N_2840,N_2849);
and U2991 (N_2991,N_2885,N_2836);
and U2992 (N_2992,N_2868,N_2850);
nor U2993 (N_2993,N_2849,N_2836);
or U2994 (N_2994,N_2865,N_2861);
nor U2995 (N_2995,N_2840,N_2831);
or U2996 (N_2996,N_2814,N_2886);
xnor U2997 (N_2997,N_2810,N_2835);
nor U2998 (N_2998,N_2803,N_2890);
xnor U2999 (N_2999,N_2848,N_2894);
nor U3000 (N_3000,N_2928,N_2915);
nor U3001 (N_3001,N_2964,N_2972);
or U3002 (N_3002,N_2983,N_2918);
nor U3003 (N_3003,N_2981,N_2906);
nor U3004 (N_3004,N_2989,N_2969);
and U3005 (N_3005,N_2910,N_2999);
xor U3006 (N_3006,N_2976,N_2952);
and U3007 (N_3007,N_2908,N_2948);
nor U3008 (N_3008,N_2987,N_2951);
nand U3009 (N_3009,N_2943,N_2991);
or U3010 (N_3010,N_2922,N_2960);
or U3011 (N_3011,N_2916,N_2900);
nand U3012 (N_3012,N_2958,N_2944);
nor U3013 (N_3013,N_2978,N_2947);
or U3014 (N_3014,N_2998,N_2901);
nand U3015 (N_3015,N_2936,N_2946);
nand U3016 (N_3016,N_2970,N_2933);
and U3017 (N_3017,N_2974,N_2979);
nor U3018 (N_3018,N_2977,N_2965);
or U3019 (N_3019,N_2907,N_2990);
nor U3020 (N_3020,N_2919,N_2996);
nor U3021 (N_3021,N_2993,N_2961);
and U3022 (N_3022,N_2911,N_2945);
nor U3023 (N_3023,N_2992,N_2938);
or U3024 (N_3024,N_2927,N_2931);
or U3025 (N_3025,N_2929,N_2917);
nor U3026 (N_3026,N_2966,N_2980);
nor U3027 (N_3027,N_2973,N_2937);
and U3028 (N_3028,N_2967,N_2953);
nor U3029 (N_3029,N_2984,N_2985);
nor U3030 (N_3030,N_2913,N_2940);
or U3031 (N_3031,N_2971,N_2941);
nor U3032 (N_3032,N_2986,N_2904);
or U3033 (N_3033,N_2935,N_2950);
or U3034 (N_3034,N_2954,N_2924);
and U3035 (N_3035,N_2975,N_2956);
and U3036 (N_3036,N_2939,N_2903);
or U3037 (N_3037,N_2914,N_2997);
nor U3038 (N_3038,N_2921,N_2923);
and U3039 (N_3039,N_2902,N_2925);
and U3040 (N_3040,N_2920,N_2957);
and U3041 (N_3041,N_2932,N_2905);
nor U3042 (N_3042,N_2988,N_2926);
nor U3043 (N_3043,N_2942,N_2968);
nor U3044 (N_3044,N_2959,N_2909);
or U3045 (N_3045,N_2995,N_2955);
or U3046 (N_3046,N_2930,N_2963);
nor U3047 (N_3047,N_2962,N_2949);
nand U3048 (N_3048,N_2994,N_2934);
and U3049 (N_3049,N_2982,N_2912);
nand U3050 (N_3050,N_2977,N_2912);
nor U3051 (N_3051,N_2922,N_2951);
and U3052 (N_3052,N_2946,N_2999);
xnor U3053 (N_3053,N_2947,N_2975);
nand U3054 (N_3054,N_2988,N_2975);
or U3055 (N_3055,N_2919,N_2917);
or U3056 (N_3056,N_2979,N_2998);
and U3057 (N_3057,N_2962,N_2977);
nor U3058 (N_3058,N_2990,N_2930);
nand U3059 (N_3059,N_2971,N_2934);
xnor U3060 (N_3060,N_2921,N_2948);
and U3061 (N_3061,N_2976,N_2951);
nor U3062 (N_3062,N_2928,N_2961);
and U3063 (N_3063,N_2948,N_2982);
nor U3064 (N_3064,N_2996,N_2905);
xnor U3065 (N_3065,N_2920,N_2950);
xor U3066 (N_3066,N_2999,N_2986);
and U3067 (N_3067,N_2946,N_2916);
xnor U3068 (N_3068,N_2942,N_2987);
nor U3069 (N_3069,N_2982,N_2923);
xnor U3070 (N_3070,N_2951,N_2911);
nor U3071 (N_3071,N_2900,N_2999);
and U3072 (N_3072,N_2973,N_2914);
nor U3073 (N_3073,N_2930,N_2956);
nand U3074 (N_3074,N_2978,N_2990);
nand U3075 (N_3075,N_2922,N_2995);
or U3076 (N_3076,N_2953,N_2901);
and U3077 (N_3077,N_2952,N_2963);
or U3078 (N_3078,N_2988,N_2971);
nand U3079 (N_3079,N_2988,N_2962);
xnor U3080 (N_3080,N_2957,N_2995);
nand U3081 (N_3081,N_2919,N_2907);
nand U3082 (N_3082,N_2913,N_2930);
nand U3083 (N_3083,N_2913,N_2958);
xnor U3084 (N_3084,N_2961,N_2919);
and U3085 (N_3085,N_2906,N_2989);
nor U3086 (N_3086,N_2968,N_2931);
nor U3087 (N_3087,N_2974,N_2960);
nand U3088 (N_3088,N_2942,N_2911);
nor U3089 (N_3089,N_2974,N_2936);
and U3090 (N_3090,N_2993,N_2977);
nand U3091 (N_3091,N_2977,N_2917);
nor U3092 (N_3092,N_2981,N_2985);
or U3093 (N_3093,N_2976,N_2900);
nor U3094 (N_3094,N_2974,N_2981);
nor U3095 (N_3095,N_2960,N_2950);
nor U3096 (N_3096,N_2946,N_2919);
nand U3097 (N_3097,N_2914,N_2998);
nor U3098 (N_3098,N_2948,N_2936);
nand U3099 (N_3099,N_2986,N_2993);
nand U3100 (N_3100,N_3069,N_3038);
xor U3101 (N_3101,N_3031,N_3019);
and U3102 (N_3102,N_3018,N_3045);
or U3103 (N_3103,N_3003,N_3088);
nor U3104 (N_3104,N_3042,N_3005);
nand U3105 (N_3105,N_3048,N_3077);
nand U3106 (N_3106,N_3057,N_3040);
or U3107 (N_3107,N_3079,N_3051);
or U3108 (N_3108,N_3059,N_3063);
and U3109 (N_3109,N_3035,N_3036);
xnor U3110 (N_3110,N_3078,N_3013);
nand U3111 (N_3111,N_3027,N_3037);
nor U3112 (N_3112,N_3023,N_3039);
nand U3113 (N_3113,N_3058,N_3009);
nor U3114 (N_3114,N_3007,N_3074);
nor U3115 (N_3115,N_3070,N_3004);
or U3116 (N_3116,N_3091,N_3084);
xnor U3117 (N_3117,N_3030,N_3064);
and U3118 (N_3118,N_3028,N_3002);
or U3119 (N_3119,N_3010,N_3098);
xor U3120 (N_3120,N_3034,N_3089);
and U3121 (N_3121,N_3053,N_3072);
or U3122 (N_3122,N_3006,N_3021);
nor U3123 (N_3123,N_3015,N_3054);
xnor U3124 (N_3124,N_3050,N_3000);
or U3125 (N_3125,N_3087,N_3062);
nand U3126 (N_3126,N_3055,N_3076);
and U3127 (N_3127,N_3067,N_3043);
nand U3128 (N_3128,N_3032,N_3041);
or U3129 (N_3129,N_3099,N_3029);
or U3130 (N_3130,N_3094,N_3044);
nand U3131 (N_3131,N_3008,N_3090);
nand U3132 (N_3132,N_3014,N_3068);
and U3133 (N_3133,N_3024,N_3052);
nor U3134 (N_3134,N_3086,N_3097);
xor U3135 (N_3135,N_3022,N_3025);
nand U3136 (N_3136,N_3085,N_3011);
nand U3137 (N_3137,N_3075,N_3047);
and U3138 (N_3138,N_3061,N_3017);
and U3139 (N_3139,N_3096,N_3020);
nand U3140 (N_3140,N_3012,N_3073);
nand U3141 (N_3141,N_3081,N_3093);
nand U3142 (N_3142,N_3080,N_3065);
xnor U3143 (N_3143,N_3092,N_3016);
xnor U3144 (N_3144,N_3083,N_3060);
nor U3145 (N_3145,N_3026,N_3082);
nand U3146 (N_3146,N_3049,N_3046);
nor U3147 (N_3147,N_3001,N_3066);
nand U3148 (N_3148,N_3033,N_3095);
nor U3149 (N_3149,N_3056,N_3071);
nand U3150 (N_3150,N_3035,N_3009);
or U3151 (N_3151,N_3026,N_3009);
xor U3152 (N_3152,N_3043,N_3052);
nand U3153 (N_3153,N_3060,N_3086);
nor U3154 (N_3154,N_3045,N_3013);
and U3155 (N_3155,N_3079,N_3017);
and U3156 (N_3156,N_3070,N_3098);
nor U3157 (N_3157,N_3054,N_3003);
or U3158 (N_3158,N_3017,N_3099);
xor U3159 (N_3159,N_3009,N_3061);
nor U3160 (N_3160,N_3054,N_3057);
or U3161 (N_3161,N_3019,N_3067);
nor U3162 (N_3162,N_3066,N_3099);
or U3163 (N_3163,N_3093,N_3087);
nand U3164 (N_3164,N_3098,N_3053);
nand U3165 (N_3165,N_3081,N_3070);
nand U3166 (N_3166,N_3086,N_3063);
and U3167 (N_3167,N_3017,N_3055);
xor U3168 (N_3168,N_3082,N_3054);
nand U3169 (N_3169,N_3063,N_3057);
and U3170 (N_3170,N_3016,N_3052);
nor U3171 (N_3171,N_3016,N_3071);
or U3172 (N_3172,N_3009,N_3030);
nand U3173 (N_3173,N_3024,N_3075);
xnor U3174 (N_3174,N_3009,N_3006);
or U3175 (N_3175,N_3052,N_3061);
nand U3176 (N_3176,N_3009,N_3067);
or U3177 (N_3177,N_3031,N_3096);
xor U3178 (N_3178,N_3018,N_3095);
xor U3179 (N_3179,N_3029,N_3001);
nor U3180 (N_3180,N_3073,N_3089);
nand U3181 (N_3181,N_3090,N_3093);
or U3182 (N_3182,N_3020,N_3045);
and U3183 (N_3183,N_3057,N_3008);
nor U3184 (N_3184,N_3096,N_3015);
nor U3185 (N_3185,N_3073,N_3076);
or U3186 (N_3186,N_3075,N_3009);
or U3187 (N_3187,N_3045,N_3024);
xor U3188 (N_3188,N_3093,N_3070);
nor U3189 (N_3189,N_3040,N_3004);
and U3190 (N_3190,N_3043,N_3020);
xnor U3191 (N_3191,N_3007,N_3060);
xnor U3192 (N_3192,N_3039,N_3010);
nor U3193 (N_3193,N_3040,N_3065);
and U3194 (N_3194,N_3011,N_3096);
nand U3195 (N_3195,N_3094,N_3029);
and U3196 (N_3196,N_3053,N_3004);
nand U3197 (N_3197,N_3043,N_3042);
nand U3198 (N_3198,N_3048,N_3025);
nor U3199 (N_3199,N_3060,N_3041);
nor U3200 (N_3200,N_3161,N_3137);
or U3201 (N_3201,N_3192,N_3176);
xor U3202 (N_3202,N_3174,N_3177);
and U3203 (N_3203,N_3140,N_3104);
nand U3204 (N_3204,N_3189,N_3110);
nor U3205 (N_3205,N_3190,N_3120);
nor U3206 (N_3206,N_3107,N_3170);
nor U3207 (N_3207,N_3159,N_3133);
and U3208 (N_3208,N_3103,N_3151);
xor U3209 (N_3209,N_3135,N_3166);
nor U3210 (N_3210,N_3112,N_3165);
nand U3211 (N_3211,N_3187,N_3118);
nor U3212 (N_3212,N_3191,N_3119);
or U3213 (N_3213,N_3109,N_3129);
nor U3214 (N_3214,N_3155,N_3163);
or U3215 (N_3215,N_3132,N_3167);
nor U3216 (N_3216,N_3149,N_3100);
nand U3217 (N_3217,N_3168,N_3193);
xor U3218 (N_3218,N_3182,N_3127);
xnor U3219 (N_3219,N_3123,N_3144);
nor U3220 (N_3220,N_3136,N_3117);
nand U3221 (N_3221,N_3160,N_3181);
or U3222 (N_3222,N_3156,N_3121);
or U3223 (N_3223,N_3195,N_3124);
or U3224 (N_3224,N_3186,N_3134);
xnor U3225 (N_3225,N_3116,N_3102);
nand U3226 (N_3226,N_3194,N_3146);
or U3227 (N_3227,N_3115,N_3130);
or U3228 (N_3228,N_3114,N_3180);
nand U3229 (N_3229,N_3175,N_3122);
or U3230 (N_3230,N_3164,N_3172);
or U3231 (N_3231,N_3185,N_3128);
or U3232 (N_3232,N_3150,N_3162);
nor U3233 (N_3233,N_3153,N_3188);
or U3234 (N_3234,N_3173,N_3199);
nand U3235 (N_3235,N_3152,N_3111);
nor U3236 (N_3236,N_3178,N_3105);
nor U3237 (N_3237,N_3108,N_3197);
or U3238 (N_3238,N_3184,N_3198);
or U3239 (N_3239,N_3113,N_3147);
nand U3240 (N_3240,N_3196,N_3125);
or U3241 (N_3241,N_3101,N_3126);
and U3242 (N_3242,N_3171,N_3158);
nor U3243 (N_3243,N_3148,N_3143);
xor U3244 (N_3244,N_3138,N_3179);
or U3245 (N_3245,N_3183,N_3169);
nor U3246 (N_3246,N_3131,N_3106);
nand U3247 (N_3247,N_3145,N_3139);
or U3248 (N_3248,N_3141,N_3154);
nand U3249 (N_3249,N_3157,N_3142);
nor U3250 (N_3250,N_3104,N_3176);
and U3251 (N_3251,N_3121,N_3131);
and U3252 (N_3252,N_3177,N_3184);
nand U3253 (N_3253,N_3105,N_3152);
or U3254 (N_3254,N_3142,N_3185);
or U3255 (N_3255,N_3134,N_3121);
nor U3256 (N_3256,N_3115,N_3155);
xor U3257 (N_3257,N_3134,N_3171);
and U3258 (N_3258,N_3186,N_3199);
and U3259 (N_3259,N_3166,N_3177);
or U3260 (N_3260,N_3105,N_3123);
and U3261 (N_3261,N_3128,N_3118);
nand U3262 (N_3262,N_3102,N_3169);
and U3263 (N_3263,N_3145,N_3104);
and U3264 (N_3264,N_3167,N_3148);
nand U3265 (N_3265,N_3199,N_3101);
and U3266 (N_3266,N_3138,N_3189);
or U3267 (N_3267,N_3161,N_3196);
and U3268 (N_3268,N_3106,N_3174);
nor U3269 (N_3269,N_3140,N_3107);
nor U3270 (N_3270,N_3189,N_3158);
xnor U3271 (N_3271,N_3176,N_3191);
and U3272 (N_3272,N_3197,N_3100);
nand U3273 (N_3273,N_3187,N_3156);
and U3274 (N_3274,N_3148,N_3116);
nor U3275 (N_3275,N_3196,N_3136);
nand U3276 (N_3276,N_3162,N_3185);
nor U3277 (N_3277,N_3110,N_3138);
and U3278 (N_3278,N_3192,N_3104);
nand U3279 (N_3279,N_3159,N_3182);
and U3280 (N_3280,N_3174,N_3105);
nand U3281 (N_3281,N_3183,N_3178);
or U3282 (N_3282,N_3196,N_3118);
nand U3283 (N_3283,N_3125,N_3116);
nor U3284 (N_3284,N_3115,N_3176);
nand U3285 (N_3285,N_3142,N_3191);
nor U3286 (N_3286,N_3195,N_3170);
and U3287 (N_3287,N_3164,N_3110);
and U3288 (N_3288,N_3177,N_3159);
nor U3289 (N_3289,N_3129,N_3193);
nand U3290 (N_3290,N_3185,N_3119);
and U3291 (N_3291,N_3136,N_3147);
and U3292 (N_3292,N_3144,N_3174);
and U3293 (N_3293,N_3124,N_3126);
or U3294 (N_3294,N_3168,N_3185);
xnor U3295 (N_3295,N_3145,N_3180);
nand U3296 (N_3296,N_3169,N_3153);
and U3297 (N_3297,N_3164,N_3153);
nand U3298 (N_3298,N_3152,N_3164);
nand U3299 (N_3299,N_3121,N_3128);
or U3300 (N_3300,N_3281,N_3272);
or U3301 (N_3301,N_3263,N_3237);
xnor U3302 (N_3302,N_3278,N_3227);
nand U3303 (N_3303,N_3239,N_3211);
xor U3304 (N_3304,N_3298,N_3257);
nand U3305 (N_3305,N_3215,N_3268);
or U3306 (N_3306,N_3259,N_3222);
nand U3307 (N_3307,N_3238,N_3212);
nor U3308 (N_3308,N_3214,N_3209);
nor U3309 (N_3309,N_3210,N_3225);
or U3310 (N_3310,N_3258,N_3203);
nor U3311 (N_3311,N_3284,N_3274);
nor U3312 (N_3312,N_3226,N_3269);
nor U3313 (N_3313,N_3293,N_3200);
nor U3314 (N_3314,N_3275,N_3283);
nor U3315 (N_3315,N_3219,N_3250);
xor U3316 (N_3316,N_3236,N_3299);
nand U3317 (N_3317,N_3246,N_3201);
nand U3318 (N_3318,N_3218,N_3213);
or U3319 (N_3319,N_3206,N_3276);
or U3320 (N_3320,N_3279,N_3229);
or U3321 (N_3321,N_3231,N_3232);
nand U3322 (N_3322,N_3234,N_3248);
xnor U3323 (N_3323,N_3296,N_3255);
and U3324 (N_3324,N_3273,N_3265);
and U3325 (N_3325,N_3251,N_3297);
and U3326 (N_3326,N_3260,N_3242);
xor U3327 (N_3327,N_3261,N_3205);
or U3328 (N_3328,N_3267,N_3271);
nor U3329 (N_3329,N_3264,N_3204);
nand U3330 (N_3330,N_3217,N_3254);
nor U3331 (N_3331,N_3266,N_3224);
or U3332 (N_3332,N_3253,N_3290);
nor U3333 (N_3333,N_3230,N_3292);
or U3334 (N_3334,N_3243,N_3286);
or U3335 (N_3335,N_3277,N_3262);
xnor U3336 (N_3336,N_3285,N_3282);
or U3337 (N_3337,N_3291,N_3287);
or U3338 (N_3338,N_3207,N_3228);
or U3339 (N_3339,N_3216,N_3240);
and U3340 (N_3340,N_3223,N_3244);
nand U3341 (N_3341,N_3247,N_3294);
or U3342 (N_3342,N_3202,N_3235);
nor U3343 (N_3343,N_3270,N_3220);
nand U3344 (N_3344,N_3208,N_3289);
or U3345 (N_3345,N_3245,N_3288);
and U3346 (N_3346,N_3221,N_3249);
or U3347 (N_3347,N_3256,N_3233);
nand U3348 (N_3348,N_3295,N_3280);
nor U3349 (N_3349,N_3252,N_3241);
nand U3350 (N_3350,N_3213,N_3298);
and U3351 (N_3351,N_3267,N_3288);
xor U3352 (N_3352,N_3274,N_3217);
nor U3353 (N_3353,N_3231,N_3282);
nand U3354 (N_3354,N_3296,N_3281);
nand U3355 (N_3355,N_3201,N_3295);
nor U3356 (N_3356,N_3242,N_3248);
and U3357 (N_3357,N_3235,N_3201);
nor U3358 (N_3358,N_3298,N_3267);
nand U3359 (N_3359,N_3282,N_3224);
nand U3360 (N_3360,N_3276,N_3293);
and U3361 (N_3361,N_3299,N_3213);
xor U3362 (N_3362,N_3215,N_3206);
and U3363 (N_3363,N_3211,N_3251);
nand U3364 (N_3364,N_3249,N_3280);
nand U3365 (N_3365,N_3228,N_3285);
or U3366 (N_3366,N_3226,N_3248);
nand U3367 (N_3367,N_3297,N_3273);
and U3368 (N_3368,N_3290,N_3217);
and U3369 (N_3369,N_3255,N_3274);
and U3370 (N_3370,N_3234,N_3246);
and U3371 (N_3371,N_3227,N_3283);
or U3372 (N_3372,N_3241,N_3240);
nor U3373 (N_3373,N_3291,N_3252);
xor U3374 (N_3374,N_3241,N_3289);
nor U3375 (N_3375,N_3214,N_3236);
nand U3376 (N_3376,N_3249,N_3283);
nand U3377 (N_3377,N_3206,N_3248);
nor U3378 (N_3378,N_3243,N_3271);
xor U3379 (N_3379,N_3212,N_3296);
nand U3380 (N_3380,N_3284,N_3211);
and U3381 (N_3381,N_3211,N_3259);
and U3382 (N_3382,N_3297,N_3212);
nor U3383 (N_3383,N_3202,N_3268);
xnor U3384 (N_3384,N_3290,N_3270);
and U3385 (N_3385,N_3245,N_3210);
or U3386 (N_3386,N_3270,N_3209);
nor U3387 (N_3387,N_3241,N_3260);
or U3388 (N_3388,N_3296,N_3239);
nand U3389 (N_3389,N_3224,N_3278);
nand U3390 (N_3390,N_3227,N_3221);
xnor U3391 (N_3391,N_3271,N_3294);
nor U3392 (N_3392,N_3258,N_3275);
or U3393 (N_3393,N_3244,N_3263);
nand U3394 (N_3394,N_3208,N_3211);
nor U3395 (N_3395,N_3246,N_3217);
nor U3396 (N_3396,N_3286,N_3275);
and U3397 (N_3397,N_3245,N_3264);
or U3398 (N_3398,N_3252,N_3287);
nor U3399 (N_3399,N_3216,N_3255);
or U3400 (N_3400,N_3304,N_3336);
and U3401 (N_3401,N_3319,N_3330);
or U3402 (N_3402,N_3369,N_3308);
xor U3403 (N_3403,N_3337,N_3340);
nor U3404 (N_3404,N_3302,N_3310);
nand U3405 (N_3405,N_3358,N_3375);
nor U3406 (N_3406,N_3339,N_3344);
nand U3407 (N_3407,N_3305,N_3354);
nand U3408 (N_3408,N_3356,N_3325);
and U3409 (N_3409,N_3388,N_3355);
nor U3410 (N_3410,N_3377,N_3360);
or U3411 (N_3411,N_3391,N_3312);
nor U3412 (N_3412,N_3342,N_3301);
nand U3413 (N_3413,N_3363,N_3353);
nor U3414 (N_3414,N_3306,N_3366);
or U3415 (N_3415,N_3365,N_3396);
nor U3416 (N_3416,N_3381,N_3364);
xnor U3417 (N_3417,N_3320,N_3303);
nor U3418 (N_3418,N_3379,N_3392);
and U3419 (N_3419,N_3347,N_3368);
nand U3420 (N_3420,N_3362,N_3359);
and U3421 (N_3421,N_3346,N_3398);
and U3422 (N_3422,N_3386,N_3328);
nand U3423 (N_3423,N_3350,N_3341);
xnor U3424 (N_3424,N_3373,N_3370);
or U3425 (N_3425,N_3329,N_3393);
nand U3426 (N_3426,N_3399,N_3390);
and U3427 (N_3427,N_3324,N_3333);
nor U3428 (N_3428,N_3385,N_3378);
or U3429 (N_3429,N_3311,N_3372);
nor U3430 (N_3430,N_3327,N_3351);
xnor U3431 (N_3431,N_3397,N_3332);
nand U3432 (N_3432,N_3309,N_3331);
nor U3433 (N_3433,N_3349,N_3321);
nand U3434 (N_3434,N_3334,N_3314);
nor U3435 (N_3435,N_3352,N_3322);
and U3436 (N_3436,N_3316,N_3361);
nor U3437 (N_3437,N_3376,N_3383);
nor U3438 (N_3438,N_3343,N_3382);
nand U3439 (N_3439,N_3318,N_3335);
or U3440 (N_3440,N_3357,N_3394);
nor U3441 (N_3441,N_3338,N_3380);
or U3442 (N_3442,N_3389,N_3367);
nand U3443 (N_3443,N_3315,N_3384);
or U3444 (N_3444,N_3348,N_3313);
or U3445 (N_3445,N_3387,N_3326);
or U3446 (N_3446,N_3395,N_3300);
nand U3447 (N_3447,N_3371,N_3317);
or U3448 (N_3448,N_3345,N_3374);
xor U3449 (N_3449,N_3307,N_3323);
or U3450 (N_3450,N_3348,N_3331);
and U3451 (N_3451,N_3391,N_3397);
nor U3452 (N_3452,N_3328,N_3303);
nor U3453 (N_3453,N_3358,N_3352);
nor U3454 (N_3454,N_3354,N_3322);
nor U3455 (N_3455,N_3321,N_3367);
or U3456 (N_3456,N_3361,N_3326);
nor U3457 (N_3457,N_3342,N_3372);
nor U3458 (N_3458,N_3315,N_3336);
or U3459 (N_3459,N_3350,N_3387);
nand U3460 (N_3460,N_3394,N_3345);
nand U3461 (N_3461,N_3334,N_3316);
nand U3462 (N_3462,N_3370,N_3361);
nor U3463 (N_3463,N_3301,N_3308);
or U3464 (N_3464,N_3389,N_3316);
or U3465 (N_3465,N_3310,N_3342);
xor U3466 (N_3466,N_3321,N_3389);
nand U3467 (N_3467,N_3302,N_3317);
nand U3468 (N_3468,N_3337,N_3333);
or U3469 (N_3469,N_3396,N_3320);
nor U3470 (N_3470,N_3367,N_3394);
nand U3471 (N_3471,N_3361,N_3378);
and U3472 (N_3472,N_3340,N_3350);
nor U3473 (N_3473,N_3388,N_3387);
and U3474 (N_3474,N_3381,N_3350);
and U3475 (N_3475,N_3368,N_3322);
or U3476 (N_3476,N_3353,N_3311);
nor U3477 (N_3477,N_3373,N_3367);
or U3478 (N_3478,N_3394,N_3365);
nor U3479 (N_3479,N_3303,N_3354);
nor U3480 (N_3480,N_3377,N_3382);
nor U3481 (N_3481,N_3397,N_3305);
nor U3482 (N_3482,N_3322,N_3357);
or U3483 (N_3483,N_3375,N_3322);
and U3484 (N_3484,N_3349,N_3372);
and U3485 (N_3485,N_3369,N_3325);
nand U3486 (N_3486,N_3374,N_3396);
nand U3487 (N_3487,N_3339,N_3365);
nand U3488 (N_3488,N_3399,N_3338);
or U3489 (N_3489,N_3399,N_3314);
or U3490 (N_3490,N_3309,N_3306);
nand U3491 (N_3491,N_3335,N_3370);
or U3492 (N_3492,N_3331,N_3379);
nor U3493 (N_3493,N_3367,N_3378);
and U3494 (N_3494,N_3321,N_3335);
and U3495 (N_3495,N_3363,N_3328);
nand U3496 (N_3496,N_3382,N_3327);
nor U3497 (N_3497,N_3376,N_3359);
nand U3498 (N_3498,N_3319,N_3382);
nor U3499 (N_3499,N_3380,N_3358);
and U3500 (N_3500,N_3484,N_3454);
nand U3501 (N_3501,N_3445,N_3467);
or U3502 (N_3502,N_3490,N_3450);
nand U3503 (N_3503,N_3459,N_3400);
xor U3504 (N_3504,N_3478,N_3469);
nand U3505 (N_3505,N_3429,N_3472);
nand U3506 (N_3506,N_3499,N_3458);
and U3507 (N_3507,N_3434,N_3456);
nor U3508 (N_3508,N_3479,N_3406);
and U3509 (N_3509,N_3482,N_3480);
nor U3510 (N_3510,N_3465,N_3404);
xnor U3511 (N_3511,N_3495,N_3417);
xnor U3512 (N_3512,N_3420,N_3428);
nor U3513 (N_3513,N_3460,N_3413);
nand U3514 (N_3514,N_3475,N_3438);
or U3515 (N_3515,N_3470,N_3442);
nand U3516 (N_3516,N_3453,N_3443);
nand U3517 (N_3517,N_3447,N_3405);
nand U3518 (N_3518,N_3486,N_3426);
xor U3519 (N_3519,N_3457,N_3449);
or U3520 (N_3520,N_3435,N_3489);
and U3521 (N_3521,N_3410,N_3473);
nand U3522 (N_3522,N_3487,N_3485);
and U3523 (N_3523,N_3463,N_3461);
or U3524 (N_3524,N_3421,N_3431);
or U3525 (N_3525,N_3481,N_3476);
nand U3526 (N_3526,N_3407,N_3418);
nor U3527 (N_3527,N_3462,N_3441);
nor U3528 (N_3528,N_3436,N_3412);
nand U3529 (N_3529,N_3409,N_3493);
nor U3530 (N_3530,N_3464,N_3433);
or U3531 (N_3531,N_3422,N_3403);
nand U3532 (N_3532,N_3466,N_3419);
xor U3533 (N_3533,N_3492,N_3427);
and U3534 (N_3534,N_3483,N_3411);
nand U3535 (N_3535,N_3401,N_3451);
nor U3536 (N_3536,N_3477,N_3416);
and U3537 (N_3537,N_3402,N_3474);
and U3538 (N_3538,N_3491,N_3468);
nor U3539 (N_3539,N_3430,N_3446);
or U3540 (N_3540,N_3471,N_3497);
nand U3541 (N_3541,N_3424,N_3444);
nor U3542 (N_3542,N_3439,N_3452);
and U3543 (N_3543,N_3408,N_3423);
or U3544 (N_3544,N_3425,N_3432);
xor U3545 (N_3545,N_3415,N_3414);
and U3546 (N_3546,N_3437,N_3455);
and U3547 (N_3547,N_3448,N_3498);
nor U3548 (N_3548,N_3494,N_3488);
and U3549 (N_3549,N_3496,N_3440);
nand U3550 (N_3550,N_3458,N_3401);
nor U3551 (N_3551,N_3473,N_3496);
and U3552 (N_3552,N_3425,N_3458);
or U3553 (N_3553,N_3401,N_3497);
xnor U3554 (N_3554,N_3429,N_3480);
nand U3555 (N_3555,N_3404,N_3421);
and U3556 (N_3556,N_3411,N_3420);
nand U3557 (N_3557,N_3486,N_3408);
nor U3558 (N_3558,N_3448,N_3497);
nand U3559 (N_3559,N_3433,N_3427);
nand U3560 (N_3560,N_3477,N_3452);
nor U3561 (N_3561,N_3434,N_3438);
and U3562 (N_3562,N_3410,N_3443);
nor U3563 (N_3563,N_3472,N_3443);
and U3564 (N_3564,N_3427,N_3456);
and U3565 (N_3565,N_3488,N_3433);
or U3566 (N_3566,N_3449,N_3482);
and U3567 (N_3567,N_3490,N_3415);
xnor U3568 (N_3568,N_3467,N_3488);
nand U3569 (N_3569,N_3476,N_3445);
or U3570 (N_3570,N_3430,N_3486);
nor U3571 (N_3571,N_3419,N_3488);
nand U3572 (N_3572,N_3407,N_3492);
xor U3573 (N_3573,N_3440,N_3464);
or U3574 (N_3574,N_3441,N_3400);
or U3575 (N_3575,N_3429,N_3417);
nand U3576 (N_3576,N_3416,N_3493);
nor U3577 (N_3577,N_3410,N_3486);
or U3578 (N_3578,N_3402,N_3410);
or U3579 (N_3579,N_3454,N_3435);
and U3580 (N_3580,N_3411,N_3484);
or U3581 (N_3581,N_3435,N_3467);
xor U3582 (N_3582,N_3490,N_3484);
nor U3583 (N_3583,N_3412,N_3459);
nor U3584 (N_3584,N_3452,N_3447);
and U3585 (N_3585,N_3498,N_3467);
xnor U3586 (N_3586,N_3447,N_3401);
nand U3587 (N_3587,N_3414,N_3497);
and U3588 (N_3588,N_3446,N_3475);
xor U3589 (N_3589,N_3425,N_3484);
nand U3590 (N_3590,N_3454,N_3406);
or U3591 (N_3591,N_3404,N_3464);
nand U3592 (N_3592,N_3447,N_3437);
or U3593 (N_3593,N_3433,N_3489);
or U3594 (N_3594,N_3487,N_3430);
and U3595 (N_3595,N_3408,N_3496);
xnor U3596 (N_3596,N_3407,N_3454);
and U3597 (N_3597,N_3470,N_3423);
nor U3598 (N_3598,N_3420,N_3458);
nor U3599 (N_3599,N_3444,N_3435);
nand U3600 (N_3600,N_3548,N_3569);
nor U3601 (N_3601,N_3572,N_3522);
or U3602 (N_3602,N_3588,N_3502);
nand U3603 (N_3603,N_3560,N_3583);
nor U3604 (N_3604,N_3562,N_3516);
and U3605 (N_3605,N_3526,N_3556);
nand U3606 (N_3606,N_3571,N_3555);
or U3607 (N_3607,N_3520,N_3557);
nand U3608 (N_3608,N_3512,N_3515);
nor U3609 (N_3609,N_3552,N_3500);
nor U3610 (N_3610,N_3517,N_3518);
nor U3611 (N_3611,N_3582,N_3590);
and U3612 (N_3612,N_3544,N_3508);
or U3613 (N_3613,N_3550,N_3598);
and U3614 (N_3614,N_3510,N_3573);
nand U3615 (N_3615,N_3570,N_3514);
nor U3616 (N_3616,N_3545,N_3533);
nand U3617 (N_3617,N_3568,N_3593);
nand U3618 (N_3618,N_3575,N_3595);
nor U3619 (N_3619,N_3592,N_3524);
and U3620 (N_3620,N_3535,N_3509);
or U3621 (N_3621,N_3576,N_3561);
nor U3622 (N_3622,N_3580,N_3534);
and U3623 (N_3623,N_3519,N_3530);
nand U3624 (N_3624,N_3536,N_3585);
nor U3625 (N_3625,N_3577,N_3551);
and U3626 (N_3626,N_3527,N_3532);
nand U3627 (N_3627,N_3559,N_3506);
and U3628 (N_3628,N_3540,N_3566);
and U3629 (N_3629,N_3538,N_3529);
and U3630 (N_3630,N_3589,N_3541);
nor U3631 (N_3631,N_3504,N_3521);
nor U3632 (N_3632,N_3581,N_3507);
nor U3633 (N_3633,N_3554,N_3505);
nor U3634 (N_3634,N_3564,N_3525);
or U3635 (N_3635,N_3543,N_3539);
and U3636 (N_3636,N_3537,N_3511);
or U3637 (N_3637,N_3547,N_3546);
nor U3638 (N_3638,N_3599,N_3563);
and U3639 (N_3639,N_3594,N_3565);
nor U3640 (N_3640,N_3596,N_3587);
or U3641 (N_3641,N_3567,N_3584);
and U3642 (N_3642,N_3523,N_3597);
or U3643 (N_3643,N_3586,N_3549);
and U3644 (N_3644,N_3528,N_3579);
or U3645 (N_3645,N_3558,N_3513);
nor U3646 (N_3646,N_3531,N_3574);
nand U3647 (N_3647,N_3503,N_3542);
nor U3648 (N_3648,N_3578,N_3591);
and U3649 (N_3649,N_3501,N_3553);
and U3650 (N_3650,N_3546,N_3552);
and U3651 (N_3651,N_3536,N_3513);
or U3652 (N_3652,N_3516,N_3510);
nor U3653 (N_3653,N_3505,N_3592);
nand U3654 (N_3654,N_3583,N_3596);
nand U3655 (N_3655,N_3520,N_3523);
nor U3656 (N_3656,N_3592,N_3526);
and U3657 (N_3657,N_3547,N_3574);
xnor U3658 (N_3658,N_3510,N_3595);
and U3659 (N_3659,N_3584,N_3556);
or U3660 (N_3660,N_3566,N_3541);
and U3661 (N_3661,N_3548,N_3527);
nor U3662 (N_3662,N_3517,N_3506);
and U3663 (N_3663,N_3542,N_3597);
nor U3664 (N_3664,N_3550,N_3545);
or U3665 (N_3665,N_3502,N_3562);
nor U3666 (N_3666,N_3508,N_3583);
nor U3667 (N_3667,N_3599,N_3590);
and U3668 (N_3668,N_3546,N_3537);
xnor U3669 (N_3669,N_3544,N_3532);
or U3670 (N_3670,N_3518,N_3593);
nor U3671 (N_3671,N_3544,N_3536);
xor U3672 (N_3672,N_3573,N_3506);
nor U3673 (N_3673,N_3568,N_3523);
nor U3674 (N_3674,N_3526,N_3572);
nand U3675 (N_3675,N_3514,N_3534);
and U3676 (N_3676,N_3535,N_3511);
or U3677 (N_3677,N_3554,N_3537);
nand U3678 (N_3678,N_3534,N_3577);
nand U3679 (N_3679,N_3532,N_3592);
xor U3680 (N_3680,N_3502,N_3520);
and U3681 (N_3681,N_3513,N_3509);
and U3682 (N_3682,N_3551,N_3503);
xnor U3683 (N_3683,N_3577,N_3545);
xor U3684 (N_3684,N_3528,N_3543);
nor U3685 (N_3685,N_3506,N_3584);
or U3686 (N_3686,N_3554,N_3592);
nand U3687 (N_3687,N_3511,N_3583);
nor U3688 (N_3688,N_3588,N_3511);
xnor U3689 (N_3689,N_3520,N_3525);
or U3690 (N_3690,N_3539,N_3574);
or U3691 (N_3691,N_3549,N_3512);
nor U3692 (N_3692,N_3572,N_3528);
nand U3693 (N_3693,N_3532,N_3579);
or U3694 (N_3694,N_3503,N_3548);
and U3695 (N_3695,N_3500,N_3532);
nor U3696 (N_3696,N_3578,N_3531);
or U3697 (N_3697,N_3537,N_3595);
xnor U3698 (N_3698,N_3510,N_3597);
nand U3699 (N_3699,N_3570,N_3590);
xnor U3700 (N_3700,N_3649,N_3638);
xor U3701 (N_3701,N_3617,N_3600);
nor U3702 (N_3702,N_3667,N_3615);
or U3703 (N_3703,N_3616,N_3634);
or U3704 (N_3704,N_3627,N_3613);
nand U3705 (N_3705,N_3620,N_3640);
or U3706 (N_3706,N_3693,N_3670);
or U3707 (N_3707,N_3607,N_3653);
or U3708 (N_3708,N_3671,N_3680);
nand U3709 (N_3709,N_3602,N_3659);
or U3710 (N_3710,N_3677,N_3655);
xor U3711 (N_3711,N_3631,N_3665);
nor U3712 (N_3712,N_3623,N_3682);
nor U3713 (N_3713,N_3699,N_3645);
xor U3714 (N_3714,N_3619,N_3611);
nor U3715 (N_3715,N_3635,N_3652);
or U3716 (N_3716,N_3674,N_3637);
nand U3717 (N_3717,N_3633,N_3609);
or U3718 (N_3718,N_3664,N_3606);
and U3719 (N_3719,N_3698,N_3610);
nand U3720 (N_3720,N_3690,N_3605);
nor U3721 (N_3721,N_3668,N_3678);
and U3722 (N_3722,N_3644,N_3647);
and U3723 (N_3723,N_3662,N_3642);
nor U3724 (N_3724,N_3684,N_3650);
xnor U3725 (N_3725,N_3604,N_3639);
nand U3726 (N_3726,N_3681,N_3679);
and U3727 (N_3727,N_3694,N_3622);
xnor U3728 (N_3728,N_3603,N_3695);
or U3729 (N_3729,N_3646,N_3641);
nor U3730 (N_3730,N_3657,N_3656);
nand U3731 (N_3731,N_3686,N_3621);
nor U3732 (N_3732,N_3687,N_3643);
and U3733 (N_3733,N_3660,N_3692);
xor U3734 (N_3734,N_3654,N_3636);
nor U3735 (N_3735,N_3697,N_3629);
and U3736 (N_3736,N_3632,N_3663);
nand U3737 (N_3737,N_3651,N_3628);
nand U3738 (N_3738,N_3688,N_3691);
xor U3739 (N_3739,N_3658,N_3672);
and U3740 (N_3740,N_3685,N_3648);
nor U3741 (N_3741,N_3608,N_3624);
nand U3742 (N_3742,N_3618,N_3614);
nand U3743 (N_3743,N_3625,N_3661);
and U3744 (N_3744,N_3612,N_3666);
nand U3745 (N_3745,N_3601,N_3673);
or U3746 (N_3746,N_3689,N_3676);
nor U3747 (N_3747,N_3630,N_3683);
nand U3748 (N_3748,N_3675,N_3626);
nand U3749 (N_3749,N_3696,N_3669);
and U3750 (N_3750,N_3660,N_3675);
nand U3751 (N_3751,N_3683,N_3676);
or U3752 (N_3752,N_3643,N_3636);
nor U3753 (N_3753,N_3692,N_3601);
or U3754 (N_3754,N_3670,N_3698);
or U3755 (N_3755,N_3604,N_3658);
nor U3756 (N_3756,N_3628,N_3658);
or U3757 (N_3757,N_3618,N_3694);
or U3758 (N_3758,N_3633,N_3630);
nand U3759 (N_3759,N_3652,N_3601);
xor U3760 (N_3760,N_3659,N_3655);
xnor U3761 (N_3761,N_3699,N_3647);
or U3762 (N_3762,N_3690,N_3677);
and U3763 (N_3763,N_3600,N_3639);
nand U3764 (N_3764,N_3646,N_3688);
nand U3765 (N_3765,N_3636,N_3648);
or U3766 (N_3766,N_3671,N_3693);
nor U3767 (N_3767,N_3698,N_3621);
nand U3768 (N_3768,N_3649,N_3680);
nor U3769 (N_3769,N_3642,N_3648);
or U3770 (N_3770,N_3627,N_3628);
and U3771 (N_3771,N_3690,N_3603);
nand U3772 (N_3772,N_3627,N_3636);
nor U3773 (N_3773,N_3663,N_3603);
or U3774 (N_3774,N_3622,N_3695);
or U3775 (N_3775,N_3603,N_3687);
or U3776 (N_3776,N_3695,N_3683);
and U3777 (N_3777,N_3663,N_3669);
nor U3778 (N_3778,N_3602,N_3601);
nand U3779 (N_3779,N_3634,N_3612);
nand U3780 (N_3780,N_3600,N_3681);
nor U3781 (N_3781,N_3605,N_3641);
xor U3782 (N_3782,N_3623,N_3672);
or U3783 (N_3783,N_3690,N_3647);
nand U3784 (N_3784,N_3613,N_3655);
and U3785 (N_3785,N_3645,N_3670);
and U3786 (N_3786,N_3633,N_3623);
and U3787 (N_3787,N_3649,N_3659);
and U3788 (N_3788,N_3642,N_3601);
nor U3789 (N_3789,N_3625,N_3624);
nor U3790 (N_3790,N_3673,N_3657);
nor U3791 (N_3791,N_3623,N_3649);
nor U3792 (N_3792,N_3645,N_3616);
or U3793 (N_3793,N_3667,N_3682);
nor U3794 (N_3794,N_3652,N_3689);
and U3795 (N_3795,N_3666,N_3644);
and U3796 (N_3796,N_3609,N_3671);
and U3797 (N_3797,N_3616,N_3682);
or U3798 (N_3798,N_3699,N_3612);
nand U3799 (N_3799,N_3623,N_3698);
or U3800 (N_3800,N_3751,N_3720);
or U3801 (N_3801,N_3737,N_3733);
xnor U3802 (N_3802,N_3748,N_3764);
or U3803 (N_3803,N_3740,N_3734);
nor U3804 (N_3804,N_3796,N_3779);
nor U3805 (N_3805,N_3707,N_3762);
nor U3806 (N_3806,N_3758,N_3787);
xnor U3807 (N_3807,N_3799,N_3708);
nand U3808 (N_3808,N_3716,N_3702);
and U3809 (N_3809,N_3760,N_3772);
and U3810 (N_3810,N_3745,N_3790);
nor U3811 (N_3811,N_3797,N_3725);
nand U3812 (N_3812,N_3715,N_3739);
nor U3813 (N_3813,N_3742,N_3718);
and U3814 (N_3814,N_3724,N_3798);
and U3815 (N_3815,N_3730,N_3775);
or U3816 (N_3816,N_3791,N_3759);
nor U3817 (N_3817,N_3756,N_3765);
nor U3818 (N_3818,N_3723,N_3738);
nand U3819 (N_3819,N_3789,N_3731);
and U3820 (N_3820,N_3719,N_3774);
nand U3821 (N_3821,N_3754,N_3729);
nand U3822 (N_3822,N_3769,N_3700);
or U3823 (N_3823,N_3744,N_3712);
or U3824 (N_3824,N_3705,N_3750);
and U3825 (N_3825,N_3757,N_3781);
nor U3826 (N_3826,N_3735,N_3721);
or U3827 (N_3827,N_3785,N_3728);
xor U3828 (N_3828,N_3755,N_3709);
or U3829 (N_3829,N_3782,N_3780);
and U3830 (N_3830,N_3793,N_3722);
nand U3831 (N_3831,N_3746,N_3726);
nand U3832 (N_3832,N_3777,N_3770);
or U3833 (N_3833,N_3703,N_3773);
xor U3834 (N_3834,N_3778,N_3783);
and U3835 (N_3835,N_3752,N_3794);
and U3836 (N_3836,N_3776,N_3714);
and U3837 (N_3837,N_3786,N_3741);
nand U3838 (N_3838,N_3767,N_3717);
nand U3839 (N_3839,N_3736,N_3788);
nor U3840 (N_3840,N_3771,N_3743);
or U3841 (N_3841,N_3768,N_3732);
nor U3842 (N_3842,N_3704,N_3747);
nand U3843 (N_3843,N_3713,N_3766);
nand U3844 (N_3844,N_3784,N_3749);
nand U3845 (N_3845,N_3706,N_3792);
nand U3846 (N_3846,N_3701,N_3753);
and U3847 (N_3847,N_3711,N_3763);
nand U3848 (N_3848,N_3795,N_3761);
nor U3849 (N_3849,N_3710,N_3727);
nor U3850 (N_3850,N_3735,N_3776);
or U3851 (N_3851,N_3701,N_3784);
and U3852 (N_3852,N_3766,N_3764);
and U3853 (N_3853,N_3778,N_3792);
nor U3854 (N_3854,N_3713,N_3743);
nor U3855 (N_3855,N_3753,N_3772);
or U3856 (N_3856,N_3790,N_3720);
nor U3857 (N_3857,N_3735,N_3709);
and U3858 (N_3858,N_3749,N_3716);
nand U3859 (N_3859,N_3751,N_3721);
xor U3860 (N_3860,N_3750,N_3773);
nor U3861 (N_3861,N_3702,N_3781);
and U3862 (N_3862,N_3725,N_3732);
nand U3863 (N_3863,N_3771,N_3711);
nor U3864 (N_3864,N_3756,N_3775);
or U3865 (N_3865,N_3759,N_3778);
and U3866 (N_3866,N_3714,N_3710);
nand U3867 (N_3867,N_3777,N_3782);
nor U3868 (N_3868,N_3714,N_3706);
nand U3869 (N_3869,N_3734,N_3724);
or U3870 (N_3870,N_3780,N_3791);
nor U3871 (N_3871,N_3738,N_3717);
and U3872 (N_3872,N_3772,N_3759);
nand U3873 (N_3873,N_3732,N_3716);
nor U3874 (N_3874,N_3713,N_3761);
or U3875 (N_3875,N_3738,N_3775);
or U3876 (N_3876,N_3770,N_3704);
nor U3877 (N_3877,N_3763,N_3722);
and U3878 (N_3878,N_3774,N_3775);
or U3879 (N_3879,N_3762,N_3795);
or U3880 (N_3880,N_3715,N_3732);
nand U3881 (N_3881,N_3798,N_3736);
and U3882 (N_3882,N_3718,N_3789);
and U3883 (N_3883,N_3779,N_3785);
xnor U3884 (N_3884,N_3763,N_3739);
nor U3885 (N_3885,N_3763,N_3784);
and U3886 (N_3886,N_3745,N_3738);
and U3887 (N_3887,N_3741,N_3750);
and U3888 (N_3888,N_3722,N_3704);
nand U3889 (N_3889,N_3776,N_3786);
nand U3890 (N_3890,N_3766,N_3799);
nand U3891 (N_3891,N_3757,N_3759);
and U3892 (N_3892,N_3767,N_3718);
nand U3893 (N_3893,N_3746,N_3749);
or U3894 (N_3894,N_3716,N_3798);
or U3895 (N_3895,N_3741,N_3755);
nor U3896 (N_3896,N_3773,N_3746);
nor U3897 (N_3897,N_3725,N_3716);
or U3898 (N_3898,N_3706,N_3739);
and U3899 (N_3899,N_3744,N_3735);
and U3900 (N_3900,N_3885,N_3842);
and U3901 (N_3901,N_3849,N_3892);
or U3902 (N_3902,N_3850,N_3840);
nand U3903 (N_3903,N_3867,N_3868);
and U3904 (N_3904,N_3855,N_3845);
nand U3905 (N_3905,N_3812,N_3835);
nor U3906 (N_3906,N_3854,N_3824);
nand U3907 (N_3907,N_3873,N_3809);
nand U3908 (N_3908,N_3884,N_3851);
and U3909 (N_3909,N_3862,N_3820);
or U3910 (N_3910,N_3804,N_3847);
xnor U3911 (N_3911,N_3801,N_3837);
nor U3912 (N_3912,N_3827,N_3870);
nand U3913 (N_3913,N_3833,N_3841);
and U3914 (N_3914,N_3880,N_3803);
nor U3915 (N_3915,N_3881,N_3856);
or U3916 (N_3916,N_3857,N_3896);
and U3917 (N_3917,N_3866,N_3836);
nand U3918 (N_3918,N_3871,N_3826);
nor U3919 (N_3919,N_3839,N_3834);
or U3920 (N_3920,N_3811,N_3898);
nor U3921 (N_3921,N_3808,N_3879);
xnor U3922 (N_3922,N_3865,N_3838);
nand U3923 (N_3923,N_3858,N_3846);
and U3924 (N_3924,N_3878,N_3806);
nand U3925 (N_3925,N_3844,N_3861);
nor U3926 (N_3926,N_3889,N_3817);
nor U3927 (N_3927,N_3831,N_3853);
nand U3928 (N_3928,N_3877,N_3815);
nor U3929 (N_3929,N_3832,N_3895);
or U3930 (N_3930,N_3882,N_3807);
and U3931 (N_3931,N_3802,N_3843);
or U3932 (N_3932,N_3848,N_3897);
xnor U3933 (N_3933,N_3859,N_3819);
or U3934 (N_3934,N_3823,N_3800);
or U3935 (N_3935,N_3822,N_3872);
nand U3936 (N_3936,N_3864,N_3891);
nor U3937 (N_3937,N_3888,N_3860);
nand U3938 (N_3938,N_3810,N_3886);
and U3939 (N_3939,N_3875,N_3814);
nand U3940 (N_3940,N_3813,N_3883);
nand U3941 (N_3941,N_3863,N_3821);
or U3942 (N_3942,N_3805,N_3887);
nor U3943 (N_3943,N_3816,N_3874);
nand U3944 (N_3944,N_3852,N_3818);
nor U3945 (N_3945,N_3890,N_3899);
xor U3946 (N_3946,N_3830,N_3893);
nor U3947 (N_3947,N_3876,N_3825);
and U3948 (N_3948,N_3869,N_3828);
or U3949 (N_3949,N_3829,N_3894);
and U3950 (N_3950,N_3816,N_3873);
nand U3951 (N_3951,N_3882,N_3827);
and U3952 (N_3952,N_3841,N_3817);
and U3953 (N_3953,N_3857,N_3880);
or U3954 (N_3954,N_3864,N_3897);
nand U3955 (N_3955,N_3810,N_3833);
nand U3956 (N_3956,N_3829,N_3846);
nand U3957 (N_3957,N_3866,N_3852);
nor U3958 (N_3958,N_3850,N_3871);
nor U3959 (N_3959,N_3820,N_3888);
and U3960 (N_3960,N_3800,N_3805);
nor U3961 (N_3961,N_3832,N_3884);
or U3962 (N_3962,N_3866,N_3845);
nor U3963 (N_3963,N_3833,N_3891);
nand U3964 (N_3964,N_3844,N_3841);
or U3965 (N_3965,N_3875,N_3885);
or U3966 (N_3966,N_3809,N_3801);
xnor U3967 (N_3967,N_3875,N_3872);
nor U3968 (N_3968,N_3878,N_3825);
nor U3969 (N_3969,N_3885,N_3832);
or U3970 (N_3970,N_3830,N_3864);
xnor U3971 (N_3971,N_3871,N_3821);
nor U3972 (N_3972,N_3802,N_3881);
nand U3973 (N_3973,N_3880,N_3866);
nand U3974 (N_3974,N_3873,N_3892);
xnor U3975 (N_3975,N_3894,N_3820);
and U3976 (N_3976,N_3885,N_3840);
or U3977 (N_3977,N_3866,N_3871);
and U3978 (N_3978,N_3862,N_3807);
and U3979 (N_3979,N_3872,N_3840);
nor U3980 (N_3980,N_3895,N_3866);
and U3981 (N_3981,N_3882,N_3813);
or U3982 (N_3982,N_3862,N_3877);
or U3983 (N_3983,N_3832,N_3891);
and U3984 (N_3984,N_3866,N_3898);
nand U3985 (N_3985,N_3841,N_3852);
nand U3986 (N_3986,N_3891,N_3812);
or U3987 (N_3987,N_3882,N_3834);
or U3988 (N_3988,N_3889,N_3844);
nand U3989 (N_3989,N_3865,N_3814);
nand U3990 (N_3990,N_3867,N_3866);
or U3991 (N_3991,N_3810,N_3809);
nand U3992 (N_3992,N_3835,N_3877);
or U3993 (N_3993,N_3869,N_3856);
and U3994 (N_3994,N_3820,N_3832);
or U3995 (N_3995,N_3859,N_3852);
nand U3996 (N_3996,N_3830,N_3852);
and U3997 (N_3997,N_3846,N_3896);
xnor U3998 (N_3998,N_3856,N_3830);
xor U3999 (N_3999,N_3846,N_3834);
nor U4000 (N_4000,N_3960,N_3953);
nand U4001 (N_4001,N_3937,N_3984);
and U4002 (N_4002,N_3916,N_3943);
or U4003 (N_4003,N_3987,N_3947);
nor U4004 (N_4004,N_3956,N_3949);
nor U4005 (N_4005,N_3931,N_3918);
and U4006 (N_4006,N_3904,N_3913);
nor U4007 (N_4007,N_3985,N_3983);
or U4008 (N_4008,N_3975,N_3974);
nand U4009 (N_4009,N_3912,N_3940);
and U4010 (N_4010,N_3934,N_3932);
xnor U4011 (N_4011,N_3998,N_3922);
nand U4012 (N_4012,N_3958,N_3991);
nand U4013 (N_4013,N_3915,N_3939);
or U4014 (N_4014,N_3973,N_3968);
nor U4015 (N_4015,N_3925,N_3923);
or U4016 (N_4016,N_3924,N_3977);
or U4017 (N_4017,N_3952,N_3957);
and U4018 (N_4018,N_3900,N_3936);
xnor U4019 (N_4019,N_3906,N_3944);
nor U4020 (N_4020,N_3962,N_3935);
nand U4021 (N_4021,N_3914,N_3971);
nor U4022 (N_4022,N_3926,N_3917);
or U4023 (N_4023,N_3948,N_3967);
nor U4024 (N_4024,N_3997,N_3963);
nor U4025 (N_4025,N_3905,N_3907);
nand U4026 (N_4026,N_3979,N_3990);
or U4027 (N_4027,N_3989,N_3982);
or U4028 (N_4028,N_3955,N_3969);
or U4029 (N_4029,N_3910,N_3978);
nor U4030 (N_4030,N_3928,N_3988);
and U4031 (N_4031,N_3938,N_3950);
nand U4032 (N_4032,N_3945,N_3995);
nor U4033 (N_4033,N_3933,N_3930);
nor U4034 (N_4034,N_3920,N_3980);
nor U4035 (N_4035,N_3965,N_3954);
and U4036 (N_4036,N_3929,N_3986);
xor U4037 (N_4037,N_3966,N_3996);
nand U4038 (N_4038,N_3901,N_3911);
and U4039 (N_4039,N_3999,N_3976);
nand U4040 (N_4040,N_3970,N_3921);
and U4041 (N_4041,N_3993,N_3908);
xor U4042 (N_4042,N_3919,N_3964);
nand U4043 (N_4043,N_3927,N_3994);
nor U4044 (N_4044,N_3902,N_3903);
nand U4045 (N_4045,N_3946,N_3959);
xor U4046 (N_4046,N_3942,N_3981);
nand U4047 (N_4047,N_3909,N_3992);
nor U4048 (N_4048,N_3972,N_3951);
nand U4049 (N_4049,N_3941,N_3961);
nor U4050 (N_4050,N_3984,N_3903);
and U4051 (N_4051,N_3961,N_3920);
and U4052 (N_4052,N_3980,N_3975);
nor U4053 (N_4053,N_3910,N_3914);
xor U4054 (N_4054,N_3952,N_3926);
nand U4055 (N_4055,N_3939,N_3955);
nor U4056 (N_4056,N_3957,N_3917);
and U4057 (N_4057,N_3960,N_3955);
nand U4058 (N_4058,N_3938,N_3953);
nand U4059 (N_4059,N_3994,N_3991);
and U4060 (N_4060,N_3905,N_3984);
or U4061 (N_4061,N_3945,N_3972);
nand U4062 (N_4062,N_3952,N_3965);
nand U4063 (N_4063,N_3933,N_3938);
or U4064 (N_4064,N_3992,N_3997);
or U4065 (N_4065,N_3955,N_3911);
nand U4066 (N_4066,N_3983,N_3921);
nor U4067 (N_4067,N_3987,N_3937);
nor U4068 (N_4068,N_3993,N_3942);
and U4069 (N_4069,N_3987,N_3970);
or U4070 (N_4070,N_3947,N_3911);
nand U4071 (N_4071,N_3905,N_3924);
nand U4072 (N_4072,N_3974,N_3963);
nand U4073 (N_4073,N_3931,N_3966);
nand U4074 (N_4074,N_3991,N_3982);
nor U4075 (N_4075,N_3961,N_3988);
or U4076 (N_4076,N_3914,N_3986);
nand U4077 (N_4077,N_3949,N_3988);
or U4078 (N_4078,N_3938,N_3925);
nor U4079 (N_4079,N_3929,N_3966);
nand U4080 (N_4080,N_3980,N_3982);
and U4081 (N_4081,N_3966,N_3926);
nor U4082 (N_4082,N_3915,N_3933);
xor U4083 (N_4083,N_3991,N_3967);
xnor U4084 (N_4084,N_3916,N_3989);
nor U4085 (N_4085,N_3958,N_3944);
or U4086 (N_4086,N_3923,N_3921);
nand U4087 (N_4087,N_3911,N_3977);
xor U4088 (N_4088,N_3979,N_3975);
nor U4089 (N_4089,N_3996,N_3949);
or U4090 (N_4090,N_3938,N_3901);
nand U4091 (N_4091,N_3966,N_3971);
nor U4092 (N_4092,N_3914,N_3977);
nor U4093 (N_4093,N_3928,N_3953);
nand U4094 (N_4094,N_3948,N_3917);
nor U4095 (N_4095,N_3949,N_3934);
nand U4096 (N_4096,N_3904,N_3912);
xor U4097 (N_4097,N_3929,N_3936);
or U4098 (N_4098,N_3910,N_3913);
nand U4099 (N_4099,N_3958,N_3908);
xor U4100 (N_4100,N_4006,N_4081);
or U4101 (N_4101,N_4091,N_4002);
xor U4102 (N_4102,N_4013,N_4057);
nand U4103 (N_4103,N_4055,N_4012);
nand U4104 (N_4104,N_4032,N_4009);
nor U4105 (N_4105,N_4028,N_4000);
or U4106 (N_4106,N_4065,N_4072);
and U4107 (N_4107,N_4097,N_4077);
nor U4108 (N_4108,N_4036,N_4025);
and U4109 (N_4109,N_4054,N_4022);
nor U4110 (N_4110,N_4047,N_4068);
nand U4111 (N_4111,N_4052,N_4043);
and U4112 (N_4112,N_4026,N_4069);
xnor U4113 (N_4113,N_4010,N_4062);
and U4114 (N_4114,N_4038,N_4041);
xor U4115 (N_4115,N_4094,N_4079);
xor U4116 (N_4116,N_4030,N_4050);
or U4117 (N_4117,N_4098,N_4086);
nand U4118 (N_4118,N_4008,N_4004);
xnor U4119 (N_4119,N_4058,N_4099);
xnor U4120 (N_4120,N_4034,N_4048);
or U4121 (N_4121,N_4024,N_4073);
nor U4122 (N_4122,N_4060,N_4020);
and U4123 (N_4123,N_4023,N_4021);
xnor U4124 (N_4124,N_4078,N_4059);
nand U4125 (N_4125,N_4033,N_4039);
or U4126 (N_4126,N_4076,N_4093);
nand U4127 (N_4127,N_4075,N_4082);
or U4128 (N_4128,N_4083,N_4087);
or U4129 (N_4129,N_4096,N_4095);
nor U4130 (N_4130,N_4070,N_4046);
or U4131 (N_4131,N_4084,N_4035);
nor U4132 (N_4132,N_4019,N_4074);
or U4133 (N_4133,N_4015,N_4017);
or U4134 (N_4134,N_4040,N_4027);
or U4135 (N_4135,N_4088,N_4056);
nor U4136 (N_4136,N_4053,N_4090);
nor U4137 (N_4137,N_4089,N_4092);
or U4138 (N_4138,N_4049,N_4066);
and U4139 (N_4139,N_4045,N_4016);
or U4140 (N_4140,N_4029,N_4080);
nand U4141 (N_4141,N_4001,N_4044);
and U4142 (N_4142,N_4064,N_4031);
and U4143 (N_4143,N_4042,N_4005);
nor U4144 (N_4144,N_4085,N_4014);
and U4145 (N_4145,N_4061,N_4007);
nand U4146 (N_4146,N_4037,N_4071);
nand U4147 (N_4147,N_4011,N_4003);
nor U4148 (N_4148,N_4051,N_4018);
or U4149 (N_4149,N_4063,N_4067);
and U4150 (N_4150,N_4062,N_4055);
nor U4151 (N_4151,N_4081,N_4062);
or U4152 (N_4152,N_4006,N_4079);
and U4153 (N_4153,N_4056,N_4081);
and U4154 (N_4154,N_4030,N_4005);
nor U4155 (N_4155,N_4022,N_4004);
nand U4156 (N_4156,N_4065,N_4053);
nor U4157 (N_4157,N_4098,N_4065);
and U4158 (N_4158,N_4050,N_4035);
xnor U4159 (N_4159,N_4084,N_4032);
nor U4160 (N_4160,N_4013,N_4055);
nor U4161 (N_4161,N_4088,N_4031);
and U4162 (N_4162,N_4071,N_4054);
and U4163 (N_4163,N_4019,N_4027);
nand U4164 (N_4164,N_4061,N_4008);
or U4165 (N_4165,N_4018,N_4044);
and U4166 (N_4166,N_4069,N_4025);
nand U4167 (N_4167,N_4038,N_4071);
and U4168 (N_4168,N_4068,N_4094);
and U4169 (N_4169,N_4019,N_4032);
nand U4170 (N_4170,N_4013,N_4069);
or U4171 (N_4171,N_4046,N_4092);
nand U4172 (N_4172,N_4053,N_4002);
or U4173 (N_4173,N_4073,N_4062);
or U4174 (N_4174,N_4013,N_4031);
and U4175 (N_4175,N_4065,N_4021);
or U4176 (N_4176,N_4089,N_4082);
nor U4177 (N_4177,N_4096,N_4023);
nor U4178 (N_4178,N_4010,N_4051);
or U4179 (N_4179,N_4097,N_4079);
nand U4180 (N_4180,N_4096,N_4039);
xor U4181 (N_4181,N_4034,N_4058);
and U4182 (N_4182,N_4048,N_4012);
nand U4183 (N_4183,N_4031,N_4025);
nor U4184 (N_4184,N_4056,N_4055);
nand U4185 (N_4185,N_4086,N_4044);
or U4186 (N_4186,N_4018,N_4030);
nand U4187 (N_4187,N_4042,N_4046);
or U4188 (N_4188,N_4074,N_4017);
and U4189 (N_4189,N_4034,N_4024);
xnor U4190 (N_4190,N_4013,N_4039);
nor U4191 (N_4191,N_4010,N_4050);
or U4192 (N_4192,N_4074,N_4094);
and U4193 (N_4193,N_4008,N_4082);
xnor U4194 (N_4194,N_4012,N_4086);
and U4195 (N_4195,N_4066,N_4089);
nor U4196 (N_4196,N_4004,N_4029);
and U4197 (N_4197,N_4003,N_4044);
and U4198 (N_4198,N_4036,N_4054);
nand U4199 (N_4199,N_4063,N_4037);
nand U4200 (N_4200,N_4187,N_4167);
xor U4201 (N_4201,N_4183,N_4171);
nor U4202 (N_4202,N_4123,N_4136);
or U4203 (N_4203,N_4151,N_4106);
nor U4204 (N_4204,N_4147,N_4111);
nor U4205 (N_4205,N_4176,N_4143);
or U4206 (N_4206,N_4197,N_4122);
nor U4207 (N_4207,N_4199,N_4163);
and U4208 (N_4208,N_4173,N_4158);
nor U4209 (N_4209,N_4149,N_4125);
or U4210 (N_4210,N_4152,N_4196);
nand U4211 (N_4211,N_4121,N_4166);
nand U4212 (N_4212,N_4115,N_4194);
nor U4213 (N_4213,N_4100,N_4112);
or U4214 (N_4214,N_4102,N_4135);
and U4215 (N_4215,N_4174,N_4138);
nand U4216 (N_4216,N_4179,N_4128);
nor U4217 (N_4217,N_4137,N_4153);
xor U4218 (N_4218,N_4127,N_4144);
and U4219 (N_4219,N_4198,N_4109);
and U4220 (N_4220,N_4103,N_4181);
nor U4221 (N_4221,N_4186,N_4157);
xor U4222 (N_4222,N_4140,N_4134);
or U4223 (N_4223,N_4120,N_4133);
xnor U4224 (N_4224,N_4178,N_4114);
nand U4225 (N_4225,N_4185,N_4105);
and U4226 (N_4226,N_4180,N_4124);
and U4227 (N_4227,N_4165,N_4156);
xnor U4228 (N_4228,N_4161,N_4191);
xor U4229 (N_4229,N_4175,N_4164);
nand U4230 (N_4230,N_4154,N_4118);
and U4231 (N_4231,N_4182,N_4110);
nand U4232 (N_4232,N_4150,N_4142);
nand U4233 (N_4233,N_4177,N_4107);
xnor U4234 (N_4234,N_4113,N_4159);
xor U4235 (N_4235,N_4108,N_4145);
and U4236 (N_4236,N_4160,N_4131);
nor U4237 (N_4237,N_4141,N_4139);
xnor U4238 (N_4238,N_4184,N_4116);
and U4239 (N_4239,N_4129,N_4190);
nand U4240 (N_4240,N_4170,N_4195);
and U4241 (N_4241,N_4188,N_4162);
or U4242 (N_4242,N_4155,N_4104);
and U4243 (N_4243,N_4192,N_4193);
nor U4244 (N_4244,N_4132,N_4172);
and U4245 (N_4245,N_4119,N_4169);
or U4246 (N_4246,N_4189,N_4148);
nor U4247 (N_4247,N_4130,N_4146);
nor U4248 (N_4248,N_4117,N_4126);
or U4249 (N_4249,N_4101,N_4168);
and U4250 (N_4250,N_4161,N_4146);
or U4251 (N_4251,N_4129,N_4151);
nor U4252 (N_4252,N_4176,N_4113);
nand U4253 (N_4253,N_4120,N_4134);
nand U4254 (N_4254,N_4126,N_4180);
nand U4255 (N_4255,N_4123,N_4141);
nor U4256 (N_4256,N_4105,N_4124);
and U4257 (N_4257,N_4135,N_4162);
xnor U4258 (N_4258,N_4131,N_4122);
or U4259 (N_4259,N_4141,N_4120);
or U4260 (N_4260,N_4142,N_4104);
and U4261 (N_4261,N_4142,N_4128);
xor U4262 (N_4262,N_4132,N_4170);
or U4263 (N_4263,N_4101,N_4110);
nor U4264 (N_4264,N_4194,N_4158);
nor U4265 (N_4265,N_4172,N_4112);
or U4266 (N_4266,N_4197,N_4192);
nor U4267 (N_4267,N_4186,N_4159);
nand U4268 (N_4268,N_4144,N_4112);
and U4269 (N_4269,N_4163,N_4117);
nor U4270 (N_4270,N_4112,N_4107);
and U4271 (N_4271,N_4126,N_4150);
xnor U4272 (N_4272,N_4122,N_4159);
nand U4273 (N_4273,N_4183,N_4162);
nor U4274 (N_4274,N_4168,N_4100);
or U4275 (N_4275,N_4140,N_4111);
nor U4276 (N_4276,N_4109,N_4107);
nor U4277 (N_4277,N_4164,N_4158);
nor U4278 (N_4278,N_4185,N_4191);
or U4279 (N_4279,N_4188,N_4134);
nand U4280 (N_4280,N_4176,N_4108);
nor U4281 (N_4281,N_4156,N_4120);
and U4282 (N_4282,N_4103,N_4183);
nand U4283 (N_4283,N_4141,N_4135);
nor U4284 (N_4284,N_4161,N_4198);
or U4285 (N_4285,N_4106,N_4135);
or U4286 (N_4286,N_4199,N_4152);
or U4287 (N_4287,N_4183,N_4119);
or U4288 (N_4288,N_4151,N_4107);
nand U4289 (N_4289,N_4176,N_4171);
or U4290 (N_4290,N_4140,N_4113);
nor U4291 (N_4291,N_4147,N_4127);
or U4292 (N_4292,N_4162,N_4198);
nor U4293 (N_4293,N_4195,N_4173);
xor U4294 (N_4294,N_4195,N_4163);
and U4295 (N_4295,N_4127,N_4138);
or U4296 (N_4296,N_4108,N_4133);
nor U4297 (N_4297,N_4156,N_4187);
or U4298 (N_4298,N_4196,N_4160);
and U4299 (N_4299,N_4106,N_4147);
nand U4300 (N_4300,N_4231,N_4264);
or U4301 (N_4301,N_4224,N_4286);
xor U4302 (N_4302,N_4217,N_4273);
and U4303 (N_4303,N_4202,N_4271);
nand U4304 (N_4304,N_4254,N_4201);
nor U4305 (N_4305,N_4268,N_4221);
nand U4306 (N_4306,N_4276,N_4256);
and U4307 (N_4307,N_4280,N_4270);
or U4308 (N_4308,N_4213,N_4265);
nor U4309 (N_4309,N_4226,N_4269);
or U4310 (N_4310,N_4262,N_4232);
nor U4311 (N_4311,N_4258,N_4242);
or U4312 (N_4312,N_4291,N_4259);
nor U4313 (N_4313,N_4284,N_4220);
or U4314 (N_4314,N_4292,N_4297);
or U4315 (N_4315,N_4206,N_4244);
or U4316 (N_4316,N_4238,N_4211);
and U4317 (N_4317,N_4229,N_4252);
nand U4318 (N_4318,N_4205,N_4293);
and U4319 (N_4319,N_4219,N_4214);
or U4320 (N_4320,N_4208,N_4239);
nor U4321 (N_4321,N_4287,N_4228);
nor U4322 (N_4322,N_4203,N_4275);
nor U4323 (N_4323,N_4204,N_4249);
nor U4324 (N_4324,N_4234,N_4263);
nand U4325 (N_4325,N_4223,N_4225);
or U4326 (N_4326,N_4285,N_4218);
nand U4327 (N_4327,N_4274,N_4243);
nor U4328 (N_4328,N_4247,N_4279);
or U4329 (N_4329,N_4235,N_4278);
nor U4330 (N_4330,N_4212,N_4215);
or U4331 (N_4331,N_4251,N_4272);
nor U4332 (N_4332,N_4248,N_4240);
nor U4333 (N_4333,N_4296,N_4289);
nor U4334 (N_4334,N_4255,N_4253);
or U4335 (N_4335,N_4294,N_4246);
or U4336 (N_4336,N_4283,N_4282);
or U4337 (N_4337,N_4245,N_4210);
nor U4338 (N_4338,N_4295,N_4236);
and U4339 (N_4339,N_4261,N_4241);
nor U4340 (N_4340,N_4209,N_4288);
and U4341 (N_4341,N_4298,N_4299);
xor U4342 (N_4342,N_4260,N_4230);
xor U4343 (N_4343,N_4233,N_4267);
xor U4344 (N_4344,N_4200,N_4216);
or U4345 (N_4345,N_4277,N_4290);
or U4346 (N_4346,N_4266,N_4237);
nand U4347 (N_4347,N_4222,N_4207);
and U4348 (N_4348,N_4227,N_4281);
and U4349 (N_4349,N_4250,N_4257);
or U4350 (N_4350,N_4200,N_4222);
and U4351 (N_4351,N_4235,N_4244);
nor U4352 (N_4352,N_4298,N_4278);
nand U4353 (N_4353,N_4266,N_4292);
or U4354 (N_4354,N_4217,N_4287);
nor U4355 (N_4355,N_4216,N_4208);
or U4356 (N_4356,N_4242,N_4297);
nor U4357 (N_4357,N_4244,N_4281);
xnor U4358 (N_4358,N_4258,N_4243);
or U4359 (N_4359,N_4261,N_4217);
and U4360 (N_4360,N_4225,N_4277);
nor U4361 (N_4361,N_4281,N_4289);
and U4362 (N_4362,N_4208,N_4251);
nor U4363 (N_4363,N_4292,N_4258);
and U4364 (N_4364,N_4231,N_4207);
and U4365 (N_4365,N_4201,N_4271);
nor U4366 (N_4366,N_4222,N_4289);
xor U4367 (N_4367,N_4233,N_4202);
nor U4368 (N_4368,N_4220,N_4227);
and U4369 (N_4369,N_4281,N_4220);
nor U4370 (N_4370,N_4208,N_4299);
and U4371 (N_4371,N_4266,N_4201);
and U4372 (N_4372,N_4282,N_4214);
nor U4373 (N_4373,N_4238,N_4221);
nor U4374 (N_4374,N_4247,N_4239);
xor U4375 (N_4375,N_4241,N_4204);
nor U4376 (N_4376,N_4237,N_4215);
nor U4377 (N_4377,N_4234,N_4299);
or U4378 (N_4378,N_4279,N_4283);
and U4379 (N_4379,N_4218,N_4229);
xor U4380 (N_4380,N_4271,N_4248);
nor U4381 (N_4381,N_4298,N_4220);
nand U4382 (N_4382,N_4241,N_4242);
and U4383 (N_4383,N_4252,N_4240);
nand U4384 (N_4384,N_4240,N_4251);
or U4385 (N_4385,N_4228,N_4273);
nand U4386 (N_4386,N_4289,N_4208);
or U4387 (N_4387,N_4238,N_4213);
nand U4388 (N_4388,N_4290,N_4292);
nor U4389 (N_4389,N_4265,N_4207);
or U4390 (N_4390,N_4240,N_4212);
nor U4391 (N_4391,N_4245,N_4212);
xor U4392 (N_4392,N_4295,N_4217);
nor U4393 (N_4393,N_4237,N_4214);
or U4394 (N_4394,N_4289,N_4223);
nand U4395 (N_4395,N_4290,N_4204);
or U4396 (N_4396,N_4286,N_4269);
or U4397 (N_4397,N_4251,N_4210);
or U4398 (N_4398,N_4273,N_4223);
or U4399 (N_4399,N_4263,N_4246);
or U4400 (N_4400,N_4346,N_4393);
or U4401 (N_4401,N_4386,N_4304);
xnor U4402 (N_4402,N_4382,N_4351);
nand U4403 (N_4403,N_4370,N_4337);
and U4404 (N_4404,N_4368,N_4363);
or U4405 (N_4405,N_4302,N_4350);
nor U4406 (N_4406,N_4389,N_4378);
or U4407 (N_4407,N_4309,N_4361);
nor U4408 (N_4408,N_4375,N_4379);
nor U4409 (N_4409,N_4301,N_4333);
or U4410 (N_4410,N_4348,N_4308);
nand U4411 (N_4411,N_4391,N_4344);
nor U4412 (N_4412,N_4399,N_4343);
nand U4413 (N_4413,N_4329,N_4377);
xor U4414 (N_4414,N_4359,N_4394);
and U4415 (N_4415,N_4387,N_4354);
or U4416 (N_4416,N_4349,N_4360);
or U4417 (N_4417,N_4385,N_4384);
and U4418 (N_4418,N_4315,N_4338);
xnor U4419 (N_4419,N_4339,N_4392);
xnor U4420 (N_4420,N_4323,N_4334);
or U4421 (N_4421,N_4380,N_4369);
and U4422 (N_4422,N_4332,N_4331);
xnor U4423 (N_4423,N_4324,N_4396);
xor U4424 (N_4424,N_4330,N_4372);
xor U4425 (N_4425,N_4327,N_4397);
nand U4426 (N_4426,N_4353,N_4347);
and U4427 (N_4427,N_4311,N_4352);
xnor U4428 (N_4428,N_4357,N_4356);
nand U4429 (N_4429,N_4367,N_4398);
and U4430 (N_4430,N_4325,N_4388);
nand U4431 (N_4431,N_4320,N_4365);
xnor U4432 (N_4432,N_4307,N_4362);
nand U4433 (N_4433,N_4316,N_4306);
or U4434 (N_4434,N_4313,N_4310);
nand U4435 (N_4435,N_4300,N_4358);
nand U4436 (N_4436,N_4381,N_4335);
nand U4437 (N_4437,N_4319,N_4374);
or U4438 (N_4438,N_4376,N_4321);
and U4439 (N_4439,N_4322,N_4366);
nand U4440 (N_4440,N_4312,N_4390);
nand U4441 (N_4441,N_4371,N_4395);
nand U4442 (N_4442,N_4336,N_4326);
xor U4443 (N_4443,N_4373,N_4340);
nor U4444 (N_4444,N_4318,N_4303);
nand U4445 (N_4445,N_4364,N_4383);
or U4446 (N_4446,N_4355,N_4317);
nand U4447 (N_4447,N_4305,N_4314);
or U4448 (N_4448,N_4341,N_4342);
nor U4449 (N_4449,N_4345,N_4328);
nor U4450 (N_4450,N_4389,N_4376);
and U4451 (N_4451,N_4338,N_4346);
nand U4452 (N_4452,N_4311,N_4372);
and U4453 (N_4453,N_4314,N_4309);
nand U4454 (N_4454,N_4304,N_4365);
nand U4455 (N_4455,N_4317,N_4329);
nor U4456 (N_4456,N_4309,N_4308);
or U4457 (N_4457,N_4346,N_4308);
nor U4458 (N_4458,N_4333,N_4347);
or U4459 (N_4459,N_4361,N_4363);
nor U4460 (N_4460,N_4363,N_4307);
or U4461 (N_4461,N_4346,N_4355);
xnor U4462 (N_4462,N_4320,N_4340);
or U4463 (N_4463,N_4353,N_4390);
or U4464 (N_4464,N_4346,N_4397);
nand U4465 (N_4465,N_4304,N_4377);
nand U4466 (N_4466,N_4376,N_4355);
nand U4467 (N_4467,N_4340,N_4388);
xor U4468 (N_4468,N_4386,N_4398);
nand U4469 (N_4469,N_4306,N_4351);
nor U4470 (N_4470,N_4333,N_4371);
nor U4471 (N_4471,N_4330,N_4338);
or U4472 (N_4472,N_4342,N_4312);
nor U4473 (N_4473,N_4310,N_4349);
and U4474 (N_4474,N_4371,N_4308);
nand U4475 (N_4475,N_4361,N_4327);
nor U4476 (N_4476,N_4376,N_4300);
and U4477 (N_4477,N_4311,N_4397);
and U4478 (N_4478,N_4399,N_4381);
nand U4479 (N_4479,N_4310,N_4384);
nand U4480 (N_4480,N_4397,N_4347);
nand U4481 (N_4481,N_4311,N_4327);
nand U4482 (N_4482,N_4363,N_4372);
or U4483 (N_4483,N_4374,N_4305);
xnor U4484 (N_4484,N_4324,N_4366);
or U4485 (N_4485,N_4371,N_4331);
or U4486 (N_4486,N_4331,N_4326);
xor U4487 (N_4487,N_4394,N_4326);
nor U4488 (N_4488,N_4372,N_4326);
nor U4489 (N_4489,N_4341,N_4329);
nand U4490 (N_4490,N_4383,N_4398);
nand U4491 (N_4491,N_4369,N_4347);
or U4492 (N_4492,N_4367,N_4336);
nand U4493 (N_4493,N_4340,N_4389);
or U4494 (N_4494,N_4319,N_4336);
nand U4495 (N_4495,N_4301,N_4362);
or U4496 (N_4496,N_4374,N_4324);
and U4497 (N_4497,N_4388,N_4347);
or U4498 (N_4498,N_4395,N_4318);
and U4499 (N_4499,N_4368,N_4329);
and U4500 (N_4500,N_4469,N_4402);
nand U4501 (N_4501,N_4472,N_4446);
or U4502 (N_4502,N_4430,N_4420);
or U4503 (N_4503,N_4476,N_4454);
nand U4504 (N_4504,N_4406,N_4428);
and U4505 (N_4505,N_4459,N_4487);
xor U4506 (N_4506,N_4473,N_4491);
and U4507 (N_4507,N_4413,N_4484);
or U4508 (N_4508,N_4404,N_4479);
or U4509 (N_4509,N_4495,N_4482);
nand U4510 (N_4510,N_4439,N_4448);
and U4511 (N_4511,N_4440,N_4494);
nor U4512 (N_4512,N_4451,N_4452);
nor U4513 (N_4513,N_4411,N_4434);
or U4514 (N_4514,N_4424,N_4471);
nor U4515 (N_4515,N_4429,N_4480);
and U4516 (N_4516,N_4435,N_4455);
or U4517 (N_4517,N_4467,N_4438);
nand U4518 (N_4518,N_4492,N_4426);
and U4519 (N_4519,N_4465,N_4407);
nor U4520 (N_4520,N_4421,N_4497);
and U4521 (N_4521,N_4450,N_4418);
and U4522 (N_4522,N_4431,N_4419);
and U4523 (N_4523,N_4457,N_4443);
or U4524 (N_4524,N_4481,N_4478);
xor U4525 (N_4525,N_4453,N_4488);
and U4526 (N_4526,N_4401,N_4475);
nor U4527 (N_4527,N_4499,N_4493);
nor U4528 (N_4528,N_4474,N_4412);
or U4529 (N_4529,N_4496,N_4403);
nor U4530 (N_4530,N_4417,N_4477);
and U4531 (N_4531,N_4415,N_4441);
or U4532 (N_4532,N_4447,N_4423);
nand U4533 (N_4533,N_4409,N_4408);
or U4534 (N_4534,N_4483,N_4422);
nand U4535 (N_4535,N_4466,N_4489);
nand U4536 (N_4536,N_4416,N_4461);
or U4537 (N_4537,N_4432,N_4414);
nand U4538 (N_4538,N_4436,N_4410);
nand U4539 (N_4539,N_4445,N_4485);
or U4540 (N_4540,N_4470,N_4490);
nor U4541 (N_4541,N_4437,N_4458);
nand U4542 (N_4542,N_4463,N_4400);
nand U4543 (N_4543,N_4486,N_4442);
and U4544 (N_4544,N_4462,N_4444);
and U4545 (N_4545,N_4498,N_4464);
nand U4546 (N_4546,N_4456,N_4433);
and U4547 (N_4547,N_4460,N_4425);
nor U4548 (N_4548,N_4405,N_4468);
and U4549 (N_4549,N_4449,N_4427);
nand U4550 (N_4550,N_4495,N_4494);
nand U4551 (N_4551,N_4479,N_4448);
and U4552 (N_4552,N_4403,N_4419);
or U4553 (N_4553,N_4441,N_4496);
and U4554 (N_4554,N_4450,N_4480);
xnor U4555 (N_4555,N_4492,N_4445);
xor U4556 (N_4556,N_4497,N_4469);
nand U4557 (N_4557,N_4424,N_4446);
or U4558 (N_4558,N_4482,N_4455);
nor U4559 (N_4559,N_4451,N_4479);
nor U4560 (N_4560,N_4470,N_4432);
nor U4561 (N_4561,N_4467,N_4419);
nand U4562 (N_4562,N_4406,N_4438);
nand U4563 (N_4563,N_4452,N_4408);
and U4564 (N_4564,N_4404,N_4424);
nor U4565 (N_4565,N_4489,N_4427);
or U4566 (N_4566,N_4454,N_4442);
nand U4567 (N_4567,N_4481,N_4456);
nor U4568 (N_4568,N_4465,N_4495);
or U4569 (N_4569,N_4481,N_4482);
nand U4570 (N_4570,N_4436,N_4480);
nand U4571 (N_4571,N_4495,N_4413);
or U4572 (N_4572,N_4466,N_4425);
and U4573 (N_4573,N_4442,N_4430);
nor U4574 (N_4574,N_4486,N_4413);
nand U4575 (N_4575,N_4423,N_4493);
nor U4576 (N_4576,N_4496,N_4421);
or U4577 (N_4577,N_4452,N_4475);
and U4578 (N_4578,N_4419,N_4413);
nor U4579 (N_4579,N_4424,N_4459);
nand U4580 (N_4580,N_4434,N_4494);
nor U4581 (N_4581,N_4418,N_4456);
and U4582 (N_4582,N_4449,N_4490);
nor U4583 (N_4583,N_4482,N_4491);
or U4584 (N_4584,N_4499,N_4407);
or U4585 (N_4585,N_4467,N_4489);
nand U4586 (N_4586,N_4443,N_4401);
nand U4587 (N_4587,N_4456,N_4492);
and U4588 (N_4588,N_4455,N_4451);
nor U4589 (N_4589,N_4401,N_4423);
and U4590 (N_4590,N_4431,N_4471);
nor U4591 (N_4591,N_4496,N_4419);
nand U4592 (N_4592,N_4441,N_4457);
or U4593 (N_4593,N_4492,N_4466);
nand U4594 (N_4594,N_4465,N_4416);
xnor U4595 (N_4595,N_4451,N_4492);
nand U4596 (N_4596,N_4441,N_4499);
nand U4597 (N_4597,N_4454,N_4448);
or U4598 (N_4598,N_4427,N_4482);
nor U4599 (N_4599,N_4497,N_4410);
nand U4600 (N_4600,N_4598,N_4550);
xor U4601 (N_4601,N_4545,N_4511);
nand U4602 (N_4602,N_4522,N_4568);
nor U4603 (N_4603,N_4529,N_4595);
nand U4604 (N_4604,N_4543,N_4584);
nor U4605 (N_4605,N_4576,N_4560);
xnor U4606 (N_4606,N_4525,N_4563);
xnor U4607 (N_4607,N_4553,N_4562);
or U4608 (N_4608,N_4585,N_4552);
or U4609 (N_4609,N_4540,N_4549);
and U4610 (N_4610,N_4532,N_4507);
nor U4611 (N_4611,N_4591,N_4593);
and U4612 (N_4612,N_4527,N_4599);
xor U4613 (N_4613,N_4567,N_4574);
xor U4614 (N_4614,N_4539,N_4537);
or U4615 (N_4615,N_4590,N_4515);
nor U4616 (N_4616,N_4514,N_4579);
nor U4617 (N_4617,N_4500,N_4534);
or U4618 (N_4618,N_4506,N_4587);
and U4619 (N_4619,N_4516,N_4573);
nand U4620 (N_4620,N_4586,N_4597);
nor U4621 (N_4621,N_4556,N_4513);
nand U4622 (N_4622,N_4581,N_4538);
and U4623 (N_4623,N_4572,N_4569);
or U4624 (N_4624,N_4501,N_4536);
xor U4625 (N_4625,N_4502,N_4588);
or U4626 (N_4626,N_4504,N_4505);
or U4627 (N_4627,N_4565,N_4548);
nor U4628 (N_4628,N_4546,N_4526);
and U4629 (N_4629,N_4530,N_4589);
or U4630 (N_4630,N_4554,N_4559);
nand U4631 (N_4631,N_4531,N_4566);
nor U4632 (N_4632,N_4503,N_4533);
xor U4633 (N_4633,N_4561,N_4523);
or U4634 (N_4634,N_4551,N_4521);
or U4635 (N_4635,N_4547,N_4582);
nand U4636 (N_4636,N_4541,N_4518);
xor U4637 (N_4637,N_4557,N_4594);
xnor U4638 (N_4638,N_4535,N_4542);
nor U4639 (N_4639,N_4580,N_4564);
nor U4640 (N_4640,N_4519,N_4520);
and U4641 (N_4641,N_4555,N_4544);
or U4642 (N_4642,N_4575,N_4578);
nor U4643 (N_4643,N_4583,N_4570);
nand U4644 (N_4644,N_4596,N_4524);
nor U4645 (N_4645,N_4517,N_4592);
and U4646 (N_4646,N_4577,N_4512);
xnor U4647 (N_4647,N_4528,N_4509);
nand U4648 (N_4648,N_4510,N_4508);
nand U4649 (N_4649,N_4558,N_4571);
and U4650 (N_4650,N_4550,N_4564);
or U4651 (N_4651,N_4555,N_4585);
nor U4652 (N_4652,N_4544,N_4554);
nor U4653 (N_4653,N_4566,N_4505);
xor U4654 (N_4654,N_4598,N_4520);
nor U4655 (N_4655,N_4533,N_4534);
nand U4656 (N_4656,N_4588,N_4524);
and U4657 (N_4657,N_4578,N_4542);
nor U4658 (N_4658,N_4518,N_4589);
nor U4659 (N_4659,N_4543,N_4555);
and U4660 (N_4660,N_4573,N_4550);
nor U4661 (N_4661,N_4582,N_4502);
and U4662 (N_4662,N_4589,N_4528);
xor U4663 (N_4663,N_4599,N_4549);
or U4664 (N_4664,N_4531,N_4568);
xor U4665 (N_4665,N_4567,N_4584);
or U4666 (N_4666,N_4512,N_4590);
nand U4667 (N_4667,N_4533,N_4558);
nand U4668 (N_4668,N_4554,N_4506);
or U4669 (N_4669,N_4510,N_4516);
nor U4670 (N_4670,N_4524,N_4531);
or U4671 (N_4671,N_4581,N_4511);
nor U4672 (N_4672,N_4594,N_4503);
nand U4673 (N_4673,N_4541,N_4588);
and U4674 (N_4674,N_4505,N_4594);
or U4675 (N_4675,N_4527,N_4563);
nor U4676 (N_4676,N_4558,N_4502);
and U4677 (N_4677,N_4547,N_4508);
nand U4678 (N_4678,N_4570,N_4543);
nor U4679 (N_4679,N_4503,N_4525);
and U4680 (N_4680,N_4534,N_4578);
nor U4681 (N_4681,N_4571,N_4570);
or U4682 (N_4682,N_4582,N_4597);
nor U4683 (N_4683,N_4527,N_4528);
and U4684 (N_4684,N_4568,N_4598);
nand U4685 (N_4685,N_4548,N_4561);
nand U4686 (N_4686,N_4513,N_4593);
nand U4687 (N_4687,N_4521,N_4537);
or U4688 (N_4688,N_4526,N_4565);
and U4689 (N_4689,N_4535,N_4578);
or U4690 (N_4690,N_4543,N_4520);
nand U4691 (N_4691,N_4547,N_4584);
and U4692 (N_4692,N_4556,N_4555);
or U4693 (N_4693,N_4506,N_4533);
nand U4694 (N_4694,N_4542,N_4559);
and U4695 (N_4695,N_4550,N_4593);
nor U4696 (N_4696,N_4546,N_4530);
nand U4697 (N_4697,N_4502,N_4547);
and U4698 (N_4698,N_4519,N_4531);
nor U4699 (N_4699,N_4533,N_4526);
nor U4700 (N_4700,N_4636,N_4684);
nor U4701 (N_4701,N_4635,N_4601);
xnor U4702 (N_4702,N_4658,N_4621);
xnor U4703 (N_4703,N_4678,N_4665);
or U4704 (N_4704,N_4602,N_4623);
or U4705 (N_4705,N_4655,N_4682);
nand U4706 (N_4706,N_4615,N_4641);
and U4707 (N_4707,N_4677,N_4680);
nand U4708 (N_4708,N_4675,N_4698);
nor U4709 (N_4709,N_4603,N_4626);
and U4710 (N_4710,N_4637,N_4673);
nand U4711 (N_4711,N_4687,N_4688);
xnor U4712 (N_4712,N_4694,N_4627);
nor U4713 (N_4713,N_4644,N_4679);
nand U4714 (N_4714,N_4681,N_4657);
and U4715 (N_4715,N_4608,N_4628);
or U4716 (N_4716,N_4653,N_4666);
or U4717 (N_4717,N_4629,N_4690);
xnor U4718 (N_4718,N_4668,N_4697);
nor U4719 (N_4719,N_4631,N_4692);
nand U4720 (N_4720,N_4607,N_4676);
nor U4721 (N_4721,N_4616,N_4620);
nor U4722 (N_4722,N_4609,N_4651);
xnor U4723 (N_4723,N_4660,N_4613);
xor U4724 (N_4724,N_4632,N_4618);
and U4725 (N_4725,N_4691,N_4634);
xor U4726 (N_4726,N_4670,N_4617);
and U4727 (N_4727,N_4664,N_4663);
nand U4728 (N_4728,N_4669,N_4689);
nor U4729 (N_4729,N_4643,N_4662);
and U4730 (N_4730,N_4696,N_4683);
nor U4731 (N_4731,N_4622,N_4647);
or U4732 (N_4732,N_4659,N_4639);
xor U4733 (N_4733,N_4610,N_4686);
and U4734 (N_4734,N_4699,N_4640);
or U4735 (N_4735,N_4638,N_4693);
nor U4736 (N_4736,N_4645,N_4612);
and U4737 (N_4737,N_4652,N_4649);
and U4738 (N_4738,N_4672,N_4633);
and U4739 (N_4739,N_4606,N_4661);
and U4740 (N_4740,N_4604,N_4619);
nand U4741 (N_4741,N_4624,N_4650);
nand U4742 (N_4742,N_4695,N_4671);
or U4743 (N_4743,N_4654,N_4667);
nor U4744 (N_4744,N_4611,N_4642);
or U4745 (N_4745,N_4614,N_4674);
nand U4746 (N_4746,N_4648,N_4625);
nor U4747 (N_4747,N_4646,N_4600);
xnor U4748 (N_4748,N_4630,N_4685);
and U4749 (N_4749,N_4605,N_4656);
nor U4750 (N_4750,N_4617,N_4692);
or U4751 (N_4751,N_4678,N_4661);
nand U4752 (N_4752,N_4694,N_4672);
nand U4753 (N_4753,N_4603,N_4664);
xor U4754 (N_4754,N_4612,N_4617);
and U4755 (N_4755,N_4690,N_4664);
or U4756 (N_4756,N_4629,N_4681);
xnor U4757 (N_4757,N_4641,N_4609);
nand U4758 (N_4758,N_4684,N_4629);
nor U4759 (N_4759,N_4687,N_4616);
nand U4760 (N_4760,N_4670,N_4693);
nor U4761 (N_4761,N_4609,N_4675);
nor U4762 (N_4762,N_4624,N_4681);
nor U4763 (N_4763,N_4693,N_4618);
nor U4764 (N_4764,N_4608,N_4603);
nand U4765 (N_4765,N_4617,N_4688);
nor U4766 (N_4766,N_4677,N_4611);
nand U4767 (N_4767,N_4623,N_4695);
nand U4768 (N_4768,N_4697,N_4616);
nand U4769 (N_4769,N_4603,N_4682);
nand U4770 (N_4770,N_4691,N_4668);
xnor U4771 (N_4771,N_4606,N_4670);
nor U4772 (N_4772,N_4619,N_4636);
or U4773 (N_4773,N_4603,N_4632);
nor U4774 (N_4774,N_4650,N_4622);
and U4775 (N_4775,N_4651,N_4683);
or U4776 (N_4776,N_4674,N_4627);
xnor U4777 (N_4777,N_4659,N_4664);
and U4778 (N_4778,N_4605,N_4652);
nand U4779 (N_4779,N_4630,N_4614);
xor U4780 (N_4780,N_4688,N_4690);
or U4781 (N_4781,N_4666,N_4626);
xnor U4782 (N_4782,N_4633,N_4629);
nand U4783 (N_4783,N_4625,N_4676);
nand U4784 (N_4784,N_4665,N_4633);
or U4785 (N_4785,N_4670,N_4625);
nor U4786 (N_4786,N_4645,N_4651);
nand U4787 (N_4787,N_4678,N_4617);
and U4788 (N_4788,N_4620,N_4641);
nand U4789 (N_4789,N_4614,N_4641);
and U4790 (N_4790,N_4696,N_4656);
or U4791 (N_4791,N_4675,N_4694);
xnor U4792 (N_4792,N_4609,N_4627);
or U4793 (N_4793,N_4634,N_4677);
nand U4794 (N_4794,N_4692,N_4620);
xnor U4795 (N_4795,N_4618,N_4601);
nor U4796 (N_4796,N_4607,N_4637);
and U4797 (N_4797,N_4600,N_4656);
or U4798 (N_4798,N_4663,N_4633);
nor U4799 (N_4799,N_4628,N_4601);
or U4800 (N_4800,N_4754,N_4772);
or U4801 (N_4801,N_4774,N_4742);
or U4802 (N_4802,N_4769,N_4767);
nand U4803 (N_4803,N_4762,N_4719);
or U4804 (N_4804,N_4779,N_4781);
nor U4805 (N_4805,N_4708,N_4747);
nor U4806 (N_4806,N_4702,N_4715);
and U4807 (N_4807,N_4763,N_4704);
and U4808 (N_4808,N_4793,N_4739);
or U4809 (N_4809,N_4780,N_4746);
nand U4810 (N_4810,N_4757,N_4741);
xnor U4811 (N_4811,N_4756,N_4731);
or U4812 (N_4812,N_4726,N_4713);
nor U4813 (N_4813,N_4786,N_4787);
and U4814 (N_4814,N_4795,N_4734);
xnor U4815 (N_4815,N_4733,N_4796);
nor U4816 (N_4816,N_4773,N_4744);
or U4817 (N_4817,N_4736,N_4760);
and U4818 (N_4818,N_4712,N_4797);
and U4819 (N_4819,N_4792,N_4706);
nand U4820 (N_4820,N_4799,N_4723);
and U4821 (N_4821,N_4791,N_4794);
or U4822 (N_4822,N_4771,N_4737);
nand U4823 (N_4823,N_4738,N_4755);
nor U4824 (N_4824,N_4710,N_4717);
nor U4825 (N_4825,N_4785,N_4750);
or U4826 (N_4826,N_4703,N_4782);
nand U4827 (N_4827,N_4718,N_4761);
nand U4828 (N_4828,N_4798,N_4721);
or U4829 (N_4829,N_4768,N_4729);
nor U4830 (N_4830,N_4728,N_4778);
and U4831 (N_4831,N_4783,N_4722);
and U4832 (N_4832,N_4735,N_4740);
nand U4833 (N_4833,N_4745,N_4789);
nor U4834 (N_4834,N_4724,N_4711);
and U4835 (N_4835,N_4749,N_4701);
nand U4836 (N_4836,N_4725,N_4752);
and U4837 (N_4837,N_4705,N_4790);
or U4838 (N_4838,N_4775,N_4759);
and U4839 (N_4839,N_4730,N_4743);
nand U4840 (N_4840,N_4788,N_4777);
or U4841 (N_4841,N_4748,N_4764);
or U4842 (N_4842,N_4770,N_4784);
and U4843 (N_4843,N_4707,N_4727);
nor U4844 (N_4844,N_4766,N_4765);
or U4845 (N_4845,N_4732,N_4751);
and U4846 (N_4846,N_4758,N_4716);
nand U4847 (N_4847,N_4753,N_4700);
or U4848 (N_4848,N_4709,N_4720);
nor U4849 (N_4849,N_4776,N_4714);
xor U4850 (N_4850,N_4716,N_4702);
or U4851 (N_4851,N_4733,N_4744);
nor U4852 (N_4852,N_4733,N_4735);
nor U4853 (N_4853,N_4794,N_4772);
or U4854 (N_4854,N_4779,N_4764);
xnor U4855 (N_4855,N_4781,N_4722);
or U4856 (N_4856,N_4719,N_4775);
and U4857 (N_4857,N_4759,N_4714);
nand U4858 (N_4858,N_4727,N_4765);
nor U4859 (N_4859,N_4775,N_4797);
or U4860 (N_4860,N_4743,N_4775);
and U4861 (N_4861,N_4711,N_4730);
and U4862 (N_4862,N_4790,N_4769);
or U4863 (N_4863,N_4742,N_4778);
or U4864 (N_4864,N_4777,N_4736);
or U4865 (N_4865,N_4762,N_4786);
nor U4866 (N_4866,N_4756,N_4701);
nor U4867 (N_4867,N_4736,N_4798);
nor U4868 (N_4868,N_4791,N_4716);
or U4869 (N_4869,N_4719,N_4763);
or U4870 (N_4870,N_4708,N_4785);
nor U4871 (N_4871,N_4798,N_4737);
nand U4872 (N_4872,N_4791,N_4704);
and U4873 (N_4873,N_4746,N_4789);
or U4874 (N_4874,N_4742,N_4757);
or U4875 (N_4875,N_4774,N_4709);
or U4876 (N_4876,N_4728,N_4717);
xor U4877 (N_4877,N_4793,N_4719);
and U4878 (N_4878,N_4737,N_4790);
nand U4879 (N_4879,N_4790,N_4782);
or U4880 (N_4880,N_4764,N_4758);
and U4881 (N_4881,N_4703,N_4754);
nor U4882 (N_4882,N_4738,N_4760);
or U4883 (N_4883,N_4781,N_4700);
and U4884 (N_4884,N_4737,N_4796);
xor U4885 (N_4885,N_4709,N_4737);
nor U4886 (N_4886,N_4712,N_4780);
nand U4887 (N_4887,N_4760,N_4722);
nor U4888 (N_4888,N_4778,N_4708);
and U4889 (N_4889,N_4795,N_4799);
nand U4890 (N_4890,N_4739,N_4729);
and U4891 (N_4891,N_4790,N_4732);
nor U4892 (N_4892,N_4718,N_4783);
nand U4893 (N_4893,N_4796,N_4743);
nor U4894 (N_4894,N_4785,N_4753);
or U4895 (N_4895,N_4795,N_4704);
and U4896 (N_4896,N_4701,N_4788);
xnor U4897 (N_4897,N_4754,N_4777);
xnor U4898 (N_4898,N_4746,N_4752);
or U4899 (N_4899,N_4714,N_4720);
nand U4900 (N_4900,N_4833,N_4841);
nor U4901 (N_4901,N_4801,N_4826);
nand U4902 (N_4902,N_4858,N_4805);
xor U4903 (N_4903,N_4851,N_4883);
nand U4904 (N_4904,N_4844,N_4806);
or U4905 (N_4905,N_4896,N_4863);
nor U4906 (N_4906,N_4840,N_4864);
and U4907 (N_4907,N_4868,N_4809);
or U4908 (N_4908,N_4859,N_4848);
and U4909 (N_4909,N_4847,N_4817);
and U4910 (N_4910,N_4865,N_4852);
nor U4911 (N_4911,N_4845,N_4846);
nor U4912 (N_4912,N_4876,N_4842);
and U4913 (N_4913,N_4814,N_4853);
nand U4914 (N_4914,N_4886,N_4836);
xnor U4915 (N_4915,N_4810,N_4870);
nor U4916 (N_4916,N_4877,N_4856);
nor U4917 (N_4917,N_4889,N_4820);
nor U4918 (N_4918,N_4831,N_4812);
xnor U4919 (N_4919,N_4861,N_4880);
nand U4920 (N_4920,N_4803,N_4871);
or U4921 (N_4921,N_4829,N_4874);
or U4922 (N_4922,N_4895,N_4894);
and U4923 (N_4923,N_4899,N_4827);
nor U4924 (N_4924,N_4811,N_4873);
and U4925 (N_4925,N_4890,N_4867);
and U4926 (N_4926,N_4825,N_4808);
or U4927 (N_4927,N_4888,N_4875);
nand U4928 (N_4928,N_4884,N_4854);
nor U4929 (N_4929,N_4893,N_4892);
or U4930 (N_4930,N_4855,N_4838);
or U4931 (N_4931,N_4866,N_4898);
and U4932 (N_4932,N_4837,N_4882);
and U4933 (N_4933,N_4872,N_4822);
and U4934 (N_4934,N_4832,N_4860);
or U4935 (N_4935,N_4897,N_4823);
nor U4936 (N_4936,N_4849,N_4891);
nand U4937 (N_4937,N_4830,N_4828);
nand U4938 (N_4938,N_4881,N_4800);
nor U4939 (N_4939,N_4887,N_4824);
and U4940 (N_4940,N_4813,N_4819);
nand U4941 (N_4941,N_4839,N_4857);
nor U4942 (N_4942,N_4850,N_4818);
xor U4943 (N_4943,N_4869,N_4834);
and U4944 (N_4944,N_4804,N_4885);
nor U4945 (N_4945,N_4802,N_4807);
and U4946 (N_4946,N_4816,N_4815);
xnor U4947 (N_4947,N_4821,N_4835);
nand U4948 (N_4948,N_4878,N_4879);
and U4949 (N_4949,N_4843,N_4862);
or U4950 (N_4950,N_4831,N_4854);
nor U4951 (N_4951,N_4880,N_4827);
xor U4952 (N_4952,N_4818,N_4806);
nor U4953 (N_4953,N_4812,N_4827);
or U4954 (N_4954,N_4836,N_4854);
or U4955 (N_4955,N_4887,N_4842);
or U4956 (N_4956,N_4870,N_4885);
xor U4957 (N_4957,N_4861,N_4801);
and U4958 (N_4958,N_4838,N_4823);
xnor U4959 (N_4959,N_4864,N_4890);
nand U4960 (N_4960,N_4821,N_4862);
nand U4961 (N_4961,N_4842,N_4827);
or U4962 (N_4962,N_4866,N_4878);
nor U4963 (N_4963,N_4804,N_4882);
and U4964 (N_4964,N_4851,N_4846);
or U4965 (N_4965,N_4870,N_4809);
or U4966 (N_4966,N_4811,N_4836);
and U4967 (N_4967,N_4802,N_4859);
xor U4968 (N_4968,N_4821,N_4848);
xor U4969 (N_4969,N_4871,N_4855);
and U4970 (N_4970,N_4840,N_4867);
nand U4971 (N_4971,N_4843,N_4895);
and U4972 (N_4972,N_4884,N_4824);
or U4973 (N_4973,N_4869,N_4804);
or U4974 (N_4974,N_4892,N_4870);
or U4975 (N_4975,N_4881,N_4837);
nand U4976 (N_4976,N_4845,N_4884);
or U4977 (N_4977,N_4891,N_4879);
xnor U4978 (N_4978,N_4864,N_4846);
nand U4979 (N_4979,N_4804,N_4815);
and U4980 (N_4980,N_4824,N_4811);
nand U4981 (N_4981,N_4839,N_4877);
nor U4982 (N_4982,N_4885,N_4822);
xor U4983 (N_4983,N_4813,N_4839);
and U4984 (N_4984,N_4819,N_4855);
nor U4985 (N_4985,N_4869,N_4813);
nand U4986 (N_4986,N_4873,N_4856);
nor U4987 (N_4987,N_4848,N_4865);
nand U4988 (N_4988,N_4843,N_4852);
nor U4989 (N_4989,N_4808,N_4841);
nor U4990 (N_4990,N_4838,N_4870);
and U4991 (N_4991,N_4835,N_4864);
or U4992 (N_4992,N_4899,N_4876);
nor U4993 (N_4993,N_4842,N_4889);
and U4994 (N_4994,N_4858,N_4812);
nor U4995 (N_4995,N_4801,N_4895);
nand U4996 (N_4996,N_4809,N_4816);
or U4997 (N_4997,N_4878,N_4873);
nand U4998 (N_4998,N_4864,N_4891);
or U4999 (N_4999,N_4843,N_4863);
or UO_0 (O_0,N_4998,N_4983);
nor UO_1 (O_1,N_4937,N_4906);
nor UO_2 (O_2,N_4965,N_4936);
and UO_3 (O_3,N_4934,N_4927);
and UO_4 (O_4,N_4943,N_4931);
and UO_5 (O_5,N_4991,N_4990);
and UO_6 (O_6,N_4969,N_4902);
nor UO_7 (O_7,N_4904,N_4984);
nor UO_8 (O_8,N_4978,N_4935);
nor UO_9 (O_9,N_4948,N_4908);
or UO_10 (O_10,N_4919,N_4954);
nor UO_11 (O_11,N_4925,N_4961);
nor UO_12 (O_12,N_4939,N_4938);
nand UO_13 (O_13,N_4945,N_4999);
or UO_14 (O_14,N_4955,N_4903);
nand UO_15 (O_15,N_4989,N_4975);
nand UO_16 (O_16,N_4952,N_4979);
nor UO_17 (O_17,N_4995,N_4950);
nor UO_18 (O_18,N_4933,N_4926);
or UO_19 (O_19,N_4977,N_4900);
and UO_20 (O_20,N_4930,N_4996);
or UO_21 (O_21,N_4959,N_4992);
nor UO_22 (O_22,N_4973,N_4957);
nand UO_23 (O_23,N_4923,N_4953);
or UO_24 (O_24,N_4918,N_4905);
or UO_25 (O_25,N_4994,N_4976);
nand UO_26 (O_26,N_4942,N_4951);
xnor UO_27 (O_27,N_4949,N_4916);
xor UO_28 (O_28,N_4972,N_4928);
and UO_29 (O_29,N_4929,N_4914);
or UO_30 (O_30,N_4956,N_4963);
and UO_31 (O_31,N_4966,N_4947);
nor UO_32 (O_32,N_4987,N_4981);
nor UO_33 (O_33,N_4967,N_4985);
or UO_34 (O_34,N_4960,N_4940);
nand UO_35 (O_35,N_4910,N_4974);
and UO_36 (O_36,N_4907,N_4911);
xor UO_37 (O_37,N_4982,N_4932);
nor UO_38 (O_38,N_4993,N_4920);
nor UO_39 (O_39,N_4922,N_4962);
xnor UO_40 (O_40,N_4968,N_4970);
nor UO_41 (O_41,N_4980,N_4944);
or UO_42 (O_42,N_4913,N_4997);
nand UO_43 (O_43,N_4986,N_4909);
nor UO_44 (O_44,N_4912,N_4901);
xnor UO_45 (O_45,N_4964,N_4924);
nand UO_46 (O_46,N_4958,N_4915);
and UO_47 (O_47,N_4917,N_4946);
nor UO_48 (O_48,N_4988,N_4971);
or UO_49 (O_49,N_4941,N_4921);
xor UO_50 (O_50,N_4976,N_4984);
or UO_51 (O_51,N_4974,N_4992);
nor UO_52 (O_52,N_4944,N_4917);
nand UO_53 (O_53,N_4961,N_4993);
nand UO_54 (O_54,N_4941,N_4923);
and UO_55 (O_55,N_4960,N_4929);
and UO_56 (O_56,N_4991,N_4913);
nor UO_57 (O_57,N_4913,N_4998);
nor UO_58 (O_58,N_4997,N_4959);
and UO_59 (O_59,N_4968,N_4928);
and UO_60 (O_60,N_4924,N_4992);
nand UO_61 (O_61,N_4999,N_4956);
nor UO_62 (O_62,N_4911,N_4974);
or UO_63 (O_63,N_4937,N_4933);
or UO_64 (O_64,N_4981,N_4974);
or UO_65 (O_65,N_4986,N_4972);
or UO_66 (O_66,N_4900,N_4970);
nand UO_67 (O_67,N_4964,N_4933);
nand UO_68 (O_68,N_4936,N_4905);
nand UO_69 (O_69,N_4982,N_4950);
nor UO_70 (O_70,N_4931,N_4977);
or UO_71 (O_71,N_4940,N_4926);
nor UO_72 (O_72,N_4902,N_4919);
and UO_73 (O_73,N_4911,N_4986);
nand UO_74 (O_74,N_4940,N_4931);
nor UO_75 (O_75,N_4984,N_4913);
nand UO_76 (O_76,N_4970,N_4955);
nand UO_77 (O_77,N_4940,N_4949);
or UO_78 (O_78,N_4973,N_4997);
and UO_79 (O_79,N_4987,N_4933);
nor UO_80 (O_80,N_4960,N_4921);
or UO_81 (O_81,N_4927,N_4965);
nor UO_82 (O_82,N_4995,N_4901);
or UO_83 (O_83,N_4966,N_4926);
or UO_84 (O_84,N_4938,N_4996);
or UO_85 (O_85,N_4937,N_4919);
or UO_86 (O_86,N_4997,N_4983);
nand UO_87 (O_87,N_4994,N_4940);
nor UO_88 (O_88,N_4999,N_4921);
nor UO_89 (O_89,N_4904,N_4987);
nor UO_90 (O_90,N_4978,N_4908);
and UO_91 (O_91,N_4961,N_4945);
nand UO_92 (O_92,N_4925,N_4970);
nor UO_93 (O_93,N_4917,N_4977);
xnor UO_94 (O_94,N_4928,N_4951);
nand UO_95 (O_95,N_4905,N_4978);
nor UO_96 (O_96,N_4972,N_4938);
nor UO_97 (O_97,N_4910,N_4934);
or UO_98 (O_98,N_4948,N_4964);
and UO_99 (O_99,N_4910,N_4998);
nand UO_100 (O_100,N_4903,N_4933);
and UO_101 (O_101,N_4984,N_4903);
nand UO_102 (O_102,N_4970,N_4996);
or UO_103 (O_103,N_4961,N_4997);
and UO_104 (O_104,N_4932,N_4959);
nor UO_105 (O_105,N_4961,N_4990);
and UO_106 (O_106,N_4996,N_4916);
or UO_107 (O_107,N_4974,N_4959);
nor UO_108 (O_108,N_4956,N_4981);
and UO_109 (O_109,N_4974,N_4920);
or UO_110 (O_110,N_4985,N_4994);
or UO_111 (O_111,N_4963,N_4925);
and UO_112 (O_112,N_4904,N_4969);
nor UO_113 (O_113,N_4951,N_4998);
and UO_114 (O_114,N_4943,N_4958);
xnor UO_115 (O_115,N_4965,N_4903);
nor UO_116 (O_116,N_4943,N_4947);
and UO_117 (O_117,N_4984,N_4991);
and UO_118 (O_118,N_4936,N_4970);
nor UO_119 (O_119,N_4925,N_4910);
xor UO_120 (O_120,N_4956,N_4953);
nor UO_121 (O_121,N_4945,N_4955);
and UO_122 (O_122,N_4944,N_4955);
or UO_123 (O_123,N_4991,N_4976);
and UO_124 (O_124,N_4945,N_4925);
nor UO_125 (O_125,N_4987,N_4994);
nand UO_126 (O_126,N_4958,N_4993);
and UO_127 (O_127,N_4973,N_4924);
nand UO_128 (O_128,N_4919,N_4927);
nor UO_129 (O_129,N_4962,N_4905);
or UO_130 (O_130,N_4974,N_4998);
nand UO_131 (O_131,N_4991,N_4988);
nor UO_132 (O_132,N_4976,N_4922);
nor UO_133 (O_133,N_4999,N_4972);
xor UO_134 (O_134,N_4981,N_4942);
or UO_135 (O_135,N_4937,N_4904);
nand UO_136 (O_136,N_4981,N_4920);
nor UO_137 (O_137,N_4948,N_4921);
nor UO_138 (O_138,N_4986,N_4961);
nand UO_139 (O_139,N_4962,N_4984);
or UO_140 (O_140,N_4979,N_4949);
nand UO_141 (O_141,N_4936,N_4955);
nand UO_142 (O_142,N_4959,N_4990);
and UO_143 (O_143,N_4987,N_4926);
or UO_144 (O_144,N_4976,N_4924);
nand UO_145 (O_145,N_4995,N_4999);
and UO_146 (O_146,N_4908,N_4939);
nand UO_147 (O_147,N_4914,N_4948);
xor UO_148 (O_148,N_4986,N_4904);
nor UO_149 (O_149,N_4923,N_4927);
xor UO_150 (O_150,N_4993,N_4995);
and UO_151 (O_151,N_4963,N_4955);
and UO_152 (O_152,N_4971,N_4977);
or UO_153 (O_153,N_4966,N_4955);
nand UO_154 (O_154,N_4976,N_4919);
nand UO_155 (O_155,N_4902,N_4930);
nor UO_156 (O_156,N_4959,N_4986);
and UO_157 (O_157,N_4911,N_4938);
nor UO_158 (O_158,N_4922,N_4939);
or UO_159 (O_159,N_4983,N_4996);
or UO_160 (O_160,N_4904,N_4993);
nand UO_161 (O_161,N_4985,N_4941);
and UO_162 (O_162,N_4970,N_4922);
xor UO_163 (O_163,N_4916,N_4951);
and UO_164 (O_164,N_4905,N_4954);
nand UO_165 (O_165,N_4971,N_4945);
xor UO_166 (O_166,N_4971,N_4964);
nor UO_167 (O_167,N_4960,N_4991);
and UO_168 (O_168,N_4956,N_4917);
and UO_169 (O_169,N_4991,N_4940);
nor UO_170 (O_170,N_4922,N_4961);
nand UO_171 (O_171,N_4975,N_4957);
and UO_172 (O_172,N_4922,N_4910);
xor UO_173 (O_173,N_4979,N_4919);
and UO_174 (O_174,N_4926,N_4919);
or UO_175 (O_175,N_4907,N_4988);
or UO_176 (O_176,N_4922,N_4955);
or UO_177 (O_177,N_4935,N_4902);
nand UO_178 (O_178,N_4935,N_4932);
or UO_179 (O_179,N_4940,N_4963);
and UO_180 (O_180,N_4979,N_4962);
and UO_181 (O_181,N_4919,N_4994);
nor UO_182 (O_182,N_4946,N_4905);
or UO_183 (O_183,N_4977,N_4925);
nand UO_184 (O_184,N_4986,N_4976);
nand UO_185 (O_185,N_4990,N_4946);
nor UO_186 (O_186,N_4966,N_4935);
and UO_187 (O_187,N_4907,N_4903);
nand UO_188 (O_188,N_4989,N_4945);
nand UO_189 (O_189,N_4978,N_4973);
nand UO_190 (O_190,N_4996,N_4953);
or UO_191 (O_191,N_4971,N_4917);
nand UO_192 (O_192,N_4909,N_4903);
or UO_193 (O_193,N_4958,N_4969);
nor UO_194 (O_194,N_4981,N_4900);
xnor UO_195 (O_195,N_4923,N_4966);
xnor UO_196 (O_196,N_4986,N_4932);
nor UO_197 (O_197,N_4977,N_4995);
nor UO_198 (O_198,N_4990,N_4938);
nor UO_199 (O_199,N_4998,N_4923);
xnor UO_200 (O_200,N_4908,N_4965);
nand UO_201 (O_201,N_4902,N_4991);
or UO_202 (O_202,N_4984,N_4987);
and UO_203 (O_203,N_4956,N_4941);
or UO_204 (O_204,N_4925,N_4999);
and UO_205 (O_205,N_4962,N_4990);
nor UO_206 (O_206,N_4981,N_4934);
nor UO_207 (O_207,N_4988,N_4993);
xnor UO_208 (O_208,N_4993,N_4966);
nor UO_209 (O_209,N_4951,N_4903);
and UO_210 (O_210,N_4985,N_4966);
xor UO_211 (O_211,N_4919,N_4971);
nand UO_212 (O_212,N_4921,N_4986);
or UO_213 (O_213,N_4924,N_4917);
nand UO_214 (O_214,N_4907,N_4967);
and UO_215 (O_215,N_4928,N_4924);
nand UO_216 (O_216,N_4979,N_4960);
and UO_217 (O_217,N_4953,N_4932);
xnor UO_218 (O_218,N_4907,N_4957);
or UO_219 (O_219,N_4931,N_4982);
or UO_220 (O_220,N_4968,N_4955);
nor UO_221 (O_221,N_4975,N_4972);
nand UO_222 (O_222,N_4953,N_4942);
and UO_223 (O_223,N_4917,N_4975);
xor UO_224 (O_224,N_4978,N_4979);
nor UO_225 (O_225,N_4981,N_4949);
nor UO_226 (O_226,N_4931,N_4998);
nor UO_227 (O_227,N_4909,N_4908);
or UO_228 (O_228,N_4901,N_4970);
or UO_229 (O_229,N_4912,N_4902);
nor UO_230 (O_230,N_4931,N_4905);
or UO_231 (O_231,N_4974,N_4918);
nand UO_232 (O_232,N_4917,N_4916);
nand UO_233 (O_233,N_4916,N_4978);
nor UO_234 (O_234,N_4912,N_4979);
xnor UO_235 (O_235,N_4992,N_4930);
and UO_236 (O_236,N_4950,N_4937);
nand UO_237 (O_237,N_4979,N_4928);
or UO_238 (O_238,N_4937,N_4922);
nor UO_239 (O_239,N_4975,N_4905);
or UO_240 (O_240,N_4931,N_4976);
or UO_241 (O_241,N_4983,N_4927);
and UO_242 (O_242,N_4935,N_4972);
nor UO_243 (O_243,N_4974,N_4939);
nor UO_244 (O_244,N_4989,N_4938);
or UO_245 (O_245,N_4984,N_4945);
nor UO_246 (O_246,N_4985,N_4927);
or UO_247 (O_247,N_4933,N_4945);
and UO_248 (O_248,N_4991,N_4972);
and UO_249 (O_249,N_4932,N_4945);
nor UO_250 (O_250,N_4955,N_4991);
nand UO_251 (O_251,N_4963,N_4958);
and UO_252 (O_252,N_4966,N_4959);
nand UO_253 (O_253,N_4925,N_4901);
nand UO_254 (O_254,N_4936,N_4933);
xnor UO_255 (O_255,N_4945,N_4969);
nor UO_256 (O_256,N_4989,N_4931);
nand UO_257 (O_257,N_4902,N_4970);
nor UO_258 (O_258,N_4911,N_4985);
nor UO_259 (O_259,N_4925,N_4959);
xor UO_260 (O_260,N_4991,N_4982);
and UO_261 (O_261,N_4913,N_4976);
or UO_262 (O_262,N_4996,N_4990);
nand UO_263 (O_263,N_4919,N_4955);
and UO_264 (O_264,N_4916,N_4968);
or UO_265 (O_265,N_4999,N_4988);
nor UO_266 (O_266,N_4933,N_4910);
nor UO_267 (O_267,N_4943,N_4915);
or UO_268 (O_268,N_4902,N_4956);
or UO_269 (O_269,N_4940,N_4993);
or UO_270 (O_270,N_4955,N_4908);
and UO_271 (O_271,N_4913,N_4999);
and UO_272 (O_272,N_4917,N_4970);
xor UO_273 (O_273,N_4958,N_4996);
or UO_274 (O_274,N_4982,N_4967);
xor UO_275 (O_275,N_4958,N_4961);
nor UO_276 (O_276,N_4901,N_4949);
or UO_277 (O_277,N_4998,N_4902);
and UO_278 (O_278,N_4956,N_4934);
nand UO_279 (O_279,N_4980,N_4914);
and UO_280 (O_280,N_4966,N_4995);
or UO_281 (O_281,N_4953,N_4998);
and UO_282 (O_282,N_4951,N_4926);
nor UO_283 (O_283,N_4959,N_4930);
or UO_284 (O_284,N_4930,N_4974);
nand UO_285 (O_285,N_4971,N_4934);
nor UO_286 (O_286,N_4945,N_4993);
or UO_287 (O_287,N_4997,N_4933);
nor UO_288 (O_288,N_4929,N_4996);
nand UO_289 (O_289,N_4965,N_4955);
nor UO_290 (O_290,N_4973,N_4965);
or UO_291 (O_291,N_4934,N_4953);
or UO_292 (O_292,N_4965,N_4932);
or UO_293 (O_293,N_4992,N_4966);
nor UO_294 (O_294,N_4901,N_4961);
and UO_295 (O_295,N_4956,N_4976);
nand UO_296 (O_296,N_4987,N_4976);
xnor UO_297 (O_297,N_4948,N_4943);
nand UO_298 (O_298,N_4929,N_4970);
or UO_299 (O_299,N_4993,N_4921);
nor UO_300 (O_300,N_4924,N_4987);
nor UO_301 (O_301,N_4928,N_4985);
or UO_302 (O_302,N_4933,N_4990);
nor UO_303 (O_303,N_4931,N_4957);
and UO_304 (O_304,N_4935,N_4947);
nand UO_305 (O_305,N_4990,N_4923);
and UO_306 (O_306,N_4985,N_4945);
nor UO_307 (O_307,N_4927,N_4962);
nor UO_308 (O_308,N_4951,N_4924);
or UO_309 (O_309,N_4975,N_4962);
nor UO_310 (O_310,N_4961,N_4902);
nor UO_311 (O_311,N_4972,N_4953);
nand UO_312 (O_312,N_4986,N_4990);
and UO_313 (O_313,N_4920,N_4954);
nor UO_314 (O_314,N_4952,N_4981);
nand UO_315 (O_315,N_4953,N_4940);
nor UO_316 (O_316,N_4949,N_4936);
xor UO_317 (O_317,N_4915,N_4983);
nand UO_318 (O_318,N_4972,N_4930);
and UO_319 (O_319,N_4981,N_4908);
nor UO_320 (O_320,N_4936,N_4915);
nand UO_321 (O_321,N_4909,N_4919);
xor UO_322 (O_322,N_4914,N_4996);
nand UO_323 (O_323,N_4929,N_4930);
nor UO_324 (O_324,N_4955,N_4933);
nand UO_325 (O_325,N_4941,N_4978);
and UO_326 (O_326,N_4974,N_4987);
nand UO_327 (O_327,N_4953,N_4904);
or UO_328 (O_328,N_4963,N_4993);
nor UO_329 (O_329,N_4919,N_4993);
xor UO_330 (O_330,N_4938,N_4940);
nor UO_331 (O_331,N_4973,N_4910);
and UO_332 (O_332,N_4976,N_4977);
or UO_333 (O_333,N_4968,N_4988);
nand UO_334 (O_334,N_4989,N_4963);
and UO_335 (O_335,N_4978,N_4948);
xnor UO_336 (O_336,N_4963,N_4922);
or UO_337 (O_337,N_4930,N_4900);
nor UO_338 (O_338,N_4989,N_4920);
nand UO_339 (O_339,N_4995,N_4947);
nand UO_340 (O_340,N_4932,N_4921);
and UO_341 (O_341,N_4999,N_4976);
or UO_342 (O_342,N_4960,N_4928);
and UO_343 (O_343,N_4950,N_4939);
and UO_344 (O_344,N_4976,N_4914);
or UO_345 (O_345,N_4966,N_4969);
and UO_346 (O_346,N_4993,N_4934);
xor UO_347 (O_347,N_4974,N_4912);
nor UO_348 (O_348,N_4951,N_4947);
nand UO_349 (O_349,N_4928,N_4999);
xor UO_350 (O_350,N_4957,N_4948);
or UO_351 (O_351,N_4990,N_4985);
or UO_352 (O_352,N_4903,N_4975);
or UO_353 (O_353,N_4975,N_4941);
and UO_354 (O_354,N_4917,N_4981);
xnor UO_355 (O_355,N_4918,N_4962);
xor UO_356 (O_356,N_4999,N_4979);
or UO_357 (O_357,N_4911,N_4961);
nand UO_358 (O_358,N_4966,N_4932);
or UO_359 (O_359,N_4925,N_4966);
or UO_360 (O_360,N_4988,N_4939);
and UO_361 (O_361,N_4985,N_4937);
and UO_362 (O_362,N_4925,N_4920);
nand UO_363 (O_363,N_4999,N_4914);
or UO_364 (O_364,N_4936,N_4987);
or UO_365 (O_365,N_4913,N_4952);
and UO_366 (O_366,N_4910,N_4941);
or UO_367 (O_367,N_4966,N_4904);
or UO_368 (O_368,N_4908,N_4996);
xor UO_369 (O_369,N_4948,N_4956);
or UO_370 (O_370,N_4903,N_4972);
and UO_371 (O_371,N_4926,N_4949);
nand UO_372 (O_372,N_4952,N_4928);
and UO_373 (O_373,N_4921,N_4951);
nand UO_374 (O_374,N_4905,N_4912);
nor UO_375 (O_375,N_4990,N_4998);
nand UO_376 (O_376,N_4952,N_4972);
and UO_377 (O_377,N_4923,N_4974);
nor UO_378 (O_378,N_4975,N_4993);
and UO_379 (O_379,N_4988,N_4926);
and UO_380 (O_380,N_4907,N_4963);
or UO_381 (O_381,N_4929,N_4984);
nand UO_382 (O_382,N_4966,N_4972);
or UO_383 (O_383,N_4908,N_4928);
and UO_384 (O_384,N_4944,N_4971);
and UO_385 (O_385,N_4961,N_4938);
nor UO_386 (O_386,N_4954,N_4985);
nand UO_387 (O_387,N_4928,N_4917);
and UO_388 (O_388,N_4964,N_4956);
and UO_389 (O_389,N_4931,N_4929);
nor UO_390 (O_390,N_4914,N_4952);
and UO_391 (O_391,N_4949,N_4955);
xor UO_392 (O_392,N_4997,N_4939);
nand UO_393 (O_393,N_4923,N_4938);
nand UO_394 (O_394,N_4951,N_4965);
nand UO_395 (O_395,N_4937,N_4924);
nand UO_396 (O_396,N_4978,N_4984);
nor UO_397 (O_397,N_4903,N_4915);
and UO_398 (O_398,N_4915,N_4941);
nor UO_399 (O_399,N_4981,N_4967);
or UO_400 (O_400,N_4972,N_4932);
nor UO_401 (O_401,N_4937,N_4963);
nor UO_402 (O_402,N_4908,N_4984);
nand UO_403 (O_403,N_4962,N_4911);
nor UO_404 (O_404,N_4936,N_4929);
nor UO_405 (O_405,N_4976,N_4953);
nand UO_406 (O_406,N_4943,N_4976);
nor UO_407 (O_407,N_4967,N_4921);
and UO_408 (O_408,N_4933,N_4906);
nand UO_409 (O_409,N_4949,N_4956);
and UO_410 (O_410,N_4968,N_4948);
or UO_411 (O_411,N_4985,N_4958);
and UO_412 (O_412,N_4957,N_4974);
and UO_413 (O_413,N_4901,N_4989);
nand UO_414 (O_414,N_4965,N_4979);
and UO_415 (O_415,N_4914,N_4967);
nand UO_416 (O_416,N_4999,N_4949);
nand UO_417 (O_417,N_4996,N_4975);
and UO_418 (O_418,N_4934,N_4975);
nor UO_419 (O_419,N_4910,N_4985);
nor UO_420 (O_420,N_4943,N_4936);
nor UO_421 (O_421,N_4966,N_4996);
nor UO_422 (O_422,N_4927,N_4911);
nand UO_423 (O_423,N_4915,N_4963);
or UO_424 (O_424,N_4983,N_4988);
xnor UO_425 (O_425,N_4987,N_4991);
and UO_426 (O_426,N_4999,N_4982);
or UO_427 (O_427,N_4906,N_4940);
nor UO_428 (O_428,N_4957,N_4939);
nand UO_429 (O_429,N_4920,N_4987);
and UO_430 (O_430,N_4988,N_4918);
or UO_431 (O_431,N_4901,N_4917);
or UO_432 (O_432,N_4924,N_4977);
xnor UO_433 (O_433,N_4966,N_4973);
and UO_434 (O_434,N_4936,N_4939);
xor UO_435 (O_435,N_4942,N_4900);
and UO_436 (O_436,N_4908,N_4954);
or UO_437 (O_437,N_4912,N_4977);
nand UO_438 (O_438,N_4984,N_4924);
and UO_439 (O_439,N_4902,N_4907);
xor UO_440 (O_440,N_4955,N_4900);
and UO_441 (O_441,N_4994,N_4944);
and UO_442 (O_442,N_4932,N_4997);
or UO_443 (O_443,N_4987,N_4971);
nand UO_444 (O_444,N_4917,N_4943);
and UO_445 (O_445,N_4948,N_4972);
nor UO_446 (O_446,N_4961,N_4963);
nor UO_447 (O_447,N_4943,N_4945);
nand UO_448 (O_448,N_4941,N_4962);
nand UO_449 (O_449,N_4935,N_4989);
and UO_450 (O_450,N_4906,N_4975);
xnor UO_451 (O_451,N_4986,N_4927);
nand UO_452 (O_452,N_4935,N_4998);
nand UO_453 (O_453,N_4978,N_4983);
nand UO_454 (O_454,N_4959,N_4924);
and UO_455 (O_455,N_4912,N_4949);
nor UO_456 (O_456,N_4978,N_4975);
nand UO_457 (O_457,N_4970,N_4956);
nand UO_458 (O_458,N_4948,N_4970);
nand UO_459 (O_459,N_4914,N_4964);
xor UO_460 (O_460,N_4983,N_4973);
nand UO_461 (O_461,N_4960,N_4908);
nor UO_462 (O_462,N_4903,N_4999);
and UO_463 (O_463,N_4905,N_4952);
or UO_464 (O_464,N_4929,N_4994);
xnor UO_465 (O_465,N_4931,N_4939);
nand UO_466 (O_466,N_4916,N_4954);
nor UO_467 (O_467,N_4943,N_4973);
nand UO_468 (O_468,N_4990,N_4992);
or UO_469 (O_469,N_4914,N_4931);
or UO_470 (O_470,N_4998,N_4925);
nor UO_471 (O_471,N_4915,N_4949);
nand UO_472 (O_472,N_4962,N_4997);
or UO_473 (O_473,N_4945,N_4975);
xor UO_474 (O_474,N_4919,N_4961);
or UO_475 (O_475,N_4925,N_4996);
xor UO_476 (O_476,N_4900,N_4921);
or UO_477 (O_477,N_4937,N_4968);
or UO_478 (O_478,N_4963,N_4904);
and UO_479 (O_479,N_4907,N_4986);
nor UO_480 (O_480,N_4953,N_4926);
nand UO_481 (O_481,N_4964,N_4992);
xor UO_482 (O_482,N_4984,N_4958);
nor UO_483 (O_483,N_4914,N_4900);
nand UO_484 (O_484,N_4967,N_4959);
xor UO_485 (O_485,N_4913,N_4963);
nor UO_486 (O_486,N_4924,N_4914);
and UO_487 (O_487,N_4942,N_4959);
nand UO_488 (O_488,N_4952,N_4937);
or UO_489 (O_489,N_4992,N_4978);
or UO_490 (O_490,N_4939,N_4951);
or UO_491 (O_491,N_4984,N_4909);
nand UO_492 (O_492,N_4930,N_4984);
nor UO_493 (O_493,N_4937,N_4934);
and UO_494 (O_494,N_4906,N_4972);
and UO_495 (O_495,N_4926,N_4955);
nor UO_496 (O_496,N_4981,N_4954);
nor UO_497 (O_497,N_4938,N_4985);
nand UO_498 (O_498,N_4941,N_4926);
or UO_499 (O_499,N_4983,N_4908);
or UO_500 (O_500,N_4924,N_4966);
nor UO_501 (O_501,N_4913,N_4917);
nand UO_502 (O_502,N_4987,N_4942);
xnor UO_503 (O_503,N_4950,N_4928);
or UO_504 (O_504,N_4909,N_4948);
xnor UO_505 (O_505,N_4921,N_4979);
nand UO_506 (O_506,N_4942,N_4920);
nand UO_507 (O_507,N_4979,N_4976);
nand UO_508 (O_508,N_4974,N_4900);
nor UO_509 (O_509,N_4907,N_4964);
xnor UO_510 (O_510,N_4901,N_4930);
or UO_511 (O_511,N_4999,N_4955);
and UO_512 (O_512,N_4938,N_4931);
nand UO_513 (O_513,N_4909,N_4912);
nand UO_514 (O_514,N_4978,N_4993);
nand UO_515 (O_515,N_4923,N_4930);
and UO_516 (O_516,N_4934,N_4925);
and UO_517 (O_517,N_4901,N_4964);
or UO_518 (O_518,N_4936,N_4914);
nor UO_519 (O_519,N_4936,N_4902);
nand UO_520 (O_520,N_4954,N_4953);
and UO_521 (O_521,N_4993,N_4953);
and UO_522 (O_522,N_4990,N_4970);
or UO_523 (O_523,N_4957,N_4924);
xnor UO_524 (O_524,N_4949,N_4911);
nand UO_525 (O_525,N_4988,N_4930);
xor UO_526 (O_526,N_4992,N_4985);
or UO_527 (O_527,N_4945,N_4924);
or UO_528 (O_528,N_4943,N_4995);
and UO_529 (O_529,N_4987,N_4985);
and UO_530 (O_530,N_4913,N_4910);
and UO_531 (O_531,N_4947,N_4925);
and UO_532 (O_532,N_4957,N_4920);
or UO_533 (O_533,N_4963,N_4923);
nor UO_534 (O_534,N_4929,N_4998);
nand UO_535 (O_535,N_4958,N_4926);
nor UO_536 (O_536,N_4978,N_4929);
or UO_537 (O_537,N_4965,N_4975);
or UO_538 (O_538,N_4908,N_4963);
or UO_539 (O_539,N_4920,N_4973);
xor UO_540 (O_540,N_4912,N_4955);
nor UO_541 (O_541,N_4917,N_4980);
or UO_542 (O_542,N_4999,N_4924);
nor UO_543 (O_543,N_4990,N_4948);
nor UO_544 (O_544,N_4986,N_4974);
and UO_545 (O_545,N_4904,N_4978);
xnor UO_546 (O_546,N_4953,N_4984);
xor UO_547 (O_547,N_4941,N_4991);
and UO_548 (O_548,N_4995,N_4926);
xnor UO_549 (O_549,N_4901,N_4938);
nor UO_550 (O_550,N_4992,N_4941);
or UO_551 (O_551,N_4973,N_4969);
xnor UO_552 (O_552,N_4911,N_4934);
nor UO_553 (O_553,N_4966,N_4906);
and UO_554 (O_554,N_4946,N_4944);
nand UO_555 (O_555,N_4961,N_4924);
nand UO_556 (O_556,N_4989,N_4900);
or UO_557 (O_557,N_4909,N_4915);
or UO_558 (O_558,N_4978,N_4971);
or UO_559 (O_559,N_4907,N_4927);
nor UO_560 (O_560,N_4967,N_4918);
and UO_561 (O_561,N_4907,N_4978);
nand UO_562 (O_562,N_4942,N_4918);
and UO_563 (O_563,N_4943,N_4994);
nor UO_564 (O_564,N_4942,N_4923);
nand UO_565 (O_565,N_4939,N_4944);
xor UO_566 (O_566,N_4986,N_4917);
nor UO_567 (O_567,N_4983,N_4974);
nor UO_568 (O_568,N_4996,N_4982);
xor UO_569 (O_569,N_4964,N_4966);
nand UO_570 (O_570,N_4901,N_4998);
and UO_571 (O_571,N_4922,N_4959);
nor UO_572 (O_572,N_4971,N_4940);
nand UO_573 (O_573,N_4911,N_4983);
nand UO_574 (O_574,N_4907,N_4918);
nand UO_575 (O_575,N_4991,N_4927);
and UO_576 (O_576,N_4955,N_4996);
nand UO_577 (O_577,N_4957,N_4989);
nand UO_578 (O_578,N_4977,N_4909);
nor UO_579 (O_579,N_4970,N_4966);
xor UO_580 (O_580,N_4939,N_4955);
or UO_581 (O_581,N_4950,N_4998);
nand UO_582 (O_582,N_4916,N_4943);
nand UO_583 (O_583,N_4900,N_4937);
nand UO_584 (O_584,N_4946,N_4952);
or UO_585 (O_585,N_4924,N_4993);
nand UO_586 (O_586,N_4925,N_4974);
or UO_587 (O_587,N_4976,N_4949);
or UO_588 (O_588,N_4914,N_4990);
and UO_589 (O_589,N_4933,N_4998);
nand UO_590 (O_590,N_4934,N_4968);
and UO_591 (O_591,N_4923,N_4964);
or UO_592 (O_592,N_4998,N_4948);
xnor UO_593 (O_593,N_4943,N_4982);
and UO_594 (O_594,N_4978,N_4960);
xor UO_595 (O_595,N_4904,N_4954);
nor UO_596 (O_596,N_4991,N_4999);
nand UO_597 (O_597,N_4975,N_4914);
nand UO_598 (O_598,N_4928,N_4961);
nor UO_599 (O_599,N_4989,N_4976);
nor UO_600 (O_600,N_4931,N_4937);
nand UO_601 (O_601,N_4971,N_4923);
or UO_602 (O_602,N_4954,N_4938);
nand UO_603 (O_603,N_4977,N_4987);
nand UO_604 (O_604,N_4916,N_4925);
and UO_605 (O_605,N_4931,N_4968);
nand UO_606 (O_606,N_4900,N_4945);
nand UO_607 (O_607,N_4958,N_4992);
and UO_608 (O_608,N_4920,N_4991);
and UO_609 (O_609,N_4910,N_4995);
and UO_610 (O_610,N_4958,N_4994);
xnor UO_611 (O_611,N_4939,N_4920);
or UO_612 (O_612,N_4968,N_4962);
nor UO_613 (O_613,N_4922,N_4917);
nor UO_614 (O_614,N_4958,N_4991);
or UO_615 (O_615,N_4945,N_4977);
nand UO_616 (O_616,N_4911,N_4917);
and UO_617 (O_617,N_4964,N_4925);
nor UO_618 (O_618,N_4901,N_4977);
or UO_619 (O_619,N_4910,N_4980);
nand UO_620 (O_620,N_4965,N_4957);
and UO_621 (O_621,N_4967,N_4938);
nand UO_622 (O_622,N_4950,N_4977);
nor UO_623 (O_623,N_4943,N_4968);
or UO_624 (O_624,N_4905,N_4915);
nor UO_625 (O_625,N_4985,N_4977);
and UO_626 (O_626,N_4959,N_4911);
or UO_627 (O_627,N_4953,N_4922);
and UO_628 (O_628,N_4922,N_4996);
or UO_629 (O_629,N_4930,N_4948);
and UO_630 (O_630,N_4906,N_4912);
nor UO_631 (O_631,N_4998,N_4918);
xor UO_632 (O_632,N_4983,N_4922);
nand UO_633 (O_633,N_4995,N_4983);
nand UO_634 (O_634,N_4909,N_4934);
or UO_635 (O_635,N_4992,N_4953);
xor UO_636 (O_636,N_4940,N_4941);
nand UO_637 (O_637,N_4948,N_4916);
nor UO_638 (O_638,N_4959,N_4945);
nand UO_639 (O_639,N_4939,N_4968);
xnor UO_640 (O_640,N_4918,N_4972);
and UO_641 (O_641,N_4906,N_4978);
nor UO_642 (O_642,N_4922,N_4982);
nor UO_643 (O_643,N_4983,N_4921);
nor UO_644 (O_644,N_4919,N_4903);
nand UO_645 (O_645,N_4951,N_4945);
or UO_646 (O_646,N_4954,N_4966);
and UO_647 (O_647,N_4965,N_4993);
xnor UO_648 (O_648,N_4932,N_4924);
or UO_649 (O_649,N_4994,N_4947);
nand UO_650 (O_650,N_4906,N_4926);
and UO_651 (O_651,N_4987,N_4929);
or UO_652 (O_652,N_4946,N_4920);
xor UO_653 (O_653,N_4918,N_4997);
xnor UO_654 (O_654,N_4999,N_4905);
and UO_655 (O_655,N_4985,N_4929);
and UO_656 (O_656,N_4954,N_4977);
nand UO_657 (O_657,N_4945,N_4904);
nor UO_658 (O_658,N_4942,N_4980);
nor UO_659 (O_659,N_4915,N_4935);
and UO_660 (O_660,N_4941,N_4934);
and UO_661 (O_661,N_4905,N_4997);
or UO_662 (O_662,N_4995,N_4938);
nor UO_663 (O_663,N_4904,N_4955);
nor UO_664 (O_664,N_4915,N_4966);
nor UO_665 (O_665,N_4960,N_4924);
or UO_666 (O_666,N_4941,N_4995);
nand UO_667 (O_667,N_4958,N_4948);
nor UO_668 (O_668,N_4934,N_4916);
nand UO_669 (O_669,N_4964,N_4983);
or UO_670 (O_670,N_4933,N_4920);
nor UO_671 (O_671,N_4900,N_4996);
or UO_672 (O_672,N_4954,N_4939);
xnor UO_673 (O_673,N_4906,N_4956);
and UO_674 (O_674,N_4951,N_4923);
nand UO_675 (O_675,N_4993,N_4987);
or UO_676 (O_676,N_4936,N_4997);
xnor UO_677 (O_677,N_4980,N_4960);
and UO_678 (O_678,N_4914,N_4916);
and UO_679 (O_679,N_4904,N_4907);
and UO_680 (O_680,N_4918,N_4954);
nand UO_681 (O_681,N_4942,N_4943);
or UO_682 (O_682,N_4994,N_4964);
nand UO_683 (O_683,N_4947,N_4911);
nor UO_684 (O_684,N_4977,N_4940);
nor UO_685 (O_685,N_4973,N_4988);
nor UO_686 (O_686,N_4952,N_4984);
nand UO_687 (O_687,N_4998,N_4995);
xor UO_688 (O_688,N_4912,N_4990);
or UO_689 (O_689,N_4927,N_4969);
or UO_690 (O_690,N_4979,N_4918);
nor UO_691 (O_691,N_4900,N_4910);
nor UO_692 (O_692,N_4995,N_4928);
nor UO_693 (O_693,N_4946,N_4945);
and UO_694 (O_694,N_4936,N_4966);
xnor UO_695 (O_695,N_4928,N_4912);
nor UO_696 (O_696,N_4978,N_4969);
and UO_697 (O_697,N_4907,N_4922);
nor UO_698 (O_698,N_4952,N_4970);
and UO_699 (O_699,N_4982,N_4945);
nor UO_700 (O_700,N_4998,N_4959);
and UO_701 (O_701,N_4954,N_4959);
nor UO_702 (O_702,N_4932,N_4928);
and UO_703 (O_703,N_4965,N_4913);
and UO_704 (O_704,N_4912,N_4945);
nand UO_705 (O_705,N_4979,N_4955);
xor UO_706 (O_706,N_4902,N_4917);
xor UO_707 (O_707,N_4911,N_4901);
and UO_708 (O_708,N_4925,N_4994);
nand UO_709 (O_709,N_4905,N_4926);
and UO_710 (O_710,N_4902,N_4948);
and UO_711 (O_711,N_4967,N_4915);
nand UO_712 (O_712,N_4991,N_4939);
or UO_713 (O_713,N_4981,N_4922);
xor UO_714 (O_714,N_4973,N_4952);
nand UO_715 (O_715,N_4931,N_4926);
and UO_716 (O_716,N_4910,N_4923);
and UO_717 (O_717,N_4965,N_4969);
xor UO_718 (O_718,N_4987,N_4964);
nand UO_719 (O_719,N_4917,N_4996);
and UO_720 (O_720,N_4979,N_4985);
nor UO_721 (O_721,N_4911,N_4900);
or UO_722 (O_722,N_4955,N_4918);
nand UO_723 (O_723,N_4948,N_4920);
nor UO_724 (O_724,N_4930,N_4926);
nor UO_725 (O_725,N_4960,N_4902);
nand UO_726 (O_726,N_4902,N_4906);
nor UO_727 (O_727,N_4948,N_4979);
xor UO_728 (O_728,N_4978,N_4910);
nor UO_729 (O_729,N_4957,N_4945);
nor UO_730 (O_730,N_4903,N_4922);
nor UO_731 (O_731,N_4979,N_4905);
nor UO_732 (O_732,N_4900,N_4929);
xor UO_733 (O_733,N_4924,N_4942);
nor UO_734 (O_734,N_4947,N_4948);
or UO_735 (O_735,N_4918,N_4958);
nand UO_736 (O_736,N_4950,N_4900);
and UO_737 (O_737,N_4904,N_4951);
and UO_738 (O_738,N_4919,N_4939);
or UO_739 (O_739,N_4961,N_4982);
or UO_740 (O_740,N_4931,N_4923);
nand UO_741 (O_741,N_4950,N_4926);
nor UO_742 (O_742,N_4990,N_4916);
and UO_743 (O_743,N_4993,N_4918);
or UO_744 (O_744,N_4977,N_4964);
nor UO_745 (O_745,N_4936,N_4918);
and UO_746 (O_746,N_4932,N_4995);
nor UO_747 (O_747,N_4954,N_4952);
nand UO_748 (O_748,N_4944,N_4992);
and UO_749 (O_749,N_4997,N_4931);
or UO_750 (O_750,N_4994,N_4974);
or UO_751 (O_751,N_4955,N_4916);
nor UO_752 (O_752,N_4996,N_4903);
and UO_753 (O_753,N_4942,N_4971);
and UO_754 (O_754,N_4931,N_4927);
and UO_755 (O_755,N_4941,N_4958);
nor UO_756 (O_756,N_4954,N_4937);
nor UO_757 (O_757,N_4951,N_4929);
and UO_758 (O_758,N_4938,N_4946);
and UO_759 (O_759,N_4943,N_4922);
and UO_760 (O_760,N_4926,N_4964);
and UO_761 (O_761,N_4967,N_4999);
xor UO_762 (O_762,N_4980,N_4923);
nand UO_763 (O_763,N_4902,N_4900);
and UO_764 (O_764,N_4916,N_4959);
nor UO_765 (O_765,N_4986,N_4993);
xor UO_766 (O_766,N_4986,N_4936);
and UO_767 (O_767,N_4995,N_4924);
nand UO_768 (O_768,N_4941,N_4967);
or UO_769 (O_769,N_4981,N_4909);
nor UO_770 (O_770,N_4952,N_4951);
nor UO_771 (O_771,N_4938,N_4945);
nor UO_772 (O_772,N_4997,N_4930);
xor UO_773 (O_773,N_4909,N_4921);
xnor UO_774 (O_774,N_4908,N_4998);
nand UO_775 (O_775,N_4974,N_4905);
nand UO_776 (O_776,N_4914,N_4940);
or UO_777 (O_777,N_4946,N_4984);
or UO_778 (O_778,N_4992,N_4902);
nand UO_779 (O_779,N_4927,N_4974);
xor UO_780 (O_780,N_4911,N_4958);
nand UO_781 (O_781,N_4997,N_4924);
nand UO_782 (O_782,N_4967,N_4947);
or UO_783 (O_783,N_4991,N_4936);
or UO_784 (O_784,N_4905,N_4942);
nand UO_785 (O_785,N_4929,N_4968);
nand UO_786 (O_786,N_4941,N_4996);
nand UO_787 (O_787,N_4963,N_4967);
or UO_788 (O_788,N_4939,N_4940);
or UO_789 (O_789,N_4943,N_4907);
nor UO_790 (O_790,N_4916,N_4927);
nand UO_791 (O_791,N_4901,N_4903);
or UO_792 (O_792,N_4970,N_4910);
and UO_793 (O_793,N_4924,N_4922);
xnor UO_794 (O_794,N_4982,N_4912);
nor UO_795 (O_795,N_4967,N_4925);
or UO_796 (O_796,N_4912,N_4946);
nand UO_797 (O_797,N_4938,N_4920);
nand UO_798 (O_798,N_4905,N_4956);
and UO_799 (O_799,N_4944,N_4923);
and UO_800 (O_800,N_4955,N_4981);
nand UO_801 (O_801,N_4940,N_4983);
nand UO_802 (O_802,N_4949,N_4986);
and UO_803 (O_803,N_4925,N_4904);
or UO_804 (O_804,N_4977,N_4963);
nand UO_805 (O_805,N_4992,N_4999);
or UO_806 (O_806,N_4992,N_4911);
nand UO_807 (O_807,N_4929,N_4947);
and UO_808 (O_808,N_4979,N_4966);
nand UO_809 (O_809,N_4958,N_4952);
or UO_810 (O_810,N_4960,N_4968);
and UO_811 (O_811,N_4987,N_4999);
nand UO_812 (O_812,N_4959,N_4934);
nor UO_813 (O_813,N_4941,N_4948);
and UO_814 (O_814,N_4968,N_4907);
or UO_815 (O_815,N_4983,N_4960);
nor UO_816 (O_816,N_4925,N_4985);
nor UO_817 (O_817,N_4964,N_4981);
or UO_818 (O_818,N_4985,N_4949);
xor UO_819 (O_819,N_4919,N_4952);
or UO_820 (O_820,N_4963,N_4990);
nor UO_821 (O_821,N_4980,N_4932);
nor UO_822 (O_822,N_4970,N_4954);
xnor UO_823 (O_823,N_4909,N_4923);
and UO_824 (O_824,N_4954,N_4906);
nand UO_825 (O_825,N_4972,N_4905);
or UO_826 (O_826,N_4926,N_4990);
and UO_827 (O_827,N_4987,N_4905);
or UO_828 (O_828,N_4919,N_4942);
and UO_829 (O_829,N_4900,N_4997);
nand UO_830 (O_830,N_4996,N_4910);
nand UO_831 (O_831,N_4966,N_4952);
and UO_832 (O_832,N_4985,N_4930);
and UO_833 (O_833,N_4957,N_4909);
xor UO_834 (O_834,N_4962,N_4996);
xnor UO_835 (O_835,N_4941,N_4937);
and UO_836 (O_836,N_4938,N_4991);
xnor UO_837 (O_837,N_4954,N_4901);
nor UO_838 (O_838,N_4932,N_4906);
and UO_839 (O_839,N_4954,N_4935);
nand UO_840 (O_840,N_4974,N_4926);
or UO_841 (O_841,N_4930,N_4942);
or UO_842 (O_842,N_4921,N_4905);
nand UO_843 (O_843,N_4904,N_4932);
and UO_844 (O_844,N_4900,N_4924);
or UO_845 (O_845,N_4917,N_4948);
xor UO_846 (O_846,N_4987,N_4900);
or UO_847 (O_847,N_4947,N_4955);
nor UO_848 (O_848,N_4912,N_4985);
and UO_849 (O_849,N_4924,N_4985);
and UO_850 (O_850,N_4926,N_4924);
nand UO_851 (O_851,N_4956,N_4933);
and UO_852 (O_852,N_4945,N_4936);
nor UO_853 (O_853,N_4954,N_4971);
xnor UO_854 (O_854,N_4929,N_4938);
or UO_855 (O_855,N_4989,N_4906);
xnor UO_856 (O_856,N_4996,N_4921);
nor UO_857 (O_857,N_4996,N_4993);
and UO_858 (O_858,N_4994,N_4962);
or UO_859 (O_859,N_4921,N_4952);
nand UO_860 (O_860,N_4936,N_4930);
nand UO_861 (O_861,N_4933,N_4932);
and UO_862 (O_862,N_4921,N_4980);
nand UO_863 (O_863,N_4910,N_4926);
nor UO_864 (O_864,N_4916,N_4930);
or UO_865 (O_865,N_4947,N_4975);
and UO_866 (O_866,N_4968,N_4986);
xnor UO_867 (O_867,N_4945,N_4968);
and UO_868 (O_868,N_4908,N_4945);
and UO_869 (O_869,N_4950,N_4913);
and UO_870 (O_870,N_4910,N_4952);
or UO_871 (O_871,N_4998,N_4982);
nor UO_872 (O_872,N_4982,N_4914);
nand UO_873 (O_873,N_4906,N_4946);
nor UO_874 (O_874,N_4960,N_4957);
nand UO_875 (O_875,N_4970,N_4989);
or UO_876 (O_876,N_4970,N_4905);
or UO_877 (O_877,N_4932,N_4951);
nor UO_878 (O_878,N_4968,N_4910);
nor UO_879 (O_879,N_4973,N_4972);
or UO_880 (O_880,N_4974,N_4977);
and UO_881 (O_881,N_4921,N_4940);
and UO_882 (O_882,N_4996,N_4931);
or UO_883 (O_883,N_4974,N_4963);
nor UO_884 (O_884,N_4903,N_4979);
or UO_885 (O_885,N_4947,N_4920);
or UO_886 (O_886,N_4989,N_4998);
or UO_887 (O_887,N_4991,N_4924);
nand UO_888 (O_888,N_4993,N_4933);
nor UO_889 (O_889,N_4984,N_4966);
or UO_890 (O_890,N_4981,N_4904);
xnor UO_891 (O_891,N_4934,N_4982);
nand UO_892 (O_892,N_4935,N_4970);
and UO_893 (O_893,N_4917,N_4915);
nor UO_894 (O_894,N_4973,N_4961);
nor UO_895 (O_895,N_4942,N_4966);
nor UO_896 (O_896,N_4964,N_4945);
nand UO_897 (O_897,N_4982,N_4980);
and UO_898 (O_898,N_4989,N_4985);
nor UO_899 (O_899,N_4956,N_4912);
and UO_900 (O_900,N_4986,N_4942);
and UO_901 (O_901,N_4983,N_4948);
or UO_902 (O_902,N_4911,N_4929);
nand UO_903 (O_903,N_4906,N_4995);
nand UO_904 (O_904,N_4920,N_4988);
nor UO_905 (O_905,N_4961,N_4918);
or UO_906 (O_906,N_4962,N_4952);
and UO_907 (O_907,N_4913,N_4918);
nand UO_908 (O_908,N_4958,N_4990);
xor UO_909 (O_909,N_4911,N_4936);
nand UO_910 (O_910,N_4979,N_4941);
or UO_911 (O_911,N_4985,N_4907);
or UO_912 (O_912,N_4933,N_4991);
nand UO_913 (O_913,N_4921,N_4907);
nand UO_914 (O_914,N_4961,N_4921);
or UO_915 (O_915,N_4969,N_4930);
nor UO_916 (O_916,N_4937,N_4927);
and UO_917 (O_917,N_4951,N_4996);
or UO_918 (O_918,N_4902,N_4979);
nand UO_919 (O_919,N_4953,N_4989);
and UO_920 (O_920,N_4950,N_4972);
or UO_921 (O_921,N_4932,N_4988);
or UO_922 (O_922,N_4983,N_4943);
nand UO_923 (O_923,N_4987,N_4988);
nor UO_924 (O_924,N_4914,N_4917);
and UO_925 (O_925,N_4926,N_4992);
nor UO_926 (O_926,N_4937,N_4997);
nor UO_927 (O_927,N_4958,N_4929);
nor UO_928 (O_928,N_4910,N_4928);
xor UO_929 (O_929,N_4901,N_4944);
nor UO_930 (O_930,N_4907,N_4974);
nor UO_931 (O_931,N_4957,N_4950);
and UO_932 (O_932,N_4906,N_4959);
nand UO_933 (O_933,N_4954,N_4945);
or UO_934 (O_934,N_4933,N_4931);
and UO_935 (O_935,N_4986,N_4967);
nor UO_936 (O_936,N_4990,N_4925);
nor UO_937 (O_937,N_4954,N_4976);
xnor UO_938 (O_938,N_4904,N_4957);
xnor UO_939 (O_939,N_4947,N_4902);
and UO_940 (O_940,N_4914,N_4960);
and UO_941 (O_941,N_4903,N_4963);
and UO_942 (O_942,N_4951,N_4931);
xnor UO_943 (O_943,N_4972,N_4914);
nor UO_944 (O_944,N_4971,N_4993);
nand UO_945 (O_945,N_4961,N_4953);
nand UO_946 (O_946,N_4944,N_4915);
or UO_947 (O_947,N_4900,N_4957);
and UO_948 (O_948,N_4912,N_4920);
nand UO_949 (O_949,N_4932,N_4990);
and UO_950 (O_950,N_4944,N_4956);
nand UO_951 (O_951,N_4984,N_4970);
and UO_952 (O_952,N_4954,N_4997);
nand UO_953 (O_953,N_4996,N_4988);
xor UO_954 (O_954,N_4906,N_4908);
and UO_955 (O_955,N_4922,N_4915);
or UO_956 (O_956,N_4904,N_4979);
and UO_957 (O_957,N_4997,N_4927);
or UO_958 (O_958,N_4903,N_4900);
or UO_959 (O_959,N_4922,N_4973);
and UO_960 (O_960,N_4964,N_4947);
nor UO_961 (O_961,N_4979,N_4943);
and UO_962 (O_962,N_4975,N_4954);
and UO_963 (O_963,N_4903,N_4985);
nor UO_964 (O_964,N_4957,N_4976);
nand UO_965 (O_965,N_4912,N_4919);
nand UO_966 (O_966,N_4977,N_4939);
nand UO_967 (O_967,N_4934,N_4995);
nor UO_968 (O_968,N_4987,N_4980);
xor UO_969 (O_969,N_4959,N_4908);
nor UO_970 (O_970,N_4911,N_4915);
and UO_971 (O_971,N_4900,N_4936);
nor UO_972 (O_972,N_4921,N_4930);
or UO_973 (O_973,N_4963,N_4998);
or UO_974 (O_974,N_4941,N_4984);
nor UO_975 (O_975,N_4973,N_4963);
nand UO_976 (O_976,N_4921,N_4926);
or UO_977 (O_977,N_4960,N_4913);
xnor UO_978 (O_978,N_4985,N_4995);
nor UO_979 (O_979,N_4960,N_4923);
xnor UO_980 (O_980,N_4915,N_4916);
nor UO_981 (O_981,N_4933,N_4928);
nand UO_982 (O_982,N_4947,N_4952);
or UO_983 (O_983,N_4970,N_4938);
nor UO_984 (O_984,N_4987,N_4931);
nor UO_985 (O_985,N_4905,N_4940);
nor UO_986 (O_986,N_4976,N_4955);
nor UO_987 (O_987,N_4995,N_4978);
and UO_988 (O_988,N_4902,N_4972);
or UO_989 (O_989,N_4989,N_4941);
nand UO_990 (O_990,N_4984,N_4906);
and UO_991 (O_991,N_4938,N_4957);
or UO_992 (O_992,N_4989,N_4983);
nor UO_993 (O_993,N_4964,N_4965);
or UO_994 (O_994,N_4939,N_4925);
or UO_995 (O_995,N_4961,N_4995);
or UO_996 (O_996,N_4958,N_4938);
nand UO_997 (O_997,N_4983,N_4968);
nor UO_998 (O_998,N_4927,N_4947);
nor UO_999 (O_999,N_4902,N_4901);
endmodule