module basic_1500_15000_2000_10_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_86,In_710);
and U1 (N_1,In_471,In_1482);
or U2 (N_2,In_641,In_1471);
and U3 (N_3,In_906,In_420);
or U4 (N_4,In_237,In_1344);
or U5 (N_5,In_566,In_610);
or U6 (N_6,In_1372,In_624);
nor U7 (N_7,In_1468,In_495);
and U8 (N_8,In_1031,In_1097);
nand U9 (N_9,In_1219,In_3);
nand U10 (N_10,In_21,In_1360);
nor U11 (N_11,In_274,In_694);
or U12 (N_12,In_1241,In_850);
and U13 (N_13,In_857,In_130);
nand U14 (N_14,In_1042,In_1083);
nand U15 (N_15,In_1200,In_1492);
nand U16 (N_16,In_639,In_398);
or U17 (N_17,In_760,In_1285);
or U18 (N_18,In_133,In_393);
nor U19 (N_19,In_1393,In_308);
nand U20 (N_20,In_517,In_339);
or U21 (N_21,In_273,In_178);
nor U22 (N_22,In_1239,In_942);
and U23 (N_23,In_7,In_464);
nor U24 (N_24,In_1428,In_93);
xor U25 (N_25,In_43,In_985);
or U26 (N_26,In_1040,In_1397);
nor U27 (N_27,In_194,In_895);
nand U28 (N_28,In_190,In_1033);
nand U29 (N_29,In_235,In_536);
xnor U30 (N_30,In_980,In_307);
xor U31 (N_31,In_672,In_356);
or U32 (N_32,In_423,In_685);
or U33 (N_33,In_12,In_426);
nand U34 (N_34,In_68,In_733);
nor U35 (N_35,In_452,In_1401);
or U36 (N_36,In_1298,In_1170);
or U37 (N_37,In_199,In_472);
or U38 (N_38,In_1044,In_1423);
nand U39 (N_39,In_684,In_1497);
and U40 (N_40,In_166,In_458);
nor U41 (N_41,In_80,In_1457);
and U42 (N_42,In_1391,In_643);
nand U43 (N_43,In_395,In_888);
and U44 (N_44,In_795,In_279);
xor U45 (N_45,In_1163,In_303);
or U46 (N_46,In_413,In_174);
nand U47 (N_47,In_1375,In_848);
and U48 (N_48,In_820,In_616);
xor U49 (N_49,In_439,In_160);
and U50 (N_50,In_329,In_1351);
nand U51 (N_51,In_534,In_1355);
nand U52 (N_52,In_1187,In_498);
and U53 (N_53,In_1151,In_100);
or U54 (N_54,In_778,In_103);
nand U55 (N_55,In_409,In_1362);
and U56 (N_56,In_1314,In_1158);
xnor U57 (N_57,In_806,In_392);
nor U58 (N_58,In_1070,In_1150);
nor U59 (N_59,In_667,In_1093);
nand U60 (N_60,In_76,In_868);
and U61 (N_61,In_1244,In_1107);
nor U62 (N_62,In_1307,In_350);
nor U63 (N_63,In_847,In_61);
xor U64 (N_64,In_309,In_703);
nor U65 (N_65,In_430,In_1133);
or U66 (N_66,In_262,In_1126);
nor U67 (N_67,In_825,In_33);
nand U68 (N_68,In_553,In_151);
nand U69 (N_69,In_922,In_280);
nor U70 (N_70,In_1231,In_225);
and U71 (N_71,In_571,In_975);
nor U72 (N_72,In_1395,In_111);
or U73 (N_73,In_819,In_348);
nor U74 (N_74,In_527,In_1335);
and U75 (N_75,In_289,In_1090);
and U76 (N_76,In_700,In_1232);
nand U77 (N_77,In_1342,In_1384);
nand U78 (N_78,In_351,In_1488);
and U79 (N_79,In_1218,In_45);
and U80 (N_80,In_406,In_572);
nor U81 (N_81,In_1141,In_758);
and U82 (N_82,In_154,In_243);
nor U83 (N_83,In_335,In_810);
nor U84 (N_84,In_278,In_405);
and U85 (N_85,In_805,In_46);
or U86 (N_86,In_401,In_1011);
nor U87 (N_87,In_1356,In_1332);
or U88 (N_88,In_705,In_345);
or U89 (N_89,In_604,In_854);
and U90 (N_90,In_821,In_164);
xor U91 (N_91,In_418,In_1366);
and U92 (N_92,In_427,In_696);
and U93 (N_93,In_182,In_124);
nand U94 (N_94,In_1319,In_42);
nand U95 (N_95,In_484,In_1398);
xor U96 (N_96,In_1123,In_925);
nand U97 (N_97,In_780,In_1006);
nand U98 (N_98,In_853,In_287);
or U99 (N_99,In_1131,In_1414);
and U100 (N_100,In_263,In_669);
nor U101 (N_101,In_1444,In_569);
and U102 (N_102,In_429,In_374);
nand U103 (N_103,In_1212,In_1075);
and U104 (N_104,In_217,In_739);
nand U105 (N_105,In_533,In_4);
or U106 (N_106,In_294,In_869);
or U107 (N_107,In_1230,In_1221);
and U108 (N_108,In_658,In_1422);
and U109 (N_109,In_707,In_276);
or U110 (N_110,In_1092,In_593);
nand U111 (N_111,In_1207,In_69);
xnor U112 (N_112,In_1122,In_1143);
nor U113 (N_113,In_1287,In_1016);
nand U114 (N_114,In_603,In_607);
nor U115 (N_115,In_500,In_874);
or U116 (N_116,In_1279,In_875);
and U117 (N_117,In_355,In_927);
nor U118 (N_118,In_878,In_1328);
nor U119 (N_119,In_1273,In_1050);
and U120 (N_120,In_488,In_838);
or U121 (N_121,In_1118,In_862);
nor U122 (N_122,In_336,In_908);
nor U123 (N_123,In_267,In_621);
or U124 (N_124,In_631,In_301);
and U125 (N_125,In_911,In_383);
or U126 (N_126,In_288,In_552);
nand U127 (N_127,In_1369,In_620);
and U128 (N_128,In_1357,In_724);
nor U129 (N_129,In_41,In_1448);
or U130 (N_130,In_670,In_866);
nand U131 (N_131,In_731,In_1078);
nor U132 (N_132,In_944,In_952);
or U133 (N_133,In_318,In_40);
and U134 (N_134,In_1409,In_656);
or U135 (N_135,In_735,In_636);
nor U136 (N_136,In_1489,In_1301);
nand U137 (N_137,In_186,In_719);
nor U138 (N_138,In_883,In_919);
nand U139 (N_139,In_1140,In_998);
and U140 (N_140,In_408,In_1115);
nor U141 (N_141,In_327,In_491);
nand U142 (N_142,In_1108,In_1077);
or U143 (N_143,In_1173,In_157);
nor U144 (N_144,In_203,In_972);
or U145 (N_145,In_1379,In_389);
or U146 (N_146,In_1034,In_489);
or U147 (N_147,In_118,In_814);
or U148 (N_148,In_994,In_1449);
or U149 (N_149,In_894,In_990);
nand U150 (N_150,In_1165,In_150);
and U151 (N_151,In_1308,In_940);
nand U152 (N_152,In_1076,In_1343);
nand U153 (N_153,In_297,In_730);
nand U154 (N_154,In_1100,In_1396);
or U155 (N_155,In_549,In_991);
or U156 (N_156,In_417,In_982);
nand U157 (N_157,In_1333,In_57);
or U158 (N_158,In_956,In_372);
nor U159 (N_159,In_729,In_767);
and U160 (N_160,In_1464,In_1469);
or U161 (N_161,In_269,In_958);
or U162 (N_162,In_817,In_465);
or U163 (N_163,In_367,In_320);
nor U164 (N_164,In_496,In_775);
and U165 (N_165,In_912,In_1121);
and U166 (N_166,In_554,In_611);
and U167 (N_167,In_822,In_451);
nor U168 (N_168,In_434,In_468);
and U169 (N_169,In_1089,In_959);
nand U170 (N_170,In_248,In_896);
and U171 (N_171,In_1327,In_415);
and U172 (N_172,In_1256,In_380);
nand U173 (N_173,In_1224,In_26);
and U174 (N_174,In_793,In_523);
or U175 (N_175,In_547,In_1295);
and U176 (N_176,In_1446,In_357);
and U177 (N_177,In_1094,In_1196);
and U178 (N_178,In_622,In_844);
xor U179 (N_179,In_699,In_1250);
or U180 (N_180,In_1254,In_1443);
nand U181 (N_181,In_75,In_1168);
nor U182 (N_182,In_1450,In_67);
and U183 (N_183,In_1157,In_938);
or U184 (N_184,In_747,In_158);
and U185 (N_185,In_926,In_344);
nand U186 (N_186,In_1037,In_663);
nand U187 (N_187,In_843,In_1381);
nor U188 (N_188,In_1420,In_1211);
nor U189 (N_189,In_575,In_1405);
nor U190 (N_190,In_626,In_24);
or U191 (N_191,In_200,In_1080);
nand U192 (N_192,In_286,In_752);
nand U193 (N_193,In_1260,In_183);
or U194 (N_194,In_613,In_1478);
and U195 (N_195,In_6,In_1098);
nor U196 (N_196,In_1205,In_1291);
or U197 (N_197,In_461,In_347);
nand U198 (N_198,In_1208,In_826);
or U199 (N_199,In_70,In_846);
nand U200 (N_200,In_1074,In_394);
and U201 (N_201,In_411,In_445);
or U202 (N_202,In_818,In_1172);
or U203 (N_203,In_708,In_419);
nand U204 (N_204,In_591,In_1104);
nor U205 (N_205,In_646,In_233);
nor U206 (N_206,In_598,In_628);
nor U207 (N_207,In_156,In_44);
or U208 (N_208,In_997,In_904);
and U209 (N_209,In_755,In_58);
nor U210 (N_210,In_644,In_1311);
nor U211 (N_211,In_510,In_1102);
nand U212 (N_212,In_1462,In_686);
and U213 (N_213,In_521,In_13);
or U214 (N_214,In_258,In_1043);
nor U215 (N_215,In_893,In_1303);
nor U216 (N_216,In_424,In_910);
and U217 (N_217,In_1214,In_65);
nand U218 (N_218,In_1029,In_1310);
and U219 (N_219,In_1290,In_447);
and U220 (N_220,In_1154,In_737);
or U221 (N_221,In_298,In_1277);
nand U222 (N_222,In_711,In_785);
nor U223 (N_223,In_790,In_1371);
nand U224 (N_224,In_1062,In_712);
nand U225 (N_225,In_583,In_1321);
xor U226 (N_226,In_941,In_541);
or U227 (N_227,In_1215,In_32);
or U228 (N_228,In_291,In_1058);
nand U229 (N_229,In_49,In_1156);
xor U230 (N_230,In_833,In_625);
xor U231 (N_231,In_535,In_513);
and U232 (N_232,In_104,In_860);
or U233 (N_233,In_977,In_689);
and U234 (N_234,In_2,In_511);
nor U235 (N_235,In_1025,In_1024);
nor U236 (N_236,In_797,In_698);
nand U237 (N_237,In_789,In_403);
and U238 (N_238,In_1278,In_487);
nor U239 (N_239,In_619,In_1480);
and U240 (N_240,In_1179,In_1174);
nor U241 (N_241,In_1269,In_665);
or U242 (N_242,In_829,In_691);
or U243 (N_243,In_1383,In_1368);
xor U244 (N_244,In_1353,In_1010);
or U245 (N_245,In_664,In_1286);
nand U246 (N_246,In_141,In_635);
and U247 (N_247,In_390,In_282);
or U248 (N_248,In_249,In_581);
or U249 (N_249,In_907,In_108);
or U250 (N_250,In_518,In_1474);
nor U251 (N_251,In_470,In_1068);
xor U252 (N_252,In_211,In_317);
nor U253 (N_253,In_845,In_1385);
and U254 (N_254,In_192,In_1316);
nor U255 (N_255,In_978,In_1106);
nand U256 (N_256,In_202,In_361);
or U257 (N_257,In_281,In_650);
and U258 (N_258,In_792,In_557);
nor U259 (N_259,In_695,In_1326);
nor U260 (N_260,In_531,In_90);
and U261 (N_261,In_1159,In_768);
nor U262 (N_262,In_1268,In_1477);
or U263 (N_263,In_1441,In_51);
and U264 (N_264,In_1201,In_1417);
nor U265 (N_265,In_476,In_1236);
nor U266 (N_266,In_1117,In_1394);
and U267 (N_267,In_1112,In_834);
nor U268 (N_268,In_1467,In_765);
nor U269 (N_269,In_220,In_384);
and U270 (N_270,In_928,In_995);
nand U271 (N_271,In_609,In_921);
xnor U272 (N_272,In_74,In_503);
nor U273 (N_273,In_1387,In_1087);
nand U274 (N_274,In_1247,In_453);
nor U275 (N_275,In_1007,In_891);
or U276 (N_276,In_378,In_195);
and U277 (N_277,In_1051,In_1354);
or U278 (N_278,In_126,In_497);
nand U279 (N_279,In_968,In_1005);
nand U280 (N_280,In_1041,In_1145);
nor U281 (N_281,In_647,In_584);
nand U282 (N_282,In_270,In_1341);
nand U283 (N_283,In_1063,In_1408);
nand U284 (N_284,In_448,In_128);
nand U285 (N_285,In_828,In_467);
nand U286 (N_286,In_1252,In_608);
and U287 (N_287,In_746,In_543);
or U288 (N_288,In_1323,In_596);
and U289 (N_289,In_537,In_592);
and U290 (N_290,In_1389,In_201);
and U291 (N_291,In_138,In_240);
and U292 (N_292,In_1125,In_936);
nand U293 (N_293,In_149,In_221);
nand U294 (N_294,In_1082,In_94);
or U295 (N_295,In_957,In_119);
xnor U296 (N_296,In_78,In_736);
nand U297 (N_297,In_1110,In_121);
nand U298 (N_298,In_771,In_824);
or U299 (N_299,In_769,In_87);
nand U300 (N_300,In_1484,In_479);
or U301 (N_301,In_1410,In_565);
or U302 (N_302,In_1223,In_1259);
or U303 (N_303,In_349,In_473);
nand U304 (N_304,In_1237,In_98);
nor U305 (N_305,In_244,In_526);
or U306 (N_306,In_839,In_1304);
and U307 (N_307,In_198,In_1160);
nor U308 (N_308,In_153,In_1403);
nand U309 (N_309,In_723,In_882);
nand U310 (N_310,In_1442,In_811);
and U311 (N_311,In_62,In_807);
nand U312 (N_312,In_568,In_377);
nor U313 (N_313,In_1209,In_1400);
and U314 (N_314,In_1284,In_946);
or U315 (N_315,In_683,In_677);
nor U316 (N_316,In_227,In_343);
or U317 (N_317,In_82,In_779);
nor U318 (N_318,In_594,In_1348);
nand U319 (N_319,In_1014,In_1280);
or U320 (N_320,In_18,In_903);
and U321 (N_321,In_776,In_340);
nand U322 (N_322,In_1137,In_81);
or U323 (N_323,In_326,In_1459);
nand U324 (N_324,In_673,In_1128);
nand U325 (N_325,In_823,In_512);
nand U326 (N_326,In_1318,In_1465);
xnor U327 (N_327,In_1032,In_319);
nor U328 (N_328,In_931,In_97);
nand U329 (N_329,In_1048,In_802);
or U330 (N_330,In_1195,In_561);
nor U331 (N_331,In_163,In_987);
nor U332 (N_332,In_1296,In_214);
or U333 (N_333,In_1021,In_144);
nor U334 (N_334,In_1003,In_1091);
xnor U335 (N_335,In_352,In_1086);
and U336 (N_336,In_905,In_983);
nand U337 (N_337,In_1057,In_272);
nand U338 (N_338,In_546,In_618);
nor U339 (N_339,In_979,In_1015);
nor U340 (N_340,In_1073,In_1175);
nand U341 (N_341,In_713,In_757);
and U342 (N_342,In_1222,In_122);
nand U343 (N_343,In_1146,In_1220);
or U344 (N_344,In_212,In_1018);
xnor U345 (N_345,In_586,In_105);
nor U346 (N_346,In_358,In_84);
or U347 (N_347,In_697,In_191);
nand U348 (N_348,In_544,In_659);
nand U349 (N_349,In_271,In_816);
nor U350 (N_350,In_1065,In_169);
xnor U351 (N_351,In_582,In_1498);
nand U352 (N_352,In_52,In_1402);
nor U353 (N_353,In_387,In_754);
or U354 (N_354,In_359,In_332);
or U355 (N_355,In_83,In_64);
nor U356 (N_356,In_766,In_187);
nand U357 (N_357,In_316,In_442);
nand U358 (N_358,In_481,In_889);
and U359 (N_359,In_1424,In_11);
and U360 (N_360,In_375,In_478);
nand U361 (N_361,In_1352,In_662);
xnor U362 (N_362,In_168,In_241);
and U363 (N_363,In_1056,In_396);
and U364 (N_364,In_1204,In_1197);
nand U365 (N_365,In_1322,In_1300);
or U366 (N_366,In_1105,In_558);
and U367 (N_367,In_578,In_796);
nand U368 (N_368,In_1476,In_132);
and U369 (N_369,In_1390,In_856);
and U370 (N_370,In_443,In_1475);
nor U371 (N_371,In_388,In_1120);
nand U372 (N_372,In_969,In_490);
nand U373 (N_373,In_599,In_999);
and U374 (N_374,In_750,In_330);
or U375 (N_375,In_175,In_836);
nor U376 (N_376,In_1161,In_916);
or U377 (N_377,In_264,In_277);
nand U378 (N_378,In_1242,In_89);
and U379 (N_379,In_266,In_890);
nor U380 (N_380,In_1113,In_653);
or U381 (N_381,In_1178,In_171);
nand U382 (N_382,In_293,In_1367);
or U383 (N_383,In_371,In_1049);
nor U384 (N_384,In_668,In_177);
and U385 (N_385,In_933,In_831);
nand U386 (N_386,In_1186,In_1176);
or U387 (N_387,In_1499,In_433);
nand U388 (N_388,In_25,In_315);
or U389 (N_389,In_295,In_803);
or U390 (N_390,In_1210,In_887);
nand U391 (N_391,In_849,In_612);
nor U392 (N_392,In_1004,In_897);
or U393 (N_393,In_1067,In_386);
nand U394 (N_394,In_542,In_1181);
nand U395 (N_395,In_462,In_466);
and U396 (N_396,In_363,In_1350);
nand U397 (N_397,In_1226,In_1432);
and U398 (N_398,In_48,In_679);
nor U399 (N_399,In_1217,In_842);
and U400 (N_400,In_954,In_59);
nor U401 (N_401,In_63,In_1228);
and U402 (N_402,In_189,In_1486);
or U403 (N_403,In_743,In_728);
nand U404 (N_404,In_254,In_184);
or U405 (N_405,In_9,In_23);
nand U406 (N_406,In_321,In_1382);
and U407 (N_407,In_455,In_324);
or U408 (N_408,In_1361,In_342);
and U409 (N_409,In_801,In_597);
nand U410 (N_410,In_1061,In_872);
nor U411 (N_411,In_92,In_437);
or U412 (N_412,In_901,In_988);
nand U413 (N_413,In_1138,In_483);
nand U414 (N_414,In_1265,In_870);
or U415 (N_415,In_1017,In_915);
nor U416 (N_416,In_1246,In_1169);
nand U417 (N_417,In_66,In_120);
and U418 (N_418,In_129,In_1233);
nand U419 (N_419,In_170,In_1436);
or U420 (N_420,In_1294,In_617);
and U421 (N_421,In_1306,In_861);
and U422 (N_422,In_222,In_773);
and U423 (N_423,In_140,In_431);
nand U424 (N_424,In_965,In_1243);
nor U425 (N_425,In_1213,In_172);
nor U426 (N_426,In_1270,In_950);
nand U427 (N_427,In_633,In_1225);
or U428 (N_428,In_1136,In_1184);
or U429 (N_429,In_1483,In_210);
or U430 (N_430,In_209,In_207);
or U431 (N_431,In_219,In_595);
or U432 (N_432,In_943,In_475);
or U433 (N_433,In_984,In_346);
or U434 (N_434,In_322,In_146);
or U435 (N_435,In_328,In_955);
or U436 (N_436,In_1292,In_606);
nand U437 (N_437,In_110,In_1199);
and U438 (N_438,In_334,In_204);
and U439 (N_439,In_1251,In_148);
or U440 (N_440,In_223,In_761);
and U441 (N_441,In_1192,In_1008);
and U442 (N_442,In_858,In_962);
and U443 (N_443,In_369,In_506);
or U444 (N_444,In_1188,In_718);
nor U445 (N_445,In_614,In_1490);
xor U446 (N_446,In_36,In_1054);
or U447 (N_447,In_123,In_840);
and U448 (N_448,In_813,In_1019);
and U449 (N_449,In_1142,In_284);
and U450 (N_450,In_1055,In_96);
and U451 (N_451,In_577,In_764);
and U452 (N_452,In_1363,In_841);
or U453 (N_453,In_745,In_333);
and U454 (N_454,In_1426,In_421);
nand U455 (N_455,In_800,In_185);
or U456 (N_456,In_970,In_1012);
nor U457 (N_457,In_937,In_310);
nor U458 (N_458,In_28,In_1013);
or U459 (N_459,In_1203,In_247);
nor U460 (N_460,In_362,In_725);
nor U461 (N_461,In_550,In_717);
nor U462 (N_462,In_116,In_337);
nor U463 (N_463,In_242,In_1191);
nand U464 (N_464,In_1494,In_173);
nand U465 (N_465,In_1144,In_967);
and U466 (N_466,In_304,In_519);
nand U467 (N_467,In_704,In_382);
nor U468 (N_468,In_1466,In_1338);
nand U469 (N_469,In_1315,In_687);
and U470 (N_470,In_1334,In_112);
nor U471 (N_471,In_311,In_1289);
and U472 (N_472,In_645,In_1447);
and U473 (N_473,In_208,In_1458);
or U474 (N_474,In_682,In_1072);
xnor U475 (N_475,In_1404,In_1376);
nor U476 (N_476,In_366,In_145);
nand U477 (N_477,In_1309,In_1111);
nor U478 (N_478,In_1276,In_562);
or U479 (N_479,In_215,In_640);
xnor U480 (N_480,In_226,In_630);
xor U481 (N_481,In_530,In_532);
and U482 (N_482,In_1202,In_155);
nand U483 (N_483,In_1109,In_134);
and U484 (N_484,In_863,In_1132);
nand U485 (N_485,In_989,In_589);
or U486 (N_486,In_935,In_1116);
nand U487 (N_487,In_524,In_229);
nor U488 (N_488,In_22,In_1238);
nand U489 (N_489,In_1491,In_1487);
or U490 (N_490,In_181,In_678);
and U491 (N_491,In_520,In_1267);
or U492 (N_492,In_236,In_1358);
nand U493 (N_493,In_1234,In_325);
nand U494 (N_494,In_886,In_152);
or U495 (N_495,In_162,In_265);
or U496 (N_496,In_545,In_218);
nand U497 (N_497,In_477,In_1419);
and U498 (N_498,In_939,In_974);
nand U499 (N_499,In_1461,In_101);
nor U500 (N_500,In_877,In_1340);
nand U501 (N_501,In_91,In_1027);
or U502 (N_502,In_1472,In_590);
nand U503 (N_503,In_1271,In_331);
or U504 (N_504,In_1299,In_446);
and U505 (N_505,In_1095,In_399);
and U506 (N_506,In_1413,In_1139);
nor U507 (N_507,In_1039,In_734);
and U508 (N_508,In_1127,In_16);
nand U509 (N_509,In_693,In_19);
nand U510 (N_510,In_1365,In_716);
nor U511 (N_511,In_1378,In_53);
nor U512 (N_512,In_79,In_688);
nand U513 (N_513,In_1189,In_1364);
or U514 (N_514,In_1452,In_1114);
xnor U515 (N_515,In_60,In_300);
and U516 (N_516,In_1023,In_1481);
nand U517 (N_517,In_283,In_1135);
and U518 (N_518,In_953,In_1071);
nor U519 (N_519,In_456,In_238);
nand U520 (N_520,In_660,In_1324);
and U521 (N_521,In_986,In_159);
nand U522 (N_522,In_314,In_798);
nor U523 (N_523,In_107,In_548);
nand U524 (N_524,In_246,In_864);
or U525 (N_525,In_425,In_353);
nor U526 (N_526,In_275,In_804);
nand U527 (N_527,In_815,In_250);
and U528 (N_528,In_1028,In_256);
and U529 (N_529,In_323,In_1066);
nor U530 (N_530,In_95,In_951);
nand U531 (N_531,In_117,In_753);
or U532 (N_532,In_923,In_701);
nor U533 (N_533,In_898,In_976);
or U534 (N_534,In_136,In_528);
nand U535 (N_535,In_5,In_1255);
nand U536 (N_536,In_782,In_559);
or U537 (N_537,In_234,In_884);
nor U538 (N_538,In_486,In_900);
and U539 (N_539,In_412,In_585);
or U540 (N_540,In_827,In_1418);
or U541 (N_541,In_774,In_1281);
nand U542 (N_542,In_1313,In_502);
nor U543 (N_543,In_1001,In_188);
or U544 (N_544,In_1425,In_230);
and U545 (N_545,In_924,In_715);
or U546 (N_546,In_748,In_852);
or U547 (N_547,In_391,In_99);
and U548 (N_548,In_909,In_368);
or U549 (N_549,In_1479,In_114);
nor U550 (N_550,In_570,In_1263);
and U551 (N_551,In_115,In_1272);
nor U552 (N_552,In_1193,In_253);
nand U553 (N_553,In_224,In_1099);
nand U554 (N_554,In_1359,In_784);
nor U555 (N_555,In_0,In_261);
or U556 (N_556,In_1336,In_702);
nor U557 (N_557,In_1274,In_1282);
or U558 (N_558,In_1171,In_137);
nand U559 (N_559,In_259,In_564);
nand U560 (N_560,In_493,In_574);
nand U561 (N_561,In_27,In_1297);
nand U562 (N_562,In_1496,In_1293);
and U563 (N_563,In_726,In_1406);
nor U564 (N_564,In_759,In_404);
or U565 (N_565,In_1038,In_588);
nand U566 (N_566,In_556,In_1262);
and U567 (N_567,In_690,In_34);
and U568 (N_568,In_666,In_742);
or U569 (N_569,In_1339,In_142);
and U570 (N_570,In_859,In_1386);
and U571 (N_571,In_1264,In_1445);
nor U572 (N_572,In_1248,In_1134);
or U573 (N_573,In_313,In_960);
nand U574 (N_574,In_167,In_1152);
nor U575 (N_575,In_1149,In_381);
and U576 (N_576,In_1317,In_1198);
or U577 (N_577,In_920,In_260);
and U578 (N_578,In_964,In_1435);
and U579 (N_579,In_772,In_463);
or U580 (N_580,In_1421,In_1047);
and U581 (N_581,In_749,In_648);
and U582 (N_582,In_1312,In_540);
and U583 (N_583,In_661,In_929);
or U584 (N_584,In_966,In_934);
and U585 (N_585,In_1069,In_837);
or U586 (N_586,In_539,In_15);
nand U587 (N_587,In_1349,In_881);
and U588 (N_588,In_436,In_1124);
nor U589 (N_589,In_1380,In_1103);
nand U590 (N_590,In_602,In_855);
and U591 (N_591,In_671,In_1216);
nor U592 (N_592,In_741,In_1374);
nor U593 (N_593,In_637,In_913);
nand U594 (N_594,In_783,In_449);
and U595 (N_595,In_55,In_1463);
nor U596 (N_596,In_379,In_385);
nand U597 (N_597,In_257,In_763);
nand U598 (N_598,In_799,In_255);
nand U599 (N_599,In_147,In_509);
nand U600 (N_600,In_1437,In_125);
nand U601 (N_601,In_948,In_1257);
and U602 (N_602,In_835,In_674);
nor U603 (N_603,In_996,In_56);
and U604 (N_604,In_971,In_1275);
or U605 (N_605,In_1045,In_623);
or U606 (N_606,In_1495,In_341);
or U607 (N_607,In_1182,In_8);
nor U608 (N_608,In_947,In_1206);
or U609 (N_609,In_1081,In_1431);
or U610 (N_610,In_1183,In_35);
nand U611 (N_611,In_507,In_370);
and U612 (N_612,In_460,In_1235);
nand U613 (N_613,In_1407,In_268);
or U614 (N_614,In_651,In_516);
nor U615 (N_615,In_1053,In_1331);
nor U616 (N_616,In_17,In_1302);
nor U617 (N_617,In_851,In_1325);
or U618 (N_618,In_680,In_10);
nor U619 (N_619,In_579,In_1392);
and U620 (N_620,In_1130,In_450);
nand U621 (N_621,In_196,In_1485);
and U622 (N_622,In_871,In_504);
nor U623 (N_623,In_1266,In_652);
xnor U624 (N_624,In_338,In_808);
and U625 (N_625,In_692,In_1);
and U626 (N_626,In_1227,In_1433);
or U627 (N_627,In_1415,In_529);
or U628 (N_628,In_1288,In_1020);
nand U629 (N_629,In_981,In_312);
or U630 (N_630,In_732,In_299);
and U631 (N_631,In_469,In_1470);
and U632 (N_632,In_400,In_1434);
nand U633 (N_633,In_830,In_601);
and U634 (N_634,In_627,In_364);
and U635 (N_635,In_482,In_252);
or U636 (N_636,In_407,In_961);
or U637 (N_637,In_1347,In_832);
nand U638 (N_638,In_39,In_72);
nor U639 (N_639,In_1473,In_435);
or U640 (N_640,In_494,In_681);
or U641 (N_641,In_567,In_576);
nor U642 (N_642,In_786,In_727);
or U643 (N_643,In_722,In_1060);
nand U644 (N_644,In_251,In_285);
and U645 (N_645,In_1022,In_161);
nand U646 (N_646,In_20,In_580);
nor U647 (N_647,In_193,In_867);
nand U648 (N_648,In_37,In_85);
or U649 (N_649,In_245,In_744);
nor U650 (N_650,In_1153,In_993);
nor U651 (N_651,In_638,In_1190);
and U652 (N_652,In_902,In_777);
and U653 (N_653,In_1346,In_525);
nor U654 (N_654,In_1249,In_1194);
nand U655 (N_655,In_180,In_77);
nand U656 (N_656,In_410,In_441);
or U657 (N_657,In_1283,In_113);
nor U658 (N_658,In_14,In_397);
or U659 (N_659,In_873,In_714);
nand U660 (N_660,In_365,In_1129);
nor U661 (N_661,In_1456,In_38);
and U662 (N_662,In_1000,In_973);
or U663 (N_663,In_1026,In_501);
and U664 (N_664,In_1253,In_1438);
nand U665 (N_665,In_791,In_879);
and U666 (N_666,In_655,In_740);
or U667 (N_667,In_1009,In_102);
nor U668 (N_668,In_457,In_135);
nor U669 (N_669,In_918,In_454);
and U670 (N_670,In_605,In_756);
nand U671 (N_671,In_1052,In_1411);
and U672 (N_672,In_376,In_876);
nand U673 (N_673,In_216,In_522);
nand U674 (N_674,In_492,In_654);
or U675 (N_675,In_1261,In_917);
or U676 (N_676,In_165,In_73);
nand U677 (N_677,In_885,In_1096);
or U678 (N_678,In_1155,In_1148);
or U679 (N_679,In_1454,In_880);
nor U680 (N_680,In_1245,In_709);
nand U681 (N_681,In_538,In_1453);
or U682 (N_682,In_1030,In_914);
and U683 (N_683,In_47,In_945);
and U684 (N_684,In_1373,In_1084);
or U685 (N_685,In_560,In_1059);
and U686 (N_686,In_1416,In_1166);
and U687 (N_687,In_505,In_373);
or U688 (N_688,In_1337,In_1330);
nand U689 (N_689,In_551,In_1388);
and U690 (N_690,In_634,In_563);
nor U691 (N_691,In_143,In_205);
and U692 (N_692,In_1440,In_127);
nand U693 (N_693,In_474,In_1429);
nand U694 (N_694,In_438,In_1412);
xnor U695 (N_695,In_402,In_179);
nor U696 (N_696,In_963,In_71);
and U697 (N_697,In_1035,In_932);
xor U698 (N_698,In_1185,In_892);
or U699 (N_699,In_1088,In_508);
or U700 (N_700,In_360,In_213);
nand U701 (N_701,In_1046,In_1167);
nand U702 (N_702,In_1427,In_228);
or U703 (N_703,In_1430,In_480);
or U704 (N_704,In_29,In_197);
xor U705 (N_705,In_296,In_306);
nand U706 (N_706,In_239,In_88);
nand U707 (N_707,In_1320,In_514);
and U708 (N_708,In_292,In_1229);
nor U709 (N_709,In_762,In_899);
or U710 (N_710,In_781,In_31);
and U711 (N_711,In_600,In_632);
and U712 (N_712,In_499,In_706);
nand U713 (N_713,In_788,In_1345);
nor U714 (N_714,In_720,In_573);
and U715 (N_715,In_555,In_1451);
or U716 (N_716,In_770,In_812);
or U717 (N_717,In_649,In_414);
nor U718 (N_718,In_1064,In_1493);
nand U719 (N_719,In_1240,In_206);
nor U720 (N_720,In_139,In_676);
nor U721 (N_721,In_232,In_1329);
or U722 (N_722,In_1180,In_290);
nor U723 (N_723,In_615,In_1162);
or U724 (N_724,In_1370,In_721);
nand U725 (N_725,In_1460,In_1119);
nor U726 (N_726,In_1079,In_1085);
and U727 (N_727,In_416,In_1002);
nand U728 (N_728,In_1439,In_949);
xnor U729 (N_729,In_1177,In_432);
nand U730 (N_730,In_675,In_440);
nand U731 (N_731,In_106,In_50);
nand U732 (N_732,In_738,In_1305);
and U733 (N_733,In_1455,In_428);
and U734 (N_734,In_422,In_30);
or U735 (N_735,In_485,In_794);
nor U736 (N_736,In_629,In_231);
nor U737 (N_737,In_1377,In_1036);
or U738 (N_738,In_444,In_657);
or U739 (N_739,In_1164,In_176);
nand U740 (N_740,In_587,In_1399);
nand U741 (N_741,In_1258,In_751);
nor U742 (N_742,In_865,In_1101);
nor U743 (N_743,In_305,In_54);
and U744 (N_744,In_787,In_354);
or U745 (N_745,In_992,In_809);
or U746 (N_746,In_109,In_131);
and U747 (N_747,In_515,In_459);
and U748 (N_748,In_930,In_1147);
or U749 (N_749,In_642,In_302);
nand U750 (N_750,In_685,In_168);
nor U751 (N_751,In_618,In_1223);
and U752 (N_752,In_664,In_591);
and U753 (N_753,In_1089,In_526);
nand U754 (N_754,In_418,In_404);
or U755 (N_755,In_127,In_941);
nor U756 (N_756,In_1161,In_974);
and U757 (N_757,In_883,In_1019);
nand U758 (N_758,In_245,In_833);
nor U759 (N_759,In_446,In_1492);
or U760 (N_760,In_159,In_958);
xnor U761 (N_761,In_39,In_1182);
and U762 (N_762,In_1299,In_53);
nor U763 (N_763,In_353,In_870);
nor U764 (N_764,In_336,In_803);
nor U765 (N_765,In_1376,In_988);
or U766 (N_766,In_295,In_1152);
nor U767 (N_767,In_605,In_1043);
or U768 (N_768,In_1365,In_521);
nand U769 (N_769,In_18,In_731);
and U770 (N_770,In_462,In_724);
or U771 (N_771,In_1107,In_1392);
nor U772 (N_772,In_1106,In_629);
or U773 (N_773,In_83,In_1442);
and U774 (N_774,In_1490,In_568);
or U775 (N_775,In_44,In_216);
and U776 (N_776,In_970,In_1223);
and U777 (N_777,In_743,In_1256);
or U778 (N_778,In_1062,In_278);
and U779 (N_779,In_1391,In_1142);
nand U780 (N_780,In_733,In_1422);
nor U781 (N_781,In_498,In_277);
and U782 (N_782,In_148,In_492);
nand U783 (N_783,In_882,In_963);
or U784 (N_784,In_962,In_995);
nand U785 (N_785,In_167,In_1336);
nand U786 (N_786,In_1073,In_997);
and U787 (N_787,In_1113,In_1406);
nand U788 (N_788,In_495,In_1321);
xor U789 (N_789,In_698,In_893);
nor U790 (N_790,In_1239,In_207);
nand U791 (N_791,In_250,In_374);
and U792 (N_792,In_345,In_1188);
and U793 (N_793,In_817,In_745);
or U794 (N_794,In_1371,In_982);
and U795 (N_795,In_1314,In_484);
nand U796 (N_796,In_126,In_1193);
and U797 (N_797,In_576,In_97);
and U798 (N_798,In_1193,In_6);
xnor U799 (N_799,In_872,In_902);
or U800 (N_800,In_345,In_726);
or U801 (N_801,In_1478,In_1058);
nor U802 (N_802,In_1290,In_1214);
nand U803 (N_803,In_87,In_257);
nor U804 (N_804,In_498,In_18);
and U805 (N_805,In_1115,In_128);
xnor U806 (N_806,In_1339,In_575);
nor U807 (N_807,In_1462,In_205);
and U808 (N_808,In_1370,In_1008);
nand U809 (N_809,In_1334,In_752);
nand U810 (N_810,In_243,In_669);
xnor U811 (N_811,In_737,In_936);
or U812 (N_812,In_1099,In_1177);
nor U813 (N_813,In_704,In_1167);
and U814 (N_814,In_620,In_739);
nand U815 (N_815,In_1328,In_1490);
and U816 (N_816,In_629,In_649);
and U817 (N_817,In_1426,In_298);
nand U818 (N_818,In_1464,In_532);
and U819 (N_819,In_1016,In_756);
nand U820 (N_820,In_970,In_10);
nor U821 (N_821,In_298,In_1498);
nor U822 (N_822,In_1250,In_839);
nand U823 (N_823,In_1002,In_1393);
nand U824 (N_824,In_1051,In_1150);
and U825 (N_825,In_1159,In_696);
or U826 (N_826,In_139,In_1047);
xnor U827 (N_827,In_1471,In_1299);
nor U828 (N_828,In_105,In_399);
nor U829 (N_829,In_376,In_516);
nand U830 (N_830,In_212,In_1089);
nor U831 (N_831,In_426,In_1422);
nor U832 (N_832,In_884,In_241);
or U833 (N_833,In_1427,In_982);
or U834 (N_834,In_901,In_786);
and U835 (N_835,In_806,In_363);
nor U836 (N_836,In_405,In_290);
nor U837 (N_837,In_884,In_496);
or U838 (N_838,In_1329,In_354);
nor U839 (N_839,In_56,In_1348);
and U840 (N_840,In_898,In_1045);
nand U841 (N_841,In_429,In_1212);
nand U842 (N_842,In_1455,In_999);
and U843 (N_843,In_1484,In_882);
nand U844 (N_844,In_158,In_342);
nand U845 (N_845,In_1149,In_756);
and U846 (N_846,In_181,In_365);
nand U847 (N_847,In_900,In_1409);
nand U848 (N_848,In_211,In_1319);
nand U849 (N_849,In_424,In_1196);
nand U850 (N_850,In_1159,In_932);
nor U851 (N_851,In_218,In_444);
nor U852 (N_852,In_1179,In_577);
or U853 (N_853,In_1045,In_1466);
or U854 (N_854,In_1429,In_1044);
nor U855 (N_855,In_414,In_132);
nor U856 (N_856,In_158,In_1045);
nor U857 (N_857,In_1322,In_932);
and U858 (N_858,In_848,In_47);
and U859 (N_859,In_169,In_1428);
nand U860 (N_860,In_1109,In_883);
nor U861 (N_861,In_976,In_889);
and U862 (N_862,In_1249,In_339);
or U863 (N_863,In_763,In_538);
nor U864 (N_864,In_1493,In_287);
nand U865 (N_865,In_881,In_342);
and U866 (N_866,In_1206,In_1298);
and U867 (N_867,In_108,In_1314);
nor U868 (N_868,In_1339,In_815);
or U869 (N_869,In_1330,In_134);
or U870 (N_870,In_646,In_1315);
and U871 (N_871,In_57,In_125);
and U872 (N_872,In_29,In_1176);
nor U873 (N_873,In_1083,In_1457);
and U874 (N_874,In_31,In_132);
nor U875 (N_875,In_401,In_625);
nand U876 (N_876,In_310,In_1074);
nor U877 (N_877,In_424,In_1364);
or U878 (N_878,In_1172,In_1176);
nor U879 (N_879,In_1197,In_895);
nor U880 (N_880,In_1361,In_1271);
and U881 (N_881,In_1353,In_1);
nor U882 (N_882,In_799,In_649);
nor U883 (N_883,In_1107,In_1127);
nor U884 (N_884,In_1030,In_652);
xnor U885 (N_885,In_862,In_449);
nand U886 (N_886,In_1102,In_389);
nor U887 (N_887,In_523,In_490);
and U888 (N_888,In_675,In_106);
or U889 (N_889,In_778,In_321);
and U890 (N_890,In_1144,In_192);
or U891 (N_891,In_1051,In_1168);
nor U892 (N_892,In_939,In_1302);
nor U893 (N_893,In_249,In_1027);
nor U894 (N_894,In_1439,In_254);
nand U895 (N_895,In_62,In_694);
nor U896 (N_896,In_1274,In_837);
or U897 (N_897,In_1173,In_690);
and U898 (N_898,In_1339,In_5);
and U899 (N_899,In_1206,In_960);
and U900 (N_900,In_173,In_277);
nor U901 (N_901,In_343,In_11);
nor U902 (N_902,In_220,In_1259);
or U903 (N_903,In_910,In_931);
and U904 (N_904,In_307,In_1448);
nor U905 (N_905,In_1416,In_134);
nor U906 (N_906,In_1197,In_1020);
or U907 (N_907,In_203,In_1411);
or U908 (N_908,In_1407,In_1222);
or U909 (N_909,In_1347,In_655);
nor U910 (N_910,In_946,In_48);
and U911 (N_911,In_942,In_468);
or U912 (N_912,In_602,In_532);
and U913 (N_913,In_321,In_889);
nor U914 (N_914,In_97,In_727);
or U915 (N_915,In_1246,In_27);
and U916 (N_916,In_202,In_1050);
and U917 (N_917,In_738,In_453);
or U918 (N_918,In_16,In_905);
nor U919 (N_919,In_982,In_1051);
and U920 (N_920,In_1067,In_813);
or U921 (N_921,In_1031,In_1491);
nor U922 (N_922,In_118,In_111);
nor U923 (N_923,In_242,In_1427);
or U924 (N_924,In_353,In_458);
nand U925 (N_925,In_1449,In_1440);
nor U926 (N_926,In_1273,In_1007);
or U927 (N_927,In_1030,In_400);
or U928 (N_928,In_569,In_756);
and U929 (N_929,In_211,In_492);
nand U930 (N_930,In_873,In_1158);
nor U931 (N_931,In_1064,In_1011);
nand U932 (N_932,In_1354,In_774);
nand U933 (N_933,In_1105,In_125);
or U934 (N_934,In_1419,In_728);
or U935 (N_935,In_836,In_1021);
and U936 (N_936,In_319,In_163);
nor U937 (N_937,In_707,In_711);
or U938 (N_938,In_1008,In_371);
nor U939 (N_939,In_939,In_1291);
or U940 (N_940,In_1066,In_152);
or U941 (N_941,In_1445,In_542);
nand U942 (N_942,In_188,In_177);
or U943 (N_943,In_525,In_67);
and U944 (N_944,In_1296,In_745);
and U945 (N_945,In_64,In_427);
nand U946 (N_946,In_1494,In_862);
or U947 (N_947,In_1048,In_1046);
and U948 (N_948,In_399,In_637);
nand U949 (N_949,In_1465,In_1187);
nor U950 (N_950,In_940,In_759);
and U951 (N_951,In_22,In_497);
and U952 (N_952,In_732,In_916);
and U953 (N_953,In_559,In_1160);
and U954 (N_954,In_597,In_1365);
nor U955 (N_955,In_941,In_1219);
nor U956 (N_956,In_693,In_357);
or U957 (N_957,In_1153,In_1066);
nor U958 (N_958,In_68,In_1431);
or U959 (N_959,In_1322,In_475);
and U960 (N_960,In_624,In_540);
or U961 (N_961,In_1374,In_504);
nor U962 (N_962,In_993,In_892);
nor U963 (N_963,In_374,In_39);
xor U964 (N_964,In_611,In_255);
nand U965 (N_965,In_1235,In_156);
nor U966 (N_966,In_239,In_621);
nor U967 (N_967,In_1111,In_259);
nor U968 (N_968,In_909,In_1035);
nor U969 (N_969,In_718,In_817);
or U970 (N_970,In_1321,In_182);
nand U971 (N_971,In_142,In_471);
nand U972 (N_972,In_1211,In_390);
nand U973 (N_973,In_835,In_356);
and U974 (N_974,In_1256,In_647);
and U975 (N_975,In_387,In_572);
and U976 (N_976,In_344,In_920);
or U977 (N_977,In_1455,In_1469);
nand U978 (N_978,In_983,In_217);
or U979 (N_979,In_1223,In_1471);
or U980 (N_980,In_1305,In_256);
nand U981 (N_981,In_1062,In_93);
and U982 (N_982,In_953,In_1321);
nand U983 (N_983,In_415,In_715);
or U984 (N_984,In_944,In_756);
nor U985 (N_985,In_732,In_1058);
or U986 (N_986,In_20,In_157);
or U987 (N_987,In_120,In_166);
nor U988 (N_988,In_1258,In_1171);
nor U989 (N_989,In_796,In_1240);
and U990 (N_990,In_707,In_872);
nand U991 (N_991,In_996,In_898);
xor U992 (N_992,In_611,In_1235);
nor U993 (N_993,In_12,In_79);
nand U994 (N_994,In_74,In_2);
nor U995 (N_995,In_235,In_99);
or U996 (N_996,In_1006,In_370);
nand U997 (N_997,In_783,In_1109);
or U998 (N_998,In_452,In_295);
nor U999 (N_999,In_1233,In_814);
xor U1000 (N_1000,In_41,In_121);
and U1001 (N_1001,In_703,In_853);
and U1002 (N_1002,In_274,In_1206);
nand U1003 (N_1003,In_5,In_512);
or U1004 (N_1004,In_20,In_1040);
nand U1005 (N_1005,In_249,In_206);
or U1006 (N_1006,In_897,In_936);
nand U1007 (N_1007,In_490,In_1130);
or U1008 (N_1008,In_815,In_773);
nand U1009 (N_1009,In_1049,In_1428);
nand U1010 (N_1010,In_843,In_371);
or U1011 (N_1011,In_1343,In_1104);
or U1012 (N_1012,In_517,In_368);
nand U1013 (N_1013,In_204,In_179);
nor U1014 (N_1014,In_356,In_754);
and U1015 (N_1015,In_1305,In_1493);
nor U1016 (N_1016,In_1390,In_1331);
or U1017 (N_1017,In_1429,In_24);
or U1018 (N_1018,In_272,In_936);
and U1019 (N_1019,In_3,In_589);
nand U1020 (N_1020,In_984,In_665);
nor U1021 (N_1021,In_554,In_462);
nand U1022 (N_1022,In_522,In_530);
nor U1023 (N_1023,In_1165,In_531);
nor U1024 (N_1024,In_315,In_225);
nand U1025 (N_1025,In_243,In_505);
nor U1026 (N_1026,In_1312,In_22);
nor U1027 (N_1027,In_1473,In_1421);
or U1028 (N_1028,In_862,In_352);
nand U1029 (N_1029,In_247,In_110);
and U1030 (N_1030,In_832,In_84);
or U1031 (N_1031,In_901,In_133);
and U1032 (N_1032,In_1146,In_351);
nor U1033 (N_1033,In_1389,In_1166);
or U1034 (N_1034,In_1267,In_1020);
nand U1035 (N_1035,In_758,In_380);
and U1036 (N_1036,In_1204,In_1227);
nor U1037 (N_1037,In_1443,In_1457);
nor U1038 (N_1038,In_829,In_658);
or U1039 (N_1039,In_1206,In_433);
or U1040 (N_1040,In_1270,In_44);
or U1041 (N_1041,In_820,In_1232);
or U1042 (N_1042,In_1315,In_455);
nor U1043 (N_1043,In_265,In_1138);
and U1044 (N_1044,In_1172,In_139);
nor U1045 (N_1045,In_1330,In_883);
nand U1046 (N_1046,In_1489,In_215);
xor U1047 (N_1047,In_1045,In_1258);
nand U1048 (N_1048,In_718,In_1125);
and U1049 (N_1049,In_1497,In_1250);
and U1050 (N_1050,In_960,In_689);
or U1051 (N_1051,In_1476,In_833);
nor U1052 (N_1052,In_1170,In_1488);
or U1053 (N_1053,In_507,In_477);
nor U1054 (N_1054,In_217,In_329);
and U1055 (N_1055,In_616,In_106);
and U1056 (N_1056,In_943,In_689);
nor U1057 (N_1057,In_286,In_1452);
nand U1058 (N_1058,In_604,In_622);
nor U1059 (N_1059,In_1403,In_1073);
and U1060 (N_1060,In_1124,In_1247);
nor U1061 (N_1061,In_384,In_725);
or U1062 (N_1062,In_874,In_335);
nor U1063 (N_1063,In_699,In_1358);
nand U1064 (N_1064,In_974,In_1142);
or U1065 (N_1065,In_1156,In_76);
and U1066 (N_1066,In_1190,In_1116);
or U1067 (N_1067,In_71,In_709);
and U1068 (N_1068,In_943,In_1297);
nor U1069 (N_1069,In_1090,In_1054);
nor U1070 (N_1070,In_195,In_518);
or U1071 (N_1071,In_114,In_689);
or U1072 (N_1072,In_70,In_294);
and U1073 (N_1073,In_1161,In_414);
nand U1074 (N_1074,In_20,In_994);
xnor U1075 (N_1075,In_680,In_111);
nor U1076 (N_1076,In_842,In_5);
or U1077 (N_1077,In_218,In_1150);
and U1078 (N_1078,In_737,In_516);
nor U1079 (N_1079,In_423,In_716);
nor U1080 (N_1080,In_83,In_733);
or U1081 (N_1081,In_1453,In_447);
nor U1082 (N_1082,In_823,In_217);
nor U1083 (N_1083,In_594,In_392);
xnor U1084 (N_1084,In_890,In_164);
nand U1085 (N_1085,In_1427,In_1015);
or U1086 (N_1086,In_557,In_962);
nor U1087 (N_1087,In_127,In_1229);
nor U1088 (N_1088,In_611,In_999);
nand U1089 (N_1089,In_4,In_779);
nand U1090 (N_1090,In_409,In_248);
and U1091 (N_1091,In_1332,In_1415);
or U1092 (N_1092,In_1183,In_1381);
nor U1093 (N_1093,In_162,In_620);
nand U1094 (N_1094,In_483,In_1147);
nor U1095 (N_1095,In_484,In_495);
or U1096 (N_1096,In_1002,In_443);
nor U1097 (N_1097,In_1065,In_696);
or U1098 (N_1098,In_736,In_1244);
or U1099 (N_1099,In_882,In_935);
xnor U1100 (N_1100,In_68,In_118);
nand U1101 (N_1101,In_600,In_776);
nand U1102 (N_1102,In_1206,In_899);
or U1103 (N_1103,In_1336,In_703);
nor U1104 (N_1104,In_270,In_1252);
nand U1105 (N_1105,In_431,In_101);
nand U1106 (N_1106,In_689,In_946);
nor U1107 (N_1107,In_68,In_641);
or U1108 (N_1108,In_1053,In_951);
and U1109 (N_1109,In_292,In_545);
and U1110 (N_1110,In_1239,In_355);
xor U1111 (N_1111,In_1043,In_582);
or U1112 (N_1112,In_66,In_725);
nor U1113 (N_1113,In_974,In_990);
nand U1114 (N_1114,In_27,In_1391);
nand U1115 (N_1115,In_832,In_530);
nand U1116 (N_1116,In_1048,In_219);
nand U1117 (N_1117,In_242,In_1304);
nand U1118 (N_1118,In_1382,In_587);
nand U1119 (N_1119,In_576,In_811);
nand U1120 (N_1120,In_528,In_1399);
nor U1121 (N_1121,In_351,In_1210);
nor U1122 (N_1122,In_1298,In_1153);
nor U1123 (N_1123,In_1168,In_822);
or U1124 (N_1124,In_205,In_172);
nand U1125 (N_1125,In_123,In_144);
nand U1126 (N_1126,In_1429,In_274);
nor U1127 (N_1127,In_241,In_1175);
and U1128 (N_1128,In_1152,In_195);
or U1129 (N_1129,In_682,In_1472);
nor U1130 (N_1130,In_195,In_1046);
nand U1131 (N_1131,In_370,In_136);
nand U1132 (N_1132,In_639,In_664);
nor U1133 (N_1133,In_1140,In_696);
or U1134 (N_1134,In_232,In_819);
nor U1135 (N_1135,In_503,In_123);
and U1136 (N_1136,In_618,In_550);
or U1137 (N_1137,In_669,In_1497);
and U1138 (N_1138,In_1358,In_191);
and U1139 (N_1139,In_643,In_714);
nor U1140 (N_1140,In_693,In_723);
xor U1141 (N_1141,In_1486,In_1171);
nand U1142 (N_1142,In_226,In_341);
and U1143 (N_1143,In_701,In_1007);
nand U1144 (N_1144,In_851,In_248);
nor U1145 (N_1145,In_240,In_135);
nand U1146 (N_1146,In_7,In_136);
or U1147 (N_1147,In_866,In_1387);
nand U1148 (N_1148,In_743,In_637);
xnor U1149 (N_1149,In_1389,In_1112);
and U1150 (N_1150,In_87,In_320);
nor U1151 (N_1151,In_1153,In_280);
and U1152 (N_1152,In_1190,In_977);
nand U1153 (N_1153,In_1220,In_769);
and U1154 (N_1154,In_127,In_163);
nand U1155 (N_1155,In_295,In_1383);
and U1156 (N_1156,In_1179,In_1170);
or U1157 (N_1157,In_635,In_866);
nand U1158 (N_1158,In_1212,In_780);
or U1159 (N_1159,In_1161,In_650);
nand U1160 (N_1160,In_1352,In_1133);
or U1161 (N_1161,In_335,In_1111);
and U1162 (N_1162,In_1083,In_953);
and U1163 (N_1163,In_597,In_62);
and U1164 (N_1164,In_924,In_267);
and U1165 (N_1165,In_1477,In_527);
nor U1166 (N_1166,In_542,In_391);
nand U1167 (N_1167,In_1417,In_1329);
xnor U1168 (N_1168,In_1192,In_552);
and U1169 (N_1169,In_434,In_1194);
nor U1170 (N_1170,In_255,In_1213);
and U1171 (N_1171,In_1033,In_1283);
or U1172 (N_1172,In_1239,In_1335);
or U1173 (N_1173,In_954,In_594);
or U1174 (N_1174,In_812,In_232);
nand U1175 (N_1175,In_1357,In_648);
nand U1176 (N_1176,In_122,In_14);
nor U1177 (N_1177,In_150,In_631);
and U1178 (N_1178,In_1423,In_586);
and U1179 (N_1179,In_115,In_926);
or U1180 (N_1180,In_112,In_1443);
or U1181 (N_1181,In_1248,In_219);
and U1182 (N_1182,In_119,In_1258);
nand U1183 (N_1183,In_923,In_567);
nand U1184 (N_1184,In_296,In_890);
and U1185 (N_1185,In_754,In_116);
and U1186 (N_1186,In_1072,In_793);
or U1187 (N_1187,In_1187,In_205);
nor U1188 (N_1188,In_780,In_1226);
or U1189 (N_1189,In_1357,In_1464);
nor U1190 (N_1190,In_796,In_482);
and U1191 (N_1191,In_1251,In_1294);
and U1192 (N_1192,In_542,In_196);
nand U1193 (N_1193,In_686,In_31);
nand U1194 (N_1194,In_229,In_266);
nor U1195 (N_1195,In_1103,In_14);
xnor U1196 (N_1196,In_842,In_854);
or U1197 (N_1197,In_1227,In_1225);
nor U1198 (N_1198,In_1425,In_1396);
nand U1199 (N_1199,In_629,In_1480);
or U1200 (N_1200,In_1143,In_510);
or U1201 (N_1201,In_1172,In_523);
or U1202 (N_1202,In_168,In_692);
and U1203 (N_1203,In_673,In_559);
and U1204 (N_1204,In_1154,In_733);
or U1205 (N_1205,In_1315,In_1317);
nand U1206 (N_1206,In_569,In_904);
nand U1207 (N_1207,In_113,In_127);
and U1208 (N_1208,In_1172,In_554);
nand U1209 (N_1209,In_14,In_1109);
nand U1210 (N_1210,In_500,In_648);
nor U1211 (N_1211,In_666,In_1078);
and U1212 (N_1212,In_184,In_508);
or U1213 (N_1213,In_33,In_381);
nor U1214 (N_1214,In_1457,In_356);
xnor U1215 (N_1215,In_213,In_707);
and U1216 (N_1216,In_1095,In_1067);
nor U1217 (N_1217,In_490,In_1398);
nand U1218 (N_1218,In_586,In_1206);
nand U1219 (N_1219,In_929,In_867);
and U1220 (N_1220,In_638,In_561);
nor U1221 (N_1221,In_565,In_61);
nor U1222 (N_1222,In_1055,In_1386);
nor U1223 (N_1223,In_644,In_96);
nand U1224 (N_1224,In_940,In_756);
nor U1225 (N_1225,In_1229,In_545);
or U1226 (N_1226,In_1491,In_883);
nor U1227 (N_1227,In_1205,In_1332);
or U1228 (N_1228,In_383,In_517);
and U1229 (N_1229,In_953,In_1227);
xnor U1230 (N_1230,In_1397,In_582);
or U1231 (N_1231,In_973,In_749);
nand U1232 (N_1232,In_1202,In_272);
and U1233 (N_1233,In_238,In_764);
and U1234 (N_1234,In_1228,In_1102);
and U1235 (N_1235,In_223,In_1380);
nor U1236 (N_1236,In_716,In_137);
nor U1237 (N_1237,In_1310,In_1007);
nor U1238 (N_1238,In_65,In_537);
and U1239 (N_1239,In_1449,In_914);
or U1240 (N_1240,In_1293,In_561);
or U1241 (N_1241,In_664,In_759);
and U1242 (N_1242,In_831,In_1097);
or U1243 (N_1243,In_1216,In_828);
or U1244 (N_1244,In_177,In_1139);
nor U1245 (N_1245,In_282,In_685);
or U1246 (N_1246,In_140,In_1265);
and U1247 (N_1247,In_955,In_787);
or U1248 (N_1248,In_688,In_343);
nand U1249 (N_1249,In_4,In_601);
nor U1250 (N_1250,In_1381,In_1181);
nor U1251 (N_1251,In_1287,In_838);
nand U1252 (N_1252,In_989,In_905);
nand U1253 (N_1253,In_442,In_1067);
or U1254 (N_1254,In_491,In_1452);
nand U1255 (N_1255,In_446,In_906);
or U1256 (N_1256,In_457,In_126);
and U1257 (N_1257,In_653,In_802);
nor U1258 (N_1258,In_1211,In_194);
nand U1259 (N_1259,In_891,In_119);
and U1260 (N_1260,In_132,In_144);
or U1261 (N_1261,In_755,In_48);
or U1262 (N_1262,In_411,In_1096);
nor U1263 (N_1263,In_1473,In_1320);
and U1264 (N_1264,In_806,In_730);
nand U1265 (N_1265,In_400,In_489);
nand U1266 (N_1266,In_1408,In_604);
nand U1267 (N_1267,In_999,In_629);
or U1268 (N_1268,In_880,In_1014);
nand U1269 (N_1269,In_363,In_489);
xnor U1270 (N_1270,In_1120,In_381);
nor U1271 (N_1271,In_1002,In_1432);
and U1272 (N_1272,In_552,In_562);
or U1273 (N_1273,In_534,In_1351);
or U1274 (N_1274,In_721,In_300);
or U1275 (N_1275,In_886,In_312);
nand U1276 (N_1276,In_524,In_881);
and U1277 (N_1277,In_481,In_1057);
or U1278 (N_1278,In_1446,In_49);
nand U1279 (N_1279,In_1120,In_429);
nand U1280 (N_1280,In_1461,In_275);
nand U1281 (N_1281,In_202,In_1262);
and U1282 (N_1282,In_1361,In_473);
and U1283 (N_1283,In_1340,In_461);
and U1284 (N_1284,In_1187,In_1396);
nor U1285 (N_1285,In_449,In_731);
or U1286 (N_1286,In_642,In_1161);
nand U1287 (N_1287,In_420,In_325);
or U1288 (N_1288,In_53,In_1476);
or U1289 (N_1289,In_335,In_1342);
nand U1290 (N_1290,In_93,In_680);
and U1291 (N_1291,In_1209,In_687);
or U1292 (N_1292,In_452,In_198);
or U1293 (N_1293,In_1190,In_1);
xnor U1294 (N_1294,In_114,In_997);
and U1295 (N_1295,In_1124,In_1424);
nand U1296 (N_1296,In_505,In_896);
and U1297 (N_1297,In_171,In_479);
and U1298 (N_1298,In_810,In_368);
nor U1299 (N_1299,In_1241,In_908);
nand U1300 (N_1300,In_835,In_1090);
nor U1301 (N_1301,In_814,In_1220);
or U1302 (N_1302,In_1272,In_1126);
and U1303 (N_1303,In_172,In_299);
or U1304 (N_1304,In_1101,In_551);
nor U1305 (N_1305,In_557,In_36);
nand U1306 (N_1306,In_444,In_394);
and U1307 (N_1307,In_897,In_778);
or U1308 (N_1308,In_847,In_1080);
and U1309 (N_1309,In_213,In_987);
nor U1310 (N_1310,In_1313,In_214);
and U1311 (N_1311,In_339,In_1333);
and U1312 (N_1312,In_1319,In_1030);
nand U1313 (N_1313,In_1184,In_375);
or U1314 (N_1314,In_1218,In_1192);
nand U1315 (N_1315,In_1117,In_1066);
or U1316 (N_1316,In_906,In_219);
nor U1317 (N_1317,In_66,In_793);
or U1318 (N_1318,In_307,In_210);
or U1319 (N_1319,In_263,In_1290);
and U1320 (N_1320,In_165,In_989);
or U1321 (N_1321,In_453,In_354);
and U1322 (N_1322,In_834,In_799);
and U1323 (N_1323,In_826,In_1079);
nor U1324 (N_1324,In_793,In_1027);
or U1325 (N_1325,In_1339,In_1152);
nor U1326 (N_1326,In_1266,In_538);
nand U1327 (N_1327,In_432,In_306);
nand U1328 (N_1328,In_253,In_494);
nor U1329 (N_1329,In_1221,In_817);
nand U1330 (N_1330,In_1110,In_499);
and U1331 (N_1331,In_430,In_1432);
or U1332 (N_1332,In_575,In_731);
nand U1333 (N_1333,In_1202,In_1197);
and U1334 (N_1334,In_1064,In_317);
nand U1335 (N_1335,In_1444,In_1107);
xnor U1336 (N_1336,In_740,In_1291);
nor U1337 (N_1337,In_537,In_479);
or U1338 (N_1338,In_327,In_481);
nand U1339 (N_1339,In_1182,In_1314);
or U1340 (N_1340,In_526,In_412);
nand U1341 (N_1341,In_600,In_1291);
or U1342 (N_1342,In_61,In_596);
nand U1343 (N_1343,In_1222,In_86);
nand U1344 (N_1344,In_993,In_339);
or U1345 (N_1345,In_651,In_559);
and U1346 (N_1346,In_802,In_1321);
and U1347 (N_1347,In_341,In_757);
and U1348 (N_1348,In_409,In_1240);
and U1349 (N_1349,In_1194,In_1196);
nand U1350 (N_1350,In_1160,In_883);
or U1351 (N_1351,In_717,In_1145);
nor U1352 (N_1352,In_1048,In_776);
nor U1353 (N_1353,In_507,In_1308);
or U1354 (N_1354,In_166,In_528);
or U1355 (N_1355,In_460,In_461);
or U1356 (N_1356,In_994,In_573);
or U1357 (N_1357,In_1027,In_1225);
xor U1358 (N_1358,In_1408,In_248);
nor U1359 (N_1359,In_399,In_495);
nand U1360 (N_1360,In_109,In_47);
nand U1361 (N_1361,In_326,In_1313);
or U1362 (N_1362,In_684,In_610);
and U1363 (N_1363,In_731,In_698);
and U1364 (N_1364,In_72,In_569);
or U1365 (N_1365,In_268,In_339);
or U1366 (N_1366,In_1391,In_331);
nor U1367 (N_1367,In_1200,In_1462);
nand U1368 (N_1368,In_664,In_406);
nor U1369 (N_1369,In_455,In_192);
and U1370 (N_1370,In_528,In_79);
or U1371 (N_1371,In_772,In_910);
or U1372 (N_1372,In_1392,In_272);
or U1373 (N_1373,In_781,In_635);
nor U1374 (N_1374,In_1096,In_4);
nand U1375 (N_1375,In_601,In_908);
or U1376 (N_1376,In_191,In_491);
and U1377 (N_1377,In_501,In_1465);
and U1378 (N_1378,In_1283,In_1173);
nor U1379 (N_1379,In_1457,In_1390);
nor U1380 (N_1380,In_1049,In_254);
or U1381 (N_1381,In_195,In_1195);
xor U1382 (N_1382,In_893,In_1099);
nor U1383 (N_1383,In_1429,In_366);
or U1384 (N_1384,In_491,In_1039);
and U1385 (N_1385,In_1465,In_1310);
nand U1386 (N_1386,In_1254,In_1000);
nand U1387 (N_1387,In_908,In_1186);
nand U1388 (N_1388,In_1038,In_368);
nand U1389 (N_1389,In_1039,In_351);
nor U1390 (N_1390,In_345,In_236);
and U1391 (N_1391,In_125,In_1350);
and U1392 (N_1392,In_1222,In_1176);
nand U1393 (N_1393,In_749,In_17);
nor U1394 (N_1394,In_1299,In_1172);
or U1395 (N_1395,In_502,In_884);
nor U1396 (N_1396,In_1176,In_247);
or U1397 (N_1397,In_1330,In_903);
and U1398 (N_1398,In_821,In_1309);
nand U1399 (N_1399,In_59,In_1161);
or U1400 (N_1400,In_901,In_1062);
nand U1401 (N_1401,In_682,In_147);
nor U1402 (N_1402,In_678,In_167);
nor U1403 (N_1403,In_1362,In_1374);
nor U1404 (N_1404,In_407,In_1396);
nand U1405 (N_1405,In_594,In_1394);
xor U1406 (N_1406,In_877,In_1413);
or U1407 (N_1407,In_91,In_281);
and U1408 (N_1408,In_99,In_37);
and U1409 (N_1409,In_1326,In_1222);
and U1410 (N_1410,In_552,In_814);
nor U1411 (N_1411,In_1456,In_1317);
and U1412 (N_1412,In_1072,In_1208);
and U1413 (N_1413,In_177,In_80);
or U1414 (N_1414,In_1080,In_348);
nand U1415 (N_1415,In_175,In_326);
nor U1416 (N_1416,In_1416,In_208);
or U1417 (N_1417,In_1213,In_1139);
nand U1418 (N_1418,In_286,In_154);
nor U1419 (N_1419,In_1348,In_1403);
and U1420 (N_1420,In_38,In_581);
nand U1421 (N_1421,In_1223,In_1057);
nand U1422 (N_1422,In_946,In_679);
or U1423 (N_1423,In_1250,In_365);
nor U1424 (N_1424,In_1480,In_809);
xnor U1425 (N_1425,In_1370,In_307);
nand U1426 (N_1426,In_596,In_776);
or U1427 (N_1427,In_806,In_479);
nor U1428 (N_1428,In_688,In_663);
nor U1429 (N_1429,In_447,In_1495);
or U1430 (N_1430,In_39,In_357);
or U1431 (N_1431,In_176,In_1231);
nand U1432 (N_1432,In_773,In_253);
nor U1433 (N_1433,In_854,In_1150);
nand U1434 (N_1434,In_621,In_1482);
or U1435 (N_1435,In_353,In_1187);
nand U1436 (N_1436,In_26,In_1212);
nand U1437 (N_1437,In_424,In_948);
xnor U1438 (N_1438,In_559,In_1236);
nor U1439 (N_1439,In_1220,In_1000);
and U1440 (N_1440,In_951,In_595);
or U1441 (N_1441,In_221,In_890);
and U1442 (N_1442,In_903,In_327);
or U1443 (N_1443,In_320,In_941);
nand U1444 (N_1444,In_724,In_68);
or U1445 (N_1445,In_1493,In_617);
and U1446 (N_1446,In_458,In_1354);
or U1447 (N_1447,In_907,In_1399);
and U1448 (N_1448,In_186,In_85);
nor U1449 (N_1449,In_303,In_325);
nor U1450 (N_1450,In_1004,In_974);
and U1451 (N_1451,In_312,In_1468);
or U1452 (N_1452,In_987,In_771);
nand U1453 (N_1453,In_1146,In_744);
or U1454 (N_1454,In_1271,In_921);
or U1455 (N_1455,In_500,In_269);
and U1456 (N_1456,In_620,In_220);
and U1457 (N_1457,In_839,In_1000);
nor U1458 (N_1458,In_188,In_519);
xnor U1459 (N_1459,In_1363,In_1332);
or U1460 (N_1460,In_1396,In_206);
nor U1461 (N_1461,In_273,In_179);
nor U1462 (N_1462,In_246,In_1098);
and U1463 (N_1463,In_269,In_50);
nand U1464 (N_1464,In_303,In_1161);
nand U1465 (N_1465,In_382,In_507);
nor U1466 (N_1466,In_534,In_812);
nand U1467 (N_1467,In_1106,In_43);
nand U1468 (N_1468,In_125,In_1287);
and U1469 (N_1469,In_789,In_663);
or U1470 (N_1470,In_1078,In_1445);
nor U1471 (N_1471,In_652,In_69);
or U1472 (N_1472,In_290,In_1068);
or U1473 (N_1473,In_479,In_540);
nand U1474 (N_1474,In_867,In_1231);
or U1475 (N_1475,In_284,In_175);
or U1476 (N_1476,In_1069,In_923);
or U1477 (N_1477,In_93,In_288);
nor U1478 (N_1478,In_77,In_1005);
nand U1479 (N_1479,In_270,In_1302);
or U1480 (N_1480,In_1275,In_289);
xor U1481 (N_1481,In_1020,In_18);
or U1482 (N_1482,In_716,In_96);
or U1483 (N_1483,In_1112,In_788);
nor U1484 (N_1484,In_584,In_1097);
xor U1485 (N_1485,In_1016,In_1103);
and U1486 (N_1486,In_1268,In_1031);
and U1487 (N_1487,In_593,In_320);
nand U1488 (N_1488,In_825,In_569);
nand U1489 (N_1489,In_1083,In_1331);
nor U1490 (N_1490,In_646,In_911);
nor U1491 (N_1491,In_1135,In_512);
nand U1492 (N_1492,In_370,In_1324);
nand U1493 (N_1493,In_675,In_1228);
nor U1494 (N_1494,In_1320,In_1435);
nand U1495 (N_1495,In_666,In_420);
or U1496 (N_1496,In_253,In_1038);
and U1497 (N_1497,In_122,In_744);
nor U1498 (N_1498,In_1162,In_571);
nand U1499 (N_1499,In_1425,In_1329);
or U1500 (N_1500,N_1473,N_185);
or U1501 (N_1501,N_787,N_567);
or U1502 (N_1502,N_773,N_1417);
and U1503 (N_1503,N_777,N_1028);
nand U1504 (N_1504,N_476,N_436);
and U1505 (N_1505,N_848,N_130);
and U1506 (N_1506,N_232,N_7);
and U1507 (N_1507,N_393,N_1057);
nand U1508 (N_1508,N_702,N_122);
or U1509 (N_1509,N_499,N_1455);
nand U1510 (N_1510,N_779,N_1405);
and U1511 (N_1511,N_263,N_1182);
and U1512 (N_1512,N_139,N_798);
or U1513 (N_1513,N_1420,N_886);
or U1514 (N_1514,N_1226,N_656);
nor U1515 (N_1515,N_233,N_547);
or U1516 (N_1516,N_754,N_218);
and U1517 (N_1517,N_936,N_1498);
nor U1518 (N_1518,N_181,N_343);
and U1519 (N_1519,N_831,N_1428);
or U1520 (N_1520,N_178,N_76);
nand U1521 (N_1521,N_1131,N_1499);
nor U1522 (N_1522,N_960,N_1221);
and U1523 (N_1523,N_387,N_266);
and U1524 (N_1524,N_316,N_138);
or U1525 (N_1525,N_160,N_1042);
and U1526 (N_1526,N_549,N_957);
and U1527 (N_1527,N_1059,N_1462);
nand U1528 (N_1528,N_1483,N_1084);
nand U1529 (N_1529,N_850,N_448);
or U1530 (N_1530,N_261,N_764);
nor U1531 (N_1531,N_906,N_1312);
nor U1532 (N_1532,N_1010,N_134);
and U1533 (N_1533,N_1271,N_257);
and U1534 (N_1534,N_362,N_1393);
nand U1535 (N_1535,N_370,N_1295);
nor U1536 (N_1536,N_125,N_718);
and U1537 (N_1537,N_518,N_1021);
or U1538 (N_1538,N_962,N_98);
nor U1539 (N_1539,N_1469,N_827);
or U1540 (N_1540,N_509,N_1032);
or U1541 (N_1541,N_825,N_398);
nor U1542 (N_1542,N_673,N_482);
or U1543 (N_1543,N_841,N_1470);
and U1544 (N_1544,N_1305,N_1381);
or U1545 (N_1545,N_33,N_483);
and U1546 (N_1546,N_103,N_378);
and U1547 (N_1547,N_692,N_96);
or U1548 (N_1548,N_1121,N_1164);
or U1549 (N_1549,N_1110,N_124);
nand U1550 (N_1550,N_585,N_81);
nor U1551 (N_1551,N_1245,N_516);
xnor U1552 (N_1552,N_657,N_437);
or U1553 (N_1553,N_756,N_438);
and U1554 (N_1554,N_872,N_965);
nor U1555 (N_1555,N_1339,N_87);
nor U1556 (N_1556,N_1460,N_1017);
or U1557 (N_1557,N_180,N_268);
or U1558 (N_1558,N_1457,N_1387);
nor U1559 (N_1559,N_1297,N_898);
and U1560 (N_1560,N_220,N_15);
and U1561 (N_1561,N_1426,N_1014);
xnor U1562 (N_1562,N_128,N_341);
nand U1563 (N_1563,N_915,N_1015);
nand U1564 (N_1564,N_1187,N_1119);
xnor U1565 (N_1565,N_1256,N_586);
nand U1566 (N_1566,N_56,N_1061);
and U1567 (N_1567,N_633,N_1421);
nand U1568 (N_1568,N_135,N_1442);
or U1569 (N_1569,N_1168,N_302);
or U1570 (N_1570,N_857,N_1482);
nand U1571 (N_1571,N_1434,N_1128);
nand U1572 (N_1572,N_276,N_1214);
or U1573 (N_1573,N_59,N_861);
nand U1574 (N_1574,N_1094,N_496);
or U1575 (N_1575,N_750,N_1325);
nor U1576 (N_1576,N_1103,N_1144);
nor U1577 (N_1577,N_802,N_1250);
and U1578 (N_1578,N_819,N_1415);
nand U1579 (N_1579,N_522,N_838);
and U1580 (N_1580,N_293,N_259);
nand U1581 (N_1581,N_104,N_769);
or U1582 (N_1582,N_623,N_752);
nand U1583 (N_1583,N_1461,N_654);
nand U1584 (N_1584,N_1396,N_1464);
nor U1585 (N_1585,N_258,N_1353);
or U1586 (N_1586,N_94,N_315);
or U1587 (N_1587,N_1324,N_666);
or U1588 (N_1588,N_205,N_412);
nor U1589 (N_1589,N_1326,N_1006);
nand U1590 (N_1590,N_198,N_118);
nor U1591 (N_1591,N_305,N_71);
nor U1592 (N_1592,N_1279,N_1019);
or U1593 (N_1593,N_369,N_294);
or U1594 (N_1594,N_597,N_588);
nor U1595 (N_1595,N_53,N_368);
nor U1596 (N_1596,N_16,N_735);
or U1597 (N_1597,N_1120,N_469);
nand U1598 (N_1598,N_93,N_431);
or U1599 (N_1599,N_176,N_1292);
or U1600 (N_1600,N_373,N_274);
or U1601 (N_1601,N_870,N_703);
or U1602 (N_1602,N_1441,N_256);
nor U1603 (N_1603,N_35,N_515);
and U1604 (N_1604,N_760,N_574);
and U1605 (N_1605,N_1007,N_154);
nand U1606 (N_1606,N_641,N_1359);
nor U1607 (N_1607,N_569,N_1385);
nand U1608 (N_1608,N_449,N_609);
nand U1609 (N_1609,N_358,N_646);
xor U1610 (N_1610,N_572,N_1113);
and U1611 (N_1611,N_955,N_168);
and U1612 (N_1612,N_332,N_847);
nand U1613 (N_1613,N_1070,N_171);
nor U1614 (N_1614,N_821,N_1156);
nand U1615 (N_1615,N_1223,N_203);
or U1616 (N_1616,N_1356,N_658);
nor U1617 (N_1617,N_240,N_64);
and U1618 (N_1618,N_615,N_91);
and U1619 (N_1619,N_1489,N_705);
nand U1620 (N_1620,N_61,N_980);
or U1621 (N_1621,N_77,N_650);
and U1622 (N_1622,N_1270,N_298);
or U1623 (N_1623,N_282,N_434);
and U1624 (N_1624,N_190,N_65);
and U1625 (N_1625,N_297,N_795);
and U1626 (N_1626,N_206,N_301);
nor U1627 (N_1627,N_595,N_1117);
or U1628 (N_1628,N_565,N_262);
and U1629 (N_1629,N_1150,N_275);
and U1630 (N_1630,N_824,N_918);
or U1631 (N_1631,N_504,N_521);
and U1632 (N_1632,N_867,N_1471);
nand U1633 (N_1633,N_107,N_680);
and U1634 (N_1634,N_1307,N_461);
nor U1635 (N_1635,N_1155,N_1308);
nand U1636 (N_1636,N_440,N_892);
nand U1637 (N_1637,N_1481,N_291);
nand U1638 (N_1638,N_445,N_51);
and U1639 (N_1639,N_1285,N_334);
and U1640 (N_1640,N_204,N_1003);
or U1641 (N_1641,N_622,N_531);
nor U1642 (N_1642,N_342,N_645);
or U1643 (N_1643,N_468,N_1450);
or U1644 (N_1644,N_1105,N_662);
and U1645 (N_1645,N_555,N_115);
and U1646 (N_1646,N_1443,N_243);
nor U1647 (N_1647,N_1332,N_1300);
nor U1648 (N_1648,N_1304,N_1310);
nor U1649 (N_1649,N_1497,N_4);
and U1650 (N_1650,N_1472,N_1244);
or U1651 (N_1651,N_1108,N_937);
and U1652 (N_1652,N_757,N_348);
nand U1653 (N_1653,N_149,N_740);
nand U1654 (N_1654,N_1188,N_881);
nor U1655 (N_1655,N_260,N_14);
nand U1656 (N_1656,N_634,N_1234);
nor U1657 (N_1657,N_505,N_1404);
and U1658 (N_1658,N_1357,N_269);
nand U1659 (N_1659,N_1152,N_1439);
nor U1660 (N_1660,N_459,N_264);
nor U1661 (N_1661,N_45,N_941);
nor U1662 (N_1662,N_354,N_166);
nand U1663 (N_1663,N_690,N_808);
and U1664 (N_1664,N_1181,N_123);
or U1665 (N_1665,N_250,N_1317);
or U1666 (N_1666,N_991,N_54);
or U1667 (N_1667,N_1224,N_247);
or U1668 (N_1668,N_1153,N_92);
and U1669 (N_1669,N_57,N_381);
or U1670 (N_1670,N_1468,N_920);
or U1671 (N_1671,N_1334,N_1252);
xnor U1672 (N_1672,N_217,N_869);
nor U1673 (N_1673,N_1186,N_932);
nand U1674 (N_1674,N_1086,N_116);
nor U1675 (N_1675,N_671,N_678);
and U1676 (N_1676,N_860,N_1448);
xnor U1677 (N_1677,N_1001,N_385);
nor U1678 (N_1678,N_1363,N_1076);
and U1679 (N_1679,N_241,N_1248);
nor U1680 (N_1680,N_349,N_1302);
or U1681 (N_1681,N_1491,N_183);
nor U1682 (N_1682,N_1342,N_391);
nor U1683 (N_1683,N_143,N_495);
and U1684 (N_1684,N_788,N_1133);
and U1685 (N_1685,N_834,N_1406);
or U1686 (N_1686,N_909,N_24);
nor U1687 (N_1687,N_292,N_995);
nor U1688 (N_1688,N_308,N_653);
nand U1689 (N_1689,N_535,N_903);
or U1690 (N_1690,N_314,N_1060);
or U1691 (N_1691,N_684,N_768);
and U1692 (N_1692,N_525,N_770);
or U1693 (N_1693,N_1219,N_1165);
or U1694 (N_1694,N_435,N_663);
and U1695 (N_1695,N_949,N_296);
or U1696 (N_1696,N_471,N_1095);
or U1697 (N_1697,N_621,N_548);
nor U1698 (N_1698,N_748,N_1080);
nand U1699 (N_1699,N_743,N_1000);
and U1700 (N_1700,N_643,N_484);
nand U1701 (N_1701,N_737,N_1413);
or U1702 (N_1702,N_1477,N_86);
and U1703 (N_1703,N_1132,N_1400);
nor U1704 (N_1704,N_720,N_173);
and U1705 (N_1705,N_244,N_163);
and U1706 (N_1706,N_1447,N_938);
nor U1707 (N_1707,N_877,N_714);
nor U1708 (N_1708,N_774,N_473);
or U1709 (N_1709,N_1116,N_771);
and U1710 (N_1710,N_111,N_971);
and U1711 (N_1711,N_1126,N_829);
and U1712 (N_1712,N_590,N_497);
nor U1713 (N_1713,N_953,N_1034);
nor U1714 (N_1714,N_189,N_359);
nor U1715 (N_1715,N_912,N_202);
or U1716 (N_1716,N_1196,N_562);
nor U1717 (N_1717,N_883,N_223);
and U1718 (N_1718,N_871,N_1137);
nor U1719 (N_1719,N_456,N_225);
nand U1720 (N_1720,N_1484,N_933);
and U1721 (N_1721,N_674,N_429);
and U1722 (N_1722,N_12,N_558);
nor U1723 (N_1723,N_1286,N_1220);
and U1724 (N_1724,N_1102,N_986);
nor U1725 (N_1725,N_415,N_74);
and U1726 (N_1726,N_213,N_1067);
and U1727 (N_1727,N_1232,N_318);
and U1728 (N_1728,N_1435,N_227);
or U1729 (N_1729,N_186,N_401);
nor U1730 (N_1730,N_1369,N_324);
nand U1731 (N_1731,N_801,N_1268);
and U1732 (N_1732,N_512,N_396);
and U1733 (N_1733,N_447,N_1492);
nor U1734 (N_1734,N_1044,N_69);
or U1735 (N_1735,N_1337,N_410);
nor U1736 (N_1736,N_1386,N_1159);
nand U1737 (N_1737,N_158,N_1225);
nand U1738 (N_1738,N_810,N_405);
nor U1739 (N_1739,N_1111,N_630);
or U1740 (N_1740,N_849,N_546);
or U1741 (N_1741,N_323,N_1348);
nor U1742 (N_1742,N_889,N_207);
and U1743 (N_1743,N_1373,N_668);
nand U1744 (N_1744,N_228,N_667);
or U1745 (N_1745,N_785,N_1329);
and U1746 (N_1746,N_534,N_664);
and U1747 (N_1747,N_1454,N_686);
nor U1748 (N_1748,N_1020,N_846);
nand U1749 (N_1749,N_843,N_501);
and U1750 (N_1750,N_806,N_44);
nand U1751 (N_1751,N_999,N_1176);
or U1752 (N_1752,N_1029,N_983);
or U1753 (N_1753,N_1146,N_1394);
nand U1754 (N_1754,N_563,N_188);
and U1755 (N_1755,N_352,N_472);
and U1756 (N_1756,N_1030,N_1431);
and U1757 (N_1757,N_778,N_811);
or U1758 (N_1758,N_627,N_853);
and U1759 (N_1759,N_1241,N_60);
or U1760 (N_1760,N_851,N_729);
or U1761 (N_1761,N_70,N_648);
and U1762 (N_1762,N_551,N_164);
and U1763 (N_1763,N_1124,N_245);
nor U1764 (N_1764,N_1183,N_27);
or U1765 (N_1765,N_979,N_408);
or U1766 (N_1766,N_1079,N_837);
or U1767 (N_1767,N_356,N_1005);
or U1768 (N_1768,N_172,N_989);
nor U1769 (N_1769,N_187,N_744);
or U1770 (N_1770,N_557,N_375);
or U1771 (N_1771,N_721,N_175);
xnor U1772 (N_1772,N_707,N_1284);
and U1773 (N_1773,N_84,N_592);
or U1774 (N_1774,N_379,N_679);
or U1775 (N_1775,N_520,N_611);
and U1776 (N_1776,N_532,N_1192);
or U1777 (N_1777,N_1136,N_1040);
or U1778 (N_1778,N_450,N_467);
nand U1779 (N_1779,N_593,N_289);
and U1780 (N_1780,N_922,N_329);
and U1781 (N_1781,N_1148,N_950);
and U1782 (N_1782,N_1138,N_1098);
and U1783 (N_1783,N_844,N_1344);
nand U1784 (N_1784,N_568,N_1422);
nor U1785 (N_1785,N_481,N_765);
or U1786 (N_1786,N_22,N_1238);
nor U1787 (N_1787,N_114,N_865);
and U1788 (N_1788,N_1264,N_746);
nand U1789 (N_1789,N_85,N_1139);
or U1790 (N_1790,N_1206,N_1217);
or U1791 (N_1791,N_1254,N_564);
nand U1792 (N_1792,N_41,N_1267);
or U1793 (N_1793,N_975,N_199);
nor U1794 (N_1794,N_1041,N_1197);
and U1795 (N_1795,N_508,N_1349);
and U1796 (N_1796,N_487,N_596);
nand U1797 (N_1797,N_1303,N_336);
and U1798 (N_1798,N_2,N_312);
or U1799 (N_1799,N_694,N_677);
nand U1800 (N_1800,N_1210,N_835);
xor U1801 (N_1801,N_251,N_617);
nand U1802 (N_1802,N_845,N_407);
nand U1803 (N_1803,N_1328,N_577);
and U1804 (N_1804,N_1350,N_1418);
nand U1805 (N_1805,N_1388,N_1173);
nor U1806 (N_1806,N_864,N_1036);
nor U1807 (N_1807,N_685,N_576);
nand U1808 (N_1808,N_193,N_836);
nor U1809 (N_1809,N_1376,N_331);
or U1810 (N_1810,N_129,N_1424);
nand U1811 (N_1811,N_1236,N_210);
nor U1812 (N_1812,N_165,N_340);
nand U1813 (N_1813,N_1486,N_78);
or U1814 (N_1814,N_573,N_1311);
nor U1815 (N_1815,N_1051,N_1008);
nand U1816 (N_1816,N_947,N_360);
and U1817 (N_1817,N_613,N_614);
nor U1818 (N_1818,N_201,N_194);
and U1819 (N_1819,N_1179,N_1354);
nor U1820 (N_1820,N_1365,N_1446);
nand U1821 (N_1821,N_700,N_709);
nor U1822 (N_1822,N_783,N_552);
or U1823 (N_1823,N_826,N_523);
nand U1824 (N_1824,N_1115,N_1172);
nand U1825 (N_1825,N_1475,N_868);
nand U1826 (N_1826,N_1237,N_1247);
or U1827 (N_1827,N_287,N_990);
nor U1828 (N_1828,N_676,N_1294);
nand U1829 (N_1829,N_959,N_761);
or U1830 (N_1830,N_1467,N_1033);
nor U1831 (N_1831,N_161,N_325);
nand U1832 (N_1832,N_1425,N_647);
or U1833 (N_1833,N_58,N_581);
or U1834 (N_1834,N_1011,N_1260);
nand U1835 (N_1835,N_109,N_878);
nand U1836 (N_1836,N_863,N_599);
nor U1837 (N_1837,N_1440,N_575);
or U1838 (N_1838,N_1058,N_451);
or U1839 (N_1839,N_722,N_730);
or U1840 (N_1840,N_1200,N_610);
and U1841 (N_1841,N_330,N_304);
nand U1842 (N_1842,N_582,N_1211);
or U1843 (N_1843,N_681,N_376);
nor U1844 (N_1844,N_772,N_1062);
nor U1845 (N_1845,N_63,N_169);
nand U1846 (N_1846,N_642,N_1026);
or U1847 (N_1847,N_733,N_432);
nor U1848 (N_1848,N_140,N_591);
nor U1849 (N_1849,N_283,N_537);
or U1850 (N_1850,N_333,N_279);
or U1851 (N_1851,N_894,N_366);
nor U1852 (N_1852,N_736,N_956);
nor U1853 (N_1853,N_67,N_1130);
and U1854 (N_1854,N_421,N_963);
nand U1855 (N_1855,N_1199,N_891);
nor U1856 (N_1856,N_776,N_350);
or U1857 (N_1857,N_89,N_1180);
nand U1858 (N_1858,N_659,N_607);
nor U1859 (N_1859,N_660,N_655);
nor U1860 (N_1860,N_1056,N_209);
nor U1861 (N_1861,N_1031,N_823);
or U1862 (N_1862,N_510,N_34);
or U1863 (N_1863,N_226,N_905);
nor U1864 (N_1864,N_285,N_306);
nand U1865 (N_1865,N_885,N_1242);
nand U1866 (N_1866,N_661,N_1129);
nor U1867 (N_1867,N_786,N_605);
or U1868 (N_1868,N_120,N_101);
and U1869 (N_1869,N_954,N_338);
nor U1870 (N_1870,N_598,N_1075);
nor U1871 (N_1871,N_904,N_719);
nand U1872 (N_1872,N_513,N_1262);
or U1873 (N_1873,N_793,N_277);
nand U1874 (N_1874,N_751,N_403);
xor U1875 (N_1875,N_1087,N_131);
xor U1876 (N_1876,N_1330,N_420);
nand U1877 (N_1877,N_529,N_446);
or U1878 (N_1878,N_457,N_689);
and U1879 (N_1879,N_422,N_82);
and U1880 (N_1880,N_1215,N_90);
or U1881 (N_1881,N_926,N_998);
and U1882 (N_1882,N_619,N_528);
or U1883 (N_1883,N_159,N_443);
nand U1884 (N_1884,N_5,N_214);
nor U1885 (N_1885,N_498,N_763);
nand U1886 (N_1886,N_1261,N_254);
and U1887 (N_1887,N_462,N_479);
nand U1888 (N_1888,N_606,N_253);
nor U1889 (N_1889,N_1390,N_1178);
and U1890 (N_1890,N_1368,N_934);
nand U1891 (N_1891,N_1380,N_1283);
and U1892 (N_1892,N_583,N_1258);
nor U1893 (N_1893,N_1313,N_1175);
and U1894 (N_1894,N_618,N_1169);
nor U1895 (N_1895,N_784,N_1118);
or U1896 (N_1896,N_625,N_1208);
nand U1897 (N_1897,N_231,N_939);
nor U1898 (N_1898,N_1071,N_48);
xor U1899 (N_1899,N_40,N_862);
and U1900 (N_1900,N_580,N_797);
or U1901 (N_1901,N_682,N_976);
or U1902 (N_1902,N_977,N_1403);
or U1903 (N_1903,N_388,N_803);
nor U1904 (N_1904,N_1054,N_13);
xor U1905 (N_1905,N_273,N_1053);
and U1906 (N_1906,N_9,N_514);
or U1907 (N_1907,N_364,N_1218);
or U1908 (N_1908,N_465,N_1338);
or U1909 (N_1909,N_1273,N_1383);
nand U1910 (N_1910,N_288,N_126);
nor U1911 (N_1911,N_488,N_967);
nor U1912 (N_1912,N_632,N_1035);
nand U1913 (N_1913,N_427,N_300);
or U1914 (N_1914,N_23,N_156);
nand U1915 (N_1915,N_1487,N_252);
or U1916 (N_1916,N_179,N_47);
or U1917 (N_1917,N_1419,N_530);
and U1918 (N_1918,N_1433,N_477);
nor U1919 (N_1919,N_389,N_1101);
or U1920 (N_1920,N_1407,N_917);
or U1921 (N_1921,N_1193,N_1163);
nand U1922 (N_1922,N_439,N_1201);
nor U1923 (N_1923,N_974,N_755);
nor U1924 (N_1924,N_141,N_1203);
and U1925 (N_1925,N_899,N_696);
nand U1926 (N_1926,N_353,N_229);
and U1927 (N_1927,N_1239,N_1287);
nor U1928 (N_1928,N_800,N_620);
and U1929 (N_1929,N_928,N_1272);
nor U1930 (N_1930,N_1023,N_815);
nand U1931 (N_1931,N_970,N_742);
or U1932 (N_1932,N_42,N_1235);
and U1933 (N_1933,N_527,N_460);
or U1934 (N_1934,N_587,N_75);
or U1935 (N_1935,N_672,N_399);
and U1936 (N_1936,N_1145,N_698);
nand U1937 (N_1937,N_644,N_6);
nand U1938 (N_1938,N_1490,N_708);
and U1939 (N_1939,N_1083,N_1104);
or U1940 (N_1940,N_1351,N_1107);
nand U1941 (N_1941,N_1466,N_470);
xnor U1942 (N_1942,N_147,N_931);
and U1943 (N_1943,N_1065,N_1476);
and U1944 (N_1944,N_1174,N_1397);
xor U1945 (N_1945,N_923,N_706);
or U1946 (N_1946,N_322,N_1290);
nor U1947 (N_1947,N_167,N_968);
nand U1948 (N_1948,N_913,N_1047);
and U1949 (N_1949,N_1,N_278);
xnor U1950 (N_1950,N_713,N_855);
nor U1951 (N_1951,N_72,N_946);
and U1952 (N_1952,N_781,N_790);
and U1953 (N_1953,N_219,N_675);
or U1954 (N_1954,N_1227,N_68);
and U1955 (N_1955,N_1316,N_317);
and U1956 (N_1956,N_326,N_153);
or U1957 (N_1957,N_545,N_910);
and U1958 (N_1958,N_884,N_1233);
nand U1959 (N_1959,N_365,N_1358);
nor U1960 (N_1960,N_1456,N_602);
and U1961 (N_1961,N_486,N_1372);
or U1962 (N_1962,N_444,N_566);
nand U1963 (N_1963,N_616,N_726);
nor U1964 (N_1964,N_1314,N_8);
or U1965 (N_1965,N_1251,N_1438);
nand U1966 (N_1966,N_1444,N_38);
nor U1967 (N_1967,N_455,N_411);
nand U1968 (N_1968,N_856,N_822);
nor U1969 (N_1969,N_571,N_1166);
nand U1970 (N_1970,N_1209,N_952);
nand U1971 (N_1971,N_1016,N_1228);
and U1972 (N_1972,N_265,N_544);
nand U1973 (N_1973,N_320,N_978);
nor U1974 (N_1974,N_1263,N_897);
or U1975 (N_1975,N_816,N_170);
or U1976 (N_1976,N_414,N_775);
nor U1977 (N_1977,N_1122,N_321);
or U1978 (N_1978,N_249,N_930);
or U1979 (N_1979,N_148,N_400);
nand U1980 (N_1980,N_1158,N_888);
nor U1981 (N_1981,N_902,N_919);
nor U1982 (N_1982,N_712,N_560);
and U1983 (N_1983,N_1402,N_425);
nand U1984 (N_1984,N_710,N_242);
or U1985 (N_1985,N_119,N_818);
or U1986 (N_1986,N_1205,N_255);
or U1987 (N_1987,N_1157,N_1391);
or U1988 (N_1988,N_517,N_1085);
nor U1989 (N_1989,N_1408,N_895);
and U1990 (N_1990,N_945,N_907);
and U1991 (N_1991,N_809,N_839);
nand U1992 (N_1992,N_286,N_151);
nand U1993 (N_1993,N_882,N_1333);
and U1994 (N_1994,N_1384,N_1171);
or U1995 (N_1995,N_1198,N_600);
or U1996 (N_1996,N_490,N_224);
xor U1997 (N_1997,N_196,N_1322);
or U1998 (N_1998,N_441,N_921);
xnor U1999 (N_1999,N_1125,N_550);
nor U2000 (N_2000,N_1052,N_840);
nand U2001 (N_2001,N_1022,N_235);
nor U2002 (N_2002,N_1063,N_1082);
nand U2003 (N_2003,N_1414,N_875);
and U2004 (N_2004,N_397,N_0);
nor U2005 (N_2005,N_1037,N_452);
xor U2006 (N_2006,N_346,N_311);
nand U2007 (N_2007,N_1213,N_105);
nor U2008 (N_2008,N_1392,N_1301);
and U2009 (N_2009,N_1412,N_426);
and U2010 (N_2010,N_380,N_344);
nor U2011 (N_2011,N_541,N_1154);
or U2012 (N_2012,N_1463,N_418);
nor U2013 (N_2013,N_236,N_1092);
or U2014 (N_2014,N_328,N_270);
nor U2015 (N_2015,N_11,N_908);
nor U2016 (N_2016,N_966,N_416);
or U2017 (N_2017,N_36,N_624);
and U2018 (N_2018,N_1143,N_295);
nand U2019 (N_2019,N_208,N_25);
nor U2020 (N_2020,N_1449,N_30);
and U2021 (N_2021,N_942,N_762);
nor U2022 (N_2022,N_792,N_1336);
nor U2023 (N_2023,N_789,N_1025);
nand U2024 (N_2024,N_1485,N_997);
nand U2025 (N_2025,N_1410,N_1194);
nand U2026 (N_2026,N_1379,N_1012);
nor U2027 (N_2027,N_688,N_1049);
or U2028 (N_2028,N_1013,N_1480);
nand U2029 (N_2029,N_1255,N_281);
and U2030 (N_2030,N_940,N_108);
and U2031 (N_2031,N_683,N_1320);
nand U2032 (N_2032,N_1068,N_1370);
and U2033 (N_2033,N_993,N_1341);
or U2034 (N_2034,N_842,N_935);
and U2035 (N_2035,N_1002,N_972);
nor U2036 (N_2036,N_395,N_858);
or U2037 (N_2037,N_299,N_695);
xor U2038 (N_2038,N_394,N_339);
nand U2039 (N_2039,N_239,N_944);
and U2040 (N_2040,N_1343,N_1050);
nand U2041 (N_2041,N_794,N_533);
or U2042 (N_2042,N_43,N_1382);
or U2043 (N_2043,N_876,N_271);
and U2044 (N_2044,N_327,N_1112);
or U2045 (N_2045,N_37,N_1432);
and U2046 (N_2046,N_914,N_10);
nor U2047 (N_2047,N_1277,N_152);
and U2048 (N_2048,N_820,N_1240);
and U2049 (N_2049,N_1162,N_854);
or U2050 (N_2050,N_31,N_594);
nor U2051 (N_2051,N_1375,N_1478);
or U2052 (N_2052,N_637,N_1281);
or U2053 (N_2053,N_1366,N_1114);
nor U2054 (N_2054,N_1371,N_99);
or U2055 (N_2055,N_561,N_1436);
nor U2056 (N_2056,N_32,N_608);
and U2057 (N_2057,N_478,N_200);
and U2058 (N_2058,N_636,N_1099);
and U2059 (N_2059,N_433,N_916);
and U2060 (N_2060,N_1204,N_494);
or U2061 (N_2061,N_466,N_699);
and U2062 (N_2062,N_374,N_195);
or U2063 (N_2063,N_651,N_969);
nand U2064 (N_2064,N_753,N_749);
nor U2065 (N_2065,N_1185,N_900);
nor U2066 (N_2066,N_500,N_1275);
and U2067 (N_2067,N_502,N_691);
nor U2068 (N_2068,N_1072,N_693);
nor U2069 (N_2069,N_1190,N_50);
nor U2070 (N_2070,N_1027,N_1321);
and U2071 (N_2071,N_117,N_727);
nor U2072 (N_2072,N_1465,N_759);
nand U2073 (N_2073,N_503,N_911);
nor U2074 (N_2074,N_559,N_1409);
nand U2075 (N_2075,N_812,N_924);
nand U2076 (N_2076,N_234,N_987);
and U2077 (N_2077,N_402,N_475);
and U2078 (N_2078,N_543,N_1142);
nand U2079 (N_2079,N_1494,N_1055);
nor U2080 (N_2080,N_1355,N_984);
and U2081 (N_2081,N_1202,N_1398);
or U2082 (N_2082,N_734,N_893);
and U2083 (N_2083,N_1048,N_807);
and U2084 (N_2084,N_524,N_150);
nor U2085 (N_2085,N_79,N_1109);
or U2086 (N_2086,N_182,N_127);
or U2087 (N_2087,N_631,N_994);
or U2088 (N_2088,N_1289,N_1495);
nor U2089 (N_2089,N_890,N_39);
nand U2090 (N_2090,N_191,N_145);
nor U2091 (N_2091,N_1074,N_1004);
or U2092 (N_2092,N_948,N_1282);
nand U2093 (N_2093,N_670,N_1451);
nand U2094 (N_2094,N_1299,N_1018);
nand U2095 (N_2095,N_1266,N_1043);
nor U2096 (N_2096,N_506,N_382);
and U2097 (N_2097,N_828,N_973);
and U2098 (N_2098,N_1291,N_1090);
nor U2099 (N_2099,N_1323,N_1306);
or U2100 (N_2100,N_1140,N_428);
nand U2101 (N_2101,N_626,N_1046);
and U2102 (N_2102,N_372,N_556);
nand U2103 (N_2103,N_28,N_347);
and U2104 (N_2104,N_1377,N_136);
nand U2105 (N_2105,N_1445,N_1257);
or U2106 (N_2106,N_964,N_1216);
nor U2107 (N_2107,N_725,N_1298);
or U2108 (N_2108,N_747,N_303);
or U2109 (N_2109,N_638,N_799);
nand U2110 (N_2110,N_1318,N_174);
nor U2111 (N_2111,N_704,N_1151);
nand U2112 (N_2112,N_489,N_1045);
nand U2113 (N_2113,N_1315,N_1453);
nor U2114 (N_2114,N_758,N_491);
or U2115 (N_2115,N_519,N_782);
nand U2116 (N_2116,N_66,N_738);
nor U2117 (N_2117,N_669,N_1474);
and U2118 (N_2118,N_1149,N_1458);
and U2119 (N_2119,N_1089,N_1346);
or U2120 (N_2120,N_1452,N_814);
nand U2121 (N_2121,N_1064,N_1259);
or U2122 (N_2122,N_386,N_1127);
nand U2123 (N_2123,N_49,N_539);
nand U2124 (N_2124,N_1374,N_106);
nor U2125 (N_2125,N_589,N_371);
nor U2126 (N_2126,N_511,N_1331);
nor U2127 (N_2127,N_526,N_833);
nand U2128 (N_2128,N_1278,N_97);
xor U2129 (N_2129,N_137,N_1161);
nor U2130 (N_2130,N_237,N_791);
or U2131 (N_2131,N_830,N_248);
or U2132 (N_2132,N_961,N_601);
nand U2133 (N_2133,N_355,N_1069);
and U2134 (N_2134,N_1401,N_1077);
or U2135 (N_2135,N_1361,N_728);
or U2136 (N_2136,N_313,N_804);
nand U2137 (N_2137,N_197,N_1493);
nor U2138 (N_2138,N_1496,N_1243);
nand U2139 (N_2139,N_767,N_406);
and U2140 (N_2140,N_1073,N_859);
nand U2141 (N_2141,N_817,N_351);
nand U2142 (N_2142,N_981,N_553);
and U2143 (N_2143,N_17,N_925);
and U2144 (N_2144,N_982,N_221);
nor U2145 (N_2145,N_390,N_1269);
nand U2146 (N_2146,N_1340,N_901);
nand U2147 (N_2147,N_1093,N_46);
and U2148 (N_2148,N_635,N_1411);
nor U2149 (N_2149,N_162,N_887);
and U2150 (N_2150,N_419,N_1230);
nor U2151 (N_2151,N_1430,N_492);
or U2152 (N_2152,N_874,N_780);
and U2153 (N_2153,N_716,N_80);
or U2154 (N_2154,N_1367,N_211);
nand U2155 (N_2155,N_927,N_1309);
or U2156 (N_2156,N_216,N_603);
nand U2157 (N_2157,N_423,N_579);
or U2158 (N_2158,N_157,N_701);
or U2159 (N_2159,N_988,N_1364);
or U2160 (N_2160,N_852,N_1360);
or U2161 (N_2161,N_873,N_404);
and U2162 (N_2162,N_584,N_424);
or U2163 (N_2163,N_1024,N_307);
nand U2164 (N_2164,N_215,N_1347);
nand U2165 (N_2165,N_417,N_272);
and U2166 (N_2166,N_1345,N_1423);
and U2167 (N_2167,N_1106,N_1231);
and U2168 (N_2168,N_832,N_246);
nand U2169 (N_2169,N_1184,N_357);
nand U2170 (N_2170,N_485,N_1088);
nor U2171 (N_2171,N_1229,N_1246);
nor U2172 (N_2172,N_142,N_1274);
and U2173 (N_2173,N_230,N_1191);
and U2174 (N_2174,N_1207,N_796);
nand U2175 (N_2175,N_1160,N_629);
and U2176 (N_2176,N_538,N_88);
and U2177 (N_2177,N_62,N_409);
or U2178 (N_2178,N_83,N_392);
or U2179 (N_2179,N_1009,N_493);
nor U2180 (N_2180,N_363,N_55);
or U2181 (N_2181,N_1081,N_604);
or U2182 (N_2182,N_102,N_1170);
or U2183 (N_2183,N_1167,N_711);
nand U2184 (N_2184,N_1212,N_1097);
nor U2185 (N_2185,N_1189,N_383);
or U2186 (N_2186,N_21,N_1265);
nand U2187 (N_2187,N_724,N_184);
or U2188 (N_2188,N_1416,N_95);
nor U2189 (N_2189,N_1066,N_687);
nand U2190 (N_2190,N_361,N_20);
nand U2191 (N_2191,N_717,N_337);
or U2192 (N_2192,N_813,N_1288);
nand U2193 (N_2193,N_1039,N_73);
and U2194 (N_2194,N_652,N_805);
nor U2195 (N_2195,N_1399,N_192);
and U2196 (N_2196,N_110,N_1437);
nand U2197 (N_2197,N_951,N_1319);
xor U2198 (N_2198,N_649,N_121);
nor U2199 (N_2199,N_319,N_1222);
or U2200 (N_2200,N_1296,N_430);
nand U2201 (N_2201,N_1195,N_985);
and U2202 (N_2202,N_413,N_1100);
nand U2203 (N_2203,N_1276,N_463);
xor U2204 (N_2204,N_100,N_290);
nor U2205 (N_2205,N_280,N_1078);
nand U2206 (N_2206,N_1488,N_18);
or U2207 (N_2207,N_943,N_480);
nand U2208 (N_2208,N_578,N_310);
nand U2209 (N_2209,N_1249,N_1427);
or U2210 (N_2210,N_1253,N_238);
nand U2211 (N_2211,N_536,N_554);
nand U2212 (N_2212,N_1389,N_146);
nor U2213 (N_2213,N_1429,N_739);
and U2214 (N_2214,N_177,N_112);
or U2215 (N_2215,N_992,N_1135);
nor U2216 (N_2216,N_454,N_377);
nor U2217 (N_2217,N_474,N_144);
or U2218 (N_2218,N_458,N_1096);
or U2219 (N_2219,N_284,N_26);
or U2220 (N_2220,N_665,N_866);
nor U2221 (N_2221,N_507,N_267);
and U2222 (N_2222,N_335,N_222);
and U2223 (N_2223,N_1378,N_766);
nor U2224 (N_2224,N_132,N_1335);
and U2225 (N_2225,N_929,N_741);
xnor U2226 (N_2226,N_639,N_880);
and U2227 (N_2227,N_1091,N_367);
nand U2228 (N_2228,N_133,N_1479);
or U2229 (N_2229,N_958,N_731);
or U2230 (N_2230,N_640,N_29);
nand U2231 (N_2231,N_1352,N_996);
or U2232 (N_2232,N_345,N_715);
or U2233 (N_2233,N_732,N_1362);
nor U2234 (N_2234,N_309,N_1147);
nor U2235 (N_2235,N_453,N_464);
or U2236 (N_2236,N_628,N_879);
nor U2237 (N_2237,N_570,N_113);
nor U2238 (N_2238,N_384,N_1280);
nor U2239 (N_2239,N_212,N_896);
and U2240 (N_2240,N_1327,N_155);
or U2241 (N_2241,N_1395,N_1038);
nor U2242 (N_2242,N_542,N_1177);
and U2243 (N_2243,N_612,N_697);
xnor U2244 (N_2244,N_3,N_723);
or U2245 (N_2245,N_1123,N_745);
and U2246 (N_2246,N_1293,N_1141);
or U2247 (N_2247,N_1134,N_19);
nand U2248 (N_2248,N_442,N_1459);
and U2249 (N_2249,N_52,N_540);
or U2250 (N_2250,N_1304,N_425);
and U2251 (N_2251,N_1153,N_176);
or U2252 (N_2252,N_1131,N_1431);
or U2253 (N_2253,N_92,N_266);
nor U2254 (N_2254,N_1323,N_1180);
and U2255 (N_2255,N_434,N_1470);
nor U2256 (N_2256,N_967,N_171);
nor U2257 (N_2257,N_308,N_408);
xnor U2258 (N_2258,N_631,N_1304);
nand U2259 (N_2259,N_493,N_228);
or U2260 (N_2260,N_469,N_880);
nor U2261 (N_2261,N_245,N_445);
nand U2262 (N_2262,N_805,N_90);
or U2263 (N_2263,N_1329,N_353);
nand U2264 (N_2264,N_1272,N_179);
or U2265 (N_2265,N_181,N_214);
or U2266 (N_2266,N_734,N_944);
or U2267 (N_2267,N_1412,N_1399);
nand U2268 (N_2268,N_756,N_264);
or U2269 (N_2269,N_1425,N_1154);
and U2270 (N_2270,N_4,N_225);
nor U2271 (N_2271,N_207,N_1402);
and U2272 (N_2272,N_994,N_1001);
or U2273 (N_2273,N_42,N_40);
nor U2274 (N_2274,N_5,N_1119);
and U2275 (N_2275,N_362,N_793);
and U2276 (N_2276,N_345,N_1152);
and U2277 (N_2277,N_455,N_1148);
xnor U2278 (N_2278,N_171,N_300);
nand U2279 (N_2279,N_537,N_844);
nor U2280 (N_2280,N_470,N_1463);
and U2281 (N_2281,N_665,N_672);
or U2282 (N_2282,N_977,N_1188);
nand U2283 (N_2283,N_1029,N_569);
nor U2284 (N_2284,N_571,N_1360);
nand U2285 (N_2285,N_1234,N_1446);
xnor U2286 (N_2286,N_635,N_1341);
or U2287 (N_2287,N_1366,N_1190);
nor U2288 (N_2288,N_602,N_872);
nand U2289 (N_2289,N_1427,N_1260);
and U2290 (N_2290,N_959,N_1318);
nor U2291 (N_2291,N_176,N_1066);
and U2292 (N_2292,N_270,N_926);
or U2293 (N_2293,N_1486,N_1198);
and U2294 (N_2294,N_414,N_526);
nand U2295 (N_2295,N_131,N_827);
and U2296 (N_2296,N_1435,N_1414);
or U2297 (N_2297,N_1206,N_643);
nor U2298 (N_2298,N_770,N_365);
nor U2299 (N_2299,N_536,N_614);
nand U2300 (N_2300,N_1433,N_1122);
xor U2301 (N_2301,N_504,N_677);
or U2302 (N_2302,N_10,N_1197);
or U2303 (N_2303,N_909,N_663);
nor U2304 (N_2304,N_667,N_208);
and U2305 (N_2305,N_583,N_739);
or U2306 (N_2306,N_562,N_668);
nor U2307 (N_2307,N_174,N_114);
and U2308 (N_2308,N_1185,N_180);
nand U2309 (N_2309,N_807,N_847);
nor U2310 (N_2310,N_952,N_1488);
and U2311 (N_2311,N_1359,N_1427);
nor U2312 (N_2312,N_1151,N_178);
nor U2313 (N_2313,N_1105,N_352);
and U2314 (N_2314,N_306,N_163);
xor U2315 (N_2315,N_797,N_356);
and U2316 (N_2316,N_265,N_47);
and U2317 (N_2317,N_478,N_30);
or U2318 (N_2318,N_991,N_1230);
nor U2319 (N_2319,N_929,N_904);
and U2320 (N_2320,N_875,N_1003);
or U2321 (N_2321,N_296,N_72);
xor U2322 (N_2322,N_1473,N_113);
nor U2323 (N_2323,N_1476,N_1013);
nor U2324 (N_2324,N_1165,N_566);
nand U2325 (N_2325,N_17,N_865);
and U2326 (N_2326,N_65,N_1407);
nand U2327 (N_2327,N_1350,N_366);
or U2328 (N_2328,N_973,N_1413);
nand U2329 (N_2329,N_679,N_1469);
nor U2330 (N_2330,N_708,N_988);
and U2331 (N_2331,N_1380,N_1439);
and U2332 (N_2332,N_443,N_847);
or U2333 (N_2333,N_321,N_210);
nand U2334 (N_2334,N_940,N_833);
nor U2335 (N_2335,N_673,N_1424);
nand U2336 (N_2336,N_885,N_1351);
nand U2337 (N_2337,N_752,N_1270);
xor U2338 (N_2338,N_108,N_272);
or U2339 (N_2339,N_311,N_1446);
nor U2340 (N_2340,N_433,N_287);
and U2341 (N_2341,N_395,N_1372);
nand U2342 (N_2342,N_1375,N_723);
and U2343 (N_2343,N_768,N_536);
nand U2344 (N_2344,N_333,N_468);
nand U2345 (N_2345,N_206,N_568);
nor U2346 (N_2346,N_1063,N_590);
or U2347 (N_2347,N_364,N_640);
nor U2348 (N_2348,N_1034,N_865);
nand U2349 (N_2349,N_1136,N_1107);
nor U2350 (N_2350,N_559,N_1337);
nor U2351 (N_2351,N_404,N_813);
xor U2352 (N_2352,N_883,N_921);
nor U2353 (N_2353,N_12,N_348);
nor U2354 (N_2354,N_905,N_590);
nand U2355 (N_2355,N_625,N_1119);
or U2356 (N_2356,N_344,N_928);
and U2357 (N_2357,N_1328,N_252);
nor U2358 (N_2358,N_452,N_899);
nor U2359 (N_2359,N_65,N_1198);
nor U2360 (N_2360,N_223,N_921);
nor U2361 (N_2361,N_1114,N_637);
and U2362 (N_2362,N_1442,N_211);
nand U2363 (N_2363,N_937,N_2);
and U2364 (N_2364,N_644,N_182);
nand U2365 (N_2365,N_161,N_1114);
nand U2366 (N_2366,N_949,N_111);
nand U2367 (N_2367,N_114,N_699);
or U2368 (N_2368,N_560,N_649);
nand U2369 (N_2369,N_1447,N_1117);
nor U2370 (N_2370,N_411,N_485);
nand U2371 (N_2371,N_1373,N_1007);
and U2372 (N_2372,N_889,N_559);
nor U2373 (N_2373,N_736,N_1386);
xor U2374 (N_2374,N_101,N_1488);
and U2375 (N_2375,N_508,N_1381);
or U2376 (N_2376,N_772,N_474);
nand U2377 (N_2377,N_1307,N_1429);
nand U2378 (N_2378,N_466,N_197);
or U2379 (N_2379,N_179,N_1453);
and U2380 (N_2380,N_1123,N_1079);
or U2381 (N_2381,N_316,N_211);
nand U2382 (N_2382,N_1327,N_535);
or U2383 (N_2383,N_107,N_255);
nor U2384 (N_2384,N_1087,N_1411);
nor U2385 (N_2385,N_733,N_361);
nor U2386 (N_2386,N_1294,N_306);
nand U2387 (N_2387,N_672,N_304);
or U2388 (N_2388,N_1116,N_1205);
or U2389 (N_2389,N_806,N_459);
nand U2390 (N_2390,N_1489,N_283);
nand U2391 (N_2391,N_444,N_1277);
nand U2392 (N_2392,N_690,N_476);
nand U2393 (N_2393,N_373,N_494);
nor U2394 (N_2394,N_826,N_688);
nand U2395 (N_2395,N_1437,N_945);
or U2396 (N_2396,N_1437,N_232);
nor U2397 (N_2397,N_1140,N_328);
or U2398 (N_2398,N_887,N_1079);
nor U2399 (N_2399,N_597,N_1052);
nand U2400 (N_2400,N_44,N_1267);
nor U2401 (N_2401,N_23,N_1202);
nor U2402 (N_2402,N_1234,N_1179);
nor U2403 (N_2403,N_223,N_495);
or U2404 (N_2404,N_642,N_1304);
and U2405 (N_2405,N_1148,N_577);
nor U2406 (N_2406,N_218,N_1058);
and U2407 (N_2407,N_362,N_668);
or U2408 (N_2408,N_1484,N_101);
nand U2409 (N_2409,N_935,N_1082);
or U2410 (N_2410,N_942,N_353);
and U2411 (N_2411,N_1448,N_438);
or U2412 (N_2412,N_1288,N_1265);
nor U2413 (N_2413,N_1375,N_979);
or U2414 (N_2414,N_1013,N_789);
xor U2415 (N_2415,N_905,N_571);
and U2416 (N_2416,N_724,N_356);
nand U2417 (N_2417,N_1189,N_513);
nor U2418 (N_2418,N_683,N_388);
or U2419 (N_2419,N_968,N_438);
or U2420 (N_2420,N_351,N_722);
nor U2421 (N_2421,N_1134,N_1333);
nand U2422 (N_2422,N_208,N_41);
or U2423 (N_2423,N_903,N_769);
nand U2424 (N_2424,N_1387,N_953);
and U2425 (N_2425,N_249,N_1059);
and U2426 (N_2426,N_137,N_1187);
nand U2427 (N_2427,N_1428,N_558);
or U2428 (N_2428,N_1494,N_1109);
or U2429 (N_2429,N_554,N_588);
or U2430 (N_2430,N_836,N_1127);
nor U2431 (N_2431,N_1362,N_682);
xor U2432 (N_2432,N_719,N_0);
or U2433 (N_2433,N_838,N_151);
or U2434 (N_2434,N_343,N_795);
xor U2435 (N_2435,N_631,N_260);
nor U2436 (N_2436,N_743,N_1152);
nand U2437 (N_2437,N_1355,N_89);
or U2438 (N_2438,N_674,N_1450);
and U2439 (N_2439,N_394,N_931);
and U2440 (N_2440,N_242,N_1354);
and U2441 (N_2441,N_300,N_1490);
or U2442 (N_2442,N_132,N_476);
or U2443 (N_2443,N_1482,N_473);
nor U2444 (N_2444,N_1421,N_1458);
nand U2445 (N_2445,N_1489,N_279);
xnor U2446 (N_2446,N_27,N_1299);
nand U2447 (N_2447,N_1167,N_161);
and U2448 (N_2448,N_1055,N_977);
or U2449 (N_2449,N_982,N_505);
nand U2450 (N_2450,N_892,N_666);
nand U2451 (N_2451,N_1081,N_1467);
nand U2452 (N_2452,N_1191,N_223);
nor U2453 (N_2453,N_166,N_425);
and U2454 (N_2454,N_751,N_1225);
xnor U2455 (N_2455,N_1434,N_1440);
nand U2456 (N_2456,N_1196,N_552);
or U2457 (N_2457,N_1419,N_602);
nand U2458 (N_2458,N_716,N_335);
and U2459 (N_2459,N_1295,N_1021);
nand U2460 (N_2460,N_1084,N_1448);
nand U2461 (N_2461,N_343,N_1031);
or U2462 (N_2462,N_683,N_1449);
or U2463 (N_2463,N_947,N_543);
nand U2464 (N_2464,N_480,N_1279);
nor U2465 (N_2465,N_49,N_1022);
and U2466 (N_2466,N_1191,N_1242);
nor U2467 (N_2467,N_846,N_532);
and U2468 (N_2468,N_603,N_241);
nand U2469 (N_2469,N_852,N_681);
and U2470 (N_2470,N_1140,N_1425);
nand U2471 (N_2471,N_728,N_177);
and U2472 (N_2472,N_133,N_185);
and U2473 (N_2473,N_1141,N_286);
xor U2474 (N_2474,N_841,N_39);
and U2475 (N_2475,N_291,N_272);
nor U2476 (N_2476,N_1444,N_314);
nand U2477 (N_2477,N_765,N_1355);
or U2478 (N_2478,N_17,N_438);
and U2479 (N_2479,N_1496,N_1062);
nand U2480 (N_2480,N_1030,N_1181);
and U2481 (N_2481,N_993,N_1441);
nor U2482 (N_2482,N_973,N_32);
nand U2483 (N_2483,N_941,N_374);
and U2484 (N_2484,N_993,N_1300);
nand U2485 (N_2485,N_931,N_754);
and U2486 (N_2486,N_786,N_915);
xnor U2487 (N_2487,N_967,N_1114);
nand U2488 (N_2488,N_90,N_460);
nor U2489 (N_2489,N_11,N_375);
nor U2490 (N_2490,N_624,N_430);
or U2491 (N_2491,N_183,N_1138);
and U2492 (N_2492,N_941,N_1036);
nor U2493 (N_2493,N_872,N_410);
nor U2494 (N_2494,N_1136,N_307);
and U2495 (N_2495,N_924,N_1275);
or U2496 (N_2496,N_1096,N_665);
and U2497 (N_2497,N_417,N_231);
nand U2498 (N_2498,N_1482,N_732);
nand U2499 (N_2499,N_963,N_321);
and U2500 (N_2500,N_699,N_183);
nand U2501 (N_2501,N_656,N_1184);
and U2502 (N_2502,N_896,N_1088);
nor U2503 (N_2503,N_1347,N_1094);
nor U2504 (N_2504,N_195,N_109);
or U2505 (N_2505,N_1012,N_936);
or U2506 (N_2506,N_914,N_1027);
or U2507 (N_2507,N_347,N_1286);
or U2508 (N_2508,N_1016,N_1217);
nor U2509 (N_2509,N_128,N_935);
nor U2510 (N_2510,N_1315,N_219);
or U2511 (N_2511,N_40,N_567);
nand U2512 (N_2512,N_1066,N_1043);
nor U2513 (N_2513,N_1224,N_1030);
nand U2514 (N_2514,N_1169,N_346);
nand U2515 (N_2515,N_830,N_398);
and U2516 (N_2516,N_146,N_898);
and U2517 (N_2517,N_894,N_225);
nand U2518 (N_2518,N_1419,N_1245);
nor U2519 (N_2519,N_572,N_872);
nand U2520 (N_2520,N_161,N_544);
or U2521 (N_2521,N_11,N_1079);
nor U2522 (N_2522,N_249,N_197);
or U2523 (N_2523,N_163,N_921);
xor U2524 (N_2524,N_941,N_294);
or U2525 (N_2525,N_159,N_66);
nor U2526 (N_2526,N_546,N_693);
or U2527 (N_2527,N_1384,N_72);
nor U2528 (N_2528,N_1082,N_485);
and U2529 (N_2529,N_704,N_414);
nor U2530 (N_2530,N_291,N_315);
and U2531 (N_2531,N_417,N_221);
nor U2532 (N_2532,N_609,N_77);
or U2533 (N_2533,N_1314,N_261);
nand U2534 (N_2534,N_1386,N_1021);
or U2535 (N_2535,N_1031,N_750);
and U2536 (N_2536,N_1434,N_1493);
or U2537 (N_2537,N_440,N_1415);
nor U2538 (N_2538,N_348,N_233);
and U2539 (N_2539,N_14,N_718);
or U2540 (N_2540,N_149,N_1432);
and U2541 (N_2541,N_1211,N_834);
nor U2542 (N_2542,N_410,N_1086);
and U2543 (N_2543,N_1389,N_1022);
xor U2544 (N_2544,N_1235,N_180);
nor U2545 (N_2545,N_908,N_312);
nor U2546 (N_2546,N_651,N_756);
nand U2547 (N_2547,N_735,N_33);
and U2548 (N_2548,N_1495,N_61);
nor U2549 (N_2549,N_506,N_889);
or U2550 (N_2550,N_928,N_1465);
nand U2551 (N_2551,N_120,N_364);
nand U2552 (N_2552,N_1027,N_325);
nor U2553 (N_2553,N_1433,N_749);
xor U2554 (N_2554,N_1187,N_383);
or U2555 (N_2555,N_338,N_472);
nand U2556 (N_2556,N_1403,N_264);
nand U2557 (N_2557,N_150,N_938);
or U2558 (N_2558,N_474,N_950);
nand U2559 (N_2559,N_946,N_1143);
nand U2560 (N_2560,N_64,N_1418);
nor U2561 (N_2561,N_1352,N_390);
or U2562 (N_2562,N_1213,N_922);
nand U2563 (N_2563,N_268,N_1276);
and U2564 (N_2564,N_1034,N_1200);
nor U2565 (N_2565,N_1306,N_1388);
nor U2566 (N_2566,N_1087,N_938);
or U2567 (N_2567,N_205,N_1083);
xnor U2568 (N_2568,N_373,N_20);
nand U2569 (N_2569,N_93,N_764);
nor U2570 (N_2570,N_79,N_1078);
nor U2571 (N_2571,N_737,N_806);
and U2572 (N_2572,N_445,N_1329);
or U2573 (N_2573,N_603,N_961);
nand U2574 (N_2574,N_1236,N_1305);
xnor U2575 (N_2575,N_595,N_1236);
or U2576 (N_2576,N_525,N_937);
nand U2577 (N_2577,N_334,N_704);
and U2578 (N_2578,N_1410,N_1359);
nand U2579 (N_2579,N_868,N_297);
nor U2580 (N_2580,N_1458,N_602);
and U2581 (N_2581,N_957,N_67);
nor U2582 (N_2582,N_314,N_328);
and U2583 (N_2583,N_542,N_885);
nand U2584 (N_2584,N_668,N_783);
or U2585 (N_2585,N_533,N_1456);
nor U2586 (N_2586,N_45,N_415);
or U2587 (N_2587,N_1216,N_321);
or U2588 (N_2588,N_460,N_142);
and U2589 (N_2589,N_1407,N_1390);
nand U2590 (N_2590,N_709,N_823);
nor U2591 (N_2591,N_711,N_248);
nand U2592 (N_2592,N_497,N_1024);
nand U2593 (N_2593,N_281,N_869);
or U2594 (N_2594,N_1218,N_1236);
or U2595 (N_2595,N_975,N_938);
nor U2596 (N_2596,N_123,N_1166);
or U2597 (N_2597,N_1488,N_755);
nand U2598 (N_2598,N_223,N_1122);
or U2599 (N_2599,N_274,N_627);
nor U2600 (N_2600,N_969,N_1142);
nand U2601 (N_2601,N_977,N_1236);
and U2602 (N_2602,N_408,N_1306);
and U2603 (N_2603,N_1048,N_902);
or U2604 (N_2604,N_849,N_198);
and U2605 (N_2605,N_1418,N_1280);
nand U2606 (N_2606,N_423,N_190);
or U2607 (N_2607,N_92,N_787);
and U2608 (N_2608,N_298,N_563);
and U2609 (N_2609,N_620,N_791);
or U2610 (N_2610,N_1079,N_391);
or U2611 (N_2611,N_1008,N_685);
nor U2612 (N_2612,N_1028,N_1267);
or U2613 (N_2613,N_387,N_154);
nor U2614 (N_2614,N_1118,N_377);
or U2615 (N_2615,N_729,N_733);
nand U2616 (N_2616,N_1136,N_305);
or U2617 (N_2617,N_409,N_821);
nand U2618 (N_2618,N_672,N_866);
or U2619 (N_2619,N_933,N_1450);
nand U2620 (N_2620,N_862,N_242);
or U2621 (N_2621,N_301,N_936);
nand U2622 (N_2622,N_1280,N_857);
or U2623 (N_2623,N_97,N_749);
nor U2624 (N_2624,N_444,N_885);
nor U2625 (N_2625,N_1284,N_1227);
and U2626 (N_2626,N_239,N_936);
nor U2627 (N_2627,N_230,N_267);
and U2628 (N_2628,N_86,N_1202);
nor U2629 (N_2629,N_1456,N_1384);
and U2630 (N_2630,N_730,N_897);
and U2631 (N_2631,N_874,N_201);
nor U2632 (N_2632,N_1254,N_1495);
nand U2633 (N_2633,N_593,N_643);
or U2634 (N_2634,N_762,N_1053);
or U2635 (N_2635,N_1309,N_1258);
nor U2636 (N_2636,N_1170,N_772);
nor U2637 (N_2637,N_179,N_1063);
nand U2638 (N_2638,N_1491,N_1489);
and U2639 (N_2639,N_925,N_1016);
or U2640 (N_2640,N_466,N_1313);
and U2641 (N_2641,N_1124,N_873);
or U2642 (N_2642,N_1201,N_275);
nand U2643 (N_2643,N_353,N_1177);
nor U2644 (N_2644,N_444,N_1061);
nand U2645 (N_2645,N_900,N_410);
nor U2646 (N_2646,N_1109,N_1170);
nor U2647 (N_2647,N_854,N_1390);
nand U2648 (N_2648,N_845,N_390);
nor U2649 (N_2649,N_555,N_991);
nand U2650 (N_2650,N_632,N_941);
nor U2651 (N_2651,N_1336,N_1487);
nand U2652 (N_2652,N_1299,N_275);
nand U2653 (N_2653,N_1391,N_586);
or U2654 (N_2654,N_705,N_1123);
nor U2655 (N_2655,N_1483,N_452);
and U2656 (N_2656,N_583,N_3);
or U2657 (N_2657,N_167,N_619);
nand U2658 (N_2658,N_633,N_301);
nor U2659 (N_2659,N_365,N_62);
or U2660 (N_2660,N_603,N_963);
nand U2661 (N_2661,N_453,N_808);
or U2662 (N_2662,N_1327,N_651);
or U2663 (N_2663,N_1317,N_138);
or U2664 (N_2664,N_1490,N_740);
or U2665 (N_2665,N_82,N_485);
nor U2666 (N_2666,N_418,N_1264);
or U2667 (N_2667,N_711,N_1145);
or U2668 (N_2668,N_143,N_872);
nor U2669 (N_2669,N_631,N_663);
nor U2670 (N_2670,N_868,N_1133);
or U2671 (N_2671,N_1060,N_852);
and U2672 (N_2672,N_1459,N_258);
nand U2673 (N_2673,N_570,N_1219);
nand U2674 (N_2674,N_543,N_448);
and U2675 (N_2675,N_1391,N_340);
and U2676 (N_2676,N_747,N_1284);
nand U2677 (N_2677,N_1350,N_374);
and U2678 (N_2678,N_232,N_1423);
or U2679 (N_2679,N_571,N_561);
nand U2680 (N_2680,N_108,N_1118);
nand U2681 (N_2681,N_302,N_552);
nand U2682 (N_2682,N_1135,N_526);
nor U2683 (N_2683,N_24,N_394);
or U2684 (N_2684,N_717,N_744);
nand U2685 (N_2685,N_526,N_1088);
nor U2686 (N_2686,N_1116,N_95);
nand U2687 (N_2687,N_698,N_61);
and U2688 (N_2688,N_1071,N_1164);
and U2689 (N_2689,N_1038,N_687);
nor U2690 (N_2690,N_1390,N_1262);
nand U2691 (N_2691,N_90,N_419);
nor U2692 (N_2692,N_802,N_496);
nor U2693 (N_2693,N_800,N_193);
or U2694 (N_2694,N_1080,N_1291);
nand U2695 (N_2695,N_477,N_1179);
nand U2696 (N_2696,N_802,N_316);
or U2697 (N_2697,N_444,N_249);
nor U2698 (N_2698,N_1351,N_543);
and U2699 (N_2699,N_720,N_407);
or U2700 (N_2700,N_195,N_276);
and U2701 (N_2701,N_502,N_764);
or U2702 (N_2702,N_1176,N_202);
nor U2703 (N_2703,N_1122,N_1);
nor U2704 (N_2704,N_1024,N_544);
nor U2705 (N_2705,N_489,N_216);
and U2706 (N_2706,N_480,N_1332);
nor U2707 (N_2707,N_927,N_660);
nand U2708 (N_2708,N_1287,N_631);
nand U2709 (N_2709,N_1270,N_111);
or U2710 (N_2710,N_1015,N_324);
nand U2711 (N_2711,N_500,N_590);
nand U2712 (N_2712,N_1372,N_1400);
nand U2713 (N_2713,N_605,N_58);
nand U2714 (N_2714,N_967,N_668);
nor U2715 (N_2715,N_213,N_1232);
or U2716 (N_2716,N_643,N_99);
or U2717 (N_2717,N_196,N_877);
or U2718 (N_2718,N_1068,N_1193);
or U2719 (N_2719,N_995,N_512);
nor U2720 (N_2720,N_448,N_1129);
or U2721 (N_2721,N_1263,N_983);
nor U2722 (N_2722,N_294,N_29);
or U2723 (N_2723,N_194,N_1491);
nand U2724 (N_2724,N_1268,N_1128);
nor U2725 (N_2725,N_887,N_101);
nand U2726 (N_2726,N_1135,N_1311);
or U2727 (N_2727,N_1322,N_124);
and U2728 (N_2728,N_696,N_429);
nand U2729 (N_2729,N_839,N_1282);
and U2730 (N_2730,N_45,N_871);
or U2731 (N_2731,N_745,N_348);
or U2732 (N_2732,N_543,N_1201);
and U2733 (N_2733,N_1243,N_254);
and U2734 (N_2734,N_1312,N_55);
nor U2735 (N_2735,N_1114,N_595);
nor U2736 (N_2736,N_1147,N_793);
xor U2737 (N_2737,N_259,N_911);
and U2738 (N_2738,N_1233,N_1104);
and U2739 (N_2739,N_230,N_176);
or U2740 (N_2740,N_245,N_593);
or U2741 (N_2741,N_1449,N_719);
and U2742 (N_2742,N_488,N_1376);
or U2743 (N_2743,N_572,N_302);
and U2744 (N_2744,N_1296,N_1014);
or U2745 (N_2745,N_894,N_619);
nand U2746 (N_2746,N_771,N_1364);
and U2747 (N_2747,N_394,N_886);
nand U2748 (N_2748,N_1250,N_425);
nand U2749 (N_2749,N_1444,N_1404);
nand U2750 (N_2750,N_913,N_101);
and U2751 (N_2751,N_526,N_141);
or U2752 (N_2752,N_1306,N_62);
or U2753 (N_2753,N_1159,N_218);
or U2754 (N_2754,N_1392,N_298);
nand U2755 (N_2755,N_97,N_606);
and U2756 (N_2756,N_224,N_919);
nand U2757 (N_2757,N_358,N_135);
nand U2758 (N_2758,N_1049,N_1454);
nor U2759 (N_2759,N_489,N_661);
or U2760 (N_2760,N_754,N_1133);
or U2761 (N_2761,N_635,N_1043);
or U2762 (N_2762,N_621,N_1393);
or U2763 (N_2763,N_1114,N_347);
and U2764 (N_2764,N_989,N_769);
and U2765 (N_2765,N_70,N_1330);
xor U2766 (N_2766,N_1080,N_348);
nand U2767 (N_2767,N_1065,N_24);
or U2768 (N_2768,N_595,N_137);
and U2769 (N_2769,N_965,N_464);
nor U2770 (N_2770,N_753,N_352);
nand U2771 (N_2771,N_304,N_1296);
xor U2772 (N_2772,N_1482,N_355);
nand U2773 (N_2773,N_922,N_891);
or U2774 (N_2774,N_210,N_697);
and U2775 (N_2775,N_163,N_1374);
and U2776 (N_2776,N_1264,N_600);
nand U2777 (N_2777,N_1096,N_559);
nor U2778 (N_2778,N_1097,N_1016);
nor U2779 (N_2779,N_31,N_34);
nor U2780 (N_2780,N_628,N_141);
nor U2781 (N_2781,N_74,N_904);
nor U2782 (N_2782,N_1191,N_1129);
or U2783 (N_2783,N_440,N_73);
or U2784 (N_2784,N_1331,N_666);
nor U2785 (N_2785,N_907,N_154);
xor U2786 (N_2786,N_1158,N_393);
and U2787 (N_2787,N_927,N_1457);
or U2788 (N_2788,N_922,N_927);
or U2789 (N_2789,N_759,N_1266);
and U2790 (N_2790,N_817,N_687);
nor U2791 (N_2791,N_1362,N_814);
and U2792 (N_2792,N_1119,N_1185);
nand U2793 (N_2793,N_1497,N_1140);
nor U2794 (N_2794,N_906,N_505);
or U2795 (N_2795,N_1497,N_1204);
and U2796 (N_2796,N_1288,N_664);
nand U2797 (N_2797,N_1013,N_115);
nor U2798 (N_2798,N_542,N_1395);
and U2799 (N_2799,N_324,N_781);
nor U2800 (N_2800,N_158,N_302);
nor U2801 (N_2801,N_576,N_608);
or U2802 (N_2802,N_1390,N_93);
nor U2803 (N_2803,N_945,N_223);
nor U2804 (N_2804,N_1036,N_675);
nand U2805 (N_2805,N_1414,N_292);
and U2806 (N_2806,N_210,N_97);
nor U2807 (N_2807,N_844,N_1345);
and U2808 (N_2808,N_391,N_415);
xnor U2809 (N_2809,N_1265,N_714);
or U2810 (N_2810,N_1272,N_552);
nor U2811 (N_2811,N_1487,N_595);
and U2812 (N_2812,N_362,N_379);
nor U2813 (N_2813,N_1383,N_1278);
or U2814 (N_2814,N_522,N_696);
or U2815 (N_2815,N_737,N_730);
nand U2816 (N_2816,N_1290,N_286);
nor U2817 (N_2817,N_470,N_979);
nor U2818 (N_2818,N_1203,N_564);
or U2819 (N_2819,N_89,N_671);
or U2820 (N_2820,N_1209,N_741);
or U2821 (N_2821,N_1106,N_964);
or U2822 (N_2822,N_569,N_1386);
nand U2823 (N_2823,N_406,N_1234);
xnor U2824 (N_2824,N_421,N_241);
or U2825 (N_2825,N_925,N_852);
and U2826 (N_2826,N_689,N_219);
nand U2827 (N_2827,N_205,N_649);
and U2828 (N_2828,N_1294,N_1261);
or U2829 (N_2829,N_376,N_475);
nand U2830 (N_2830,N_1373,N_215);
nor U2831 (N_2831,N_781,N_925);
nor U2832 (N_2832,N_818,N_458);
or U2833 (N_2833,N_522,N_1021);
or U2834 (N_2834,N_669,N_899);
and U2835 (N_2835,N_681,N_1029);
and U2836 (N_2836,N_893,N_1037);
and U2837 (N_2837,N_390,N_130);
and U2838 (N_2838,N_244,N_1391);
or U2839 (N_2839,N_777,N_1226);
and U2840 (N_2840,N_565,N_1086);
nor U2841 (N_2841,N_1220,N_215);
nand U2842 (N_2842,N_859,N_301);
nor U2843 (N_2843,N_553,N_181);
nor U2844 (N_2844,N_758,N_769);
and U2845 (N_2845,N_672,N_1209);
or U2846 (N_2846,N_1140,N_1336);
nor U2847 (N_2847,N_785,N_1353);
nor U2848 (N_2848,N_294,N_1322);
nor U2849 (N_2849,N_755,N_819);
and U2850 (N_2850,N_657,N_507);
nor U2851 (N_2851,N_658,N_885);
or U2852 (N_2852,N_846,N_877);
nand U2853 (N_2853,N_1460,N_35);
and U2854 (N_2854,N_255,N_125);
and U2855 (N_2855,N_1368,N_757);
nand U2856 (N_2856,N_142,N_565);
and U2857 (N_2857,N_178,N_1459);
nor U2858 (N_2858,N_1124,N_9);
and U2859 (N_2859,N_211,N_356);
or U2860 (N_2860,N_228,N_561);
or U2861 (N_2861,N_154,N_1197);
nand U2862 (N_2862,N_498,N_695);
and U2863 (N_2863,N_107,N_914);
or U2864 (N_2864,N_753,N_1406);
or U2865 (N_2865,N_1157,N_1091);
and U2866 (N_2866,N_402,N_588);
or U2867 (N_2867,N_432,N_1255);
nor U2868 (N_2868,N_490,N_570);
and U2869 (N_2869,N_504,N_547);
nor U2870 (N_2870,N_1020,N_1336);
nor U2871 (N_2871,N_1431,N_847);
or U2872 (N_2872,N_367,N_1113);
nor U2873 (N_2873,N_569,N_1324);
nand U2874 (N_2874,N_1349,N_1055);
nor U2875 (N_2875,N_1446,N_242);
nor U2876 (N_2876,N_31,N_1185);
nand U2877 (N_2877,N_1178,N_513);
or U2878 (N_2878,N_129,N_742);
or U2879 (N_2879,N_870,N_370);
nor U2880 (N_2880,N_1075,N_473);
and U2881 (N_2881,N_372,N_1283);
nand U2882 (N_2882,N_1204,N_872);
and U2883 (N_2883,N_54,N_208);
or U2884 (N_2884,N_138,N_769);
and U2885 (N_2885,N_891,N_609);
nor U2886 (N_2886,N_411,N_871);
nor U2887 (N_2887,N_799,N_335);
or U2888 (N_2888,N_739,N_1057);
nor U2889 (N_2889,N_90,N_357);
or U2890 (N_2890,N_528,N_341);
nand U2891 (N_2891,N_619,N_6);
nor U2892 (N_2892,N_559,N_474);
and U2893 (N_2893,N_181,N_1402);
nand U2894 (N_2894,N_1465,N_579);
and U2895 (N_2895,N_81,N_236);
or U2896 (N_2896,N_1243,N_161);
or U2897 (N_2897,N_1461,N_530);
nand U2898 (N_2898,N_1,N_1119);
or U2899 (N_2899,N_1321,N_567);
nand U2900 (N_2900,N_191,N_1099);
nand U2901 (N_2901,N_352,N_26);
nand U2902 (N_2902,N_1340,N_1342);
or U2903 (N_2903,N_329,N_266);
nor U2904 (N_2904,N_230,N_1244);
nand U2905 (N_2905,N_1189,N_1085);
and U2906 (N_2906,N_1379,N_822);
and U2907 (N_2907,N_252,N_941);
nand U2908 (N_2908,N_183,N_952);
nand U2909 (N_2909,N_1309,N_647);
and U2910 (N_2910,N_337,N_741);
or U2911 (N_2911,N_318,N_811);
or U2912 (N_2912,N_724,N_1413);
and U2913 (N_2913,N_1181,N_1474);
and U2914 (N_2914,N_939,N_382);
nand U2915 (N_2915,N_414,N_1174);
nand U2916 (N_2916,N_414,N_626);
nand U2917 (N_2917,N_183,N_631);
nand U2918 (N_2918,N_998,N_1392);
xor U2919 (N_2919,N_186,N_224);
and U2920 (N_2920,N_836,N_833);
or U2921 (N_2921,N_132,N_324);
and U2922 (N_2922,N_819,N_980);
or U2923 (N_2923,N_575,N_514);
or U2924 (N_2924,N_1096,N_1371);
nand U2925 (N_2925,N_331,N_544);
nor U2926 (N_2926,N_1298,N_421);
xor U2927 (N_2927,N_365,N_472);
and U2928 (N_2928,N_205,N_840);
and U2929 (N_2929,N_1328,N_357);
nand U2930 (N_2930,N_41,N_844);
or U2931 (N_2931,N_648,N_176);
nand U2932 (N_2932,N_953,N_466);
or U2933 (N_2933,N_67,N_250);
nor U2934 (N_2934,N_615,N_282);
nand U2935 (N_2935,N_713,N_1082);
nand U2936 (N_2936,N_291,N_541);
nor U2937 (N_2937,N_881,N_907);
nor U2938 (N_2938,N_1112,N_1113);
or U2939 (N_2939,N_839,N_730);
nand U2940 (N_2940,N_1459,N_1164);
nor U2941 (N_2941,N_617,N_465);
or U2942 (N_2942,N_416,N_417);
or U2943 (N_2943,N_939,N_280);
nor U2944 (N_2944,N_1434,N_634);
or U2945 (N_2945,N_269,N_707);
nor U2946 (N_2946,N_39,N_1278);
and U2947 (N_2947,N_85,N_994);
nor U2948 (N_2948,N_762,N_285);
nor U2949 (N_2949,N_254,N_280);
and U2950 (N_2950,N_223,N_368);
and U2951 (N_2951,N_13,N_756);
nand U2952 (N_2952,N_667,N_449);
nor U2953 (N_2953,N_703,N_1122);
nor U2954 (N_2954,N_493,N_939);
nor U2955 (N_2955,N_1099,N_1457);
or U2956 (N_2956,N_1164,N_695);
and U2957 (N_2957,N_966,N_1152);
nand U2958 (N_2958,N_843,N_824);
or U2959 (N_2959,N_581,N_367);
nor U2960 (N_2960,N_1324,N_918);
and U2961 (N_2961,N_568,N_117);
nand U2962 (N_2962,N_495,N_1426);
and U2963 (N_2963,N_695,N_280);
nand U2964 (N_2964,N_176,N_1086);
or U2965 (N_2965,N_987,N_1415);
and U2966 (N_2966,N_438,N_379);
nor U2967 (N_2967,N_342,N_1276);
xnor U2968 (N_2968,N_1204,N_305);
and U2969 (N_2969,N_880,N_328);
nand U2970 (N_2970,N_1146,N_184);
and U2971 (N_2971,N_739,N_1123);
and U2972 (N_2972,N_513,N_914);
or U2973 (N_2973,N_282,N_252);
nand U2974 (N_2974,N_659,N_147);
nor U2975 (N_2975,N_374,N_912);
nor U2976 (N_2976,N_1405,N_1227);
and U2977 (N_2977,N_872,N_469);
nand U2978 (N_2978,N_882,N_671);
nand U2979 (N_2979,N_372,N_1118);
nor U2980 (N_2980,N_222,N_855);
and U2981 (N_2981,N_1117,N_880);
nor U2982 (N_2982,N_385,N_177);
nor U2983 (N_2983,N_921,N_603);
nand U2984 (N_2984,N_105,N_296);
nor U2985 (N_2985,N_579,N_1357);
nand U2986 (N_2986,N_546,N_922);
and U2987 (N_2987,N_487,N_181);
and U2988 (N_2988,N_122,N_301);
and U2989 (N_2989,N_1225,N_275);
and U2990 (N_2990,N_166,N_656);
nand U2991 (N_2991,N_1418,N_1088);
or U2992 (N_2992,N_869,N_393);
nand U2993 (N_2993,N_389,N_652);
or U2994 (N_2994,N_1178,N_294);
and U2995 (N_2995,N_102,N_696);
and U2996 (N_2996,N_1169,N_733);
nor U2997 (N_2997,N_398,N_968);
nand U2998 (N_2998,N_1453,N_51);
nor U2999 (N_2999,N_463,N_687);
or U3000 (N_3000,N_1693,N_1845);
nand U3001 (N_3001,N_2727,N_1515);
and U3002 (N_3002,N_2637,N_1547);
nor U3003 (N_3003,N_2776,N_2736);
and U3004 (N_3004,N_1781,N_2651);
nor U3005 (N_3005,N_2300,N_2977);
nor U3006 (N_3006,N_1881,N_2225);
nor U3007 (N_3007,N_2660,N_2648);
and U3008 (N_3008,N_2869,N_1996);
nand U3009 (N_3009,N_1862,N_2572);
nand U3010 (N_3010,N_2939,N_2148);
and U3011 (N_3011,N_1920,N_2583);
nand U3012 (N_3012,N_2042,N_2859);
nor U3013 (N_3013,N_1840,N_2856);
nand U3014 (N_3014,N_2622,N_2885);
nor U3015 (N_3015,N_2232,N_1827);
and U3016 (N_3016,N_2849,N_2184);
nand U3017 (N_3017,N_2697,N_2355);
nand U3018 (N_3018,N_2101,N_2076);
or U3019 (N_3019,N_2255,N_2978);
nand U3020 (N_3020,N_2009,N_2417);
and U3021 (N_3021,N_2965,N_2383);
nand U3022 (N_3022,N_2201,N_2274);
nor U3023 (N_3023,N_1697,N_2593);
or U3024 (N_3024,N_2342,N_2025);
nor U3025 (N_3025,N_2372,N_1835);
and U3026 (N_3026,N_1832,N_2610);
or U3027 (N_3027,N_1704,N_2751);
or U3028 (N_3028,N_2282,N_1662);
nor U3029 (N_3029,N_2813,N_1619);
or U3030 (N_3030,N_2035,N_1877);
or U3031 (N_3031,N_2334,N_2363);
nand U3032 (N_3032,N_2411,N_1533);
and U3033 (N_3033,N_1570,N_2457);
and U3034 (N_3034,N_1931,N_1673);
nand U3035 (N_3035,N_2440,N_2008);
nor U3036 (N_3036,N_1701,N_2698);
nand U3037 (N_3037,N_1597,N_1789);
nand U3038 (N_3038,N_2799,N_2481);
nor U3039 (N_3039,N_1512,N_2022);
nor U3040 (N_3040,N_1698,N_1988);
nor U3041 (N_3041,N_2190,N_2807);
and U3042 (N_3042,N_2812,N_1747);
nor U3043 (N_3043,N_2345,N_1984);
or U3044 (N_3044,N_2344,N_1696);
nand U3045 (N_3045,N_1623,N_2012);
nand U3046 (N_3046,N_2587,N_2559);
or U3047 (N_3047,N_2681,N_2360);
nand U3048 (N_3048,N_2853,N_2191);
xor U3049 (N_3049,N_2915,N_2724);
and U3050 (N_3050,N_2186,N_1686);
nand U3051 (N_3051,N_1678,N_1858);
and U3052 (N_3052,N_2485,N_2100);
nand U3053 (N_3053,N_1782,N_2600);
and U3054 (N_3054,N_2316,N_2424);
nor U3055 (N_3055,N_1598,N_2384);
and U3056 (N_3056,N_2074,N_2983);
nand U3057 (N_3057,N_1586,N_2889);
or U3058 (N_3058,N_2548,N_2431);
and U3059 (N_3059,N_1962,N_2606);
and U3060 (N_3060,N_2828,N_2373);
or U3061 (N_3061,N_2228,N_2013);
and U3062 (N_3062,N_1687,N_1897);
or U3063 (N_3063,N_2341,N_2421);
and U3064 (N_3064,N_1502,N_2140);
or U3065 (N_3065,N_1611,N_2602);
and U3066 (N_3066,N_1749,N_1960);
or U3067 (N_3067,N_2445,N_1938);
nor U3068 (N_3068,N_1946,N_1581);
or U3069 (N_3069,N_2735,N_2864);
nand U3070 (N_3070,N_2541,N_2033);
or U3071 (N_3071,N_1596,N_2638);
or U3072 (N_3072,N_2375,N_2512);
or U3073 (N_3073,N_2410,N_2798);
or U3074 (N_3074,N_2197,N_2540);
or U3075 (N_3075,N_2204,N_2497);
xnor U3076 (N_3076,N_1552,N_2888);
nor U3077 (N_3077,N_2611,N_2487);
nor U3078 (N_3078,N_1731,N_2133);
or U3079 (N_3079,N_2361,N_2507);
or U3080 (N_3080,N_2510,N_1806);
nor U3081 (N_3081,N_2745,N_1944);
or U3082 (N_3082,N_1794,N_1854);
and U3083 (N_3083,N_2332,N_2787);
nand U3084 (N_3084,N_2784,N_2774);
nand U3085 (N_3085,N_2967,N_2783);
or U3086 (N_3086,N_1966,N_2832);
nor U3087 (N_3087,N_2511,N_1913);
and U3088 (N_3088,N_2021,N_2295);
xor U3089 (N_3089,N_2720,N_2272);
nand U3090 (N_3090,N_2508,N_2224);
nand U3091 (N_3091,N_2716,N_2974);
or U3092 (N_3092,N_1742,N_1824);
nor U3093 (N_3093,N_1764,N_2273);
xor U3094 (N_3094,N_2881,N_1648);
nor U3095 (N_3095,N_2119,N_1868);
nor U3096 (N_3096,N_2525,N_1879);
nor U3097 (N_3097,N_2390,N_2396);
nand U3098 (N_3098,N_1580,N_2820);
nand U3099 (N_3099,N_2044,N_2125);
or U3100 (N_3100,N_2609,N_1819);
or U3101 (N_3101,N_2934,N_1923);
and U3102 (N_3102,N_2114,N_2176);
and U3103 (N_3103,N_2854,N_2712);
and U3104 (N_3104,N_2909,N_2839);
nand U3105 (N_3105,N_2953,N_2605);
nand U3106 (N_3106,N_2115,N_2924);
nand U3107 (N_3107,N_1539,N_2450);
and U3108 (N_3108,N_2922,N_2601);
nand U3109 (N_3109,N_2654,N_2566);
nor U3110 (N_3110,N_2756,N_1573);
or U3111 (N_3111,N_2208,N_2171);
nor U3112 (N_3112,N_2950,N_1759);
or U3113 (N_3113,N_2290,N_2704);
nor U3114 (N_3114,N_1892,N_1994);
or U3115 (N_3115,N_2092,N_1884);
or U3116 (N_3116,N_1604,N_2349);
or U3117 (N_3117,N_2781,N_2629);
nand U3118 (N_3118,N_2843,N_2452);
nor U3119 (N_3119,N_2242,N_2183);
or U3120 (N_3120,N_1963,N_2376);
nand U3121 (N_3121,N_2442,N_2683);
nor U3122 (N_3122,N_2049,N_2509);
nor U3123 (N_3123,N_2659,N_2011);
nor U3124 (N_3124,N_2844,N_2283);
nor U3125 (N_3125,N_2136,N_1836);
nand U3126 (N_3126,N_1980,N_2918);
and U3127 (N_3127,N_2858,N_2573);
or U3128 (N_3128,N_2796,N_1737);
nor U3129 (N_3129,N_2210,N_2019);
nand U3130 (N_3130,N_2625,N_1866);
nor U3131 (N_3131,N_2589,N_2229);
xnor U3132 (N_3132,N_1636,N_2066);
nand U3133 (N_3133,N_1997,N_2879);
or U3134 (N_3134,N_2532,N_2718);
nand U3135 (N_3135,N_2180,N_2563);
and U3136 (N_3136,N_2945,N_2205);
and U3137 (N_3137,N_2760,N_2526);
or U3138 (N_3138,N_1642,N_1799);
nor U3139 (N_3139,N_1633,N_1930);
nor U3140 (N_3140,N_1525,N_2514);
or U3141 (N_3141,N_1763,N_2122);
or U3142 (N_3142,N_2539,N_2579);
or U3143 (N_3143,N_2407,N_2494);
xor U3144 (N_3144,N_2673,N_2112);
nand U3145 (N_3145,N_2169,N_1788);
or U3146 (N_3146,N_1550,N_1865);
nor U3147 (N_3147,N_2362,N_2422);
or U3148 (N_3148,N_2144,N_2182);
nand U3149 (N_3149,N_2824,N_2585);
nand U3150 (N_3150,N_1720,N_2623);
and U3151 (N_3151,N_1715,N_2595);
nor U3152 (N_3152,N_2391,N_2527);
and U3153 (N_3153,N_1625,N_1891);
nor U3154 (N_3154,N_2126,N_2364);
or U3155 (N_3155,N_1679,N_2482);
and U3156 (N_3156,N_2367,N_2048);
nor U3157 (N_3157,N_2250,N_2430);
nand U3158 (N_3158,N_2470,N_1758);
nor U3159 (N_3159,N_1851,N_1902);
nand U3160 (N_3160,N_1668,N_2840);
and U3161 (N_3161,N_1766,N_2314);
xnor U3162 (N_3162,N_1707,N_1859);
nand U3163 (N_3163,N_2371,N_2468);
nand U3164 (N_3164,N_1807,N_1989);
nand U3165 (N_3165,N_1834,N_2218);
nand U3166 (N_3166,N_2018,N_2956);
and U3167 (N_3167,N_2621,N_1936);
nor U3168 (N_3168,N_1875,N_2071);
nor U3169 (N_3169,N_2663,N_2203);
or U3170 (N_3170,N_1755,N_1712);
nand U3171 (N_3171,N_2435,N_1510);
nor U3172 (N_3172,N_2002,N_2645);
or U3173 (N_3173,N_2237,N_2121);
or U3174 (N_3174,N_2646,N_2343);
or U3175 (N_3175,N_2916,N_1922);
nand U3176 (N_3176,N_1926,N_2976);
and U3177 (N_3177,N_2175,N_2168);
and U3178 (N_3178,N_2240,N_2016);
or U3179 (N_3179,N_2780,N_1503);
nor U3180 (N_3180,N_2634,N_1752);
or U3181 (N_3181,N_2165,N_1878);
nand U3182 (N_3182,N_2249,N_2519);
and U3183 (N_3183,N_2238,N_1847);
nor U3184 (N_3184,N_1864,N_1762);
or U3185 (N_3185,N_1514,N_2528);
nor U3186 (N_3186,N_2944,N_2617);
and U3187 (N_3187,N_2065,N_2664);
nand U3188 (N_3188,N_1815,N_1703);
nor U3189 (N_3189,N_2878,N_2117);
or U3190 (N_3190,N_2192,N_2919);
and U3191 (N_3191,N_2586,N_1725);
nand U3192 (N_3192,N_1925,N_2198);
or U3193 (N_3193,N_2116,N_2836);
nor U3194 (N_3194,N_1757,N_1970);
nor U3195 (N_3195,N_2801,N_1684);
and U3196 (N_3196,N_2301,N_2276);
or U3197 (N_3197,N_2159,N_1695);
nor U3198 (N_3198,N_2336,N_1956);
or U3199 (N_3199,N_1869,N_2303);
and U3200 (N_3200,N_1813,N_1765);
nor U3201 (N_3201,N_2026,N_2231);
nor U3202 (N_3202,N_1903,N_2340);
or U3203 (N_3203,N_2725,N_2335);
or U3204 (N_3204,N_2694,N_2177);
or U3205 (N_3205,N_2767,N_1831);
nand U3206 (N_3206,N_2489,N_2146);
or U3207 (N_3207,N_2568,N_2642);
and U3208 (N_3208,N_2439,N_1537);
nor U3209 (N_3209,N_2739,N_2810);
nand U3210 (N_3210,N_2260,N_2848);
nor U3211 (N_3211,N_2505,N_2469);
and U3212 (N_3212,N_1805,N_1954);
and U3213 (N_3213,N_1846,N_2317);
nor U3214 (N_3214,N_2678,N_2748);
or U3215 (N_3215,N_2986,N_2731);
and U3216 (N_3216,N_1981,N_1932);
or U3217 (N_3217,N_2216,N_1711);
nand U3218 (N_3218,N_1561,N_2661);
or U3219 (N_3219,N_1934,N_2128);
xor U3220 (N_3220,N_1803,N_1928);
nor U3221 (N_3221,N_1850,N_1738);
nand U3222 (N_3222,N_2746,N_2754);
and U3223 (N_3223,N_2517,N_2102);
nor U3224 (N_3224,N_2105,N_2196);
nor U3225 (N_3225,N_2211,N_1826);
nand U3226 (N_3226,N_2814,N_2688);
and U3227 (N_3227,N_2329,N_2571);
nand U3228 (N_3228,N_2912,N_1706);
nor U3229 (N_3229,N_2130,N_2368);
or U3230 (N_3230,N_1540,N_2577);
nor U3231 (N_3231,N_1509,N_2719);
nand U3232 (N_3232,N_1993,N_2486);
nor U3233 (N_3233,N_1987,N_2330);
and U3234 (N_3234,N_2474,N_2775);
or U3235 (N_3235,N_2996,N_1553);
and U3236 (N_3236,N_2394,N_2941);
or U3237 (N_3237,N_2308,N_2374);
or U3238 (N_3238,N_2319,N_1820);
and U3239 (N_3239,N_2138,N_2312);
nand U3240 (N_3240,N_2952,N_1817);
or U3241 (N_3241,N_2728,N_2914);
nor U3242 (N_3242,N_2834,N_1556);
and U3243 (N_3243,N_1841,N_1719);
nand U3244 (N_3244,N_2706,N_2428);
nor U3245 (N_3245,N_1554,N_1739);
nor U3246 (N_3246,N_2294,N_2451);
xnor U3247 (N_3247,N_2955,N_1535);
xnor U3248 (N_3248,N_2655,N_2679);
or U3249 (N_3249,N_1965,N_2045);
nor U3250 (N_3250,N_2292,N_2789);
nand U3251 (N_3251,N_2931,N_2630);
xor U3252 (N_3252,N_2772,N_1898);
nand U3253 (N_3253,N_1669,N_1816);
and U3254 (N_3254,N_1584,N_2705);
and U3255 (N_3255,N_1685,N_2708);
nor U3256 (N_3256,N_1671,N_2369);
nor U3257 (N_3257,N_1768,N_2682);
and U3258 (N_3258,N_1917,N_2553);
or U3259 (N_3259,N_1880,N_2433);
and U3260 (N_3260,N_2825,N_1951);
nor U3261 (N_3261,N_2929,N_2555);
or U3262 (N_3262,N_1750,N_2506);
and U3263 (N_3263,N_1569,N_2263);
or U3264 (N_3264,N_2271,N_2173);
or U3265 (N_3265,N_2790,N_2741);
nor U3266 (N_3266,N_2906,N_2010);
or U3267 (N_3267,N_2608,N_2419);
or U3268 (N_3268,N_2083,N_2932);
and U3269 (N_3269,N_1772,N_2040);
nand U3270 (N_3270,N_2281,N_2722);
and U3271 (N_3271,N_2403,N_2730);
nor U3272 (N_3272,N_1661,N_2323);
nand U3273 (N_3273,N_2529,N_2804);
or U3274 (N_3274,N_1773,N_1656);
nor U3275 (N_3275,N_1716,N_2518);
nor U3276 (N_3276,N_1967,N_1896);
nand U3277 (N_3277,N_2172,N_1577);
and U3278 (N_3278,N_1982,N_2296);
nor U3279 (N_3279,N_2782,N_1635);
and U3280 (N_3280,N_2761,N_2723);
and U3281 (N_3281,N_2446,N_1943);
nor U3282 (N_3282,N_1659,N_2588);
nor U3283 (N_3283,N_2581,N_2786);
or U3284 (N_3284,N_2151,N_1558);
and U3285 (N_3285,N_1791,N_2027);
nand U3286 (N_3286,N_2620,N_1974);
or U3287 (N_3287,N_2055,N_2147);
and U3288 (N_3288,N_2244,N_2466);
nand U3289 (N_3289,N_2545,N_2594);
or U3290 (N_3290,N_2239,N_1822);
or U3291 (N_3291,N_2656,N_1918);
and U3292 (N_3292,N_1905,N_2156);
nor U3293 (N_3293,N_1948,N_2139);
or U3294 (N_3294,N_2023,N_1955);
and U3295 (N_3295,N_2356,N_2867);
nor U3296 (N_3296,N_2217,N_2614);
or U3297 (N_3297,N_2189,N_2947);
or U3298 (N_3298,N_1833,N_1613);
and U3299 (N_3299,N_1672,N_2456);
nor U3300 (N_3300,N_2835,N_2808);
nor U3301 (N_3301,N_2940,N_2591);
and U3302 (N_3302,N_2079,N_2093);
or U3303 (N_3303,N_2488,N_2596);
nor U3304 (N_3304,N_2875,N_2269);
and U3305 (N_3305,N_1590,N_1830);
nand U3306 (N_3306,N_2465,N_2770);
nor U3307 (N_3307,N_1732,N_2408);
nand U3308 (N_3308,N_2543,N_2521);
nand U3309 (N_3309,N_2153,N_1876);
or U3310 (N_3310,N_2170,N_2414);
or U3311 (N_3311,N_2616,N_1863);
or U3312 (N_3312,N_1904,N_2865);
nor U3313 (N_3313,N_2964,N_1631);
nor U3314 (N_3314,N_1968,N_1802);
nand U3315 (N_3315,N_2366,N_2309);
nor U3316 (N_3316,N_1576,N_1734);
and U3317 (N_3317,N_2546,N_2680);
or U3318 (N_3318,N_2155,N_2973);
nor U3319 (N_3319,N_1658,N_1572);
nor U3320 (N_3320,N_1630,N_2711);
nor U3321 (N_3321,N_1796,N_2753);
nand U3322 (N_3322,N_1829,N_1536);
nand U3323 (N_3323,N_2624,N_2757);
or U3324 (N_3324,N_2473,N_1721);
nand U3325 (N_3325,N_1914,N_1628);
nand U3326 (N_3326,N_2631,N_2351);
and U3327 (N_3327,N_2887,N_2709);
or U3328 (N_3328,N_2851,N_2460);
nand U3329 (N_3329,N_1828,N_2358);
nor U3330 (N_3330,N_1991,N_2993);
nor U3331 (N_3331,N_2975,N_2876);
or U3332 (N_3332,N_1689,N_2462);
or U3333 (N_3333,N_2047,N_1618);
nor U3334 (N_3334,N_1814,N_1614);
nor U3335 (N_3335,N_2202,N_2059);
and U3336 (N_3336,N_2946,N_2406);
or U3337 (N_3337,N_1521,N_2206);
or U3338 (N_3338,N_2884,N_2959);
nand U3339 (N_3339,N_2458,N_1691);
and U3340 (N_3340,N_1971,N_2324);
or U3341 (N_3341,N_1741,N_2693);
or U3342 (N_3342,N_2084,N_2024);
nand U3343 (N_3343,N_1842,N_2253);
nand U3344 (N_3344,N_2692,N_2123);
or U3345 (N_3345,N_2318,N_1637);
or U3346 (N_3346,N_2264,N_1756);
or U3347 (N_3347,N_1735,N_2350);
or U3348 (N_3348,N_1601,N_2393);
nand U3349 (N_3349,N_2998,N_2051);
and U3350 (N_3350,N_1753,N_1795);
and U3351 (N_3351,N_2141,N_1990);
and U3352 (N_3352,N_1651,N_2038);
and U3353 (N_3353,N_1665,N_2326);
or U3354 (N_3354,N_2647,N_2726);
or U3355 (N_3355,N_2615,N_2037);
and U3356 (N_3356,N_2304,N_2041);
nor U3357 (N_3357,N_1770,N_1629);
and U3358 (N_3358,N_2030,N_1513);
nand U3359 (N_3359,N_2972,N_2963);
and U3360 (N_3360,N_1945,N_1942);
nor U3361 (N_3361,N_2277,N_1952);
or U3362 (N_3362,N_2392,N_2522);
and U3363 (N_3363,N_2053,N_2747);
nor U3364 (N_3364,N_2580,N_2826);
nand U3365 (N_3365,N_2467,N_1774);
and U3366 (N_3366,N_1726,N_2052);
or U3367 (N_3367,N_2298,N_2069);
nor U3368 (N_3368,N_2903,N_2305);
and U3369 (N_3369,N_2379,N_1587);
and U3370 (N_3370,N_2299,N_2454);
nand U3371 (N_3371,N_2057,N_2425);
or U3372 (N_3372,N_2199,N_1787);
nand U3373 (N_3373,N_1871,N_2564);
nor U3374 (N_3374,N_1893,N_2310);
nand U3375 (N_3375,N_2759,N_2043);
and U3376 (N_3376,N_1517,N_2890);
nand U3377 (N_3377,N_2385,N_2984);
or U3378 (N_3378,N_1728,N_2740);
nor U3379 (N_3379,N_1873,N_2797);
nand U3380 (N_3380,N_2297,N_2805);
and U3381 (N_3381,N_1560,N_2833);
and U3382 (N_3382,N_2247,N_2056);
and U3383 (N_3383,N_2054,N_2788);
nand U3384 (N_3384,N_1844,N_2426);
nand U3385 (N_3385,N_2910,N_2504);
nor U3386 (N_3386,N_1593,N_2088);
nand U3387 (N_3387,N_1940,N_2448);
nor U3388 (N_3388,N_2951,N_1837);
or U3389 (N_3389,N_2386,N_2491);
xnor U3390 (N_3390,N_2090,N_2077);
nor U3391 (N_3391,N_2652,N_2311);
and U3392 (N_3392,N_1627,N_2154);
or U3393 (N_3393,N_2185,N_2671);
nor U3394 (N_3394,N_2464,N_2662);
or U3395 (N_3395,N_2028,N_2721);
nand U3396 (N_3396,N_1575,N_1709);
nor U3397 (N_3397,N_2653,N_2738);
nand U3398 (N_3398,N_2000,N_1699);
and U3399 (N_3399,N_2483,N_2007);
and U3400 (N_3400,N_2558,N_2937);
nand U3401 (N_3401,N_1592,N_2388);
nand U3402 (N_3402,N_2847,N_1626);
nand U3403 (N_3403,N_1692,N_1901);
nand U3404 (N_3404,N_2067,N_2215);
nor U3405 (N_3405,N_2778,N_2503);
nand U3406 (N_3406,N_2819,N_2441);
nor U3407 (N_3407,N_2872,N_2178);
and U3408 (N_3408,N_2135,N_2870);
nor U3409 (N_3409,N_2905,N_1911);
nor U3410 (N_3410,N_2640,N_2883);
or U3411 (N_3411,N_2766,N_2167);
or U3412 (N_3412,N_2811,N_1978);
or U3413 (N_3413,N_2412,N_2017);
xor U3414 (N_3414,N_2471,N_1999);
nand U3415 (N_3415,N_2286,N_2562);
nor U3416 (N_3416,N_2534,N_1571);
or U3417 (N_3417,N_2254,N_2357);
and U3418 (N_3418,N_2744,N_2124);
or U3419 (N_3419,N_2632,N_2081);
nand U3420 (N_3420,N_2771,N_2795);
nor U3421 (N_3421,N_2677,N_2098);
nor U3422 (N_3422,N_2992,N_2703);
xnor U3423 (N_3423,N_2475,N_1717);
or U3424 (N_3424,N_2911,N_2143);
xnor U3425 (N_3425,N_1508,N_2064);
nor U3426 (N_3426,N_2533,N_1736);
nand U3427 (N_3427,N_2863,N_1524);
or U3428 (N_3428,N_2707,N_2520);
or U3429 (N_3429,N_1983,N_2150);
and U3430 (N_3430,N_1501,N_2821);
and U3431 (N_3431,N_1640,N_2267);
and U3432 (N_3432,N_2641,N_1568);
and U3433 (N_3433,N_2668,N_2644);
nor U3434 (N_3434,N_1910,N_2399);
or U3435 (N_3435,N_1975,N_2603);
and U3436 (N_3436,N_1664,N_2927);
and U3437 (N_3437,N_2499,N_2800);
and U3438 (N_3438,N_2014,N_2338);
and U3439 (N_3439,N_1563,N_2085);
nor U3440 (N_3440,N_1555,N_2275);
nand U3441 (N_3441,N_2188,N_2039);
nand U3442 (N_3442,N_2938,N_1958);
or U3443 (N_3443,N_1793,N_1722);
or U3444 (N_3444,N_2674,N_2315);
nand U3445 (N_3445,N_1634,N_1744);
nand U3446 (N_3446,N_1595,N_1751);
nand U3447 (N_3447,N_2220,N_2666);
or U3448 (N_3448,N_2613,N_2429);
nand U3449 (N_3449,N_2339,N_1780);
or U3450 (N_3450,N_1677,N_1825);
or U3451 (N_3451,N_2401,N_1953);
nor U3452 (N_3452,N_2160,N_2127);
nor U3453 (N_3453,N_2714,N_2221);
and U3454 (N_3454,N_2971,N_2219);
nand U3455 (N_3455,N_2498,N_2930);
and U3456 (N_3456,N_2111,N_2933);
nor U3457 (N_3457,N_2359,N_2413);
and U3458 (N_3458,N_2524,N_2370);
or U3459 (N_3459,N_2427,N_2831);
and U3460 (N_3460,N_2097,N_2104);
or U3461 (N_3461,N_1786,N_1582);
or U3462 (N_3462,N_2068,N_2892);
nand U3463 (N_3463,N_2670,N_2437);
and U3464 (N_3464,N_2248,N_2265);
and U3465 (N_3465,N_2961,N_2841);
or U3466 (N_3466,N_2868,N_2003);
nand U3467 (N_3467,N_1655,N_1972);
nand U3468 (N_3468,N_2837,N_2968);
nand U3469 (N_3469,N_2162,N_1608);
or U3470 (N_3470,N_2762,N_1771);
nor U3471 (N_3471,N_2791,N_2096);
nand U3472 (N_3472,N_2382,N_2434);
nand U3473 (N_3473,N_2346,N_2734);
and U3474 (N_3474,N_2404,N_1516);
or U3475 (N_3475,N_2194,N_2899);
nand U3476 (N_3476,N_1632,N_1578);
or U3477 (N_3477,N_1969,N_1688);
and U3478 (N_3478,N_1700,N_1964);
nor U3479 (N_3479,N_2715,N_1888);
and U3480 (N_3480,N_1562,N_2699);
and U3481 (N_3481,N_2480,N_2236);
or U3482 (N_3482,N_2633,N_1605);
and U3483 (N_3483,N_2389,N_1927);
and U3484 (N_3484,N_1992,N_2113);
xnor U3485 (N_3485,N_1838,N_1589);
nand U3486 (N_3486,N_2377,N_1921);
and U3487 (N_3487,N_1933,N_2894);
or U3488 (N_3488,N_2060,N_2904);
nor U3489 (N_3489,N_1895,N_2686);
and U3490 (N_3490,N_2251,N_1804);
nor U3491 (N_3491,N_2327,N_2307);
nor U3492 (N_3492,N_2597,N_2958);
and U3493 (N_3493,N_2980,N_2667);
nand U3494 (N_3494,N_2880,N_1647);
or U3495 (N_3495,N_2592,N_2561);
nor U3496 (N_3496,N_2365,N_2001);
nor U3497 (N_3497,N_2405,N_1929);
nand U3498 (N_3498,N_1522,N_1823);
nand U3499 (N_3499,N_2179,N_1843);
nor U3500 (N_3500,N_1663,N_2152);
or U3501 (N_3501,N_2502,N_2278);
nand U3502 (N_3502,N_2166,N_2578);
and U3503 (N_3503,N_2322,N_1708);
or U3504 (N_3504,N_2802,N_2006);
nand U3505 (N_3505,N_1542,N_1935);
nand U3506 (N_3506,N_2477,N_1549);
xor U3507 (N_3507,N_1899,N_2855);
nor U3508 (N_3508,N_1616,N_2669);
nor U3509 (N_3509,N_1779,N_2495);
nor U3510 (N_3510,N_1870,N_2628);
or U3511 (N_3511,N_2209,N_2873);
and U3512 (N_3512,N_2400,N_1666);
or U3513 (N_3513,N_2755,N_2779);
or U3514 (N_3514,N_2960,N_2845);
nor U3515 (N_3515,N_2020,N_2576);
or U3516 (N_3516,N_2737,N_2966);
nor U3517 (N_3517,N_2987,N_2957);
nor U3518 (N_3518,N_1546,N_2455);
and U3519 (N_3519,N_2928,N_2157);
nand U3520 (N_3520,N_2423,N_2005);
and U3521 (N_3521,N_2717,N_1585);
or U3522 (N_3522,N_1602,N_1683);
nand U3523 (N_3523,N_2936,N_1518);
or U3524 (N_3524,N_2262,N_1924);
or U3525 (N_3525,N_1775,N_1784);
or U3526 (N_3526,N_2538,N_2823);
nor U3527 (N_3527,N_2773,N_1579);
and U3528 (N_3528,N_1849,N_2015);
nor U3529 (N_3529,N_2459,N_2523);
nor U3530 (N_3530,N_2750,N_2492);
nand U3531 (N_3531,N_1801,N_2550);
or U3532 (N_3532,N_2943,N_1638);
nand U3533 (N_3533,N_2598,N_2061);
and U3534 (N_3534,N_2866,N_1889);
nand U3535 (N_3535,N_1594,N_2073);
nor U3536 (N_3536,N_2891,N_1882);
and U3537 (N_3537,N_1909,N_2710);
or U3538 (N_3538,N_1976,N_2241);
or U3539 (N_3539,N_2920,N_2484);
or U3540 (N_3540,N_1714,N_2266);
xnor U3541 (N_3541,N_2742,N_2627);
and U3542 (N_3542,N_1622,N_1748);
nand U3543 (N_3543,N_1760,N_2415);
and U3544 (N_3544,N_1527,N_1500);
or U3545 (N_3545,N_1855,N_2072);
nor U3546 (N_3546,N_2164,N_1810);
or U3547 (N_3547,N_1519,N_2969);
or U3548 (N_3548,N_1852,N_2676);
or U3549 (N_3549,N_2258,N_2145);
or U3550 (N_3550,N_2650,N_2701);
or U3551 (N_3551,N_2213,N_2733);
and U3552 (N_3552,N_2691,N_1912);
nor U3553 (N_3553,N_1530,N_1643);
and U3554 (N_3554,N_2672,N_1532);
and U3555 (N_3555,N_1937,N_2935);
or U3556 (N_3556,N_1681,N_2395);
or U3557 (N_3557,N_2695,N_1785);
or U3558 (N_3558,N_2226,N_2619);
nor U3559 (N_3559,N_1545,N_2444);
or U3560 (N_3560,N_2900,N_1506);
and U3561 (N_3561,N_2575,N_2129);
and U3562 (N_3562,N_1538,N_1551);
nor U3563 (N_3563,N_2347,N_2768);
and U3564 (N_3564,N_1606,N_1667);
or U3565 (N_3565,N_2142,N_2348);
nor U3566 (N_3566,N_1740,N_2328);
nand U3567 (N_3567,N_2163,N_1727);
nor U3568 (N_3568,N_2785,N_2793);
nor U3569 (N_3569,N_2599,N_2842);
nand U3570 (N_3570,N_2817,N_2689);
xor U3571 (N_3571,N_2861,N_2897);
xor U3572 (N_3572,N_2985,N_1811);
nor U3573 (N_3573,N_2846,N_2063);
nor U3574 (N_3574,N_2942,N_2354);
or U3575 (N_3575,N_2535,N_2320);
or U3576 (N_3576,N_2078,N_2214);
xor U3577 (N_3577,N_2658,N_1950);
or U3578 (N_3578,N_1861,N_1529);
and U3579 (N_3579,N_2569,N_2991);
and U3580 (N_3580,N_2874,N_1653);
and U3581 (N_3581,N_2643,N_1985);
nor U3582 (N_3582,N_1857,N_2871);
xor U3583 (N_3583,N_1541,N_1797);
and U3584 (N_3584,N_2095,N_2416);
nand U3585 (N_3585,N_1557,N_2472);
xnor U3586 (N_3586,N_2252,N_2816);
nor U3587 (N_3587,N_2582,N_1690);
nand U3588 (N_3588,N_2031,N_1959);
and U3589 (N_3589,N_2635,N_2700);
nand U3590 (N_3590,N_2665,N_2261);
xor U3591 (N_3591,N_2554,N_1915);
and U3592 (N_3592,N_2161,N_1949);
or U3593 (N_3593,N_2516,N_2402);
nand U3594 (N_3594,N_2418,N_2898);
or U3595 (N_3595,N_2995,N_2657);
and U3596 (N_3596,N_2907,N_1544);
nand U3597 (N_3597,N_2397,N_2496);
nor U3598 (N_3598,N_2574,N_1961);
or U3599 (N_3599,N_1676,N_2230);
nand U3600 (N_3600,N_1853,N_2752);
nand U3601 (N_3601,N_2926,N_1565);
nand U3602 (N_3602,N_2313,N_2877);
nand U3603 (N_3603,N_1890,N_2565);
nor U3604 (N_3604,N_1939,N_1730);
or U3605 (N_3605,N_2449,N_2536);
and U3606 (N_3606,N_2908,N_2687);
and U3607 (N_3607,N_2062,N_2994);
nand U3608 (N_3608,N_2882,N_1652);
and U3609 (N_3609,N_1543,N_2158);
or U3610 (N_3610,N_2432,N_2438);
and U3611 (N_3611,N_2285,N_1588);
or U3612 (N_3612,N_2109,N_2765);
or U3613 (N_3613,N_1848,N_1523);
nand U3614 (N_3614,N_2988,N_2461);
and U3615 (N_3615,N_1723,N_2193);
nand U3616 (N_3616,N_1887,N_1710);
and U3617 (N_3617,N_1798,N_2763);
nor U3618 (N_3618,N_1610,N_1507);
or U3619 (N_3619,N_1599,N_1657);
or U3620 (N_3620,N_1660,N_1743);
nor U3621 (N_3621,N_2212,N_2293);
and U3622 (N_3622,N_2187,N_2551);
and U3623 (N_3623,N_2749,N_1977);
and U3624 (N_3624,N_2256,N_2381);
nand U3625 (N_3625,N_2029,N_1624);
and U3626 (N_3626,N_1505,N_2792);
and U3627 (N_3627,N_1761,N_1607);
or U3628 (N_3628,N_1800,N_2639);
xnor U3629 (N_3629,N_1729,N_2050);
and U3630 (N_3630,N_2259,N_2769);
xnor U3631 (N_3631,N_1867,N_2557);
and U3632 (N_3632,N_2758,N_2447);
xnor U3633 (N_3633,N_2902,N_2962);
or U3634 (N_3634,N_2531,N_1941);
and U3635 (N_3635,N_2106,N_2118);
nand U3636 (N_3636,N_2378,N_2058);
or U3637 (N_3637,N_1705,N_2289);
or U3638 (N_3638,N_1907,N_2732);
or U3639 (N_3639,N_1548,N_1776);
and U3640 (N_3640,N_1564,N_2291);
and U3641 (N_3641,N_1674,N_2436);
nand U3642 (N_3642,N_1600,N_2590);
nand U3643 (N_3643,N_2091,N_2181);
xnor U3644 (N_3644,N_2777,N_2530);
nor U3645 (N_3645,N_2584,N_2893);
nor U3646 (N_3646,N_1526,N_2453);
nand U3647 (N_3647,N_2287,N_2333);
nand U3648 (N_3648,N_2829,N_1724);
nor U3649 (N_3649,N_2103,N_1769);
nor U3650 (N_3650,N_2479,N_2004);
or U3651 (N_3651,N_2636,N_2321);
and U3652 (N_3652,N_1947,N_2850);
nand U3653 (N_3653,N_2923,N_2982);
or U3654 (N_3654,N_2949,N_1621);
nand U3655 (N_3655,N_2860,N_2702);
or U3656 (N_3656,N_2537,N_1649);
nor U3657 (N_3657,N_1808,N_1583);
or U3658 (N_3658,N_1620,N_1792);
or U3659 (N_3659,N_2852,N_2420);
nor U3660 (N_3660,N_1654,N_1745);
or U3661 (N_3661,N_1998,N_2794);
nor U3662 (N_3662,N_2547,N_1591);
nand U3663 (N_3663,N_1574,N_2925);
or U3664 (N_3664,N_2838,N_2556);
and U3665 (N_3665,N_2567,N_1818);
nand U3666 (N_3666,N_2607,N_2222);
nand U3667 (N_3667,N_2549,N_2094);
nand U3668 (N_3668,N_2207,N_1645);
or U3669 (N_3669,N_2696,N_2743);
and U3670 (N_3670,N_2806,N_2075);
nor U3671 (N_3671,N_2685,N_2087);
and U3672 (N_3672,N_2288,N_1718);
or U3673 (N_3673,N_2352,N_2729);
nor U3674 (N_3674,N_2476,N_2954);
nor U3675 (N_3675,N_2896,N_2513);
or U3676 (N_3676,N_2353,N_1754);
nor U3677 (N_3677,N_2082,N_1872);
or U3678 (N_3678,N_2080,N_1995);
and U3679 (N_3679,N_2764,N_2200);
and U3680 (N_3680,N_2137,N_1839);
nand U3681 (N_3681,N_2233,N_2107);
and U3682 (N_3682,N_2331,N_2544);
nand U3683 (N_3683,N_2120,N_1567);
nor U3684 (N_3684,N_2070,N_1812);
nand U3685 (N_3685,N_2443,N_2234);
and U3686 (N_3686,N_2818,N_2235);
and U3687 (N_3687,N_2246,N_1919);
nand U3688 (N_3688,N_2195,N_1809);
and U3689 (N_3689,N_1986,N_2895);
nor U3690 (N_3690,N_1531,N_2604);
nor U3691 (N_3691,N_2970,N_1680);
nand U3692 (N_3692,N_1746,N_2223);
nor U3693 (N_3693,N_1778,N_2913);
nand U3694 (N_3694,N_2989,N_2257);
or U3695 (N_3695,N_2981,N_2046);
and U3696 (N_3696,N_1520,N_2032);
nor U3697 (N_3697,N_1767,N_1783);
and U3698 (N_3698,N_1566,N_2500);
and U3699 (N_3699,N_2089,N_2245);
nand U3700 (N_3700,N_1639,N_1615);
nand U3701 (N_3701,N_1609,N_2999);
or U3702 (N_3702,N_2570,N_2675);
nand U3703 (N_3703,N_1883,N_1617);
nor U3704 (N_3704,N_2552,N_2132);
or U3705 (N_3705,N_2280,N_1900);
nand U3706 (N_3706,N_1528,N_1957);
and U3707 (N_3707,N_2901,N_2110);
or U3708 (N_3708,N_1894,N_1682);
nor U3709 (N_3709,N_2649,N_1973);
nor U3710 (N_3710,N_2243,N_2990);
and U3711 (N_3711,N_2886,N_2490);
or U3712 (N_3712,N_2917,N_2862);
or U3713 (N_3713,N_2036,N_2387);
nor U3714 (N_3714,N_1713,N_2822);
nor U3715 (N_3715,N_1504,N_1644);
and U3716 (N_3716,N_1641,N_2515);
and U3717 (N_3717,N_2268,N_2149);
nand U3718 (N_3718,N_2134,N_2618);
nor U3719 (N_3719,N_1511,N_1856);
or U3720 (N_3720,N_1733,N_2560);
and U3721 (N_3721,N_2827,N_2398);
nand U3722 (N_3722,N_2325,N_2270);
nand U3723 (N_3723,N_2612,N_2997);
nand U3724 (N_3724,N_1670,N_2086);
and U3725 (N_3725,N_2463,N_2131);
nand U3726 (N_3726,N_2302,N_1790);
or U3727 (N_3727,N_2337,N_2099);
and U3728 (N_3728,N_2108,N_2279);
nor U3729 (N_3729,N_1860,N_1821);
nand U3730 (N_3730,N_2809,N_2478);
and U3731 (N_3731,N_1874,N_2830);
nand U3732 (N_3732,N_2306,N_1603);
or U3733 (N_3733,N_2174,N_1916);
and U3734 (N_3734,N_2626,N_1646);
or U3735 (N_3735,N_1559,N_1885);
nand U3736 (N_3736,N_2690,N_1534);
and U3737 (N_3737,N_2684,N_1908);
nor U3738 (N_3738,N_2815,N_2501);
or U3739 (N_3739,N_2803,N_2857);
nor U3740 (N_3740,N_2713,N_2493);
nor U3741 (N_3741,N_2542,N_1702);
nor U3742 (N_3742,N_2409,N_1979);
or U3743 (N_3743,N_1906,N_1694);
nand U3744 (N_3744,N_2921,N_1612);
xnor U3745 (N_3745,N_2227,N_2284);
xor U3746 (N_3746,N_2380,N_1650);
or U3747 (N_3747,N_1777,N_2979);
or U3748 (N_3748,N_2948,N_1675);
nor U3749 (N_3749,N_2034,N_1886);
and U3750 (N_3750,N_2255,N_2117);
nor U3751 (N_3751,N_1630,N_1711);
nor U3752 (N_3752,N_2820,N_2090);
nor U3753 (N_3753,N_1562,N_1870);
nand U3754 (N_3754,N_2701,N_2728);
nand U3755 (N_3755,N_2287,N_2776);
and U3756 (N_3756,N_2343,N_2052);
and U3757 (N_3757,N_2136,N_1956);
nand U3758 (N_3758,N_1711,N_2301);
nand U3759 (N_3759,N_1966,N_2526);
or U3760 (N_3760,N_1714,N_1947);
or U3761 (N_3761,N_2515,N_2025);
or U3762 (N_3762,N_1629,N_2189);
nand U3763 (N_3763,N_1927,N_2010);
or U3764 (N_3764,N_2802,N_2040);
nand U3765 (N_3765,N_1641,N_1783);
and U3766 (N_3766,N_2926,N_2321);
or U3767 (N_3767,N_1938,N_1762);
nor U3768 (N_3768,N_2334,N_2495);
and U3769 (N_3769,N_1607,N_1907);
nand U3770 (N_3770,N_2380,N_2741);
and U3771 (N_3771,N_1900,N_2840);
nor U3772 (N_3772,N_2463,N_2857);
nor U3773 (N_3773,N_2660,N_2981);
and U3774 (N_3774,N_2693,N_2334);
nor U3775 (N_3775,N_1783,N_2651);
or U3776 (N_3776,N_1553,N_1554);
nor U3777 (N_3777,N_1990,N_2736);
nor U3778 (N_3778,N_2289,N_1774);
or U3779 (N_3779,N_2943,N_1716);
nand U3780 (N_3780,N_2981,N_1961);
and U3781 (N_3781,N_2562,N_1839);
and U3782 (N_3782,N_2997,N_2955);
and U3783 (N_3783,N_2401,N_2848);
nand U3784 (N_3784,N_2523,N_2275);
nand U3785 (N_3785,N_2564,N_2061);
nor U3786 (N_3786,N_2277,N_2127);
nor U3787 (N_3787,N_1760,N_2340);
nor U3788 (N_3788,N_2120,N_2806);
and U3789 (N_3789,N_2809,N_1978);
and U3790 (N_3790,N_1545,N_1955);
or U3791 (N_3791,N_1670,N_2059);
nand U3792 (N_3792,N_1806,N_2402);
or U3793 (N_3793,N_2888,N_2021);
or U3794 (N_3794,N_1782,N_2108);
and U3795 (N_3795,N_1502,N_1722);
and U3796 (N_3796,N_1793,N_2615);
or U3797 (N_3797,N_2315,N_2844);
or U3798 (N_3798,N_1557,N_1848);
and U3799 (N_3799,N_1596,N_2828);
nor U3800 (N_3800,N_1733,N_2078);
nand U3801 (N_3801,N_2303,N_2708);
nor U3802 (N_3802,N_2414,N_2240);
nand U3803 (N_3803,N_1716,N_2477);
and U3804 (N_3804,N_2349,N_2127);
nor U3805 (N_3805,N_2367,N_1599);
nor U3806 (N_3806,N_2168,N_2117);
and U3807 (N_3807,N_1977,N_1533);
and U3808 (N_3808,N_1708,N_1571);
or U3809 (N_3809,N_2157,N_2665);
or U3810 (N_3810,N_2111,N_2466);
and U3811 (N_3811,N_2980,N_2454);
and U3812 (N_3812,N_1677,N_1582);
or U3813 (N_3813,N_1770,N_2415);
or U3814 (N_3814,N_2197,N_2642);
or U3815 (N_3815,N_2360,N_1640);
nor U3816 (N_3816,N_1599,N_1719);
and U3817 (N_3817,N_2708,N_2061);
nor U3818 (N_3818,N_2528,N_2027);
or U3819 (N_3819,N_1532,N_2450);
nand U3820 (N_3820,N_2597,N_2456);
or U3821 (N_3821,N_2972,N_2905);
and U3822 (N_3822,N_2062,N_2150);
nand U3823 (N_3823,N_1566,N_1548);
nand U3824 (N_3824,N_2252,N_2623);
and U3825 (N_3825,N_2538,N_2475);
nand U3826 (N_3826,N_2811,N_2789);
nor U3827 (N_3827,N_1781,N_2189);
nor U3828 (N_3828,N_2892,N_2662);
nor U3829 (N_3829,N_2741,N_1529);
nand U3830 (N_3830,N_1783,N_2904);
nor U3831 (N_3831,N_1833,N_1685);
or U3832 (N_3832,N_1945,N_1755);
and U3833 (N_3833,N_2582,N_2710);
and U3834 (N_3834,N_2432,N_2014);
or U3835 (N_3835,N_2685,N_1902);
and U3836 (N_3836,N_2837,N_1889);
or U3837 (N_3837,N_2333,N_2366);
and U3838 (N_3838,N_2500,N_1785);
nand U3839 (N_3839,N_1717,N_1530);
nor U3840 (N_3840,N_2020,N_1792);
nor U3841 (N_3841,N_2155,N_2987);
or U3842 (N_3842,N_2462,N_2541);
xor U3843 (N_3843,N_1518,N_2273);
and U3844 (N_3844,N_2472,N_2187);
and U3845 (N_3845,N_2535,N_2663);
nor U3846 (N_3846,N_2603,N_2719);
nand U3847 (N_3847,N_1732,N_2081);
and U3848 (N_3848,N_2772,N_2729);
nor U3849 (N_3849,N_1764,N_2191);
and U3850 (N_3850,N_1692,N_2180);
and U3851 (N_3851,N_1893,N_2552);
nand U3852 (N_3852,N_1840,N_2551);
or U3853 (N_3853,N_2649,N_2827);
nor U3854 (N_3854,N_2087,N_2886);
or U3855 (N_3855,N_2505,N_2415);
or U3856 (N_3856,N_1646,N_2221);
nand U3857 (N_3857,N_2359,N_2042);
nor U3858 (N_3858,N_2436,N_1541);
and U3859 (N_3859,N_2648,N_1673);
and U3860 (N_3860,N_2832,N_2401);
and U3861 (N_3861,N_2921,N_1737);
nor U3862 (N_3862,N_2025,N_1993);
or U3863 (N_3863,N_2550,N_2174);
and U3864 (N_3864,N_2825,N_2018);
nor U3865 (N_3865,N_2728,N_2427);
nor U3866 (N_3866,N_1608,N_2834);
nor U3867 (N_3867,N_2815,N_2619);
and U3868 (N_3868,N_2444,N_2689);
nor U3869 (N_3869,N_2345,N_2821);
xor U3870 (N_3870,N_1927,N_2286);
nand U3871 (N_3871,N_2273,N_2839);
or U3872 (N_3872,N_2163,N_1681);
and U3873 (N_3873,N_2523,N_1743);
nor U3874 (N_3874,N_2485,N_2354);
and U3875 (N_3875,N_2926,N_2824);
nor U3876 (N_3876,N_1883,N_1748);
nor U3877 (N_3877,N_1985,N_1551);
nor U3878 (N_3878,N_1810,N_2954);
and U3879 (N_3879,N_1522,N_2816);
and U3880 (N_3880,N_2784,N_2170);
nand U3881 (N_3881,N_2463,N_2519);
or U3882 (N_3882,N_2187,N_2206);
nor U3883 (N_3883,N_2333,N_2152);
nand U3884 (N_3884,N_2315,N_2775);
or U3885 (N_3885,N_2960,N_2710);
nand U3886 (N_3886,N_2552,N_1544);
nand U3887 (N_3887,N_2929,N_2444);
xnor U3888 (N_3888,N_2674,N_1697);
nor U3889 (N_3889,N_2577,N_2715);
nor U3890 (N_3890,N_1699,N_2694);
nor U3891 (N_3891,N_2547,N_1536);
nand U3892 (N_3892,N_2867,N_1759);
nand U3893 (N_3893,N_2306,N_2073);
nand U3894 (N_3894,N_2997,N_2419);
nor U3895 (N_3895,N_2109,N_2783);
nand U3896 (N_3896,N_2485,N_1964);
nor U3897 (N_3897,N_2178,N_2460);
and U3898 (N_3898,N_1953,N_2061);
nand U3899 (N_3899,N_2563,N_2600);
nand U3900 (N_3900,N_1613,N_2193);
and U3901 (N_3901,N_2452,N_2801);
or U3902 (N_3902,N_2588,N_1839);
or U3903 (N_3903,N_1747,N_1545);
and U3904 (N_3904,N_2005,N_2685);
nor U3905 (N_3905,N_2169,N_2702);
and U3906 (N_3906,N_2124,N_2030);
nand U3907 (N_3907,N_2964,N_1941);
and U3908 (N_3908,N_1712,N_2135);
nor U3909 (N_3909,N_2625,N_2384);
or U3910 (N_3910,N_2470,N_2663);
nor U3911 (N_3911,N_2780,N_2345);
nand U3912 (N_3912,N_2792,N_1812);
or U3913 (N_3913,N_2535,N_1715);
nor U3914 (N_3914,N_2740,N_1516);
and U3915 (N_3915,N_2822,N_2356);
and U3916 (N_3916,N_2192,N_1934);
or U3917 (N_3917,N_2490,N_1804);
and U3918 (N_3918,N_2948,N_1916);
or U3919 (N_3919,N_2746,N_2470);
xor U3920 (N_3920,N_1505,N_2009);
or U3921 (N_3921,N_2205,N_1645);
or U3922 (N_3922,N_2213,N_1847);
or U3923 (N_3923,N_2181,N_2749);
or U3924 (N_3924,N_2409,N_2117);
nand U3925 (N_3925,N_2926,N_2058);
nand U3926 (N_3926,N_2097,N_1969);
or U3927 (N_3927,N_1579,N_2546);
and U3928 (N_3928,N_1711,N_1644);
nor U3929 (N_3929,N_2677,N_2829);
nor U3930 (N_3930,N_1955,N_1500);
nor U3931 (N_3931,N_2099,N_2518);
and U3932 (N_3932,N_2086,N_1767);
or U3933 (N_3933,N_2141,N_2083);
nor U3934 (N_3934,N_2627,N_2282);
and U3935 (N_3935,N_1582,N_2931);
nor U3936 (N_3936,N_2129,N_2540);
or U3937 (N_3937,N_1953,N_1722);
nor U3938 (N_3938,N_2343,N_2328);
nor U3939 (N_3939,N_2794,N_2759);
nand U3940 (N_3940,N_2312,N_2258);
nand U3941 (N_3941,N_1868,N_2650);
nor U3942 (N_3942,N_2962,N_2646);
and U3943 (N_3943,N_2480,N_1945);
and U3944 (N_3944,N_2822,N_2681);
nor U3945 (N_3945,N_1626,N_2797);
nor U3946 (N_3946,N_2316,N_2080);
nand U3947 (N_3947,N_1654,N_1686);
nand U3948 (N_3948,N_2947,N_2512);
and U3949 (N_3949,N_2988,N_1731);
and U3950 (N_3950,N_2060,N_2259);
nor U3951 (N_3951,N_1993,N_1753);
nand U3952 (N_3952,N_2659,N_2534);
and U3953 (N_3953,N_2571,N_1754);
nand U3954 (N_3954,N_2343,N_2348);
or U3955 (N_3955,N_2796,N_2119);
or U3956 (N_3956,N_2361,N_1523);
and U3957 (N_3957,N_2867,N_1800);
nand U3958 (N_3958,N_1599,N_1543);
or U3959 (N_3959,N_2447,N_1547);
or U3960 (N_3960,N_1589,N_2469);
xor U3961 (N_3961,N_2009,N_2603);
nand U3962 (N_3962,N_2811,N_1852);
and U3963 (N_3963,N_2337,N_2081);
or U3964 (N_3964,N_2897,N_2893);
nor U3965 (N_3965,N_2567,N_2141);
nor U3966 (N_3966,N_2269,N_2144);
and U3967 (N_3967,N_1943,N_1990);
nand U3968 (N_3968,N_2332,N_2593);
and U3969 (N_3969,N_2270,N_1984);
nand U3970 (N_3970,N_1763,N_2464);
xnor U3971 (N_3971,N_2272,N_2285);
nand U3972 (N_3972,N_1757,N_2714);
nor U3973 (N_3973,N_2403,N_2895);
and U3974 (N_3974,N_1994,N_2406);
and U3975 (N_3975,N_2852,N_1941);
nand U3976 (N_3976,N_2369,N_2608);
and U3977 (N_3977,N_1860,N_2657);
or U3978 (N_3978,N_2130,N_2980);
nand U3979 (N_3979,N_1835,N_2579);
nand U3980 (N_3980,N_2242,N_2467);
nor U3981 (N_3981,N_1733,N_1892);
and U3982 (N_3982,N_2362,N_2905);
nor U3983 (N_3983,N_2869,N_1896);
or U3984 (N_3984,N_2785,N_1762);
and U3985 (N_3985,N_2682,N_2231);
nand U3986 (N_3986,N_1962,N_1792);
or U3987 (N_3987,N_1592,N_2921);
and U3988 (N_3988,N_2229,N_2854);
or U3989 (N_3989,N_2778,N_1521);
nand U3990 (N_3990,N_1744,N_1610);
and U3991 (N_3991,N_1901,N_2186);
nand U3992 (N_3992,N_2350,N_2072);
or U3993 (N_3993,N_2878,N_2839);
and U3994 (N_3994,N_1790,N_2690);
and U3995 (N_3995,N_2364,N_1777);
nand U3996 (N_3996,N_2328,N_2248);
and U3997 (N_3997,N_1540,N_1779);
nand U3998 (N_3998,N_1663,N_2131);
and U3999 (N_3999,N_1569,N_2078);
or U4000 (N_4000,N_2423,N_1531);
nand U4001 (N_4001,N_2624,N_1701);
nand U4002 (N_4002,N_1856,N_2928);
nor U4003 (N_4003,N_2050,N_1747);
nor U4004 (N_4004,N_2612,N_2783);
or U4005 (N_4005,N_2104,N_2093);
nor U4006 (N_4006,N_1929,N_2887);
nand U4007 (N_4007,N_1596,N_1508);
nor U4008 (N_4008,N_2399,N_2926);
nand U4009 (N_4009,N_2819,N_2294);
and U4010 (N_4010,N_2285,N_2326);
nand U4011 (N_4011,N_2125,N_1963);
nand U4012 (N_4012,N_2105,N_1723);
or U4013 (N_4013,N_2648,N_2096);
nand U4014 (N_4014,N_2707,N_2469);
nand U4015 (N_4015,N_2417,N_2171);
or U4016 (N_4016,N_2840,N_1707);
and U4017 (N_4017,N_2260,N_2138);
and U4018 (N_4018,N_1942,N_2470);
xnor U4019 (N_4019,N_2345,N_2384);
or U4020 (N_4020,N_1695,N_1918);
nand U4021 (N_4021,N_2836,N_1872);
or U4022 (N_4022,N_1689,N_1772);
nor U4023 (N_4023,N_1637,N_2574);
or U4024 (N_4024,N_1630,N_1695);
and U4025 (N_4025,N_2072,N_1953);
nand U4026 (N_4026,N_2660,N_2186);
nor U4027 (N_4027,N_1780,N_2487);
or U4028 (N_4028,N_2024,N_1535);
or U4029 (N_4029,N_1696,N_2189);
and U4030 (N_4030,N_2823,N_1669);
and U4031 (N_4031,N_1876,N_2833);
and U4032 (N_4032,N_2750,N_2826);
and U4033 (N_4033,N_2855,N_2914);
xnor U4034 (N_4034,N_2430,N_1648);
and U4035 (N_4035,N_2034,N_2961);
and U4036 (N_4036,N_2944,N_2565);
nor U4037 (N_4037,N_1924,N_1713);
or U4038 (N_4038,N_2342,N_2894);
nor U4039 (N_4039,N_1641,N_2157);
nand U4040 (N_4040,N_2676,N_1793);
nand U4041 (N_4041,N_2018,N_2820);
nand U4042 (N_4042,N_1804,N_2025);
or U4043 (N_4043,N_2300,N_1723);
and U4044 (N_4044,N_2915,N_2612);
nand U4045 (N_4045,N_2596,N_2960);
and U4046 (N_4046,N_2900,N_2552);
or U4047 (N_4047,N_2287,N_1917);
and U4048 (N_4048,N_1571,N_2905);
or U4049 (N_4049,N_1941,N_2759);
or U4050 (N_4050,N_1750,N_2266);
and U4051 (N_4051,N_1711,N_1892);
nand U4052 (N_4052,N_1886,N_2794);
or U4053 (N_4053,N_2981,N_1619);
nand U4054 (N_4054,N_1626,N_2482);
and U4055 (N_4055,N_2970,N_1995);
nor U4056 (N_4056,N_2241,N_2399);
or U4057 (N_4057,N_1579,N_2340);
nor U4058 (N_4058,N_2602,N_2772);
or U4059 (N_4059,N_2191,N_2811);
and U4060 (N_4060,N_2426,N_2820);
nor U4061 (N_4061,N_2291,N_2691);
and U4062 (N_4062,N_2431,N_2913);
and U4063 (N_4063,N_1779,N_1979);
or U4064 (N_4064,N_2660,N_1784);
nand U4065 (N_4065,N_2768,N_2248);
or U4066 (N_4066,N_2465,N_2461);
nand U4067 (N_4067,N_2002,N_2578);
or U4068 (N_4068,N_2520,N_2350);
or U4069 (N_4069,N_1602,N_1531);
nor U4070 (N_4070,N_2848,N_2343);
and U4071 (N_4071,N_1600,N_2156);
xor U4072 (N_4072,N_1969,N_1755);
or U4073 (N_4073,N_1889,N_1792);
xnor U4074 (N_4074,N_2797,N_2229);
or U4075 (N_4075,N_2794,N_2946);
or U4076 (N_4076,N_2202,N_2041);
nor U4077 (N_4077,N_1541,N_2528);
nand U4078 (N_4078,N_2126,N_2712);
and U4079 (N_4079,N_1518,N_1870);
nand U4080 (N_4080,N_2967,N_1810);
or U4081 (N_4081,N_2892,N_2128);
nor U4082 (N_4082,N_1708,N_1848);
or U4083 (N_4083,N_1548,N_2314);
xor U4084 (N_4084,N_2916,N_1666);
and U4085 (N_4085,N_1780,N_1867);
or U4086 (N_4086,N_1519,N_2494);
and U4087 (N_4087,N_1678,N_2649);
xor U4088 (N_4088,N_2891,N_2718);
nand U4089 (N_4089,N_1689,N_2704);
nor U4090 (N_4090,N_1530,N_2229);
nor U4091 (N_4091,N_2473,N_1918);
and U4092 (N_4092,N_2134,N_2065);
nand U4093 (N_4093,N_1527,N_2191);
nor U4094 (N_4094,N_1721,N_2764);
nor U4095 (N_4095,N_2805,N_2357);
or U4096 (N_4096,N_2256,N_2604);
or U4097 (N_4097,N_1560,N_2671);
or U4098 (N_4098,N_1787,N_2740);
and U4099 (N_4099,N_1863,N_1562);
or U4100 (N_4100,N_1609,N_2937);
nor U4101 (N_4101,N_2612,N_1635);
xnor U4102 (N_4102,N_2661,N_2532);
or U4103 (N_4103,N_1967,N_1642);
nor U4104 (N_4104,N_1812,N_2970);
and U4105 (N_4105,N_1861,N_2660);
nor U4106 (N_4106,N_2244,N_2990);
nand U4107 (N_4107,N_2477,N_2226);
and U4108 (N_4108,N_2450,N_1848);
nor U4109 (N_4109,N_2132,N_1780);
and U4110 (N_4110,N_2063,N_2123);
or U4111 (N_4111,N_2687,N_2241);
nor U4112 (N_4112,N_2558,N_2473);
nand U4113 (N_4113,N_1506,N_1614);
nand U4114 (N_4114,N_2538,N_2307);
and U4115 (N_4115,N_1895,N_1501);
or U4116 (N_4116,N_2706,N_2822);
or U4117 (N_4117,N_2817,N_2328);
or U4118 (N_4118,N_1952,N_2385);
or U4119 (N_4119,N_1740,N_2526);
or U4120 (N_4120,N_2910,N_2188);
and U4121 (N_4121,N_1945,N_2994);
nor U4122 (N_4122,N_1687,N_2903);
and U4123 (N_4123,N_1857,N_2061);
nor U4124 (N_4124,N_2804,N_2944);
nand U4125 (N_4125,N_2546,N_2215);
nand U4126 (N_4126,N_2043,N_2997);
nand U4127 (N_4127,N_2053,N_2606);
or U4128 (N_4128,N_2649,N_2217);
or U4129 (N_4129,N_2518,N_2823);
nor U4130 (N_4130,N_2608,N_2641);
nor U4131 (N_4131,N_2637,N_2218);
or U4132 (N_4132,N_1927,N_1826);
nor U4133 (N_4133,N_2239,N_2829);
xor U4134 (N_4134,N_1552,N_2702);
nand U4135 (N_4135,N_1631,N_1854);
nor U4136 (N_4136,N_2069,N_2089);
nand U4137 (N_4137,N_2813,N_1799);
nor U4138 (N_4138,N_2692,N_2149);
nand U4139 (N_4139,N_2180,N_2886);
nor U4140 (N_4140,N_1509,N_2992);
nand U4141 (N_4141,N_2764,N_2991);
xor U4142 (N_4142,N_1514,N_2964);
and U4143 (N_4143,N_2311,N_2535);
or U4144 (N_4144,N_2213,N_2847);
nor U4145 (N_4145,N_2242,N_1530);
nand U4146 (N_4146,N_2890,N_1899);
or U4147 (N_4147,N_2596,N_2638);
nor U4148 (N_4148,N_2518,N_1801);
or U4149 (N_4149,N_2637,N_1743);
nand U4150 (N_4150,N_2633,N_2535);
or U4151 (N_4151,N_2209,N_1825);
and U4152 (N_4152,N_2512,N_2180);
or U4153 (N_4153,N_2933,N_2461);
nand U4154 (N_4154,N_2267,N_2630);
and U4155 (N_4155,N_1516,N_2469);
or U4156 (N_4156,N_1717,N_2666);
or U4157 (N_4157,N_2201,N_1744);
or U4158 (N_4158,N_1645,N_1632);
and U4159 (N_4159,N_2408,N_1987);
or U4160 (N_4160,N_2123,N_1882);
nor U4161 (N_4161,N_2990,N_1545);
and U4162 (N_4162,N_2646,N_1519);
nor U4163 (N_4163,N_2018,N_2318);
or U4164 (N_4164,N_2119,N_2687);
or U4165 (N_4165,N_2377,N_2980);
and U4166 (N_4166,N_2970,N_1525);
xor U4167 (N_4167,N_2442,N_2703);
nor U4168 (N_4168,N_1647,N_1814);
and U4169 (N_4169,N_2868,N_2032);
and U4170 (N_4170,N_2507,N_1909);
nor U4171 (N_4171,N_1924,N_1950);
or U4172 (N_4172,N_1711,N_2370);
nand U4173 (N_4173,N_2337,N_2783);
xor U4174 (N_4174,N_1535,N_2626);
or U4175 (N_4175,N_2284,N_1666);
nor U4176 (N_4176,N_2458,N_2105);
nor U4177 (N_4177,N_1676,N_2326);
nor U4178 (N_4178,N_2411,N_2419);
and U4179 (N_4179,N_2184,N_1873);
nand U4180 (N_4180,N_1857,N_2103);
and U4181 (N_4181,N_1501,N_2164);
and U4182 (N_4182,N_1709,N_2975);
nand U4183 (N_4183,N_2883,N_2426);
nand U4184 (N_4184,N_2966,N_2679);
nor U4185 (N_4185,N_2565,N_2553);
nor U4186 (N_4186,N_2051,N_2710);
nand U4187 (N_4187,N_2907,N_2729);
and U4188 (N_4188,N_1941,N_2630);
or U4189 (N_4189,N_2538,N_2873);
and U4190 (N_4190,N_2073,N_2681);
nor U4191 (N_4191,N_1699,N_2512);
nor U4192 (N_4192,N_1714,N_2632);
nand U4193 (N_4193,N_2306,N_2782);
nor U4194 (N_4194,N_2609,N_2533);
nand U4195 (N_4195,N_2153,N_2123);
and U4196 (N_4196,N_2197,N_2631);
nand U4197 (N_4197,N_2010,N_2615);
and U4198 (N_4198,N_1886,N_1597);
and U4199 (N_4199,N_2497,N_2189);
nor U4200 (N_4200,N_2600,N_2805);
nor U4201 (N_4201,N_2289,N_2185);
or U4202 (N_4202,N_1511,N_2006);
or U4203 (N_4203,N_1831,N_2129);
and U4204 (N_4204,N_2543,N_2510);
nand U4205 (N_4205,N_1646,N_2295);
nor U4206 (N_4206,N_2289,N_2040);
and U4207 (N_4207,N_2314,N_2903);
and U4208 (N_4208,N_2294,N_2912);
and U4209 (N_4209,N_2863,N_2416);
or U4210 (N_4210,N_2958,N_2868);
nand U4211 (N_4211,N_1685,N_1694);
and U4212 (N_4212,N_2111,N_2093);
nand U4213 (N_4213,N_2369,N_2870);
nor U4214 (N_4214,N_2090,N_2721);
nand U4215 (N_4215,N_2047,N_1637);
nor U4216 (N_4216,N_2852,N_2478);
nor U4217 (N_4217,N_1697,N_2143);
nand U4218 (N_4218,N_2908,N_2169);
nor U4219 (N_4219,N_2665,N_2976);
nand U4220 (N_4220,N_1804,N_2976);
nor U4221 (N_4221,N_2686,N_2771);
and U4222 (N_4222,N_2364,N_2540);
nand U4223 (N_4223,N_2017,N_2774);
nor U4224 (N_4224,N_2047,N_2439);
nand U4225 (N_4225,N_2861,N_2761);
or U4226 (N_4226,N_2175,N_2341);
or U4227 (N_4227,N_2812,N_2359);
nor U4228 (N_4228,N_2627,N_2762);
nand U4229 (N_4229,N_1790,N_2563);
nand U4230 (N_4230,N_1790,N_2541);
nor U4231 (N_4231,N_2400,N_1771);
nand U4232 (N_4232,N_2790,N_2212);
or U4233 (N_4233,N_2470,N_2370);
and U4234 (N_4234,N_2971,N_2337);
nor U4235 (N_4235,N_2442,N_2387);
nand U4236 (N_4236,N_2283,N_2898);
or U4237 (N_4237,N_2573,N_2966);
and U4238 (N_4238,N_2156,N_2447);
nor U4239 (N_4239,N_2522,N_2605);
nand U4240 (N_4240,N_2768,N_2763);
or U4241 (N_4241,N_2644,N_1977);
nand U4242 (N_4242,N_2652,N_2847);
nor U4243 (N_4243,N_2326,N_1552);
or U4244 (N_4244,N_1525,N_2857);
nand U4245 (N_4245,N_2910,N_1594);
and U4246 (N_4246,N_2663,N_1642);
xnor U4247 (N_4247,N_2658,N_2661);
xnor U4248 (N_4248,N_1701,N_2478);
xor U4249 (N_4249,N_1780,N_2981);
and U4250 (N_4250,N_2139,N_2351);
and U4251 (N_4251,N_2241,N_2576);
and U4252 (N_4252,N_1553,N_1967);
and U4253 (N_4253,N_1726,N_2672);
nor U4254 (N_4254,N_2021,N_1945);
nand U4255 (N_4255,N_2925,N_2550);
or U4256 (N_4256,N_1910,N_1987);
nor U4257 (N_4257,N_2115,N_1833);
nor U4258 (N_4258,N_1579,N_2142);
or U4259 (N_4259,N_1614,N_2779);
nor U4260 (N_4260,N_1590,N_1515);
and U4261 (N_4261,N_2121,N_2664);
or U4262 (N_4262,N_2841,N_2891);
nor U4263 (N_4263,N_1946,N_2504);
and U4264 (N_4264,N_1786,N_2712);
nor U4265 (N_4265,N_2954,N_2224);
and U4266 (N_4266,N_1921,N_2223);
or U4267 (N_4267,N_1690,N_1908);
nor U4268 (N_4268,N_1948,N_2457);
or U4269 (N_4269,N_1836,N_1905);
or U4270 (N_4270,N_1670,N_2116);
nor U4271 (N_4271,N_1621,N_1795);
xor U4272 (N_4272,N_2756,N_2327);
or U4273 (N_4273,N_1725,N_2897);
nand U4274 (N_4274,N_1615,N_1544);
and U4275 (N_4275,N_1621,N_2348);
or U4276 (N_4276,N_2398,N_2893);
nor U4277 (N_4277,N_2349,N_1833);
nand U4278 (N_4278,N_2899,N_1815);
and U4279 (N_4279,N_2058,N_2347);
or U4280 (N_4280,N_2228,N_2158);
and U4281 (N_4281,N_2185,N_1624);
and U4282 (N_4282,N_2483,N_1631);
and U4283 (N_4283,N_2189,N_2547);
nand U4284 (N_4284,N_2591,N_1916);
or U4285 (N_4285,N_2591,N_2755);
or U4286 (N_4286,N_1819,N_2335);
nor U4287 (N_4287,N_2474,N_1779);
nor U4288 (N_4288,N_2695,N_1631);
nor U4289 (N_4289,N_2828,N_2386);
or U4290 (N_4290,N_1502,N_1879);
and U4291 (N_4291,N_1505,N_2336);
nand U4292 (N_4292,N_2275,N_1817);
nand U4293 (N_4293,N_2693,N_2065);
and U4294 (N_4294,N_2394,N_2996);
or U4295 (N_4295,N_2882,N_2914);
nor U4296 (N_4296,N_2778,N_2812);
nand U4297 (N_4297,N_1809,N_2440);
or U4298 (N_4298,N_1769,N_1563);
or U4299 (N_4299,N_1918,N_2440);
xor U4300 (N_4300,N_1991,N_2612);
nor U4301 (N_4301,N_1885,N_2719);
nand U4302 (N_4302,N_1518,N_1939);
and U4303 (N_4303,N_2123,N_2072);
nand U4304 (N_4304,N_2103,N_2027);
nor U4305 (N_4305,N_2378,N_2855);
or U4306 (N_4306,N_1630,N_2283);
nor U4307 (N_4307,N_1742,N_2693);
or U4308 (N_4308,N_1872,N_1750);
xor U4309 (N_4309,N_2081,N_2868);
and U4310 (N_4310,N_2570,N_2875);
nand U4311 (N_4311,N_2411,N_1558);
or U4312 (N_4312,N_1790,N_2776);
nand U4313 (N_4313,N_1667,N_2134);
or U4314 (N_4314,N_1922,N_2986);
nand U4315 (N_4315,N_2999,N_2780);
nand U4316 (N_4316,N_1522,N_2065);
and U4317 (N_4317,N_2315,N_2482);
nand U4318 (N_4318,N_1582,N_2383);
nor U4319 (N_4319,N_1634,N_2625);
nor U4320 (N_4320,N_2153,N_1591);
or U4321 (N_4321,N_1862,N_1653);
nand U4322 (N_4322,N_1640,N_1888);
and U4323 (N_4323,N_1667,N_2594);
nand U4324 (N_4324,N_2055,N_2158);
and U4325 (N_4325,N_2861,N_1895);
and U4326 (N_4326,N_1592,N_1830);
nand U4327 (N_4327,N_1964,N_2205);
nand U4328 (N_4328,N_2781,N_2312);
or U4329 (N_4329,N_2088,N_2022);
nor U4330 (N_4330,N_2727,N_2202);
and U4331 (N_4331,N_1707,N_1972);
nand U4332 (N_4332,N_2514,N_2485);
or U4333 (N_4333,N_1880,N_2794);
or U4334 (N_4334,N_2143,N_2305);
and U4335 (N_4335,N_2326,N_2242);
nand U4336 (N_4336,N_2460,N_2646);
nor U4337 (N_4337,N_2812,N_1799);
nand U4338 (N_4338,N_2431,N_2115);
nand U4339 (N_4339,N_2547,N_2709);
or U4340 (N_4340,N_2279,N_1713);
nand U4341 (N_4341,N_1714,N_2655);
nor U4342 (N_4342,N_2899,N_1716);
nor U4343 (N_4343,N_2481,N_2479);
nand U4344 (N_4344,N_2923,N_2431);
and U4345 (N_4345,N_1771,N_2916);
and U4346 (N_4346,N_1984,N_1527);
nand U4347 (N_4347,N_2495,N_2386);
and U4348 (N_4348,N_1646,N_1861);
and U4349 (N_4349,N_2086,N_1771);
nand U4350 (N_4350,N_2085,N_2060);
or U4351 (N_4351,N_2219,N_2323);
or U4352 (N_4352,N_2438,N_2123);
nand U4353 (N_4353,N_1641,N_2722);
or U4354 (N_4354,N_1616,N_1709);
nand U4355 (N_4355,N_2540,N_2969);
and U4356 (N_4356,N_2227,N_2059);
nor U4357 (N_4357,N_2914,N_2936);
and U4358 (N_4358,N_2319,N_2961);
nor U4359 (N_4359,N_1988,N_2846);
and U4360 (N_4360,N_1841,N_1737);
or U4361 (N_4361,N_2063,N_2226);
or U4362 (N_4362,N_2998,N_1904);
nor U4363 (N_4363,N_1592,N_2831);
and U4364 (N_4364,N_2512,N_2428);
and U4365 (N_4365,N_2777,N_2041);
nand U4366 (N_4366,N_2788,N_2357);
or U4367 (N_4367,N_1982,N_2370);
or U4368 (N_4368,N_2776,N_2387);
or U4369 (N_4369,N_2927,N_2407);
or U4370 (N_4370,N_2074,N_2939);
nand U4371 (N_4371,N_1995,N_2513);
nand U4372 (N_4372,N_2851,N_1850);
nand U4373 (N_4373,N_2408,N_2686);
and U4374 (N_4374,N_1799,N_1779);
and U4375 (N_4375,N_2046,N_1689);
nand U4376 (N_4376,N_2664,N_2071);
or U4377 (N_4377,N_1785,N_1841);
and U4378 (N_4378,N_2639,N_1840);
nand U4379 (N_4379,N_2605,N_2240);
nor U4380 (N_4380,N_2774,N_2985);
or U4381 (N_4381,N_1712,N_2778);
or U4382 (N_4382,N_1776,N_1924);
or U4383 (N_4383,N_2821,N_2660);
and U4384 (N_4384,N_1897,N_2045);
nor U4385 (N_4385,N_1917,N_2606);
nand U4386 (N_4386,N_1519,N_1822);
nand U4387 (N_4387,N_1971,N_1864);
xnor U4388 (N_4388,N_2855,N_2140);
nor U4389 (N_4389,N_2286,N_2612);
or U4390 (N_4390,N_1584,N_2204);
nor U4391 (N_4391,N_2615,N_2839);
and U4392 (N_4392,N_2851,N_1638);
nand U4393 (N_4393,N_2529,N_1670);
and U4394 (N_4394,N_2607,N_2976);
xnor U4395 (N_4395,N_2529,N_2332);
and U4396 (N_4396,N_1954,N_2816);
or U4397 (N_4397,N_1917,N_1806);
nor U4398 (N_4398,N_2059,N_1732);
xor U4399 (N_4399,N_2688,N_2700);
nand U4400 (N_4400,N_2494,N_1691);
and U4401 (N_4401,N_2555,N_1616);
or U4402 (N_4402,N_2699,N_1609);
and U4403 (N_4403,N_2131,N_2557);
xnor U4404 (N_4404,N_2944,N_2186);
nor U4405 (N_4405,N_2470,N_2640);
nor U4406 (N_4406,N_2769,N_2592);
or U4407 (N_4407,N_1923,N_2875);
nand U4408 (N_4408,N_2432,N_2499);
nor U4409 (N_4409,N_1627,N_2151);
and U4410 (N_4410,N_2210,N_2209);
nor U4411 (N_4411,N_2577,N_2355);
nand U4412 (N_4412,N_2190,N_2110);
nand U4413 (N_4413,N_2304,N_2384);
nor U4414 (N_4414,N_2116,N_1657);
nor U4415 (N_4415,N_1843,N_1824);
nor U4416 (N_4416,N_2885,N_1647);
nand U4417 (N_4417,N_1913,N_2049);
and U4418 (N_4418,N_2006,N_1502);
nor U4419 (N_4419,N_2906,N_1835);
or U4420 (N_4420,N_2954,N_1844);
and U4421 (N_4421,N_2593,N_1603);
and U4422 (N_4422,N_2924,N_2912);
nand U4423 (N_4423,N_2170,N_2819);
nor U4424 (N_4424,N_2883,N_2030);
nand U4425 (N_4425,N_2911,N_1714);
or U4426 (N_4426,N_2639,N_2815);
nand U4427 (N_4427,N_1570,N_2817);
nand U4428 (N_4428,N_2207,N_1665);
and U4429 (N_4429,N_2220,N_2443);
or U4430 (N_4430,N_1792,N_2493);
nor U4431 (N_4431,N_1661,N_1809);
and U4432 (N_4432,N_2001,N_1611);
nand U4433 (N_4433,N_2118,N_2042);
or U4434 (N_4434,N_2569,N_2989);
nor U4435 (N_4435,N_2723,N_1908);
nor U4436 (N_4436,N_2593,N_2674);
or U4437 (N_4437,N_2636,N_1629);
or U4438 (N_4438,N_2387,N_2711);
nand U4439 (N_4439,N_2604,N_1532);
xor U4440 (N_4440,N_2088,N_2027);
and U4441 (N_4441,N_2844,N_2434);
and U4442 (N_4442,N_2667,N_2015);
or U4443 (N_4443,N_2490,N_2781);
or U4444 (N_4444,N_1777,N_1745);
or U4445 (N_4445,N_1737,N_1947);
nor U4446 (N_4446,N_1931,N_1786);
and U4447 (N_4447,N_2792,N_2026);
and U4448 (N_4448,N_1986,N_2196);
and U4449 (N_4449,N_1650,N_2499);
and U4450 (N_4450,N_2404,N_1676);
and U4451 (N_4451,N_2696,N_2146);
nor U4452 (N_4452,N_1823,N_2813);
nor U4453 (N_4453,N_1609,N_2191);
or U4454 (N_4454,N_1762,N_2958);
nor U4455 (N_4455,N_2598,N_2649);
nor U4456 (N_4456,N_1595,N_1794);
or U4457 (N_4457,N_2467,N_2259);
or U4458 (N_4458,N_2182,N_2218);
nor U4459 (N_4459,N_1631,N_2242);
and U4460 (N_4460,N_2783,N_2098);
nand U4461 (N_4461,N_2770,N_2813);
xnor U4462 (N_4462,N_2141,N_1813);
xnor U4463 (N_4463,N_2568,N_2516);
and U4464 (N_4464,N_2437,N_2203);
nor U4465 (N_4465,N_2826,N_2100);
nand U4466 (N_4466,N_2531,N_2343);
or U4467 (N_4467,N_1634,N_2229);
or U4468 (N_4468,N_1692,N_1675);
xor U4469 (N_4469,N_1800,N_1617);
and U4470 (N_4470,N_1750,N_2617);
nor U4471 (N_4471,N_1696,N_2144);
nand U4472 (N_4472,N_2384,N_1640);
and U4473 (N_4473,N_1642,N_1684);
and U4474 (N_4474,N_2095,N_2479);
or U4475 (N_4475,N_1581,N_2791);
and U4476 (N_4476,N_2869,N_1727);
nand U4477 (N_4477,N_2145,N_2044);
nor U4478 (N_4478,N_2271,N_1619);
nand U4479 (N_4479,N_2390,N_1518);
and U4480 (N_4480,N_2986,N_1976);
and U4481 (N_4481,N_2932,N_2453);
nor U4482 (N_4482,N_2136,N_1610);
and U4483 (N_4483,N_2649,N_2967);
and U4484 (N_4484,N_2246,N_2309);
and U4485 (N_4485,N_2875,N_2973);
xor U4486 (N_4486,N_2401,N_2087);
nand U4487 (N_4487,N_1835,N_2180);
nor U4488 (N_4488,N_2317,N_2377);
and U4489 (N_4489,N_2710,N_1921);
and U4490 (N_4490,N_2505,N_2393);
nand U4491 (N_4491,N_2014,N_1716);
and U4492 (N_4492,N_1521,N_2117);
and U4493 (N_4493,N_1635,N_2208);
and U4494 (N_4494,N_2231,N_2790);
and U4495 (N_4495,N_2679,N_1902);
nor U4496 (N_4496,N_2659,N_1895);
and U4497 (N_4497,N_2495,N_2951);
nand U4498 (N_4498,N_2014,N_2947);
or U4499 (N_4499,N_2764,N_2624);
nor U4500 (N_4500,N_3161,N_4115);
nand U4501 (N_4501,N_4467,N_3292);
or U4502 (N_4502,N_4003,N_3203);
or U4503 (N_4503,N_3676,N_3268);
or U4504 (N_4504,N_3307,N_3218);
nand U4505 (N_4505,N_3394,N_4478);
nand U4506 (N_4506,N_4389,N_3931);
nand U4507 (N_4507,N_4350,N_3908);
and U4508 (N_4508,N_4498,N_3088);
nand U4509 (N_4509,N_3255,N_3191);
or U4510 (N_4510,N_4370,N_4172);
or U4511 (N_4511,N_3983,N_4394);
nand U4512 (N_4512,N_3787,N_3456);
nor U4513 (N_4513,N_4265,N_4450);
or U4514 (N_4514,N_3228,N_3419);
and U4515 (N_4515,N_3576,N_4220);
nor U4516 (N_4516,N_4169,N_3339);
nand U4517 (N_4517,N_4249,N_3310);
and U4518 (N_4518,N_4330,N_3572);
nor U4519 (N_4519,N_3170,N_3683);
xor U4520 (N_4520,N_4002,N_3362);
nor U4521 (N_4521,N_3723,N_4023);
nand U4522 (N_4522,N_3820,N_4399);
and U4523 (N_4523,N_3167,N_4475);
nor U4524 (N_4524,N_3123,N_4014);
nor U4525 (N_4525,N_3960,N_3017);
xnor U4526 (N_4526,N_3797,N_3776);
or U4527 (N_4527,N_3597,N_3485);
or U4528 (N_4528,N_3948,N_3095);
and U4529 (N_4529,N_3637,N_3254);
and U4530 (N_4530,N_4223,N_4455);
or U4531 (N_4531,N_3925,N_3032);
or U4532 (N_4532,N_3096,N_3087);
and U4533 (N_4533,N_4055,N_4361);
nand U4534 (N_4534,N_3938,N_4188);
or U4535 (N_4535,N_4388,N_4251);
nor U4536 (N_4536,N_3208,N_4494);
and U4537 (N_4537,N_3305,N_3091);
and U4538 (N_4538,N_3370,N_3805);
and U4539 (N_4539,N_3318,N_4336);
nand U4540 (N_4540,N_4377,N_3759);
xnor U4541 (N_4541,N_3186,N_3730);
and U4542 (N_4542,N_3371,N_3578);
xor U4543 (N_4543,N_3320,N_4136);
and U4544 (N_4544,N_3888,N_3501);
nor U4545 (N_4545,N_3617,N_3051);
and U4546 (N_4546,N_4064,N_3952);
xnor U4547 (N_4547,N_4380,N_3285);
nor U4548 (N_4548,N_3898,N_3978);
nand U4549 (N_4549,N_3242,N_3233);
nor U4550 (N_4550,N_3591,N_3804);
nor U4551 (N_4551,N_4154,N_3418);
or U4552 (N_4552,N_4191,N_3024);
or U4553 (N_4553,N_3355,N_4238);
nand U4554 (N_4554,N_3330,N_4319);
nor U4555 (N_4555,N_3574,N_3048);
nand U4556 (N_4556,N_4213,N_3199);
or U4557 (N_4557,N_3620,N_4061);
or U4558 (N_4558,N_3140,N_3302);
and U4559 (N_4559,N_4021,N_4116);
or U4560 (N_4560,N_3402,N_3593);
and U4561 (N_4561,N_3442,N_3621);
nand U4562 (N_4562,N_3841,N_4199);
nand U4563 (N_4563,N_3426,N_4221);
nor U4564 (N_4564,N_3265,N_3935);
nor U4565 (N_4565,N_3890,N_4292);
xnor U4566 (N_4566,N_3178,N_3136);
and U4567 (N_4567,N_3369,N_4229);
nor U4568 (N_4568,N_3876,N_3860);
xor U4569 (N_4569,N_3072,N_3642);
nor U4570 (N_4570,N_3177,N_3245);
nor U4571 (N_4571,N_3459,N_3436);
or U4572 (N_4572,N_3201,N_3571);
nor U4573 (N_4573,N_3342,N_3594);
and U4574 (N_4574,N_3223,N_3774);
or U4575 (N_4575,N_4086,N_3545);
and U4576 (N_4576,N_3751,N_3517);
or U4577 (N_4577,N_3352,N_3650);
or U4578 (N_4578,N_3216,N_4446);
xor U4579 (N_4579,N_3530,N_3964);
and U4580 (N_4580,N_4282,N_3691);
and U4581 (N_4581,N_3811,N_3915);
or U4582 (N_4582,N_3602,N_4344);
nor U4583 (N_4583,N_3070,N_3120);
nor U4584 (N_4584,N_4009,N_3356);
nor U4585 (N_4585,N_4395,N_4484);
or U4586 (N_4586,N_3147,N_3509);
nand U4587 (N_4587,N_3084,N_3390);
and U4588 (N_4588,N_3328,N_4174);
nand U4589 (N_4589,N_3643,N_3891);
and U4590 (N_4590,N_3118,N_3117);
nor U4591 (N_4591,N_4190,N_3899);
xor U4592 (N_4592,N_3605,N_3026);
nor U4593 (N_4593,N_3664,N_4122);
nor U4594 (N_4594,N_3793,N_4333);
or U4595 (N_4595,N_3555,N_3071);
or U4596 (N_4596,N_3634,N_3060);
nand U4597 (N_4597,N_4070,N_3102);
and U4598 (N_4598,N_3174,N_3798);
or U4599 (N_4599,N_3552,N_3556);
nor U4600 (N_4600,N_3973,N_3999);
or U4601 (N_4601,N_4392,N_3554);
or U4602 (N_4602,N_3225,N_3912);
and U4603 (N_4603,N_4153,N_3412);
or U4604 (N_4604,N_3611,N_4385);
or U4605 (N_4605,N_3796,N_3050);
and U4606 (N_4606,N_3705,N_4075);
and U4607 (N_4607,N_3654,N_4060);
or U4608 (N_4608,N_3407,N_4131);
and U4609 (N_4609,N_3564,N_3904);
or U4610 (N_4610,N_3439,N_3281);
and U4611 (N_4611,N_4499,N_3403);
and U4612 (N_4612,N_4464,N_3706);
or U4613 (N_4613,N_3346,N_3969);
xnor U4614 (N_4614,N_3162,N_3303);
nor U4615 (N_4615,N_3236,N_4027);
and U4616 (N_4616,N_3493,N_4274);
or U4617 (N_4617,N_3470,N_4375);
or U4618 (N_4618,N_3893,N_3910);
nor U4619 (N_4619,N_4216,N_4417);
nor U4620 (N_4620,N_3538,N_3513);
and U4621 (N_4621,N_3648,N_3041);
nand U4622 (N_4622,N_3979,N_3042);
nor U4623 (N_4623,N_4204,N_4017);
nand U4624 (N_4624,N_3153,N_3894);
and U4625 (N_4625,N_3599,N_3704);
or U4626 (N_4626,N_3901,N_4365);
nor U4627 (N_4627,N_3840,N_4077);
and U4628 (N_4628,N_3139,N_3647);
and U4629 (N_4629,N_3731,N_3458);
nor U4630 (N_4630,N_3395,N_3406);
or U4631 (N_4631,N_4052,N_3966);
or U4632 (N_4632,N_4285,N_3815);
and U4633 (N_4633,N_4295,N_4324);
nand U4634 (N_4634,N_4401,N_3372);
nor U4635 (N_4635,N_3306,N_3974);
and U4636 (N_4636,N_3756,N_4124);
nor U4637 (N_4637,N_3638,N_4428);
nor U4638 (N_4638,N_3663,N_4102);
nand U4639 (N_4639,N_3007,N_4215);
nor U4640 (N_4640,N_3331,N_3504);
or U4641 (N_4641,N_3563,N_3018);
xnor U4642 (N_4642,N_4101,N_4327);
nor U4643 (N_4643,N_3625,N_4167);
nand U4644 (N_4644,N_3852,N_4130);
nand U4645 (N_4645,N_3404,N_4314);
nor U4646 (N_4646,N_4203,N_3019);
nand U4647 (N_4647,N_4486,N_3166);
and U4648 (N_4648,N_3172,N_4279);
nand U4649 (N_4649,N_4218,N_3188);
and U4650 (N_4650,N_3669,N_4110);
or U4651 (N_4651,N_4390,N_3657);
or U4652 (N_4652,N_3057,N_3833);
or U4653 (N_4653,N_4125,N_4449);
or U4654 (N_4654,N_3416,N_3760);
nand U4655 (N_4655,N_4193,N_3525);
nor U4656 (N_4656,N_3692,N_4054);
and U4657 (N_4657,N_4171,N_3639);
or U4658 (N_4658,N_3202,N_3719);
or U4659 (N_4659,N_4278,N_3918);
or U4660 (N_4660,N_3524,N_3856);
and U4661 (N_4661,N_3333,N_3741);
or U4662 (N_4662,N_3844,N_3336);
nand U4663 (N_4663,N_3825,N_3008);
or U4664 (N_4664,N_3849,N_4407);
or U4665 (N_4665,N_4043,N_3434);
and U4666 (N_4666,N_3635,N_3884);
nor U4667 (N_4667,N_3353,N_3921);
nand U4668 (N_4668,N_3733,N_4089);
or U4669 (N_4669,N_3887,N_4178);
nor U4670 (N_4670,N_3121,N_3247);
nand U4671 (N_4671,N_3762,N_4198);
or U4672 (N_4672,N_4097,N_4264);
nor U4673 (N_4673,N_4187,N_4414);
nor U4674 (N_4674,N_3702,N_3049);
or U4675 (N_4675,N_4042,N_4090);
or U4676 (N_4676,N_3113,N_3110);
nand U4677 (N_4677,N_3993,N_3401);
or U4678 (N_4678,N_3343,N_4160);
nand U4679 (N_4679,N_3949,N_4420);
and U4680 (N_4680,N_4355,N_4255);
nor U4681 (N_4681,N_3782,N_3035);
and U4682 (N_4682,N_4304,N_3073);
and U4683 (N_4683,N_3780,N_3322);
and U4684 (N_4684,N_3528,N_4049);
nor U4685 (N_4685,N_3507,N_3799);
or U4686 (N_4686,N_3765,N_3963);
nand U4687 (N_4687,N_3266,N_3772);
nand U4688 (N_4688,N_4242,N_4105);
nand U4689 (N_4689,N_3861,N_3445);
and U4690 (N_4690,N_3257,N_3359);
or U4691 (N_4691,N_4474,N_4138);
and U4692 (N_4692,N_3956,N_3607);
nor U4693 (N_4693,N_3671,N_3503);
nand U4694 (N_4694,N_3274,N_3033);
nand U4695 (N_4695,N_4100,N_3261);
and U4696 (N_4696,N_3766,N_4312);
or U4697 (N_4697,N_3827,N_3784);
and U4698 (N_4698,N_3540,N_4010);
or U4699 (N_4699,N_3532,N_4032);
nor U4700 (N_4700,N_3689,N_3011);
nand U4701 (N_4701,N_3075,N_3865);
or U4702 (N_4702,N_3697,N_4020);
and U4703 (N_4703,N_3002,N_3606);
and U4704 (N_4704,N_3249,N_3151);
nand U4705 (N_4705,N_4140,N_3258);
or U4706 (N_4706,N_3644,N_3809);
nand U4707 (N_4707,N_3830,N_3344);
or U4708 (N_4708,N_3488,N_4041);
nor U4709 (N_4709,N_4277,N_4487);
nor U4710 (N_4710,N_3149,N_3924);
or U4711 (N_4711,N_3325,N_4128);
nor U4712 (N_4712,N_4033,N_3690);
or U4713 (N_4713,N_3029,N_3821);
and U4714 (N_4714,N_3735,N_4416);
or U4715 (N_4715,N_3460,N_4400);
nand U4716 (N_4716,N_4293,N_4079);
and U4717 (N_4717,N_3196,N_3626);
and U4718 (N_4718,N_4311,N_4306);
nor U4719 (N_4719,N_3045,N_4240);
nand U4720 (N_4720,N_4429,N_3038);
nor U4721 (N_4721,N_4461,N_3400);
nor U4722 (N_4722,N_3946,N_3666);
nor U4723 (N_4723,N_3609,N_4479);
and U4724 (N_4724,N_3059,N_4107);
and U4725 (N_4725,N_3750,N_3491);
or U4726 (N_4726,N_4076,N_3655);
or U4727 (N_4727,N_3708,N_4029);
or U4728 (N_4728,N_4351,N_3679);
nor U4729 (N_4729,N_4335,N_4113);
nand U4730 (N_4730,N_4485,N_3848);
and U4731 (N_4731,N_4197,N_3577);
nor U4732 (N_4732,N_3729,N_4241);
and U4733 (N_4733,N_3596,N_4157);
xor U4734 (N_4734,N_4248,N_3929);
or U4735 (N_4735,N_3832,N_3985);
or U4736 (N_4736,N_4004,N_4127);
or U4737 (N_4737,N_3573,N_4452);
nand U4738 (N_4738,N_3585,N_3349);
and U4739 (N_4739,N_4129,N_4173);
nand U4740 (N_4740,N_3089,N_4145);
nand U4741 (N_4741,N_3997,N_4256);
nor U4742 (N_4742,N_3659,N_3211);
nand U4743 (N_4743,N_4120,N_3864);
and U4744 (N_4744,N_3478,N_4262);
or U4745 (N_4745,N_3662,N_4210);
nand U4746 (N_4746,N_3850,N_3695);
nand U4747 (N_4747,N_4258,N_3616);
or U4748 (N_4748,N_3364,N_4337);
nand U4749 (N_4749,N_3463,N_3300);
nor U4750 (N_4750,N_4393,N_4137);
or U4751 (N_4751,N_3119,N_3788);
nand U4752 (N_4752,N_3632,N_3630);
nor U4753 (N_4753,N_3219,N_3747);
nand U4754 (N_4754,N_3064,N_4068);
or U4755 (N_4755,N_3030,N_3080);
nor U4756 (N_4756,N_3358,N_4159);
nand U4757 (N_4757,N_4074,N_3975);
and U4758 (N_4758,N_3013,N_4423);
and U4759 (N_4759,N_3000,N_3467);
and U4760 (N_4760,N_3361,N_4315);
nor U4761 (N_4761,N_4189,N_4175);
nand U4762 (N_4762,N_4362,N_4364);
and U4763 (N_4763,N_3745,N_3843);
and U4764 (N_4764,N_4237,N_4371);
or U4765 (N_4765,N_3489,N_4334);
and U4766 (N_4766,N_3466,N_4287);
nor U4767 (N_4767,N_3673,N_3127);
and U4768 (N_4768,N_4007,N_4382);
or U4769 (N_4769,N_4270,N_3476);
or U4770 (N_4770,N_3264,N_3243);
or U4771 (N_4771,N_3173,N_4266);
and U4772 (N_4772,N_3256,N_3699);
or U4773 (N_4773,N_4104,N_3396);
nor U4774 (N_4774,N_4451,N_3549);
xnor U4775 (N_4775,N_3083,N_3180);
nor U4776 (N_4776,N_4212,N_4272);
or U4777 (N_4777,N_3753,N_3758);
nor U4778 (N_4778,N_4226,N_4252);
or U4779 (N_4779,N_3934,N_3781);
nand U4780 (N_4780,N_4263,N_3791);
or U4781 (N_4781,N_3304,N_3619);
and U4782 (N_4782,N_3871,N_3134);
nor U4783 (N_4783,N_3092,N_4348);
nand U4784 (N_4784,N_4083,N_3831);
nand U4785 (N_4785,N_3099,N_4245);
or U4786 (N_4786,N_3814,N_3794);
nand U4787 (N_4787,N_4069,N_4239);
nand U4788 (N_4788,N_3138,N_3276);
or U4789 (N_4789,N_3360,N_3877);
nand U4790 (N_4790,N_3338,N_4123);
nand U4791 (N_4791,N_3293,N_3646);
nor U4792 (N_4792,N_3828,N_4180);
and U4793 (N_4793,N_3942,N_4006);
nand U4794 (N_4794,N_3299,N_3472);
nor U4795 (N_4795,N_4040,N_4297);
or U4796 (N_4796,N_3937,N_4307);
nand U4797 (N_4797,N_3115,N_3449);
and U4798 (N_4798,N_3015,N_3768);
nand U4799 (N_4799,N_4481,N_3347);
nor U4800 (N_4800,N_3451,N_3253);
or U4801 (N_4801,N_4268,N_4179);
or U4802 (N_4802,N_3580,N_3713);
or U4803 (N_4803,N_3622,N_4425);
nor U4804 (N_4804,N_3195,N_3498);
nand U4805 (N_4805,N_3584,N_3853);
nor U4806 (N_4806,N_3283,N_3326);
nor U4807 (N_4807,N_4437,N_3623);
nand U4808 (N_4808,N_4384,N_4254);
nor U4809 (N_4809,N_3693,N_3785);
nand U4810 (N_4810,N_3204,N_3461);
or U4811 (N_4811,N_3640,N_3238);
nor U4812 (N_4812,N_3239,N_3490);
or U4813 (N_4813,N_4201,N_3327);
nand U4814 (N_4814,N_3357,N_4084);
nand U4815 (N_4815,N_3440,N_3475);
nand U4816 (N_4816,N_3754,N_3561);
or U4817 (N_4817,N_3221,N_3278);
and U4818 (N_4818,N_4477,N_3156);
nand U4819 (N_4819,N_3749,N_3539);
or U4820 (N_4820,N_3510,N_3259);
or U4821 (N_4821,N_4080,N_3824);
or U4822 (N_4822,N_3200,N_3570);
nor U4823 (N_4823,N_3900,N_4343);
or U4824 (N_4824,N_4466,N_3389);
or U4825 (N_4825,N_3380,N_4422);
xnor U4826 (N_4826,N_4402,N_3542);
nand U4827 (N_4827,N_4360,N_4030);
and U4828 (N_4828,N_3421,N_4099);
nand U4829 (N_4829,N_3222,N_3157);
and U4830 (N_4830,N_4339,N_4424);
or U4831 (N_4831,N_3520,N_3728);
and U4832 (N_4832,N_3977,N_4290);
or U4833 (N_4833,N_4207,N_3308);
and U4834 (N_4834,N_4170,N_3232);
or U4835 (N_4835,N_4396,N_3529);
or U4836 (N_4836,N_3712,N_4168);
nor U4837 (N_4837,N_3939,N_4313);
nand U4838 (N_4838,N_3755,N_3565);
or U4839 (N_4839,N_3567,N_4194);
or U4840 (N_4840,N_4296,N_3003);
or U4841 (N_4841,N_3348,N_3779);
or U4842 (N_4842,N_4353,N_3615);
nand U4843 (N_4843,N_3526,N_3618);
nor U4844 (N_4844,N_3430,N_3968);
and U4845 (N_4845,N_3290,N_4271);
and U4846 (N_4846,N_4026,N_4374);
and U4847 (N_4847,N_3629,N_4063);
nor U4848 (N_4848,N_3537,N_4412);
nor U4849 (N_4849,N_3911,N_3739);
or U4850 (N_4850,N_3280,N_3062);
or U4851 (N_4851,N_3313,N_3688);
nor U4852 (N_4852,N_3464,N_3012);
nand U4853 (N_4853,N_3989,N_4456);
nand U4854 (N_4854,N_3427,N_3531);
nor U4855 (N_4855,N_4162,N_3453);
or U4856 (N_4856,N_4284,N_4469);
and U4857 (N_4857,N_3586,N_4085);
and U4858 (N_4858,N_4118,N_3919);
nand U4859 (N_4859,N_4121,N_4244);
or U4860 (N_4860,N_3082,N_3835);
or U4861 (N_4861,N_3014,N_4146);
or U4862 (N_4862,N_3077,N_3727);
nand U4863 (N_4863,N_4236,N_3614);
xnor U4864 (N_4864,N_4067,N_4000);
nor U4865 (N_4865,N_4317,N_3954);
nor U4866 (N_4866,N_4460,N_3743);
and U4867 (N_4867,N_4430,N_3022);
or U4868 (N_4868,N_3652,N_4381);
nor U4869 (N_4869,N_3016,N_3725);
or U4870 (N_4870,N_3732,N_4098);
nor U4871 (N_4871,N_3129,N_3335);
or U4872 (N_4872,N_3958,N_3250);
and U4873 (N_4873,N_3587,N_3111);
and U4874 (N_4874,N_3943,N_3234);
or U4875 (N_4875,N_3496,N_3345);
nand U4876 (N_4876,N_3980,N_4294);
nand U4877 (N_4877,N_3066,N_3624);
nor U4878 (N_4878,N_3514,N_3499);
or U4879 (N_4879,N_3763,N_3267);
or U4880 (N_4880,N_3608,N_3044);
nor U4881 (N_4881,N_4413,N_3090);
nand U4882 (N_4882,N_3990,N_4016);
nor U4883 (N_4883,N_4147,N_3036);
or U4884 (N_4884,N_3382,N_3961);
or U4885 (N_4885,N_3773,N_3740);
or U4886 (N_4886,N_3229,N_3056);
and U4887 (N_4887,N_3481,N_3431);
or U4888 (N_4888,N_4117,N_3145);
or U4889 (N_4889,N_4039,N_4427);
or U4890 (N_4890,N_3193,N_3058);
and U4891 (N_4891,N_4303,N_4139);
and U4892 (N_4892,N_3321,N_3546);
and U4893 (N_4893,N_3883,N_3213);
nor U4894 (N_4894,N_3681,N_3107);
and U4895 (N_4895,N_3895,N_3583);
nor U4896 (N_4896,N_4209,N_4051);
or U4897 (N_4897,N_3922,N_3685);
or U4898 (N_4898,N_3423,N_4112);
or U4899 (N_4899,N_3209,N_3387);
or U4900 (N_4900,N_3137,N_3757);
nor U4901 (N_4901,N_3473,N_3164);
and U4902 (N_4902,N_3428,N_3736);
nor U4903 (N_4903,N_3296,N_3154);
nand U4904 (N_4904,N_3721,N_3738);
or U4905 (N_4905,N_3926,N_4114);
or U4906 (N_4906,N_4433,N_4024);
nor U4907 (N_4907,N_4059,N_3950);
or U4908 (N_4908,N_4096,N_3649);
nand U4909 (N_4909,N_4322,N_3198);
and U4910 (N_4910,N_3377,N_4291);
and U4911 (N_4911,N_3192,N_3636);
or U4912 (N_4912,N_3886,N_3786);
or U4913 (N_4913,N_4232,N_3881);
or U4914 (N_4914,N_3711,N_4246);
nand U4915 (N_4915,N_4230,N_3160);
or U4916 (N_4916,N_3857,N_3764);
nand U4917 (N_4917,N_3873,N_3734);
or U4918 (N_4918,N_3604,N_3397);
and U4919 (N_4919,N_3350,N_4163);
or U4920 (N_4920,N_3519,N_3437);
nand U4921 (N_4921,N_3866,N_3432);
nor U4922 (N_4922,N_3462,N_3516);
nor U4923 (N_4923,N_3068,N_4471);
nand U4924 (N_4924,N_3955,N_3903);
nand U4925 (N_4925,N_4135,N_3581);
nand U4926 (N_4926,N_3506,N_3933);
and U4927 (N_4927,N_3645,N_3052);
or U4928 (N_4928,N_4144,N_4359);
nand U4929 (N_4929,N_4045,N_3131);
nand U4930 (N_4930,N_3592,N_4091);
or U4931 (N_4931,N_4298,N_4259);
nand U4932 (N_4932,N_4345,N_4426);
nand U4933 (N_4933,N_3896,N_4225);
nor U4934 (N_4934,N_3744,N_4493);
or U4935 (N_4935,N_4342,N_4058);
and U4936 (N_4936,N_3559,N_4034);
or U4937 (N_4937,N_4286,N_4320);
nor U4938 (N_4938,N_3703,N_3874);
or U4939 (N_4939,N_4288,N_3778);
nor U4940 (N_4940,N_4148,N_3409);
nand U4941 (N_4941,N_3527,N_3595);
nor U4942 (N_4942,N_3309,N_3771);
or U4943 (N_4943,N_3424,N_3813);
or U4944 (N_4944,N_4195,N_3373);
nand U4945 (N_4945,N_4050,N_3363);
and U4946 (N_4946,N_3672,N_3812);
nand U4947 (N_4947,N_3882,N_3047);
nand U4948 (N_4948,N_4326,N_3568);
and U4949 (N_4949,N_3315,N_3709);
or U4950 (N_4950,N_4141,N_3190);
or U4951 (N_4951,N_4358,N_3135);
nor U4952 (N_4952,N_3670,N_4177);
nor U4953 (N_4953,N_3631,N_4106);
nand U4954 (N_4954,N_4011,N_4149);
or U4955 (N_4955,N_3078,N_3823);
nor U4956 (N_4956,N_4418,N_3125);
and U4957 (N_4957,N_4346,N_4235);
nor U4958 (N_4958,N_4005,N_3025);
and U4959 (N_4959,N_3505,N_3067);
nor U4960 (N_4960,N_3181,N_3142);
or U4961 (N_4961,N_3471,N_4458);
nor U4962 (N_4962,N_4489,N_3547);
nand U4963 (N_4963,N_3179,N_3085);
nor U4964 (N_4964,N_4301,N_4328);
and U4965 (N_4965,N_3737,N_3448);
or U4966 (N_4966,N_3905,N_3790);
nand U4967 (N_4967,N_3996,N_3103);
xor U4968 (N_4968,N_4028,N_4386);
nand U4969 (N_4969,N_4442,N_3720);
nand U4970 (N_4970,N_3548,N_4176);
nor U4971 (N_4971,N_3512,N_3589);
nor U4972 (N_4972,N_3917,N_3109);
and U4973 (N_4973,N_3674,N_3108);
or U4974 (N_4974,N_3536,N_4445);
nor U4975 (N_4975,N_4357,N_3405);
or U4976 (N_4976,N_3194,N_4152);
nor U4977 (N_4977,N_3701,N_4289);
and U4978 (N_4978,N_3101,N_3859);
and U4979 (N_4979,N_3523,N_3959);
or U4980 (N_4980,N_4062,N_3144);
or U4981 (N_4981,N_3947,N_3834);
nor U4982 (N_4982,N_3722,N_3433);
nand U4983 (N_4983,N_4308,N_3301);
or U4984 (N_4984,N_3425,N_3061);
or U4985 (N_4985,N_3858,N_3130);
nor U4986 (N_4986,N_3212,N_3240);
or U4987 (N_4987,N_4081,N_3970);
or U4988 (N_4988,N_3992,N_4419);
or U4989 (N_4989,N_3665,N_4234);
and U4990 (N_4990,N_3716,N_4132);
nand U4991 (N_4991,N_4283,N_4073);
or U4992 (N_4992,N_4454,N_4186);
nor U4993 (N_4993,N_4480,N_3141);
or U4994 (N_4994,N_3368,N_4228);
nor U4995 (N_4995,N_3682,N_4387);
or U4996 (N_4996,N_3579,N_4373);
nor U4997 (N_4997,N_3340,N_4224);
nor U4998 (N_4998,N_3446,N_3575);
and U4999 (N_4999,N_4253,N_3783);
or U5000 (N_5000,N_3230,N_4495);
or U5001 (N_5001,N_3217,N_4276);
nand U5002 (N_5002,N_4404,N_3100);
nor U5003 (N_5003,N_4088,N_4181);
and U5004 (N_5004,N_3189,N_4094);
or U5005 (N_5005,N_4447,N_4119);
or U5006 (N_5006,N_3653,N_3566);
nor U5007 (N_5007,N_3714,N_3168);
nor U5008 (N_5008,N_4305,N_3414);
nand U5009 (N_5009,N_4111,N_3271);
nand U5010 (N_5010,N_3184,N_3452);
nand U5011 (N_5011,N_4182,N_3122);
or U5012 (N_5012,N_3220,N_4184);
xnor U5013 (N_5013,N_3847,N_3656);
or U5014 (N_5014,N_3494,N_4164);
and U5015 (N_5015,N_3889,N_4453);
or U5016 (N_5016,N_4463,N_3541);
nor U5017 (N_5017,N_3839,N_4161);
or U5018 (N_5018,N_3367,N_3601);
nor U5019 (N_5019,N_3319,N_3287);
or U5020 (N_5020,N_4151,N_4309);
or U5021 (N_5021,N_3962,N_3916);
or U5022 (N_5022,N_3133,N_4347);
nand U5023 (N_5023,N_3284,N_3295);
xor U5024 (N_5024,N_3098,N_4367);
or U5025 (N_5025,N_4352,N_4219);
nand U5026 (N_5026,N_4332,N_3913);
or U5027 (N_5027,N_4403,N_4038);
nor U5028 (N_5028,N_3880,N_4165);
or U5029 (N_5029,N_4095,N_3429);
or U5030 (N_5030,N_3224,N_4299);
nor U5031 (N_5031,N_3930,N_3998);
nor U5032 (N_5032,N_4325,N_3867);
nor U5033 (N_5033,N_4378,N_3386);
or U5034 (N_5034,N_4468,N_3715);
nand U5035 (N_5035,N_3104,N_3497);
nand U5036 (N_5036,N_4441,N_4397);
and U5037 (N_5037,N_3752,N_4376);
nor U5038 (N_5038,N_3231,N_3063);
or U5039 (N_5039,N_4166,N_3515);
nor U5040 (N_5040,N_3846,N_4492);
or U5041 (N_5041,N_3972,N_4323);
nor U5042 (N_5042,N_3312,N_4217);
nor U5043 (N_5043,N_3251,N_3097);
and U5044 (N_5044,N_3043,N_3408);
or U5045 (N_5045,N_4280,N_3422);
nand U5046 (N_5046,N_3795,N_3272);
nand U5047 (N_5047,N_3399,N_3633);
nor U5048 (N_5048,N_4250,N_3094);
xnor U5049 (N_5049,N_4318,N_3661);
nor U5050 (N_5050,N_3582,N_3398);
and U5051 (N_5051,N_3872,N_3870);
nor U5052 (N_5052,N_3028,N_3598);
and U5053 (N_5053,N_4354,N_4103);
or U5054 (N_5054,N_3694,N_3957);
nor U5055 (N_5055,N_3411,N_4331);
nand U5056 (N_5056,N_3388,N_3443);
or U5057 (N_5057,N_3158,N_3660);
xnor U5058 (N_5058,N_4338,N_3802);
nor U5059 (N_5059,N_3005,N_4363);
nand U5060 (N_5060,N_4108,N_3726);
nor U5061 (N_5061,N_4434,N_3855);
and U5062 (N_5062,N_3337,N_3678);
or U5063 (N_5063,N_3376,N_3246);
nor U5064 (N_5064,N_3769,N_3329);
or U5065 (N_5065,N_3215,N_4302);
or U5066 (N_5066,N_4415,N_4497);
or U5067 (N_5067,N_4214,N_3001);
and U5068 (N_5068,N_3909,N_4227);
and U5069 (N_5069,N_4044,N_3550);
xor U5070 (N_5070,N_3105,N_3165);
or U5071 (N_5071,N_3522,N_4202);
nor U5072 (N_5072,N_3502,N_3324);
nand U5073 (N_5073,N_4001,N_3126);
nor U5074 (N_5074,N_3603,N_3535);
nand U5075 (N_5075,N_3183,N_3037);
or U5076 (N_5076,N_3334,N_3612);
nand U5077 (N_5077,N_3819,N_3967);
nand U5078 (N_5078,N_3534,N_3065);
or U5079 (N_5079,N_3384,N_3175);
nand U5080 (N_5080,N_4379,N_3684);
nor U5081 (N_5081,N_3055,N_4018);
nor U5082 (N_5082,N_3914,N_3869);
or U5083 (N_5083,N_3862,N_3020);
and U5084 (N_5084,N_3341,N_3810);
nor U5085 (N_5085,N_4443,N_3093);
nand U5086 (N_5086,N_3486,N_3323);
and U5087 (N_5087,N_4008,N_3988);
and U5088 (N_5088,N_4448,N_4012);
or U5089 (N_5089,N_3482,N_4465);
nor U5090 (N_5090,N_4222,N_3558);
nand U5091 (N_5091,N_3484,N_4019);
nor U5092 (N_5092,N_4126,N_4022);
or U5093 (N_5093,N_3907,N_4158);
and U5094 (N_5094,N_3641,N_3986);
and U5095 (N_5095,N_3878,N_4391);
and U5096 (N_5096,N_4490,N_3379);
nor U5097 (N_5097,N_4093,N_4247);
or U5098 (N_5098,N_4071,N_3269);
and U5099 (N_5099,N_3474,N_4142);
or U5100 (N_5100,N_4133,N_3441);
or U5101 (N_5101,N_4438,N_3053);
and U5102 (N_5102,N_3438,N_3590);
nand U5103 (N_5103,N_3995,N_4340);
xnor U5104 (N_5104,N_3816,N_4047);
and U5105 (N_5105,N_4411,N_4369);
or U5106 (N_5106,N_4269,N_3868);
nand U5107 (N_5107,N_4072,N_3455);
nand U5108 (N_5108,N_3767,N_4349);
nand U5109 (N_5109,N_3851,N_3508);
or U5110 (N_5110,N_3553,N_4473);
or U5111 (N_5111,N_3205,N_3818);
nand U5112 (N_5112,N_3976,N_3836);
nand U5113 (N_5113,N_3842,N_3700);
and U5114 (N_5114,N_3206,N_4457);
xnor U5115 (N_5115,N_3235,N_4267);
nor U5116 (N_5116,N_3314,N_4491);
nand U5117 (N_5117,N_3981,N_3366);
nand U5118 (N_5118,N_4483,N_3351);
nor U5119 (N_5119,N_3081,N_4134);
or U5120 (N_5120,N_3410,N_3710);
and U5121 (N_5121,N_3273,N_3588);
nor U5122 (N_5122,N_4439,N_3457);
or U5123 (N_5123,N_3148,N_3707);
nand U5124 (N_5124,N_3469,N_3696);
nor U5125 (N_5125,N_3317,N_3454);
or U5126 (N_5126,N_3447,N_4233);
or U5127 (N_5127,N_4053,N_4109);
xor U5128 (N_5128,N_3518,N_3444);
nand U5129 (N_5129,N_3171,N_3822);
or U5130 (N_5130,N_4150,N_3748);
or U5131 (N_5131,N_3544,N_3500);
or U5132 (N_5132,N_3074,N_3854);
nor U5133 (N_5133,N_4013,N_4356);
or U5134 (N_5134,N_3724,N_3492);
nor U5135 (N_5135,N_3237,N_3863);
nand U5136 (N_5136,N_4341,N_3932);
nor U5137 (N_5137,N_4472,N_3717);
or U5138 (N_5138,N_3477,N_4155);
and U5139 (N_5139,N_3885,N_3906);
nor U5140 (N_5140,N_4273,N_3613);
nand U5141 (N_5141,N_3248,N_3241);
nor U5142 (N_5142,N_3210,N_3027);
nor U5143 (N_5143,N_3667,N_3829);
and U5144 (N_5144,N_3375,N_3761);
nand U5145 (N_5145,N_3374,N_3465);
or U5146 (N_5146,N_3106,N_3944);
and U5147 (N_5147,N_3079,N_3383);
nand U5148 (N_5148,N_3040,N_3808);
xnor U5149 (N_5149,N_3483,N_3069);
nor U5150 (N_5150,N_3610,N_3479);
nand U5151 (N_5151,N_4408,N_4057);
or U5152 (N_5152,N_3054,N_4092);
and U5153 (N_5153,N_4048,N_3817);
nand U5154 (N_5154,N_3034,N_3270);
and U5155 (N_5155,N_4488,N_3845);
nand U5156 (N_5156,N_4459,N_4257);
or U5157 (N_5157,N_4436,N_3086);
and U5158 (N_5158,N_3551,N_3803);
nor U5159 (N_5159,N_3297,N_3227);
or U5160 (N_5160,N_4405,N_3468);
nand U5161 (N_5161,N_3480,N_4421);
nor U5162 (N_5162,N_3923,N_3936);
nor U5163 (N_5163,N_4368,N_3185);
nor U5164 (N_5164,N_3381,N_4015);
nand U5165 (N_5165,N_3046,N_3777);
or U5166 (N_5166,N_3920,N_3675);
or U5167 (N_5167,N_3146,N_4409);
or U5168 (N_5168,N_3965,N_3982);
or U5169 (N_5169,N_3039,N_3543);
nand U5170 (N_5170,N_4143,N_3837);
and U5171 (N_5171,N_3332,N_3262);
nor U5172 (N_5172,N_4036,N_4275);
and U5173 (N_5173,N_4211,N_4482);
or U5174 (N_5174,N_4231,N_3112);
nor U5175 (N_5175,N_3282,N_4037);
or U5176 (N_5176,N_3114,N_3392);
nor U5177 (N_5177,N_3354,N_4183);
or U5178 (N_5178,N_3021,N_3187);
or U5179 (N_5179,N_3150,N_3277);
or U5180 (N_5180,N_3994,N_4261);
or U5181 (N_5181,N_4470,N_3627);
nor U5182 (N_5182,N_3940,N_4310);
and U5183 (N_5183,N_3838,N_4065);
nor U5184 (N_5184,N_3316,N_3420);
or U5185 (N_5185,N_4205,N_3807);
and U5186 (N_5186,N_3987,N_4462);
and U5187 (N_5187,N_4444,N_4260);
or U5188 (N_5188,N_4206,N_3792);
or U5189 (N_5189,N_4185,N_3004);
nand U5190 (N_5190,N_4406,N_3533);
and U5191 (N_5191,N_3687,N_3176);
nor U5192 (N_5192,N_3742,N_3562);
and U5193 (N_5193,N_3677,N_3557);
nand U5194 (N_5194,N_3826,N_3718);
and U5195 (N_5195,N_4321,N_3875);
nor U5196 (N_5196,N_3971,N_3628);
nand U5197 (N_5197,N_4496,N_3775);
or U5198 (N_5198,N_3152,N_4435);
nor U5199 (N_5199,N_3132,N_3006);
nand U5200 (N_5200,N_3252,N_3801);
and U5201 (N_5201,N_3770,N_3560);
nand U5202 (N_5202,N_3031,N_3686);
and U5203 (N_5203,N_3289,N_4196);
xnor U5204 (N_5204,N_4208,N_3155);
nor U5205 (N_5205,N_3169,N_3879);
or U5206 (N_5206,N_4078,N_4281);
nor U5207 (N_5207,N_4383,N_3941);
xor U5208 (N_5208,N_4440,N_3393);
or U5209 (N_5209,N_4410,N_3511);
and U5210 (N_5210,N_3163,N_3984);
or U5211 (N_5211,N_3600,N_3286);
and U5212 (N_5212,N_3263,N_3450);
and U5213 (N_5213,N_3275,N_3698);
and U5214 (N_5214,N_3116,N_3009);
xor U5215 (N_5215,N_3159,N_3143);
nand U5216 (N_5216,N_3288,N_4082);
and U5217 (N_5217,N_3311,N_3226);
and U5218 (N_5218,N_4046,N_3789);
nor U5219 (N_5219,N_3417,N_4025);
or U5220 (N_5220,N_3680,N_4243);
nand U5221 (N_5221,N_4432,N_3658);
nand U5222 (N_5222,N_3413,N_3521);
nand U5223 (N_5223,N_4476,N_3951);
nand U5224 (N_5224,N_3076,N_3298);
and U5225 (N_5225,N_4398,N_3244);
or U5226 (N_5226,N_3291,N_4156);
and U5227 (N_5227,N_4366,N_3897);
nand U5228 (N_5228,N_3945,N_4329);
and U5229 (N_5229,N_3182,N_4316);
nand U5230 (N_5230,N_3415,N_3746);
and U5231 (N_5231,N_3928,N_4056);
xnor U5232 (N_5232,N_3487,N_4035);
nor U5233 (N_5233,N_3207,N_4200);
or U5234 (N_5234,N_3385,N_4066);
nor U5235 (N_5235,N_3124,N_4431);
nand U5236 (N_5236,N_3495,N_3365);
nor U5237 (N_5237,N_4087,N_3902);
xnor U5238 (N_5238,N_3214,N_3023);
nand U5239 (N_5239,N_3435,N_4192);
nand U5240 (N_5240,N_3197,N_3010);
nand U5241 (N_5241,N_3800,N_3391);
or U5242 (N_5242,N_3991,N_3927);
nand U5243 (N_5243,N_4372,N_3279);
nor U5244 (N_5244,N_3569,N_3128);
or U5245 (N_5245,N_3892,N_3378);
xor U5246 (N_5246,N_3294,N_3806);
nor U5247 (N_5247,N_3651,N_3953);
or U5248 (N_5248,N_3260,N_4300);
or U5249 (N_5249,N_3668,N_4031);
nand U5250 (N_5250,N_4006,N_3510);
nor U5251 (N_5251,N_3031,N_3802);
and U5252 (N_5252,N_3443,N_3936);
nand U5253 (N_5253,N_3341,N_3775);
nand U5254 (N_5254,N_3219,N_3562);
nand U5255 (N_5255,N_3263,N_3962);
nand U5256 (N_5256,N_3439,N_3272);
or U5257 (N_5257,N_3024,N_3382);
nor U5258 (N_5258,N_4281,N_4092);
nand U5259 (N_5259,N_3165,N_3979);
xor U5260 (N_5260,N_3112,N_3656);
and U5261 (N_5261,N_3879,N_3855);
nor U5262 (N_5262,N_3135,N_3317);
or U5263 (N_5263,N_4373,N_3994);
nand U5264 (N_5264,N_3192,N_3047);
nor U5265 (N_5265,N_3022,N_3308);
and U5266 (N_5266,N_3145,N_4456);
or U5267 (N_5267,N_3086,N_3986);
and U5268 (N_5268,N_4114,N_4331);
nand U5269 (N_5269,N_3242,N_4473);
nand U5270 (N_5270,N_3166,N_3349);
and U5271 (N_5271,N_3508,N_4204);
nor U5272 (N_5272,N_3813,N_4240);
nor U5273 (N_5273,N_3715,N_3476);
nand U5274 (N_5274,N_3805,N_3976);
and U5275 (N_5275,N_3424,N_3112);
nor U5276 (N_5276,N_3595,N_4430);
and U5277 (N_5277,N_3415,N_3775);
and U5278 (N_5278,N_3102,N_3836);
nand U5279 (N_5279,N_3781,N_3505);
or U5280 (N_5280,N_4041,N_3739);
and U5281 (N_5281,N_3733,N_3605);
nor U5282 (N_5282,N_3174,N_3387);
nand U5283 (N_5283,N_3048,N_4175);
and U5284 (N_5284,N_3031,N_4476);
and U5285 (N_5285,N_3474,N_3802);
and U5286 (N_5286,N_3224,N_3909);
nand U5287 (N_5287,N_3348,N_4327);
or U5288 (N_5288,N_3069,N_4359);
and U5289 (N_5289,N_3041,N_4146);
or U5290 (N_5290,N_3842,N_3775);
nand U5291 (N_5291,N_4336,N_3915);
and U5292 (N_5292,N_3260,N_4222);
nor U5293 (N_5293,N_4336,N_4150);
nor U5294 (N_5294,N_3475,N_3625);
nor U5295 (N_5295,N_4258,N_3301);
or U5296 (N_5296,N_3342,N_4207);
nor U5297 (N_5297,N_3224,N_4268);
nand U5298 (N_5298,N_3590,N_4181);
nor U5299 (N_5299,N_4178,N_4118);
or U5300 (N_5300,N_4316,N_4205);
nor U5301 (N_5301,N_4030,N_3473);
nand U5302 (N_5302,N_3192,N_3680);
nor U5303 (N_5303,N_4487,N_3520);
and U5304 (N_5304,N_4036,N_4493);
and U5305 (N_5305,N_3481,N_3075);
or U5306 (N_5306,N_4022,N_3852);
and U5307 (N_5307,N_3012,N_3566);
nand U5308 (N_5308,N_3856,N_3478);
and U5309 (N_5309,N_3425,N_3736);
nor U5310 (N_5310,N_3090,N_3241);
nand U5311 (N_5311,N_4224,N_3178);
or U5312 (N_5312,N_4201,N_4141);
or U5313 (N_5313,N_3306,N_4064);
nand U5314 (N_5314,N_4318,N_3659);
or U5315 (N_5315,N_4118,N_4258);
xor U5316 (N_5316,N_4143,N_3835);
or U5317 (N_5317,N_3515,N_3600);
xor U5318 (N_5318,N_3075,N_4424);
and U5319 (N_5319,N_3319,N_3692);
and U5320 (N_5320,N_3383,N_3629);
nor U5321 (N_5321,N_3543,N_3813);
and U5322 (N_5322,N_4141,N_3058);
nor U5323 (N_5323,N_3002,N_3902);
and U5324 (N_5324,N_4031,N_3213);
nor U5325 (N_5325,N_4286,N_4259);
or U5326 (N_5326,N_3244,N_3392);
or U5327 (N_5327,N_4122,N_4029);
and U5328 (N_5328,N_3816,N_3287);
or U5329 (N_5329,N_4199,N_4090);
and U5330 (N_5330,N_3878,N_3345);
nand U5331 (N_5331,N_4311,N_3716);
xor U5332 (N_5332,N_3705,N_3636);
nor U5333 (N_5333,N_4466,N_3463);
nand U5334 (N_5334,N_3918,N_3808);
and U5335 (N_5335,N_3924,N_4266);
or U5336 (N_5336,N_4129,N_3386);
nor U5337 (N_5337,N_3635,N_4324);
and U5338 (N_5338,N_4268,N_3943);
nor U5339 (N_5339,N_3062,N_3263);
and U5340 (N_5340,N_4010,N_4113);
and U5341 (N_5341,N_3683,N_3010);
nand U5342 (N_5342,N_3847,N_4217);
nand U5343 (N_5343,N_3119,N_3626);
or U5344 (N_5344,N_3473,N_3715);
and U5345 (N_5345,N_3535,N_4197);
and U5346 (N_5346,N_3888,N_3122);
or U5347 (N_5347,N_3978,N_3799);
and U5348 (N_5348,N_3187,N_3374);
or U5349 (N_5349,N_4421,N_3241);
or U5350 (N_5350,N_4441,N_4156);
or U5351 (N_5351,N_3227,N_3622);
xnor U5352 (N_5352,N_3573,N_3680);
nand U5353 (N_5353,N_4079,N_3060);
or U5354 (N_5354,N_4146,N_3337);
nor U5355 (N_5355,N_3847,N_4277);
nand U5356 (N_5356,N_3015,N_4171);
nand U5357 (N_5357,N_3756,N_4050);
and U5358 (N_5358,N_4202,N_3565);
nor U5359 (N_5359,N_3936,N_3582);
and U5360 (N_5360,N_3508,N_3568);
or U5361 (N_5361,N_3410,N_3127);
nor U5362 (N_5362,N_3519,N_4247);
nor U5363 (N_5363,N_3316,N_3126);
and U5364 (N_5364,N_3913,N_3672);
or U5365 (N_5365,N_4008,N_4049);
nand U5366 (N_5366,N_3088,N_3806);
nand U5367 (N_5367,N_3975,N_4246);
and U5368 (N_5368,N_4155,N_3828);
nand U5369 (N_5369,N_3429,N_3457);
nor U5370 (N_5370,N_4214,N_4375);
nor U5371 (N_5371,N_3776,N_3634);
nor U5372 (N_5372,N_4097,N_4061);
and U5373 (N_5373,N_3808,N_4020);
and U5374 (N_5374,N_3202,N_4030);
or U5375 (N_5375,N_3285,N_4104);
nand U5376 (N_5376,N_4203,N_3790);
or U5377 (N_5377,N_3063,N_3548);
nor U5378 (N_5378,N_3224,N_4317);
xnor U5379 (N_5379,N_3182,N_3614);
nor U5380 (N_5380,N_3896,N_3995);
nand U5381 (N_5381,N_4321,N_3287);
and U5382 (N_5382,N_3695,N_4141);
nand U5383 (N_5383,N_4380,N_3792);
nand U5384 (N_5384,N_3182,N_3545);
or U5385 (N_5385,N_4096,N_3742);
or U5386 (N_5386,N_3923,N_3887);
nor U5387 (N_5387,N_4405,N_3911);
and U5388 (N_5388,N_4279,N_3121);
nor U5389 (N_5389,N_3602,N_3670);
and U5390 (N_5390,N_3053,N_3209);
nand U5391 (N_5391,N_3987,N_3998);
and U5392 (N_5392,N_3648,N_3268);
nand U5393 (N_5393,N_4121,N_3644);
or U5394 (N_5394,N_4368,N_3680);
nor U5395 (N_5395,N_4094,N_4446);
or U5396 (N_5396,N_3750,N_3290);
nor U5397 (N_5397,N_3542,N_3067);
nand U5398 (N_5398,N_3350,N_3330);
nand U5399 (N_5399,N_3620,N_3444);
and U5400 (N_5400,N_3745,N_3656);
nor U5401 (N_5401,N_3380,N_3347);
nor U5402 (N_5402,N_3144,N_3118);
or U5403 (N_5403,N_3105,N_3591);
or U5404 (N_5404,N_4176,N_3143);
nand U5405 (N_5405,N_3180,N_4113);
xnor U5406 (N_5406,N_3865,N_4145);
or U5407 (N_5407,N_3882,N_4208);
and U5408 (N_5408,N_3582,N_3982);
or U5409 (N_5409,N_3310,N_3551);
and U5410 (N_5410,N_4240,N_4046);
nand U5411 (N_5411,N_3857,N_3537);
nor U5412 (N_5412,N_3508,N_4266);
xor U5413 (N_5413,N_4013,N_3220);
nor U5414 (N_5414,N_4484,N_3118);
nand U5415 (N_5415,N_4290,N_3710);
nor U5416 (N_5416,N_4112,N_3159);
nor U5417 (N_5417,N_3750,N_4037);
or U5418 (N_5418,N_3872,N_3429);
or U5419 (N_5419,N_3632,N_3143);
and U5420 (N_5420,N_3880,N_3538);
nand U5421 (N_5421,N_3530,N_4249);
or U5422 (N_5422,N_3404,N_3550);
and U5423 (N_5423,N_4024,N_3544);
and U5424 (N_5424,N_4472,N_3633);
and U5425 (N_5425,N_3127,N_3434);
or U5426 (N_5426,N_3514,N_4390);
nor U5427 (N_5427,N_3952,N_4109);
nor U5428 (N_5428,N_3409,N_3235);
and U5429 (N_5429,N_3717,N_3483);
nand U5430 (N_5430,N_3993,N_3523);
nand U5431 (N_5431,N_3367,N_4152);
nand U5432 (N_5432,N_3378,N_3397);
xor U5433 (N_5433,N_4215,N_4483);
nor U5434 (N_5434,N_3860,N_3932);
nand U5435 (N_5435,N_3210,N_3484);
nand U5436 (N_5436,N_3684,N_3181);
nand U5437 (N_5437,N_3149,N_4426);
nor U5438 (N_5438,N_3727,N_4101);
xnor U5439 (N_5439,N_3348,N_4123);
and U5440 (N_5440,N_4487,N_4316);
and U5441 (N_5441,N_3214,N_3653);
nor U5442 (N_5442,N_3060,N_3486);
nor U5443 (N_5443,N_3013,N_4299);
or U5444 (N_5444,N_3501,N_3278);
nand U5445 (N_5445,N_3016,N_3974);
or U5446 (N_5446,N_3053,N_4329);
or U5447 (N_5447,N_3289,N_3038);
nor U5448 (N_5448,N_3551,N_3687);
nand U5449 (N_5449,N_3349,N_4354);
nand U5450 (N_5450,N_4083,N_3857);
nand U5451 (N_5451,N_3141,N_3034);
or U5452 (N_5452,N_3226,N_3385);
nor U5453 (N_5453,N_3711,N_3452);
nor U5454 (N_5454,N_3033,N_3288);
and U5455 (N_5455,N_3201,N_3897);
and U5456 (N_5456,N_3274,N_4144);
or U5457 (N_5457,N_3149,N_3325);
nor U5458 (N_5458,N_4478,N_3039);
xnor U5459 (N_5459,N_4058,N_4214);
and U5460 (N_5460,N_3577,N_3837);
nor U5461 (N_5461,N_3392,N_3671);
nor U5462 (N_5462,N_3884,N_3959);
and U5463 (N_5463,N_4121,N_4169);
nor U5464 (N_5464,N_4441,N_4260);
nor U5465 (N_5465,N_3210,N_4109);
nand U5466 (N_5466,N_4370,N_4359);
and U5467 (N_5467,N_3296,N_3604);
or U5468 (N_5468,N_3108,N_3648);
and U5469 (N_5469,N_3793,N_3965);
nor U5470 (N_5470,N_3458,N_4273);
nor U5471 (N_5471,N_4037,N_3218);
or U5472 (N_5472,N_3364,N_3335);
nor U5473 (N_5473,N_4053,N_4156);
nand U5474 (N_5474,N_3548,N_3275);
or U5475 (N_5475,N_3210,N_4471);
nand U5476 (N_5476,N_3771,N_4372);
xnor U5477 (N_5477,N_4329,N_3328);
nand U5478 (N_5478,N_3629,N_3335);
and U5479 (N_5479,N_3955,N_4080);
nor U5480 (N_5480,N_3536,N_3797);
nand U5481 (N_5481,N_4483,N_4232);
and U5482 (N_5482,N_3207,N_3844);
and U5483 (N_5483,N_4032,N_4191);
and U5484 (N_5484,N_3984,N_3948);
or U5485 (N_5485,N_3226,N_3924);
nor U5486 (N_5486,N_3461,N_3915);
nand U5487 (N_5487,N_3285,N_3939);
or U5488 (N_5488,N_4354,N_3299);
or U5489 (N_5489,N_4082,N_3113);
and U5490 (N_5490,N_4180,N_3341);
xnor U5491 (N_5491,N_3296,N_3110);
nand U5492 (N_5492,N_4437,N_3065);
nand U5493 (N_5493,N_3162,N_3697);
and U5494 (N_5494,N_3744,N_3978);
and U5495 (N_5495,N_3368,N_3647);
and U5496 (N_5496,N_3012,N_3787);
nor U5497 (N_5497,N_3927,N_4051);
or U5498 (N_5498,N_3594,N_4163);
nand U5499 (N_5499,N_3988,N_3304);
or U5500 (N_5500,N_3192,N_4221);
or U5501 (N_5501,N_3181,N_3812);
or U5502 (N_5502,N_3033,N_3241);
and U5503 (N_5503,N_3846,N_4130);
nand U5504 (N_5504,N_3479,N_3090);
and U5505 (N_5505,N_3618,N_3572);
nand U5506 (N_5506,N_3543,N_3728);
or U5507 (N_5507,N_3724,N_3691);
or U5508 (N_5508,N_3846,N_4110);
nor U5509 (N_5509,N_3878,N_3402);
or U5510 (N_5510,N_3275,N_4108);
and U5511 (N_5511,N_4089,N_4321);
nor U5512 (N_5512,N_3381,N_3875);
nand U5513 (N_5513,N_3801,N_3101);
nand U5514 (N_5514,N_3028,N_3126);
and U5515 (N_5515,N_3528,N_3633);
nand U5516 (N_5516,N_3859,N_3392);
and U5517 (N_5517,N_4025,N_3346);
nor U5518 (N_5518,N_3516,N_4396);
and U5519 (N_5519,N_3258,N_4122);
or U5520 (N_5520,N_3097,N_4077);
nand U5521 (N_5521,N_3121,N_4089);
nand U5522 (N_5522,N_4465,N_4096);
nand U5523 (N_5523,N_3951,N_3464);
nor U5524 (N_5524,N_3497,N_3679);
nor U5525 (N_5525,N_4146,N_3350);
nor U5526 (N_5526,N_3234,N_4489);
nor U5527 (N_5527,N_3113,N_4270);
nor U5528 (N_5528,N_3247,N_3846);
nand U5529 (N_5529,N_3666,N_3457);
or U5530 (N_5530,N_3270,N_3554);
nand U5531 (N_5531,N_3472,N_3109);
or U5532 (N_5532,N_4314,N_3099);
nor U5533 (N_5533,N_3263,N_3937);
or U5534 (N_5534,N_3339,N_3871);
or U5535 (N_5535,N_3609,N_3504);
and U5536 (N_5536,N_3668,N_4258);
nor U5537 (N_5537,N_3653,N_3318);
nor U5538 (N_5538,N_3764,N_4141);
or U5539 (N_5539,N_4341,N_4378);
or U5540 (N_5540,N_4142,N_4417);
nor U5541 (N_5541,N_3879,N_4321);
and U5542 (N_5542,N_3492,N_4267);
or U5543 (N_5543,N_3445,N_4287);
or U5544 (N_5544,N_4264,N_3285);
and U5545 (N_5545,N_3623,N_3788);
or U5546 (N_5546,N_3610,N_3913);
nand U5547 (N_5547,N_4116,N_3049);
and U5548 (N_5548,N_3036,N_4356);
and U5549 (N_5549,N_4049,N_3626);
and U5550 (N_5550,N_3620,N_4180);
or U5551 (N_5551,N_3999,N_3959);
and U5552 (N_5552,N_3424,N_3976);
nor U5553 (N_5553,N_3465,N_3913);
or U5554 (N_5554,N_4232,N_3465);
and U5555 (N_5555,N_4037,N_3225);
or U5556 (N_5556,N_3737,N_4410);
nand U5557 (N_5557,N_4338,N_4470);
xor U5558 (N_5558,N_4301,N_3397);
or U5559 (N_5559,N_4380,N_4323);
nor U5560 (N_5560,N_4399,N_4259);
and U5561 (N_5561,N_3788,N_3276);
and U5562 (N_5562,N_3367,N_3615);
or U5563 (N_5563,N_4344,N_3939);
nor U5564 (N_5564,N_3679,N_3794);
and U5565 (N_5565,N_3274,N_3283);
or U5566 (N_5566,N_4412,N_4334);
or U5567 (N_5567,N_3678,N_3200);
nor U5568 (N_5568,N_3150,N_3815);
nor U5569 (N_5569,N_4488,N_3097);
nand U5570 (N_5570,N_3536,N_3023);
or U5571 (N_5571,N_3114,N_3379);
nor U5572 (N_5572,N_3145,N_3459);
and U5573 (N_5573,N_3320,N_4096);
and U5574 (N_5574,N_4391,N_4420);
and U5575 (N_5575,N_3290,N_4423);
or U5576 (N_5576,N_4173,N_4331);
nand U5577 (N_5577,N_4247,N_3868);
and U5578 (N_5578,N_3502,N_3240);
and U5579 (N_5579,N_3689,N_3370);
and U5580 (N_5580,N_3636,N_3506);
or U5581 (N_5581,N_3931,N_4187);
or U5582 (N_5582,N_3147,N_3261);
nand U5583 (N_5583,N_3617,N_3406);
and U5584 (N_5584,N_4438,N_3709);
nor U5585 (N_5585,N_3998,N_3862);
nand U5586 (N_5586,N_3466,N_3188);
nand U5587 (N_5587,N_4032,N_4499);
and U5588 (N_5588,N_3397,N_3429);
or U5589 (N_5589,N_3404,N_3342);
nand U5590 (N_5590,N_3785,N_4364);
and U5591 (N_5591,N_3446,N_3797);
xnor U5592 (N_5592,N_4245,N_3000);
or U5593 (N_5593,N_4042,N_3944);
nand U5594 (N_5594,N_4266,N_3125);
nand U5595 (N_5595,N_4454,N_3819);
or U5596 (N_5596,N_3213,N_3185);
nand U5597 (N_5597,N_4005,N_4385);
xor U5598 (N_5598,N_3362,N_3780);
or U5599 (N_5599,N_3292,N_4391);
and U5600 (N_5600,N_4132,N_4254);
nand U5601 (N_5601,N_4180,N_3374);
and U5602 (N_5602,N_3058,N_3596);
and U5603 (N_5603,N_4077,N_4483);
nor U5604 (N_5604,N_3362,N_3917);
nand U5605 (N_5605,N_3243,N_3757);
or U5606 (N_5606,N_4044,N_4233);
and U5607 (N_5607,N_3864,N_3355);
nor U5608 (N_5608,N_4098,N_3373);
or U5609 (N_5609,N_3162,N_3081);
nand U5610 (N_5610,N_3882,N_4398);
nor U5611 (N_5611,N_3748,N_3459);
nor U5612 (N_5612,N_3414,N_3733);
and U5613 (N_5613,N_4112,N_3534);
or U5614 (N_5614,N_4355,N_3848);
nor U5615 (N_5615,N_3618,N_3991);
or U5616 (N_5616,N_4384,N_3981);
or U5617 (N_5617,N_3168,N_4033);
or U5618 (N_5618,N_3165,N_3257);
nand U5619 (N_5619,N_3329,N_3479);
or U5620 (N_5620,N_3982,N_3310);
nand U5621 (N_5621,N_3894,N_3710);
and U5622 (N_5622,N_4490,N_4168);
or U5623 (N_5623,N_3226,N_4263);
nor U5624 (N_5624,N_3896,N_3684);
nand U5625 (N_5625,N_3703,N_3139);
and U5626 (N_5626,N_3572,N_3078);
nand U5627 (N_5627,N_3337,N_4387);
or U5628 (N_5628,N_3100,N_4211);
nand U5629 (N_5629,N_3768,N_4252);
and U5630 (N_5630,N_3922,N_3936);
or U5631 (N_5631,N_3577,N_3392);
or U5632 (N_5632,N_4113,N_3085);
and U5633 (N_5633,N_3703,N_3233);
and U5634 (N_5634,N_4142,N_3797);
nand U5635 (N_5635,N_4441,N_4373);
or U5636 (N_5636,N_3261,N_4140);
nor U5637 (N_5637,N_4417,N_3602);
or U5638 (N_5638,N_3757,N_3990);
nand U5639 (N_5639,N_3533,N_3328);
or U5640 (N_5640,N_3196,N_4085);
nor U5641 (N_5641,N_3808,N_3480);
nor U5642 (N_5642,N_3945,N_3842);
or U5643 (N_5643,N_3369,N_3700);
or U5644 (N_5644,N_3120,N_4397);
and U5645 (N_5645,N_3041,N_4084);
or U5646 (N_5646,N_4073,N_4324);
and U5647 (N_5647,N_4169,N_3565);
nor U5648 (N_5648,N_3992,N_3168);
nor U5649 (N_5649,N_3333,N_3140);
nand U5650 (N_5650,N_3446,N_3311);
nand U5651 (N_5651,N_3725,N_3642);
and U5652 (N_5652,N_3999,N_4399);
nand U5653 (N_5653,N_3605,N_4463);
nor U5654 (N_5654,N_3235,N_3559);
and U5655 (N_5655,N_4024,N_3118);
nand U5656 (N_5656,N_3068,N_3864);
and U5657 (N_5657,N_3946,N_4296);
nand U5658 (N_5658,N_3933,N_3132);
and U5659 (N_5659,N_3732,N_3317);
and U5660 (N_5660,N_3138,N_3327);
nor U5661 (N_5661,N_3609,N_3390);
and U5662 (N_5662,N_3741,N_4034);
and U5663 (N_5663,N_3472,N_3051);
nand U5664 (N_5664,N_3129,N_3313);
nor U5665 (N_5665,N_3361,N_3251);
xnor U5666 (N_5666,N_3762,N_3155);
and U5667 (N_5667,N_3863,N_3455);
nand U5668 (N_5668,N_3154,N_3702);
nand U5669 (N_5669,N_3262,N_3886);
or U5670 (N_5670,N_3116,N_3664);
or U5671 (N_5671,N_4483,N_3006);
nand U5672 (N_5672,N_3646,N_3509);
and U5673 (N_5673,N_4222,N_3109);
nand U5674 (N_5674,N_3594,N_4036);
or U5675 (N_5675,N_3721,N_4318);
nand U5676 (N_5676,N_4208,N_3447);
or U5677 (N_5677,N_4092,N_3886);
xnor U5678 (N_5678,N_4362,N_3281);
nand U5679 (N_5679,N_3781,N_4221);
nor U5680 (N_5680,N_4068,N_4402);
nor U5681 (N_5681,N_3095,N_3824);
or U5682 (N_5682,N_3291,N_4111);
nand U5683 (N_5683,N_4289,N_4279);
nor U5684 (N_5684,N_3492,N_3023);
or U5685 (N_5685,N_3086,N_3176);
nand U5686 (N_5686,N_3685,N_3631);
nand U5687 (N_5687,N_3350,N_3956);
nor U5688 (N_5688,N_3793,N_4370);
nand U5689 (N_5689,N_3193,N_3592);
or U5690 (N_5690,N_3900,N_3004);
or U5691 (N_5691,N_4268,N_3598);
or U5692 (N_5692,N_4296,N_4348);
nor U5693 (N_5693,N_4422,N_3006);
nor U5694 (N_5694,N_4133,N_3096);
and U5695 (N_5695,N_4233,N_3153);
nor U5696 (N_5696,N_3398,N_3109);
nor U5697 (N_5697,N_4154,N_3360);
nor U5698 (N_5698,N_3584,N_4485);
or U5699 (N_5699,N_3693,N_3357);
or U5700 (N_5700,N_3546,N_4071);
and U5701 (N_5701,N_4262,N_4250);
nand U5702 (N_5702,N_4332,N_3379);
nand U5703 (N_5703,N_4341,N_3433);
nand U5704 (N_5704,N_3676,N_4025);
nand U5705 (N_5705,N_4444,N_4448);
and U5706 (N_5706,N_4162,N_4260);
nand U5707 (N_5707,N_3083,N_4220);
and U5708 (N_5708,N_3791,N_3080);
nand U5709 (N_5709,N_3233,N_4077);
and U5710 (N_5710,N_3792,N_4158);
and U5711 (N_5711,N_4010,N_3314);
nor U5712 (N_5712,N_3138,N_4495);
nand U5713 (N_5713,N_4219,N_4166);
nor U5714 (N_5714,N_3133,N_3930);
or U5715 (N_5715,N_4009,N_4324);
or U5716 (N_5716,N_4291,N_3730);
and U5717 (N_5717,N_3644,N_3707);
or U5718 (N_5718,N_3927,N_4169);
or U5719 (N_5719,N_4300,N_3906);
nand U5720 (N_5720,N_3378,N_4327);
nor U5721 (N_5721,N_3194,N_4326);
nand U5722 (N_5722,N_3354,N_3735);
and U5723 (N_5723,N_3253,N_3387);
xnor U5724 (N_5724,N_3490,N_3756);
nand U5725 (N_5725,N_3807,N_4440);
xor U5726 (N_5726,N_3984,N_4256);
xor U5727 (N_5727,N_4162,N_3788);
nand U5728 (N_5728,N_3114,N_4061);
nor U5729 (N_5729,N_4437,N_3932);
or U5730 (N_5730,N_3353,N_3879);
xor U5731 (N_5731,N_3790,N_3766);
nand U5732 (N_5732,N_3617,N_3818);
nand U5733 (N_5733,N_3171,N_3978);
and U5734 (N_5734,N_3386,N_3778);
nor U5735 (N_5735,N_3111,N_3600);
nor U5736 (N_5736,N_3202,N_4151);
or U5737 (N_5737,N_4177,N_3906);
nand U5738 (N_5738,N_3492,N_4062);
or U5739 (N_5739,N_4490,N_3626);
or U5740 (N_5740,N_3071,N_3750);
and U5741 (N_5741,N_4294,N_4292);
nor U5742 (N_5742,N_4063,N_3213);
and U5743 (N_5743,N_4164,N_3928);
nand U5744 (N_5744,N_3244,N_3848);
or U5745 (N_5745,N_4056,N_4072);
nand U5746 (N_5746,N_3187,N_4016);
or U5747 (N_5747,N_4166,N_3488);
xor U5748 (N_5748,N_3512,N_4065);
nor U5749 (N_5749,N_3003,N_3658);
and U5750 (N_5750,N_3221,N_3749);
nand U5751 (N_5751,N_4408,N_4062);
or U5752 (N_5752,N_3241,N_3204);
and U5753 (N_5753,N_3446,N_3597);
and U5754 (N_5754,N_3903,N_3142);
or U5755 (N_5755,N_3438,N_4373);
nor U5756 (N_5756,N_3629,N_4328);
nand U5757 (N_5757,N_3928,N_3232);
nor U5758 (N_5758,N_4189,N_3680);
or U5759 (N_5759,N_3861,N_3006);
and U5760 (N_5760,N_3064,N_3587);
and U5761 (N_5761,N_3531,N_4466);
and U5762 (N_5762,N_3120,N_4117);
and U5763 (N_5763,N_3541,N_4475);
or U5764 (N_5764,N_4141,N_4499);
nor U5765 (N_5765,N_3937,N_3238);
and U5766 (N_5766,N_3018,N_3632);
and U5767 (N_5767,N_3445,N_3884);
nand U5768 (N_5768,N_4257,N_3841);
nor U5769 (N_5769,N_3415,N_3567);
nor U5770 (N_5770,N_3783,N_4048);
nor U5771 (N_5771,N_3442,N_3864);
nor U5772 (N_5772,N_4478,N_4289);
xor U5773 (N_5773,N_3505,N_4164);
and U5774 (N_5774,N_3965,N_4322);
nor U5775 (N_5775,N_4236,N_3607);
and U5776 (N_5776,N_3417,N_4148);
or U5777 (N_5777,N_3948,N_3534);
nor U5778 (N_5778,N_3410,N_3405);
nand U5779 (N_5779,N_3830,N_3283);
nand U5780 (N_5780,N_4233,N_4055);
nor U5781 (N_5781,N_3702,N_4064);
nor U5782 (N_5782,N_3611,N_3993);
nand U5783 (N_5783,N_3011,N_3920);
or U5784 (N_5784,N_3927,N_3868);
nor U5785 (N_5785,N_3610,N_3343);
and U5786 (N_5786,N_4140,N_4091);
and U5787 (N_5787,N_4353,N_4032);
and U5788 (N_5788,N_3120,N_4009);
or U5789 (N_5789,N_3328,N_3744);
nor U5790 (N_5790,N_3634,N_3783);
nor U5791 (N_5791,N_4283,N_3849);
or U5792 (N_5792,N_4341,N_3860);
nand U5793 (N_5793,N_4159,N_3780);
xnor U5794 (N_5794,N_3263,N_4015);
xnor U5795 (N_5795,N_3360,N_3802);
nor U5796 (N_5796,N_3872,N_3286);
and U5797 (N_5797,N_3958,N_3179);
or U5798 (N_5798,N_3584,N_3915);
nor U5799 (N_5799,N_3109,N_4103);
nor U5800 (N_5800,N_4038,N_3608);
nor U5801 (N_5801,N_4229,N_3657);
nor U5802 (N_5802,N_3936,N_3296);
nand U5803 (N_5803,N_3166,N_4029);
nor U5804 (N_5804,N_3288,N_3372);
nand U5805 (N_5805,N_4423,N_3538);
nor U5806 (N_5806,N_3819,N_3393);
nand U5807 (N_5807,N_3744,N_3121);
and U5808 (N_5808,N_3059,N_3382);
or U5809 (N_5809,N_4493,N_4495);
nor U5810 (N_5810,N_4162,N_3577);
and U5811 (N_5811,N_3021,N_3317);
or U5812 (N_5812,N_3629,N_3156);
and U5813 (N_5813,N_4026,N_3476);
and U5814 (N_5814,N_3061,N_4349);
nand U5815 (N_5815,N_3290,N_3457);
or U5816 (N_5816,N_4073,N_4113);
nor U5817 (N_5817,N_3645,N_3791);
and U5818 (N_5818,N_3350,N_3551);
nor U5819 (N_5819,N_4244,N_4164);
or U5820 (N_5820,N_4461,N_3590);
and U5821 (N_5821,N_3998,N_3753);
or U5822 (N_5822,N_3855,N_4013);
nand U5823 (N_5823,N_3886,N_3062);
or U5824 (N_5824,N_3411,N_3109);
or U5825 (N_5825,N_3075,N_3804);
nand U5826 (N_5826,N_4128,N_3932);
or U5827 (N_5827,N_3595,N_3545);
nand U5828 (N_5828,N_4146,N_4306);
xor U5829 (N_5829,N_4203,N_3472);
and U5830 (N_5830,N_3909,N_4021);
or U5831 (N_5831,N_3963,N_4294);
nor U5832 (N_5832,N_3377,N_3120);
nor U5833 (N_5833,N_4466,N_4029);
or U5834 (N_5834,N_3731,N_3989);
nand U5835 (N_5835,N_3874,N_3153);
nor U5836 (N_5836,N_4264,N_3661);
nor U5837 (N_5837,N_3639,N_3426);
or U5838 (N_5838,N_4474,N_3258);
xor U5839 (N_5839,N_3992,N_3998);
nor U5840 (N_5840,N_3678,N_4195);
or U5841 (N_5841,N_3707,N_3514);
nand U5842 (N_5842,N_3482,N_4051);
or U5843 (N_5843,N_3775,N_4140);
and U5844 (N_5844,N_3979,N_3894);
nand U5845 (N_5845,N_4461,N_3068);
and U5846 (N_5846,N_3854,N_3188);
and U5847 (N_5847,N_3131,N_3333);
and U5848 (N_5848,N_4209,N_3106);
or U5849 (N_5849,N_3689,N_4277);
nor U5850 (N_5850,N_3939,N_4024);
nor U5851 (N_5851,N_3892,N_4370);
nand U5852 (N_5852,N_3901,N_4197);
or U5853 (N_5853,N_3022,N_3360);
and U5854 (N_5854,N_4162,N_3770);
nand U5855 (N_5855,N_4111,N_3044);
or U5856 (N_5856,N_4110,N_3607);
and U5857 (N_5857,N_3455,N_3914);
nor U5858 (N_5858,N_3198,N_3866);
nand U5859 (N_5859,N_4066,N_4477);
and U5860 (N_5860,N_4041,N_3336);
nand U5861 (N_5861,N_3208,N_3512);
and U5862 (N_5862,N_4302,N_4061);
and U5863 (N_5863,N_4119,N_4368);
nand U5864 (N_5864,N_3008,N_3066);
nand U5865 (N_5865,N_4416,N_4414);
and U5866 (N_5866,N_3711,N_3182);
nand U5867 (N_5867,N_3024,N_4120);
or U5868 (N_5868,N_4169,N_3428);
and U5869 (N_5869,N_4480,N_3278);
nand U5870 (N_5870,N_3334,N_3489);
or U5871 (N_5871,N_3350,N_3512);
nor U5872 (N_5872,N_3881,N_4009);
nand U5873 (N_5873,N_3515,N_3050);
and U5874 (N_5874,N_3140,N_3202);
and U5875 (N_5875,N_3688,N_3591);
and U5876 (N_5876,N_4224,N_4052);
nand U5877 (N_5877,N_4066,N_3711);
or U5878 (N_5878,N_3546,N_3587);
nor U5879 (N_5879,N_3315,N_3749);
or U5880 (N_5880,N_4370,N_3278);
nor U5881 (N_5881,N_3373,N_3550);
nand U5882 (N_5882,N_4438,N_3865);
nor U5883 (N_5883,N_3599,N_3665);
nand U5884 (N_5884,N_4236,N_4304);
and U5885 (N_5885,N_3190,N_3135);
nand U5886 (N_5886,N_4494,N_3160);
nand U5887 (N_5887,N_3777,N_3273);
nand U5888 (N_5888,N_3872,N_3427);
nand U5889 (N_5889,N_4330,N_4441);
nor U5890 (N_5890,N_3005,N_3227);
nand U5891 (N_5891,N_3662,N_3040);
nand U5892 (N_5892,N_3442,N_3243);
nand U5893 (N_5893,N_3342,N_3065);
or U5894 (N_5894,N_4064,N_3095);
and U5895 (N_5895,N_3876,N_4227);
nand U5896 (N_5896,N_3938,N_3551);
or U5897 (N_5897,N_4345,N_4378);
nor U5898 (N_5898,N_4313,N_4022);
nor U5899 (N_5899,N_3911,N_4381);
nor U5900 (N_5900,N_3232,N_4357);
and U5901 (N_5901,N_3616,N_4124);
nand U5902 (N_5902,N_3904,N_4200);
and U5903 (N_5903,N_3061,N_4072);
and U5904 (N_5904,N_3368,N_4398);
and U5905 (N_5905,N_3097,N_3372);
and U5906 (N_5906,N_3279,N_4094);
or U5907 (N_5907,N_3843,N_4437);
nand U5908 (N_5908,N_3830,N_4129);
nor U5909 (N_5909,N_3508,N_3004);
and U5910 (N_5910,N_4150,N_4106);
nand U5911 (N_5911,N_4400,N_3926);
or U5912 (N_5912,N_3562,N_3567);
nand U5913 (N_5913,N_3374,N_3242);
or U5914 (N_5914,N_3552,N_3377);
nor U5915 (N_5915,N_3834,N_3589);
nand U5916 (N_5916,N_3809,N_4470);
or U5917 (N_5917,N_3104,N_4099);
nand U5918 (N_5918,N_4062,N_3905);
nand U5919 (N_5919,N_3125,N_3594);
nor U5920 (N_5920,N_3173,N_3315);
nand U5921 (N_5921,N_4275,N_3295);
nor U5922 (N_5922,N_3607,N_3610);
nand U5923 (N_5923,N_3879,N_4145);
and U5924 (N_5924,N_3461,N_3504);
nor U5925 (N_5925,N_3678,N_3941);
or U5926 (N_5926,N_4471,N_3044);
nand U5927 (N_5927,N_4086,N_3343);
and U5928 (N_5928,N_4292,N_4298);
and U5929 (N_5929,N_3992,N_3065);
or U5930 (N_5930,N_3017,N_4324);
nor U5931 (N_5931,N_4109,N_3108);
and U5932 (N_5932,N_4126,N_3116);
nor U5933 (N_5933,N_3138,N_4083);
or U5934 (N_5934,N_3837,N_4020);
nor U5935 (N_5935,N_3999,N_3216);
or U5936 (N_5936,N_3850,N_3008);
nor U5937 (N_5937,N_4124,N_3863);
or U5938 (N_5938,N_4129,N_4488);
or U5939 (N_5939,N_4061,N_3130);
xnor U5940 (N_5940,N_4436,N_3527);
nor U5941 (N_5941,N_4056,N_3041);
and U5942 (N_5942,N_3380,N_4230);
nand U5943 (N_5943,N_3593,N_4494);
and U5944 (N_5944,N_3917,N_3806);
nand U5945 (N_5945,N_3886,N_3531);
nand U5946 (N_5946,N_4403,N_4094);
nand U5947 (N_5947,N_3788,N_4354);
nand U5948 (N_5948,N_3026,N_4139);
and U5949 (N_5949,N_3415,N_3723);
and U5950 (N_5950,N_4376,N_3094);
nor U5951 (N_5951,N_3559,N_3588);
nand U5952 (N_5952,N_4114,N_3717);
and U5953 (N_5953,N_4128,N_4421);
nor U5954 (N_5954,N_4191,N_3541);
and U5955 (N_5955,N_4451,N_3008);
xor U5956 (N_5956,N_4495,N_3861);
nor U5957 (N_5957,N_3346,N_4187);
nand U5958 (N_5958,N_3266,N_4178);
nand U5959 (N_5959,N_4229,N_3400);
nor U5960 (N_5960,N_3872,N_3539);
nor U5961 (N_5961,N_4388,N_3908);
and U5962 (N_5962,N_3497,N_3087);
or U5963 (N_5963,N_4070,N_4264);
nand U5964 (N_5964,N_4450,N_3245);
or U5965 (N_5965,N_3237,N_3063);
nor U5966 (N_5966,N_4467,N_3516);
or U5967 (N_5967,N_4356,N_4426);
and U5968 (N_5968,N_3977,N_3480);
and U5969 (N_5969,N_4029,N_4393);
nand U5970 (N_5970,N_4462,N_3876);
nor U5971 (N_5971,N_3680,N_3493);
and U5972 (N_5972,N_4431,N_4165);
nand U5973 (N_5973,N_3635,N_4293);
nand U5974 (N_5974,N_4037,N_3184);
nand U5975 (N_5975,N_3253,N_3191);
or U5976 (N_5976,N_3040,N_3542);
xor U5977 (N_5977,N_4318,N_3354);
nor U5978 (N_5978,N_3842,N_4409);
xnor U5979 (N_5979,N_3768,N_3311);
nor U5980 (N_5980,N_3413,N_3247);
xnor U5981 (N_5981,N_3235,N_3600);
nand U5982 (N_5982,N_3216,N_4187);
nand U5983 (N_5983,N_3362,N_3573);
nand U5984 (N_5984,N_4279,N_3574);
and U5985 (N_5985,N_3667,N_3081);
nor U5986 (N_5986,N_3901,N_3319);
nor U5987 (N_5987,N_4364,N_3262);
and U5988 (N_5988,N_3435,N_4373);
nor U5989 (N_5989,N_3578,N_4134);
or U5990 (N_5990,N_3133,N_4483);
or U5991 (N_5991,N_3709,N_3524);
nand U5992 (N_5992,N_4424,N_3319);
nor U5993 (N_5993,N_3552,N_3202);
and U5994 (N_5994,N_3796,N_3730);
nor U5995 (N_5995,N_3112,N_3271);
and U5996 (N_5996,N_4391,N_4469);
nand U5997 (N_5997,N_3215,N_3740);
nor U5998 (N_5998,N_4201,N_3833);
nor U5999 (N_5999,N_4310,N_3097);
nand U6000 (N_6000,N_4849,N_4599);
nand U6001 (N_6001,N_5696,N_5365);
nor U6002 (N_6002,N_4559,N_5420);
or U6003 (N_6003,N_5908,N_5688);
nand U6004 (N_6004,N_5863,N_5473);
nor U6005 (N_6005,N_5046,N_5303);
or U6006 (N_6006,N_4706,N_5251);
or U6007 (N_6007,N_5650,N_5555);
or U6008 (N_6008,N_5659,N_4628);
and U6009 (N_6009,N_5063,N_5539);
nor U6010 (N_6010,N_4756,N_5166);
and U6011 (N_6011,N_5865,N_5891);
nand U6012 (N_6012,N_4968,N_5322);
and U6013 (N_6013,N_5220,N_4592);
and U6014 (N_6014,N_4570,N_5866);
nor U6015 (N_6015,N_4778,N_4869);
nand U6016 (N_6016,N_4531,N_4518);
and U6017 (N_6017,N_5733,N_5988);
nor U6018 (N_6018,N_4743,N_5032);
nor U6019 (N_6019,N_4741,N_4703);
nand U6020 (N_6020,N_5557,N_5190);
and U6021 (N_6021,N_5577,N_5961);
nand U6022 (N_6022,N_5771,N_5153);
or U6023 (N_6023,N_4511,N_5631);
and U6024 (N_6024,N_5802,N_5358);
or U6025 (N_6025,N_4950,N_4631);
or U6026 (N_6026,N_5123,N_5242);
nor U6027 (N_6027,N_4597,N_5324);
and U6028 (N_6028,N_4530,N_5091);
or U6029 (N_6029,N_4609,N_5695);
and U6030 (N_6030,N_4677,N_5947);
nor U6031 (N_6031,N_5637,N_5413);
and U6032 (N_6032,N_5878,N_4739);
nor U6033 (N_6033,N_5183,N_4520);
nand U6034 (N_6034,N_5393,N_5478);
nand U6035 (N_6035,N_5277,N_5972);
or U6036 (N_6036,N_4918,N_5974);
nor U6037 (N_6037,N_5664,N_5548);
nand U6038 (N_6038,N_4765,N_5300);
nor U6039 (N_6039,N_5172,N_5169);
nand U6040 (N_6040,N_4845,N_5052);
and U6041 (N_6041,N_5202,N_5390);
and U6042 (N_6042,N_5313,N_4943);
and U6043 (N_6043,N_4789,N_5188);
or U6044 (N_6044,N_4563,N_5389);
or U6045 (N_6045,N_4678,N_5429);
nand U6046 (N_6046,N_5376,N_5682);
or U6047 (N_6047,N_5149,N_5828);
nand U6048 (N_6048,N_5725,N_4864);
or U6049 (N_6049,N_5129,N_4780);
nor U6050 (N_6050,N_5477,N_5714);
nand U6051 (N_6051,N_5775,N_5247);
nand U6052 (N_6052,N_5084,N_5041);
and U6053 (N_6053,N_4745,N_4601);
nor U6054 (N_6054,N_5993,N_5923);
or U6055 (N_6055,N_4852,N_4876);
or U6056 (N_6056,N_4596,N_5273);
and U6057 (N_6057,N_5118,N_5753);
and U6058 (N_6058,N_5261,N_4643);
xnor U6059 (N_6059,N_5464,N_5872);
nand U6060 (N_6060,N_5731,N_5163);
and U6061 (N_6061,N_5575,N_5827);
and U6062 (N_6062,N_5285,N_4565);
and U6063 (N_6063,N_5094,N_4528);
nor U6064 (N_6064,N_4552,N_4836);
nand U6065 (N_6065,N_5338,N_5799);
nor U6066 (N_6066,N_5022,N_5136);
and U6067 (N_6067,N_4718,N_4818);
nand U6068 (N_6068,N_4546,N_5965);
and U6069 (N_6069,N_5004,N_5369);
or U6070 (N_6070,N_4701,N_5435);
nand U6071 (N_6071,N_5919,N_5984);
nand U6072 (N_6072,N_5522,N_5640);
or U6073 (N_6073,N_4670,N_4908);
or U6074 (N_6074,N_5994,N_4660);
nor U6075 (N_6075,N_5050,N_5228);
nor U6076 (N_6076,N_5434,N_5109);
nor U6077 (N_6077,N_5598,N_4867);
or U6078 (N_6078,N_4621,N_4783);
nand U6079 (N_6079,N_5955,N_5959);
xor U6080 (N_6080,N_4988,N_4535);
nor U6081 (N_6081,N_5850,N_4659);
nor U6082 (N_6082,N_5969,N_4506);
xor U6083 (N_6083,N_5068,N_4909);
and U6084 (N_6084,N_5493,N_5895);
nor U6085 (N_6085,N_5877,N_5777);
nor U6086 (N_6086,N_5938,N_5099);
nor U6087 (N_6087,N_4995,N_4692);
nand U6088 (N_6088,N_4676,N_5312);
or U6089 (N_6089,N_4714,N_4771);
nor U6090 (N_6090,N_5170,N_4638);
nand U6091 (N_6091,N_5027,N_5811);
and U6092 (N_6092,N_5119,N_5311);
and U6093 (N_6093,N_4833,N_5465);
or U6094 (N_6094,N_5352,N_5504);
nand U6095 (N_6095,N_5067,N_5034);
and U6096 (N_6096,N_5418,N_5846);
and U6097 (N_6097,N_4913,N_5956);
and U6098 (N_6098,N_5213,N_5713);
and U6099 (N_6099,N_5812,N_5168);
nand U6100 (N_6100,N_5441,N_5658);
nor U6101 (N_6101,N_4607,N_5888);
and U6102 (N_6102,N_5737,N_4807);
and U6103 (N_6103,N_4547,N_5019);
or U6104 (N_6104,N_4564,N_5342);
nand U6105 (N_6105,N_5049,N_4572);
or U6106 (N_6106,N_4610,N_4773);
and U6107 (N_6107,N_4779,N_4814);
nand U6108 (N_6108,N_4812,N_5121);
and U6109 (N_6109,N_4664,N_5954);
and U6110 (N_6110,N_5578,N_5087);
and U6111 (N_6111,N_4951,N_4720);
and U6112 (N_6112,N_5910,N_5419);
nand U6113 (N_6113,N_5964,N_4612);
and U6114 (N_6114,N_5529,N_5256);
nor U6115 (N_6115,N_5932,N_5037);
or U6116 (N_6116,N_5667,N_5968);
or U6117 (N_6117,N_4748,N_4509);
nor U6118 (N_6118,N_5901,N_5134);
or U6119 (N_6119,N_5233,N_4661);
and U6120 (N_6120,N_4777,N_5951);
nor U6121 (N_6121,N_5368,N_5038);
nand U6122 (N_6122,N_5144,N_5699);
nand U6123 (N_6123,N_4666,N_4872);
and U6124 (N_6124,N_5158,N_5662);
nand U6125 (N_6125,N_5054,N_5366);
and U6126 (N_6126,N_5613,N_4976);
xor U6127 (N_6127,N_4573,N_4713);
nand U6128 (N_6128,N_5421,N_5105);
nand U6129 (N_6129,N_5702,N_4768);
nor U6130 (N_6130,N_5933,N_5440);
or U6131 (N_6131,N_5761,N_5056);
and U6132 (N_6132,N_4965,N_4927);
or U6133 (N_6133,N_5388,N_5013);
and U6134 (N_6134,N_4616,N_5830);
nand U6135 (N_6135,N_5375,N_4603);
and U6136 (N_6136,N_5058,N_5395);
nand U6137 (N_6137,N_5849,N_5679);
nor U6138 (N_6138,N_4964,N_5140);
and U6139 (N_6139,N_5654,N_5276);
nand U6140 (N_6140,N_5122,N_5918);
nand U6141 (N_6141,N_5031,N_5454);
nor U6142 (N_6142,N_5357,N_5182);
nand U6143 (N_6143,N_4665,N_5927);
and U6144 (N_6144,N_5622,N_4853);
nor U6145 (N_6145,N_4625,N_4650);
nor U6146 (N_6146,N_4928,N_5683);
or U6147 (N_6147,N_5044,N_4969);
and U6148 (N_6148,N_5779,N_5469);
nand U6149 (N_6149,N_5206,N_5618);
or U6150 (N_6150,N_5344,N_4809);
and U6151 (N_6151,N_5098,N_4878);
nand U6152 (N_6152,N_5047,N_4949);
nor U6153 (N_6153,N_4711,N_5345);
or U6154 (N_6154,N_4758,N_4737);
nand U6155 (N_6155,N_4593,N_4827);
nor U6156 (N_6156,N_4558,N_5936);
nor U6157 (N_6157,N_5139,N_5581);
nor U6158 (N_6158,N_5296,N_5398);
and U6159 (N_6159,N_4545,N_5571);
and U6160 (N_6160,N_4668,N_4887);
or U6161 (N_6161,N_5281,N_5962);
nand U6162 (N_6162,N_5893,N_5298);
nand U6163 (N_6163,N_5000,N_5576);
nand U6164 (N_6164,N_5997,N_5958);
nor U6165 (N_6165,N_4623,N_5001);
nor U6166 (N_6166,N_5948,N_5360);
or U6167 (N_6167,N_4734,N_5826);
xor U6168 (N_6168,N_5708,N_4891);
or U6169 (N_6169,N_5379,N_4899);
xnor U6170 (N_6170,N_4846,N_5354);
nor U6171 (N_6171,N_5619,N_4691);
or U6172 (N_6172,N_5309,N_4514);
or U6173 (N_6173,N_5766,N_4639);
and U6174 (N_6174,N_4751,N_4548);
nor U6175 (N_6175,N_5535,N_5339);
nor U6176 (N_6176,N_5847,N_4742);
nor U6177 (N_6177,N_5490,N_5728);
or U6178 (N_6178,N_5852,N_5361);
and U6179 (N_6179,N_4747,N_5267);
nor U6180 (N_6180,N_5154,N_5781);
nand U6181 (N_6181,N_4662,N_5402);
nand U6182 (N_6182,N_4694,N_5095);
nor U6183 (N_6183,N_5939,N_5743);
xnor U6184 (N_6184,N_5007,N_5861);
nor U6185 (N_6185,N_4679,N_4920);
or U6186 (N_6186,N_4884,N_5999);
and U6187 (N_6187,N_4917,N_5859);
nor U6188 (N_6188,N_5732,N_5758);
or U6189 (N_6189,N_5468,N_5148);
and U6190 (N_6190,N_5211,N_5186);
and U6191 (N_6191,N_4681,N_5727);
and U6192 (N_6192,N_5293,N_5108);
nand U6193 (N_6193,N_4774,N_5840);
or U6194 (N_6194,N_4635,N_5600);
or U6195 (N_6195,N_5567,N_4571);
and U6196 (N_6196,N_4655,N_5515);
nor U6197 (N_6197,N_5081,N_4895);
or U6198 (N_6198,N_4693,N_4823);
and U6199 (N_6199,N_5266,N_5518);
and U6200 (N_6200,N_5334,N_5632);
or U6201 (N_6201,N_5252,N_5350);
and U6202 (N_6202,N_5784,N_5832);
xnor U6203 (N_6203,N_5718,N_5432);
nor U6204 (N_6204,N_4562,N_5330);
nor U6205 (N_6205,N_5125,N_5160);
or U6206 (N_6206,N_5656,N_5075);
xnor U6207 (N_6207,N_5572,N_4697);
or U6208 (N_6208,N_4654,N_4859);
nor U6209 (N_6209,N_5137,N_4804);
or U6210 (N_6210,N_5808,N_5701);
or U6211 (N_6211,N_5981,N_5533);
and U6212 (N_6212,N_5983,N_5184);
and U6213 (N_6213,N_5980,N_4501);
xnor U6214 (N_6214,N_5782,N_5584);
xnor U6215 (N_6215,N_4721,N_4996);
nor U6216 (N_6216,N_5016,N_4508);
nor U6217 (N_6217,N_5989,N_5605);
nor U6218 (N_6218,N_4510,N_4502);
xor U6219 (N_6219,N_4841,N_5762);
nand U6220 (N_6220,N_5255,N_5531);
nor U6221 (N_6221,N_4525,N_4544);
or U6222 (N_6222,N_5258,N_5175);
nor U6223 (N_6223,N_5985,N_5804);
nor U6224 (N_6224,N_5077,N_4642);
nor U6225 (N_6225,N_5355,N_4857);
or U6226 (N_6226,N_5466,N_5425);
nand U6227 (N_6227,N_5043,N_5165);
or U6228 (N_6228,N_4978,N_5614);
and U6229 (N_6229,N_5716,N_4519);
or U6230 (N_6230,N_4822,N_4803);
nand U6231 (N_6231,N_4667,N_5909);
nor U6232 (N_6232,N_5929,N_5249);
nand U6233 (N_6233,N_4802,N_4960);
nor U6234 (N_6234,N_5018,N_5500);
and U6235 (N_6235,N_4794,N_4750);
nor U6236 (N_6236,N_5809,N_5209);
or U6237 (N_6237,N_5672,N_5460);
or U6238 (N_6238,N_5039,N_5689);
or U6239 (N_6239,N_4591,N_5083);
nor U6240 (N_6240,N_5076,N_4837);
or U6241 (N_6241,N_5192,N_5214);
and U6242 (N_6242,N_5411,N_4850);
nor U6243 (N_6243,N_5250,N_4815);
nand U6244 (N_6244,N_5684,N_4940);
nand U6245 (N_6245,N_5457,N_5686);
nor U6246 (N_6246,N_5364,N_5232);
nand U6247 (N_6247,N_5604,N_4790);
nand U6248 (N_6248,N_5196,N_5208);
xnor U6249 (N_6249,N_5596,N_4663);
nor U6250 (N_6250,N_4992,N_5191);
nand U6251 (N_6251,N_5200,N_4839);
and U6252 (N_6252,N_4984,N_5127);
nor U6253 (N_6253,N_4991,N_5528);
nor U6254 (N_6254,N_4730,N_4578);
or U6255 (N_6255,N_5234,N_5815);
and U6256 (N_6256,N_4817,N_4608);
or U6257 (N_6257,N_5957,N_5316);
nor U6258 (N_6258,N_5128,N_4763);
nor U6259 (N_6259,N_4647,N_4675);
and U6260 (N_6260,N_5270,N_4543);
and U6261 (N_6261,N_5800,N_5476);
nor U6262 (N_6262,N_5057,N_5422);
or U6263 (N_6263,N_5289,N_4974);
or U6264 (N_6264,N_4579,N_5795);
nand U6265 (N_6265,N_4819,N_4957);
or U6266 (N_6266,N_5132,N_4848);
xor U6267 (N_6267,N_4998,N_4844);
or U6268 (N_6268,N_4994,N_4652);
nor U6269 (N_6269,N_5253,N_5643);
and U6270 (N_6270,N_5445,N_5433);
nor U6271 (N_6271,N_4522,N_5582);
or U6272 (N_6272,N_4504,N_4952);
and U6273 (N_6273,N_5769,N_5587);
and U6274 (N_6274,N_5294,N_4929);
nand U6275 (N_6275,N_5212,N_5221);
nand U6276 (N_6276,N_4955,N_5855);
nor U6277 (N_6277,N_5374,N_5554);
and U6278 (N_6278,N_5561,N_4914);
or U6279 (N_6279,N_4617,N_5020);
nor U6280 (N_6280,N_5813,N_5331);
nor U6281 (N_6281,N_5979,N_4533);
and U6282 (N_6282,N_5586,N_4605);
nand U6283 (N_6283,N_4566,N_5945);
and U6284 (N_6284,N_4854,N_4633);
or U6285 (N_6285,N_5479,N_5973);
nor U6286 (N_6286,N_4521,N_4981);
nand U6287 (N_6287,N_4970,N_5496);
nor U6288 (N_6288,N_4786,N_4568);
or U6289 (N_6289,N_5491,N_4586);
nor U6290 (N_6290,N_5349,N_5502);
and U6291 (N_6291,N_4507,N_5824);
xnor U6292 (N_6292,N_5215,N_4885);
and U6293 (N_6293,N_5755,N_4934);
nand U6294 (N_6294,N_4557,N_5438);
and U6295 (N_6295,N_5792,N_4813);
nor U6296 (N_6296,N_5097,N_5562);
or U6297 (N_6297,N_5328,N_4658);
nor U6298 (N_6298,N_5135,N_5002);
or U6299 (N_6299,N_5693,N_5765);
nand U6300 (N_6300,N_4785,N_4740);
nor U6301 (N_6301,N_4816,N_5171);
and U6302 (N_6302,N_5065,N_5503);
nor U6303 (N_6303,N_5394,N_5726);
nand U6304 (N_6304,N_5793,N_4759);
and U6305 (N_6305,N_4875,N_5426);
nor U6306 (N_6306,N_5514,N_5543);
nand U6307 (N_6307,N_5382,N_5151);
and U6308 (N_6308,N_4580,N_4641);
nand U6309 (N_6309,N_4792,N_4843);
or U6310 (N_6310,N_5615,N_5715);
and U6311 (N_6311,N_4523,N_5982);
or U6312 (N_6312,N_5078,N_5082);
nand U6313 (N_6313,N_5794,N_4880);
nand U6314 (N_6314,N_4744,N_5963);
nand U6315 (N_6315,N_4584,N_5589);
nand U6316 (N_6316,N_4728,N_5508);
nand U6317 (N_6317,N_4731,N_5120);
nor U6318 (N_6318,N_5788,N_5048);
or U6319 (N_6319,N_5101,N_4726);
nor U6320 (N_6320,N_5308,N_5159);
nand U6321 (N_6321,N_5807,N_4733);
nand U6322 (N_6322,N_5602,N_4683);
nor U6323 (N_6323,N_5942,N_5926);
or U6324 (N_6324,N_5569,N_5621);
or U6325 (N_6325,N_5472,N_5371);
and U6326 (N_6326,N_5524,N_5745);
nand U6327 (N_6327,N_5236,N_5185);
and U6328 (N_6328,N_5690,N_5451);
and U6329 (N_6329,N_5042,N_4987);
nor U6330 (N_6330,N_5279,N_5275);
nor U6331 (N_6331,N_5976,N_5329);
and U6332 (N_6332,N_4907,N_5756);
nand U6333 (N_6333,N_5952,N_5593);
or U6334 (N_6334,N_5486,N_5673);
or U6335 (N_6335,N_4997,N_5990);
nand U6336 (N_6336,N_5162,N_5222);
xor U6337 (N_6337,N_5456,N_5116);
nor U6338 (N_6338,N_5397,N_5879);
nand U6339 (N_6339,N_5623,N_5911);
or U6340 (N_6340,N_5564,N_5953);
nor U6341 (N_6341,N_4611,N_5407);
nand U6342 (N_6342,N_5676,N_5829);
and U6343 (N_6343,N_5302,N_5723);
and U6344 (N_6344,N_4690,N_4515);
or U6345 (N_6345,N_4553,N_4561);
nor U6346 (N_6346,N_5885,N_5288);
and U6347 (N_6347,N_5239,N_4871);
nand U6348 (N_6348,N_5534,N_5437);
and U6349 (N_6349,N_5040,N_5260);
nor U6350 (N_6350,N_4863,N_4700);
and U6351 (N_6351,N_5385,N_5060);
nor U6352 (N_6352,N_5106,N_5157);
and U6353 (N_6353,N_5960,N_5883);
nand U6354 (N_6354,N_5899,N_5317);
and U6355 (N_6355,N_5921,N_5343);
nand U6356 (N_6356,N_5513,N_4873);
nand U6357 (N_6357,N_5017,N_5588);
nor U6358 (N_6358,N_5553,N_5864);
xnor U6359 (N_6359,N_5821,N_5178);
nor U6360 (N_6360,N_4512,N_4999);
nor U6361 (N_6361,N_5680,N_4787);
and U6362 (N_6362,N_5741,N_5203);
and U6363 (N_6363,N_5594,N_5523);
nand U6364 (N_6364,N_5970,N_4725);
or U6365 (N_6365,N_4986,N_5387);
nand U6366 (N_6366,N_5573,N_5340);
and U6367 (N_6367,N_5071,N_5197);
and U6368 (N_6368,N_5341,N_5744);
xnor U6369 (N_6369,N_5946,N_4784);
nor U6370 (N_6370,N_5131,N_4526);
nand U6371 (N_6371,N_4674,N_5112);
nor U6372 (N_6372,N_5995,N_4699);
nand U6373 (N_6373,N_4808,N_5991);
or U6374 (N_6374,N_5996,N_4932);
nor U6375 (N_6375,N_5180,N_5264);
and U6376 (N_6376,N_5532,N_5559);
xor U6377 (N_6377,N_4944,N_4587);
and U6378 (N_6378,N_5896,N_5648);
or U6379 (N_6379,N_5545,N_4961);
nand U6380 (N_6380,N_4979,N_4838);
or U6381 (N_6381,N_5704,N_5494);
nor U6382 (N_6382,N_5754,N_5412);
nor U6383 (N_6383,N_4772,N_5915);
or U6384 (N_6384,N_4904,N_4855);
nor U6385 (N_6385,N_5805,N_5607);
nor U6386 (N_6386,N_5114,N_4629);
nor U6387 (N_6387,N_5912,N_5870);
nor U6388 (N_6388,N_5674,N_5698);
and U6389 (N_6389,N_5843,N_4626);
nand U6390 (N_6390,N_4529,N_5721);
or U6391 (N_6391,N_5336,N_4901);
and U6392 (N_6392,N_5014,N_4735);
nor U6393 (N_6393,N_5367,N_5785);
and U6394 (N_6394,N_5636,N_5563);
or U6395 (N_6395,N_5868,N_5484);
nor U6396 (N_6396,N_5565,N_5776);
or U6397 (N_6397,N_4856,N_5069);
nand U6398 (N_6398,N_4959,N_4912);
or U6399 (N_6399,N_5750,N_5971);
xor U6400 (N_6400,N_4769,N_5625);
nor U6401 (N_6401,N_5644,N_5226);
and U6402 (N_6402,N_5138,N_5579);
nor U6403 (N_6403,N_5304,N_4541);
and U6404 (N_6404,N_5620,N_5797);
and U6405 (N_6405,N_4866,N_4942);
nor U6406 (N_6406,N_4749,N_4933);
or U6407 (N_6407,N_5501,N_5820);
nand U6408 (N_6408,N_5892,N_4554);
or U6409 (N_6409,N_4618,N_5113);
nor U6410 (N_6410,N_5703,N_5488);
nor U6411 (N_6411,N_5405,N_5786);
and U6412 (N_6412,N_4671,N_5416);
and U6413 (N_6413,N_4902,N_5665);
nand U6414 (N_6414,N_5225,N_4761);
nand U6415 (N_6415,N_4835,N_5838);
and U6416 (N_6416,N_5527,N_5663);
nand U6417 (N_6417,N_5949,N_5482);
nor U6418 (N_6418,N_5035,N_4931);
and U6419 (N_6419,N_4595,N_5585);
nor U6420 (N_6420,N_5819,N_4555);
nand U6421 (N_6421,N_5229,N_5126);
nor U6422 (N_6422,N_5759,N_5373);
nor U6423 (N_6423,N_5526,N_5530);
or U6424 (N_6424,N_4972,N_5876);
and U6425 (N_6425,N_5924,N_5380);
nand U6426 (N_6426,N_4600,N_4897);
xor U6427 (N_6427,N_5730,N_5327);
and U6428 (N_6428,N_4954,N_5845);
nor U6429 (N_6429,N_5117,N_4963);
xnor U6430 (N_6430,N_4536,N_4860);
and U6431 (N_6431,N_5006,N_5790);
and U6432 (N_6432,N_4698,N_5150);
nand U6433 (N_6433,N_5757,N_5301);
nand U6434 (N_6434,N_5645,N_4834);
nor U6435 (N_6435,N_5803,N_5124);
nand U6436 (N_6436,N_5992,N_5104);
nand U6437 (N_6437,N_5719,N_4702);
xor U6438 (N_6438,N_5066,N_5931);
nand U6439 (N_6439,N_4695,N_5778);
and U6440 (N_6440,N_5238,N_5337);
nor U6441 (N_6441,N_5740,N_5320);
or U6442 (N_6442,N_4911,N_5363);
and U6443 (N_6443,N_4762,N_4889);
nand U6444 (N_6444,N_5902,N_5459);
nor U6445 (N_6445,N_5487,N_4613);
nand U6446 (N_6446,N_5384,N_4842);
nand U6447 (N_6447,N_5709,N_5635);
or U6448 (N_6448,N_5021,N_5986);
nand U6449 (N_6449,N_5452,N_5710);
or U6450 (N_6450,N_4851,N_5742);
nand U6451 (N_6451,N_5661,N_4729);
nand U6452 (N_6452,N_4684,N_5089);
nand U6453 (N_6453,N_5310,N_4637);
or U6454 (N_6454,N_5568,N_5837);
nor U6455 (N_6455,N_4505,N_4882);
nand U6456 (N_6456,N_5817,N_5318);
nor U6457 (N_6457,N_5152,N_5248);
nor U6458 (N_6458,N_4615,N_5763);
nor U6459 (N_6459,N_5045,N_5096);
and U6460 (N_6460,N_4791,N_5284);
nand U6461 (N_6461,N_5566,N_5107);
and U6462 (N_6462,N_5133,N_5760);
nor U6463 (N_6463,N_5935,N_5711);
and U6464 (N_6464,N_4798,N_5351);
or U6465 (N_6465,N_4537,N_5415);
and U6466 (N_6466,N_5480,N_5485);
nor U6467 (N_6467,N_5519,N_4598);
nor U6468 (N_6468,N_5386,N_4716);
or U6469 (N_6469,N_5218,N_4921);
nor U6470 (N_6470,N_4513,N_5347);
nand U6471 (N_6471,N_5550,N_5599);
and U6472 (N_6472,N_5825,N_5399);
and U6473 (N_6473,N_5198,N_5130);
and U6474 (N_6474,N_5431,N_5102);
nand U6475 (N_6475,N_4644,N_5442);
nand U6476 (N_6476,N_5498,N_4766);
nor U6477 (N_6477,N_4705,N_5254);
xor U6478 (N_6478,N_5404,N_5278);
nor U6479 (N_6479,N_4648,N_5439);
or U6480 (N_6480,N_5205,N_5280);
or U6481 (N_6481,N_4538,N_5903);
nand U6482 (N_6482,N_4636,N_4906);
and U6483 (N_6483,N_5536,N_5008);
nor U6484 (N_6484,N_5629,N_4905);
or U6485 (N_6485,N_5244,N_5889);
nor U6486 (N_6486,N_5207,N_4862);
or U6487 (N_6487,N_5074,N_4982);
nor U6488 (N_6488,N_5542,N_4619);
and U6489 (N_6489,N_5842,N_5257);
nand U6490 (N_6490,N_5174,N_4832);
nand U6491 (N_6491,N_5237,N_4946);
nand U6492 (N_6492,N_5796,N_5103);
and U6493 (N_6493,N_5430,N_5462);
or U6494 (N_6494,N_5219,N_5854);
or U6495 (N_6495,N_5287,N_4622);
nand U6496 (N_6496,N_5230,N_5780);
and U6497 (N_6497,N_4985,N_4646);
nand U6498 (N_6498,N_5646,N_4977);
or U6499 (N_6499,N_5142,N_4673);
and U6500 (N_6500,N_4606,N_5898);
nor U6501 (N_6501,N_4517,N_4567);
and U6502 (N_6502,N_5446,N_5217);
nor U6503 (N_6503,N_4935,N_5179);
nand U6504 (N_6504,N_5381,N_5752);
and U6505 (N_6505,N_5541,N_5647);
or U6506 (N_6506,N_4594,N_5540);
nand U6507 (N_6507,N_4656,N_4799);
or U6508 (N_6508,N_4868,N_5146);
and U6509 (N_6509,N_5141,N_4724);
nand U6510 (N_6510,N_5332,N_5323);
nor U6511 (N_6511,N_5609,N_4503);
xor U6512 (N_6512,N_5511,N_4962);
or U6513 (N_6513,N_5590,N_5499);
or U6514 (N_6514,N_5070,N_4582);
or U6515 (N_6515,N_4956,N_5470);
nor U6516 (N_6516,N_5639,N_5560);
and U6517 (N_6517,N_4993,N_5240);
nor U6518 (N_6518,N_5978,N_5836);
or U6519 (N_6519,N_5720,N_5143);
and U6520 (N_6520,N_5475,N_5290);
nand U6521 (N_6521,N_5286,N_5739);
and U6522 (N_6522,N_5610,N_4886);
nor U6523 (N_6523,N_5033,N_4983);
and U6524 (N_6524,N_4975,N_5269);
nor U6525 (N_6525,N_5977,N_4915);
nor U6526 (N_6526,N_5145,N_5314);
xnor U6527 (N_6527,N_4709,N_5922);
or U6528 (N_6528,N_5930,N_5768);
or U6529 (N_6529,N_5633,N_4624);
nor U6530 (N_6530,N_5423,N_5410);
nand U6531 (N_6531,N_5556,N_4923);
nand U6532 (N_6532,N_4500,N_5920);
nor U6533 (N_6533,N_5080,N_4630);
or U6534 (N_6534,N_4685,N_5950);
and U6535 (N_6535,N_5608,N_5497);
and U6536 (N_6536,N_4569,N_5616);
or U6537 (N_6537,N_5801,N_5092);
nor U6538 (N_6538,N_5875,N_4556);
nor U6539 (N_6539,N_5914,N_5156);
xor U6540 (N_6540,N_4990,N_4589);
nand U6541 (N_6541,N_4903,N_5934);
and U6542 (N_6542,N_4781,N_5862);
and U6543 (N_6543,N_4925,N_5967);
or U6544 (N_6544,N_5634,N_4861);
and U6545 (N_6545,N_5164,N_5770);
and U6546 (N_6546,N_5235,N_5428);
nor U6547 (N_6547,N_4576,N_5841);
nand U6548 (N_6548,N_5641,N_5774);
nor U6549 (N_6549,N_5271,N_5406);
or U6550 (N_6550,N_5583,N_5873);
nand U6551 (N_6551,N_5505,N_4649);
nor U6552 (N_6552,N_5424,N_4881);
nand U6553 (N_6553,N_5735,N_5890);
nand U6554 (N_6554,N_5291,N_5734);
nand U6555 (N_6555,N_4945,N_4532);
or U6556 (N_6556,N_5467,N_5444);
and U6557 (N_6557,N_5816,N_5814);
and U6558 (N_6558,N_4980,N_5155);
and U6559 (N_6559,N_4967,N_5798);
nand U6560 (N_6560,N_5907,N_4840);
and U6561 (N_6561,N_4760,N_5263);
and U6562 (N_6562,N_4825,N_5677);
xor U6563 (N_6563,N_4893,N_4971);
nand U6564 (N_6564,N_4604,N_5652);
nor U6565 (N_6565,N_4755,N_4549);
nand U6566 (N_6566,N_5061,N_5193);
or U6567 (N_6567,N_5917,N_5111);
and U6568 (N_6568,N_4764,N_5245);
nand U6569 (N_6569,N_4797,N_5086);
xnor U6570 (N_6570,N_5724,N_5558);
or U6571 (N_6571,N_5201,N_5326);
and U6572 (N_6572,N_5595,N_4811);
or U6573 (N_6573,N_5005,N_4829);
and U6574 (N_6574,N_5516,N_4746);
nor U6575 (N_6575,N_4948,N_4828);
nor U6576 (N_6576,N_5011,N_5904);
nand U6577 (N_6577,N_5224,N_4651);
nor U6578 (N_6578,N_5746,N_5210);
or U6579 (N_6579,N_4574,N_5940);
nand U6580 (N_6580,N_4588,N_4719);
and U6581 (N_6581,N_4870,N_4686);
or U6582 (N_6582,N_5305,N_4910);
nand U6583 (N_6583,N_5272,N_5705);
and U6584 (N_6584,N_4539,N_5447);
xor U6585 (N_6585,N_5030,N_5881);
nand U6586 (N_6586,N_5292,N_5941);
nor U6587 (N_6587,N_5806,N_5749);
nor U6588 (N_6588,N_4575,N_5570);
and U6589 (N_6589,N_5023,N_5194);
and U6590 (N_6590,N_5887,N_5844);
nand U6591 (N_6591,N_5026,N_5913);
nor U6592 (N_6592,N_5871,N_5823);
nand U6593 (N_6593,N_5666,N_5333);
and U6594 (N_6594,N_4722,N_5880);
or U6595 (N_6595,N_5628,N_5937);
or U6596 (N_6596,N_4645,N_5391);
nand U6597 (N_6597,N_4715,N_5853);
and U6598 (N_6598,N_5449,N_5408);
xor U6599 (N_6599,N_5461,N_5546);
nand U6600 (N_6600,N_5738,N_5717);
or U6601 (N_6601,N_5262,N_4776);
and U6602 (N_6602,N_4653,N_5072);
nor U6603 (N_6603,N_5525,N_5681);
or U6604 (N_6604,N_5736,N_5547);
or U6605 (N_6605,N_5010,N_5818);
and U6606 (N_6606,N_5009,N_4708);
and U6607 (N_6607,N_5858,N_4926);
and U6608 (N_6608,N_5897,N_5362);
nor U6609 (N_6609,N_5706,N_5216);
or U6610 (N_6610,N_5204,N_5268);
or U6611 (N_6611,N_5507,N_5093);
and U6612 (N_6612,N_4551,N_5177);
and U6613 (N_6613,N_4717,N_5998);
xor U6614 (N_6614,N_4939,N_4801);
or U6615 (N_6615,N_4788,N_5851);
xor U6616 (N_6616,N_5024,N_5712);
and U6617 (N_6617,N_5243,N_4736);
nand U6618 (N_6618,N_4682,N_4805);
nor U6619 (N_6619,N_4824,N_4821);
or U6620 (N_6620,N_5521,N_5603);
and U6621 (N_6621,N_5495,N_5685);
or U6622 (N_6622,N_5789,N_5671);
nor U6623 (N_6623,N_5678,N_5670);
and U6624 (N_6624,N_5265,N_5592);
or U6625 (N_6625,N_4775,N_5675);
nor U6626 (N_6626,N_5580,N_5860);
and U6627 (N_6627,N_5544,N_5869);
nand U6628 (N_6628,N_4930,N_4577);
nor U6629 (N_6629,N_5856,N_5414);
nand U6630 (N_6630,N_5471,N_5729);
nor U6631 (N_6631,N_5894,N_5307);
or U6632 (N_6632,N_5181,N_5448);
and U6633 (N_6633,N_4688,N_4896);
or U6634 (N_6634,N_5651,N_4634);
nand U6635 (N_6635,N_4820,N_5783);
nand U6636 (N_6636,N_5687,N_5147);
or U6637 (N_6637,N_4858,N_5085);
nor U6638 (N_6638,N_5517,N_5900);
nand U6639 (N_6639,N_5538,N_4966);
and U6640 (N_6640,N_5700,N_5319);
and U6641 (N_6641,N_5400,N_4534);
and U6642 (N_6642,N_5401,N_4689);
nand U6643 (N_6643,N_4585,N_5348);
nor U6644 (N_6644,N_5624,N_5638);
nand U6645 (N_6645,N_5834,N_5173);
and U6646 (N_6646,N_4770,N_4704);
nand U6647 (N_6647,N_5356,N_5297);
nand U6648 (N_6648,N_5321,N_5916);
and U6649 (N_6649,N_5335,N_5246);
and U6650 (N_6650,N_4865,N_5436);
nand U6651 (N_6651,N_5520,N_5055);
or U6652 (N_6652,N_4894,N_5669);
nand U6653 (N_6653,N_4712,N_4753);
nor U6654 (N_6654,N_5657,N_5591);
nor U6655 (N_6655,N_5747,N_4936);
nor U6656 (N_6656,N_4602,N_5697);
nor U6657 (N_6657,N_5187,N_4560);
nor U6658 (N_6658,N_5295,N_5626);
and U6659 (N_6659,N_5722,N_5325);
and U6660 (N_6660,N_5668,N_4810);
or U6661 (N_6661,N_4958,N_5458);
nor U6662 (N_6662,N_4847,N_5403);
or U6663 (N_6663,N_4924,N_4874);
nor U6664 (N_6664,N_5025,N_5928);
nor U6665 (N_6665,N_4632,N_5100);
and U6666 (N_6666,N_5392,N_4793);
and U6667 (N_6667,N_5692,N_5259);
nor U6668 (N_6668,N_5831,N_5617);
or U6669 (N_6669,N_5537,N_5029);
or U6670 (N_6670,N_5073,N_5906);
and U6671 (N_6671,N_5370,N_5606);
nand U6672 (N_6672,N_5966,N_5611);
and U6673 (N_6673,N_5707,N_4680);
nor U6674 (N_6674,N_4888,N_5767);
and U6675 (N_6675,N_5417,N_5839);
and U6676 (N_6676,N_4540,N_5833);
or U6677 (N_6677,N_5882,N_4516);
and U6678 (N_6678,N_5549,N_5383);
or U6679 (N_6679,N_5810,N_4524);
or U6680 (N_6680,N_5372,N_4581);
or U6681 (N_6681,N_5751,N_5649);
nand U6682 (N_6682,N_4738,N_4800);
and U6683 (N_6683,N_4796,N_4727);
or U6684 (N_6684,N_4627,N_5359);
or U6685 (N_6685,N_5655,N_4542);
and U6686 (N_6686,N_5176,N_5627);
and U6687 (N_6687,N_5653,N_5450);
and U6688 (N_6688,N_5353,N_5378);
and U6689 (N_6689,N_4898,N_5346);
or U6690 (N_6690,N_5088,N_5975);
nand U6691 (N_6691,N_4947,N_5791);
or U6692 (N_6692,N_4614,N_5886);
nand U6693 (N_6693,N_4883,N_5691);
or U6694 (N_6694,N_4754,N_5377);
nor U6695 (N_6695,N_4938,N_4767);
or U6696 (N_6696,N_4922,N_5787);
and U6697 (N_6697,N_5987,N_5161);
and U6698 (N_6698,N_5110,N_5283);
nand U6699 (N_6699,N_5227,N_4640);
or U6700 (N_6700,N_4795,N_4890);
and U6701 (N_6701,N_5905,N_5481);
nor U6702 (N_6702,N_4752,N_5506);
and U6703 (N_6703,N_4669,N_5453);
nand U6704 (N_6704,N_4831,N_4806);
nor U6705 (N_6705,N_5189,N_4973);
and U6706 (N_6706,N_5874,N_5601);
nor U6707 (N_6707,N_5694,N_4696);
nor U6708 (N_6708,N_4723,N_5396);
and U6709 (N_6709,N_4707,N_4710);
nor U6710 (N_6710,N_5167,N_4757);
nor U6711 (N_6711,N_5274,N_4892);
or U6712 (N_6712,N_5015,N_5772);
nand U6713 (N_6713,N_4877,N_5199);
nand U6714 (N_6714,N_4620,N_4672);
nor U6715 (N_6715,N_4989,N_5064);
and U6716 (N_6716,N_5455,N_5642);
or U6717 (N_6717,N_5764,N_5773);
or U6718 (N_6718,N_5492,N_4826);
nor U6719 (N_6719,N_5003,N_4900);
and U6720 (N_6720,N_5463,N_4782);
nand U6721 (N_6721,N_5282,N_4657);
nand U6722 (N_6722,N_5053,N_5483);
nor U6723 (N_6723,N_4879,N_5315);
and U6724 (N_6724,N_4953,N_5051);
nor U6725 (N_6725,N_5231,N_5748);
nand U6726 (N_6726,N_5090,N_5443);
or U6727 (N_6727,N_4937,N_5062);
nor U6728 (N_6728,N_4916,N_5427);
or U6729 (N_6729,N_5489,N_5660);
or U6730 (N_6730,N_5884,N_5552);
nor U6731 (N_6731,N_5512,N_4687);
and U6732 (N_6732,N_4941,N_5195);
and U6733 (N_6733,N_5028,N_5822);
or U6734 (N_6734,N_5857,N_5306);
xor U6735 (N_6735,N_5079,N_5943);
nor U6736 (N_6736,N_5059,N_4590);
or U6737 (N_6737,N_5551,N_5115);
or U6738 (N_6738,N_5944,N_5630);
xor U6739 (N_6739,N_5509,N_5012);
and U6740 (N_6740,N_5597,N_5510);
nor U6741 (N_6741,N_4732,N_4550);
nand U6742 (N_6742,N_4527,N_5474);
nor U6743 (N_6743,N_5867,N_5299);
or U6744 (N_6744,N_5241,N_4583);
nand U6745 (N_6745,N_5612,N_5036);
nor U6746 (N_6746,N_5574,N_5835);
nand U6747 (N_6747,N_4830,N_5848);
or U6748 (N_6748,N_4919,N_5223);
or U6749 (N_6749,N_5925,N_5409);
nand U6750 (N_6750,N_5596,N_4858);
or U6751 (N_6751,N_5752,N_5905);
and U6752 (N_6752,N_5510,N_5243);
and U6753 (N_6753,N_5970,N_4968);
nor U6754 (N_6754,N_5802,N_5336);
and U6755 (N_6755,N_4521,N_4758);
or U6756 (N_6756,N_4723,N_5800);
and U6757 (N_6757,N_5370,N_5016);
xnor U6758 (N_6758,N_5491,N_5723);
nand U6759 (N_6759,N_5515,N_4814);
nor U6760 (N_6760,N_5984,N_4815);
nor U6761 (N_6761,N_5893,N_4838);
and U6762 (N_6762,N_4983,N_4720);
nand U6763 (N_6763,N_5539,N_4931);
and U6764 (N_6764,N_4577,N_4685);
or U6765 (N_6765,N_4540,N_5028);
and U6766 (N_6766,N_5324,N_4800);
nand U6767 (N_6767,N_5828,N_5679);
or U6768 (N_6768,N_5783,N_4608);
or U6769 (N_6769,N_4707,N_4850);
and U6770 (N_6770,N_4937,N_5894);
or U6771 (N_6771,N_5129,N_4766);
or U6772 (N_6772,N_4714,N_5503);
and U6773 (N_6773,N_5558,N_5864);
and U6774 (N_6774,N_5051,N_5674);
or U6775 (N_6775,N_5133,N_4964);
nand U6776 (N_6776,N_5028,N_4785);
nor U6777 (N_6777,N_5104,N_4925);
nand U6778 (N_6778,N_5322,N_4774);
or U6779 (N_6779,N_4855,N_4549);
nor U6780 (N_6780,N_5242,N_5234);
and U6781 (N_6781,N_4758,N_5328);
and U6782 (N_6782,N_5084,N_4922);
and U6783 (N_6783,N_4775,N_5177);
nand U6784 (N_6784,N_5210,N_5168);
or U6785 (N_6785,N_5605,N_4736);
or U6786 (N_6786,N_4889,N_4751);
xnor U6787 (N_6787,N_5809,N_5434);
and U6788 (N_6788,N_5723,N_5896);
nor U6789 (N_6789,N_5451,N_5818);
nor U6790 (N_6790,N_5575,N_5599);
and U6791 (N_6791,N_5269,N_5091);
nor U6792 (N_6792,N_5060,N_5223);
nor U6793 (N_6793,N_4701,N_5478);
or U6794 (N_6794,N_4963,N_5151);
and U6795 (N_6795,N_4721,N_4813);
or U6796 (N_6796,N_5347,N_4569);
or U6797 (N_6797,N_5921,N_5748);
and U6798 (N_6798,N_4923,N_4784);
nor U6799 (N_6799,N_5668,N_4614);
nor U6800 (N_6800,N_4597,N_4615);
and U6801 (N_6801,N_4522,N_4791);
nand U6802 (N_6802,N_4591,N_5792);
or U6803 (N_6803,N_4904,N_5002);
nor U6804 (N_6804,N_5206,N_4677);
or U6805 (N_6805,N_5782,N_5085);
or U6806 (N_6806,N_5643,N_5831);
nor U6807 (N_6807,N_4708,N_5471);
and U6808 (N_6808,N_5844,N_4654);
nand U6809 (N_6809,N_5488,N_5915);
or U6810 (N_6810,N_5112,N_5932);
and U6811 (N_6811,N_4665,N_4746);
or U6812 (N_6812,N_5981,N_5083);
nand U6813 (N_6813,N_5852,N_5572);
nand U6814 (N_6814,N_5692,N_4712);
nor U6815 (N_6815,N_4500,N_4808);
and U6816 (N_6816,N_5847,N_5784);
nor U6817 (N_6817,N_4928,N_4736);
nand U6818 (N_6818,N_5110,N_4638);
xnor U6819 (N_6819,N_4947,N_5492);
nand U6820 (N_6820,N_5374,N_4892);
nand U6821 (N_6821,N_5507,N_5938);
nor U6822 (N_6822,N_4982,N_5598);
nand U6823 (N_6823,N_4756,N_4812);
and U6824 (N_6824,N_4593,N_5605);
nor U6825 (N_6825,N_5994,N_5053);
nor U6826 (N_6826,N_4830,N_4871);
or U6827 (N_6827,N_5816,N_5334);
or U6828 (N_6828,N_4651,N_5362);
or U6829 (N_6829,N_4620,N_5481);
nand U6830 (N_6830,N_4875,N_4918);
and U6831 (N_6831,N_5872,N_5898);
nand U6832 (N_6832,N_5663,N_5846);
nor U6833 (N_6833,N_5781,N_5117);
nand U6834 (N_6834,N_4972,N_4609);
nor U6835 (N_6835,N_4965,N_5227);
and U6836 (N_6836,N_5237,N_5504);
or U6837 (N_6837,N_4786,N_5328);
or U6838 (N_6838,N_5251,N_5331);
nand U6839 (N_6839,N_5717,N_5057);
nor U6840 (N_6840,N_5616,N_5845);
and U6841 (N_6841,N_4923,N_4632);
or U6842 (N_6842,N_4954,N_5616);
nand U6843 (N_6843,N_5887,N_5563);
nand U6844 (N_6844,N_5214,N_5763);
and U6845 (N_6845,N_5971,N_5101);
or U6846 (N_6846,N_5656,N_4921);
nor U6847 (N_6847,N_5705,N_5309);
or U6848 (N_6848,N_5345,N_5903);
and U6849 (N_6849,N_4777,N_5354);
nand U6850 (N_6850,N_5480,N_5260);
nor U6851 (N_6851,N_4843,N_5196);
and U6852 (N_6852,N_5153,N_5774);
and U6853 (N_6853,N_4711,N_5722);
nand U6854 (N_6854,N_5580,N_4752);
and U6855 (N_6855,N_5722,N_4655);
or U6856 (N_6856,N_5806,N_5725);
nor U6857 (N_6857,N_4836,N_5212);
nand U6858 (N_6858,N_5744,N_5050);
nor U6859 (N_6859,N_5844,N_4931);
or U6860 (N_6860,N_5776,N_4588);
and U6861 (N_6861,N_5405,N_5544);
nor U6862 (N_6862,N_4531,N_4868);
and U6863 (N_6863,N_5859,N_5547);
nor U6864 (N_6864,N_5795,N_5765);
or U6865 (N_6865,N_4626,N_5297);
nor U6866 (N_6866,N_5325,N_4547);
nor U6867 (N_6867,N_5583,N_4989);
nor U6868 (N_6868,N_5244,N_5201);
nor U6869 (N_6869,N_5289,N_5974);
and U6870 (N_6870,N_5166,N_4577);
nand U6871 (N_6871,N_5339,N_5338);
nor U6872 (N_6872,N_4914,N_5563);
and U6873 (N_6873,N_5544,N_5698);
nand U6874 (N_6874,N_4507,N_5722);
or U6875 (N_6875,N_5728,N_5578);
or U6876 (N_6876,N_4674,N_5498);
nor U6877 (N_6877,N_5888,N_4582);
nand U6878 (N_6878,N_4833,N_4956);
nor U6879 (N_6879,N_4529,N_4791);
nand U6880 (N_6880,N_4947,N_4915);
or U6881 (N_6881,N_5759,N_5843);
nor U6882 (N_6882,N_4548,N_5520);
nand U6883 (N_6883,N_5141,N_5709);
or U6884 (N_6884,N_5439,N_5720);
nor U6885 (N_6885,N_4582,N_5712);
and U6886 (N_6886,N_5933,N_4816);
or U6887 (N_6887,N_5930,N_4684);
nand U6888 (N_6888,N_4553,N_4708);
nor U6889 (N_6889,N_5636,N_5520);
or U6890 (N_6890,N_5948,N_5547);
nand U6891 (N_6891,N_4588,N_5324);
or U6892 (N_6892,N_4810,N_5007);
and U6893 (N_6893,N_5010,N_5510);
or U6894 (N_6894,N_5788,N_4773);
nand U6895 (N_6895,N_5151,N_4985);
or U6896 (N_6896,N_5768,N_5706);
xor U6897 (N_6897,N_5698,N_5008);
and U6898 (N_6898,N_4622,N_5481);
or U6899 (N_6899,N_4873,N_5362);
and U6900 (N_6900,N_4728,N_5852);
and U6901 (N_6901,N_5712,N_4877);
and U6902 (N_6902,N_5993,N_5418);
or U6903 (N_6903,N_5901,N_5905);
nor U6904 (N_6904,N_5809,N_5959);
and U6905 (N_6905,N_4965,N_4680);
and U6906 (N_6906,N_5688,N_5834);
nor U6907 (N_6907,N_5914,N_4554);
or U6908 (N_6908,N_4652,N_5529);
nand U6909 (N_6909,N_5730,N_5020);
nand U6910 (N_6910,N_4594,N_5864);
or U6911 (N_6911,N_4795,N_5539);
nand U6912 (N_6912,N_4714,N_5609);
and U6913 (N_6913,N_4563,N_5462);
or U6914 (N_6914,N_4934,N_5390);
nand U6915 (N_6915,N_5914,N_5863);
nand U6916 (N_6916,N_5702,N_4991);
or U6917 (N_6917,N_4901,N_4783);
nor U6918 (N_6918,N_4746,N_5968);
and U6919 (N_6919,N_5613,N_5838);
and U6920 (N_6920,N_4710,N_5808);
nand U6921 (N_6921,N_5179,N_4929);
nor U6922 (N_6922,N_5096,N_4700);
or U6923 (N_6923,N_5437,N_5335);
nor U6924 (N_6924,N_5340,N_4904);
nand U6925 (N_6925,N_5419,N_5859);
nand U6926 (N_6926,N_5288,N_4576);
or U6927 (N_6927,N_5150,N_4653);
nor U6928 (N_6928,N_5452,N_4561);
or U6929 (N_6929,N_5260,N_5975);
and U6930 (N_6930,N_5310,N_5116);
nor U6931 (N_6931,N_4898,N_5083);
or U6932 (N_6932,N_5139,N_5797);
nand U6933 (N_6933,N_5727,N_4712);
nor U6934 (N_6934,N_4926,N_5591);
or U6935 (N_6935,N_5893,N_5652);
nor U6936 (N_6936,N_5550,N_5101);
nand U6937 (N_6937,N_4602,N_4800);
xnor U6938 (N_6938,N_4815,N_4855);
nor U6939 (N_6939,N_5302,N_4875);
nor U6940 (N_6940,N_5644,N_5053);
xor U6941 (N_6941,N_5419,N_5275);
nor U6942 (N_6942,N_4735,N_5506);
nand U6943 (N_6943,N_5794,N_5853);
and U6944 (N_6944,N_5924,N_4540);
nor U6945 (N_6945,N_5326,N_5378);
nand U6946 (N_6946,N_5795,N_5280);
nor U6947 (N_6947,N_4898,N_5278);
and U6948 (N_6948,N_5183,N_5579);
nor U6949 (N_6949,N_5115,N_5030);
and U6950 (N_6950,N_5199,N_4562);
or U6951 (N_6951,N_4561,N_5543);
nor U6952 (N_6952,N_5698,N_4658);
nor U6953 (N_6953,N_5880,N_4613);
and U6954 (N_6954,N_5842,N_5520);
nand U6955 (N_6955,N_5679,N_4795);
nor U6956 (N_6956,N_5414,N_5557);
or U6957 (N_6957,N_5648,N_4741);
nor U6958 (N_6958,N_4670,N_4867);
and U6959 (N_6959,N_4594,N_5607);
nand U6960 (N_6960,N_4825,N_5732);
or U6961 (N_6961,N_5788,N_5134);
nand U6962 (N_6962,N_4539,N_4765);
nor U6963 (N_6963,N_5101,N_4861);
nand U6964 (N_6964,N_5997,N_5493);
nand U6965 (N_6965,N_4700,N_4679);
or U6966 (N_6966,N_5099,N_5982);
or U6967 (N_6967,N_4747,N_5291);
or U6968 (N_6968,N_4738,N_5603);
and U6969 (N_6969,N_5401,N_4559);
nand U6970 (N_6970,N_5624,N_5098);
and U6971 (N_6971,N_5974,N_5894);
xnor U6972 (N_6972,N_5504,N_5539);
nand U6973 (N_6973,N_4763,N_5554);
or U6974 (N_6974,N_5539,N_4670);
and U6975 (N_6975,N_5133,N_5089);
and U6976 (N_6976,N_4960,N_4994);
and U6977 (N_6977,N_4659,N_4613);
nand U6978 (N_6978,N_4951,N_5264);
nand U6979 (N_6979,N_4707,N_5916);
or U6980 (N_6980,N_5414,N_5389);
or U6981 (N_6981,N_5184,N_5253);
nand U6982 (N_6982,N_5709,N_5851);
nor U6983 (N_6983,N_4968,N_5083);
and U6984 (N_6984,N_4787,N_5317);
or U6985 (N_6985,N_5046,N_5194);
nor U6986 (N_6986,N_4698,N_5316);
and U6987 (N_6987,N_5965,N_5703);
nand U6988 (N_6988,N_4699,N_4803);
nand U6989 (N_6989,N_4843,N_5691);
and U6990 (N_6990,N_4766,N_4517);
or U6991 (N_6991,N_5564,N_4603);
nor U6992 (N_6992,N_5161,N_5793);
nor U6993 (N_6993,N_5219,N_5022);
and U6994 (N_6994,N_5972,N_5770);
xnor U6995 (N_6995,N_4686,N_5019);
nor U6996 (N_6996,N_5499,N_5266);
nand U6997 (N_6997,N_5488,N_4772);
or U6998 (N_6998,N_4896,N_5614);
nand U6999 (N_6999,N_5107,N_5907);
nor U7000 (N_7000,N_5396,N_5992);
xnor U7001 (N_7001,N_5490,N_4597);
or U7002 (N_7002,N_5965,N_4788);
nor U7003 (N_7003,N_5316,N_4958);
nand U7004 (N_7004,N_4767,N_4978);
or U7005 (N_7005,N_5664,N_4822);
and U7006 (N_7006,N_4782,N_5700);
nor U7007 (N_7007,N_4846,N_5452);
nand U7008 (N_7008,N_5218,N_5458);
and U7009 (N_7009,N_5026,N_5498);
or U7010 (N_7010,N_4648,N_5091);
or U7011 (N_7011,N_5484,N_5549);
nand U7012 (N_7012,N_5553,N_4563);
nor U7013 (N_7013,N_5637,N_4640);
or U7014 (N_7014,N_5027,N_5068);
nand U7015 (N_7015,N_4934,N_5079);
and U7016 (N_7016,N_5830,N_5924);
or U7017 (N_7017,N_5575,N_5348);
and U7018 (N_7018,N_4870,N_5179);
nor U7019 (N_7019,N_4657,N_5189);
nor U7020 (N_7020,N_5338,N_5445);
nand U7021 (N_7021,N_5617,N_5388);
nand U7022 (N_7022,N_4954,N_4600);
and U7023 (N_7023,N_5450,N_4758);
and U7024 (N_7024,N_4593,N_5357);
or U7025 (N_7025,N_4931,N_5590);
nand U7026 (N_7026,N_5671,N_4878);
or U7027 (N_7027,N_4583,N_4884);
nand U7028 (N_7028,N_4707,N_5842);
and U7029 (N_7029,N_5980,N_5247);
nand U7030 (N_7030,N_5127,N_5728);
nand U7031 (N_7031,N_5592,N_5495);
nand U7032 (N_7032,N_5914,N_4946);
and U7033 (N_7033,N_5083,N_5049);
and U7034 (N_7034,N_5563,N_4687);
and U7035 (N_7035,N_4937,N_4530);
nor U7036 (N_7036,N_5157,N_5646);
or U7037 (N_7037,N_5735,N_5496);
and U7038 (N_7038,N_5332,N_4986);
and U7039 (N_7039,N_5818,N_5315);
and U7040 (N_7040,N_5685,N_4838);
or U7041 (N_7041,N_4625,N_4832);
nand U7042 (N_7042,N_4990,N_4843);
or U7043 (N_7043,N_4815,N_5080);
nor U7044 (N_7044,N_4558,N_5374);
nor U7045 (N_7045,N_5214,N_4833);
and U7046 (N_7046,N_4926,N_4578);
nand U7047 (N_7047,N_4924,N_4599);
nand U7048 (N_7048,N_4759,N_4773);
nand U7049 (N_7049,N_5664,N_5987);
or U7050 (N_7050,N_4876,N_5192);
or U7051 (N_7051,N_5980,N_4575);
nand U7052 (N_7052,N_5032,N_4553);
and U7053 (N_7053,N_5315,N_5271);
nand U7054 (N_7054,N_4700,N_5751);
nor U7055 (N_7055,N_5889,N_4791);
or U7056 (N_7056,N_5689,N_5553);
xnor U7057 (N_7057,N_5097,N_5915);
nand U7058 (N_7058,N_5108,N_4505);
nor U7059 (N_7059,N_5042,N_5796);
nor U7060 (N_7060,N_5851,N_5043);
nor U7061 (N_7061,N_5468,N_4716);
nor U7062 (N_7062,N_5887,N_5435);
nand U7063 (N_7063,N_5369,N_5955);
and U7064 (N_7064,N_5859,N_5532);
nor U7065 (N_7065,N_4736,N_4579);
nor U7066 (N_7066,N_5339,N_5490);
or U7067 (N_7067,N_5226,N_4703);
nor U7068 (N_7068,N_5097,N_4931);
nor U7069 (N_7069,N_4867,N_5597);
nor U7070 (N_7070,N_5767,N_5449);
xor U7071 (N_7071,N_5651,N_5431);
or U7072 (N_7072,N_4991,N_4827);
and U7073 (N_7073,N_4986,N_5905);
nand U7074 (N_7074,N_5177,N_5595);
or U7075 (N_7075,N_4927,N_4822);
and U7076 (N_7076,N_5125,N_5672);
or U7077 (N_7077,N_4797,N_4706);
or U7078 (N_7078,N_4918,N_5712);
or U7079 (N_7079,N_5803,N_5710);
nor U7080 (N_7080,N_5240,N_4858);
and U7081 (N_7081,N_5871,N_5511);
nand U7082 (N_7082,N_5798,N_5903);
xor U7083 (N_7083,N_5587,N_5231);
or U7084 (N_7084,N_4721,N_5535);
or U7085 (N_7085,N_5150,N_4975);
and U7086 (N_7086,N_5135,N_5436);
or U7087 (N_7087,N_5558,N_5673);
nor U7088 (N_7088,N_5911,N_4577);
nor U7089 (N_7089,N_5148,N_4705);
nor U7090 (N_7090,N_5201,N_5735);
or U7091 (N_7091,N_5830,N_5450);
or U7092 (N_7092,N_5986,N_5508);
nor U7093 (N_7093,N_5205,N_5717);
nor U7094 (N_7094,N_5614,N_4870);
and U7095 (N_7095,N_5833,N_4505);
and U7096 (N_7096,N_5275,N_5520);
nor U7097 (N_7097,N_4538,N_5634);
nor U7098 (N_7098,N_5408,N_5004);
and U7099 (N_7099,N_5825,N_5492);
nand U7100 (N_7100,N_5945,N_4905);
and U7101 (N_7101,N_5392,N_4656);
nand U7102 (N_7102,N_5452,N_5667);
or U7103 (N_7103,N_5394,N_4698);
and U7104 (N_7104,N_5425,N_4681);
nand U7105 (N_7105,N_5690,N_5684);
nor U7106 (N_7106,N_5679,N_5996);
nor U7107 (N_7107,N_5716,N_5534);
or U7108 (N_7108,N_5703,N_5369);
nand U7109 (N_7109,N_4661,N_5928);
nor U7110 (N_7110,N_5854,N_5338);
and U7111 (N_7111,N_5110,N_5058);
and U7112 (N_7112,N_5402,N_5777);
xor U7113 (N_7113,N_4634,N_4939);
nand U7114 (N_7114,N_5259,N_5188);
nor U7115 (N_7115,N_4628,N_4842);
or U7116 (N_7116,N_4817,N_5944);
nand U7117 (N_7117,N_5096,N_4737);
nand U7118 (N_7118,N_4963,N_5824);
or U7119 (N_7119,N_4927,N_5072);
and U7120 (N_7120,N_5903,N_5256);
nand U7121 (N_7121,N_5265,N_4891);
nand U7122 (N_7122,N_4804,N_5489);
or U7123 (N_7123,N_5586,N_5425);
nor U7124 (N_7124,N_5079,N_4933);
or U7125 (N_7125,N_5478,N_5861);
or U7126 (N_7126,N_5501,N_5270);
nor U7127 (N_7127,N_4604,N_5704);
nor U7128 (N_7128,N_5233,N_4952);
or U7129 (N_7129,N_5709,N_5578);
and U7130 (N_7130,N_4789,N_4749);
xor U7131 (N_7131,N_5960,N_5826);
nor U7132 (N_7132,N_5069,N_4579);
nor U7133 (N_7133,N_4652,N_5151);
nor U7134 (N_7134,N_5275,N_4598);
nand U7135 (N_7135,N_5238,N_4850);
or U7136 (N_7136,N_5421,N_5734);
nand U7137 (N_7137,N_5540,N_4944);
nand U7138 (N_7138,N_4516,N_5808);
and U7139 (N_7139,N_5060,N_5331);
xor U7140 (N_7140,N_5452,N_4529);
nor U7141 (N_7141,N_5355,N_5073);
and U7142 (N_7142,N_4841,N_5786);
or U7143 (N_7143,N_5634,N_5787);
or U7144 (N_7144,N_5767,N_4735);
and U7145 (N_7145,N_5340,N_5138);
nor U7146 (N_7146,N_5240,N_4666);
nor U7147 (N_7147,N_5671,N_5909);
or U7148 (N_7148,N_5703,N_4839);
nand U7149 (N_7149,N_5255,N_5842);
or U7150 (N_7150,N_5417,N_5880);
nand U7151 (N_7151,N_4589,N_4987);
nor U7152 (N_7152,N_5272,N_5453);
and U7153 (N_7153,N_4719,N_5623);
nor U7154 (N_7154,N_5862,N_5922);
or U7155 (N_7155,N_5017,N_4529);
or U7156 (N_7156,N_5462,N_5191);
nor U7157 (N_7157,N_4687,N_4653);
and U7158 (N_7158,N_4800,N_4791);
nand U7159 (N_7159,N_4672,N_4518);
nor U7160 (N_7160,N_5014,N_5148);
and U7161 (N_7161,N_5278,N_5275);
nor U7162 (N_7162,N_5181,N_5066);
nor U7163 (N_7163,N_5469,N_5910);
or U7164 (N_7164,N_4577,N_5979);
nor U7165 (N_7165,N_5825,N_5298);
nand U7166 (N_7166,N_5529,N_5546);
or U7167 (N_7167,N_5849,N_5700);
and U7168 (N_7168,N_5118,N_4548);
nor U7169 (N_7169,N_5654,N_4750);
nand U7170 (N_7170,N_5530,N_4911);
and U7171 (N_7171,N_5195,N_5322);
and U7172 (N_7172,N_4510,N_5134);
or U7173 (N_7173,N_4930,N_5136);
or U7174 (N_7174,N_5677,N_4977);
and U7175 (N_7175,N_5210,N_5980);
and U7176 (N_7176,N_5401,N_5046);
or U7177 (N_7177,N_5445,N_4646);
and U7178 (N_7178,N_5821,N_5561);
or U7179 (N_7179,N_5708,N_5148);
nor U7180 (N_7180,N_5044,N_5312);
and U7181 (N_7181,N_5507,N_4796);
xor U7182 (N_7182,N_5058,N_4645);
nand U7183 (N_7183,N_5991,N_5628);
nand U7184 (N_7184,N_5690,N_5155);
or U7185 (N_7185,N_5696,N_4760);
or U7186 (N_7186,N_4550,N_5701);
nand U7187 (N_7187,N_5671,N_4979);
and U7188 (N_7188,N_4813,N_5976);
nand U7189 (N_7189,N_5172,N_4806);
nor U7190 (N_7190,N_4716,N_5401);
and U7191 (N_7191,N_5433,N_4845);
nand U7192 (N_7192,N_5454,N_5941);
and U7193 (N_7193,N_5183,N_5588);
nand U7194 (N_7194,N_4582,N_5303);
or U7195 (N_7195,N_5634,N_4939);
or U7196 (N_7196,N_4548,N_5089);
and U7197 (N_7197,N_5449,N_5264);
and U7198 (N_7198,N_5361,N_4620);
and U7199 (N_7199,N_5175,N_5317);
nand U7200 (N_7200,N_5730,N_5871);
and U7201 (N_7201,N_4953,N_5429);
or U7202 (N_7202,N_5689,N_5405);
and U7203 (N_7203,N_4624,N_4525);
and U7204 (N_7204,N_5528,N_4735);
nand U7205 (N_7205,N_5130,N_4672);
and U7206 (N_7206,N_4871,N_5998);
nand U7207 (N_7207,N_5192,N_5781);
nor U7208 (N_7208,N_4608,N_5436);
or U7209 (N_7209,N_4604,N_5098);
xor U7210 (N_7210,N_5760,N_4889);
nor U7211 (N_7211,N_5820,N_4801);
and U7212 (N_7212,N_4707,N_5365);
nor U7213 (N_7213,N_5530,N_5734);
nor U7214 (N_7214,N_5611,N_5413);
and U7215 (N_7215,N_4534,N_4974);
nand U7216 (N_7216,N_4637,N_4933);
and U7217 (N_7217,N_5271,N_5623);
nand U7218 (N_7218,N_4816,N_5126);
nand U7219 (N_7219,N_4549,N_5425);
nor U7220 (N_7220,N_5556,N_4602);
nor U7221 (N_7221,N_4700,N_5345);
nor U7222 (N_7222,N_4861,N_4855);
or U7223 (N_7223,N_4780,N_4939);
and U7224 (N_7224,N_5792,N_4569);
and U7225 (N_7225,N_5935,N_4526);
nor U7226 (N_7226,N_5790,N_5936);
nor U7227 (N_7227,N_5362,N_4503);
or U7228 (N_7228,N_5632,N_4879);
nor U7229 (N_7229,N_4828,N_4759);
nor U7230 (N_7230,N_4715,N_4589);
nor U7231 (N_7231,N_5168,N_4825);
nor U7232 (N_7232,N_5904,N_5118);
and U7233 (N_7233,N_5660,N_5966);
and U7234 (N_7234,N_4686,N_4548);
and U7235 (N_7235,N_5056,N_5960);
nand U7236 (N_7236,N_4737,N_5500);
or U7237 (N_7237,N_5569,N_5095);
and U7238 (N_7238,N_5315,N_5932);
nor U7239 (N_7239,N_5049,N_5024);
nor U7240 (N_7240,N_5031,N_4513);
nand U7241 (N_7241,N_4986,N_5250);
nor U7242 (N_7242,N_5274,N_5965);
and U7243 (N_7243,N_5543,N_4884);
and U7244 (N_7244,N_4868,N_5625);
and U7245 (N_7245,N_4672,N_5426);
nor U7246 (N_7246,N_5735,N_5803);
and U7247 (N_7247,N_4892,N_5737);
or U7248 (N_7248,N_4807,N_5567);
nor U7249 (N_7249,N_5107,N_4888);
nand U7250 (N_7250,N_4930,N_4665);
or U7251 (N_7251,N_4923,N_4554);
nor U7252 (N_7252,N_4728,N_5790);
nor U7253 (N_7253,N_4528,N_5075);
xor U7254 (N_7254,N_5017,N_5701);
or U7255 (N_7255,N_5161,N_5860);
xor U7256 (N_7256,N_4857,N_4747);
xor U7257 (N_7257,N_4592,N_4638);
xnor U7258 (N_7258,N_5793,N_5834);
or U7259 (N_7259,N_4576,N_5431);
nor U7260 (N_7260,N_5623,N_5257);
nor U7261 (N_7261,N_4601,N_5847);
nor U7262 (N_7262,N_5785,N_4820);
or U7263 (N_7263,N_5596,N_5125);
nor U7264 (N_7264,N_5076,N_4745);
nand U7265 (N_7265,N_5876,N_4990);
or U7266 (N_7266,N_5117,N_5608);
nor U7267 (N_7267,N_5260,N_4512);
nor U7268 (N_7268,N_4855,N_5233);
or U7269 (N_7269,N_5569,N_5914);
nand U7270 (N_7270,N_5593,N_4708);
or U7271 (N_7271,N_5925,N_4807);
nor U7272 (N_7272,N_4845,N_5064);
or U7273 (N_7273,N_4796,N_5766);
nor U7274 (N_7274,N_4890,N_5165);
nand U7275 (N_7275,N_5140,N_5357);
or U7276 (N_7276,N_5323,N_5079);
or U7277 (N_7277,N_4863,N_5268);
or U7278 (N_7278,N_5629,N_4599);
xor U7279 (N_7279,N_5203,N_5030);
and U7280 (N_7280,N_4512,N_5993);
and U7281 (N_7281,N_5966,N_4602);
nor U7282 (N_7282,N_5530,N_5149);
and U7283 (N_7283,N_4653,N_4742);
nor U7284 (N_7284,N_4926,N_5953);
nand U7285 (N_7285,N_5032,N_5744);
or U7286 (N_7286,N_5063,N_5934);
and U7287 (N_7287,N_5869,N_5204);
nand U7288 (N_7288,N_4702,N_4759);
nor U7289 (N_7289,N_4578,N_5682);
nand U7290 (N_7290,N_5415,N_5174);
nor U7291 (N_7291,N_5226,N_5511);
and U7292 (N_7292,N_5483,N_5237);
or U7293 (N_7293,N_4906,N_4816);
nand U7294 (N_7294,N_4882,N_4983);
or U7295 (N_7295,N_4816,N_5877);
or U7296 (N_7296,N_4865,N_5398);
and U7297 (N_7297,N_5811,N_5702);
nor U7298 (N_7298,N_5696,N_5359);
nand U7299 (N_7299,N_5467,N_5816);
nand U7300 (N_7300,N_5763,N_4954);
or U7301 (N_7301,N_5124,N_5543);
or U7302 (N_7302,N_5365,N_4870);
or U7303 (N_7303,N_5005,N_4749);
or U7304 (N_7304,N_5769,N_5056);
and U7305 (N_7305,N_4699,N_5253);
and U7306 (N_7306,N_4580,N_5480);
nand U7307 (N_7307,N_5420,N_5174);
nor U7308 (N_7308,N_4908,N_5423);
and U7309 (N_7309,N_4614,N_5184);
and U7310 (N_7310,N_4644,N_4824);
or U7311 (N_7311,N_4877,N_4830);
nor U7312 (N_7312,N_5380,N_4833);
nor U7313 (N_7313,N_5758,N_5403);
nor U7314 (N_7314,N_5443,N_5502);
nor U7315 (N_7315,N_4569,N_5316);
or U7316 (N_7316,N_5970,N_5444);
or U7317 (N_7317,N_5718,N_4786);
or U7318 (N_7318,N_5243,N_5879);
nor U7319 (N_7319,N_4714,N_4500);
nor U7320 (N_7320,N_5846,N_5618);
and U7321 (N_7321,N_4631,N_4847);
nor U7322 (N_7322,N_5127,N_5970);
nor U7323 (N_7323,N_5484,N_5008);
nor U7324 (N_7324,N_5218,N_5195);
nor U7325 (N_7325,N_4895,N_5334);
and U7326 (N_7326,N_4779,N_4937);
or U7327 (N_7327,N_5374,N_5880);
or U7328 (N_7328,N_5587,N_4652);
or U7329 (N_7329,N_5094,N_5673);
nand U7330 (N_7330,N_5868,N_4941);
nand U7331 (N_7331,N_5746,N_5466);
or U7332 (N_7332,N_4824,N_5569);
and U7333 (N_7333,N_5118,N_5382);
nand U7334 (N_7334,N_4915,N_5276);
xor U7335 (N_7335,N_5321,N_4999);
or U7336 (N_7336,N_4900,N_4634);
nand U7337 (N_7337,N_4856,N_4804);
and U7338 (N_7338,N_5207,N_4593);
nand U7339 (N_7339,N_5418,N_5340);
or U7340 (N_7340,N_4829,N_4637);
nor U7341 (N_7341,N_4882,N_5206);
or U7342 (N_7342,N_5624,N_5971);
or U7343 (N_7343,N_5381,N_4916);
nand U7344 (N_7344,N_4641,N_4769);
nor U7345 (N_7345,N_5476,N_5629);
or U7346 (N_7346,N_5993,N_5660);
or U7347 (N_7347,N_5648,N_4738);
nand U7348 (N_7348,N_5746,N_4825);
or U7349 (N_7349,N_5568,N_4632);
and U7350 (N_7350,N_5533,N_4629);
or U7351 (N_7351,N_4678,N_4851);
nand U7352 (N_7352,N_5310,N_4543);
xor U7353 (N_7353,N_4769,N_5018);
and U7354 (N_7354,N_5367,N_5561);
nor U7355 (N_7355,N_5983,N_5018);
or U7356 (N_7356,N_4804,N_4565);
or U7357 (N_7357,N_5896,N_5303);
xnor U7358 (N_7358,N_5835,N_5077);
or U7359 (N_7359,N_4719,N_5438);
nand U7360 (N_7360,N_4886,N_5367);
and U7361 (N_7361,N_5048,N_5504);
nand U7362 (N_7362,N_5997,N_4746);
nand U7363 (N_7363,N_5551,N_5365);
nand U7364 (N_7364,N_5934,N_4934);
nand U7365 (N_7365,N_5037,N_4607);
and U7366 (N_7366,N_4837,N_4698);
nor U7367 (N_7367,N_5384,N_5908);
or U7368 (N_7368,N_5388,N_5608);
nand U7369 (N_7369,N_5571,N_5340);
or U7370 (N_7370,N_5088,N_4956);
nor U7371 (N_7371,N_5882,N_5052);
nand U7372 (N_7372,N_4957,N_5520);
nand U7373 (N_7373,N_4702,N_4724);
and U7374 (N_7374,N_4831,N_5593);
or U7375 (N_7375,N_5653,N_5436);
or U7376 (N_7376,N_4985,N_5522);
nor U7377 (N_7377,N_5568,N_5026);
nand U7378 (N_7378,N_5321,N_4974);
nor U7379 (N_7379,N_5575,N_4572);
and U7380 (N_7380,N_4567,N_4873);
or U7381 (N_7381,N_5099,N_5266);
nor U7382 (N_7382,N_5262,N_5184);
or U7383 (N_7383,N_5010,N_4698);
or U7384 (N_7384,N_5607,N_5139);
nor U7385 (N_7385,N_5376,N_5549);
nor U7386 (N_7386,N_5572,N_5118);
nand U7387 (N_7387,N_5602,N_5860);
or U7388 (N_7388,N_5720,N_5890);
and U7389 (N_7389,N_5159,N_4669);
and U7390 (N_7390,N_5339,N_5236);
nor U7391 (N_7391,N_4815,N_5024);
xor U7392 (N_7392,N_5859,N_5704);
or U7393 (N_7393,N_4507,N_5147);
or U7394 (N_7394,N_5180,N_5474);
nand U7395 (N_7395,N_5091,N_5323);
nor U7396 (N_7396,N_4657,N_4801);
or U7397 (N_7397,N_5453,N_5594);
nor U7398 (N_7398,N_5675,N_4990);
nand U7399 (N_7399,N_4620,N_5256);
nand U7400 (N_7400,N_5502,N_4661);
and U7401 (N_7401,N_5074,N_4716);
nand U7402 (N_7402,N_5645,N_5805);
and U7403 (N_7403,N_4625,N_4549);
nor U7404 (N_7404,N_5256,N_5826);
and U7405 (N_7405,N_5302,N_5831);
or U7406 (N_7406,N_5129,N_5108);
or U7407 (N_7407,N_5055,N_5133);
and U7408 (N_7408,N_5890,N_5694);
or U7409 (N_7409,N_4954,N_5376);
nand U7410 (N_7410,N_5571,N_5967);
nor U7411 (N_7411,N_4927,N_5671);
nor U7412 (N_7412,N_4806,N_4702);
nor U7413 (N_7413,N_5212,N_5678);
nand U7414 (N_7414,N_5830,N_4923);
nand U7415 (N_7415,N_5432,N_5159);
or U7416 (N_7416,N_5871,N_5313);
or U7417 (N_7417,N_4827,N_5678);
nand U7418 (N_7418,N_4503,N_5161);
nand U7419 (N_7419,N_5331,N_5110);
nand U7420 (N_7420,N_5787,N_5179);
or U7421 (N_7421,N_5905,N_5156);
nor U7422 (N_7422,N_5411,N_4904);
or U7423 (N_7423,N_4576,N_5063);
nor U7424 (N_7424,N_4751,N_5344);
nand U7425 (N_7425,N_4554,N_5723);
nor U7426 (N_7426,N_5285,N_5831);
nor U7427 (N_7427,N_4652,N_5601);
and U7428 (N_7428,N_4621,N_5062);
nor U7429 (N_7429,N_5314,N_5753);
nand U7430 (N_7430,N_5678,N_5945);
or U7431 (N_7431,N_5837,N_5212);
nand U7432 (N_7432,N_5414,N_4662);
nor U7433 (N_7433,N_5518,N_5136);
or U7434 (N_7434,N_4971,N_4714);
nand U7435 (N_7435,N_5078,N_5571);
nor U7436 (N_7436,N_4958,N_4659);
or U7437 (N_7437,N_5933,N_4758);
nor U7438 (N_7438,N_5711,N_4910);
and U7439 (N_7439,N_4889,N_5590);
nand U7440 (N_7440,N_5979,N_5851);
and U7441 (N_7441,N_5233,N_4878);
and U7442 (N_7442,N_4537,N_4789);
nand U7443 (N_7443,N_5254,N_5972);
nand U7444 (N_7444,N_5052,N_5942);
and U7445 (N_7445,N_5541,N_4590);
nor U7446 (N_7446,N_5317,N_5068);
or U7447 (N_7447,N_5581,N_5738);
or U7448 (N_7448,N_5417,N_5074);
and U7449 (N_7449,N_5097,N_5973);
and U7450 (N_7450,N_5742,N_5662);
and U7451 (N_7451,N_5274,N_4975);
nor U7452 (N_7452,N_5033,N_4928);
or U7453 (N_7453,N_4569,N_4751);
or U7454 (N_7454,N_5607,N_5884);
nand U7455 (N_7455,N_4601,N_4839);
xnor U7456 (N_7456,N_4794,N_5118);
and U7457 (N_7457,N_5589,N_5621);
and U7458 (N_7458,N_5032,N_5587);
nor U7459 (N_7459,N_4808,N_5542);
nand U7460 (N_7460,N_4746,N_5235);
or U7461 (N_7461,N_4879,N_4603);
nor U7462 (N_7462,N_5161,N_5739);
nor U7463 (N_7463,N_4957,N_4770);
nor U7464 (N_7464,N_4745,N_4519);
nor U7465 (N_7465,N_4840,N_5082);
nand U7466 (N_7466,N_5085,N_4734);
and U7467 (N_7467,N_4745,N_4738);
and U7468 (N_7468,N_5993,N_5704);
nor U7469 (N_7469,N_4515,N_5415);
or U7470 (N_7470,N_4525,N_5096);
and U7471 (N_7471,N_5920,N_5466);
and U7472 (N_7472,N_5623,N_4811);
or U7473 (N_7473,N_5438,N_5961);
nor U7474 (N_7474,N_4752,N_4588);
and U7475 (N_7475,N_5559,N_5611);
nand U7476 (N_7476,N_4614,N_4691);
nand U7477 (N_7477,N_4740,N_4752);
or U7478 (N_7478,N_5978,N_4854);
or U7479 (N_7479,N_4822,N_5808);
and U7480 (N_7480,N_4819,N_5792);
nand U7481 (N_7481,N_4788,N_4730);
or U7482 (N_7482,N_4694,N_4779);
or U7483 (N_7483,N_4780,N_5922);
nor U7484 (N_7484,N_4540,N_5728);
or U7485 (N_7485,N_4590,N_5423);
nand U7486 (N_7486,N_5354,N_5336);
and U7487 (N_7487,N_4623,N_4809);
nand U7488 (N_7488,N_4557,N_5054);
and U7489 (N_7489,N_5724,N_5753);
nor U7490 (N_7490,N_5195,N_5957);
or U7491 (N_7491,N_5704,N_5268);
and U7492 (N_7492,N_5251,N_5627);
and U7493 (N_7493,N_5171,N_4529);
and U7494 (N_7494,N_5420,N_4845);
nor U7495 (N_7495,N_4593,N_5548);
nor U7496 (N_7496,N_4714,N_4665);
and U7497 (N_7497,N_5450,N_5854);
or U7498 (N_7498,N_5797,N_5698);
and U7499 (N_7499,N_5920,N_5641);
or U7500 (N_7500,N_7011,N_6899);
and U7501 (N_7501,N_7389,N_6403);
or U7502 (N_7502,N_6630,N_6238);
nand U7503 (N_7503,N_6093,N_7299);
nand U7504 (N_7504,N_7210,N_7426);
and U7505 (N_7505,N_6404,N_6506);
nand U7506 (N_7506,N_7310,N_6074);
and U7507 (N_7507,N_6741,N_6863);
nor U7508 (N_7508,N_7280,N_6384);
or U7509 (N_7509,N_7209,N_6826);
nor U7510 (N_7510,N_6964,N_7436);
nor U7511 (N_7511,N_7019,N_6066);
nand U7512 (N_7512,N_7242,N_6619);
nor U7513 (N_7513,N_6381,N_6905);
nor U7514 (N_7514,N_6646,N_6064);
and U7515 (N_7515,N_7112,N_6200);
or U7516 (N_7516,N_6819,N_7109);
nand U7517 (N_7517,N_6166,N_7415);
nor U7518 (N_7518,N_6120,N_7330);
and U7519 (N_7519,N_7337,N_6022);
and U7520 (N_7520,N_6608,N_7043);
nor U7521 (N_7521,N_6903,N_6694);
nand U7522 (N_7522,N_6040,N_6125);
nor U7523 (N_7523,N_6735,N_7143);
nor U7524 (N_7524,N_6462,N_7049);
nand U7525 (N_7525,N_6188,N_7339);
nor U7526 (N_7526,N_6544,N_6292);
and U7527 (N_7527,N_6456,N_6326);
and U7528 (N_7528,N_6033,N_7003);
or U7529 (N_7529,N_6647,N_6334);
or U7530 (N_7530,N_6807,N_7156);
or U7531 (N_7531,N_6138,N_6657);
and U7532 (N_7532,N_6717,N_7127);
and U7533 (N_7533,N_6164,N_6416);
and U7534 (N_7534,N_6050,N_6568);
xor U7535 (N_7535,N_7317,N_6285);
nand U7536 (N_7536,N_6284,N_6765);
or U7537 (N_7537,N_7223,N_7478);
and U7538 (N_7538,N_7321,N_7148);
nor U7539 (N_7539,N_7167,N_6140);
nand U7540 (N_7540,N_6180,N_7084);
nand U7541 (N_7541,N_6096,N_6108);
nor U7542 (N_7542,N_6952,N_6419);
nand U7543 (N_7543,N_6283,N_7336);
and U7544 (N_7544,N_6759,N_6049);
and U7545 (N_7545,N_6303,N_6435);
nor U7546 (N_7546,N_6366,N_6895);
or U7547 (N_7547,N_7149,N_6159);
nand U7548 (N_7548,N_6039,N_6565);
and U7549 (N_7549,N_6612,N_6222);
nand U7550 (N_7550,N_6913,N_6989);
and U7551 (N_7551,N_6362,N_7166);
nand U7552 (N_7552,N_7183,N_6012);
or U7553 (N_7553,N_7273,N_7423);
and U7554 (N_7554,N_7191,N_7081);
nand U7555 (N_7555,N_6958,N_6978);
nor U7556 (N_7556,N_6850,N_6882);
and U7557 (N_7557,N_7364,N_6331);
and U7558 (N_7558,N_6136,N_7298);
or U7559 (N_7559,N_6249,N_7018);
or U7560 (N_7560,N_6473,N_7147);
nand U7561 (N_7561,N_6153,N_7390);
and U7562 (N_7562,N_6686,N_6708);
or U7563 (N_7563,N_6367,N_6428);
and U7564 (N_7564,N_7160,N_6814);
and U7565 (N_7565,N_6221,N_6339);
and U7566 (N_7566,N_6982,N_6868);
or U7567 (N_7567,N_6747,N_7383);
or U7568 (N_7568,N_7228,N_6811);
nor U7569 (N_7569,N_6205,N_6310);
nor U7570 (N_7570,N_7353,N_6547);
or U7571 (N_7571,N_6231,N_6349);
and U7572 (N_7572,N_7044,N_7474);
or U7573 (N_7573,N_7134,N_6282);
nor U7574 (N_7574,N_7168,N_7224);
xnor U7575 (N_7575,N_6970,N_6554);
and U7576 (N_7576,N_6699,N_6206);
or U7577 (N_7577,N_7301,N_7494);
or U7578 (N_7578,N_7370,N_7468);
nand U7579 (N_7579,N_6635,N_6208);
nand U7580 (N_7580,N_6347,N_7486);
or U7581 (N_7581,N_6896,N_6689);
nor U7582 (N_7582,N_6408,N_6385);
nor U7583 (N_7583,N_7063,N_6395);
and U7584 (N_7584,N_6135,N_7358);
and U7585 (N_7585,N_6571,N_6492);
nor U7586 (N_7586,N_7200,N_6682);
or U7587 (N_7587,N_6969,N_7296);
nor U7588 (N_7588,N_6626,N_6676);
and U7589 (N_7589,N_6329,N_6348);
nand U7590 (N_7590,N_6019,N_7028);
nand U7591 (N_7591,N_6241,N_6578);
or U7592 (N_7592,N_6115,N_6237);
nand U7593 (N_7593,N_6388,N_6976);
or U7594 (N_7594,N_6059,N_6352);
nand U7595 (N_7595,N_6902,N_7135);
nand U7596 (N_7596,N_6225,N_7379);
nor U7597 (N_7597,N_6307,N_6121);
nor U7598 (N_7598,N_7195,N_6530);
and U7599 (N_7599,N_6667,N_6800);
nand U7600 (N_7600,N_7214,N_7110);
nand U7601 (N_7601,N_7289,N_6762);
and U7602 (N_7602,N_6269,N_7244);
nand U7603 (N_7603,N_6965,N_6170);
nand U7604 (N_7604,N_6939,N_6534);
nand U7605 (N_7605,N_7247,N_7107);
nand U7606 (N_7606,N_6393,N_6112);
nand U7607 (N_7607,N_6559,N_6212);
nor U7608 (N_7608,N_6668,N_6770);
nand U7609 (N_7609,N_7085,N_6184);
nor U7610 (N_7610,N_6058,N_6055);
nand U7611 (N_7611,N_7307,N_7026);
nor U7612 (N_7612,N_6321,N_6157);
or U7613 (N_7613,N_6070,N_6109);
nor U7614 (N_7614,N_7188,N_7464);
and U7615 (N_7615,N_7329,N_7231);
nand U7616 (N_7616,N_7420,N_7089);
nand U7617 (N_7617,N_6802,N_6972);
nor U7618 (N_7618,N_7221,N_6088);
nand U7619 (N_7619,N_6204,N_7295);
or U7620 (N_7620,N_6207,N_6161);
nand U7621 (N_7621,N_6609,N_6673);
xor U7622 (N_7622,N_6061,N_6234);
and U7623 (N_7623,N_7216,N_6971);
nand U7624 (N_7624,N_7281,N_6721);
nand U7625 (N_7625,N_6894,N_7311);
or U7626 (N_7626,N_6185,N_7103);
and U7627 (N_7627,N_6029,N_7461);
and U7628 (N_7628,N_6703,N_7344);
and U7629 (N_7629,N_6740,N_6364);
or U7630 (N_7630,N_7090,N_6401);
nor U7631 (N_7631,N_6943,N_6444);
nand U7632 (N_7632,N_7233,N_6974);
nand U7633 (N_7633,N_6585,N_7171);
nor U7634 (N_7634,N_6091,N_6431);
nor U7635 (N_7635,N_7190,N_6529);
or U7636 (N_7636,N_7159,N_7041);
or U7637 (N_7637,N_6084,N_6134);
or U7638 (N_7638,N_7249,N_6515);
or U7639 (N_7639,N_6177,N_7498);
nor U7640 (N_7640,N_6178,N_6528);
nor U7641 (N_7641,N_7125,N_7055);
and U7642 (N_7642,N_6202,N_6195);
nand U7643 (N_7643,N_7454,N_7154);
nand U7644 (N_7644,N_7095,N_6675);
and U7645 (N_7645,N_6817,N_7239);
nand U7646 (N_7646,N_6541,N_7456);
or U7647 (N_7647,N_6598,N_7386);
and U7648 (N_7648,N_7203,N_6302);
and U7649 (N_7649,N_7172,N_7179);
nand U7650 (N_7650,N_7104,N_6575);
and U7651 (N_7651,N_7335,N_6360);
or U7652 (N_7652,N_6550,N_7056);
nor U7653 (N_7653,N_6869,N_7004);
nor U7654 (N_7654,N_6254,N_6591);
nand U7655 (N_7655,N_6753,N_7162);
nor U7656 (N_7656,N_6097,N_6083);
or U7657 (N_7657,N_7328,N_6704);
nand U7658 (N_7658,N_7388,N_6773);
nor U7659 (N_7659,N_6354,N_6546);
and U7660 (N_7660,N_6137,N_7485);
nor U7661 (N_7661,N_6918,N_6931);
nand U7662 (N_7662,N_6616,N_6990);
and U7663 (N_7663,N_7073,N_6955);
nand U7664 (N_7664,N_6464,N_6825);
and U7665 (N_7665,N_6552,N_6638);
or U7666 (N_7666,N_6828,N_6163);
nand U7667 (N_7667,N_6469,N_7067);
and U7668 (N_7668,N_7009,N_6183);
and U7669 (N_7669,N_6507,N_6294);
nor U7670 (N_7670,N_6458,N_6436);
nand U7671 (N_7671,N_6176,N_6441);
and U7672 (N_7672,N_7293,N_6235);
and U7673 (N_7673,N_6984,N_6004);
nor U7674 (N_7674,N_6684,N_6094);
nor U7675 (N_7675,N_6917,N_6837);
or U7676 (N_7676,N_6308,N_6579);
and U7677 (N_7677,N_7031,N_6291);
nor U7678 (N_7678,N_6930,N_7215);
nand U7679 (N_7679,N_7375,N_7439);
or U7680 (N_7680,N_6526,N_6259);
and U7681 (N_7681,N_6804,N_6831);
nor U7682 (N_7682,N_6181,N_7139);
nor U7683 (N_7683,N_6472,N_6119);
nor U7684 (N_7684,N_6037,N_7097);
and U7685 (N_7685,N_6196,N_7106);
nor U7686 (N_7686,N_6025,N_7177);
or U7687 (N_7687,N_6588,N_7080);
nand U7688 (N_7688,N_6509,N_6981);
xor U7689 (N_7689,N_6962,N_6244);
xnor U7690 (N_7690,N_6365,N_6967);
nor U7691 (N_7691,N_6483,N_7380);
nor U7692 (N_7692,N_6147,N_6764);
nor U7693 (N_7693,N_6489,N_6398);
and U7694 (N_7694,N_7155,N_6468);
nor U7695 (N_7695,N_6286,N_6928);
nor U7696 (N_7696,N_7122,N_6169);
nand U7697 (N_7697,N_6780,N_6624);
nand U7698 (N_7698,N_6320,N_6324);
and U7699 (N_7699,N_6340,N_6690);
nand U7700 (N_7700,N_6938,N_7238);
xnor U7701 (N_7701,N_6323,N_7445);
or U7702 (N_7702,N_7037,N_6306);
and U7703 (N_7703,N_7213,N_7045);
nor U7704 (N_7704,N_7184,N_7120);
or U7705 (N_7705,N_7432,N_7240);
nor U7706 (N_7706,N_7258,N_6520);
or U7707 (N_7707,N_7479,N_6841);
nand U7708 (N_7708,N_6343,N_7441);
xnor U7709 (N_7709,N_6809,N_6046);
nor U7710 (N_7710,N_7354,N_6570);
and U7711 (N_7711,N_6957,N_6688);
or U7712 (N_7712,N_6650,N_6038);
nand U7713 (N_7713,N_7022,N_7150);
nor U7714 (N_7714,N_6143,N_6835);
nand U7715 (N_7715,N_6081,N_6229);
nor U7716 (N_7716,N_6449,N_6236);
nor U7717 (N_7717,N_7256,N_7181);
nand U7718 (N_7718,N_6071,N_6144);
nand U7719 (N_7719,N_7250,N_6482);
or U7720 (N_7720,N_6775,N_6133);
xor U7721 (N_7721,N_6999,N_6662);
and U7722 (N_7722,N_6274,N_6830);
or U7723 (N_7723,N_6445,N_6386);
nand U7724 (N_7724,N_6150,N_6726);
xnor U7725 (N_7725,N_7092,N_7382);
nand U7726 (N_7726,N_6884,N_6715);
and U7727 (N_7727,N_6087,N_6854);
or U7728 (N_7728,N_6461,N_7254);
nand U7729 (N_7729,N_6371,N_6574);
and U7730 (N_7730,N_6281,N_6333);
and U7731 (N_7731,N_6782,N_7023);
and U7732 (N_7732,N_6769,N_6062);
and U7733 (N_7733,N_6027,N_7477);
or U7734 (N_7734,N_6750,N_7248);
or U7735 (N_7735,N_6211,N_6977);
and U7736 (N_7736,N_6808,N_7381);
or U7737 (N_7737,N_6466,N_7008);
or U7738 (N_7738,N_7169,N_6023);
nor U7739 (N_7739,N_6068,N_6516);
and U7740 (N_7740,N_6090,N_6165);
nor U7741 (N_7741,N_6132,N_7284);
or U7742 (N_7742,N_7323,N_7393);
nor U7743 (N_7743,N_6653,N_6251);
and U7744 (N_7744,N_6746,N_6590);
and U7745 (N_7745,N_6774,N_7163);
nor U7746 (N_7746,N_6906,N_6866);
nor U7747 (N_7747,N_6197,N_6243);
and U7748 (N_7748,N_6532,N_7099);
nand U7749 (N_7749,N_6815,N_7218);
and U7750 (N_7750,N_6611,N_6128);
nand U7751 (N_7751,N_7356,N_6172);
nor U7752 (N_7752,N_6123,N_7411);
or U7753 (N_7753,N_7185,N_6605);
and U7754 (N_7754,N_6649,N_6543);
or U7755 (N_7755,N_6031,N_7002);
or U7756 (N_7756,N_7421,N_6380);
or U7757 (N_7757,N_6793,N_6829);
or U7758 (N_7758,N_7053,N_6947);
and U7759 (N_7759,N_7006,N_6217);
or U7760 (N_7760,N_6305,N_6402);
and U7761 (N_7761,N_6003,N_6853);
or U7762 (N_7762,N_6660,N_7476);
and U7763 (N_7763,N_7487,N_7027);
or U7764 (N_7764,N_6790,N_6680);
xor U7765 (N_7765,N_6495,N_6685);
nor U7766 (N_7766,N_7189,N_6505);
nor U7767 (N_7767,N_7433,N_6414);
or U7768 (N_7768,N_6954,N_6337);
or U7769 (N_7769,N_6430,N_7373);
nor U7770 (N_7770,N_7040,N_7268);
xnor U7771 (N_7771,N_7227,N_7402);
xnor U7772 (N_7772,N_7391,N_7394);
nand U7773 (N_7773,N_6420,N_7261);
or U7774 (N_7774,N_6390,N_6997);
nor U7775 (N_7775,N_7271,N_6335);
and U7776 (N_7776,N_7352,N_7131);
nand U7777 (N_7777,N_7338,N_6034);
and U7778 (N_7778,N_7392,N_6168);
nand U7779 (N_7779,N_7157,N_6415);
nand U7780 (N_7780,N_6114,N_7235);
xnor U7781 (N_7781,N_6020,N_7052);
or U7782 (N_7782,N_6261,N_7208);
nor U7783 (N_7783,N_6493,N_6102);
or U7784 (N_7784,N_7133,N_6763);
xor U7785 (N_7785,N_6862,N_6179);
and U7786 (N_7786,N_6533,N_6936);
and U7787 (N_7787,N_6149,N_7292);
nand U7788 (N_7788,N_6018,N_6299);
or U7789 (N_7789,N_7276,N_7098);
nand U7790 (N_7790,N_6915,N_6073);
and U7791 (N_7791,N_6054,N_7061);
xor U7792 (N_7792,N_6563,N_7158);
nand U7793 (N_7793,N_6599,N_6739);
and U7794 (N_7794,N_6410,N_6778);
or U7795 (N_7795,N_6433,N_6309);
and U7796 (N_7796,N_6785,N_6139);
nand U7797 (N_7797,N_6514,N_6490);
nand U7798 (N_7798,N_6870,N_6459);
and U7799 (N_7799,N_6949,N_7257);
nand U7800 (N_7800,N_7400,N_7059);
and U7801 (N_7801,N_7038,N_6889);
nor U7802 (N_7802,N_6476,N_7422);
nand U7803 (N_7803,N_6110,N_6890);
and U7804 (N_7804,N_7174,N_6101);
and U7805 (N_7805,N_7079,N_6501);
nor U7806 (N_7806,N_7032,N_6572);
nand U7807 (N_7807,N_7197,N_6524);
or U7808 (N_7808,N_7277,N_7260);
and U7809 (N_7809,N_6754,N_6396);
nor U7810 (N_7810,N_6883,N_6898);
and U7811 (N_7811,N_7326,N_6344);
nor U7812 (N_7812,N_6838,N_6710);
and U7813 (N_7813,N_6481,N_6583);
nor U7814 (N_7814,N_6615,N_7121);
and U7815 (N_7815,N_6988,N_7320);
or U7816 (N_7816,N_7291,N_6142);
nand U7817 (N_7817,N_6963,N_6713);
nand U7818 (N_7818,N_6701,N_6443);
nor U7819 (N_7819,N_6538,N_6028);
nand U7820 (N_7820,N_6692,N_6712);
and U7821 (N_7821,N_6056,N_7105);
nor U7822 (N_7822,N_7452,N_7449);
or U7823 (N_7823,N_6772,N_6678);
and U7824 (N_7824,N_7444,N_6214);
nor U7825 (N_7825,N_6045,N_6914);
nand U7826 (N_7826,N_6698,N_6993);
nand U7827 (N_7827,N_6151,N_6080);
or U7828 (N_7828,N_6322,N_6983);
and U7829 (N_7829,N_6296,N_6842);
nor U7830 (N_7830,N_6935,N_6655);
and U7831 (N_7831,N_6907,N_7302);
and U7832 (N_7832,N_6758,N_7137);
nor U7833 (N_7833,N_6358,N_6287);
or U7834 (N_7834,N_7165,N_6519);
nand U7835 (N_7835,N_6266,N_6175);
or U7836 (N_7836,N_7451,N_7252);
or U7837 (N_7837,N_6210,N_6318);
and U7838 (N_7838,N_6173,N_6904);
nand U7839 (N_7839,N_6162,N_6932);
and U7840 (N_7840,N_7453,N_6779);
nor U7841 (N_7841,N_6876,N_6409);
or U7842 (N_7842,N_6986,N_6794);
and U7843 (N_7843,N_6942,N_6720);
and U7844 (N_7844,N_6154,N_7232);
nor U7845 (N_7845,N_7132,N_7404);
or U7846 (N_7846,N_6397,N_6399);
nor U7847 (N_7847,N_6560,N_7230);
or U7848 (N_7848,N_7237,N_6558);
or U7849 (N_7849,N_6130,N_6766);
nor U7850 (N_7850,N_6671,N_6540);
or U7851 (N_7851,N_6451,N_7030);
and U7852 (N_7852,N_6191,N_6155);
nor U7853 (N_7853,N_6706,N_6992);
nor U7854 (N_7854,N_7303,N_6711);
nand U7855 (N_7855,N_7115,N_7078);
or U7856 (N_7856,N_7412,N_6851);
nor U7857 (N_7857,N_6363,N_6350);
nor U7858 (N_7858,N_6141,N_6312);
nor U7859 (N_7859,N_7316,N_7319);
or U7860 (N_7860,N_6002,N_7014);
nor U7861 (N_7861,N_7499,N_6586);
and U7862 (N_7862,N_6219,N_6319);
nor U7863 (N_7863,N_6304,N_6536);
and U7864 (N_7864,N_6961,N_6351);
nand U7865 (N_7865,N_7142,N_6453);
nor U7866 (N_7866,N_6593,N_7243);
and U7867 (N_7867,N_7241,N_6761);
or U7868 (N_7868,N_7251,N_7192);
or U7869 (N_7869,N_6691,N_7202);
nor U7870 (N_7870,N_6672,N_6767);
nand U7871 (N_7871,N_6317,N_6233);
and U7872 (N_7872,N_6374,N_6457);
and U7873 (N_7873,N_6878,N_7126);
xor U7874 (N_7874,N_7117,N_7017);
nor U7875 (N_7875,N_6788,N_6199);
nand U7876 (N_7876,N_6665,N_6255);
nor U7877 (N_7877,N_6338,N_7385);
and U7878 (N_7878,N_7417,N_6875);
and U7879 (N_7879,N_7425,N_6623);
or U7880 (N_7880,N_6921,N_6893);
and U7881 (N_7881,N_6953,N_6258);
nand U7882 (N_7882,N_7459,N_6478);
nor U7883 (N_7883,N_7124,N_6987);
or U7884 (N_7884,N_7489,N_7398);
nor U7885 (N_7885,N_6497,N_6724);
or U7886 (N_7886,N_6827,N_7482);
or U7887 (N_7887,N_6268,N_7480);
nand U7888 (N_7888,N_6858,N_6683);
and U7889 (N_7889,N_6485,N_6355);
nor U7890 (N_7890,N_6107,N_7367);
and U7891 (N_7891,N_6744,N_6816);
nand U7892 (N_7892,N_6645,N_6230);
or U7893 (N_7893,N_7318,N_6263);
and U7894 (N_7894,N_6146,N_7345);
xor U7895 (N_7895,N_6542,N_6127);
and U7896 (N_7896,N_7333,N_7282);
or U7897 (N_7897,N_7334,N_7229);
and U7898 (N_7898,N_6877,N_7173);
or U7899 (N_7899,N_7259,N_7151);
nor U7900 (N_7900,N_6228,N_7493);
nor U7901 (N_7901,N_6298,N_7051);
nand U7902 (N_7902,N_6418,N_6941);
or U7903 (N_7903,N_6874,N_7272);
or U7904 (N_7904,N_6634,N_6968);
nor U7905 (N_7905,N_7463,N_6480);
and U7906 (N_7906,N_6951,N_6881);
or U7907 (N_7907,N_7343,N_6777);
nor U7908 (N_7908,N_7010,N_6860);
nand U7909 (N_7909,N_7123,N_7068);
nand U7910 (N_7910,N_6632,N_7064);
nor U7911 (N_7911,N_7024,N_6695);
nor U7912 (N_7912,N_6330,N_6803);
nor U7913 (N_7913,N_7286,N_7076);
or U7914 (N_7914,N_6085,N_7217);
or U7915 (N_7915,N_7245,N_6063);
nor U7916 (N_7916,N_6250,N_6786);
and U7917 (N_7917,N_6189,N_7384);
nor U7918 (N_7918,N_7341,N_6067);
and U7919 (N_7919,N_6567,N_6082);
or U7920 (N_7920,N_7048,N_6582);
nor U7921 (N_7921,N_7082,N_7427);
nor U7922 (N_7922,N_6674,N_7094);
nor U7923 (N_7923,N_6240,N_6372);
nor U7924 (N_7924,N_7012,N_6412);
nand U7925 (N_7925,N_6924,N_7377);
nor U7926 (N_7926,N_6871,N_6226);
and U7927 (N_7927,N_7365,N_7178);
nor U7928 (N_7928,N_6290,N_6193);
nor U7929 (N_7929,N_6922,N_6810);
or U7930 (N_7930,N_6737,N_6836);
nand U7931 (N_7931,N_6232,N_6617);
xnor U7932 (N_7932,N_6887,N_6669);
and U7933 (N_7933,N_7187,N_6512);
nor U7934 (N_7934,N_7294,N_7327);
xor U7935 (N_7935,N_7366,N_6723);
nor U7936 (N_7936,N_6659,N_6477);
nand U7937 (N_7937,N_7495,N_7397);
nand U7938 (N_7938,N_6945,N_6919);
nor U7939 (N_7939,N_6171,N_7435);
and U7940 (N_7940,N_6709,N_6834);
nor U7941 (N_7941,N_7070,N_7013);
nand U7942 (N_7942,N_6569,N_6220);
xnor U7943 (N_7943,N_7096,N_6537);
and U7944 (N_7944,N_6719,N_7413);
and U7945 (N_7945,N_6032,N_6086);
and U7946 (N_7946,N_6092,N_6407);
nand U7947 (N_7947,N_7473,N_6979);
nor U7948 (N_7948,N_6846,N_7363);
and U7949 (N_7949,N_6927,N_6116);
and U7950 (N_7950,N_6929,N_6280);
nor U7951 (N_7951,N_7088,N_6589);
or U7952 (N_7952,N_6702,N_6900);
or U7953 (N_7953,N_6768,N_6378);
or U7954 (N_7954,N_6687,N_6089);
nor U7955 (N_7955,N_6357,N_6447);
nor U7956 (N_7956,N_7290,N_6722);
nor U7957 (N_7957,N_6783,N_6152);
and U7958 (N_7958,N_6491,N_6361);
nand U7959 (N_7959,N_7025,N_7164);
nand U7960 (N_7960,N_7368,N_6106);
or U7961 (N_7961,N_7180,N_7399);
or U7962 (N_7962,N_6824,N_7491);
and U7963 (N_7963,N_7351,N_6311);
and U7964 (N_7964,N_6278,N_6429);
nand U7965 (N_7965,N_6376,N_7042);
nand U7966 (N_7966,N_6535,N_6700);
nor U7967 (N_7967,N_6242,N_7199);
nor U7968 (N_7968,N_6332,N_6610);
nor U7969 (N_7969,N_7315,N_6382);
nor U7970 (N_7970,N_6859,N_6751);
nor U7971 (N_7971,N_6198,N_7246);
or U7972 (N_7972,N_6053,N_6276);
nor U7973 (N_7973,N_7182,N_7219);
nand U7974 (N_7974,N_7058,N_6267);
nor U7975 (N_7975,N_7308,N_6422);
nand U7976 (N_7976,N_6628,N_6805);
or U7977 (N_7977,N_6223,N_6888);
or U7978 (N_7978,N_6182,N_6861);
nor U7979 (N_7979,N_6908,N_6345);
nand U7980 (N_7980,N_6257,N_7407);
nor U7981 (N_7981,N_6434,N_7462);
nor U7982 (N_7982,N_6095,N_7414);
or U7983 (N_7983,N_7305,N_6400);
or U7984 (N_7984,N_6048,N_6314);
and U7985 (N_7985,N_7410,N_6577);
or U7986 (N_7986,N_7253,N_7304);
nand U7987 (N_7987,N_6174,N_6991);
and U7988 (N_7988,N_6592,N_6985);
nor U7989 (N_7989,N_7362,N_6912);
nor U7990 (N_7990,N_6622,N_6375);
nor U7991 (N_7991,N_6901,N_6015);
nand U7992 (N_7992,N_7450,N_6849);
or U7993 (N_7993,N_7409,N_7255);
and U7994 (N_7994,N_7020,N_7265);
and U7995 (N_7995,N_6756,N_7262);
or U7996 (N_7996,N_7087,N_7467);
nor U7997 (N_7997,N_6525,N_7270);
nand U7998 (N_7998,N_6771,N_6911);
nor U7999 (N_7999,N_6677,N_6379);
or U8000 (N_8000,N_6203,N_6603);
nand U8001 (N_8001,N_6789,N_7116);
nor U8002 (N_8002,N_7015,N_7455);
nor U8003 (N_8003,N_6748,N_7484);
or U8004 (N_8004,N_7047,N_7405);
nand U8005 (N_8005,N_7201,N_6432);
nor U8006 (N_8006,N_6007,N_6995);
nor U8007 (N_8007,N_6812,N_7340);
and U8008 (N_8008,N_6052,N_6644);
nor U8009 (N_8009,N_6618,N_6394);
xor U8010 (N_8010,N_6417,N_6389);
and U8011 (N_8011,N_6131,N_6855);
nand U8012 (N_8012,N_7138,N_6272);
nor U8013 (N_8013,N_7000,N_7469);
nand U8014 (N_8014,N_7346,N_7349);
and U8015 (N_8015,N_6369,N_6795);
or U8016 (N_8016,N_6729,N_7324);
and U8017 (N_8017,N_6471,N_6446);
and U8018 (N_8018,N_6940,N_6960);
nor U8019 (N_8019,N_7153,N_6539);
nand U8020 (N_8020,N_7236,N_6562);
and U8021 (N_8021,N_6216,N_7350);
and U8022 (N_8022,N_7470,N_6406);
and U8023 (N_8023,N_6948,N_6602);
nand U8024 (N_8024,N_6891,N_6100);
nand U8025 (N_8025,N_6731,N_6463);
or U8026 (N_8026,N_7141,N_6342);
and U8027 (N_8027,N_6359,N_6897);
and U8028 (N_8028,N_6663,N_6279);
nor U8029 (N_8029,N_7408,N_7046);
and U8030 (N_8030,N_7442,N_6732);
nand U8031 (N_8031,N_6848,N_6213);
and U8032 (N_8032,N_6923,N_6531);
or U8033 (N_8033,N_6806,N_6346);
or U8034 (N_8034,N_6024,N_6821);
or U8035 (N_8035,N_6581,N_6122);
nand U8036 (N_8036,N_7269,N_6822);
nand U8037 (N_8037,N_6607,N_7481);
nand U8038 (N_8038,N_6818,N_6487);
and U8039 (N_8039,N_6757,N_7176);
nand U8040 (N_8040,N_7447,N_6427);
or U8041 (N_8041,N_6099,N_6555);
nor U8042 (N_8042,N_7376,N_6705);
nor U8043 (N_8043,N_6648,N_6511);
nand U8044 (N_8044,N_6595,N_7186);
and U8045 (N_8045,N_7492,N_7387);
and U8046 (N_8046,N_6124,N_7206);
nand U8047 (N_8047,N_6111,N_6021);
nor U8048 (N_8048,N_6448,N_6642);
nor U8049 (N_8049,N_6718,N_6014);
and U8050 (N_8050,N_6502,N_6270);
and U8051 (N_8051,N_6933,N_6275);
or U8052 (N_8052,N_6370,N_6749);
nand U8053 (N_8053,N_6580,N_6118);
nor U8054 (N_8054,N_6813,N_6934);
and U8055 (N_8055,N_6734,N_6631);
nand U8056 (N_8056,N_6696,N_6613);
nor U8057 (N_8057,N_6392,N_6844);
nand U8058 (N_8058,N_6265,N_6098);
and U8059 (N_8059,N_6486,N_7288);
nand U8060 (N_8060,N_7431,N_6411);
and U8061 (N_8061,N_7086,N_6865);
and U8062 (N_8062,N_6105,N_6035);
nor U8063 (N_8063,N_6845,N_6077);
or U8064 (N_8064,N_6005,N_6716);
or U8065 (N_8065,N_6556,N_6892);
or U8066 (N_8066,N_6792,N_7226);
and U8067 (N_8067,N_6545,N_6373);
or U8068 (N_8068,N_6423,N_6745);
nor U8069 (N_8069,N_6190,N_6224);
nand U8070 (N_8070,N_7145,N_7140);
nand U8071 (N_8071,N_6295,N_7029);
nand U8072 (N_8072,N_7113,N_7325);
or U8073 (N_8073,N_7152,N_6658);
or U8074 (N_8074,N_6640,N_6513);
or U8075 (N_8075,N_7355,N_6956);
nor U8076 (N_8076,N_6288,N_7374);
and U8077 (N_8077,N_7401,N_7471);
or U8078 (N_8078,N_7274,N_6518);
or U8079 (N_8079,N_7266,N_6438);
and U8080 (N_8080,N_6273,N_7136);
and U8081 (N_8081,N_7416,N_6011);
or U8082 (N_8082,N_6186,N_6484);
nand U8083 (N_8083,N_6656,N_6633);
nand U8084 (N_8084,N_6510,N_6670);
and U8085 (N_8085,N_7300,N_6654);
or U8086 (N_8086,N_7065,N_7193);
and U8087 (N_8087,N_7403,N_6215);
nand U8088 (N_8088,N_6145,N_7438);
and U8089 (N_8089,N_7074,N_6553);
nand U8090 (N_8090,N_7312,N_7129);
nor U8091 (N_8091,N_6614,N_6727);
or U8092 (N_8092,N_6980,N_6426);
nor U8093 (N_8093,N_7313,N_7225);
nor U8094 (N_8094,N_7287,N_6076);
and U8095 (N_8095,N_7101,N_6728);
or U8096 (N_8096,N_6641,N_6439);
and U8097 (N_8097,N_7434,N_6327);
nand U8098 (N_8098,N_7050,N_6156);
nand U8099 (N_8099,N_6065,N_6043);
and U8100 (N_8100,N_6148,N_7035);
and U8101 (N_8101,N_6325,N_7443);
xor U8102 (N_8102,N_7144,N_6442);
xnor U8103 (N_8103,N_6781,N_6738);
and U8104 (N_8104,N_6297,N_6460);
nand U8105 (N_8105,N_7488,N_7114);
nand U8106 (N_8106,N_7360,N_6880);
and U8107 (N_8107,N_6966,N_6925);
and U8108 (N_8108,N_6627,N_6078);
or U8109 (N_8109,N_7108,N_7297);
nand U8110 (N_8110,N_6879,N_6248);
and U8111 (N_8111,N_7357,N_7306);
nand U8112 (N_8112,N_7496,N_7060);
nand U8113 (N_8113,N_6527,N_6017);
and U8114 (N_8114,N_7448,N_7283);
nand U8115 (N_8115,N_7175,N_7093);
and U8116 (N_8116,N_6103,N_6194);
and U8117 (N_8117,N_7170,N_6104);
and U8118 (N_8118,N_7222,N_6652);
and U8119 (N_8119,N_7429,N_6551);
or U8120 (N_8120,N_6117,N_6636);
nor U8121 (N_8121,N_6975,N_6639);
nand U8122 (N_8122,N_6252,N_6158);
or U8123 (N_8123,N_7437,N_6470);
or U8124 (N_8124,N_6508,N_6606);
nor U8125 (N_8125,N_7075,N_6799);
nand U8126 (N_8126,N_6069,N_6126);
and U8127 (N_8127,N_6523,N_6253);
nand U8128 (N_8128,N_7007,N_6503);
and U8129 (N_8129,N_6289,N_6847);
or U8130 (N_8130,N_6886,N_6368);
or U8131 (N_8131,N_7119,N_7083);
or U8132 (N_8132,N_6548,N_6260);
and U8133 (N_8133,N_6264,N_7036);
and U8134 (N_8134,N_6504,N_6852);
and U8135 (N_8135,N_6391,N_7062);
and U8136 (N_8136,N_6167,N_6113);
or U8137 (N_8137,N_6316,N_7033);
or U8138 (N_8138,N_6499,N_6561);
and U8139 (N_8139,N_7072,N_6383);
or U8140 (N_8140,N_6001,N_6833);
nor U8141 (N_8141,N_6625,N_6760);
or U8142 (N_8142,N_6437,N_7039);
nand U8143 (N_8143,N_7347,N_6566);
or U8144 (N_8144,N_6755,N_6454);
nor U8145 (N_8145,N_7418,N_7465);
and U8146 (N_8146,N_6300,N_7057);
nor U8147 (N_8147,N_6661,N_6450);
or U8148 (N_8148,N_7361,N_6820);
nor U8149 (N_8149,N_7458,N_7211);
or U8150 (N_8150,N_7396,N_6725);
or U8151 (N_8151,N_6465,N_6239);
and U8152 (N_8152,N_6959,N_6651);
nand U8153 (N_8153,N_6864,N_7371);
and U8154 (N_8154,N_6637,N_6293);
nand U8155 (N_8155,N_6832,N_6823);
or U8156 (N_8156,N_6600,N_6474);
or U8157 (N_8157,N_6564,N_6336);
xor U8158 (N_8158,N_6839,N_7005);
xor U8159 (N_8159,N_6714,N_7054);
and U8160 (N_8160,N_6909,N_6072);
nor U8161 (N_8161,N_7161,N_6377);
and U8162 (N_8162,N_6742,N_6629);
nand U8163 (N_8163,N_6405,N_6643);
and U8164 (N_8164,N_6787,N_6885);
or U8165 (N_8165,N_7483,N_6801);
nand U8166 (N_8166,N_6743,N_6946);
nor U8167 (N_8167,N_7069,N_6498);
nor U8168 (N_8168,N_6475,N_7285);
nor U8169 (N_8169,N_7001,N_7021);
or U8170 (N_8170,N_7369,N_7111);
or U8171 (N_8171,N_6950,N_6044);
nand U8172 (N_8172,N_6752,N_6621);
nor U8173 (N_8173,N_6681,N_6920);
and U8174 (N_8174,N_6494,N_7275);
nand U8175 (N_8175,N_6856,N_7220);
nor U8176 (N_8176,N_6425,N_6421);
xnor U8177 (N_8177,N_6872,N_6797);
nor U8178 (N_8178,N_7204,N_6341);
and U8179 (N_8179,N_6424,N_6549);
and U8180 (N_8180,N_7314,N_6679);
nor U8181 (N_8181,N_6666,N_7372);
and U8182 (N_8182,N_7066,N_6262);
nand U8183 (N_8183,N_7430,N_7475);
nor U8184 (N_8184,N_6051,N_7034);
nor U8185 (N_8185,N_6736,N_6201);
nand U8186 (N_8186,N_6604,N_7332);
nand U8187 (N_8187,N_7406,N_6697);
and U8188 (N_8188,N_6664,N_6452);
or U8189 (N_8189,N_6192,N_6041);
nand U8190 (N_8190,N_6521,N_6584);
nand U8191 (N_8191,N_6596,N_6016);
nand U8192 (N_8192,N_6328,N_6008);
nor U8193 (N_8193,N_6733,N_6353);
or U8194 (N_8194,N_6227,N_6047);
nand U8195 (N_8195,N_6857,N_7348);
or U8196 (N_8196,N_7212,N_7100);
xor U8197 (N_8197,N_6247,N_7342);
nand U8198 (N_8198,N_7196,N_6006);
nand U8199 (N_8199,N_7378,N_6926);
or U8200 (N_8200,N_7446,N_6973);
nand U8201 (N_8201,N_6620,N_6455);
or U8202 (N_8202,N_6776,N_6075);
nand U8203 (N_8203,N_6009,N_6030);
and U8204 (N_8204,N_6707,N_6479);
xor U8205 (N_8205,N_6496,N_6916);
and U8206 (N_8206,N_6245,N_7395);
nand U8207 (N_8207,N_6798,N_7322);
and U8208 (N_8208,N_6042,N_7077);
nand U8209 (N_8209,N_7091,N_6500);
and U8210 (N_8210,N_6301,N_7264);
nor U8211 (N_8211,N_6000,N_7128);
nor U8212 (N_8212,N_6843,N_6277);
and U8213 (N_8213,N_6522,N_6937);
or U8214 (N_8214,N_6998,N_6576);
nand U8215 (N_8215,N_6730,N_6013);
or U8216 (N_8216,N_7198,N_6840);
or U8217 (N_8217,N_6796,N_6996);
nor U8218 (N_8218,N_7428,N_7130);
xor U8219 (N_8219,N_7071,N_6209);
nor U8220 (N_8220,N_7440,N_7016);
nand U8221 (N_8221,N_7359,N_6557);
or U8222 (N_8222,N_6060,N_6587);
and U8223 (N_8223,N_6944,N_7267);
nor U8224 (N_8224,N_7118,N_7234);
nor U8225 (N_8225,N_6873,N_6246);
nor U8226 (N_8226,N_7194,N_7309);
or U8227 (N_8227,N_6057,N_7146);
and U8228 (N_8228,N_7424,N_7457);
and U8229 (N_8229,N_7419,N_6256);
nand U8230 (N_8230,N_7102,N_6218);
and U8231 (N_8231,N_6079,N_6467);
and U8232 (N_8232,N_6791,N_6026);
nor U8233 (N_8233,N_7278,N_6187);
nor U8234 (N_8234,N_6601,N_6440);
nor U8235 (N_8235,N_7460,N_6693);
or U8236 (N_8236,N_7205,N_6271);
and U8237 (N_8237,N_7466,N_6313);
nor U8238 (N_8238,N_7331,N_6597);
nand U8239 (N_8239,N_6910,N_6160);
and U8240 (N_8240,N_6488,N_7207);
nand U8241 (N_8241,N_7490,N_7497);
and U8242 (N_8242,N_6784,N_6867);
and U8243 (N_8243,N_7472,N_6594);
and U8244 (N_8244,N_7279,N_6517);
nand U8245 (N_8245,N_6356,N_6994);
nand U8246 (N_8246,N_6036,N_6387);
and U8247 (N_8247,N_6129,N_7263);
nor U8248 (N_8248,N_6573,N_6010);
nand U8249 (N_8249,N_6413,N_6315);
nand U8250 (N_8250,N_7007,N_6398);
nor U8251 (N_8251,N_6237,N_6757);
xnor U8252 (N_8252,N_7247,N_7414);
nand U8253 (N_8253,N_7347,N_6196);
nand U8254 (N_8254,N_6423,N_7346);
or U8255 (N_8255,N_6500,N_6031);
nand U8256 (N_8256,N_6915,N_7027);
nor U8257 (N_8257,N_7053,N_6198);
nand U8258 (N_8258,N_7309,N_6003);
nor U8259 (N_8259,N_6589,N_7087);
nand U8260 (N_8260,N_6264,N_6688);
nor U8261 (N_8261,N_6086,N_6770);
nand U8262 (N_8262,N_6793,N_6307);
and U8263 (N_8263,N_7043,N_6097);
or U8264 (N_8264,N_6663,N_6099);
and U8265 (N_8265,N_6886,N_6190);
nor U8266 (N_8266,N_7096,N_6686);
or U8267 (N_8267,N_7251,N_7090);
nor U8268 (N_8268,N_6070,N_6764);
xor U8269 (N_8269,N_6764,N_6270);
and U8270 (N_8270,N_6325,N_6767);
nand U8271 (N_8271,N_6822,N_6652);
and U8272 (N_8272,N_6294,N_6330);
nor U8273 (N_8273,N_7422,N_6348);
and U8274 (N_8274,N_7388,N_7394);
nand U8275 (N_8275,N_6172,N_7292);
nor U8276 (N_8276,N_6467,N_7369);
and U8277 (N_8277,N_6986,N_6346);
nor U8278 (N_8278,N_6358,N_7131);
nor U8279 (N_8279,N_6667,N_7236);
nand U8280 (N_8280,N_7470,N_6932);
or U8281 (N_8281,N_6222,N_6756);
nand U8282 (N_8282,N_6240,N_7133);
or U8283 (N_8283,N_6882,N_6528);
or U8284 (N_8284,N_6451,N_7205);
nor U8285 (N_8285,N_7487,N_6565);
xnor U8286 (N_8286,N_7469,N_7109);
and U8287 (N_8287,N_7240,N_7010);
and U8288 (N_8288,N_7323,N_7436);
and U8289 (N_8289,N_6486,N_6124);
and U8290 (N_8290,N_6189,N_7317);
and U8291 (N_8291,N_6431,N_6894);
xnor U8292 (N_8292,N_6804,N_6761);
nand U8293 (N_8293,N_6390,N_6861);
nor U8294 (N_8294,N_6386,N_7250);
nor U8295 (N_8295,N_7165,N_6817);
nand U8296 (N_8296,N_6907,N_6570);
xor U8297 (N_8297,N_6763,N_6122);
nor U8298 (N_8298,N_6553,N_6431);
nand U8299 (N_8299,N_6531,N_6783);
or U8300 (N_8300,N_7058,N_7292);
nor U8301 (N_8301,N_7069,N_6302);
and U8302 (N_8302,N_7496,N_6364);
nor U8303 (N_8303,N_6129,N_7231);
and U8304 (N_8304,N_7196,N_7101);
and U8305 (N_8305,N_6663,N_6169);
or U8306 (N_8306,N_6068,N_6445);
nand U8307 (N_8307,N_6779,N_6243);
or U8308 (N_8308,N_6257,N_6296);
xnor U8309 (N_8309,N_7108,N_6533);
or U8310 (N_8310,N_7194,N_7255);
or U8311 (N_8311,N_6156,N_7135);
or U8312 (N_8312,N_6482,N_6461);
nand U8313 (N_8313,N_7394,N_6048);
nor U8314 (N_8314,N_6620,N_6671);
xnor U8315 (N_8315,N_6499,N_6784);
nand U8316 (N_8316,N_6997,N_6336);
nor U8317 (N_8317,N_6702,N_6758);
or U8318 (N_8318,N_6828,N_6609);
nor U8319 (N_8319,N_6571,N_7119);
and U8320 (N_8320,N_7474,N_6408);
and U8321 (N_8321,N_6974,N_6709);
nand U8322 (N_8322,N_7232,N_7484);
nand U8323 (N_8323,N_7441,N_6406);
nor U8324 (N_8324,N_7315,N_7171);
nor U8325 (N_8325,N_6873,N_6611);
nor U8326 (N_8326,N_6620,N_6907);
nand U8327 (N_8327,N_7122,N_6772);
and U8328 (N_8328,N_6328,N_7074);
nand U8329 (N_8329,N_6889,N_6281);
nand U8330 (N_8330,N_7456,N_7430);
nand U8331 (N_8331,N_6775,N_6925);
nand U8332 (N_8332,N_7012,N_6847);
nor U8333 (N_8333,N_6625,N_6140);
and U8334 (N_8334,N_7091,N_6368);
and U8335 (N_8335,N_6011,N_7121);
or U8336 (N_8336,N_6301,N_7073);
nand U8337 (N_8337,N_6036,N_7352);
nor U8338 (N_8338,N_6199,N_6120);
nand U8339 (N_8339,N_7363,N_6021);
or U8340 (N_8340,N_7331,N_6446);
nor U8341 (N_8341,N_6819,N_7303);
or U8342 (N_8342,N_6416,N_6145);
and U8343 (N_8343,N_6749,N_6161);
nor U8344 (N_8344,N_6764,N_6473);
nor U8345 (N_8345,N_6106,N_6069);
nand U8346 (N_8346,N_6574,N_7444);
or U8347 (N_8347,N_7448,N_7350);
and U8348 (N_8348,N_6883,N_6390);
nand U8349 (N_8349,N_7015,N_6536);
and U8350 (N_8350,N_6580,N_6035);
and U8351 (N_8351,N_6828,N_6981);
nand U8352 (N_8352,N_6147,N_7282);
nor U8353 (N_8353,N_7221,N_6611);
nor U8354 (N_8354,N_6149,N_7294);
xor U8355 (N_8355,N_6823,N_6780);
nand U8356 (N_8356,N_6612,N_7068);
nand U8357 (N_8357,N_6090,N_6189);
and U8358 (N_8358,N_6351,N_6696);
xnor U8359 (N_8359,N_6442,N_6609);
xnor U8360 (N_8360,N_7266,N_6280);
nand U8361 (N_8361,N_7126,N_6123);
nand U8362 (N_8362,N_6382,N_6127);
nand U8363 (N_8363,N_6575,N_6523);
and U8364 (N_8364,N_6340,N_6914);
nand U8365 (N_8365,N_6522,N_6138);
or U8366 (N_8366,N_6058,N_6368);
and U8367 (N_8367,N_6438,N_6207);
or U8368 (N_8368,N_7026,N_6597);
and U8369 (N_8369,N_6617,N_6021);
and U8370 (N_8370,N_6979,N_6342);
nor U8371 (N_8371,N_6730,N_7295);
nand U8372 (N_8372,N_7329,N_6285);
and U8373 (N_8373,N_6475,N_6213);
nand U8374 (N_8374,N_7231,N_7225);
and U8375 (N_8375,N_7019,N_7374);
and U8376 (N_8376,N_7408,N_6553);
or U8377 (N_8377,N_7304,N_7349);
or U8378 (N_8378,N_7066,N_6535);
or U8379 (N_8379,N_6725,N_6602);
and U8380 (N_8380,N_6557,N_6924);
and U8381 (N_8381,N_6786,N_7355);
nand U8382 (N_8382,N_6830,N_7012);
or U8383 (N_8383,N_6240,N_6364);
nor U8384 (N_8384,N_7304,N_6328);
nor U8385 (N_8385,N_6923,N_7330);
or U8386 (N_8386,N_7185,N_7109);
or U8387 (N_8387,N_6134,N_7288);
and U8388 (N_8388,N_6699,N_6926);
nand U8389 (N_8389,N_7315,N_6332);
and U8390 (N_8390,N_7473,N_6401);
nand U8391 (N_8391,N_6968,N_6019);
nand U8392 (N_8392,N_7277,N_7354);
nor U8393 (N_8393,N_7121,N_6283);
nor U8394 (N_8394,N_7147,N_6643);
or U8395 (N_8395,N_7311,N_7483);
nor U8396 (N_8396,N_6318,N_7025);
or U8397 (N_8397,N_6323,N_6097);
or U8398 (N_8398,N_6488,N_7230);
xor U8399 (N_8399,N_7466,N_6876);
nand U8400 (N_8400,N_6901,N_7030);
or U8401 (N_8401,N_6888,N_6381);
or U8402 (N_8402,N_7499,N_7351);
nor U8403 (N_8403,N_6666,N_7199);
nor U8404 (N_8404,N_6223,N_6139);
nor U8405 (N_8405,N_7474,N_6555);
or U8406 (N_8406,N_6101,N_7491);
nor U8407 (N_8407,N_6528,N_7069);
nor U8408 (N_8408,N_6475,N_6405);
nand U8409 (N_8409,N_7017,N_6364);
nand U8410 (N_8410,N_6874,N_6510);
and U8411 (N_8411,N_6220,N_7159);
nor U8412 (N_8412,N_6099,N_6591);
and U8413 (N_8413,N_7232,N_6932);
or U8414 (N_8414,N_6163,N_6837);
and U8415 (N_8415,N_6109,N_7041);
and U8416 (N_8416,N_6011,N_6319);
nor U8417 (N_8417,N_6310,N_6696);
or U8418 (N_8418,N_6509,N_7391);
or U8419 (N_8419,N_6920,N_7374);
nand U8420 (N_8420,N_6479,N_7282);
or U8421 (N_8421,N_6837,N_6227);
or U8422 (N_8422,N_7452,N_6293);
nor U8423 (N_8423,N_7354,N_6509);
or U8424 (N_8424,N_6154,N_7413);
or U8425 (N_8425,N_7363,N_7336);
and U8426 (N_8426,N_7195,N_7051);
nor U8427 (N_8427,N_6231,N_6575);
nand U8428 (N_8428,N_7434,N_6517);
and U8429 (N_8429,N_6546,N_6791);
or U8430 (N_8430,N_7453,N_6280);
nand U8431 (N_8431,N_6703,N_6108);
nand U8432 (N_8432,N_6982,N_6674);
and U8433 (N_8433,N_6288,N_6057);
nand U8434 (N_8434,N_7172,N_7499);
nor U8435 (N_8435,N_6363,N_7222);
or U8436 (N_8436,N_7391,N_6348);
nand U8437 (N_8437,N_6115,N_6758);
xor U8438 (N_8438,N_7379,N_6130);
or U8439 (N_8439,N_7046,N_6957);
nand U8440 (N_8440,N_7479,N_6627);
xnor U8441 (N_8441,N_6271,N_6911);
nor U8442 (N_8442,N_6937,N_6852);
nand U8443 (N_8443,N_6520,N_7233);
nand U8444 (N_8444,N_6177,N_6397);
nand U8445 (N_8445,N_7423,N_7213);
nand U8446 (N_8446,N_7145,N_7100);
and U8447 (N_8447,N_7248,N_7156);
nor U8448 (N_8448,N_7298,N_6020);
nor U8449 (N_8449,N_6977,N_6726);
nor U8450 (N_8450,N_6312,N_6617);
or U8451 (N_8451,N_7072,N_6316);
xnor U8452 (N_8452,N_6123,N_6392);
nor U8453 (N_8453,N_6704,N_6424);
nand U8454 (N_8454,N_7086,N_7038);
or U8455 (N_8455,N_7043,N_7489);
nand U8456 (N_8456,N_6028,N_7368);
and U8457 (N_8457,N_6304,N_7493);
nand U8458 (N_8458,N_7182,N_7391);
or U8459 (N_8459,N_7288,N_7031);
and U8460 (N_8460,N_6890,N_6298);
nand U8461 (N_8461,N_6509,N_6125);
nor U8462 (N_8462,N_7117,N_6435);
and U8463 (N_8463,N_6313,N_7418);
and U8464 (N_8464,N_6028,N_6694);
nand U8465 (N_8465,N_7192,N_6463);
nor U8466 (N_8466,N_6001,N_6610);
and U8467 (N_8467,N_7183,N_7477);
and U8468 (N_8468,N_6363,N_6099);
or U8469 (N_8469,N_6412,N_6207);
nand U8470 (N_8470,N_6572,N_6054);
nor U8471 (N_8471,N_6035,N_6097);
nand U8472 (N_8472,N_6788,N_6478);
or U8473 (N_8473,N_6866,N_7247);
nand U8474 (N_8474,N_6120,N_7401);
nor U8475 (N_8475,N_6111,N_6822);
nand U8476 (N_8476,N_6323,N_6894);
nor U8477 (N_8477,N_6068,N_7051);
nand U8478 (N_8478,N_6686,N_7491);
and U8479 (N_8479,N_6092,N_7119);
nor U8480 (N_8480,N_7335,N_7017);
and U8481 (N_8481,N_6754,N_7196);
nor U8482 (N_8482,N_7287,N_6289);
nand U8483 (N_8483,N_7202,N_7168);
nand U8484 (N_8484,N_7181,N_7485);
nand U8485 (N_8485,N_6440,N_6781);
nand U8486 (N_8486,N_6674,N_6539);
and U8487 (N_8487,N_6588,N_6424);
nand U8488 (N_8488,N_6735,N_6198);
nor U8489 (N_8489,N_6106,N_6864);
nand U8490 (N_8490,N_6370,N_6424);
nand U8491 (N_8491,N_6864,N_6092);
nor U8492 (N_8492,N_6983,N_7441);
nand U8493 (N_8493,N_7443,N_6001);
and U8494 (N_8494,N_7161,N_7164);
or U8495 (N_8495,N_6587,N_6320);
nand U8496 (N_8496,N_6984,N_6514);
nand U8497 (N_8497,N_6027,N_6941);
or U8498 (N_8498,N_6992,N_7413);
and U8499 (N_8499,N_7278,N_6492);
and U8500 (N_8500,N_6773,N_7348);
or U8501 (N_8501,N_6778,N_7114);
and U8502 (N_8502,N_7252,N_6895);
nand U8503 (N_8503,N_6158,N_7306);
or U8504 (N_8504,N_7253,N_6959);
or U8505 (N_8505,N_6152,N_6385);
nor U8506 (N_8506,N_6327,N_6006);
or U8507 (N_8507,N_7365,N_6559);
or U8508 (N_8508,N_7018,N_6694);
and U8509 (N_8509,N_6941,N_6311);
or U8510 (N_8510,N_7192,N_7172);
and U8511 (N_8511,N_6612,N_7289);
or U8512 (N_8512,N_6311,N_6140);
nand U8513 (N_8513,N_6155,N_6890);
or U8514 (N_8514,N_7112,N_6135);
and U8515 (N_8515,N_6958,N_7263);
and U8516 (N_8516,N_6375,N_7032);
nand U8517 (N_8517,N_6354,N_6572);
nand U8518 (N_8518,N_7032,N_6664);
nand U8519 (N_8519,N_6503,N_7127);
nand U8520 (N_8520,N_7159,N_7480);
nand U8521 (N_8521,N_6147,N_6334);
xnor U8522 (N_8522,N_7310,N_7284);
nor U8523 (N_8523,N_6826,N_6214);
or U8524 (N_8524,N_7171,N_7047);
nor U8525 (N_8525,N_7481,N_6395);
nand U8526 (N_8526,N_7025,N_7098);
and U8527 (N_8527,N_6629,N_6578);
and U8528 (N_8528,N_6672,N_7133);
nand U8529 (N_8529,N_6808,N_6099);
nor U8530 (N_8530,N_6690,N_6583);
xor U8531 (N_8531,N_7382,N_6799);
nand U8532 (N_8532,N_6844,N_6878);
or U8533 (N_8533,N_7412,N_6092);
and U8534 (N_8534,N_6488,N_6963);
and U8535 (N_8535,N_6944,N_6317);
nor U8536 (N_8536,N_7436,N_6117);
or U8537 (N_8537,N_6282,N_6012);
nor U8538 (N_8538,N_6219,N_6782);
and U8539 (N_8539,N_6786,N_6872);
and U8540 (N_8540,N_6402,N_7465);
and U8541 (N_8541,N_7201,N_6674);
nand U8542 (N_8542,N_6735,N_6227);
nor U8543 (N_8543,N_7213,N_6569);
nand U8544 (N_8544,N_6340,N_6177);
nand U8545 (N_8545,N_6520,N_6004);
nor U8546 (N_8546,N_6695,N_6629);
nor U8547 (N_8547,N_6989,N_7164);
and U8548 (N_8548,N_7366,N_6901);
nand U8549 (N_8549,N_6897,N_6630);
or U8550 (N_8550,N_6515,N_7121);
nor U8551 (N_8551,N_7186,N_6164);
nand U8552 (N_8552,N_6122,N_7476);
or U8553 (N_8553,N_6922,N_6127);
nand U8554 (N_8554,N_7034,N_7297);
and U8555 (N_8555,N_6391,N_7018);
and U8556 (N_8556,N_7387,N_7001);
and U8557 (N_8557,N_6347,N_7284);
xnor U8558 (N_8558,N_7407,N_6812);
and U8559 (N_8559,N_6626,N_7494);
and U8560 (N_8560,N_6171,N_6271);
and U8561 (N_8561,N_6917,N_6466);
and U8562 (N_8562,N_6394,N_6300);
nand U8563 (N_8563,N_6531,N_7175);
and U8564 (N_8564,N_6827,N_7365);
nand U8565 (N_8565,N_6354,N_7169);
nand U8566 (N_8566,N_7023,N_6026);
or U8567 (N_8567,N_7402,N_7488);
nand U8568 (N_8568,N_7495,N_6748);
nand U8569 (N_8569,N_6742,N_7117);
and U8570 (N_8570,N_6982,N_7436);
and U8571 (N_8571,N_6080,N_7404);
xor U8572 (N_8572,N_6865,N_7097);
nor U8573 (N_8573,N_6504,N_6792);
nor U8574 (N_8574,N_6394,N_7043);
nor U8575 (N_8575,N_6512,N_7328);
xnor U8576 (N_8576,N_6822,N_7126);
nor U8577 (N_8577,N_6255,N_6858);
nand U8578 (N_8578,N_6413,N_7187);
and U8579 (N_8579,N_6276,N_6085);
nand U8580 (N_8580,N_7088,N_6581);
and U8581 (N_8581,N_6170,N_6024);
nand U8582 (N_8582,N_7078,N_6400);
nor U8583 (N_8583,N_6046,N_6516);
nor U8584 (N_8584,N_6172,N_7067);
nand U8585 (N_8585,N_6012,N_7410);
nand U8586 (N_8586,N_6810,N_6338);
nand U8587 (N_8587,N_6878,N_6486);
and U8588 (N_8588,N_6145,N_6526);
and U8589 (N_8589,N_6208,N_6350);
nand U8590 (N_8590,N_6743,N_6025);
and U8591 (N_8591,N_6993,N_7256);
nor U8592 (N_8592,N_6769,N_7450);
nand U8593 (N_8593,N_7193,N_6554);
and U8594 (N_8594,N_7018,N_7034);
nor U8595 (N_8595,N_7078,N_7034);
and U8596 (N_8596,N_7395,N_7161);
or U8597 (N_8597,N_7433,N_6258);
nand U8598 (N_8598,N_6297,N_6665);
nor U8599 (N_8599,N_6117,N_6215);
and U8600 (N_8600,N_6329,N_6331);
nor U8601 (N_8601,N_7176,N_7487);
xor U8602 (N_8602,N_6101,N_6712);
and U8603 (N_8603,N_6973,N_6619);
xor U8604 (N_8604,N_6313,N_6410);
or U8605 (N_8605,N_6584,N_7142);
nand U8606 (N_8606,N_7414,N_7080);
and U8607 (N_8607,N_6652,N_6130);
nor U8608 (N_8608,N_6701,N_7248);
or U8609 (N_8609,N_6333,N_6305);
nor U8610 (N_8610,N_7244,N_7424);
or U8611 (N_8611,N_7234,N_6040);
nor U8612 (N_8612,N_6351,N_7318);
and U8613 (N_8613,N_6884,N_6229);
xnor U8614 (N_8614,N_7303,N_6735);
and U8615 (N_8615,N_6144,N_6596);
and U8616 (N_8616,N_7350,N_6881);
and U8617 (N_8617,N_6075,N_6673);
and U8618 (N_8618,N_6444,N_6048);
and U8619 (N_8619,N_6250,N_6207);
or U8620 (N_8620,N_7041,N_6929);
nand U8621 (N_8621,N_6933,N_6940);
nor U8622 (N_8622,N_6320,N_7365);
or U8623 (N_8623,N_7314,N_6677);
nand U8624 (N_8624,N_6075,N_6871);
or U8625 (N_8625,N_6154,N_6488);
nor U8626 (N_8626,N_7091,N_6803);
or U8627 (N_8627,N_6131,N_6976);
nand U8628 (N_8628,N_7357,N_6149);
nor U8629 (N_8629,N_6430,N_6965);
or U8630 (N_8630,N_6951,N_7230);
and U8631 (N_8631,N_7455,N_7134);
nor U8632 (N_8632,N_6895,N_6493);
and U8633 (N_8633,N_6367,N_6520);
nor U8634 (N_8634,N_6878,N_6419);
nor U8635 (N_8635,N_6469,N_6173);
nand U8636 (N_8636,N_6730,N_6948);
and U8637 (N_8637,N_6718,N_6397);
and U8638 (N_8638,N_7049,N_6594);
nand U8639 (N_8639,N_7499,N_7073);
xor U8640 (N_8640,N_6854,N_6358);
nor U8641 (N_8641,N_7257,N_6467);
nand U8642 (N_8642,N_6030,N_6965);
and U8643 (N_8643,N_6111,N_6300);
or U8644 (N_8644,N_6338,N_6873);
nand U8645 (N_8645,N_6795,N_7474);
or U8646 (N_8646,N_7261,N_6437);
nor U8647 (N_8647,N_6736,N_6958);
or U8648 (N_8648,N_6222,N_6121);
and U8649 (N_8649,N_6118,N_6841);
and U8650 (N_8650,N_6584,N_6204);
nor U8651 (N_8651,N_7359,N_6429);
nor U8652 (N_8652,N_6269,N_7218);
nor U8653 (N_8653,N_7102,N_6661);
or U8654 (N_8654,N_7192,N_6235);
and U8655 (N_8655,N_7020,N_6761);
and U8656 (N_8656,N_7228,N_6669);
or U8657 (N_8657,N_6750,N_6765);
nand U8658 (N_8658,N_7295,N_6250);
or U8659 (N_8659,N_7339,N_7234);
or U8660 (N_8660,N_7128,N_6570);
nor U8661 (N_8661,N_6541,N_7363);
and U8662 (N_8662,N_7419,N_7059);
nand U8663 (N_8663,N_6100,N_6012);
nor U8664 (N_8664,N_6843,N_6801);
nand U8665 (N_8665,N_6294,N_7341);
nand U8666 (N_8666,N_6103,N_6057);
nand U8667 (N_8667,N_6067,N_7282);
or U8668 (N_8668,N_6239,N_6058);
nand U8669 (N_8669,N_6033,N_6157);
nand U8670 (N_8670,N_6855,N_7400);
nor U8671 (N_8671,N_7492,N_6916);
nand U8672 (N_8672,N_6268,N_6754);
and U8673 (N_8673,N_6784,N_6048);
nor U8674 (N_8674,N_6026,N_6217);
or U8675 (N_8675,N_6365,N_7346);
xnor U8676 (N_8676,N_6124,N_6540);
or U8677 (N_8677,N_7356,N_6950);
nand U8678 (N_8678,N_6706,N_6878);
nor U8679 (N_8679,N_7298,N_6699);
nor U8680 (N_8680,N_6190,N_6428);
nand U8681 (N_8681,N_6659,N_7065);
nand U8682 (N_8682,N_7414,N_6185);
or U8683 (N_8683,N_6233,N_6270);
or U8684 (N_8684,N_7219,N_6505);
nor U8685 (N_8685,N_6331,N_6593);
or U8686 (N_8686,N_6882,N_6331);
and U8687 (N_8687,N_7473,N_6578);
and U8688 (N_8688,N_6846,N_7258);
xnor U8689 (N_8689,N_6726,N_6599);
nand U8690 (N_8690,N_6619,N_7208);
nor U8691 (N_8691,N_6840,N_7176);
or U8692 (N_8692,N_7151,N_6604);
nand U8693 (N_8693,N_6384,N_7341);
nor U8694 (N_8694,N_6894,N_6942);
nand U8695 (N_8695,N_7106,N_6701);
nand U8696 (N_8696,N_7363,N_6668);
nand U8697 (N_8697,N_6321,N_6713);
nor U8698 (N_8698,N_6364,N_6604);
nand U8699 (N_8699,N_6985,N_6130);
nand U8700 (N_8700,N_6159,N_6087);
or U8701 (N_8701,N_6256,N_6764);
and U8702 (N_8702,N_6465,N_6527);
or U8703 (N_8703,N_6440,N_6177);
or U8704 (N_8704,N_6010,N_6976);
nor U8705 (N_8705,N_6435,N_6431);
nand U8706 (N_8706,N_6388,N_6571);
or U8707 (N_8707,N_7453,N_7389);
xor U8708 (N_8708,N_7410,N_6593);
nor U8709 (N_8709,N_7357,N_6630);
nand U8710 (N_8710,N_6862,N_6962);
nand U8711 (N_8711,N_6633,N_6472);
nor U8712 (N_8712,N_6360,N_6399);
and U8713 (N_8713,N_6138,N_7169);
or U8714 (N_8714,N_7329,N_6200);
nand U8715 (N_8715,N_7164,N_6991);
nand U8716 (N_8716,N_6388,N_6701);
or U8717 (N_8717,N_6265,N_7197);
nor U8718 (N_8718,N_7263,N_7119);
nor U8719 (N_8719,N_7198,N_6842);
or U8720 (N_8720,N_6671,N_6755);
nand U8721 (N_8721,N_6155,N_6928);
nand U8722 (N_8722,N_6293,N_6476);
or U8723 (N_8723,N_6305,N_6555);
nand U8724 (N_8724,N_7482,N_6202);
or U8725 (N_8725,N_6858,N_6904);
nand U8726 (N_8726,N_7286,N_7365);
nor U8727 (N_8727,N_6240,N_6824);
or U8728 (N_8728,N_6846,N_6584);
xor U8729 (N_8729,N_6555,N_7410);
or U8730 (N_8730,N_7322,N_6736);
or U8731 (N_8731,N_6593,N_6848);
or U8732 (N_8732,N_6305,N_6606);
or U8733 (N_8733,N_6492,N_6069);
and U8734 (N_8734,N_6298,N_6098);
nor U8735 (N_8735,N_6343,N_7052);
or U8736 (N_8736,N_7072,N_6141);
nor U8737 (N_8737,N_6265,N_6156);
nor U8738 (N_8738,N_6383,N_6501);
nand U8739 (N_8739,N_6600,N_6551);
and U8740 (N_8740,N_6226,N_7468);
xnor U8741 (N_8741,N_6625,N_6225);
and U8742 (N_8742,N_6573,N_7101);
or U8743 (N_8743,N_7333,N_6428);
and U8744 (N_8744,N_7353,N_7345);
nand U8745 (N_8745,N_7092,N_6053);
nand U8746 (N_8746,N_6966,N_6522);
and U8747 (N_8747,N_6645,N_6881);
and U8748 (N_8748,N_6732,N_6944);
nor U8749 (N_8749,N_6644,N_6428);
and U8750 (N_8750,N_7038,N_7390);
nand U8751 (N_8751,N_6457,N_7474);
nand U8752 (N_8752,N_7337,N_6532);
and U8753 (N_8753,N_6335,N_6925);
and U8754 (N_8754,N_7101,N_6896);
nand U8755 (N_8755,N_6203,N_6809);
and U8756 (N_8756,N_7338,N_6544);
and U8757 (N_8757,N_6012,N_6905);
and U8758 (N_8758,N_6228,N_6724);
and U8759 (N_8759,N_6354,N_6052);
nand U8760 (N_8760,N_6884,N_7379);
nor U8761 (N_8761,N_6094,N_6298);
nor U8762 (N_8762,N_7162,N_7337);
or U8763 (N_8763,N_7062,N_6511);
nand U8764 (N_8764,N_6462,N_7084);
nand U8765 (N_8765,N_6064,N_7022);
and U8766 (N_8766,N_7345,N_7159);
nand U8767 (N_8767,N_7004,N_6470);
nand U8768 (N_8768,N_6270,N_6615);
nand U8769 (N_8769,N_7092,N_7398);
or U8770 (N_8770,N_6421,N_6036);
or U8771 (N_8771,N_6907,N_6420);
or U8772 (N_8772,N_6083,N_6740);
and U8773 (N_8773,N_6728,N_6985);
or U8774 (N_8774,N_7092,N_6629);
nor U8775 (N_8775,N_7038,N_7433);
nand U8776 (N_8776,N_6491,N_6135);
or U8777 (N_8777,N_7421,N_6934);
nor U8778 (N_8778,N_6667,N_6037);
nor U8779 (N_8779,N_6121,N_6290);
xor U8780 (N_8780,N_6096,N_6317);
or U8781 (N_8781,N_6757,N_7023);
nand U8782 (N_8782,N_7116,N_7404);
nor U8783 (N_8783,N_6116,N_6134);
nor U8784 (N_8784,N_7139,N_7086);
nor U8785 (N_8785,N_6585,N_7197);
xor U8786 (N_8786,N_7298,N_6014);
nor U8787 (N_8787,N_6260,N_6820);
nand U8788 (N_8788,N_6605,N_6800);
nor U8789 (N_8789,N_7305,N_6646);
and U8790 (N_8790,N_6837,N_6276);
nand U8791 (N_8791,N_6766,N_6413);
or U8792 (N_8792,N_7450,N_6047);
or U8793 (N_8793,N_7254,N_6261);
and U8794 (N_8794,N_6808,N_6913);
nand U8795 (N_8795,N_6344,N_7154);
nor U8796 (N_8796,N_6228,N_6138);
and U8797 (N_8797,N_6680,N_6123);
nand U8798 (N_8798,N_6784,N_6697);
nor U8799 (N_8799,N_6883,N_7444);
nand U8800 (N_8800,N_7360,N_7254);
or U8801 (N_8801,N_6708,N_6339);
nand U8802 (N_8802,N_6757,N_7339);
and U8803 (N_8803,N_6915,N_6474);
nor U8804 (N_8804,N_7486,N_6072);
nor U8805 (N_8805,N_6321,N_6683);
or U8806 (N_8806,N_6308,N_6361);
or U8807 (N_8807,N_6105,N_6842);
nor U8808 (N_8808,N_6079,N_6024);
or U8809 (N_8809,N_6955,N_6753);
nand U8810 (N_8810,N_7204,N_6788);
xor U8811 (N_8811,N_7053,N_6080);
xor U8812 (N_8812,N_6116,N_6170);
and U8813 (N_8813,N_6307,N_6001);
nand U8814 (N_8814,N_6910,N_7172);
and U8815 (N_8815,N_7022,N_7475);
or U8816 (N_8816,N_7255,N_7319);
and U8817 (N_8817,N_6458,N_7115);
and U8818 (N_8818,N_6280,N_6984);
nand U8819 (N_8819,N_6471,N_6008);
and U8820 (N_8820,N_7386,N_6690);
and U8821 (N_8821,N_7204,N_7351);
and U8822 (N_8822,N_6298,N_6285);
or U8823 (N_8823,N_7019,N_6728);
nand U8824 (N_8824,N_7086,N_6597);
and U8825 (N_8825,N_7451,N_6680);
or U8826 (N_8826,N_6689,N_7236);
xor U8827 (N_8827,N_6311,N_6606);
and U8828 (N_8828,N_7425,N_7368);
nand U8829 (N_8829,N_7362,N_7113);
nor U8830 (N_8830,N_6214,N_6660);
or U8831 (N_8831,N_6205,N_6320);
nand U8832 (N_8832,N_6268,N_6319);
nor U8833 (N_8833,N_6132,N_6089);
and U8834 (N_8834,N_6873,N_6318);
nand U8835 (N_8835,N_6148,N_6173);
or U8836 (N_8836,N_7498,N_6532);
or U8837 (N_8837,N_7180,N_6050);
and U8838 (N_8838,N_7479,N_6428);
nand U8839 (N_8839,N_7141,N_6843);
or U8840 (N_8840,N_7498,N_6376);
nand U8841 (N_8841,N_7093,N_6499);
nor U8842 (N_8842,N_7084,N_6078);
and U8843 (N_8843,N_7075,N_6596);
and U8844 (N_8844,N_6522,N_6720);
xnor U8845 (N_8845,N_7326,N_7279);
nand U8846 (N_8846,N_6387,N_6589);
and U8847 (N_8847,N_6007,N_6749);
or U8848 (N_8848,N_6111,N_7273);
nand U8849 (N_8849,N_6694,N_6738);
or U8850 (N_8850,N_7120,N_7113);
nor U8851 (N_8851,N_6668,N_6738);
and U8852 (N_8852,N_6825,N_7309);
or U8853 (N_8853,N_7130,N_6785);
and U8854 (N_8854,N_7083,N_6595);
and U8855 (N_8855,N_6001,N_6509);
nor U8856 (N_8856,N_7252,N_7007);
and U8857 (N_8857,N_7018,N_6648);
nand U8858 (N_8858,N_7451,N_6926);
nor U8859 (N_8859,N_7039,N_7236);
nand U8860 (N_8860,N_7320,N_6538);
nand U8861 (N_8861,N_6663,N_7460);
nand U8862 (N_8862,N_6118,N_6473);
xnor U8863 (N_8863,N_6223,N_6450);
xor U8864 (N_8864,N_6967,N_6263);
nand U8865 (N_8865,N_7458,N_6542);
and U8866 (N_8866,N_6692,N_6980);
or U8867 (N_8867,N_7134,N_7331);
and U8868 (N_8868,N_6065,N_6734);
nor U8869 (N_8869,N_6405,N_6839);
xnor U8870 (N_8870,N_7061,N_6925);
nor U8871 (N_8871,N_7037,N_7430);
or U8872 (N_8872,N_6893,N_6738);
nor U8873 (N_8873,N_6183,N_6602);
and U8874 (N_8874,N_6452,N_7122);
and U8875 (N_8875,N_6209,N_6247);
nor U8876 (N_8876,N_7341,N_7413);
or U8877 (N_8877,N_6406,N_6616);
nand U8878 (N_8878,N_6857,N_7242);
or U8879 (N_8879,N_6111,N_6167);
nor U8880 (N_8880,N_6545,N_6455);
nand U8881 (N_8881,N_6630,N_6742);
nand U8882 (N_8882,N_6121,N_6230);
nand U8883 (N_8883,N_6428,N_6445);
nand U8884 (N_8884,N_7373,N_6736);
nor U8885 (N_8885,N_6268,N_6919);
nand U8886 (N_8886,N_6482,N_6090);
and U8887 (N_8887,N_6920,N_7132);
nand U8888 (N_8888,N_6100,N_7303);
or U8889 (N_8889,N_7237,N_6175);
or U8890 (N_8890,N_6997,N_6274);
and U8891 (N_8891,N_6131,N_6270);
or U8892 (N_8892,N_6138,N_6722);
or U8893 (N_8893,N_6377,N_7253);
nand U8894 (N_8894,N_7280,N_7001);
and U8895 (N_8895,N_6661,N_6556);
nor U8896 (N_8896,N_6629,N_7042);
nand U8897 (N_8897,N_7139,N_6990);
nand U8898 (N_8898,N_6233,N_6530);
nand U8899 (N_8899,N_6975,N_6202);
and U8900 (N_8900,N_6093,N_6025);
xnor U8901 (N_8901,N_6751,N_6622);
nand U8902 (N_8902,N_7456,N_7065);
nand U8903 (N_8903,N_6043,N_6974);
and U8904 (N_8904,N_6761,N_6067);
or U8905 (N_8905,N_7246,N_6679);
and U8906 (N_8906,N_6937,N_6302);
nand U8907 (N_8907,N_6778,N_7074);
or U8908 (N_8908,N_6801,N_6154);
and U8909 (N_8909,N_6131,N_6235);
nand U8910 (N_8910,N_6644,N_6501);
and U8911 (N_8911,N_6966,N_6309);
and U8912 (N_8912,N_6450,N_6542);
and U8913 (N_8913,N_6680,N_6983);
nand U8914 (N_8914,N_6428,N_7459);
nor U8915 (N_8915,N_6774,N_6935);
and U8916 (N_8916,N_6918,N_7481);
and U8917 (N_8917,N_6619,N_7397);
nand U8918 (N_8918,N_6550,N_6456);
nand U8919 (N_8919,N_6736,N_6141);
nor U8920 (N_8920,N_6896,N_6278);
nand U8921 (N_8921,N_7341,N_6473);
nor U8922 (N_8922,N_6787,N_6194);
nand U8923 (N_8923,N_6434,N_7397);
and U8924 (N_8924,N_6892,N_6688);
nand U8925 (N_8925,N_6161,N_6785);
nor U8926 (N_8926,N_6907,N_6521);
or U8927 (N_8927,N_6096,N_6524);
nor U8928 (N_8928,N_7241,N_7042);
nand U8929 (N_8929,N_6488,N_6092);
or U8930 (N_8930,N_6934,N_6592);
or U8931 (N_8931,N_6680,N_7069);
nand U8932 (N_8932,N_7265,N_7057);
nor U8933 (N_8933,N_7228,N_6403);
nand U8934 (N_8934,N_6846,N_6920);
nor U8935 (N_8935,N_6094,N_6242);
nand U8936 (N_8936,N_6705,N_6281);
and U8937 (N_8937,N_6316,N_7006);
or U8938 (N_8938,N_7009,N_7368);
and U8939 (N_8939,N_7113,N_6394);
nor U8940 (N_8940,N_7110,N_7035);
or U8941 (N_8941,N_6871,N_6478);
nor U8942 (N_8942,N_6056,N_6845);
nand U8943 (N_8943,N_6550,N_6645);
or U8944 (N_8944,N_7389,N_6134);
nor U8945 (N_8945,N_6382,N_6063);
nor U8946 (N_8946,N_6084,N_6295);
and U8947 (N_8947,N_6817,N_6004);
and U8948 (N_8948,N_6867,N_6341);
nor U8949 (N_8949,N_6808,N_6338);
xor U8950 (N_8950,N_6999,N_6924);
nand U8951 (N_8951,N_7351,N_6169);
and U8952 (N_8952,N_6375,N_6658);
nand U8953 (N_8953,N_6260,N_6047);
and U8954 (N_8954,N_6375,N_6347);
nor U8955 (N_8955,N_7002,N_7396);
and U8956 (N_8956,N_7030,N_7003);
nor U8957 (N_8957,N_6330,N_6036);
or U8958 (N_8958,N_6036,N_7162);
nor U8959 (N_8959,N_6611,N_6926);
and U8960 (N_8960,N_7428,N_6470);
nor U8961 (N_8961,N_7429,N_6286);
and U8962 (N_8962,N_6065,N_6446);
xor U8963 (N_8963,N_6955,N_7297);
nand U8964 (N_8964,N_6573,N_7148);
and U8965 (N_8965,N_6042,N_6238);
or U8966 (N_8966,N_6709,N_6150);
nand U8967 (N_8967,N_7407,N_6133);
or U8968 (N_8968,N_6216,N_6824);
nor U8969 (N_8969,N_6501,N_6001);
and U8970 (N_8970,N_6266,N_6747);
and U8971 (N_8971,N_6285,N_7412);
or U8972 (N_8972,N_6128,N_6478);
nand U8973 (N_8973,N_6933,N_7495);
nand U8974 (N_8974,N_6819,N_6190);
nand U8975 (N_8975,N_6777,N_6123);
nand U8976 (N_8976,N_6510,N_6779);
or U8977 (N_8977,N_7022,N_6566);
xor U8978 (N_8978,N_6722,N_7352);
and U8979 (N_8979,N_6145,N_6009);
nand U8980 (N_8980,N_6705,N_6233);
and U8981 (N_8981,N_6746,N_6248);
nor U8982 (N_8982,N_6400,N_6556);
or U8983 (N_8983,N_7071,N_6489);
nor U8984 (N_8984,N_7180,N_6378);
nand U8985 (N_8985,N_6567,N_6408);
or U8986 (N_8986,N_6353,N_7009);
or U8987 (N_8987,N_7358,N_6669);
xnor U8988 (N_8988,N_6357,N_6051);
nor U8989 (N_8989,N_7042,N_6345);
nor U8990 (N_8990,N_6667,N_7134);
and U8991 (N_8991,N_6096,N_6519);
or U8992 (N_8992,N_6377,N_6567);
nand U8993 (N_8993,N_6351,N_6954);
or U8994 (N_8994,N_6247,N_7402);
nor U8995 (N_8995,N_6860,N_7080);
or U8996 (N_8996,N_6748,N_6201);
nor U8997 (N_8997,N_7085,N_7456);
nor U8998 (N_8998,N_6374,N_6219);
nand U8999 (N_8999,N_6895,N_7240);
nor U9000 (N_9000,N_7504,N_8170);
nand U9001 (N_9001,N_8911,N_8960);
and U9002 (N_9002,N_7744,N_7646);
nand U9003 (N_9003,N_8383,N_8281);
and U9004 (N_9004,N_7885,N_8063);
or U9005 (N_9005,N_8958,N_8735);
xor U9006 (N_9006,N_7692,N_7774);
nand U9007 (N_9007,N_8458,N_7570);
nor U9008 (N_9008,N_7811,N_8250);
nor U9009 (N_9009,N_8898,N_8892);
or U9010 (N_9010,N_8502,N_8326);
nand U9011 (N_9011,N_8932,N_7889);
and U9012 (N_9012,N_8470,N_8738);
and U9013 (N_9013,N_8726,N_7933);
nand U9014 (N_9014,N_8113,N_7729);
or U9015 (N_9015,N_8890,N_8607);
nor U9016 (N_9016,N_8151,N_7622);
nand U9017 (N_9017,N_7952,N_8159);
or U9018 (N_9018,N_7942,N_7664);
nor U9019 (N_9019,N_7777,N_7533);
xnor U9020 (N_9020,N_8843,N_8328);
or U9021 (N_9021,N_7545,N_7963);
and U9022 (N_9022,N_8247,N_8036);
xnor U9023 (N_9023,N_7608,N_8216);
or U9024 (N_9024,N_8256,N_8736);
nor U9025 (N_9025,N_7542,N_7937);
or U9026 (N_9026,N_8220,N_7939);
and U9027 (N_9027,N_7629,N_7865);
nor U9028 (N_9028,N_8079,N_8525);
nand U9029 (N_9029,N_8972,N_7965);
nor U9030 (N_9030,N_7678,N_8287);
and U9031 (N_9031,N_8872,N_8059);
nand U9032 (N_9032,N_8871,N_8436);
or U9033 (N_9033,N_7881,N_8765);
nand U9034 (N_9034,N_8424,N_8795);
and U9035 (N_9035,N_8303,N_8939);
and U9036 (N_9036,N_7901,N_7649);
or U9037 (N_9037,N_8663,N_8096);
or U9038 (N_9038,N_8002,N_7945);
nand U9039 (N_9039,N_8650,N_7958);
or U9040 (N_9040,N_7872,N_8676);
nand U9041 (N_9041,N_7663,N_8563);
or U9042 (N_9042,N_8329,N_7908);
nor U9043 (N_9043,N_8373,N_8507);
nor U9044 (N_9044,N_7603,N_8123);
and U9045 (N_9045,N_8009,N_8644);
nor U9046 (N_9046,N_7943,N_7920);
nor U9047 (N_9047,N_7696,N_8488);
or U9048 (N_9048,N_8440,N_8249);
nor U9049 (N_9049,N_8949,N_8666);
and U9050 (N_9050,N_8980,N_8512);
nand U9051 (N_9051,N_7589,N_8131);
nand U9052 (N_9052,N_8395,N_7806);
nand U9053 (N_9053,N_8837,N_8201);
and U9054 (N_9054,N_8610,N_8711);
nor U9055 (N_9055,N_7707,N_8126);
or U9056 (N_9056,N_8906,N_7807);
and U9057 (N_9057,N_8990,N_8446);
nand U9058 (N_9058,N_8978,N_8881);
and U9059 (N_9059,N_7572,N_7667);
nand U9060 (N_9060,N_7548,N_8192);
or U9061 (N_9061,N_8882,N_8724);
or U9062 (N_9062,N_8380,N_7668);
nor U9063 (N_9063,N_7553,N_8116);
and U9064 (N_9064,N_7932,N_8412);
nand U9065 (N_9065,N_8087,N_8697);
nor U9066 (N_9066,N_7573,N_8677);
nor U9067 (N_9067,N_7623,N_8127);
nor U9068 (N_9068,N_8505,N_7565);
xor U9069 (N_9069,N_7611,N_7948);
and U9070 (N_9070,N_8439,N_7618);
and U9071 (N_9071,N_8879,N_7754);
and U9072 (N_9072,N_8323,N_8503);
and U9073 (N_9073,N_8908,N_7673);
or U9074 (N_9074,N_8902,N_8771);
nand U9075 (N_9075,N_7640,N_7964);
and U9076 (N_9076,N_8518,N_8717);
nor U9077 (N_9077,N_7561,N_8046);
nand U9078 (N_9078,N_8073,N_8917);
or U9079 (N_9079,N_8385,N_8211);
nand U9080 (N_9080,N_8108,N_8386);
and U9081 (N_9081,N_8802,N_8365);
nand U9082 (N_9082,N_8334,N_8179);
or U9083 (N_9083,N_7656,N_8751);
nor U9084 (N_9084,N_8725,N_8915);
and U9085 (N_9085,N_8613,N_8234);
nand U9086 (N_9086,N_8188,N_7802);
and U9087 (N_9087,N_8407,N_7600);
nor U9088 (N_9088,N_8855,N_8927);
nand U9089 (N_9089,N_8072,N_8346);
nand U9090 (N_9090,N_8943,N_7816);
and U9091 (N_9091,N_7812,N_8950);
and U9092 (N_9092,N_8683,N_8461);
nand U9093 (N_9093,N_8444,N_8348);
or U9094 (N_9094,N_8402,N_8624);
or U9095 (N_9095,N_8698,N_8769);
or U9096 (N_9096,N_8430,N_7680);
nand U9097 (N_9097,N_7796,N_8028);
nand U9098 (N_9098,N_8626,N_7890);
and U9099 (N_9099,N_8618,N_8081);
and U9100 (N_9100,N_8900,N_8681);
or U9101 (N_9101,N_8712,N_8934);
nand U9102 (N_9102,N_7984,N_7539);
and U9103 (N_9103,N_8038,N_8224);
and U9104 (N_9104,N_7610,N_8543);
or U9105 (N_9105,N_8530,N_7502);
or U9106 (N_9106,N_8416,N_7687);
and U9107 (N_9107,N_8589,N_8526);
nor U9108 (N_9108,N_8965,N_8953);
or U9109 (N_9109,N_8789,N_8309);
nand U9110 (N_9110,N_8275,N_8272);
nor U9111 (N_9111,N_7973,N_7571);
xor U9112 (N_9112,N_7830,N_8846);
or U9113 (N_9113,N_8199,N_8568);
and U9114 (N_9114,N_7645,N_8556);
nand U9115 (N_9115,N_8686,N_7927);
nand U9116 (N_9116,N_8245,N_7977);
nor U9117 (N_9117,N_8017,N_8174);
nand U9118 (N_9118,N_8217,N_8236);
nand U9119 (N_9119,N_8119,N_8860);
nor U9120 (N_9120,N_8664,N_7925);
nand U9121 (N_9121,N_8779,N_8672);
nor U9122 (N_9122,N_8075,N_8080);
nand U9123 (N_9123,N_8710,N_8052);
nand U9124 (N_9124,N_8393,N_7913);
nand U9125 (N_9125,N_8106,N_8111);
or U9126 (N_9126,N_7768,N_8661);
nand U9127 (N_9127,N_8457,N_8428);
or U9128 (N_9128,N_7652,N_7863);
or U9129 (N_9129,N_8273,N_7994);
and U9130 (N_9130,N_8930,N_8109);
and U9131 (N_9131,N_7910,N_8190);
nand U9132 (N_9132,N_8371,N_7594);
or U9133 (N_9133,N_7512,N_8582);
and U9134 (N_9134,N_7563,N_8094);
and U9135 (N_9135,N_8757,N_7718);
and U9136 (N_9136,N_7951,N_7922);
nor U9137 (N_9137,N_7771,N_8668);
nor U9138 (N_9138,N_7789,N_8074);
or U9139 (N_9139,N_8714,N_8870);
nor U9140 (N_9140,N_8225,N_7794);
or U9141 (N_9141,N_7755,N_8619);
or U9142 (N_9142,N_8448,N_8172);
nand U9143 (N_9143,N_7826,N_7828);
nor U9144 (N_9144,N_7967,N_8606);
nand U9145 (N_9145,N_8764,N_7800);
nand U9146 (N_9146,N_7624,N_8925);
and U9147 (N_9147,N_8991,N_7627);
nor U9148 (N_9148,N_8102,N_7938);
nor U9149 (N_9149,N_8042,N_7982);
nor U9150 (N_9150,N_8948,N_8579);
and U9151 (N_9151,N_7597,N_8340);
xnor U9152 (N_9152,N_8665,N_8995);
nand U9153 (N_9153,N_8180,N_8228);
and U9154 (N_9154,N_7527,N_8193);
nor U9155 (N_9155,N_8977,N_7787);
or U9156 (N_9156,N_7598,N_8352);
nand U9157 (N_9157,N_7947,N_8358);
and U9158 (N_9158,N_8051,N_7891);
nand U9159 (N_9159,N_8585,N_8308);
xor U9160 (N_9160,N_8071,N_8586);
nand U9161 (N_9161,N_8744,N_7798);
nor U9162 (N_9162,N_7778,N_8477);
and U9163 (N_9163,N_8214,N_7924);
or U9164 (N_9164,N_7625,N_7862);
or U9165 (N_9165,N_7660,N_7887);
and U9166 (N_9166,N_8797,N_7556);
nand U9167 (N_9167,N_8291,N_8219);
and U9168 (N_9168,N_8670,N_7520);
nand U9169 (N_9169,N_7934,N_8780);
and U9170 (N_9170,N_7953,N_8445);
and U9171 (N_9171,N_8226,N_8460);
nor U9172 (N_9172,N_8982,N_8547);
nand U9173 (N_9173,N_7564,N_7847);
or U9174 (N_9174,N_8025,N_8527);
nor U9175 (N_9175,N_8791,N_8629);
and U9176 (N_9176,N_8367,N_7985);
nand U9177 (N_9177,N_8330,N_8667);
nor U9178 (N_9178,N_8705,N_8739);
nand U9179 (N_9179,N_8561,N_8316);
or U9180 (N_9180,N_7983,N_8647);
and U9181 (N_9181,N_7543,N_8023);
or U9182 (N_9182,N_8867,N_8615);
or U9183 (N_9183,N_8198,N_8021);
nand U9184 (N_9184,N_8857,N_7851);
nand U9185 (N_9185,N_8104,N_8907);
and U9186 (N_9186,N_8508,N_8775);
or U9187 (N_9187,N_8999,N_8150);
nand U9188 (N_9188,N_8379,N_7686);
or U9189 (N_9189,N_8053,N_8824);
nand U9190 (N_9190,N_8260,N_7711);
nor U9191 (N_9191,N_7503,N_8064);
xor U9192 (N_9192,N_7683,N_7892);
and U9193 (N_9193,N_8163,N_7767);
nand U9194 (N_9194,N_8429,N_8105);
nor U9195 (N_9195,N_8821,N_8356);
or U9196 (N_9196,N_8959,N_7650);
or U9197 (N_9197,N_8913,N_8420);
or U9198 (N_9198,N_7810,N_8045);
and U9199 (N_9199,N_8142,N_8189);
nand U9200 (N_9200,N_8928,N_8363);
nand U9201 (N_9201,N_7867,N_7860);
nand U9202 (N_9202,N_8830,N_8171);
or U9203 (N_9203,N_8040,N_7861);
nor U9204 (N_9204,N_7595,N_7661);
and U9205 (N_9205,N_8899,N_8801);
nor U9206 (N_9206,N_8637,N_8265);
nor U9207 (N_9207,N_8546,N_8926);
and U9208 (N_9208,N_7791,N_8084);
and U9209 (N_9209,N_8317,N_7825);
nand U9210 (N_9210,N_8056,N_8360);
nand U9211 (N_9211,N_8516,N_7620);
nand U9212 (N_9212,N_8259,N_8874);
nand U9213 (N_9213,N_7907,N_8464);
and U9214 (N_9214,N_7501,N_8044);
nand U9215 (N_9215,N_8749,N_8120);
nor U9216 (N_9216,N_8766,N_8122);
nor U9217 (N_9217,N_7647,N_8888);
nand U9218 (N_9218,N_7829,N_8160);
and U9219 (N_9219,N_8885,N_8041);
nor U9220 (N_9220,N_8920,N_7714);
nand U9221 (N_9221,N_8774,N_8609);
nand U9222 (N_9222,N_8069,N_8572);
xor U9223 (N_9223,N_8558,N_8376);
and U9224 (N_9224,N_7786,N_8325);
and U9225 (N_9225,N_7737,N_8157);
or U9226 (N_9226,N_8447,N_7715);
nand U9227 (N_9227,N_7996,N_8758);
and U9228 (N_9228,N_8283,N_7734);
nor U9229 (N_9229,N_7720,N_8840);
nand U9230 (N_9230,N_8737,N_7790);
nand U9231 (N_9231,N_8178,N_7510);
and U9232 (N_9232,N_8060,N_8357);
and U9233 (N_9233,N_8232,N_8454);
nor U9234 (N_9234,N_7876,N_8183);
nor U9235 (N_9235,N_8509,N_7701);
nor U9236 (N_9236,N_8614,N_7721);
and U9237 (N_9237,N_8834,N_8897);
nand U9238 (N_9238,N_7773,N_8573);
nor U9239 (N_9239,N_7665,N_8481);
nor U9240 (N_9240,N_8716,N_8782);
and U9241 (N_9241,N_7975,N_7820);
nand U9242 (N_9242,N_8506,N_8603);
or U9243 (N_9243,N_7955,N_8673);
xnor U9244 (N_9244,N_8810,N_7500);
or U9245 (N_9245,N_8144,N_8989);
or U9246 (N_9246,N_7509,N_8221);
nor U9247 (N_9247,N_8583,N_8631);
nor U9248 (N_9248,N_7739,N_7582);
nor U9249 (N_9249,N_8007,N_8022);
nor U9250 (N_9250,N_8306,N_8008);
nand U9251 (N_9251,N_8628,N_7591);
nor U9252 (N_9252,N_8574,N_7602);
and U9253 (N_9253,N_8878,N_8845);
and U9254 (N_9254,N_7588,N_8320);
and U9255 (N_9255,N_7999,N_7870);
nor U9256 (N_9256,N_7926,N_8895);
nor U9257 (N_9257,N_8945,N_7762);
nor U9258 (N_9258,N_8931,N_8336);
and U9259 (N_9259,N_8450,N_7654);
nor U9260 (N_9260,N_7929,N_8649);
or U9261 (N_9261,N_8842,N_8808);
xnor U9262 (N_9262,N_8347,N_7842);
and U9263 (N_9263,N_8803,N_8242);
nand U9264 (N_9264,N_8533,N_7528);
nor U9265 (N_9265,N_8398,N_7705);
nand U9266 (N_9266,N_8315,N_8656);
and U9267 (N_9267,N_8331,N_8605);
or U9268 (N_9268,N_8415,N_8400);
and U9269 (N_9269,N_8851,N_7633);
nor U9270 (N_9270,N_8602,N_8388);
and U9271 (N_9271,N_8638,N_8727);
or U9272 (N_9272,N_8996,N_8921);
or U9273 (N_9273,N_8669,N_7848);
or U9274 (N_9274,N_8564,N_8184);
nand U9275 (N_9275,N_7526,N_8762);
and U9276 (N_9276,N_8255,N_7615);
and U9277 (N_9277,N_8029,N_8277);
nor U9278 (N_9278,N_8984,N_8252);
or U9279 (N_9279,N_8501,N_8544);
nand U9280 (N_9280,N_7717,N_8873);
or U9281 (N_9281,N_8792,N_8004);
nand U9282 (N_9282,N_8635,N_7630);
nor U9283 (N_9283,N_8034,N_7915);
or U9284 (N_9284,N_8731,N_8847);
or U9285 (N_9285,N_8825,N_7893);
or U9286 (N_9286,N_7916,N_8478);
and U9287 (N_9287,N_7560,N_8295);
or U9288 (N_9288,N_8537,N_8539);
nand U9289 (N_9289,N_7517,N_7747);
or U9290 (N_9290,N_7854,N_8186);
nand U9291 (N_9291,N_8612,N_8886);
or U9292 (N_9292,N_8055,N_7749);
and U9293 (N_9293,N_8704,N_7693);
nor U9294 (N_9294,N_8438,N_7894);
nor U9295 (N_9295,N_8729,N_8078);
nor U9296 (N_9296,N_7516,N_8473);
nor U9297 (N_9297,N_7751,N_8690);
nor U9298 (N_9298,N_8625,N_7834);
nor U9299 (N_9299,N_8132,N_8659);
or U9300 (N_9300,N_8310,N_7882);
or U9301 (N_9301,N_8422,N_7884);
nand U9302 (N_9302,N_8327,N_7575);
nand U9303 (N_9303,N_8451,N_8397);
xor U9304 (N_9304,N_7997,N_7757);
nand U9305 (N_9305,N_7580,N_8655);
nor U9306 (N_9306,N_7552,N_8682);
nor U9307 (N_9307,N_8191,N_8103);
or U9308 (N_9308,N_7764,N_8648);
xnor U9309 (N_9309,N_8086,N_8520);
or U9310 (N_9310,N_8335,N_8061);
and U9311 (N_9311,N_7655,N_8462);
nand U9312 (N_9312,N_8875,N_7710);
nor U9313 (N_9313,N_8693,N_8455);
and U9314 (N_9314,N_7682,N_8567);
xnor U9315 (N_9315,N_8597,N_8175);
or U9316 (N_9316,N_7704,N_7609);
nand U9317 (N_9317,N_8427,N_7616);
nor U9318 (N_9318,N_7850,N_7899);
nor U9319 (N_9319,N_7607,N_7869);
or U9320 (N_9320,N_7783,N_8707);
nand U9321 (N_9321,N_7671,N_7974);
and U9322 (N_9322,N_7648,N_8047);
and U9323 (N_9323,N_8253,N_8752);
nor U9324 (N_9324,N_8584,N_8257);
nor U9325 (N_9325,N_7756,N_8522);
nand U9326 (N_9326,N_7877,N_7752);
or U9327 (N_9327,N_7653,N_8679);
or U9328 (N_9328,N_7742,N_8702);
nor U9329 (N_9329,N_8196,N_8569);
or U9330 (N_9330,N_8903,N_8121);
or U9331 (N_9331,N_8777,N_8662);
nand U9332 (N_9332,N_8818,N_7827);
or U9333 (N_9333,N_7506,N_8389);
and U9334 (N_9334,N_8786,N_7840);
nand U9335 (N_9335,N_8819,N_8426);
or U9336 (N_9336,N_7628,N_8923);
or U9337 (N_9337,N_7838,N_8093);
nor U9338 (N_9338,N_8307,N_8639);
nand U9339 (N_9339,N_8550,N_7917);
xor U9340 (N_9340,N_8098,N_8964);
and U9341 (N_9341,N_8800,N_8954);
nand U9342 (N_9342,N_8399,N_8479);
and U9343 (N_9343,N_7638,N_8222);
and U9344 (N_9344,N_8804,N_8431);
nand U9345 (N_9345,N_8552,N_8169);
nor U9346 (N_9346,N_8554,N_7868);
nand U9347 (N_9347,N_7921,N_7681);
nand U9348 (N_9348,N_8298,N_8811);
nand U9349 (N_9349,N_8215,N_8973);
nand U9350 (N_9350,N_8290,N_7675);
nor U9351 (N_9351,N_7763,N_8708);
nor U9352 (N_9352,N_8529,N_7741);
nand U9353 (N_9353,N_7781,N_8014);
and U9354 (N_9354,N_7513,N_8092);
and U9355 (N_9355,N_8262,N_8849);
nand U9356 (N_9356,N_8244,N_7935);
nand U9357 (N_9357,N_8532,N_8936);
nor U9358 (N_9358,N_8570,N_8200);
nor U9359 (N_9359,N_8167,N_8381);
nand U9360 (N_9360,N_8364,N_7605);
nand U9361 (N_9361,N_8322,N_7815);
or U9362 (N_9362,N_8161,N_7803);
nor U9363 (N_9363,N_8489,N_7519);
and U9364 (N_9364,N_8684,N_8391);
nor U9365 (N_9365,N_8441,N_7601);
nor U9366 (N_9366,N_8565,N_8929);
nor U9367 (N_9367,N_7923,N_8844);
or U9368 (N_9368,N_8750,N_7736);
or U9369 (N_9369,N_8282,N_8862);
nand U9370 (N_9370,N_8692,N_8559);
or U9371 (N_9371,N_7809,N_7634);
nor U9372 (N_9372,N_7535,N_7538);
nand U9373 (N_9373,N_8778,N_8100);
and U9374 (N_9374,N_8496,N_8858);
and U9375 (N_9375,N_7919,N_8937);
nor U9376 (N_9376,N_7641,N_7593);
and U9377 (N_9377,N_8205,N_8576);
and U9378 (N_9378,N_7579,N_8299);
and U9379 (N_9379,N_7546,N_7962);
nand U9380 (N_9380,N_8442,N_8227);
or U9381 (N_9381,N_7626,N_8753);
nor U9382 (N_9382,N_8026,N_8024);
nand U9383 (N_9383,N_8536,N_7801);
nand U9384 (N_9384,N_8206,N_8696);
or U9385 (N_9385,N_7724,N_8591);
or U9386 (N_9386,N_7530,N_8620);
nor U9387 (N_9387,N_8468,N_8091);
xor U9388 (N_9388,N_8137,N_7670);
nand U9389 (N_9389,N_7900,N_8812);
nand U9390 (N_9390,N_8037,N_8054);
nand U9391 (N_9391,N_7590,N_8233);
nand U9392 (N_9392,N_7769,N_7566);
nor U9393 (N_9393,N_8213,N_7586);
or U9394 (N_9394,N_8145,N_8297);
nand U9395 (N_9395,N_8850,N_7732);
nor U9396 (N_9396,N_8300,N_8820);
and U9397 (N_9397,N_8642,N_8645);
and U9398 (N_9398,N_8831,N_8209);
and U9399 (N_9399,N_7855,N_8577);
or U9400 (N_9400,N_8433,N_7902);
nor U9401 (N_9401,N_8555,N_8793);
nand U9402 (N_9402,N_7574,N_7845);
nand U9403 (N_9403,N_8768,N_8168);
or U9404 (N_9404,N_8986,N_7875);
nor U9405 (N_9405,N_8611,N_8880);
nor U9406 (N_9406,N_7587,N_8285);
or U9407 (N_9407,N_8404,N_7753);
nand U9408 (N_9408,N_8019,N_7695);
or U9409 (N_9409,N_8301,N_7708);
xnor U9410 (N_9410,N_8378,N_8743);
and U9411 (N_9411,N_8049,N_8599);
nor U9412 (N_9412,N_8313,N_7991);
and U9413 (N_9413,N_7666,N_8414);
nand U9414 (N_9414,N_8268,N_8838);
and U9415 (N_9415,N_8798,N_8270);
nand U9416 (N_9416,N_7599,N_7635);
xnor U9417 (N_9417,N_8833,N_8238);
nor U9418 (N_9418,N_8904,N_7551);
nor U9419 (N_9419,N_7981,N_7966);
nand U9420 (N_9420,N_8274,N_8514);
nand U9421 (N_9421,N_8523,N_8646);
nor U9422 (N_9422,N_8070,N_8884);
xor U9423 (N_9423,N_8861,N_7897);
and U9424 (N_9424,N_7657,N_7822);
and U9425 (N_9425,N_7971,N_8288);
nand U9426 (N_9426,N_8202,N_8353);
nand U9427 (N_9427,N_7905,N_7978);
nor U9428 (N_9428,N_7568,N_8733);
or U9429 (N_9429,N_7703,N_7818);
nor U9430 (N_9430,N_8562,N_7954);
nor U9431 (N_9431,N_7697,N_8976);
nand U9432 (N_9432,N_8815,N_8967);
nor U9433 (N_9433,N_8018,N_8835);
or U9434 (N_9434,N_8970,N_8341);
and U9435 (N_9435,N_7976,N_7722);
nand U9436 (N_9436,N_7735,N_8115);
nand U9437 (N_9437,N_8730,N_7776);
xor U9438 (N_9438,N_8685,N_8177);
nor U9439 (N_9439,N_8891,N_7632);
or U9440 (N_9440,N_7550,N_8413);
or U9441 (N_9441,N_8557,N_7987);
and U9442 (N_9442,N_8158,N_8039);
nand U9443 (N_9443,N_7614,N_7631);
nand U9444 (N_9444,N_8836,N_8841);
and U9445 (N_9445,N_8342,N_7532);
nor U9446 (N_9446,N_8294,N_8355);
nor U9447 (N_9447,N_7772,N_8033);
nor U9448 (N_9448,N_8763,N_8595);
and U9449 (N_9449,N_8240,N_7523);
and U9450 (N_9450,N_8264,N_7567);
nand U9451 (N_9451,N_8571,N_8974);
and U9452 (N_9452,N_8254,N_7903);
nor U9453 (N_9453,N_8521,N_8601);
and U9454 (N_9454,N_8963,N_7585);
and U9455 (N_9455,N_8689,N_7866);
nand U9456 (N_9456,N_8700,N_8146);
or U9457 (N_9457,N_8652,N_8940);
or U9458 (N_9458,N_8794,N_8864);
nand U9459 (N_9459,N_7643,N_8852);
and U9460 (N_9460,N_7972,N_7672);
or U9461 (N_9461,N_8484,N_7688);
and U9462 (N_9462,N_8869,N_7529);
nor U9463 (N_9463,N_8333,N_7960);
xnor U9464 (N_9464,N_8553,N_7814);
and U9465 (N_9465,N_8293,N_7515);
nor U9466 (N_9466,N_8916,N_8944);
or U9467 (N_9467,N_7980,N_8592);
nor U9468 (N_9468,N_8487,N_7782);
nand U9469 (N_9469,N_8896,N_7541);
nand U9470 (N_9470,N_8095,N_8359);
or U9471 (N_9471,N_7669,N_8089);
and U9472 (N_9472,N_7859,N_8020);
nor U9473 (N_9473,N_8859,N_8469);
or U9474 (N_9474,N_7992,N_8012);
or U9475 (N_9475,N_8587,N_7878);
nand U9476 (N_9476,N_8790,N_8031);
or U9477 (N_9477,N_7957,N_7888);
and U9478 (N_9478,N_8745,N_8384);
nor U9479 (N_9479,N_8997,N_8776);
nor U9480 (N_9480,N_8491,N_8062);
nor U9481 (N_9481,N_8204,N_7961);
nor U9482 (N_9482,N_7895,N_8154);
nor U9483 (N_9483,N_8382,N_8418);
nor U9484 (N_9484,N_8361,N_8946);
nor U9485 (N_9485,N_8406,N_7969);
and U9486 (N_9486,N_8077,N_8868);
nand U9487 (N_9487,N_8541,N_8396);
nor U9488 (N_9488,N_7511,N_8877);
nand U9489 (N_9489,N_8754,N_8337);
and U9490 (N_9490,N_7604,N_8632);
and U9491 (N_9491,N_8678,N_8785);
xnor U9492 (N_9492,N_8992,N_8660);
or U9493 (N_9493,N_7788,N_7694);
and U9494 (N_9494,N_8097,N_8701);
or U9495 (N_9495,N_8680,N_8876);
nand U9496 (N_9496,N_7537,N_8090);
or U9497 (N_9497,N_7808,N_7728);
nand U9498 (N_9498,N_7879,N_7522);
nor U9499 (N_9499,N_8947,N_7831);
and U9500 (N_9500,N_8181,N_8278);
nand U9501 (N_9501,N_8598,N_7785);
nand U9502 (N_9502,N_8405,N_8495);
nand U9503 (N_9503,N_8806,N_8542);
and U9504 (N_9504,N_8149,N_7766);
nor U9505 (N_9505,N_8140,N_8742);
nand U9506 (N_9506,N_7578,N_7759);
nand U9507 (N_9507,N_8235,N_8370);
nor U9508 (N_9508,N_7805,N_7792);
or U9509 (N_9509,N_8651,N_7770);
nor U9510 (N_9510,N_8952,N_7821);
nor U9511 (N_9511,N_7873,N_8453);
or U9512 (N_9512,N_7819,N_8653);
or U9513 (N_9513,N_7780,N_8208);
and U9514 (N_9514,N_8814,N_8817);
nor U9515 (N_9515,N_8068,N_8362);
nand U9516 (N_9516,N_8476,N_8136);
and U9517 (N_9517,N_7849,N_8718);
or U9518 (N_9518,N_8302,N_8519);
nor U9519 (N_9519,N_7990,N_8048);
and U9520 (N_9520,N_7986,N_7760);
or U9521 (N_9521,N_8003,N_7911);
nand U9522 (N_9522,N_8694,N_8425);
or U9523 (N_9523,N_8773,N_7740);
nor U9524 (N_9524,N_8173,N_7824);
or U9525 (N_9525,N_8728,N_8305);
nand U9526 (N_9526,N_8912,N_8575);
xor U9527 (N_9527,N_8933,N_8459);
nand U9528 (N_9528,N_8593,N_8432);
nand U9529 (N_9529,N_8099,N_7761);
or U9530 (N_9530,N_8276,N_7896);
or U9531 (N_9531,N_7758,N_8258);
or U9532 (N_9532,N_7928,N_8578);
and U9533 (N_9533,N_7700,N_7745);
nor U9534 (N_9534,N_8720,N_7690);
or U9535 (N_9535,N_8230,N_8807);
or U9536 (N_9536,N_8640,N_7836);
nor U9537 (N_9537,N_8942,N_8493);
and U9538 (N_9538,N_7843,N_8630);
and U9539 (N_9539,N_8827,N_7583);
or U9540 (N_9540,N_7998,N_8286);
or U9541 (N_9541,N_8392,N_7559);
xor U9542 (N_9542,N_8813,N_7639);
nor U9543 (N_9543,N_8590,N_7837);
nor U9544 (N_9544,N_7874,N_8251);
nand U9545 (N_9545,N_8760,N_8671);
nand U9546 (N_9546,N_8463,N_7651);
or U9547 (N_9547,N_8164,N_7612);
nand U9548 (N_9548,N_7730,N_7706);
nand U9549 (N_9549,N_7797,N_8319);
nor U9550 (N_9550,N_8261,N_8165);
nor U9551 (N_9551,N_8403,N_8854);
and U9552 (N_9552,N_7558,N_8212);
or U9553 (N_9553,N_8410,N_8941);
nor U9554 (N_9554,N_8767,N_8889);
xor U9555 (N_9555,N_7858,N_8153);
or U9556 (N_9556,N_8443,N_7793);
nand U9557 (N_9557,N_8435,N_8350);
or U9558 (N_9558,N_8354,N_8210);
or U9559 (N_9559,N_8005,N_8237);
nand U9560 (N_9560,N_8703,N_8124);
or U9561 (N_9561,N_8901,N_7750);
xor U9562 (N_9562,N_8321,N_8006);
and U9563 (N_9563,N_7569,N_8975);
nand U9564 (N_9564,N_8284,N_8141);
and U9565 (N_9565,N_8456,N_7514);
and U9566 (N_9566,N_8408,N_8467);
or U9567 (N_9567,N_8182,N_7508);
and U9568 (N_9568,N_8480,N_8924);
and U9569 (N_9569,N_8499,N_7617);
nand U9570 (N_9570,N_8263,N_7959);
nor U9571 (N_9571,N_8304,N_8229);
nand U9572 (N_9572,N_8594,N_8784);
and U9573 (N_9573,N_8510,N_8551);
nand U9574 (N_9574,N_8349,N_8466);
nand U9575 (N_9575,N_8581,N_8344);
nor U9576 (N_9576,N_8083,N_7979);
nor U9577 (N_9577,N_7833,N_7702);
and U9578 (N_9578,N_8616,N_8128);
or U9579 (N_9579,N_8517,N_8856);
and U9580 (N_9580,N_7871,N_8289);
or U9581 (N_9581,N_8822,N_8674);
and U9582 (N_9582,N_7944,N_8935);
or U9583 (N_9583,N_7949,N_8600);
xor U9584 (N_9584,N_7738,N_8866);
nor U9585 (N_9585,N_7562,N_8596);
nor U9586 (N_9586,N_8483,N_7534);
nor U9587 (N_9587,N_8914,N_8312);
and U9588 (N_9588,N_8343,N_8117);
nand U9589 (N_9589,N_8713,N_7596);
nor U9590 (N_9590,N_8981,N_8770);
and U9591 (N_9591,N_8893,N_8417);
nand U9592 (N_9592,N_7904,N_8207);
and U9593 (N_9593,N_8369,N_8741);
and U9594 (N_9594,N_8010,N_7995);
or U9595 (N_9595,N_8152,N_8627);
and U9596 (N_9596,N_8394,N_8633);
nor U9597 (N_9597,N_7841,N_7857);
and U9598 (N_9598,N_8449,N_8243);
or U9599 (N_9599,N_8279,N_8636);
nand U9600 (N_9600,N_8500,N_7813);
nand U9601 (N_9601,N_8983,N_7993);
nor U9602 (N_9602,N_7691,N_8375);
nand U9603 (N_9603,N_7795,N_8515);
nor U9604 (N_9604,N_7844,N_8409);
xor U9605 (N_9605,N_8534,N_8267);
and U9606 (N_9606,N_8043,N_8734);
nor U9607 (N_9607,N_7989,N_7731);
nand U9608 (N_9608,N_7505,N_8988);
nand U9609 (N_9609,N_8076,N_8528);
xnor U9610 (N_9610,N_7658,N_8176);
or U9611 (N_9611,N_8805,N_7727);
nor U9612 (N_9612,N_8799,N_8135);
and U9613 (N_9613,N_8719,N_8148);
and U9614 (N_9614,N_8082,N_7864);
and U9615 (N_9615,N_8747,N_8883);
or U9616 (N_9616,N_7941,N_7676);
or U9617 (N_9617,N_7547,N_8566);
nand U9618 (N_9618,N_8905,N_8956);
xor U9619 (N_9619,N_8657,N_8241);
or U9620 (N_9620,N_7521,N_7709);
or U9621 (N_9621,N_8761,N_8617);
and U9622 (N_9622,N_7637,N_8715);
and U9623 (N_9623,N_8740,N_8622);
or U9624 (N_9624,N_7746,N_7940);
or U9625 (N_9625,N_8138,N_7536);
and U9626 (N_9626,N_8796,N_8118);
and U9627 (N_9627,N_7719,N_8706);
nor U9628 (N_9628,N_8979,N_8504);
nor U9629 (N_9629,N_8372,N_8623);
nand U9630 (N_9630,N_8608,N_8016);
nand U9631 (N_9631,N_7584,N_7733);
nor U9632 (N_9632,N_8166,N_8338);
nand U9633 (N_9633,N_8535,N_8266);
nand U9634 (N_9634,N_7823,N_7886);
and U9635 (N_9635,N_8919,N_8437);
or U9636 (N_9636,N_8125,N_8756);
and U9637 (N_9637,N_7936,N_7555);
nor U9638 (N_9638,N_8088,N_8691);
nor U9639 (N_9639,N_8497,N_8492);
nor U9640 (N_9640,N_7852,N_7946);
xor U9641 (N_9641,N_7576,N_8015);
nor U9642 (N_9642,N_8194,N_8271);
and U9643 (N_9643,N_7577,N_8985);
nand U9644 (N_9644,N_8134,N_8604);
nor U9645 (N_9645,N_8197,N_8269);
or U9646 (N_9646,N_8709,N_8058);
and U9647 (N_9647,N_8486,N_8809);
nand U9648 (N_9648,N_7659,N_8292);
or U9649 (N_9649,N_8248,N_8239);
xnor U9650 (N_9650,N_7832,N_7689);
or U9651 (N_9651,N_7606,N_7912);
or U9652 (N_9652,N_8688,N_8951);
nand U9653 (N_9653,N_7518,N_8368);
nor U9654 (N_9654,N_7662,N_8910);
nor U9655 (N_9655,N_8187,N_7748);
and U9656 (N_9656,N_7644,N_8961);
nor U9657 (N_9657,N_8401,N_8863);
nand U9658 (N_9658,N_7525,N_8475);
nor U9659 (N_9659,N_8482,N_8155);
or U9660 (N_9660,N_7642,N_8311);
or U9661 (N_9661,N_8969,N_7799);
nor U9662 (N_9662,N_7883,N_8366);
and U9663 (N_9663,N_7856,N_8695);
or U9664 (N_9664,N_8823,N_8816);
or U9665 (N_9665,N_8955,N_8865);
nand U9666 (N_9666,N_8032,N_8748);
xnor U9667 (N_9667,N_7931,N_8721);
or U9668 (N_9668,N_8027,N_8067);
nand U9669 (N_9669,N_8971,N_7898);
and U9670 (N_9670,N_8531,N_7906);
nor U9671 (N_9671,N_7698,N_8421);
nor U9672 (N_9672,N_7507,N_8829);
and U9673 (N_9673,N_8065,N_8434);
or U9674 (N_9674,N_8011,N_8548);
nor U9675 (N_9675,N_7765,N_8390);
nand U9676 (N_9676,N_8826,N_8723);
nor U9677 (N_9677,N_8538,N_8918);
and U9678 (N_9678,N_8580,N_8419);
xor U9679 (N_9679,N_7592,N_8314);
and U9680 (N_9680,N_8545,N_7956);
nand U9681 (N_9681,N_7544,N_8030);
nand U9682 (N_9682,N_8511,N_8994);
or U9683 (N_9683,N_8588,N_8387);
nand U9684 (N_9684,N_8035,N_7613);
nand U9685 (N_9685,N_7930,N_8658);
nor U9686 (N_9686,N_8641,N_8498);
or U9687 (N_9687,N_8909,N_7554);
or U9688 (N_9688,N_8722,N_7804);
nand U9689 (N_9689,N_7839,N_8643);
and U9690 (N_9690,N_8223,N_8993);
nand U9691 (N_9691,N_7685,N_8759);
or U9692 (N_9692,N_8218,N_7968);
nand U9693 (N_9693,N_8129,N_7684);
xnor U9694 (N_9694,N_8472,N_7540);
nor U9695 (N_9695,N_8987,N_8112);
nand U9696 (N_9696,N_8246,N_8621);
xor U9697 (N_9697,N_8687,N_8513);
or U9698 (N_9698,N_7988,N_8746);
and U9699 (N_9699,N_8828,N_8755);
nor U9700 (N_9700,N_7725,N_7699);
and U9701 (N_9701,N_7914,N_8998);
or U9702 (N_9702,N_8143,N_8832);
nand U9703 (N_9703,N_8377,N_8185);
nand U9704 (N_9704,N_8922,N_7817);
nand U9705 (N_9705,N_8057,N_7674);
nor U9706 (N_9706,N_8490,N_7723);
nor U9707 (N_9707,N_8374,N_7835);
nand U9708 (N_9708,N_8339,N_8156);
or U9709 (N_9709,N_7779,N_8938);
nor U9710 (N_9710,N_8772,N_8085);
or U9711 (N_9711,N_7846,N_7970);
or U9712 (N_9712,N_7853,N_8050);
nand U9713 (N_9713,N_7679,N_8485);
xnor U9714 (N_9714,N_7621,N_7880);
or U9715 (N_9715,N_7775,N_8066);
nor U9716 (N_9716,N_8494,N_8000);
xor U9717 (N_9717,N_8147,N_8634);
and U9718 (N_9718,N_8781,N_8195);
and U9719 (N_9719,N_8318,N_8107);
and U9720 (N_9720,N_8732,N_8788);
or U9721 (N_9721,N_8540,N_8324);
nor U9722 (N_9722,N_8332,N_8783);
nand U9723 (N_9723,N_8296,N_7581);
or U9724 (N_9724,N_7726,N_8411);
nor U9725 (N_9725,N_8130,N_8968);
xnor U9726 (N_9726,N_8894,N_7713);
and U9727 (N_9727,N_8966,N_8887);
and U9728 (N_9728,N_8962,N_7716);
or U9729 (N_9729,N_7636,N_8231);
nand U9730 (N_9730,N_8114,N_8848);
nand U9731 (N_9731,N_7712,N_8101);
or U9732 (N_9732,N_7524,N_8013);
or U9733 (N_9733,N_8699,N_8787);
nand U9734 (N_9734,N_7950,N_7557);
and U9735 (N_9735,N_7619,N_8465);
nor U9736 (N_9736,N_7743,N_8471);
nor U9737 (N_9737,N_7918,N_8839);
and U9738 (N_9738,N_8474,N_8203);
or U9739 (N_9739,N_8452,N_8133);
or U9740 (N_9740,N_8001,N_8853);
nand U9741 (N_9741,N_8423,N_8675);
nand U9742 (N_9742,N_7531,N_8549);
xnor U9743 (N_9743,N_8162,N_8345);
and U9744 (N_9744,N_8110,N_8957);
nand U9745 (N_9745,N_8280,N_8351);
or U9746 (N_9746,N_8560,N_8654);
and U9747 (N_9747,N_8139,N_8524);
or U9748 (N_9748,N_7784,N_7549);
nor U9749 (N_9749,N_7909,N_7677);
and U9750 (N_9750,N_8423,N_8432);
nor U9751 (N_9751,N_7835,N_8336);
nand U9752 (N_9752,N_8023,N_8030);
or U9753 (N_9753,N_8015,N_8039);
and U9754 (N_9754,N_7646,N_7533);
nor U9755 (N_9755,N_8942,N_8135);
nor U9756 (N_9756,N_8117,N_8820);
and U9757 (N_9757,N_8724,N_7995);
nor U9758 (N_9758,N_8127,N_7642);
nor U9759 (N_9759,N_8219,N_8261);
xor U9760 (N_9760,N_8235,N_7994);
and U9761 (N_9761,N_8367,N_8221);
or U9762 (N_9762,N_8099,N_8583);
and U9763 (N_9763,N_8712,N_8093);
and U9764 (N_9764,N_8500,N_7739);
nor U9765 (N_9765,N_7824,N_8376);
and U9766 (N_9766,N_7929,N_8740);
nand U9767 (N_9767,N_8657,N_8352);
nor U9768 (N_9768,N_8481,N_8113);
nand U9769 (N_9769,N_7543,N_8193);
nand U9770 (N_9770,N_8844,N_8549);
nor U9771 (N_9771,N_8239,N_8186);
and U9772 (N_9772,N_8144,N_8176);
and U9773 (N_9773,N_8598,N_8387);
xnor U9774 (N_9774,N_8617,N_8514);
nor U9775 (N_9775,N_8424,N_8545);
nor U9776 (N_9776,N_8330,N_7647);
and U9777 (N_9777,N_8123,N_8988);
or U9778 (N_9778,N_7659,N_8229);
nor U9779 (N_9779,N_8311,N_7806);
nor U9780 (N_9780,N_8368,N_8173);
nand U9781 (N_9781,N_7555,N_7941);
nand U9782 (N_9782,N_8029,N_8853);
and U9783 (N_9783,N_8480,N_7747);
and U9784 (N_9784,N_7841,N_8639);
or U9785 (N_9785,N_8558,N_8439);
and U9786 (N_9786,N_8283,N_8196);
or U9787 (N_9787,N_8414,N_7557);
or U9788 (N_9788,N_8127,N_8037);
nand U9789 (N_9789,N_8871,N_7816);
and U9790 (N_9790,N_7974,N_8457);
nand U9791 (N_9791,N_8508,N_8924);
nor U9792 (N_9792,N_7547,N_7759);
and U9793 (N_9793,N_7614,N_8004);
nand U9794 (N_9794,N_8636,N_8079);
or U9795 (N_9795,N_8979,N_8506);
nor U9796 (N_9796,N_8575,N_7678);
or U9797 (N_9797,N_8310,N_7728);
nor U9798 (N_9798,N_7792,N_8724);
nor U9799 (N_9799,N_8878,N_8279);
nor U9800 (N_9800,N_8172,N_8525);
nand U9801 (N_9801,N_7700,N_7892);
and U9802 (N_9802,N_8363,N_8748);
or U9803 (N_9803,N_8644,N_8854);
xor U9804 (N_9804,N_7515,N_8839);
or U9805 (N_9805,N_7617,N_8796);
nand U9806 (N_9806,N_7698,N_8044);
or U9807 (N_9807,N_8686,N_7764);
nor U9808 (N_9808,N_8375,N_8161);
and U9809 (N_9809,N_7738,N_8101);
nand U9810 (N_9810,N_8572,N_8703);
and U9811 (N_9811,N_8201,N_7782);
nor U9812 (N_9812,N_8838,N_7585);
nand U9813 (N_9813,N_8886,N_8779);
nand U9814 (N_9814,N_7746,N_8008);
or U9815 (N_9815,N_8979,N_7997);
nand U9816 (N_9816,N_7601,N_8359);
nand U9817 (N_9817,N_8768,N_8030);
or U9818 (N_9818,N_7894,N_8753);
nor U9819 (N_9819,N_8035,N_7959);
and U9820 (N_9820,N_7620,N_8469);
nand U9821 (N_9821,N_8058,N_8296);
nor U9822 (N_9822,N_7620,N_8819);
and U9823 (N_9823,N_8520,N_8393);
nor U9824 (N_9824,N_7507,N_8974);
or U9825 (N_9825,N_8334,N_8954);
and U9826 (N_9826,N_8792,N_8331);
nor U9827 (N_9827,N_8115,N_8535);
nor U9828 (N_9828,N_8233,N_8767);
nand U9829 (N_9829,N_8405,N_8436);
nor U9830 (N_9830,N_7524,N_8292);
nor U9831 (N_9831,N_8208,N_7768);
or U9832 (N_9832,N_8107,N_7660);
and U9833 (N_9833,N_8913,N_8243);
and U9834 (N_9834,N_8486,N_8140);
nand U9835 (N_9835,N_8654,N_7990);
nor U9836 (N_9836,N_8756,N_7992);
nor U9837 (N_9837,N_8170,N_8156);
nor U9838 (N_9838,N_7931,N_8334);
or U9839 (N_9839,N_8384,N_8564);
nor U9840 (N_9840,N_8716,N_8823);
and U9841 (N_9841,N_8373,N_8115);
nor U9842 (N_9842,N_8957,N_7762);
nand U9843 (N_9843,N_7845,N_7520);
and U9844 (N_9844,N_7523,N_8249);
or U9845 (N_9845,N_8771,N_8961);
nand U9846 (N_9846,N_8670,N_7607);
nand U9847 (N_9847,N_7694,N_7639);
and U9848 (N_9848,N_7689,N_8359);
nor U9849 (N_9849,N_8504,N_8134);
or U9850 (N_9850,N_8457,N_8894);
or U9851 (N_9851,N_8009,N_8578);
and U9852 (N_9852,N_7777,N_8701);
xor U9853 (N_9853,N_8806,N_7905);
and U9854 (N_9854,N_7952,N_8494);
nand U9855 (N_9855,N_8212,N_8639);
nor U9856 (N_9856,N_8996,N_8503);
and U9857 (N_9857,N_8271,N_7758);
nand U9858 (N_9858,N_7635,N_7837);
nand U9859 (N_9859,N_7596,N_7751);
and U9860 (N_9860,N_8945,N_8805);
and U9861 (N_9861,N_8868,N_8558);
nand U9862 (N_9862,N_8473,N_8096);
nand U9863 (N_9863,N_7540,N_7518);
or U9864 (N_9864,N_8942,N_8937);
nor U9865 (N_9865,N_8496,N_8348);
xnor U9866 (N_9866,N_7670,N_8547);
nor U9867 (N_9867,N_8669,N_8620);
nand U9868 (N_9868,N_8104,N_8362);
or U9869 (N_9869,N_8688,N_8424);
nor U9870 (N_9870,N_7852,N_8476);
or U9871 (N_9871,N_8718,N_8116);
or U9872 (N_9872,N_7679,N_8989);
nand U9873 (N_9873,N_7752,N_8974);
nand U9874 (N_9874,N_8773,N_7575);
nor U9875 (N_9875,N_8510,N_7744);
or U9876 (N_9876,N_7742,N_7509);
nor U9877 (N_9877,N_8822,N_8484);
or U9878 (N_9878,N_8788,N_8454);
nand U9879 (N_9879,N_8047,N_7522);
nor U9880 (N_9880,N_8762,N_7845);
and U9881 (N_9881,N_7934,N_8734);
or U9882 (N_9882,N_8878,N_8716);
and U9883 (N_9883,N_8457,N_8750);
or U9884 (N_9884,N_8917,N_8925);
nor U9885 (N_9885,N_8184,N_7548);
nand U9886 (N_9886,N_8311,N_7940);
or U9887 (N_9887,N_7524,N_7909);
and U9888 (N_9888,N_8721,N_8152);
and U9889 (N_9889,N_7575,N_8210);
nor U9890 (N_9890,N_7882,N_8979);
or U9891 (N_9891,N_8213,N_8752);
nor U9892 (N_9892,N_8128,N_7719);
or U9893 (N_9893,N_8866,N_8728);
and U9894 (N_9894,N_8806,N_7611);
and U9895 (N_9895,N_8030,N_7679);
nor U9896 (N_9896,N_8931,N_7861);
and U9897 (N_9897,N_8608,N_7831);
nand U9898 (N_9898,N_8462,N_8996);
or U9899 (N_9899,N_8758,N_8621);
nor U9900 (N_9900,N_8869,N_8080);
nand U9901 (N_9901,N_8553,N_8852);
or U9902 (N_9902,N_8139,N_8074);
and U9903 (N_9903,N_7917,N_8724);
xnor U9904 (N_9904,N_8213,N_7509);
or U9905 (N_9905,N_8692,N_8320);
or U9906 (N_9906,N_7542,N_8274);
nand U9907 (N_9907,N_7925,N_8851);
nand U9908 (N_9908,N_7994,N_8699);
nor U9909 (N_9909,N_7865,N_7764);
nor U9910 (N_9910,N_8103,N_7949);
or U9911 (N_9911,N_7986,N_8245);
nand U9912 (N_9912,N_7892,N_8555);
and U9913 (N_9913,N_7981,N_7982);
nor U9914 (N_9914,N_8813,N_8203);
or U9915 (N_9915,N_8172,N_8441);
or U9916 (N_9916,N_7551,N_8796);
nor U9917 (N_9917,N_8827,N_8672);
or U9918 (N_9918,N_8694,N_8734);
nor U9919 (N_9919,N_8781,N_7560);
xnor U9920 (N_9920,N_7838,N_8496);
nor U9921 (N_9921,N_8392,N_7796);
and U9922 (N_9922,N_8350,N_8640);
and U9923 (N_9923,N_8547,N_8028);
and U9924 (N_9924,N_8089,N_8523);
and U9925 (N_9925,N_7658,N_8712);
or U9926 (N_9926,N_8242,N_8376);
nand U9927 (N_9927,N_8892,N_8977);
nor U9928 (N_9928,N_8039,N_7932);
nor U9929 (N_9929,N_8485,N_8812);
xnor U9930 (N_9930,N_8466,N_8399);
and U9931 (N_9931,N_8308,N_8303);
and U9932 (N_9932,N_8669,N_8977);
and U9933 (N_9933,N_7813,N_7580);
or U9934 (N_9934,N_8999,N_7623);
nand U9935 (N_9935,N_8984,N_8207);
or U9936 (N_9936,N_7800,N_7761);
nand U9937 (N_9937,N_8025,N_7876);
and U9938 (N_9938,N_8669,N_8649);
nor U9939 (N_9939,N_7730,N_8062);
nand U9940 (N_9940,N_7738,N_8487);
or U9941 (N_9941,N_8958,N_8420);
nand U9942 (N_9942,N_8465,N_8133);
nand U9943 (N_9943,N_8073,N_7937);
nand U9944 (N_9944,N_7895,N_7535);
or U9945 (N_9945,N_8816,N_8745);
and U9946 (N_9946,N_7734,N_8828);
nor U9947 (N_9947,N_7749,N_7867);
or U9948 (N_9948,N_8986,N_7853);
or U9949 (N_9949,N_8514,N_8844);
nor U9950 (N_9950,N_8582,N_7716);
and U9951 (N_9951,N_8167,N_7515);
nand U9952 (N_9952,N_8712,N_7630);
and U9953 (N_9953,N_8891,N_7624);
nand U9954 (N_9954,N_8151,N_8165);
nand U9955 (N_9955,N_8016,N_8220);
nor U9956 (N_9956,N_8396,N_7526);
and U9957 (N_9957,N_7781,N_7954);
or U9958 (N_9958,N_8955,N_8474);
nor U9959 (N_9959,N_7945,N_7626);
nor U9960 (N_9960,N_8081,N_8290);
and U9961 (N_9961,N_8845,N_8547);
or U9962 (N_9962,N_8072,N_8464);
nand U9963 (N_9963,N_7575,N_8906);
nand U9964 (N_9964,N_8929,N_8342);
or U9965 (N_9965,N_7642,N_8207);
and U9966 (N_9966,N_8179,N_8137);
nor U9967 (N_9967,N_8373,N_8649);
nor U9968 (N_9968,N_8217,N_8301);
nor U9969 (N_9969,N_8400,N_7882);
nand U9970 (N_9970,N_8090,N_8852);
nand U9971 (N_9971,N_7913,N_8179);
nand U9972 (N_9972,N_8397,N_8179);
nand U9973 (N_9973,N_8783,N_7990);
or U9974 (N_9974,N_7963,N_8016);
nor U9975 (N_9975,N_8714,N_8217);
or U9976 (N_9976,N_8048,N_8503);
nor U9977 (N_9977,N_8332,N_8372);
nand U9978 (N_9978,N_8779,N_7624);
nand U9979 (N_9979,N_8428,N_8662);
and U9980 (N_9980,N_8298,N_8526);
nor U9981 (N_9981,N_8356,N_8482);
nand U9982 (N_9982,N_8340,N_8232);
nor U9983 (N_9983,N_7788,N_8480);
nand U9984 (N_9984,N_8382,N_8836);
nand U9985 (N_9985,N_8695,N_8047);
and U9986 (N_9986,N_8506,N_8099);
nor U9987 (N_9987,N_8117,N_8295);
or U9988 (N_9988,N_8011,N_8868);
and U9989 (N_9989,N_8401,N_7873);
nor U9990 (N_9990,N_8884,N_7913);
and U9991 (N_9991,N_7910,N_8483);
nor U9992 (N_9992,N_8178,N_8777);
or U9993 (N_9993,N_8577,N_7584);
nor U9994 (N_9994,N_8042,N_8697);
or U9995 (N_9995,N_7769,N_8132);
and U9996 (N_9996,N_8615,N_8486);
nand U9997 (N_9997,N_7588,N_8373);
and U9998 (N_9998,N_7933,N_8604);
nor U9999 (N_9999,N_7751,N_7630);
nor U10000 (N_10000,N_8692,N_8167);
nor U10001 (N_10001,N_8050,N_8289);
nand U10002 (N_10002,N_8798,N_8309);
nor U10003 (N_10003,N_8402,N_8493);
nor U10004 (N_10004,N_7692,N_7557);
nor U10005 (N_10005,N_8442,N_8707);
xor U10006 (N_10006,N_7943,N_8859);
nand U10007 (N_10007,N_7616,N_8989);
nand U10008 (N_10008,N_7733,N_7677);
or U10009 (N_10009,N_8037,N_8477);
nand U10010 (N_10010,N_7783,N_8836);
or U10011 (N_10011,N_8014,N_7766);
and U10012 (N_10012,N_7626,N_8313);
and U10013 (N_10013,N_8383,N_7621);
or U10014 (N_10014,N_8918,N_7721);
and U10015 (N_10015,N_7991,N_7948);
and U10016 (N_10016,N_7832,N_8464);
or U10017 (N_10017,N_7790,N_7597);
nor U10018 (N_10018,N_8650,N_7573);
or U10019 (N_10019,N_7585,N_8794);
nand U10020 (N_10020,N_7891,N_8932);
nand U10021 (N_10021,N_7610,N_7767);
and U10022 (N_10022,N_8649,N_8600);
nand U10023 (N_10023,N_8346,N_8047);
nor U10024 (N_10024,N_8045,N_8221);
nor U10025 (N_10025,N_8078,N_7758);
or U10026 (N_10026,N_8394,N_8485);
nor U10027 (N_10027,N_7882,N_8121);
xor U10028 (N_10028,N_8573,N_7869);
and U10029 (N_10029,N_8520,N_7638);
or U10030 (N_10030,N_7823,N_7694);
and U10031 (N_10031,N_8376,N_8385);
or U10032 (N_10032,N_8619,N_8280);
nand U10033 (N_10033,N_8828,N_7793);
and U10034 (N_10034,N_8452,N_8191);
or U10035 (N_10035,N_8517,N_8455);
and U10036 (N_10036,N_8412,N_8504);
nor U10037 (N_10037,N_7516,N_8831);
and U10038 (N_10038,N_8647,N_7568);
nand U10039 (N_10039,N_8668,N_8870);
and U10040 (N_10040,N_8627,N_8708);
nor U10041 (N_10041,N_8138,N_8895);
nor U10042 (N_10042,N_8578,N_7701);
or U10043 (N_10043,N_8031,N_7517);
nand U10044 (N_10044,N_7886,N_7551);
or U10045 (N_10045,N_8292,N_8530);
nor U10046 (N_10046,N_7645,N_7630);
or U10047 (N_10047,N_8419,N_8687);
nand U10048 (N_10048,N_8310,N_8911);
nor U10049 (N_10049,N_8770,N_8220);
or U10050 (N_10050,N_7890,N_7867);
nor U10051 (N_10051,N_8804,N_7824);
nand U10052 (N_10052,N_8559,N_8655);
nand U10053 (N_10053,N_8852,N_8998);
and U10054 (N_10054,N_7706,N_8779);
nand U10055 (N_10055,N_8469,N_7797);
nor U10056 (N_10056,N_8552,N_8028);
nor U10057 (N_10057,N_8612,N_7708);
or U10058 (N_10058,N_7683,N_7871);
nand U10059 (N_10059,N_8028,N_7765);
nor U10060 (N_10060,N_7547,N_8143);
or U10061 (N_10061,N_8944,N_8138);
nand U10062 (N_10062,N_8116,N_7872);
nand U10063 (N_10063,N_8205,N_8032);
xnor U10064 (N_10064,N_8039,N_8315);
nor U10065 (N_10065,N_8999,N_8587);
or U10066 (N_10066,N_8392,N_7840);
nand U10067 (N_10067,N_8811,N_7700);
nor U10068 (N_10068,N_8061,N_7660);
nand U10069 (N_10069,N_7802,N_8871);
nand U10070 (N_10070,N_8887,N_8604);
and U10071 (N_10071,N_7841,N_8030);
or U10072 (N_10072,N_7783,N_8853);
nand U10073 (N_10073,N_7693,N_7749);
and U10074 (N_10074,N_8626,N_8090);
or U10075 (N_10075,N_7828,N_7625);
and U10076 (N_10076,N_8202,N_8581);
nor U10077 (N_10077,N_8454,N_8652);
or U10078 (N_10078,N_8458,N_8669);
and U10079 (N_10079,N_8744,N_8747);
nor U10080 (N_10080,N_8598,N_8374);
nor U10081 (N_10081,N_8836,N_7640);
or U10082 (N_10082,N_8343,N_8602);
nor U10083 (N_10083,N_7838,N_8097);
and U10084 (N_10084,N_7766,N_7720);
and U10085 (N_10085,N_8809,N_7848);
and U10086 (N_10086,N_8268,N_8915);
and U10087 (N_10087,N_7721,N_7943);
nor U10088 (N_10088,N_7670,N_8672);
nor U10089 (N_10089,N_8190,N_7694);
nand U10090 (N_10090,N_7847,N_7939);
or U10091 (N_10091,N_8294,N_7733);
nand U10092 (N_10092,N_8823,N_8003);
nand U10093 (N_10093,N_8564,N_7797);
xnor U10094 (N_10094,N_7580,N_8266);
xor U10095 (N_10095,N_8401,N_8636);
and U10096 (N_10096,N_8768,N_8018);
or U10097 (N_10097,N_7800,N_8700);
and U10098 (N_10098,N_8487,N_7620);
and U10099 (N_10099,N_7810,N_8427);
nand U10100 (N_10100,N_8448,N_8193);
or U10101 (N_10101,N_7562,N_8540);
nor U10102 (N_10102,N_7959,N_8255);
and U10103 (N_10103,N_8786,N_8934);
or U10104 (N_10104,N_7815,N_8710);
nand U10105 (N_10105,N_7674,N_8908);
nor U10106 (N_10106,N_8888,N_7955);
nand U10107 (N_10107,N_8784,N_8471);
nand U10108 (N_10108,N_8943,N_8559);
nand U10109 (N_10109,N_8578,N_8269);
nor U10110 (N_10110,N_8487,N_8083);
and U10111 (N_10111,N_7744,N_8690);
nand U10112 (N_10112,N_8155,N_8733);
and U10113 (N_10113,N_7552,N_7743);
nor U10114 (N_10114,N_8933,N_7856);
and U10115 (N_10115,N_8724,N_7703);
nor U10116 (N_10116,N_8736,N_8919);
nor U10117 (N_10117,N_8172,N_8335);
and U10118 (N_10118,N_8258,N_8036);
and U10119 (N_10119,N_8271,N_7677);
nor U10120 (N_10120,N_8026,N_8206);
and U10121 (N_10121,N_7927,N_7618);
nand U10122 (N_10122,N_8960,N_7510);
nor U10123 (N_10123,N_7760,N_8777);
or U10124 (N_10124,N_8163,N_8963);
nor U10125 (N_10125,N_8683,N_8369);
nand U10126 (N_10126,N_7966,N_8335);
nor U10127 (N_10127,N_8327,N_7969);
and U10128 (N_10128,N_8936,N_8591);
nand U10129 (N_10129,N_7902,N_8378);
or U10130 (N_10130,N_8997,N_8324);
and U10131 (N_10131,N_8280,N_8390);
nor U10132 (N_10132,N_7785,N_8121);
nand U10133 (N_10133,N_8767,N_7582);
nand U10134 (N_10134,N_8719,N_8712);
nand U10135 (N_10135,N_7861,N_7549);
nor U10136 (N_10136,N_7578,N_8045);
and U10137 (N_10137,N_8038,N_8547);
and U10138 (N_10138,N_8624,N_7880);
nand U10139 (N_10139,N_7513,N_8725);
and U10140 (N_10140,N_7837,N_8626);
and U10141 (N_10141,N_7653,N_7970);
or U10142 (N_10142,N_8770,N_7960);
xnor U10143 (N_10143,N_7746,N_7811);
or U10144 (N_10144,N_8020,N_8816);
or U10145 (N_10145,N_8951,N_8703);
or U10146 (N_10146,N_8607,N_7985);
or U10147 (N_10147,N_8234,N_7618);
nand U10148 (N_10148,N_8170,N_8465);
or U10149 (N_10149,N_7909,N_8155);
and U10150 (N_10150,N_8598,N_8736);
and U10151 (N_10151,N_8887,N_8746);
nor U10152 (N_10152,N_8803,N_8886);
or U10153 (N_10153,N_8928,N_8995);
nand U10154 (N_10154,N_7514,N_8902);
nand U10155 (N_10155,N_7645,N_8839);
nand U10156 (N_10156,N_7542,N_8717);
nor U10157 (N_10157,N_8577,N_7675);
nand U10158 (N_10158,N_7911,N_8903);
or U10159 (N_10159,N_7543,N_7907);
nand U10160 (N_10160,N_8384,N_8238);
nor U10161 (N_10161,N_7820,N_8141);
and U10162 (N_10162,N_8147,N_8193);
or U10163 (N_10163,N_8818,N_8689);
and U10164 (N_10164,N_7958,N_8158);
and U10165 (N_10165,N_7636,N_8160);
nor U10166 (N_10166,N_7569,N_8152);
nor U10167 (N_10167,N_7562,N_8578);
or U10168 (N_10168,N_7643,N_8862);
nand U10169 (N_10169,N_7688,N_7949);
and U10170 (N_10170,N_8089,N_8529);
nand U10171 (N_10171,N_7534,N_8853);
nand U10172 (N_10172,N_8591,N_8595);
or U10173 (N_10173,N_8812,N_8066);
nand U10174 (N_10174,N_8970,N_7808);
nand U10175 (N_10175,N_8693,N_7790);
or U10176 (N_10176,N_8113,N_7862);
and U10177 (N_10177,N_8285,N_8415);
and U10178 (N_10178,N_8562,N_8947);
or U10179 (N_10179,N_7703,N_7810);
or U10180 (N_10180,N_7625,N_7522);
and U10181 (N_10181,N_8896,N_7926);
and U10182 (N_10182,N_8712,N_8738);
and U10183 (N_10183,N_8513,N_8886);
nand U10184 (N_10184,N_8620,N_8934);
nand U10185 (N_10185,N_8788,N_7702);
nand U10186 (N_10186,N_8951,N_8763);
nand U10187 (N_10187,N_8895,N_7641);
or U10188 (N_10188,N_8780,N_8561);
xor U10189 (N_10189,N_8264,N_8576);
and U10190 (N_10190,N_8540,N_7767);
nor U10191 (N_10191,N_7527,N_8824);
nand U10192 (N_10192,N_8362,N_8767);
and U10193 (N_10193,N_8000,N_7536);
nand U10194 (N_10194,N_8450,N_7552);
nand U10195 (N_10195,N_8944,N_8583);
nand U10196 (N_10196,N_7873,N_8091);
xor U10197 (N_10197,N_8412,N_8611);
or U10198 (N_10198,N_7590,N_7856);
or U10199 (N_10199,N_8791,N_8526);
nor U10200 (N_10200,N_8321,N_8595);
and U10201 (N_10201,N_7913,N_7624);
and U10202 (N_10202,N_8823,N_7910);
nor U10203 (N_10203,N_8622,N_8092);
and U10204 (N_10204,N_7976,N_8182);
and U10205 (N_10205,N_7842,N_7862);
nor U10206 (N_10206,N_7862,N_8309);
nor U10207 (N_10207,N_8782,N_8717);
or U10208 (N_10208,N_8942,N_7698);
nor U10209 (N_10209,N_8030,N_8656);
nor U10210 (N_10210,N_7836,N_8081);
and U10211 (N_10211,N_7879,N_8068);
nor U10212 (N_10212,N_7966,N_8248);
nor U10213 (N_10213,N_7518,N_8216);
or U10214 (N_10214,N_8160,N_8373);
nor U10215 (N_10215,N_7681,N_8973);
nand U10216 (N_10216,N_7896,N_7793);
nor U10217 (N_10217,N_8602,N_8913);
and U10218 (N_10218,N_7637,N_8993);
nor U10219 (N_10219,N_8308,N_7647);
or U10220 (N_10220,N_8620,N_7658);
and U10221 (N_10221,N_8004,N_7625);
or U10222 (N_10222,N_8004,N_8945);
nand U10223 (N_10223,N_7642,N_7771);
nand U10224 (N_10224,N_7776,N_8088);
and U10225 (N_10225,N_8524,N_8014);
nor U10226 (N_10226,N_8168,N_8669);
or U10227 (N_10227,N_8346,N_7819);
and U10228 (N_10228,N_7654,N_8834);
and U10229 (N_10229,N_8081,N_8311);
nor U10230 (N_10230,N_8312,N_8447);
and U10231 (N_10231,N_7555,N_7890);
nand U10232 (N_10232,N_8046,N_8476);
and U10233 (N_10233,N_7989,N_8982);
nand U10234 (N_10234,N_8717,N_8759);
or U10235 (N_10235,N_8171,N_7580);
or U10236 (N_10236,N_8678,N_7813);
nor U10237 (N_10237,N_8870,N_8995);
nand U10238 (N_10238,N_7682,N_8152);
and U10239 (N_10239,N_8608,N_8700);
nor U10240 (N_10240,N_7500,N_8286);
nor U10241 (N_10241,N_7831,N_7713);
nand U10242 (N_10242,N_8790,N_8994);
nand U10243 (N_10243,N_8123,N_8718);
nand U10244 (N_10244,N_8010,N_8735);
and U10245 (N_10245,N_7709,N_8950);
nor U10246 (N_10246,N_8662,N_8382);
nand U10247 (N_10247,N_7917,N_8516);
nand U10248 (N_10248,N_8679,N_8649);
and U10249 (N_10249,N_7953,N_7870);
nand U10250 (N_10250,N_8607,N_8151);
nand U10251 (N_10251,N_8424,N_7735);
nor U10252 (N_10252,N_8294,N_8070);
or U10253 (N_10253,N_7905,N_7590);
nor U10254 (N_10254,N_8175,N_8777);
nand U10255 (N_10255,N_8439,N_8778);
and U10256 (N_10256,N_8056,N_7893);
nand U10257 (N_10257,N_7660,N_7558);
nand U10258 (N_10258,N_8627,N_8390);
nor U10259 (N_10259,N_8010,N_7664);
or U10260 (N_10260,N_7906,N_8761);
or U10261 (N_10261,N_8446,N_7672);
nand U10262 (N_10262,N_7897,N_7761);
or U10263 (N_10263,N_8421,N_7745);
nand U10264 (N_10264,N_7743,N_8773);
or U10265 (N_10265,N_8149,N_7773);
and U10266 (N_10266,N_8590,N_8553);
nor U10267 (N_10267,N_7991,N_8784);
or U10268 (N_10268,N_8664,N_8403);
nor U10269 (N_10269,N_8536,N_7683);
nand U10270 (N_10270,N_7527,N_8819);
and U10271 (N_10271,N_7891,N_8581);
nand U10272 (N_10272,N_7581,N_7729);
nor U10273 (N_10273,N_8624,N_7545);
nand U10274 (N_10274,N_8065,N_7846);
or U10275 (N_10275,N_8711,N_8594);
or U10276 (N_10276,N_8658,N_8583);
and U10277 (N_10277,N_8245,N_8499);
or U10278 (N_10278,N_7690,N_7759);
and U10279 (N_10279,N_7981,N_7554);
nor U10280 (N_10280,N_8114,N_7644);
xor U10281 (N_10281,N_7843,N_8250);
nand U10282 (N_10282,N_8063,N_8652);
or U10283 (N_10283,N_7799,N_8629);
and U10284 (N_10284,N_8859,N_8564);
nand U10285 (N_10285,N_7880,N_8879);
nor U10286 (N_10286,N_7809,N_8929);
nand U10287 (N_10287,N_8667,N_7753);
nor U10288 (N_10288,N_8864,N_8894);
and U10289 (N_10289,N_8851,N_8720);
and U10290 (N_10290,N_7524,N_7853);
nor U10291 (N_10291,N_7827,N_7660);
nand U10292 (N_10292,N_8753,N_7932);
nand U10293 (N_10293,N_7789,N_7665);
and U10294 (N_10294,N_8256,N_7786);
nand U10295 (N_10295,N_8530,N_7993);
and U10296 (N_10296,N_8343,N_8878);
or U10297 (N_10297,N_8512,N_7690);
or U10298 (N_10298,N_7662,N_7940);
nand U10299 (N_10299,N_8159,N_7929);
and U10300 (N_10300,N_8832,N_8454);
nand U10301 (N_10301,N_7714,N_7949);
nand U10302 (N_10302,N_8476,N_7764);
nand U10303 (N_10303,N_8700,N_8723);
nand U10304 (N_10304,N_7917,N_8375);
nor U10305 (N_10305,N_7633,N_8895);
nand U10306 (N_10306,N_8004,N_8743);
and U10307 (N_10307,N_8141,N_8048);
or U10308 (N_10308,N_7998,N_7960);
nand U10309 (N_10309,N_8152,N_7595);
or U10310 (N_10310,N_7715,N_7997);
and U10311 (N_10311,N_8193,N_7518);
nor U10312 (N_10312,N_8478,N_8929);
and U10313 (N_10313,N_7951,N_8314);
and U10314 (N_10314,N_7583,N_8399);
and U10315 (N_10315,N_8188,N_7535);
and U10316 (N_10316,N_8098,N_7797);
nand U10317 (N_10317,N_8226,N_7592);
or U10318 (N_10318,N_7522,N_8729);
nand U10319 (N_10319,N_8730,N_8986);
nor U10320 (N_10320,N_8555,N_8755);
and U10321 (N_10321,N_8634,N_7626);
nand U10322 (N_10322,N_8149,N_8007);
or U10323 (N_10323,N_8087,N_7969);
and U10324 (N_10324,N_8754,N_8576);
nor U10325 (N_10325,N_8949,N_7559);
and U10326 (N_10326,N_8446,N_8711);
nor U10327 (N_10327,N_8490,N_7684);
nor U10328 (N_10328,N_7970,N_7704);
nand U10329 (N_10329,N_8186,N_7754);
nand U10330 (N_10330,N_7939,N_8373);
and U10331 (N_10331,N_8007,N_7871);
and U10332 (N_10332,N_8896,N_8225);
or U10333 (N_10333,N_8289,N_7962);
or U10334 (N_10334,N_8720,N_8288);
xnor U10335 (N_10335,N_8079,N_8726);
or U10336 (N_10336,N_7922,N_7733);
or U10337 (N_10337,N_7994,N_8828);
nor U10338 (N_10338,N_7572,N_8582);
nand U10339 (N_10339,N_8504,N_8743);
nand U10340 (N_10340,N_8503,N_8284);
or U10341 (N_10341,N_7958,N_8622);
or U10342 (N_10342,N_8005,N_8923);
nand U10343 (N_10343,N_8486,N_7784);
or U10344 (N_10344,N_8513,N_7611);
xnor U10345 (N_10345,N_8269,N_8627);
or U10346 (N_10346,N_7829,N_8838);
or U10347 (N_10347,N_8422,N_7500);
and U10348 (N_10348,N_7731,N_8970);
or U10349 (N_10349,N_7662,N_8790);
or U10350 (N_10350,N_8115,N_8716);
or U10351 (N_10351,N_8855,N_8534);
and U10352 (N_10352,N_8241,N_8295);
or U10353 (N_10353,N_8770,N_8256);
nand U10354 (N_10354,N_7500,N_8505);
or U10355 (N_10355,N_7760,N_8911);
or U10356 (N_10356,N_7953,N_7556);
and U10357 (N_10357,N_8114,N_8868);
or U10358 (N_10358,N_7848,N_8748);
or U10359 (N_10359,N_7972,N_8600);
or U10360 (N_10360,N_7774,N_8827);
nand U10361 (N_10361,N_7608,N_8606);
nor U10362 (N_10362,N_7802,N_8616);
nor U10363 (N_10363,N_8186,N_8020);
and U10364 (N_10364,N_7523,N_8511);
and U10365 (N_10365,N_8043,N_7792);
or U10366 (N_10366,N_8033,N_8432);
nor U10367 (N_10367,N_7879,N_8828);
nor U10368 (N_10368,N_7813,N_7509);
nor U10369 (N_10369,N_8012,N_8189);
and U10370 (N_10370,N_8699,N_8918);
and U10371 (N_10371,N_8512,N_8811);
or U10372 (N_10372,N_7720,N_7788);
and U10373 (N_10373,N_8702,N_8285);
or U10374 (N_10374,N_8931,N_8034);
nand U10375 (N_10375,N_8214,N_7506);
nor U10376 (N_10376,N_7584,N_8245);
nor U10377 (N_10377,N_8261,N_8513);
nand U10378 (N_10378,N_8717,N_8362);
and U10379 (N_10379,N_8733,N_7943);
and U10380 (N_10380,N_8159,N_8987);
nor U10381 (N_10381,N_8140,N_8247);
nor U10382 (N_10382,N_8826,N_8739);
nor U10383 (N_10383,N_7579,N_8805);
and U10384 (N_10384,N_7593,N_8106);
and U10385 (N_10385,N_8620,N_7721);
nor U10386 (N_10386,N_8791,N_7546);
nand U10387 (N_10387,N_7880,N_8445);
and U10388 (N_10388,N_8827,N_7654);
nand U10389 (N_10389,N_7580,N_7834);
or U10390 (N_10390,N_8360,N_7894);
or U10391 (N_10391,N_8527,N_8274);
and U10392 (N_10392,N_8021,N_8887);
nand U10393 (N_10393,N_8730,N_8074);
or U10394 (N_10394,N_8843,N_8787);
nand U10395 (N_10395,N_8226,N_8963);
nand U10396 (N_10396,N_8293,N_7600);
and U10397 (N_10397,N_8677,N_7912);
or U10398 (N_10398,N_8303,N_8809);
or U10399 (N_10399,N_8465,N_8380);
xnor U10400 (N_10400,N_8549,N_8764);
nor U10401 (N_10401,N_7774,N_8555);
nand U10402 (N_10402,N_8327,N_8512);
or U10403 (N_10403,N_8368,N_8165);
and U10404 (N_10404,N_8877,N_8406);
or U10405 (N_10405,N_8869,N_8610);
or U10406 (N_10406,N_7692,N_8815);
or U10407 (N_10407,N_7963,N_8404);
or U10408 (N_10408,N_8527,N_7956);
and U10409 (N_10409,N_7992,N_8365);
and U10410 (N_10410,N_8755,N_7823);
nand U10411 (N_10411,N_8249,N_8837);
or U10412 (N_10412,N_8878,N_8368);
or U10413 (N_10413,N_8300,N_8637);
nor U10414 (N_10414,N_8716,N_8904);
and U10415 (N_10415,N_8285,N_7541);
or U10416 (N_10416,N_8030,N_8825);
or U10417 (N_10417,N_7903,N_7865);
or U10418 (N_10418,N_8142,N_8113);
or U10419 (N_10419,N_8135,N_8067);
xor U10420 (N_10420,N_8653,N_7980);
nor U10421 (N_10421,N_8202,N_8605);
and U10422 (N_10422,N_8674,N_7569);
or U10423 (N_10423,N_8782,N_7781);
and U10424 (N_10424,N_7547,N_8216);
or U10425 (N_10425,N_7561,N_7946);
nor U10426 (N_10426,N_8913,N_7950);
and U10427 (N_10427,N_8408,N_8867);
xnor U10428 (N_10428,N_8368,N_8356);
or U10429 (N_10429,N_7670,N_8575);
and U10430 (N_10430,N_8533,N_7885);
nor U10431 (N_10431,N_7917,N_8619);
nand U10432 (N_10432,N_7771,N_8130);
and U10433 (N_10433,N_8650,N_8887);
nor U10434 (N_10434,N_8201,N_7663);
nand U10435 (N_10435,N_8254,N_7521);
or U10436 (N_10436,N_8174,N_8097);
nand U10437 (N_10437,N_8065,N_7799);
and U10438 (N_10438,N_8766,N_8452);
nor U10439 (N_10439,N_8543,N_8534);
nor U10440 (N_10440,N_8729,N_8680);
nand U10441 (N_10441,N_8369,N_8265);
or U10442 (N_10442,N_7661,N_8812);
and U10443 (N_10443,N_8145,N_7672);
or U10444 (N_10444,N_8797,N_8678);
nand U10445 (N_10445,N_8934,N_8204);
nor U10446 (N_10446,N_8791,N_7650);
and U10447 (N_10447,N_8357,N_7707);
and U10448 (N_10448,N_8666,N_8926);
or U10449 (N_10449,N_7747,N_7866);
and U10450 (N_10450,N_8069,N_7854);
nor U10451 (N_10451,N_8753,N_7575);
nor U10452 (N_10452,N_8410,N_8712);
nand U10453 (N_10453,N_8380,N_8370);
and U10454 (N_10454,N_8734,N_8379);
nor U10455 (N_10455,N_8817,N_7719);
nand U10456 (N_10456,N_8599,N_7742);
or U10457 (N_10457,N_8628,N_8421);
and U10458 (N_10458,N_8704,N_8125);
nand U10459 (N_10459,N_7835,N_7851);
or U10460 (N_10460,N_7812,N_8976);
nand U10461 (N_10461,N_8705,N_8346);
nand U10462 (N_10462,N_7789,N_8018);
and U10463 (N_10463,N_8401,N_8721);
nor U10464 (N_10464,N_7807,N_8848);
or U10465 (N_10465,N_8927,N_8828);
and U10466 (N_10466,N_7572,N_8566);
and U10467 (N_10467,N_7916,N_7589);
nor U10468 (N_10468,N_8772,N_8537);
nand U10469 (N_10469,N_8074,N_8151);
and U10470 (N_10470,N_8037,N_8710);
nor U10471 (N_10471,N_8358,N_8667);
and U10472 (N_10472,N_7839,N_8222);
nor U10473 (N_10473,N_7831,N_7816);
and U10474 (N_10474,N_7680,N_8890);
nand U10475 (N_10475,N_8638,N_8805);
nand U10476 (N_10476,N_8887,N_8799);
nand U10477 (N_10477,N_8836,N_8529);
nor U10478 (N_10478,N_8841,N_7883);
nand U10479 (N_10479,N_7960,N_7710);
or U10480 (N_10480,N_7710,N_8004);
xor U10481 (N_10481,N_8225,N_8422);
nor U10482 (N_10482,N_8107,N_7730);
and U10483 (N_10483,N_8061,N_8991);
and U10484 (N_10484,N_8902,N_8064);
nand U10485 (N_10485,N_8413,N_8820);
nor U10486 (N_10486,N_8673,N_8053);
and U10487 (N_10487,N_7920,N_7811);
nand U10488 (N_10488,N_8146,N_8444);
and U10489 (N_10489,N_8343,N_8142);
or U10490 (N_10490,N_8693,N_8263);
and U10491 (N_10491,N_7878,N_8014);
and U10492 (N_10492,N_8134,N_8168);
and U10493 (N_10493,N_8565,N_8522);
and U10494 (N_10494,N_7638,N_7645);
nand U10495 (N_10495,N_7818,N_8075);
and U10496 (N_10496,N_8265,N_8000);
and U10497 (N_10497,N_8693,N_7850);
nand U10498 (N_10498,N_8911,N_8640);
and U10499 (N_10499,N_8100,N_8571);
nor U10500 (N_10500,N_10373,N_10153);
nand U10501 (N_10501,N_9553,N_9756);
and U10502 (N_10502,N_10333,N_10494);
nor U10503 (N_10503,N_9549,N_9514);
or U10504 (N_10504,N_10357,N_9721);
and U10505 (N_10505,N_9273,N_9119);
nor U10506 (N_10506,N_9166,N_10330);
and U10507 (N_10507,N_9203,N_9500);
nand U10508 (N_10508,N_9853,N_10366);
and U10509 (N_10509,N_10384,N_9626);
nand U10510 (N_10510,N_10430,N_9713);
or U10511 (N_10511,N_10302,N_10012);
or U10512 (N_10512,N_9093,N_9659);
or U10513 (N_10513,N_10463,N_9785);
nand U10514 (N_10514,N_9021,N_10120);
and U10515 (N_10515,N_10404,N_9412);
and U10516 (N_10516,N_9333,N_9222);
and U10517 (N_10517,N_9368,N_9290);
nor U10518 (N_10518,N_9343,N_10247);
or U10519 (N_10519,N_10484,N_9774);
nand U10520 (N_10520,N_9895,N_9362);
or U10521 (N_10521,N_9184,N_9194);
nor U10522 (N_10522,N_9288,N_10278);
nand U10523 (N_10523,N_9998,N_9949);
nand U10524 (N_10524,N_9398,N_9267);
nor U10525 (N_10525,N_9661,N_10399);
and U10526 (N_10526,N_9728,N_9304);
nor U10527 (N_10527,N_9487,N_9211);
and U10528 (N_10528,N_9838,N_10392);
and U10529 (N_10529,N_9775,N_9481);
or U10530 (N_10530,N_10074,N_9313);
or U10531 (N_10531,N_10268,N_9479);
nor U10532 (N_10532,N_9277,N_10382);
xnor U10533 (N_10533,N_10217,N_10455);
nand U10534 (N_10534,N_9688,N_9674);
nand U10535 (N_10535,N_9972,N_10047);
nand U10536 (N_10536,N_9705,N_9421);
nand U10537 (N_10537,N_9557,N_9634);
and U10538 (N_10538,N_9723,N_9866);
or U10539 (N_10539,N_10176,N_9589);
nor U10540 (N_10540,N_10263,N_10202);
and U10541 (N_10541,N_9832,N_9735);
and U10542 (N_10542,N_9381,N_10155);
nor U10543 (N_10543,N_9305,N_10305);
or U10544 (N_10544,N_9952,N_9606);
and U10545 (N_10545,N_9174,N_10369);
nor U10546 (N_10546,N_10375,N_9591);
or U10547 (N_10547,N_10020,N_9978);
nand U10548 (N_10548,N_10477,N_10461);
xor U10549 (N_10549,N_9593,N_10239);
nor U10550 (N_10550,N_9090,N_9474);
nor U10551 (N_10551,N_9319,N_9173);
and U10552 (N_10552,N_10031,N_9827);
nor U10553 (N_10553,N_9217,N_9029);
and U10554 (N_10554,N_9725,N_9472);
nand U10555 (N_10555,N_9066,N_10150);
and U10556 (N_10556,N_9180,N_9291);
nor U10557 (N_10557,N_10209,N_9325);
or U10558 (N_10558,N_10381,N_10062);
nand U10559 (N_10559,N_9062,N_10487);
and U10560 (N_10560,N_9594,N_10024);
nand U10561 (N_10561,N_9954,N_9595);
or U10562 (N_10562,N_9434,N_9402);
or U10563 (N_10563,N_10439,N_10293);
and U10564 (N_10564,N_9657,N_9097);
nor U10565 (N_10565,N_9997,N_9161);
nor U10566 (N_10566,N_10486,N_9216);
and U10567 (N_10567,N_9048,N_9136);
or U10568 (N_10568,N_10246,N_9964);
or U10569 (N_10569,N_9238,N_9205);
nor U10570 (N_10570,N_9878,N_9641);
and U10571 (N_10571,N_9639,N_9698);
nand U10572 (N_10572,N_9407,N_10379);
nor U10573 (N_10573,N_10126,N_10470);
nand U10574 (N_10574,N_9590,N_9200);
or U10575 (N_10575,N_10460,N_9015);
nand U10576 (N_10576,N_9005,N_9079);
nor U10577 (N_10577,N_9341,N_9058);
and U10578 (N_10578,N_9669,N_9944);
nand U10579 (N_10579,N_9631,N_9787);
xor U10580 (N_10580,N_9007,N_9121);
nand U10581 (N_10581,N_9262,N_9495);
or U10582 (N_10582,N_9582,N_9030);
or U10583 (N_10583,N_9840,N_10130);
nand U10584 (N_10584,N_9215,N_9570);
nand U10585 (N_10585,N_9547,N_9017);
nand U10586 (N_10586,N_10482,N_10168);
or U10587 (N_10587,N_9771,N_10206);
or U10588 (N_10588,N_9129,N_10255);
and U10589 (N_10589,N_9815,N_9336);
nand U10590 (N_10590,N_9958,N_9406);
or U10591 (N_10591,N_10037,N_9792);
and U10592 (N_10592,N_10148,N_10426);
and U10593 (N_10593,N_9845,N_9767);
nand U10594 (N_10594,N_9176,N_9138);
and U10595 (N_10595,N_9812,N_10203);
and U10596 (N_10596,N_9706,N_9115);
nor U10597 (N_10597,N_9692,N_9051);
nand U10598 (N_10598,N_9271,N_9965);
nand U10599 (N_10599,N_9356,N_9134);
nand U10600 (N_10600,N_9403,N_9801);
and U10601 (N_10601,N_9835,N_9747);
nor U10602 (N_10602,N_9419,N_10158);
nand U10603 (N_10603,N_9940,N_9170);
nor U10604 (N_10604,N_9888,N_9491);
nor U10605 (N_10605,N_9401,N_9887);
or U10606 (N_10606,N_9159,N_9625);
nor U10607 (N_10607,N_9507,N_10266);
nor U10608 (N_10608,N_10115,N_9332);
nand U10609 (N_10609,N_9742,N_9919);
nor U10610 (N_10610,N_9187,N_9882);
nor U10611 (N_10611,N_9810,N_9683);
and U10612 (N_10612,N_10058,N_9156);
nor U10613 (N_10613,N_9921,N_9453);
nand U10614 (N_10614,N_9636,N_10456);
nand U10615 (N_10615,N_10067,N_10124);
and U10616 (N_10616,N_10006,N_9955);
nand U10617 (N_10617,N_9724,N_9351);
or U10618 (N_10618,N_9635,N_9060);
nand U10619 (N_10619,N_9183,N_9632);
nand U10620 (N_10620,N_10267,N_10110);
nor U10621 (N_10621,N_10118,N_10013);
nor U10622 (N_10622,N_10036,N_9618);
nor U10623 (N_10623,N_9772,N_9982);
nand U10624 (N_10624,N_10454,N_9254);
nor U10625 (N_10625,N_10408,N_9164);
and U10626 (N_10626,N_10133,N_9408);
and U10627 (N_10627,N_10044,N_9163);
or U10628 (N_10628,N_9498,N_9150);
nand U10629 (N_10629,N_10046,N_9755);
nor U10630 (N_10630,N_9148,N_10476);
nor U10631 (N_10631,N_10041,N_10167);
nor U10632 (N_10632,N_10114,N_10145);
nor U10633 (N_10633,N_9019,N_9936);
nor U10634 (N_10634,N_9300,N_9390);
and U10635 (N_10635,N_10332,N_10179);
or U10636 (N_10636,N_10241,N_10151);
or U10637 (N_10637,N_10339,N_9743);
or U10638 (N_10638,N_9764,N_10415);
or U10639 (N_10639,N_10019,N_9846);
nand U10640 (N_10640,N_9397,N_10273);
nor U10641 (N_10641,N_9354,N_10423);
xor U10642 (N_10642,N_10068,N_9535);
and U10643 (N_10643,N_9848,N_9744);
and U10644 (N_10644,N_10452,N_9380);
nor U10645 (N_10645,N_10225,N_9769);
or U10646 (N_10646,N_10199,N_9002);
or U10647 (N_10647,N_9046,N_9369);
nand U10648 (N_10648,N_10218,N_10223);
nand U10649 (N_10649,N_10295,N_9863);
and U10650 (N_10650,N_9602,N_10342);
or U10651 (N_10651,N_10257,N_9433);
nand U10652 (N_10652,N_10464,N_9816);
or U10653 (N_10653,N_10211,N_10403);
nor U10654 (N_10654,N_9349,N_10250);
or U10655 (N_10655,N_9577,N_10097);
or U10656 (N_10656,N_9992,N_9001);
nand U10657 (N_10657,N_9494,N_9116);
and U10658 (N_10658,N_10001,N_9579);
nor U10659 (N_10659,N_10412,N_10190);
nand U10660 (N_10660,N_9033,N_9469);
nor U10661 (N_10661,N_10023,N_10318);
nor U10662 (N_10662,N_10205,N_9670);
and U10663 (N_10663,N_9074,N_10316);
or U10664 (N_10664,N_10016,N_9685);
and U10665 (N_10665,N_9207,N_10371);
nor U10666 (N_10666,N_10060,N_9794);
nand U10667 (N_10667,N_10076,N_9569);
and U10668 (N_10668,N_9568,N_9455);
and U10669 (N_10669,N_9506,N_10304);
nor U10670 (N_10670,N_9908,N_9563);
nor U10671 (N_10671,N_9730,N_9773);
nand U10672 (N_10672,N_9283,N_9808);
or U10673 (N_10673,N_9152,N_9966);
nand U10674 (N_10674,N_10405,N_9519);
nand U10675 (N_10675,N_9399,N_9361);
nor U10676 (N_10676,N_9654,N_9752);
nor U10677 (N_10677,N_10171,N_9485);
or U10678 (N_10678,N_9647,N_9762);
nor U10679 (N_10679,N_10351,N_9665);
and U10680 (N_10680,N_10374,N_9938);
and U10681 (N_10681,N_10083,N_9127);
nor U10682 (N_10682,N_10088,N_9172);
nor U10683 (N_10683,N_9653,N_10280);
nor U10684 (N_10684,N_9040,N_10327);
and U10685 (N_10685,N_10215,N_9315);
or U10686 (N_10686,N_10372,N_9522);
and U10687 (N_10687,N_9109,N_10216);
nor U10688 (N_10688,N_10324,N_10285);
and U10689 (N_10689,N_9236,N_10222);
and U10690 (N_10690,N_9426,N_9901);
or U10691 (N_10691,N_10146,N_9517);
or U10692 (N_10692,N_10416,N_9796);
and U10693 (N_10693,N_9145,N_9210);
nand U10694 (N_10694,N_9682,N_9822);
and U10695 (N_10695,N_9658,N_9346);
and U10696 (N_10696,N_9886,N_9316);
nand U10697 (N_10697,N_10326,N_9087);
nand U10698 (N_10698,N_9352,N_9786);
or U10699 (N_10699,N_9444,N_9873);
nor U10700 (N_10700,N_9228,N_9189);
nand U10701 (N_10701,N_10035,N_10185);
nand U10702 (N_10702,N_9269,N_9169);
nor U10703 (N_10703,N_9289,N_9338);
or U10704 (N_10704,N_9611,N_9460);
nor U10705 (N_10705,N_9197,N_9142);
nand U10706 (N_10706,N_9693,N_9024);
and U10707 (N_10707,N_9247,N_10424);
nand U10708 (N_10708,N_9781,N_9096);
and U10709 (N_10709,N_9761,N_10389);
or U10710 (N_10710,N_9256,N_10029);
nand U10711 (N_10711,N_9061,N_9562);
nand U10712 (N_10712,N_10099,N_9573);
nor U10713 (N_10713,N_10492,N_10224);
nor U10714 (N_10714,N_9696,N_10243);
or U10715 (N_10715,N_9328,N_9057);
and U10716 (N_10716,N_9345,N_10499);
and U10717 (N_10717,N_9043,N_9085);
and U10718 (N_10718,N_10233,N_9310);
or U10719 (N_10719,N_9100,N_10207);
nand U10720 (N_10720,N_9923,N_9400);
or U10721 (N_10721,N_10394,N_10201);
nor U10722 (N_10722,N_10481,N_9969);
and U10723 (N_10723,N_10162,N_10063);
nand U10724 (N_10724,N_10363,N_9028);
and U10725 (N_10725,N_9107,N_9449);
nand U10726 (N_10726,N_9600,N_10090);
and U10727 (N_10727,N_9175,N_9082);
nand U10728 (N_10728,N_9975,N_10433);
or U10729 (N_10729,N_10112,N_9359);
nand U10730 (N_10730,N_9979,N_9671);
and U10731 (N_10731,N_9204,N_10457);
or U10732 (N_10732,N_10322,N_10238);
nand U10733 (N_10733,N_10100,N_9745);
or U10734 (N_10734,N_9610,N_10143);
nand U10735 (N_10735,N_10301,N_10117);
and U10736 (N_10736,N_10284,N_9282);
and U10737 (N_10737,N_10227,N_10077);
or U10738 (N_10738,N_9515,N_10249);
nand U10739 (N_10739,N_9086,N_10475);
nor U10740 (N_10740,N_10320,N_9431);
nor U10741 (N_10741,N_9864,N_9993);
and U10742 (N_10742,N_10248,N_10080);
nor U10743 (N_10743,N_9218,N_9417);
xnor U10744 (N_10744,N_9961,N_9738);
nor U10745 (N_10745,N_9650,N_10210);
nand U10746 (N_10746,N_10410,N_10358);
nand U10747 (N_10747,N_9574,N_9829);
nand U10748 (N_10748,N_9384,N_9736);
xnor U10749 (N_10749,N_9766,N_9084);
nand U10750 (N_10750,N_10376,N_9896);
or U10751 (N_10751,N_9914,N_10256);
nor U10752 (N_10752,N_10039,N_10377);
or U10753 (N_10753,N_9006,N_10490);
and U10754 (N_10754,N_9892,N_10395);
nand U10755 (N_10755,N_9836,N_10135);
and U10756 (N_10756,N_10109,N_9411);
and U10757 (N_10757,N_9396,N_9340);
and U10758 (N_10758,N_9104,N_10303);
nor U10759 (N_10759,N_9904,N_10313);
nor U10760 (N_10760,N_9244,N_10480);
or U10761 (N_10761,N_9101,N_10378);
nand U10762 (N_10762,N_10421,N_9734);
or U10763 (N_10763,N_9027,N_10467);
xor U10764 (N_10764,N_10193,N_9881);
and U10765 (N_10765,N_9684,N_9153);
or U10766 (N_10766,N_9967,N_9828);
nand U10767 (N_10767,N_9788,N_10136);
and U10768 (N_10768,N_9056,N_9372);
or U10769 (N_10769,N_9457,N_9415);
xor U10770 (N_10770,N_9675,N_9227);
and U10771 (N_10771,N_10204,N_9648);
or U10772 (N_10772,N_9946,N_9284);
nor U10773 (N_10773,N_9758,N_9414);
nor U10774 (N_10774,N_10191,N_9118);
nor U10775 (N_10775,N_9311,N_9939);
xnor U10776 (N_10776,N_10163,N_10253);
and U10777 (N_10777,N_9081,N_9375);
or U10778 (N_10778,N_9662,N_9167);
nand U10779 (N_10779,N_9286,N_9365);
nor U10780 (N_10780,N_10220,N_10123);
nand U10781 (N_10781,N_9666,N_9274);
or U10782 (N_10782,N_9893,N_10321);
and U10783 (N_10783,N_10214,N_10050);
nor U10784 (N_10784,N_10106,N_9425);
nor U10785 (N_10785,N_10187,N_9245);
nand U10786 (N_10786,N_9710,N_10312);
and U10787 (N_10787,N_9470,N_9446);
nor U10788 (N_10788,N_9091,N_9686);
or U10789 (N_10789,N_9473,N_10348);
xor U10790 (N_10790,N_10094,N_9373);
nor U10791 (N_10791,N_9850,N_9441);
or U10792 (N_10792,N_9942,N_10309);
or U10793 (N_10793,N_10105,N_9137);
xor U10794 (N_10794,N_9545,N_9996);
nor U10795 (N_10795,N_9039,N_9320);
and U10796 (N_10796,N_10497,N_9071);
and U10797 (N_10797,N_9054,N_9748);
and U10798 (N_10798,N_10010,N_9480);
or U10799 (N_10799,N_9382,N_9655);
nor U10800 (N_10800,N_10496,N_9041);
xor U10801 (N_10801,N_9592,N_9999);
nand U10802 (N_10802,N_9697,N_9022);
and U10803 (N_10803,N_10393,N_10345);
and U10804 (N_10804,N_9916,N_9977);
nor U10805 (N_10805,N_10367,N_10265);
nor U10806 (N_10806,N_9225,N_9943);
nor U10807 (N_10807,N_9149,N_9806);
xnor U10808 (N_10808,N_9571,N_10025);
or U10809 (N_10809,N_9621,N_10438);
or U10810 (N_10810,N_9428,N_9819);
or U10811 (N_10811,N_9727,N_9239);
or U10812 (N_10812,N_9567,N_9869);
nand U10813 (N_10813,N_9760,N_9374);
nor U10814 (N_10814,N_10196,N_10361);
and U10815 (N_10815,N_10445,N_10072);
or U10816 (N_10816,N_9422,N_9917);
and U10817 (N_10817,N_9912,N_10449);
nor U10818 (N_10818,N_10414,N_9672);
nor U10819 (N_10819,N_9597,N_9925);
nand U10820 (N_10820,N_9141,N_9974);
nand U10821 (N_10821,N_9139,N_9443);
nand U10822 (N_10822,N_9642,N_9813);
or U10823 (N_10823,N_10428,N_9584);
and U10824 (N_10824,N_9548,N_9157);
xor U10825 (N_10825,N_10251,N_9257);
nand U10826 (N_10826,N_9249,N_9834);
or U10827 (N_10827,N_9779,N_10420);
or U10828 (N_10828,N_10198,N_9889);
or U10829 (N_10829,N_9330,N_10432);
and U10830 (N_10830,N_10113,N_9064);
and U10831 (N_10831,N_10033,N_9209);
nand U10832 (N_10832,N_10479,N_10197);
and U10833 (N_10833,N_9782,N_9055);
or U10834 (N_10834,N_9950,N_10021);
nand U10835 (N_10835,N_9861,N_10078);
and U10836 (N_10836,N_9126,N_9504);
nand U10837 (N_10837,N_9114,N_10360);
and U10838 (N_10838,N_10434,N_9722);
nor U10839 (N_10839,N_9561,N_9404);
or U10840 (N_10840,N_9322,N_9050);
xnor U10841 (N_10841,N_9078,N_9456);
nand U10842 (N_10842,N_9379,N_10468);
and U10843 (N_10843,N_9435,N_10485);
or U10844 (N_10844,N_10003,N_9614);
or U10845 (N_10845,N_9783,N_9047);
and U10846 (N_10846,N_9070,N_10459);
and U10847 (N_10847,N_9113,N_9035);
nand U10848 (N_10848,N_9246,N_9529);
nor U10849 (N_10849,N_9376,N_10262);
xnor U10850 (N_10850,N_9663,N_9128);
nand U10851 (N_10851,N_10128,N_10419);
nand U10852 (N_10852,N_9823,N_9587);
and U10853 (N_10853,N_9044,N_10200);
nor U10854 (N_10854,N_10290,N_10057);
nand U10855 (N_10855,N_9991,N_10258);
nand U10856 (N_10856,N_10306,N_9185);
and U10857 (N_10857,N_9601,N_9413);
or U10858 (N_10858,N_9875,N_9214);
nand U10859 (N_10859,N_9691,N_9818);
and U10860 (N_10860,N_9931,N_9377);
and U10861 (N_10861,N_9757,N_10221);
or U10862 (N_10862,N_9751,N_10084);
and U10863 (N_10863,N_9447,N_10271);
or U10864 (N_10864,N_9147,N_9088);
or U10865 (N_10865,N_10356,N_9660);
or U10866 (N_10866,N_10127,N_10472);
xor U10867 (N_10867,N_10272,N_9477);
nand U10868 (N_10868,N_10129,N_9793);
or U10869 (N_10869,N_9440,N_9234);
nand U10870 (N_10870,N_9740,N_10493);
or U10871 (N_10871,N_9510,N_9484);
and U10872 (N_10872,N_10385,N_9181);
or U10873 (N_10873,N_9556,N_10331);
or U10874 (N_10874,N_9080,N_10352);
and U10875 (N_10875,N_9110,N_9820);
nor U10876 (N_10876,N_10279,N_9125);
nand U10877 (N_10877,N_10052,N_9894);
and U10878 (N_10878,N_10043,N_9392);
and U10879 (N_10879,N_9324,N_10401);
nor U10880 (N_10880,N_9623,N_9031);
nand U10881 (N_10881,N_9502,N_9532);
or U10882 (N_10882,N_9059,N_10134);
and U10883 (N_10883,N_10314,N_9701);
nand U10884 (N_10884,N_9279,N_9450);
and U10885 (N_10885,N_10140,N_9366);
or U10886 (N_10886,N_10427,N_9821);
and U10887 (N_10887,N_9937,N_10446);
nand U10888 (N_10888,N_10131,N_9191);
nor U10889 (N_10889,N_9656,N_10056);
nand U10890 (N_10890,N_9988,N_10294);
nand U10891 (N_10891,N_9907,N_9000);
or U10892 (N_10892,N_9242,N_10450);
or U10893 (N_10893,N_10045,N_9870);
nor U10894 (N_10894,N_9980,N_9266);
nand U10895 (N_10895,N_10048,N_9168);
nand U10896 (N_10896,N_9903,N_9538);
and U10897 (N_10897,N_10400,N_10089);
or U10898 (N_10898,N_10213,N_9393);
xor U10899 (N_10899,N_9018,N_10422);
or U10900 (N_10900,N_9857,N_9464);
nand U10901 (N_10901,N_9985,N_9638);
nor U10902 (N_10902,N_9603,N_9784);
nand U10903 (N_10903,N_9524,N_10390);
or U10904 (N_10904,N_9367,N_9520);
xor U10905 (N_10905,N_10355,N_10437);
and U10906 (N_10906,N_10364,N_9508);
nor U10907 (N_10907,N_9841,N_10226);
or U10908 (N_10908,N_9814,N_9883);
xor U10909 (N_10909,N_9552,N_9984);
and U10910 (N_10910,N_9489,N_10066);
nor U10911 (N_10911,N_9526,N_9466);
and U10912 (N_10912,N_9973,N_10299);
nor U10913 (N_10913,N_9689,N_10125);
or U10914 (N_10914,N_9220,N_9876);
or U10915 (N_10915,N_10275,N_9700);
nand U10916 (N_10916,N_9750,N_10409);
or U10917 (N_10917,N_10368,N_9759);
nor U10918 (N_10918,N_9409,N_9909);
or U10919 (N_10919,N_9702,N_10453);
nand U10920 (N_10920,N_9424,N_10236);
xnor U10921 (N_10921,N_9025,N_10121);
nor U10922 (N_10922,N_9436,N_9360);
or U10923 (N_10923,N_9679,N_9072);
nor U10924 (N_10924,N_9296,N_10189);
and U10925 (N_10925,N_10443,N_10245);
and U10926 (N_10926,N_9729,N_9461);
and U10927 (N_10927,N_9038,N_9709);
and U10928 (N_10928,N_10283,N_9008);
nor U10929 (N_10929,N_9492,N_10177);
nand U10930 (N_10930,N_9095,N_9957);
and U10931 (N_10931,N_9158,N_9852);
and U10932 (N_10932,N_9598,N_9445);
or U10933 (N_10933,N_9651,N_9294);
or U10934 (N_10934,N_9765,N_9012);
nor U10935 (N_10935,N_9695,N_10232);
nor U10936 (N_10936,N_9233,N_9490);
and U10937 (N_10937,N_9378,N_9664);
nor U10938 (N_10938,N_9468,N_10152);
and U10939 (N_10939,N_9927,N_10073);
and U10940 (N_10940,N_9014,N_9326);
nor U10941 (N_10941,N_10172,N_9179);
or U10942 (N_10942,N_10182,N_9036);
nor U10943 (N_10943,N_9230,N_9512);
or U10944 (N_10944,N_9963,N_10132);
nor U10945 (N_10945,N_9438,N_9699);
and U10946 (N_10946,N_9309,N_10173);
nor U10947 (N_10947,N_10488,N_9911);
and U10948 (N_10948,N_9260,N_9833);
nor U10949 (N_10949,N_9276,N_9877);
nor U10950 (N_10950,N_9165,N_10064);
nand U10951 (N_10951,N_9010,N_10288);
nand U10952 (N_10952,N_9342,N_10059);
nand U10953 (N_10953,N_9630,N_9112);
and U10954 (N_10954,N_9192,N_10362);
nor U10955 (N_10955,N_9613,N_9891);
nor U10956 (N_10956,N_9073,N_10259);
and U10957 (N_10957,N_9859,N_9023);
nand U10958 (N_10958,N_9250,N_9668);
or U10959 (N_10959,N_9627,N_9117);
and U10960 (N_10960,N_9753,N_10329);
or U10961 (N_10961,N_9212,N_9146);
and U10962 (N_10962,N_9499,N_10065);
nand U10963 (N_10963,N_9799,N_9716);
or U10964 (N_10964,N_10169,N_10370);
nand U10965 (N_10965,N_9182,N_9251);
nor U10966 (N_10966,N_9604,N_9452);
nand U10967 (N_10967,N_9968,N_10402);
nand U10968 (N_10968,N_10085,N_9198);
and U10969 (N_10969,N_9929,N_10184);
and U10970 (N_10970,N_9708,N_10298);
and U10971 (N_10971,N_10007,N_9712);
and U10972 (N_10972,N_10087,N_9899);
nand U10973 (N_10973,N_10156,N_10103);
nor U10974 (N_10974,N_9596,N_9102);
or U10975 (N_10975,N_9160,N_9317);
nand U10976 (N_10976,N_10095,N_9644);
and U10977 (N_10977,N_9559,N_9503);
or U10978 (N_10978,N_9448,N_9732);
nor U10979 (N_10979,N_10194,N_10429);
or U10980 (N_10980,N_9410,N_10435);
nand U10981 (N_10981,N_9541,N_10425);
nor U10982 (N_10982,N_9131,N_10442);
or U10983 (N_10983,N_9511,N_9371);
or U10984 (N_10984,N_9344,N_10469);
or U10985 (N_10985,N_10311,N_9265);
nand U10986 (N_10986,N_9314,N_10014);
nand U10987 (N_10987,N_9930,N_10380);
xor U10988 (N_10988,N_9089,N_9248);
and U10989 (N_10989,N_9337,N_9124);
nor U10990 (N_10990,N_10053,N_10354);
nand U10991 (N_10991,N_9451,N_9037);
or U10992 (N_10992,N_10040,N_10328);
and U10993 (N_10993,N_10030,N_9720);
nor U10994 (N_10994,N_9232,N_10447);
nand U10995 (N_10995,N_9439,N_9069);
and U10996 (N_10996,N_10325,N_9292);
and U10997 (N_10997,N_9092,N_9830);
nand U10998 (N_10998,N_9854,N_9791);
xor U10999 (N_10999,N_9358,N_9920);
or U11000 (N_11000,N_10323,N_9860);
or U11001 (N_11001,N_9364,N_9229);
or U11002 (N_11002,N_9962,N_10406);
or U11003 (N_11003,N_9947,N_10465);
or U11004 (N_11004,N_9270,N_9802);
nand U11005 (N_11005,N_9303,N_9357);
nand U11006 (N_11006,N_9501,N_10229);
or U11007 (N_11007,N_9667,N_9199);
nand U11008 (N_11008,N_9633,N_10061);
or U11009 (N_11009,N_9287,N_9551);
and U11010 (N_11010,N_9231,N_10261);
or U11011 (N_11011,N_9913,N_10353);
nor U11012 (N_11012,N_9890,N_9607);
or U11013 (N_11013,N_9133,N_10141);
nand U11014 (N_11014,N_9558,N_9459);
nand U11015 (N_11015,N_9544,N_10122);
nand U11016 (N_11016,N_9924,N_9213);
nand U11017 (N_11017,N_9640,N_9525);
nor U11018 (N_11018,N_10458,N_9855);
nand U11019 (N_11019,N_10192,N_10139);
nor U11020 (N_11020,N_9321,N_9858);
nand U11021 (N_11021,N_9004,N_10018);
nor U11022 (N_11022,N_9355,N_9994);
or U11023 (N_11023,N_9804,N_9301);
or U11024 (N_11024,N_10032,N_9554);
or U11025 (N_11025,N_9842,N_9308);
or U11026 (N_11026,N_10344,N_10391);
or U11027 (N_11027,N_9077,N_9608);
nor U11028 (N_11028,N_9798,N_9462);
or U11029 (N_11029,N_10174,N_9268);
or U11030 (N_11030,N_9795,N_9540);
nand U11031 (N_11031,N_9052,N_9386);
nor U11032 (N_11032,N_10289,N_10219);
or U11033 (N_11033,N_10495,N_9391);
and U11034 (N_11034,N_10473,N_9261);
and U11035 (N_11035,N_10448,N_9370);
nor U11036 (N_11036,N_10180,N_9418);
and U11037 (N_11037,N_9394,N_9272);
nand U11038 (N_11038,N_10101,N_10159);
xor U11039 (N_11039,N_9609,N_10160);
or U11040 (N_11040,N_10274,N_9763);
nor U11041 (N_11041,N_9839,N_10462);
nand U11042 (N_11042,N_10407,N_9905);
nor U11043 (N_11043,N_9981,N_9971);
and U11044 (N_11044,N_9976,N_10186);
nor U11045 (N_11045,N_10281,N_9318);
or U11046 (N_11046,N_10008,N_9867);
nand U11047 (N_11047,N_9235,N_9155);
nor U11048 (N_11048,N_9363,N_9193);
nand U11049 (N_11049,N_10296,N_9259);
nand U11050 (N_11050,N_9910,N_9676);
nor U11051 (N_11051,N_9983,N_9202);
nand U11052 (N_11052,N_10137,N_9144);
nor U11053 (N_11053,N_9717,N_9581);
and U11054 (N_11054,N_9624,N_9586);
and U11055 (N_11055,N_9719,N_9483);
nand U11056 (N_11056,N_10411,N_10260);
or U11057 (N_11057,N_9885,N_9186);
nor U11058 (N_11058,N_9879,N_9120);
nand U11059 (N_11059,N_10054,N_9295);
and U11060 (N_11060,N_9871,N_9546);
or U11061 (N_11061,N_9299,N_9353);
and U11062 (N_11062,N_9578,N_9704);
nand U11063 (N_11063,N_9951,N_10079);
nand U11064 (N_11064,N_9190,N_10365);
and U11065 (N_11065,N_9195,N_9646);
nand U11066 (N_11066,N_9293,N_9687);
nand U11067 (N_11067,N_9223,N_9432);
and U11068 (N_11068,N_9790,N_9776);
nand U11069 (N_11069,N_9824,N_10440);
nor U11070 (N_11070,N_9135,N_9013);
nand U11071 (N_11071,N_9348,N_10231);
nand U11072 (N_11072,N_9707,N_9329);
and U11073 (N_11073,N_9989,N_9948);
nor U11074 (N_11074,N_10270,N_9171);
or U11075 (N_11075,N_9555,N_9851);
nand U11076 (N_11076,N_10387,N_9649);
or U11077 (N_11077,N_10244,N_9902);
or U11078 (N_11078,N_9868,N_9678);
and U11079 (N_11079,N_9475,N_10359);
nand U11080 (N_11080,N_10165,N_10175);
xnor U11081 (N_11081,N_10350,N_9539);
and U11082 (N_11082,N_10228,N_10388);
or U11083 (N_11083,N_9130,N_10157);
nand U11084 (N_11084,N_9241,N_9934);
xor U11085 (N_11085,N_10478,N_10183);
nor U11086 (N_11086,N_9536,N_9162);
and U11087 (N_11087,N_9347,N_9550);
or U11088 (N_11088,N_9206,N_9437);
nand U11089 (N_11089,N_9465,N_9770);
or U11090 (N_11090,N_9099,N_9387);
nand U11091 (N_11091,N_9800,N_9389);
or U11092 (N_11092,N_10349,N_10092);
and U11093 (N_11093,N_9797,N_9612);
nand U11094 (N_11094,N_9339,N_9777);
or U11095 (N_11095,N_9652,N_10341);
nand U11096 (N_11096,N_9383,N_10282);
or U11097 (N_11097,N_9711,N_9645);
and U11098 (N_11098,N_10252,N_10276);
nand U11099 (N_11099,N_9897,N_9034);
or U11100 (N_11100,N_9298,N_9497);
and U11101 (N_11101,N_9075,N_10070);
and U11102 (N_11102,N_10170,N_9076);
nor U11103 (N_11103,N_9395,N_9331);
nand U11104 (N_11104,N_9521,N_9576);
or U11105 (N_11105,N_10396,N_10069);
nor U11106 (N_11106,N_9323,N_10237);
and U11107 (N_11107,N_9094,N_10336);
nor U11108 (N_11108,N_9731,N_10212);
nand U11109 (N_11109,N_9715,N_10181);
and U11110 (N_11110,N_10264,N_9844);
or U11111 (N_11111,N_9739,N_10398);
and U11112 (N_11112,N_9471,N_10337);
nor U11113 (N_11113,N_9177,N_9307);
and U11114 (N_11114,N_10027,N_10310);
or U11115 (N_11115,N_9537,N_9327);
nor U11116 (N_11116,N_9898,N_10254);
and U11117 (N_11117,N_10102,N_9108);
or U11118 (N_11118,N_9423,N_9768);
and U11119 (N_11119,N_10000,N_9865);
or U11120 (N_11120,N_9690,N_9849);
nor U11121 (N_11121,N_9932,N_10397);
nor U11122 (N_11122,N_9564,N_9243);
nor U11123 (N_11123,N_9572,N_10230);
nor U11124 (N_11124,N_9953,N_9302);
or U11125 (N_11125,N_9754,N_9429);
nand U11126 (N_11126,N_10154,N_10346);
nor U11127 (N_11127,N_10022,N_9143);
and U11128 (N_11128,N_9334,N_10297);
nand U11129 (N_11129,N_9467,N_9049);
or U11130 (N_11130,N_9201,N_10498);
or U11131 (N_11131,N_10082,N_9496);
or U11132 (N_11132,N_9906,N_9420);
or U11133 (N_11133,N_9523,N_9221);
nor U11134 (N_11134,N_10116,N_9140);
or U11135 (N_11135,N_9531,N_9505);
nand U11136 (N_11136,N_10188,N_9178);
and U11137 (N_11137,N_10075,N_9825);
or U11138 (N_11138,N_10093,N_9872);
nor U11139 (N_11139,N_9065,N_10051);
nor U11140 (N_11140,N_9718,N_9123);
nor U11141 (N_11141,N_10161,N_10178);
and U11142 (N_11142,N_9918,N_9083);
and U11143 (N_11143,N_9264,N_9677);
nor U11144 (N_11144,N_9263,N_10338);
or U11145 (N_11145,N_10300,N_9427);
or U11146 (N_11146,N_9566,N_9935);
nor U11147 (N_11147,N_9280,N_10466);
nand U11148 (N_11148,N_9063,N_9826);
or U11149 (N_11149,N_10319,N_9486);
nand U11150 (N_11150,N_10081,N_9959);
and U11151 (N_11151,N_10307,N_10444);
and U11152 (N_11152,N_9780,N_9053);
or U11153 (N_11153,N_9746,N_9599);
nor U11154 (N_11154,N_9105,N_9016);
nor U11155 (N_11155,N_10104,N_10234);
nor U11156 (N_11156,N_9533,N_9430);
nor U11157 (N_11157,N_9240,N_9442);
or U11158 (N_11158,N_10491,N_9629);
or U11159 (N_11159,N_10005,N_10340);
nand U11160 (N_11160,N_9281,N_10418);
nand U11161 (N_11161,N_9628,N_9454);
nor U11162 (N_11162,N_10166,N_10055);
or U11163 (N_11163,N_10413,N_9811);
and U11164 (N_11164,N_10208,N_10149);
and U11165 (N_11165,N_9862,N_9941);
or U11166 (N_11166,N_9620,N_10383);
nor U11167 (N_11167,N_9509,N_10091);
and U11168 (N_11168,N_9622,N_9275);
or U11169 (N_11169,N_9703,N_9778);
nand U11170 (N_11170,N_9518,N_9476);
nor U11171 (N_11171,N_9458,N_9416);
and U11172 (N_11172,N_9151,N_9513);
or U11173 (N_11173,N_10386,N_9312);
and U11174 (N_11174,N_10489,N_9226);
nor U11175 (N_11175,N_10347,N_9575);
nand U11176 (N_11176,N_9956,N_9306);
and U11177 (N_11177,N_9733,N_9847);
nor U11178 (N_11178,N_10474,N_9530);
nor U11179 (N_11179,N_9585,N_9856);
and U11180 (N_11180,N_9350,N_10277);
or U11181 (N_11181,N_9714,N_9809);
xnor U11182 (N_11182,N_10107,N_9637);
or U11183 (N_11183,N_9527,N_9068);
nand U11184 (N_11184,N_10471,N_9580);
and U11185 (N_11185,N_9154,N_10431);
nand U11186 (N_11186,N_9132,N_9837);
and U11187 (N_11187,N_10483,N_9335);
or U11188 (N_11188,N_9928,N_10269);
nor U11189 (N_11189,N_10038,N_9560);
nor U11190 (N_11190,N_10286,N_9493);
nand U11191 (N_11191,N_9258,N_9388);
or U11192 (N_11192,N_9297,N_10235);
nand U11193 (N_11193,N_9694,N_10098);
or U11194 (N_11194,N_9122,N_10417);
or U11195 (N_11195,N_9106,N_9067);
and U11196 (N_11196,N_9817,N_10242);
nand U11197 (N_11197,N_10287,N_10147);
and U11198 (N_11198,N_9615,N_10009);
and U11199 (N_11199,N_10451,N_9219);
nor U11200 (N_11200,N_9605,N_9990);
and U11201 (N_11201,N_9208,N_10315);
nor U11202 (N_11202,N_10108,N_9516);
and U11203 (N_11203,N_10436,N_9385);
nand U11204 (N_11204,N_10017,N_9278);
and U11205 (N_11205,N_9915,N_9933);
nor U11206 (N_11206,N_9726,N_9103);
or U11207 (N_11207,N_10195,N_9831);
nand U11208 (N_11208,N_10049,N_9528);
and U11209 (N_11209,N_10042,N_9616);
xnor U11210 (N_11210,N_9749,N_10142);
nand U11211 (N_11211,N_9737,N_10026);
and U11212 (N_11212,N_9945,N_9960);
or U11213 (N_11213,N_10343,N_9643);
nor U11214 (N_11214,N_9619,N_9534);
or U11215 (N_11215,N_9237,N_9617);
nor U11216 (N_11216,N_9803,N_9583);
nor U11217 (N_11217,N_9285,N_9478);
or U11218 (N_11218,N_9009,N_10240);
nor U11219 (N_11219,N_9020,N_9880);
nand U11220 (N_11220,N_9741,N_10317);
and U11221 (N_11221,N_9681,N_10308);
nand U11222 (N_11222,N_10071,N_10096);
and U11223 (N_11223,N_9970,N_9884);
nand U11224 (N_11224,N_9224,N_10015);
xnor U11225 (N_11225,N_10334,N_9111);
and U11226 (N_11226,N_9805,N_9680);
or U11227 (N_11227,N_10335,N_10028);
nand U11228 (N_11228,N_9032,N_9463);
or U11229 (N_11229,N_9543,N_9922);
nand U11230 (N_11230,N_9926,N_10292);
and U11231 (N_11231,N_9565,N_9542);
and U11232 (N_11232,N_9188,N_9488);
nor U11233 (N_11233,N_9255,N_9098);
nand U11234 (N_11234,N_9405,N_9986);
nor U11235 (N_11235,N_9011,N_9987);
nor U11236 (N_11236,N_9807,N_10086);
nand U11237 (N_11237,N_9995,N_9789);
nor U11238 (N_11238,N_9900,N_10002);
nor U11239 (N_11239,N_9673,N_10034);
nand U11240 (N_11240,N_9026,N_10144);
and U11241 (N_11241,N_9588,N_9843);
xor U11242 (N_11242,N_9253,N_10004);
and U11243 (N_11243,N_9045,N_9003);
nand U11244 (N_11244,N_9042,N_9874);
nand U11245 (N_11245,N_10138,N_10441);
nor U11246 (N_11246,N_9482,N_9196);
and U11247 (N_11247,N_10111,N_10011);
or U11248 (N_11248,N_10291,N_10164);
nand U11249 (N_11249,N_9252,N_10119);
or U11250 (N_11250,N_10304,N_10027);
or U11251 (N_11251,N_10489,N_9164);
nand U11252 (N_11252,N_9764,N_10287);
and U11253 (N_11253,N_9072,N_9109);
nor U11254 (N_11254,N_9477,N_9529);
nand U11255 (N_11255,N_10162,N_9816);
nand U11256 (N_11256,N_10180,N_9220);
or U11257 (N_11257,N_10064,N_10257);
nand U11258 (N_11258,N_9654,N_9505);
nand U11259 (N_11259,N_9962,N_9891);
and U11260 (N_11260,N_9270,N_10363);
and U11261 (N_11261,N_10423,N_9476);
nand U11262 (N_11262,N_10005,N_9948);
or U11263 (N_11263,N_10369,N_9709);
and U11264 (N_11264,N_9797,N_9788);
nor U11265 (N_11265,N_9954,N_10115);
and U11266 (N_11266,N_10339,N_9067);
nand U11267 (N_11267,N_9884,N_10092);
and U11268 (N_11268,N_9852,N_9894);
or U11269 (N_11269,N_9907,N_9567);
nand U11270 (N_11270,N_9342,N_9228);
or U11271 (N_11271,N_9443,N_10366);
nor U11272 (N_11272,N_9071,N_9946);
nand U11273 (N_11273,N_9785,N_10235);
nand U11274 (N_11274,N_9208,N_9380);
or U11275 (N_11275,N_9371,N_9507);
or U11276 (N_11276,N_10482,N_10135);
and U11277 (N_11277,N_9638,N_9033);
and U11278 (N_11278,N_10173,N_10353);
and U11279 (N_11279,N_9331,N_9374);
nor U11280 (N_11280,N_9678,N_9451);
xor U11281 (N_11281,N_9050,N_10102);
and U11282 (N_11282,N_9153,N_9981);
and U11283 (N_11283,N_10288,N_10426);
or U11284 (N_11284,N_9029,N_10351);
and U11285 (N_11285,N_9853,N_10472);
or U11286 (N_11286,N_9935,N_9862);
and U11287 (N_11287,N_9045,N_10082);
nor U11288 (N_11288,N_9971,N_9482);
nor U11289 (N_11289,N_9862,N_9760);
nand U11290 (N_11290,N_9430,N_10267);
nand U11291 (N_11291,N_10486,N_9980);
or U11292 (N_11292,N_10033,N_9063);
nor U11293 (N_11293,N_9799,N_10443);
or U11294 (N_11294,N_9785,N_9577);
nand U11295 (N_11295,N_9127,N_10338);
nand U11296 (N_11296,N_9295,N_9621);
and U11297 (N_11297,N_9092,N_9329);
nor U11298 (N_11298,N_9052,N_10019);
nor U11299 (N_11299,N_9586,N_10440);
nor U11300 (N_11300,N_10185,N_9519);
nor U11301 (N_11301,N_9110,N_9140);
nor U11302 (N_11302,N_9352,N_9046);
or U11303 (N_11303,N_10332,N_10342);
or U11304 (N_11304,N_9340,N_9530);
nor U11305 (N_11305,N_9058,N_9023);
nand U11306 (N_11306,N_9377,N_10371);
nand U11307 (N_11307,N_9318,N_9483);
and U11308 (N_11308,N_9325,N_9567);
and U11309 (N_11309,N_9732,N_9297);
nor U11310 (N_11310,N_10015,N_10181);
nand U11311 (N_11311,N_9696,N_9341);
xor U11312 (N_11312,N_9333,N_9912);
nor U11313 (N_11313,N_10123,N_9790);
or U11314 (N_11314,N_9845,N_10321);
nor U11315 (N_11315,N_10171,N_10312);
nor U11316 (N_11316,N_9160,N_9864);
and U11317 (N_11317,N_9426,N_10006);
and U11318 (N_11318,N_9004,N_10165);
nor U11319 (N_11319,N_9091,N_10329);
and U11320 (N_11320,N_10101,N_9728);
and U11321 (N_11321,N_9129,N_9850);
nand U11322 (N_11322,N_10282,N_9444);
nand U11323 (N_11323,N_9651,N_10310);
nand U11324 (N_11324,N_10170,N_9546);
nor U11325 (N_11325,N_10150,N_10371);
and U11326 (N_11326,N_10121,N_9142);
or U11327 (N_11327,N_9017,N_9940);
nor U11328 (N_11328,N_9893,N_9621);
nor U11329 (N_11329,N_10026,N_9537);
or U11330 (N_11330,N_10324,N_9612);
nor U11331 (N_11331,N_9745,N_10411);
nor U11332 (N_11332,N_9011,N_10265);
nor U11333 (N_11333,N_9621,N_10462);
nor U11334 (N_11334,N_9912,N_9566);
nand U11335 (N_11335,N_9012,N_10447);
and U11336 (N_11336,N_9894,N_10062);
and U11337 (N_11337,N_9186,N_10413);
or U11338 (N_11338,N_9447,N_10310);
nor U11339 (N_11339,N_9297,N_9404);
or U11340 (N_11340,N_9384,N_9808);
nor U11341 (N_11341,N_10049,N_10128);
or U11342 (N_11342,N_9560,N_9029);
nand U11343 (N_11343,N_9519,N_9745);
nor U11344 (N_11344,N_9849,N_10273);
nor U11345 (N_11345,N_10351,N_9629);
or U11346 (N_11346,N_9904,N_9767);
and U11347 (N_11347,N_10324,N_10357);
and U11348 (N_11348,N_9390,N_9519);
nand U11349 (N_11349,N_9014,N_9771);
and U11350 (N_11350,N_10209,N_9596);
and U11351 (N_11351,N_10192,N_10283);
or U11352 (N_11352,N_10218,N_10311);
or U11353 (N_11353,N_9108,N_9351);
and U11354 (N_11354,N_10093,N_9985);
nor U11355 (N_11355,N_9975,N_9157);
or U11356 (N_11356,N_9751,N_9769);
or U11357 (N_11357,N_9977,N_10204);
or U11358 (N_11358,N_10461,N_9902);
and U11359 (N_11359,N_9720,N_9020);
nand U11360 (N_11360,N_9700,N_9440);
nand U11361 (N_11361,N_9767,N_9400);
nand U11362 (N_11362,N_10478,N_10319);
nand U11363 (N_11363,N_10460,N_10244);
and U11364 (N_11364,N_9397,N_9980);
nor U11365 (N_11365,N_9153,N_9921);
or U11366 (N_11366,N_9105,N_9629);
nand U11367 (N_11367,N_10283,N_10112);
nor U11368 (N_11368,N_9873,N_10072);
or U11369 (N_11369,N_9321,N_10018);
nand U11370 (N_11370,N_9596,N_9516);
and U11371 (N_11371,N_9079,N_9336);
and U11372 (N_11372,N_9200,N_9264);
and U11373 (N_11373,N_9569,N_10398);
or U11374 (N_11374,N_9632,N_10387);
or U11375 (N_11375,N_9958,N_10205);
nand U11376 (N_11376,N_10339,N_9087);
or U11377 (N_11377,N_9877,N_9843);
nor U11378 (N_11378,N_10311,N_10177);
nand U11379 (N_11379,N_9484,N_10479);
nor U11380 (N_11380,N_9605,N_9619);
or U11381 (N_11381,N_10182,N_10214);
and U11382 (N_11382,N_9056,N_9659);
or U11383 (N_11383,N_9161,N_9268);
and U11384 (N_11384,N_9152,N_9231);
nor U11385 (N_11385,N_9815,N_9626);
nand U11386 (N_11386,N_9197,N_10119);
nand U11387 (N_11387,N_10229,N_9224);
and U11388 (N_11388,N_10397,N_9344);
nand U11389 (N_11389,N_10132,N_9176);
and U11390 (N_11390,N_10013,N_10276);
or U11391 (N_11391,N_9856,N_10250);
xnor U11392 (N_11392,N_9693,N_10409);
nand U11393 (N_11393,N_9960,N_9487);
xnor U11394 (N_11394,N_9733,N_9702);
and U11395 (N_11395,N_10330,N_9322);
and U11396 (N_11396,N_9404,N_9670);
nor U11397 (N_11397,N_9096,N_9263);
and U11398 (N_11398,N_9006,N_9576);
nor U11399 (N_11399,N_9551,N_9022);
nor U11400 (N_11400,N_9014,N_10292);
nand U11401 (N_11401,N_9203,N_9806);
nand U11402 (N_11402,N_9927,N_9330);
or U11403 (N_11403,N_9422,N_9927);
and U11404 (N_11404,N_9008,N_9730);
nor U11405 (N_11405,N_9507,N_9711);
nor U11406 (N_11406,N_9295,N_9321);
or U11407 (N_11407,N_9677,N_10226);
nor U11408 (N_11408,N_9905,N_9932);
or U11409 (N_11409,N_9400,N_9963);
and U11410 (N_11410,N_9936,N_9053);
or U11411 (N_11411,N_9495,N_10468);
nand U11412 (N_11412,N_9196,N_9508);
nand U11413 (N_11413,N_9948,N_10310);
or U11414 (N_11414,N_9047,N_10446);
nand U11415 (N_11415,N_10456,N_9024);
and U11416 (N_11416,N_10183,N_9235);
nand U11417 (N_11417,N_9300,N_9872);
nand U11418 (N_11418,N_10126,N_9365);
and U11419 (N_11419,N_9355,N_9216);
nor U11420 (N_11420,N_9906,N_9880);
nor U11421 (N_11421,N_9465,N_10316);
nand U11422 (N_11422,N_10243,N_9591);
or U11423 (N_11423,N_10304,N_9194);
nand U11424 (N_11424,N_9513,N_9088);
nor U11425 (N_11425,N_9769,N_9454);
nor U11426 (N_11426,N_9818,N_9042);
nor U11427 (N_11427,N_9843,N_9618);
and U11428 (N_11428,N_9447,N_9914);
and U11429 (N_11429,N_9385,N_9492);
nand U11430 (N_11430,N_9764,N_9301);
and U11431 (N_11431,N_9410,N_10017);
nor U11432 (N_11432,N_9981,N_10256);
nand U11433 (N_11433,N_9724,N_9864);
nand U11434 (N_11434,N_9740,N_9424);
or U11435 (N_11435,N_9273,N_10110);
nand U11436 (N_11436,N_9275,N_10349);
and U11437 (N_11437,N_9802,N_9871);
and U11438 (N_11438,N_9681,N_10443);
or U11439 (N_11439,N_9485,N_9593);
nor U11440 (N_11440,N_9367,N_10414);
and U11441 (N_11441,N_9361,N_9270);
nor U11442 (N_11442,N_9778,N_9415);
nand U11443 (N_11443,N_9538,N_10128);
nand U11444 (N_11444,N_10362,N_9154);
and U11445 (N_11445,N_10000,N_10354);
or U11446 (N_11446,N_10399,N_9796);
or U11447 (N_11447,N_10212,N_9281);
and U11448 (N_11448,N_9899,N_9066);
and U11449 (N_11449,N_9446,N_9909);
nor U11450 (N_11450,N_9060,N_9154);
nor U11451 (N_11451,N_9491,N_10073);
or U11452 (N_11452,N_9504,N_10203);
nor U11453 (N_11453,N_9537,N_9997);
nand U11454 (N_11454,N_10323,N_9150);
and U11455 (N_11455,N_9657,N_9662);
nand U11456 (N_11456,N_9923,N_9407);
or U11457 (N_11457,N_10055,N_10004);
or U11458 (N_11458,N_10304,N_9095);
nand U11459 (N_11459,N_9270,N_10091);
nor U11460 (N_11460,N_10408,N_10115);
or U11461 (N_11461,N_9644,N_9587);
nor U11462 (N_11462,N_9705,N_9503);
nor U11463 (N_11463,N_10061,N_9628);
or U11464 (N_11464,N_9798,N_9506);
nor U11465 (N_11465,N_10165,N_10077);
nor U11466 (N_11466,N_9955,N_9153);
nand U11467 (N_11467,N_10187,N_9801);
nor U11468 (N_11468,N_9688,N_9188);
or U11469 (N_11469,N_9140,N_9325);
nand U11470 (N_11470,N_9716,N_10473);
nand U11471 (N_11471,N_9257,N_9284);
nor U11472 (N_11472,N_9741,N_9957);
and U11473 (N_11473,N_10474,N_10410);
nor U11474 (N_11474,N_10434,N_10427);
nor U11475 (N_11475,N_9121,N_9604);
or U11476 (N_11476,N_10430,N_9912);
nor U11477 (N_11477,N_10474,N_10480);
or U11478 (N_11478,N_10382,N_9773);
or U11479 (N_11479,N_10372,N_10094);
and U11480 (N_11480,N_9339,N_10434);
nand U11481 (N_11481,N_9153,N_9426);
nand U11482 (N_11482,N_9657,N_9154);
nand U11483 (N_11483,N_10049,N_10363);
and U11484 (N_11484,N_9856,N_9790);
and U11485 (N_11485,N_9700,N_10364);
and U11486 (N_11486,N_9123,N_9041);
nand U11487 (N_11487,N_10216,N_9135);
nor U11488 (N_11488,N_9336,N_10206);
nand U11489 (N_11489,N_9624,N_10026);
or U11490 (N_11490,N_9715,N_9597);
nor U11491 (N_11491,N_10440,N_10363);
or U11492 (N_11492,N_9698,N_10460);
xnor U11493 (N_11493,N_10010,N_9495);
and U11494 (N_11494,N_9763,N_10003);
nor U11495 (N_11495,N_10386,N_9916);
nor U11496 (N_11496,N_9582,N_9204);
nand U11497 (N_11497,N_9353,N_10164);
and U11498 (N_11498,N_10128,N_10074);
or U11499 (N_11499,N_9951,N_10461);
and U11500 (N_11500,N_9259,N_10035);
nand U11501 (N_11501,N_9555,N_9067);
nand U11502 (N_11502,N_9314,N_10380);
nand U11503 (N_11503,N_9559,N_9638);
or U11504 (N_11504,N_9503,N_9621);
or U11505 (N_11505,N_10459,N_10171);
nor U11506 (N_11506,N_10353,N_10186);
nor U11507 (N_11507,N_10165,N_10127);
xor U11508 (N_11508,N_9484,N_9053);
or U11509 (N_11509,N_9423,N_9506);
or U11510 (N_11510,N_9544,N_9618);
or U11511 (N_11511,N_9349,N_9456);
or U11512 (N_11512,N_9479,N_9816);
nand U11513 (N_11513,N_10439,N_9880);
or U11514 (N_11514,N_9167,N_10388);
or U11515 (N_11515,N_10079,N_9383);
and U11516 (N_11516,N_9864,N_10378);
nand U11517 (N_11517,N_10225,N_9381);
nor U11518 (N_11518,N_9917,N_9566);
nand U11519 (N_11519,N_10241,N_9519);
and U11520 (N_11520,N_9885,N_9675);
or U11521 (N_11521,N_10256,N_9567);
nand U11522 (N_11522,N_10221,N_10228);
and U11523 (N_11523,N_9845,N_9714);
nor U11524 (N_11524,N_9395,N_9694);
xor U11525 (N_11525,N_10276,N_10442);
nor U11526 (N_11526,N_9973,N_9662);
and U11527 (N_11527,N_9404,N_9882);
and U11528 (N_11528,N_9077,N_9682);
xnor U11529 (N_11529,N_9712,N_10441);
or U11530 (N_11530,N_9144,N_10242);
nor U11531 (N_11531,N_9671,N_10450);
nor U11532 (N_11532,N_9755,N_9341);
nand U11533 (N_11533,N_10067,N_9221);
nor U11534 (N_11534,N_10277,N_10346);
or U11535 (N_11535,N_9000,N_9446);
xor U11536 (N_11536,N_9511,N_10435);
and U11537 (N_11537,N_10234,N_10471);
nand U11538 (N_11538,N_10062,N_10465);
or U11539 (N_11539,N_9200,N_9201);
and U11540 (N_11540,N_9638,N_9042);
xnor U11541 (N_11541,N_9555,N_9407);
xnor U11542 (N_11542,N_10216,N_9684);
nor U11543 (N_11543,N_9462,N_10445);
or U11544 (N_11544,N_9046,N_9187);
or U11545 (N_11545,N_10352,N_9974);
and U11546 (N_11546,N_9912,N_10255);
or U11547 (N_11547,N_10452,N_9847);
nor U11548 (N_11548,N_9612,N_9177);
or U11549 (N_11549,N_10278,N_9486);
nor U11550 (N_11550,N_9525,N_9781);
nand U11551 (N_11551,N_9637,N_9479);
and U11552 (N_11552,N_9511,N_9215);
nor U11553 (N_11553,N_10155,N_9901);
nor U11554 (N_11554,N_9456,N_10435);
and U11555 (N_11555,N_9353,N_9538);
nand U11556 (N_11556,N_9293,N_10411);
nor U11557 (N_11557,N_9506,N_9324);
nor U11558 (N_11558,N_10027,N_10023);
nand U11559 (N_11559,N_9523,N_9638);
xnor U11560 (N_11560,N_10232,N_9845);
or U11561 (N_11561,N_9663,N_9269);
and U11562 (N_11562,N_10210,N_9046);
nand U11563 (N_11563,N_9517,N_9701);
nor U11564 (N_11564,N_9670,N_10022);
and U11565 (N_11565,N_9506,N_9914);
and U11566 (N_11566,N_10198,N_10239);
nand U11567 (N_11567,N_9680,N_10097);
nor U11568 (N_11568,N_9398,N_9969);
or U11569 (N_11569,N_9329,N_9036);
and U11570 (N_11570,N_9636,N_9058);
xnor U11571 (N_11571,N_9808,N_10298);
or U11572 (N_11572,N_10348,N_9802);
nand U11573 (N_11573,N_9251,N_10073);
nand U11574 (N_11574,N_10093,N_9694);
nand U11575 (N_11575,N_9358,N_10159);
xor U11576 (N_11576,N_9036,N_9225);
or U11577 (N_11577,N_9495,N_10312);
nand U11578 (N_11578,N_9444,N_9603);
and U11579 (N_11579,N_10268,N_9416);
nand U11580 (N_11580,N_10074,N_9872);
and U11581 (N_11581,N_9211,N_9574);
or U11582 (N_11582,N_10131,N_9946);
nand U11583 (N_11583,N_9834,N_9561);
nor U11584 (N_11584,N_9408,N_10321);
nor U11585 (N_11585,N_9193,N_10462);
nand U11586 (N_11586,N_9052,N_9003);
nor U11587 (N_11587,N_10019,N_10091);
nor U11588 (N_11588,N_9081,N_10349);
and U11589 (N_11589,N_9655,N_9705);
nand U11590 (N_11590,N_9188,N_9933);
nand U11591 (N_11591,N_10124,N_9709);
nand U11592 (N_11592,N_9717,N_10211);
or U11593 (N_11593,N_9121,N_9178);
nand U11594 (N_11594,N_9904,N_9967);
nand U11595 (N_11595,N_9287,N_9778);
or U11596 (N_11596,N_10474,N_10297);
nand U11597 (N_11597,N_9426,N_9471);
and U11598 (N_11598,N_9403,N_9923);
nor U11599 (N_11599,N_9401,N_9200);
or U11600 (N_11600,N_9341,N_10430);
and U11601 (N_11601,N_9097,N_9686);
nand U11602 (N_11602,N_9432,N_9887);
or U11603 (N_11603,N_9359,N_10322);
or U11604 (N_11604,N_9815,N_9786);
and U11605 (N_11605,N_10231,N_10495);
or U11606 (N_11606,N_10088,N_10431);
nor U11607 (N_11607,N_9315,N_9097);
and U11608 (N_11608,N_9801,N_9355);
nor U11609 (N_11609,N_9348,N_9231);
or U11610 (N_11610,N_9769,N_10471);
and U11611 (N_11611,N_10032,N_9607);
and U11612 (N_11612,N_9368,N_9030);
xnor U11613 (N_11613,N_9928,N_9420);
and U11614 (N_11614,N_9121,N_9099);
or U11615 (N_11615,N_9806,N_9324);
or U11616 (N_11616,N_10334,N_10155);
nor U11617 (N_11617,N_10459,N_9084);
or U11618 (N_11618,N_10079,N_10284);
and U11619 (N_11619,N_9814,N_9346);
or U11620 (N_11620,N_10402,N_9128);
and U11621 (N_11621,N_9276,N_9458);
xnor U11622 (N_11622,N_9959,N_9032);
nand U11623 (N_11623,N_9340,N_9213);
and U11624 (N_11624,N_9094,N_9980);
and U11625 (N_11625,N_10304,N_9791);
nand U11626 (N_11626,N_9644,N_10244);
nor U11627 (N_11627,N_10464,N_10198);
nand U11628 (N_11628,N_10322,N_9325);
and U11629 (N_11629,N_9428,N_9182);
or U11630 (N_11630,N_10126,N_9679);
and U11631 (N_11631,N_10034,N_10101);
nor U11632 (N_11632,N_10195,N_10247);
or U11633 (N_11633,N_9314,N_9597);
and U11634 (N_11634,N_9104,N_10230);
or U11635 (N_11635,N_9163,N_10361);
or U11636 (N_11636,N_9494,N_9124);
or U11637 (N_11637,N_9231,N_9854);
nand U11638 (N_11638,N_10397,N_10033);
nand U11639 (N_11639,N_9799,N_9943);
and U11640 (N_11640,N_10142,N_9774);
nand U11641 (N_11641,N_9055,N_9181);
nand U11642 (N_11642,N_9740,N_10422);
or U11643 (N_11643,N_9527,N_9213);
and U11644 (N_11644,N_10032,N_9763);
nand U11645 (N_11645,N_9621,N_9285);
and U11646 (N_11646,N_9265,N_10029);
or U11647 (N_11647,N_10295,N_10212);
and U11648 (N_11648,N_9150,N_9688);
and U11649 (N_11649,N_10002,N_9791);
or U11650 (N_11650,N_9967,N_9452);
or U11651 (N_11651,N_10385,N_10235);
and U11652 (N_11652,N_10005,N_9117);
nor U11653 (N_11653,N_9693,N_9442);
nor U11654 (N_11654,N_9899,N_10068);
nor U11655 (N_11655,N_9678,N_9671);
or U11656 (N_11656,N_9138,N_10285);
or U11657 (N_11657,N_9118,N_10451);
nor U11658 (N_11658,N_10277,N_9628);
and U11659 (N_11659,N_9913,N_9763);
and U11660 (N_11660,N_10115,N_9620);
nor U11661 (N_11661,N_9379,N_9833);
and U11662 (N_11662,N_9263,N_9559);
or U11663 (N_11663,N_10178,N_9195);
and U11664 (N_11664,N_9795,N_9645);
nand U11665 (N_11665,N_9564,N_9525);
nand U11666 (N_11666,N_10485,N_10242);
or U11667 (N_11667,N_9396,N_10045);
nand U11668 (N_11668,N_10457,N_9205);
nand U11669 (N_11669,N_10482,N_10490);
nor U11670 (N_11670,N_9505,N_10349);
or U11671 (N_11671,N_10007,N_10411);
or U11672 (N_11672,N_9997,N_9976);
or U11673 (N_11673,N_9324,N_10392);
and U11674 (N_11674,N_10363,N_9328);
nand U11675 (N_11675,N_9652,N_10463);
or U11676 (N_11676,N_9984,N_9637);
or U11677 (N_11677,N_10470,N_9334);
nand U11678 (N_11678,N_9998,N_10291);
nand U11679 (N_11679,N_10334,N_9314);
xor U11680 (N_11680,N_9231,N_10467);
and U11681 (N_11681,N_9943,N_9481);
nand U11682 (N_11682,N_9282,N_9982);
nand U11683 (N_11683,N_10440,N_10177);
nor U11684 (N_11684,N_9353,N_9199);
and U11685 (N_11685,N_9671,N_9284);
or U11686 (N_11686,N_10216,N_9874);
nor U11687 (N_11687,N_9746,N_9964);
nand U11688 (N_11688,N_9830,N_9989);
nor U11689 (N_11689,N_10100,N_10164);
nor U11690 (N_11690,N_9424,N_9316);
and U11691 (N_11691,N_9131,N_9334);
or U11692 (N_11692,N_9232,N_9338);
or U11693 (N_11693,N_9250,N_9772);
and U11694 (N_11694,N_9485,N_9951);
or U11695 (N_11695,N_9398,N_9744);
and U11696 (N_11696,N_9365,N_9493);
and U11697 (N_11697,N_10076,N_9066);
or U11698 (N_11698,N_9264,N_9290);
or U11699 (N_11699,N_10413,N_9064);
nor U11700 (N_11700,N_9327,N_9733);
xnor U11701 (N_11701,N_9634,N_9554);
nor U11702 (N_11702,N_9909,N_10245);
nor U11703 (N_11703,N_9268,N_10436);
nand U11704 (N_11704,N_9896,N_9194);
nor U11705 (N_11705,N_10040,N_9179);
nand U11706 (N_11706,N_9225,N_9260);
and U11707 (N_11707,N_10289,N_9118);
nand U11708 (N_11708,N_9243,N_10116);
or U11709 (N_11709,N_9322,N_9664);
nor U11710 (N_11710,N_10007,N_9616);
nor U11711 (N_11711,N_9587,N_9375);
nand U11712 (N_11712,N_9783,N_9044);
or U11713 (N_11713,N_10490,N_9992);
nor U11714 (N_11714,N_10336,N_10395);
nand U11715 (N_11715,N_9185,N_9989);
and U11716 (N_11716,N_9021,N_9783);
or U11717 (N_11717,N_9111,N_9097);
nor U11718 (N_11718,N_9578,N_9001);
and U11719 (N_11719,N_9043,N_10335);
nand U11720 (N_11720,N_9203,N_10148);
nand U11721 (N_11721,N_10151,N_9698);
nand U11722 (N_11722,N_9187,N_9153);
or U11723 (N_11723,N_10210,N_9099);
nor U11724 (N_11724,N_10458,N_9833);
and U11725 (N_11725,N_9586,N_10219);
nand U11726 (N_11726,N_9545,N_9030);
nand U11727 (N_11727,N_10241,N_9893);
xor U11728 (N_11728,N_10075,N_9958);
nand U11729 (N_11729,N_9246,N_9782);
nand U11730 (N_11730,N_9220,N_9032);
and U11731 (N_11731,N_9944,N_10247);
nand U11732 (N_11732,N_10044,N_9478);
nor U11733 (N_11733,N_9218,N_9534);
nor U11734 (N_11734,N_10248,N_10057);
or U11735 (N_11735,N_9600,N_9426);
nand U11736 (N_11736,N_9794,N_10082);
nor U11737 (N_11737,N_10159,N_10102);
nand U11738 (N_11738,N_9903,N_9604);
nand U11739 (N_11739,N_9460,N_9108);
nor U11740 (N_11740,N_10399,N_10430);
nor U11741 (N_11741,N_9488,N_10298);
xnor U11742 (N_11742,N_9329,N_9502);
and U11743 (N_11743,N_9488,N_10246);
or U11744 (N_11744,N_9795,N_9704);
nor U11745 (N_11745,N_9481,N_9131);
nand U11746 (N_11746,N_9043,N_10334);
xor U11747 (N_11747,N_9984,N_9366);
or U11748 (N_11748,N_10087,N_9583);
nor U11749 (N_11749,N_9766,N_10418);
and U11750 (N_11750,N_9987,N_9044);
or U11751 (N_11751,N_10087,N_9447);
nor U11752 (N_11752,N_9585,N_10007);
nand U11753 (N_11753,N_10304,N_9860);
or U11754 (N_11754,N_9395,N_10449);
and U11755 (N_11755,N_10332,N_10372);
or U11756 (N_11756,N_10351,N_9774);
and U11757 (N_11757,N_10095,N_9790);
nor U11758 (N_11758,N_10269,N_9898);
nor U11759 (N_11759,N_10356,N_9531);
nand U11760 (N_11760,N_9411,N_10074);
and U11761 (N_11761,N_9099,N_10115);
nand U11762 (N_11762,N_9910,N_10127);
or U11763 (N_11763,N_10273,N_10004);
or U11764 (N_11764,N_9140,N_10458);
nor U11765 (N_11765,N_9671,N_9343);
and U11766 (N_11766,N_9355,N_10476);
nor U11767 (N_11767,N_9022,N_9143);
or U11768 (N_11768,N_9729,N_9594);
or U11769 (N_11769,N_9072,N_9559);
or U11770 (N_11770,N_9784,N_9022);
or U11771 (N_11771,N_9242,N_9801);
or U11772 (N_11772,N_10318,N_9457);
or U11773 (N_11773,N_9949,N_9200);
or U11774 (N_11774,N_9876,N_10342);
nand U11775 (N_11775,N_10400,N_10262);
or U11776 (N_11776,N_10330,N_9852);
nor U11777 (N_11777,N_10112,N_10238);
nor U11778 (N_11778,N_9841,N_9936);
nand U11779 (N_11779,N_9549,N_9272);
or U11780 (N_11780,N_9807,N_9255);
nor U11781 (N_11781,N_9222,N_10241);
nor U11782 (N_11782,N_9630,N_9968);
and U11783 (N_11783,N_9491,N_9104);
and U11784 (N_11784,N_9627,N_10185);
xor U11785 (N_11785,N_9886,N_9795);
nand U11786 (N_11786,N_9913,N_9574);
nand U11787 (N_11787,N_9143,N_9096);
nand U11788 (N_11788,N_9229,N_9490);
or U11789 (N_11789,N_10471,N_10210);
nor U11790 (N_11790,N_9236,N_10491);
or U11791 (N_11791,N_10103,N_9803);
or U11792 (N_11792,N_9747,N_10171);
or U11793 (N_11793,N_10355,N_9192);
and U11794 (N_11794,N_9400,N_9353);
and U11795 (N_11795,N_9975,N_9025);
and U11796 (N_11796,N_10306,N_9670);
or U11797 (N_11797,N_9443,N_10283);
and U11798 (N_11798,N_9359,N_9966);
or U11799 (N_11799,N_9660,N_9444);
or U11800 (N_11800,N_9427,N_9415);
or U11801 (N_11801,N_10440,N_9175);
nor U11802 (N_11802,N_9856,N_10464);
and U11803 (N_11803,N_9823,N_9071);
or U11804 (N_11804,N_10074,N_9483);
nand U11805 (N_11805,N_9390,N_9669);
nor U11806 (N_11806,N_10287,N_9424);
nor U11807 (N_11807,N_9905,N_9958);
nor U11808 (N_11808,N_10312,N_9259);
or U11809 (N_11809,N_9911,N_10372);
nor U11810 (N_11810,N_10356,N_9492);
and U11811 (N_11811,N_10322,N_9940);
or U11812 (N_11812,N_9975,N_9415);
nor U11813 (N_11813,N_9801,N_9553);
nand U11814 (N_11814,N_10403,N_9499);
nor U11815 (N_11815,N_9336,N_9973);
and U11816 (N_11816,N_9593,N_9318);
xnor U11817 (N_11817,N_9390,N_10489);
and U11818 (N_11818,N_9127,N_9874);
nor U11819 (N_11819,N_9982,N_9328);
xor U11820 (N_11820,N_9784,N_9087);
nand U11821 (N_11821,N_9515,N_9230);
nand U11822 (N_11822,N_9680,N_10050);
nor U11823 (N_11823,N_9720,N_9261);
or U11824 (N_11824,N_10135,N_9239);
nor U11825 (N_11825,N_9295,N_10107);
and U11826 (N_11826,N_9337,N_9440);
or U11827 (N_11827,N_9133,N_10381);
or U11828 (N_11828,N_9462,N_9338);
or U11829 (N_11829,N_9393,N_9675);
or U11830 (N_11830,N_10316,N_9091);
and U11831 (N_11831,N_10098,N_10082);
and U11832 (N_11832,N_10154,N_10242);
nand U11833 (N_11833,N_10169,N_9360);
nor U11834 (N_11834,N_9268,N_9330);
and U11835 (N_11835,N_10035,N_9269);
and U11836 (N_11836,N_9290,N_9550);
nor U11837 (N_11837,N_9238,N_9906);
nand U11838 (N_11838,N_9276,N_9050);
nor U11839 (N_11839,N_9390,N_10493);
and U11840 (N_11840,N_9966,N_10189);
or U11841 (N_11841,N_9210,N_9862);
and U11842 (N_11842,N_9021,N_9686);
nor U11843 (N_11843,N_9521,N_9704);
or U11844 (N_11844,N_9123,N_9268);
or U11845 (N_11845,N_10395,N_10110);
or U11846 (N_11846,N_10377,N_10402);
xnor U11847 (N_11847,N_9313,N_9450);
and U11848 (N_11848,N_10242,N_10499);
or U11849 (N_11849,N_9380,N_10340);
or U11850 (N_11850,N_9767,N_9023);
or U11851 (N_11851,N_9204,N_9595);
and U11852 (N_11852,N_9394,N_9428);
nor U11853 (N_11853,N_9619,N_9266);
nor U11854 (N_11854,N_10349,N_9022);
nor U11855 (N_11855,N_9565,N_9278);
nand U11856 (N_11856,N_9600,N_10419);
nor U11857 (N_11857,N_9061,N_9472);
and U11858 (N_11858,N_10390,N_9451);
nor U11859 (N_11859,N_10337,N_9402);
and U11860 (N_11860,N_9568,N_9624);
nand U11861 (N_11861,N_10363,N_9139);
nor U11862 (N_11862,N_10274,N_9688);
and U11863 (N_11863,N_9361,N_9117);
nand U11864 (N_11864,N_9100,N_9448);
nor U11865 (N_11865,N_9613,N_9029);
or U11866 (N_11866,N_9412,N_9330);
xnor U11867 (N_11867,N_10032,N_10249);
and U11868 (N_11868,N_9572,N_10186);
or U11869 (N_11869,N_10253,N_9945);
nor U11870 (N_11870,N_9129,N_9540);
nand U11871 (N_11871,N_10366,N_9126);
nand U11872 (N_11872,N_10271,N_9273);
nand U11873 (N_11873,N_10476,N_9556);
or U11874 (N_11874,N_9794,N_9377);
or U11875 (N_11875,N_9529,N_9738);
nor U11876 (N_11876,N_9251,N_10160);
nand U11877 (N_11877,N_10074,N_9838);
nor U11878 (N_11878,N_10244,N_9782);
nand U11879 (N_11879,N_9287,N_10415);
nor U11880 (N_11880,N_9798,N_10488);
nand U11881 (N_11881,N_9408,N_9311);
or U11882 (N_11882,N_9131,N_10250);
nand U11883 (N_11883,N_10497,N_9676);
nor U11884 (N_11884,N_9571,N_9300);
nor U11885 (N_11885,N_9170,N_9494);
or U11886 (N_11886,N_9648,N_10401);
or U11887 (N_11887,N_9716,N_9663);
or U11888 (N_11888,N_10267,N_10236);
and U11889 (N_11889,N_10350,N_9140);
nand U11890 (N_11890,N_9932,N_10143);
and U11891 (N_11891,N_9394,N_9205);
xnor U11892 (N_11892,N_9849,N_9598);
and U11893 (N_11893,N_9318,N_10013);
or U11894 (N_11894,N_9111,N_9205);
and U11895 (N_11895,N_9163,N_10016);
nor U11896 (N_11896,N_10123,N_9941);
and U11897 (N_11897,N_9706,N_10018);
nand U11898 (N_11898,N_9385,N_10205);
and U11899 (N_11899,N_10325,N_9256);
nand U11900 (N_11900,N_9586,N_9673);
or U11901 (N_11901,N_10328,N_9271);
nand U11902 (N_11902,N_10340,N_9212);
nand U11903 (N_11903,N_10156,N_9192);
and U11904 (N_11904,N_9003,N_9093);
or U11905 (N_11905,N_9216,N_9736);
and U11906 (N_11906,N_9063,N_9092);
and U11907 (N_11907,N_10057,N_9163);
or U11908 (N_11908,N_9082,N_9652);
and U11909 (N_11909,N_9709,N_9228);
xor U11910 (N_11910,N_9351,N_10184);
nand U11911 (N_11911,N_10166,N_9389);
nand U11912 (N_11912,N_9620,N_9197);
and U11913 (N_11913,N_9667,N_9683);
nand U11914 (N_11914,N_9223,N_10364);
or U11915 (N_11915,N_9675,N_9886);
nand U11916 (N_11916,N_9178,N_9980);
nand U11917 (N_11917,N_9276,N_10263);
nor U11918 (N_11918,N_9013,N_9014);
nor U11919 (N_11919,N_10493,N_9711);
xor U11920 (N_11920,N_9087,N_9734);
and U11921 (N_11921,N_10426,N_10032);
nand U11922 (N_11922,N_9644,N_9383);
and U11923 (N_11923,N_9268,N_10156);
or U11924 (N_11924,N_9273,N_9719);
nor U11925 (N_11925,N_9024,N_10226);
nor U11926 (N_11926,N_10032,N_9022);
or U11927 (N_11927,N_9120,N_9017);
nor U11928 (N_11928,N_10416,N_10339);
and U11929 (N_11929,N_9203,N_9057);
nand U11930 (N_11930,N_9633,N_9407);
and U11931 (N_11931,N_9230,N_10371);
or U11932 (N_11932,N_9587,N_10166);
and U11933 (N_11933,N_9371,N_9423);
or U11934 (N_11934,N_10067,N_9884);
or U11935 (N_11935,N_10293,N_9572);
or U11936 (N_11936,N_9408,N_9299);
or U11937 (N_11937,N_10320,N_10331);
nand U11938 (N_11938,N_10374,N_9723);
nand U11939 (N_11939,N_9780,N_9795);
and U11940 (N_11940,N_10218,N_10403);
nand U11941 (N_11941,N_9977,N_9621);
nand U11942 (N_11942,N_10497,N_9481);
nor U11943 (N_11943,N_9293,N_9594);
or U11944 (N_11944,N_10392,N_9405);
nand U11945 (N_11945,N_9950,N_9002);
xnor U11946 (N_11946,N_9397,N_9914);
nand U11947 (N_11947,N_10217,N_10441);
nand U11948 (N_11948,N_9535,N_9367);
or U11949 (N_11949,N_9354,N_9074);
and U11950 (N_11950,N_9967,N_9399);
xor U11951 (N_11951,N_10126,N_10242);
and U11952 (N_11952,N_10337,N_10143);
and U11953 (N_11953,N_9961,N_9989);
and U11954 (N_11954,N_9742,N_10412);
and U11955 (N_11955,N_9227,N_9333);
nand U11956 (N_11956,N_10129,N_9117);
and U11957 (N_11957,N_9056,N_9389);
and U11958 (N_11958,N_9475,N_9026);
nand U11959 (N_11959,N_9313,N_9783);
nor U11960 (N_11960,N_9992,N_10243);
nand U11961 (N_11961,N_9696,N_10096);
nor U11962 (N_11962,N_9176,N_10183);
and U11963 (N_11963,N_9984,N_9524);
nor U11964 (N_11964,N_9978,N_10343);
or U11965 (N_11965,N_9097,N_10070);
nand U11966 (N_11966,N_9714,N_10101);
or U11967 (N_11967,N_9724,N_10211);
and U11968 (N_11968,N_9106,N_9983);
xor U11969 (N_11969,N_9752,N_10425);
and U11970 (N_11970,N_9761,N_9809);
or U11971 (N_11971,N_9347,N_10317);
or U11972 (N_11972,N_9603,N_9698);
or U11973 (N_11973,N_9723,N_9118);
xor U11974 (N_11974,N_9165,N_9475);
nor U11975 (N_11975,N_9594,N_9642);
nor U11976 (N_11976,N_10119,N_9000);
nand U11977 (N_11977,N_9314,N_9834);
nand U11978 (N_11978,N_10106,N_9569);
nand U11979 (N_11979,N_9414,N_9965);
nor U11980 (N_11980,N_9717,N_9961);
or U11981 (N_11981,N_9267,N_9515);
and U11982 (N_11982,N_9733,N_9120);
or U11983 (N_11983,N_9277,N_9762);
nand U11984 (N_11984,N_9959,N_9291);
nand U11985 (N_11985,N_10075,N_9069);
nor U11986 (N_11986,N_10118,N_9932);
nand U11987 (N_11987,N_9107,N_9327);
nand U11988 (N_11988,N_10079,N_9528);
and U11989 (N_11989,N_9942,N_9217);
or U11990 (N_11990,N_9411,N_10117);
or U11991 (N_11991,N_9009,N_10033);
and U11992 (N_11992,N_10077,N_9977);
xnor U11993 (N_11993,N_9985,N_9560);
or U11994 (N_11994,N_10303,N_9976);
or U11995 (N_11995,N_10400,N_9825);
nand U11996 (N_11996,N_10008,N_9043);
and U11997 (N_11997,N_10098,N_10300);
nand U11998 (N_11998,N_9967,N_9761);
or U11999 (N_11999,N_9046,N_9256);
and U12000 (N_12000,N_10979,N_10949);
nand U12001 (N_12001,N_11760,N_10519);
and U12002 (N_12002,N_11738,N_11773);
and U12003 (N_12003,N_11411,N_10945);
nor U12004 (N_12004,N_10881,N_10757);
nand U12005 (N_12005,N_11143,N_11049);
nor U12006 (N_12006,N_11901,N_10775);
nand U12007 (N_12007,N_10729,N_10649);
nor U12008 (N_12008,N_11160,N_11612);
and U12009 (N_12009,N_11187,N_11702);
nand U12010 (N_12010,N_11636,N_11899);
nor U12011 (N_12011,N_10817,N_11585);
and U12012 (N_12012,N_11793,N_10603);
nand U12013 (N_12013,N_11964,N_11848);
nand U12014 (N_12014,N_11939,N_11279);
nor U12015 (N_12015,N_11204,N_11764);
and U12016 (N_12016,N_11463,N_11507);
or U12017 (N_12017,N_11545,N_10517);
nand U12018 (N_12018,N_10666,N_10552);
or U12019 (N_12019,N_10574,N_10963);
or U12020 (N_12020,N_11883,N_11405);
xor U12021 (N_12021,N_11308,N_11126);
nand U12022 (N_12022,N_11863,N_10950);
nor U12023 (N_12023,N_10832,N_11010);
or U12024 (N_12024,N_10710,N_10610);
nor U12025 (N_12025,N_11697,N_11805);
or U12026 (N_12026,N_11392,N_10650);
nor U12027 (N_12027,N_11814,N_10762);
nand U12028 (N_12028,N_10774,N_11567);
nor U12029 (N_12029,N_10670,N_11844);
nand U12030 (N_12030,N_11243,N_11025);
nor U12031 (N_12031,N_11448,N_10618);
and U12032 (N_12032,N_10581,N_11783);
or U12033 (N_12033,N_11840,N_11709);
or U12034 (N_12034,N_11277,N_11623);
nor U12035 (N_12035,N_10596,N_10772);
or U12036 (N_12036,N_11298,N_11048);
nor U12037 (N_12037,N_10630,N_11947);
or U12038 (N_12038,N_11089,N_10663);
or U12039 (N_12039,N_11260,N_10905);
and U12040 (N_12040,N_11787,N_11123);
or U12041 (N_12041,N_11789,N_11798);
or U12042 (N_12042,N_11186,N_11924);
and U12043 (N_12043,N_10977,N_10955);
and U12044 (N_12044,N_11889,N_11085);
nand U12045 (N_12045,N_11822,N_11181);
nor U12046 (N_12046,N_10940,N_11198);
nand U12047 (N_12047,N_11053,N_11063);
nor U12048 (N_12048,N_11843,N_11541);
nand U12049 (N_12049,N_10944,N_10564);
and U12050 (N_12050,N_11965,N_11564);
or U12051 (N_12051,N_11978,N_10628);
nor U12052 (N_12052,N_11443,N_11679);
nor U12053 (N_12053,N_11346,N_11894);
and U12054 (N_12054,N_11271,N_10681);
nor U12055 (N_12055,N_11573,N_10759);
or U12056 (N_12056,N_10820,N_11111);
nand U12057 (N_12057,N_10995,N_10608);
xor U12058 (N_12058,N_11719,N_10962);
nand U12059 (N_12059,N_10981,N_11933);
nand U12060 (N_12060,N_10993,N_10657);
and U12061 (N_12061,N_11873,N_11634);
and U12062 (N_12062,N_11452,N_11743);
nand U12063 (N_12063,N_11390,N_10859);
and U12064 (N_12064,N_11399,N_10813);
nand U12065 (N_12065,N_10588,N_11687);
and U12066 (N_12066,N_11627,N_10855);
nor U12067 (N_12067,N_11533,N_11218);
and U12068 (N_12068,N_10727,N_10957);
nand U12069 (N_12069,N_10599,N_11115);
or U12070 (N_12070,N_11625,N_10508);
nor U12071 (N_12071,N_11985,N_11436);
nor U12072 (N_12072,N_10640,N_10819);
nand U12073 (N_12073,N_10732,N_11890);
nor U12074 (N_12074,N_11992,N_11414);
or U12075 (N_12075,N_11437,N_11553);
nand U12076 (N_12076,N_11487,N_10936);
nor U12077 (N_12077,N_11846,N_11145);
and U12078 (N_12078,N_11159,N_11594);
or U12079 (N_12079,N_11895,N_11214);
nor U12080 (N_12080,N_10680,N_11715);
or U12081 (N_12081,N_10857,N_11945);
and U12082 (N_12082,N_10810,N_10792);
and U12083 (N_12083,N_10842,N_11907);
or U12084 (N_12084,N_11182,N_10569);
or U12085 (N_12085,N_11620,N_10789);
nand U12086 (N_12086,N_10948,N_11130);
nand U12087 (N_12087,N_11402,N_10753);
and U12088 (N_12088,N_10823,N_10966);
or U12089 (N_12089,N_11338,N_11774);
nand U12090 (N_12090,N_10777,N_10869);
nand U12091 (N_12091,N_10804,N_10685);
and U12092 (N_12092,N_11090,N_10559);
nor U12093 (N_12093,N_10626,N_11097);
and U12094 (N_12094,N_11489,N_11450);
xor U12095 (N_12095,N_11818,N_11231);
nor U12096 (N_12096,N_11305,N_11456);
nor U12097 (N_12097,N_11297,N_10562);
or U12098 (N_12098,N_11096,N_10746);
nand U12099 (N_12099,N_10873,N_11142);
xor U12100 (N_12100,N_11370,N_11642);
or U12101 (N_12101,N_10891,N_10744);
nor U12102 (N_12102,N_11762,N_11014);
and U12103 (N_12103,N_11953,N_11935);
nor U12104 (N_12104,N_11660,N_11575);
nor U12105 (N_12105,N_11156,N_11853);
or U12106 (N_12106,N_10637,N_11113);
and U12107 (N_12107,N_11577,N_10926);
or U12108 (N_12108,N_10512,N_11672);
nand U12109 (N_12109,N_10511,N_11395);
nand U12110 (N_12110,N_10971,N_11195);
nand U12111 (N_12111,N_11849,N_11257);
nand U12112 (N_12112,N_11815,N_11175);
and U12113 (N_12113,N_11912,N_11385);
nand U12114 (N_12114,N_11024,N_11886);
nor U12115 (N_12115,N_10654,N_11432);
or U12116 (N_12116,N_10695,N_10809);
nor U12117 (N_12117,N_11373,N_11102);
nor U12118 (N_12118,N_10551,N_11607);
or U12119 (N_12119,N_11695,N_11483);
and U12120 (N_12120,N_11066,N_11713);
nor U12121 (N_12121,N_11230,N_10540);
xnor U12122 (N_12122,N_11203,N_11251);
and U12123 (N_12123,N_11601,N_11735);
nand U12124 (N_12124,N_11957,N_11219);
nor U12125 (N_12125,N_11286,N_11800);
or U12126 (N_12126,N_10973,N_10560);
and U12127 (N_12127,N_11348,N_11602);
nor U12128 (N_12128,N_10707,N_11600);
nand U12129 (N_12129,N_11887,N_10808);
nor U12130 (N_12130,N_11670,N_11427);
and U12131 (N_12131,N_10684,N_11882);
nand U12132 (N_12132,N_10668,N_10518);
and U12133 (N_12133,N_11624,N_11301);
or U12134 (N_12134,N_11059,N_11644);
nor U12135 (N_12135,N_10754,N_10880);
or U12136 (N_12136,N_10935,N_11689);
and U12137 (N_12137,N_11942,N_11124);
and U12138 (N_12138,N_11898,N_11484);
nand U12139 (N_12139,N_11550,N_11572);
or U12140 (N_12140,N_11633,N_10565);
nand U12141 (N_12141,N_11897,N_11529);
and U12142 (N_12142,N_10954,N_10682);
or U12143 (N_12143,N_10605,N_11310);
nand U12144 (N_12144,N_11663,N_11329);
and U12145 (N_12145,N_10535,N_11710);
or U12146 (N_12146,N_11866,N_10634);
xnor U12147 (N_12147,N_10716,N_11439);
and U12148 (N_12148,N_11144,N_11613);
or U12149 (N_12149,N_11080,N_10738);
or U12150 (N_12150,N_11701,N_11556);
or U12151 (N_12151,N_11369,N_11128);
nand U12152 (N_12152,N_10805,N_11054);
nor U12153 (N_12153,N_11064,N_11692);
and U12154 (N_12154,N_10632,N_11604);
nor U12155 (N_12155,N_11970,N_11536);
and U12156 (N_12156,N_11287,N_11929);
nor U12157 (N_12157,N_11470,N_11363);
and U12158 (N_12158,N_11632,N_11176);
nor U12159 (N_12159,N_11065,N_10718);
or U12160 (N_12160,N_11311,N_11500);
nand U12161 (N_12161,N_10982,N_10943);
nor U12162 (N_12162,N_10504,N_11209);
or U12163 (N_12163,N_10725,N_11360);
or U12164 (N_12164,N_11649,N_10665);
xor U12165 (N_12165,N_11502,N_10721);
nand U12166 (N_12166,N_11611,N_11685);
nor U12167 (N_12167,N_11700,N_11676);
and U12168 (N_12168,N_10633,N_10723);
or U12169 (N_12169,N_11595,N_11727);
xor U12170 (N_12170,N_11501,N_10801);
or U12171 (N_12171,N_11269,N_11398);
xor U12172 (N_12172,N_11668,N_11121);
nand U12173 (N_12173,N_11491,N_10876);
nor U12174 (N_12174,N_11292,N_11016);
nand U12175 (N_12175,N_11998,N_11823);
nor U12176 (N_12176,N_11780,N_11629);
or U12177 (N_12177,N_11009,N_11256);
nand U12178 (N_12178,N_10697,N_11655);
and U12179 (N_12179,N_11433,N_10745);
or U12180 (N_12180,N_10699,N_10598);
or U12181 (N_12181,N_11653,N_10712);
or U12182 (N_12182,N_11605,N_10748);
or U12183 (N_12183,N_11696,N_10816);
nand U12184 (N_12184,N_11011,N_10641);
or U12185 (N_12185,N_11495,N_10829);
and U12186 (N_12186,N_11029,N_10896);
nor U12187 (N_12187,N_11261,N_11274);
nor U12188 (N_12188,N_11132,N_11309);
and U12189 (N_12189,N_11387,N_11656);
or U12190 (N_12190,N_10899,N_11751);
nand U12191 (N_12191,N_11569,N_10768);
or U12192 (N_12192,N_11313,N_11913);
nand U12193 (N_12193,N_10764,N_11083);
and U12194 (N_12194,N_10545,N_11996);
or U12195 (N_12195,N_10990,N_10514);
nor U12196 (N_12196,N_10992,N_10568);
or U12197 (N_12197,N_11919,N_11799);
and U12198 (N_12198,N_10534,N_10527);
nand U12199 (N_12199,N_11020,N_11651);
and U12200 (N_12200,N_10659,N_11834);
and U12201 (N_12201,N_10701,N_11087);
or U12202 (N_12202,N_11587,N_11878);
nor U12203 (N_12203,N_11180,N_10904);
nor U12204 (N_12204,N_10578,N_10742);
or U12205 (N_12205,N_11455,N_11961);
nor U12206 (N_12206,N_10501,N_11816);
and U12207 (N_12207,N_10509,N_10690);
or U12208 (N_12208,N_11474,N_11225);
xnor U12209 (N_12209,N_11974,N_10591);
nand U12210 (N_12210,N_11892,N_11152);
or U12211 (N_12211,N_11317,N_11103);
nor U12212 (N_12212,N_11170,N_10622);
and U12213 (N_12213,N_11384,N_10631);
nor U12214 (N_12214,N_11018,N_10909);
nor U12215 (N_12215,N_11397,N_10642);
or U12216 (N_12216,N_11986,N_11819);
nand U12217 (N_12217,N_11813,N_10576);
nor U12218 (N_12218,N_10521,N_11458);
xnor U12219 (N_12219,N_10920,N_11367);
or U12220 (N_12220,N_10629,N_11479);
nand U12221 (N_12221,N_11976,N_10667);
nor U12222 (N_12222,N_11910,N_10778);
and U12223 (N_12223,N_10892,N_11118);
or U12224 (N_12224,N_11312,N_11327);
and U12225 (N_12225,N_11721,N_11667);
and U12226 (N_12226,N_10843,N_11561);
or U12227 (N_12227,N_11802,N_11820);
and U12228 (N_12228,N_11503,N_11254);
nand U12229 (N_12229,N_10614,N_11326);
or U12230 (N_12230,N_10818,N_10612);
nand U12231 (N_12231,N_11488,N_11888);
and U12232 (N_12232,N_11422,N_11598);
nand U12233 (N_12233,N_10589,N_11467);
nor U12234 (N_12234,N_11040,N_11698);
or U12235 (N_12235,N_10836,N_11794);
and U12236 (N_12236,N_11786,N_10711);
nor U12237 (N_12237,N_11795,N_11549);
nor U12238 (N_12238,N_11275,N_10999);
or U12239 (N_12239,N_11622,N_11324);
or U12240 (N_12240,N_10870,N_10925);
or U12241 (N_12241,N_11197,N_11350);
nand U12242 (N_12242,N_11586,N_10672);
nor U12243 (N_12243,N_11002,N_10644);
xnor U12244 (N_12244,N_10752,N_11328);
or U12245 (N_12245,N_11900,N_11001);
or U12246 (N_12246,N_11043,N_10532);
nand U12247 (N_12247,N_10841,N_11683);
nor U12248 (N_12248,N_10726,N_11821);
or U12249 (N_12249,N_11266,N_11110);
nand U12250 (N_12250,N_10513,N_11646);
nor U12251 (N_12251,N_11055,N_11400);
and U12252 (N_12252,N_11658,N_10844);
xor U12253 (N_12253,N_11759,N_11968);
nand U12254 (N_12254,N_11812,N_11498);
nand U12255 (N_12255,N_10910,N_11580);
and U12256 (N_12256,N_11262,N_11937);
and U12257 (N_12257,N_10550,N_10756);
and U12258 (N_12258,N_10848,N_11711);
nor U12259 (N_12259,N_11035,N_10798);
nor U12260 (N_12260,N_11388,N_11675);
nand U12261 (N_12261,N_11505,N_11088);
or U12262 (N_12262,N_11568,N_11915);
nor U12263 (N_12263,N_11213,N_11720);
nor U12264 (N_12264,N_11127,N_11161);
and U12265 (N_12265,N_11534,N_11493);
and U12266 (N_12266,N_11962,N_10536);
nand U12267 (N_12267,N_10662,N_11979);
nand U12268 (N_12268,N_11959,N_11902);
or U12269 (N_12269,N_11099,N_11235);
and U12270 (N_12270,N_11927,N_11528);
nor U12271 (N_12271,N_11562,N_11677);
nand U12272 (N_12272,N_10720,N_11189);
and U12273 (N_12273,N_11837,N_11169);
nor U12274 (N_12274,N_10834,N_11094);
nor U12275 (N_12275,N_11183,N_10923);
or U12276 (N_12276,N_11987,N_10854);
and U12277 (N_12277,N_11278,N_11210);
nand U12278 (N_12278,N_10897,N_11446);
and U12279 (N_12279,N_11304,N_11425);
or U12280 (N_12280,N_11299,N_11833);
nand U12281 (N_12281,N_11948,N_10620);
or U12282 (N_12282,N_10524,N_11930);
and U12283 (N_12283,N_11997,N_10847);
or U12284 (N_12284,N_11856,N_10583);
nor U12285 (N_12285,N_10579,N_10827);
nor U12286 (N_12286,N_10737,N_10643);
and U12287 (N_12287,N_10906,N_10901);
or U12288 (N_12288,N_11911,N_11314);
or U12289 (N_12289,N_11988,N_10814);
and U12290 (N_12290,N_11442,N_11412);
xor U12291 (N_12291,N_10828,N_11736);
nor U12292 (N_12292,N_11158,N_10871);
nor U12293 (N_12293,N_10553,N_11177);
or U12294 (N_12294,N_11767,N_10607);
or U12295 (N_12295,N_11717,N_11841);
nand U12296 (N_12296,N_11867,N_11686);
or U12297 (N_12297,N_10557,N_11539);
or U12298 (N_12298,N_10547,N_11552);
and U12299 (N_12299,N_11227,N_10766);
or U12300 (N_12300,N_10903,N_11428);
nand U12301 (N_12301,N_11378,N_11185);
or U12302 (N_12302,N_10964,N_11086);
nand U12303 (N_12303,N_11981,N_10914);
nor U12304 (N_12304,N_10812,N_11045);
nand U12305 (N_12305,N_10915,N_11374);
or U12306 (N_12306,N_11960,N_10930);
and U12307 (N_12307,N_11877,N_11252);
and U12308 (N_12308,N_10863,N_10735);
nand U12309 (N_12309,N_11039,N_10911);
nor U12310 (N_12310,N_11909,N_10533);
nand U12311 (N_12311,N_10976,N_11989);
xor U12312 (N_12312,N_10747,N_10719);
and U12313 (N_12313,N_11782,N_10624);
and U12314 (N_12314,N_11832,N_11468);
nor U12315 (N_12315,N_11141,N_11386);
or U12316 (N_12316,N_10875,N_11396);
and U12317 (N_12317,N_10922,N_11779);
or U12318 (N_12318,N_11365,N_11641);
nor U12319 (N_12319,N_10912,N_11497);
nor U12320 (N_12320,N_11756,N_10635);
nor U12321 (N_12321,N_10683,N_11574);
nor U12322 (N_12322,N_10698,N_11831);
and U12323 (N_12323,N_11558,N_11943);
nor U12324 (N_12324,N_11726,N_10580);
xor U12325 (N_12325,N_11030,N_11074);
and U12326 (N_12326,N_11200,N_10693);
and U12327 (N_12327,N_11515,N_11264);
and U12328 (N_12328,N_10561,N_10613);
xnor U12329 (N_12329,N_10837,N_10833);
or U12330 (N_12330,N_11606,N_10749);
xor U12331 (N_12331,N_10889,N_11525);
nand U12332 (N_12332,N_11393,N_11449);
nor U12333 (N_12333,N_11616,N_11570);
nand U12334 (N_12334,N_10677,N_11647);
and U12335 (N_12335,N_11548,N_10793);
nand U12336 (N_12336,N_10786,N_11460);
nand U12337 (N_12337,N_10965,N_10840);
nor U12338 (N_12338,N_10539,N_11492);
or U12339 (N_12339,N_11718,N_11532);
or U12340 (N_12340,N_11995,N_10594);
nand U12341 (N_12341,N_10664,N_10885);
nand U12342 (N_12342,N_10573,N_10556);
or U12343 (N_12343,N_11358,N_11306);
or U12344 (N_12344,N_11364,N_10988);
or U12345 (N_12345,N_11547,N_11072);
nand U12346 (N_12346,N_10765,N_11073);
or U12347 (N_12347,N_11237,N_11216);
nand U12348 (N_12348,N_10604,N_10694);
or U12349 (N_12349,N_10794,N_11682);
or U12350 (N_12350,N_11868,N_11908);
or U12351 (N_12351,N_11920,N_11164);
nor U12352 (N_12352,N_11521,N_11971);
nor U12353 (N_12353,N_11067,N_10972);
nand U12354 (N_12354,N_10619,N_11052);
or U12355 (N_12355,N_11368,N_11201);
nor U12356 (N_12356,N_11916,N_11149);
and U12357 (N_12357,N_10590,N_11355);
and U12358 (N_12358,N_11905,N_11593);
nor U12359 (N_12359,N_11000,N_11828);
nor U12360 (N_12360,N_11588,N_11406);
and U12361 (N_12361,N_11737,N_11027);
or U12362 (N_12362,N_11120,N_11332);
and U12363 (N_12363,N_10653,N_10878);
or U12364 (N_12364,N_11105,N_10656);
nand U12365 (N_12365,N_11003,N_10679);
or U12366 (N_12366,N_11777,N_11315);
or U12367 (N_12367,N_10652,N_10704);
nand U12368 (N_12368,N_10678,N_11518);
nor U12369 (N_12369,N_10593,N_11674);
nor U12370 (N_12370,N_11084,N_10884);
nor U12371 (N_12371,N_10548,N_11409);
nand U12372 (N_12372,N_11032,N_10616);
nor U12373 (N_12373,N_10651,N_11060);
and U12374 (N_12374,N_11281,N_11731);
nor U12375 (N_12375,N_11334,N_11514);
or U12376 (N_12376,N_10645,N_11466);
or U12377 (N_12377,N_11583,N_10853);
nor U12378 (N_12378,N_10660,N_11851);
nor U12379 (N_12379,N_10606,N_10563);
or U12380 (N_12380,N_11854,N_11784);
or U12381 (N_12381,N_10597,N_11033);
or U12382 (N_12382,N_11662,N_11862);
xor U12383 (N_12383,N_11391,N_10566);
nand U12384 (N_12384,N_10928,N_10582);
or U12385 (N_12385,N_11291,N_11857);
or U12386 (N_12386,N_11781,N_11860);
nor U12387 (N_12387,N_11896,N_11842);
or U12388 (N_12388,N_10890,N_10688);
nor U12389 (N_12389,N_10714,N_10974);
nand U12390 (N_12390,N_10601,N_11839);
or U12391 (N_12391,N_11174,N_11638);
and U12392 (N_12392,N_11838,N_11690);
or U12393 (N_12393,N_11005,N_11476);
and U12394 (N_12394,N_11217,N_11808);
or U12395 (N_12395,N_11984,N_11657);
and U12396 (N_12396,N_11906,N_10731);
or U12397 (N_12397,N_11037,N_10706);
nand U12398 (N_12398,N_11116,N_11302);
or U12399 (N_12399,N_11591,N_11835);
xnor U12400 (N_12400,N_11645,N_11614);
and U12401 (N_12401,N_11050,N_11557);
nor U12402 (N_12402,N_11337,N_11323);
nand U12403 (N_12403,N_10861,N_11714);
or U12404 (N_12404,N_11163,N_11404);
and U12405 (N_12405,N_11993,N_11008);
or U12406 (N_12406,N_11325,N_11766);
and U12407 (N_12407,N_10755,N_11879);
and U12408 (N_12408,N_11730,N_11527);
nand U12409 (N_12409,N_11471,N_10761);
or U12410 (N_12410,N_11417,N_11321);
nor U12411 (N_12411,N_11704,N_11240);
nor U12412 (N_12412,N_11931,N_10609);
and U12413 (N_12413,N_11424,N_10953);
nand U12414 (N_12414,N_11967,N_11592);
and U12415 (N_12415,N_11956,N_11554);
or U12416 (N_12416,N_11797,N_11081);
nand U12417 (N_12417,N_11504,N_11950);
and U12418 (N_12418,N_11418,N_11434);
nor U12419 (N_12419,N_11630,N_10908);
nand U12420 (N_12420,N_11108,N_10941);
nor U12421 (N_12421,N_11707,N_10796);
nor U12422 (N_12422,N_10877,N_10743);
or U12423 (N_12423,N_10636,N_10831);
nand U12424 (N_12424,N_11893,N_11444);
or U12425 (N_12425,N_11140,N_11155);
or U12426 (N_12426,N_11265,N_11590);
nand U12427 (N_12427,N_11193,N_11754);
or U12428 (N_12428,N_11871,N_11772);
and U12429 (N_12429,N_11046,N_11807);
or U12430 (N_12430,N_10845,N_11168);
nand U12431 (N_12431,N_11665,N_10994);
nand U12432 (N_12432,N_10858,N_10730);
xor U12433 (N_12433,N_11283,N_11112);
nand U12434 (N_12434,N_11206,N_10830);
nand U12435 (N_12435,N_10763,N_10671);
and U12436 (N_12436,N_11233,N_11165);
or U12437 (N_12437,N_10961,N_10546);
nor U12438 (N_12438,N_10983,N_10938);
and U12439 (N_12439,N_11075,N_11336);
or U12440 (N_12440,N_11380,N_10968);
nand U12441 (N_12441,N_10967,N_11537);
nand U12442 (N_12442,N_11619,N_11104);
and U12443 (N_12443,N_11830,N_11952);
or U12444 (N_12444,N_10797,N_11510);
nand U12445 (N_12445,N_10715,N_10658);
nand U12446 (N_12446,N_11615,N_11371);
or U12447 (N_12447,N_11722,N_11914);
nor U12448 (N_12448,N_10739,N_10647);
nand U12449 (N_12449,N_11618,N_10868);
nor U12450 (N_12450,N_11117,N_11241);
and U12451 (N_12451,N_11419,N_11749);
and U12452 (N_12452,N_11119,N_11546);
and U12453 (N_12453,N_11520,N_10687);
and U12454 (N_12454,N_10520,N_11847);
and U12455 (N_12455,N_11512,N_11581);
and U12456 (N_12456,N_11589,N_11136);
nand U12457 (N_12457,N_11949,N_10713);
and U12458 (N_12458,N_11508,N_11680);
nand U12459 (N_12459,N_11980,N_10824);
or U12460 (N_12460,N_11041,N_10526);
or U12461 (N_12461,N_10741,N_11430);
or U12462 (N_12462,N_10661,N_11415);
nand U12463 (N_12463,N_11082,N_10570);
nand U12464 (N_12464,N_10617,N_10516);
nand U12465 (N_12465,N_11524,N_11459);
and U12466 (N_12466,N_11921,N_11744);
and U12467 (N_12467,N_10538,N_11253);
and U12468 (N_12468,N_11125,N_11068);
or U12469 (N_12469,N_11990,N_11864);
nand U12470 (N_12470,N_10541,N_11250);
or U12471 (N_12471,N_10916,N_10917);
or U12472 (N_12472,N_11824,N_10676);
or U12473 (N_12473,N_11870,N_10542);
and U12474 (N_12474,N_11453,N_11925);
and U12475 (N_12475,N_11440,N_11036);
or U12476 (N_12476,N_11249,N_11401);
or U12477 (N_12477,N_11845,N_11284);
nand U12478 (N_12478,N_10769,N_10985);
or U12479 (N_12479,N_11133,N_10867);
nor U12480 (N_12480,N_10627,N_10900);
nand U12481 (N_12481,N_10913,N_11416);
nand U12482 (N_12482,N_10780,N_11747);
or U12483 (N_12483,N_11114,N_11699);
or U12484 (N_12484,N_10696,N_10779);
nand U12485 (N_12485,N_11903,N_11817);
nand U12486 (N_12486,N_11379,N_10939);
xor U12487 (N_12487,N_11004,N_11429);
and U12488 (N_12488,N_11563,N_10692);
nand U12489 (N_12489,N_11669,N_11874);
or U12490 (N_12490,N_11958,N_10782);
nand U12491 (N_12491,N_10937,N_11681);
nor U12492 (N_12492,N_11639,N_10895);
nand U12493 (N_12493,N_10825,N_11922);
xnor U12494 (N_12494,N_11928,N_11285);
nand U12495 (N_12495,N_11229,N_11280);
and U12496 (N_12496,N_11289,N_11457);
and U12497 (N_12497,N_10646,N_11221);
or U12498 (N_12498,N_11473,N_11061);
or U12499 (N_12499,N_11272,N_11975);
and U12500 (N_12500,N_11540,N_11530);
xnor U12501 (N_12501,N_10623,N_11869);
or U12502 (N_12502,N_11678,N_10838);
and U12503 (N_12503,N_11062,N_11723);
and U12504 (N_12504,N_11827,N_11770);
nand U12505 (N_12505,N_11785,N_11923);
nor U12506 (N_12506,N_11007,N_11708);
xor U12507 (N_12507,N_11196,N_11172);
nand U12508 (N_12508,N_10554,N_10835);
nor U12509 (N_12509,N_11938,N_10507);
nor U12510 (N_12510,N_11056,N_11408);
nor U12511 (N_12511,N_11829,N_11944);
xnor U12512 (N_12512,N_11628,N_11666);
and U12513 (N_12513,N_11438,N_11732);
nor U12514 (N_12514,N_11626,N_11013);
nand U12515 (N_12515,N_10902,N_11423);
or U12516 (N_12516,N_11220,N_11454);
nand U12517 (N_12517,N_10639,N_11790);
and U12518 (N_12518,N_11796,N_11451);
or U12519 (N_12519,N_11725,N_10691);
and U12520 (N_12520,N_10958,N_10822);
or U12521 (N_12521,N_11752,N_10852);
or U12522 (N_12522,N_10980,N_11758);
and U12523 (N_12523,N_11106,N_11481);
and U12524 (N_12524,N_11202,N_11109);
nor U12525 (N_12525,N_11881,N_11664);
and U12526 (N_12526,N_11057,N_10933);
nor U12527 (N_12527,N_11478,N_10600);
nor U12528 (N_12528,N_11565,N_11162);
xnor U12529 (N_12529,N_11222,N_11394);
xnor U12530 (N_12530,N_11765,N_11750);
or U12531 (N_12531,N_11499,N_11093);
nor U12532 (N_12532,N_11376,N_10882);
or U12533 (N_12533,N_11643,N_10879);
or U12534 (N_12534,N_10522,N_11316);
and U12535 (N_12535,N_11768,N_11122);
or U12536 (N_12536,N_10924,N_11809);
nor U12537 (N_12537,N_11407,N_11107);
nor U12538 (N_12538,N_11691,N_11091);
nor U12539 (N_12539,N_10750,N_10866);
or U12540 (N_12540,N_10709,N_11224);
xnor U12541 (N_12541,N_11746,N_10705);
nor U12542 (N_12542,N_11028,N_11482);
and U12543 (N_12543,N_11523,N_11753);
or U12544 (N_12544,N_11858,N_11148);
nand U12545 (N_12545,N_11825,N_11319);
nor U12546 (N_12546,N_10621,N_11421);
and U12547 (N_12547,N_10791,N_10929);
nor U12548 (N_12548,N_11652,N_10585);
nand U12549 (N_12549,N_11166,N_10537);
nor U12550 (N_12550,N_11223,N_11936);
nor U12551 (N_12551,N_10700,N_11318);
and U12552 (N_12552,N_10584,N_10790);
nor U12553 (N_12553,N_11300,N_10907);
and U12554 (N_12554,N_10708,N_10784);
nand U12555 (N_12555,N_10751,N_11875);
nand U12556 (N_12556,N_11199,N_11571);
and U12557 (N_12557,N_10860,N_10592);
or U12558 (N_12558,N_11248,N_11167);
nor U12559 (N_12559,N_11245,N_10515);
nand U12560 (N_12560,N_11904,N_11740);
nor U12561 (N_12561,N_11716,N_11359);
nand U12562 (N_12562,N_11042,N_11560);
or U12563 (N_12563,N_11184,N_10502);
or U12564 (N_12564,N_10760,N_10558);
nand U12565 (N_12565,N_10998,N_11640);
nand U12566 (N_12566,N_11757,N_11955);
and U12567 (N_12567,N_10510,N_10567);
or U12568 (N_12568,N_10886,N_11349);
and U12569 (N_12569,N_11157,N_11357);
or U12570 (N_12570,N_11954,N_11852);
nor U12571 (N_12571,N_11242,N_11077);
nor U12572 (N_12572,N_10734,N_10894);
and U12573 (N_12573,N_10528,N_11584);
nand U12574 (N_12574,N_11631,N_11535);
or U12575 (N_12575,N_11884,N_10942);
nor U12576 (N_12576,N_10648,N_11506);
nor U12577 (N_12577,N_10960,N_11238);
nor U12578 (N_12578,N_11441,N_11362);
nor U12579 (N_12579,N_11188,N_10525);
or U12580 (N_12580,N_11576,N_11331);
and U12581 (N_12581,N_11803,N_11776);
nor U12582 (N_12582,N_11019,N_10850);
nor U12583 (N_12583,N_10728,N_11246);
or U12584 (N_12584,N_11179,N_11693);
or U12585 (N_12585,N_11012,N_11178);
or U12586 (N_12586,N_11034,N_11290);
nor U12587 (N_12587,N_11578,N_10571);
or U12588 (N_12588,N_11026,N_11352);
nand U12589 (N_12589,N_11098,N_10783);
nor U12590 (N_12590,N_11917,N_11296);
nand U12591 (N_12591,N_11100,N_11420);
nor U12592 (N_12592,N_11684,N_11171);
nand U12593 (N_12593,N_10500,N_11146);
and U12594 (N_12594,N_10625,N_11131);
or U12595 (N_12595,N_11486,N_10826);
nor U12596 (N_12596,N_11994,N_11192);
and U12597 (N_12597,N_11377,N_11579);
nor U12598 (N_12598,N_11775,N_11134);
nor U12599 (N_12599,N_11273,N_11239);
and U12600 (N_12600,N_11880,N_10883);
or U12601 (N_12601,N_11597,N_11340);
nand U12602 (N_12602,N_11194,N_10549);
xnor U12603 (N_12603,N_10733,N_11659);
or U12604 (N_12604,N_10686,N_11135);
and U12605 (N_12605,N_10898,N_11850);
and U12606 (N_12606,N_11769,N_11139);
nand U12607 (N_12607,N_11137,N_11372);
nand U12608 (N_12608,N_11207,N_11983);
or U12609 (N_12609,N_11509,N_11244);
or U12610 (N_12610,N_11733,N_11403);
nor U12611 (N_12611,N_11341,N_11610);
and U12612 (N_12612,N_11855,N_10523);
nor U12613 (N_12613,N_10602,N_11999);
or U12614 (N_12614,N_10724,N_10773);
and U12615 (N_12615,N_11494,N_11513);
and U12616 (N_12616,N_10978,N_10675);
and U12617 (N_12617,N_10946,N_11969);
or U12618 (N_12618,N_11215,N_11951);
nand U12619 (N_12619,N_11138,N_10893);
and U12620 (N_12620,N_11745,N_11496);
and U12621 (N_12621,N_11342,N_10703);
nand U12622 (N_12622,N_10806,N_10865);
nor U12623 (N_12623,N_10851,N_11810);
nor U12624 (N_12624,N_11788,N_11150);
and U12625 (N_12625,N_10849,N_11154);
nand U12626 (N_12626,N_10888,N_11375);
or U12627 (N_12627,N_11101,N_11477);
xor U12628 (N_12628,N_10969,N_10655);
and U12629 (N_12629,N_10572,N_11023);
or U12630 (N_12630,N_11047,N_11617);
nor U12631 (N_12631,N_11926,N_10821);
and U12632 (N_12632,N_11982,N_11648);
nor U12633 (N_12633,N_10934,N_11330);
nor U12634 (N_12634,N_11729,N_10799);
nor U12635 (N_12635,N_11190,N_11519);
nand U12636 (N_12636,N_11366,N_11977);
nand U12637 (N_12637,N_10555,N_10673);
nand U12638 (N_12638,N_11069,N_11462);
nor U12639 (N_12639,N_10951,N_11092);
nand U12640 (N_12640,N_11544,N_10947);
nand U12641 (N_12641,N_11792,N_11791);
or U12642 (N_12642,N_11282,N_10919);
or U12643 (N_12643,N_11654,N_11650);
nand U12644 (N_12644,N_11232,N_11294);
or U12645 (N_12645,N_11526,N_11076);
nand U12646 (N_12646,N_11734,N_11006);
nand U12647 (N_12647,N_11044,N_11475);
nand U12648 (N_12648,N_11706,N_10615);
or U12649 (N_12649,N_11480,N_11258);
or U12650 (N_12650,N_10921,N_10736);
or U12651 (N_12651,N_10989,N_11778);
and U12652 (N_12652,N_11021,N_11621);
or U12653 (N_12653,N_11804,N_11383);
nand U12654 (N_12654,N_10587,N_10795);
and U12655 (N_12655,N_10575,N_11413);
nor U12656 (N_12656,N_11551,N_11058);
nor U12657 (N_12657,N_10503,N_10918);
and U12658 (N_12658,N_11885,N_11445);
or U12659 (N_12659,N_11095,N_10862);
nand U12660 (N_12660,N_11946,N_11661);
nor U12661 (N_12661,N_10931,N_11435);
or U12662 (N_12662,N_11972,N_10927);
nor U12663 (N_12663,N_11191,N_11469);
and U12664 (N_12664,N_10722,N_11353);
nand U12665 (N_12665,N_10543,N_10975);
nor U12666 (N_12666,N_10505,N_11872);
nand U12667 (N_12667,N_11761,N_11771);
or U12668 (N_12668,N_11322,N_10758);
and U12669 (N_12669,N_11410,N_11211);
nor U12670 (N_12670,N_10702,N_11307);
nand U12671 (N_12671,N_11345,N_11596);
and U12672 (N_12672,N_11603,N_11356);
nand U12673 (N_12673,N_11431,N_11542);
and U12674 (N_12674,N_11865,N_11811);
or U12675 (N_12675,N_11705,N_11755);
and U12676 (N_12676,N_11555,N_10815);
nor U12677 (N_12677,N_10586,N_11671);
xor U12678 (N_12678,N_11022,N_11490);
or U12679 (N_12679,N_10872,N_11531);
or U12680 (N_12680,N_11940,N_11173);
nand U12681 (N_12681,N_11226,N_11836);
nand U12682 (N_12682,N_11295,N_11748);
nand U12683 (N_12683,N_11333,N_10987);
nor U12684 (N_12684,N_11973,N_11276);
nor U12685 (N_12685,N_11259,N_11741);
and U12686 (N_12686,N_11343,N_11234);
nand U12687 (N_12687,N_11320,N_11712);
or U12688 (N_12688,N_11472,N_10771);
or U12689 (N_12689,N_10839,N_11270);
or U12690 (N_12690,N_11288,N_11728);
nor U12691 (N_12691,N_10997,N_11151);
or U12692 (N_12692,N_11071,N_11236);
or U12693 (N_12693,N_11876,N_11017);
nor U12694 (N_12694,N_10785,N_11344);
and U12695 (N_12695,N_11806,N_11212);
nor U12696 (N_12696,N_11609,N_10674);
nand U12697 (N_12697,N_10984,N_11485);
nand U12698 (N_12698,N_11426,N_11688);
xnor U12699 (N_12699,N_10776,N_10788);
or U12700 (N_12700,N_10781,N_11447);
or U12701 (N_12701,N_10932,N_11543);
nand U12702 (N_12702,N_11516,N_11051);
and U12703 (N_12703,N_11303,N_11461);
nand U12704 (N_12704,N_10986,N_11031);
or U12705 (N_12705,N_11673,N_11694);
or U12706 (N_12706,N_11941,N_10740);
or U12707 (N_12707,N_11361,N_11801);
or U12708 (N_12708,N_11147,N_10887);
or U12709 (N_12709,N_11464,N_11381);
and U12710 (N_12710,N_11637,N_11724);
and U12711 (N_12711,N_10802,N_10956);
nor U12712 (N_12712,N_10506,N_10952);
nand U12713 (N_12713,N_11599,N_11966);
nand U12714 (N_12714,N_10803,N_11918);
nand U12715 (N_12715,N_11293,N_10787);
or U12716 (N_12716,N_11153,N_10529);
nand U12717 (N_12717,N_11859,N_11991);
nand U12718 (N_12718,N_10717,N_11739);
and U12719 (N_12719,N_11038,N_11351);
and U12720 (N_12720,N_11517,N_11934);
nor U12721 (N_12721,N_11129,N_10767);
and U12722 (N_12722,N_11582,N_11228);
or U12723 (N_12723,N_11247,N_11963);
or U12724 (N_12724,N_11354,N_11566);
nand U12725 (N_12725,N_11932,N_10531);
and U12726 (N_12726,N_11389,N_11267);
nand U12727 (N_12727,N_10689,N_10577);
nor U12728 (N_12728,N_10811,N_10970);
or U12729 (N_12729,N_10959,N_11465);
or U12730 (N_12730,N_11208,N_11763);
or U12731 (N_12731,N_11263,N_10611);
and U12732 (N_12732,N_11078,N_11511);
nand U12733 (N_12733,N_11268,N_10770);
nand U12734 (N_12734,N_11635,N_11339);
or U12735 (N_12735,N_11522,N_11861);
nand U12736 (N_12736,N_10991,N_11255);
and U12737 (N_12737,N_10996,N_11559);
and U12738 (N_12738,N_11079,N_10846);
or U12739 (N_12739,N_10638,N_10530);
nor U12740 (N_12740,N_10669,N_10595);
nor U12741 (N_12741,N_11891,N_11538);
nand U12742 (N_12742,N_11382,N_11205);
nand U12743 (N_12743,N_11608,N_10864);
or U12744 (N_12744,N_10544,N_11703);
nor U12745 (N_12745,N_11742,N_11826);
or U12746 (N_12746,N_11335,N_10856);
and U12747 (N_12747,N_10874,N_11347);
nor U12748 (N_12748,N_10807,N_11070);
nor U12749 (N_12749,N_11015,N_10800);
nor U12750 (N_12750,N_10680,N_11517);
nand U12751 (N_12751,N_10954,N_10778);
nand U12752 (N_12752,N_10598,N_11311);
nand U12753 (N_12753,N_11201,N_10919);
and U12754 (N_12754,N_10849,N_11920);
nand U12755 (N_12755,N_11263,N_11256);
nor U12756 (N_12756,N_11581,N_10551);
nand U12757 (N_12757,N_11948,N_10757);
nor U12758 (N_12758,N_11958,N_10628);
or U12759 (N_12759,N_11752,N_11851);
nor U12760 (N_12760,N_10580,N_11182);
nor U12761 (N_12761,N_11498,N_11288);
xnor U12762 (N_12762,N_11418,N_10692);
nand U12763 (N_12763,N_11208,N_11186);
or U12764 (N_12764,N_11501,N_11890);
xnor U12765 (N_12765,N_11174,N_10529);
nand U12766 (N_12766,N_10856,N_10945);
or U12767 (N_12767,N_11858,N_11089);
nand U12768 (N_12768,N_11815,N_10905);
nor U12769 (N_12769,N_11555,N_11577);
nand U12770 (N_12770,N_10581,N_11319);
nor U12771 (N_12771,N_11725,N_11764);
and U12772 (N_12772,N_11337,N_10616);
or U12773 (N_12773,N_11630,N_11840);
and U12774 (N_12774,N_11938,N_11175);
or U12775 (N_12775,N_11110,N_11877);
and U12776 (N_12776,N_11253,N_10974);
nor U12777 (N_12777,N_10826,N_10622);
nand U12778 (N_12778,N_11159,N_10801);
nand U12779 (N_12779,N_11990,N_10679);
nand U12780 (N_12780,N_10856,N_11124);
or U12781 (N_12781,N_11427,N_10952);
and U12782 (N_12782,N_11310,N_10843);
nor U12783 (N_12783,N_10671,N_11684);
nor U12784 (N_12784,N_11105,N_10867);
and U12785 (N_12785,N_11540,N_11252);
or U12786 (N_12786,N_10928,N_11069);
nand U12787 (N_12787,N_11673,N_11597);
and U12788 (N_12788,N_11091,N_11410);
nand U12789 (N_12789,N_11673,N_11064);
nand U12790 (N_12790,N_10688,N_10976);
nor U12791 (N_12791,N_11198,N_11554);
or U12792 (N_12792,N_10920,N_11346);
nand U12793 (N_12793,N_11899,N_11861);
nor U12794 (N_12794,N_10537,N_11226);
nor U12795 (N_12795,N_11210,N_11923);
nand U12796 (N_12796,N_11161,N_11381);
or U12797 (N_12797,N_10548,N_10666);
and U12798 (N_12798,N_11324,N_11437);
nand U12799 (N_12799,N_10841,N_11750);
or U12800 (N_12800,N_11288,N_11870);
nor U12801 (N_12801,N_11982,N_11006);
and U12802 (N_12802,N_11908,N_11172);
nor U12803 (N_12803,N_11050,N_11033);
nor U12804 (N_12804,N_10709,N_11558);
or U12805 (N_12805,N_10602,N_11718);
nor U12806 (N_12806,N_11420,N_11673);
nand U12807 (N_12807,N_10643,N_11197);
nor U12808 (N_12808,N_11866,N_10579);
or U12809 (N_12809,N_11828,N_10715);
nand U12810 (N_12810,N_11394,N_11271);
or U12811 (N_12811,N_11414,N_10953);
and U12812 (N_12812,N_10732,N_10832);
or U12813 (N_12813,N_11579,N_10750);
and U12814 (N_12814,N_10922,N_11200);
and U12815 (N_12815,N_11760,N_11621);
and U12816 (N_12816,N_11224,N_11534);
and U12817 (N_12817,N_11674,N_11182);
and U12818 (N_12818,N_10631,N_11067);
or U12819 (N_12819,N_10560,N_11114);
and U12820 (N_12820,N_11348,N_11628);
nor U12821 (N_12821,N_11096,N_11860);
and U12822 (N_12822,N_11969,N_10753);
and U12823 (N_12823,N_10925,N_11566);
or U12824 (N_12824,N_11921,N_11478);
and U12825 (N_12825,N_11074,N_10843);
nor U12826 (N_12826,N_10938,N_10713);
nand U12827 (N_12827,N_11788,N_11720);
nand U12828 (N_12828,N_11691,N_11713);
xnor U12829 (N_12829,N_11083,N_10836);
nand U12830 (N_12830,N_11012,N_11997);
nor U12831 (N_12831,N_10904,N_10620);
nor U12832 (N_12832,N_11195,N_10940);
nand U12833 (N_12833,N_11588,N_11105);
nor U12834 (N_12834,N_11574,N_11364);
nand U12835 (N_12835,N_11746,N_10775);
nand U12836 (N_12836,N_11032,N_11380);
or U12837 (N_12837,N_11608,N_11316);
or U12838 (N_12838,N_10520,N_11874);
nor U12839 (N_12839,N_11417,N_11693);
or U12840 (N_12840,N_11343,N_10729);
nor U12841 (N_12841,N_11144,N_11813);
or U12842 (N_12842,N_10509,N_10544);
xnor U12843 (N_12843,N_11038,N_11171);
nand U12844 (N_12844,N_11913,N_11040);
nor U12845 (N_12845,N_10841,N_11546);
xnor U12846 (N_12846,N_11426,N_10855);
nor U12847 (N_12847,N_10795,N_11868);
or U12848 (N_12848,N_11716,N_11969);
or U12849 (N_12849,N_11707,N_11677);
or U12850 (N_12850,N_10976,N_11787);
or U12851 (N_12851,N_11835,N_11608);
nand U12852 (N_12852,N_11049,N_11869);
and U12853 (N_12853,N_11453,N_10609);
or U12854 (N_12854,N_11922,N_10961);
nand U12855 (N_12855,N_11460,N_10881);
or U12856 (N_12856,N_11781,N_11180);
nand U12857 (N_12857,N_10573,N_11324);
and U12858 (N_12858,N_11633,N_10632);
nand U12859 (N_12859,N_11270,N_11354);
or U12860 (N_12860,N_11946,N_11410);
nand U12861 (N_12861,N_10834,N_10760);
nand U12862 (N_12862,N_10866,N_10922);
and U12863 (N_12863,N_11814,N_11238);
and U12864 (N_12864,N_11354,N_11272);
nand U12865 (N_12865,N_10553,N_11022);
and U12866 (N_12866,N_11007,N_11181);
and U12867 (N_12867,N_11333,N_10514);
or U12868 (N_12868,N_10531,N_10953);
nand U12869 (N_12869,N_10956,N_10657);
or U12870 (N_12870,N_11958,N_10653);
or U12871 (N_12871,N_10990,N_11766);
or U12872 (N_12872,N_11183,N_11037);
nor U12873 (N_12873,N_10522,N_11896);
or U12874 (N_12874,N_11172,N_11243);
nor U12875 (N_12875,N_11157,N_11052);
or U12876 (N_12876,N_11635,N_11931);
or U12877 (N_12877,N_11559,N_10668);
nand U12878 (N_12878,N_10763,N_11908);
nand U12879 (N_12879,N_11748,N_11081);
and U12880 (N_12880,N_11122,N_11700);
or U12881 (N_12881,N_10841,N_11575);
nand U12882 (N_12882,N_10733,N_10825);
nor U12883 (N_12883,N_11204,N_10986);
nor U12884 (N_12884,N_11734,N_11594);
nand U12885 (N_12885,N_11848,N_10865);
nand U12886 (N_12886,N_11029,N_11575);
and U12887 (N_12887,N_10704,N_10543);
or U12888 (N_12888,N_11775,N_11143);
nor U12889 (N_12889,N_11350,N_11503);
nor U12890 (N_12890,N_10693,N_10839);
and U12891 (N_12891,N_11751,N_11199);
nand U12892 (N_12892,N_10669,N_11292);
and U12893 (N_12893,N_11355,N_11149);
nand U12894 (N_12894,N_11431,N_10536);
and U12895 (N_12895,N_11595,N_11377);
nor U12896 (N_12896,N_11777,N_11788);
and U12897 (N_12897,N_11624,N_11157);
and U12898 (N_12898,N_10895,N_11375);
or U12899 (N_12899,N_10735,N_10630);
nor U12900 (N_12900,N_11515,N_10508);
nor U12901 (N_12901,N_11147,N_11014);
or U12902 (N_12902,N_11090,N_10704);
nand U12903 (N_12903,N_10749,N_11605);
and U12904 (N_12904,N_11398,N_10726);
or U12905 (N_12905,N_11557,N_11122);
or U12906 (N_12906,N_10939,N_10845);
or U12907 (N_12907,N_11802,N_11793);
or U12908 (N_12908,N_11651,N_11001);
or U12909 (N_12909,N_10962,N_10681);
nor U12910 (N_12910,N_11470,N_10793);
nand U12911 (N_12911,N_11513,N_11372);
nand U12912 (N_12912,N_11751,N_11992);
or U12913 (N_12913,N_11259,N_11677);
or U12914 (N_12914,N_11650,N_11935);
nand U12915 (N_12915,N_10566,N_11884);
or U12916 (N_12916,N_11439,N_11592);
nor U12917 (N_12917,N_10993,N_10617);
or U12918 (N_12918,N_10749,N_11417);
and U12919 (N_12919,N_10699,N_10637);
and U12920 (N_12920,N_10861,N_11868);
nor U12921 (N_12921,N_10900,N_11903);
and U12922 (N_12922,N_11467,N_11804);
and U12923 (N_12923,N_11677,N_10957);
or U12924 (N_12924,N_10902,N_10879);
or U12925 (N_12925,N_10932,N_10841);
or U12926 (N_12926,N_10706,N_11126);
nor U12927 (N_12927,N_11140,N_10977);
nor U12928 (N_12928,N_11955,N_11133);
or U12929 (N_12929,N_11368,N_11067);
and U12930 (N_12930,N_11373,N_11020);
nand U12931 (N_12931,N_11112,N_11818);
or U12932 (N_12932,N_11767,N_11253);
and U12933 (N_12933,N_11861,N_11260);
and U12934 (N_12934,N_11440,N_11911);
nand U12935 (N_12935,N_11922,N_11729);
and U12936 (N_12936,N_11941,N_10852);
nor U12937 (N_12937,N_11842,N_10838);
nor U12938 (N_12938,N_11519,N_10906);
and U12939 (N_12939,N_11852,N_10661);
nor U12940 (N_12940,N_10879,N_10949);
nor U12941 (N_12941,N_11571,N_11939);
or U12942 (N_12942,N_11031,N_10599);
nand U12943 (N_12943,N_11699,N_10504);
nor U12944 (N_12944,N_10974,N_11821);
or U12945 (N_12945,N_11194,N_10519);
and U12946 (N_12946,N_11855,N_11528);
and U12947 (N_12947,N_11545,N_11621);
or U12948 (N_12948,N_10952,N_10645);
or U12949 (N_12949,N_10655,N_11502);
nand U12950 (N_12950,N_10898,N_11505);
nor U12951 (N_12951,N_10587,N_10605);
nor U12952 (N_12952,N_11442,N_11699);
nand U12953 (N_12953,N_11964,N_11590);
or U12954 (N_12954,N_11732,N_11919);
xor U12955 (N_12955,N_11982,N_10813);
or U12956 (N_12956,N_10886,N_11633);
and U12957 (N_12957,N_10779,N_11012);
nand U12958 (N_12958,N_10552,N_11452);
nand U12959 (N_12959,N_10733,N_11903);
nor U12960 (N_12960,N_10781,N_10879);
nand U12961 (N_12961,N_11154,N_11938);
and U12962 (N_12962,N_11821,N_11742);
or U12963 (N_12963,N_11388,N_11015);
and U12964 (N_12964,N_11770,N_10787);
and U12965 (N_12965,N_11016,N_10674);
nand U12966 (N_12966,N_11285,N_10515);
and U12967 (N_12967,N_11766,N_11923);
and U12968 (N_12968,N_11295,N_11435);
or U12969 (N_12969,N_10808,N_10793);
nor U12970 (N_12970,N_11846,N_11808);
nor U12971 (N_12971,N_11415,N_11381);
and U12972 (N_12972,N_11335,N_11558);
or U12973 (N_12973,N_10513,N_11197);
nor U12974 (N_12974,N_11390,N_10677);
xnor U12975 (N_12975,N_11682,N_11156);
nor U12976 (N_12976,N_10517,N_10812);
or U12977 (N_12977,N_10986,N_11097);
and U12978 (N_12978,N_11096,N_11782);
or U12979 (N_12979,N_10601,N_11331);
or U12980 (N_12980,N_11056,N_11915);
nand U12981 (N_12981,N_11712,N_11541);
and U12982 (N_12982,N_11643,N_11197);
nand U12983 (N_12983,N_11571,N_11445);
nor U12984 (N_12984,N_10636,N_11067);
xnor U12985 (N_12985,N_10704,N_10598);
or U12986 (N_12986,N_11105,N_11002);
and U12987 (N_12987,N_11396,N_11401);
and U12988 (N_12988,N_11893,N_11583);
or U12989 (N_12989,N_10765,N_10571);
or U12990 (N_12990,N_11045,N_11595);
nor U12991 (N_12991,N_11282,N_11254);
nor U12992 (N_12992,N_11835,N_10656);
nor U12993 (N_12993,N_10749,N_10906);
and U12994 (N_12994,N_11609,N_11139);
nand U12995 (N_12995,N_10789,N_11814);
and U12996 (N_12996,N_10689,N_10696);
nor U12997 (N_12997,N_11398,N_10878);
and U12998 (N_12998,N_11753,N_11855);
and U12999 (N_12999,N_11763,N_11097);
nand U13000 (N_13000,N_10549,N_11510);
and U13001 (N_13001,N_11072,N_11945);
and U13002 (N_13002,N_11509,N_10809);
nand U13003 (N_13003,N_10695,N_10772);
and U13004 (N_13004,N_11578,N_11579);
nor U13005 (N_13005,N_11328,N_10605);
nand U13006 (N_13006,N_10887,N_10803);
and U13007 (N_13007,N_10631,N_11997);
nor U13008 (N_13008,N_11390,N_11492);
nand U13009 (N_13009,N_11730,N_11697);
and U13010 (N_13010,N_10949,N_11297);
or U13011 (N_13011,N_11601,N_11796);
and U13012 (N_13012,N_11962,N_11114);
nand U13013 (N_13013,N_11342,N_11903);
nand U13014 (N_13014,N_10902,N_11560);
nor U13015 (N_13015,N_11246,N_11089);
nor U13016 (N_13016,N_10642,N_11159);
nor U13017 (N_13017,N_10859,N_11446);
nand U13018 (N_13018,N_11429,N_10983);
nor U13019 (N_13019,N_11789,N_11662);
nand U13020 (N_13020,N_11564,N_11440);
nand U13021 (N_13021,N_11006,N_10727);
nand U13022 (N_13022,N_11679,N_11983);
nand U13023 (N_13023,N_11943,N_11901);
xnor U13024 (N_13024,N_11381,N_10678);
and U13025 (N_13025,N_11850,N_10866);
and U13026 (N_13026,N_10738,N_11061);
nor U13027 (N_13027,N_11390,N_10560);
or U13028 (N_13028,N_11534,N_11307);
nor U13029 (N_13029,N_11864,N_11238);
and U13030 (N_13030,N_11033,N_11047);
nand U13031 (N_13031,N_11931,N_11076);
and U13032 (N_13032,N_10778,N_11308);
or U13033 (N_13033,N_10615,N_11455);
and U13034 (N_13034,N_11471,N_10905);
xnor U13035 (N_13035,N_10628,N_11526);
nor U13036 (N_13036,N_11214,N_11316);
nand U13037 (N_13037,N_11852,N_11692);
or U13038 (N_13038,N_11419,N_11759);
nor U13039 (N_13039,N_10578,N_10737);
or U13040 (N_13040,N_10963,N_11710);
and U13041 (N_13041,N_11884,N_11996);
nand U13042 (N_13042,N_11093,N_11873);
nand U13043 (N_13043,N_10684,N_11967);
xor U13044 (N_13044,N_10755,N_11218);
or U13045 (N_13045,N_11671,N_11632);
nand U13046 (N_13046,N_10700,N_11288);
xnor U13047 (N_13047,N_10597,N_11329);
nand U13048 (N_13048,N_10677,N_11600);
nor U13049 (N_13049,N_11822,N_11520);
nor U13050 (N_13050,N_11966,N_11214);
and U13051 (N_13051,N_10639,N_11844);
or U13052 (N_13052,N_10582,N_11287);
nand U13053 (N_13053,N_11529,N_11717);
nor U13054 (N_13054,N_10515,N_11085);
nor U13055 (N_13055,N_11077,N_11774);
or U13056 (N_13056,N_10629,N_10697);
nor U13057 (N_13057,N_11332,N_10820);
nand U13058 (N_13058,N_11297,N_11018);
nand U13059 (N_13059,N_11027,N_11544);
nor U13060 (N_13060,N_11786,N_11438);
or U13061 (N_13061,N_10582,N_11489);
nor U13062 (N_13062,N_11707,N_10709);
or U13063 (N_13063,N_10998,N_11927);
and U13064 (N_13064,N_11648,N_10744);
nor U13065 (N_13065,N_11289,N_11636);
and U13066 (N_13066,N_10596,N_11758);
nand U13067 (N_13067,N_10969,N_10939);
nor U13068 (N_13068,N_11133,N_11875);
nand U13069 (N_13069,N_10906,N_11552);
nor U13070 (N_13070,N_10724,N_11434);
and U13071 (N_13071,N_11508,N_11412);
nand U13072 (N_13072,N_10798,N_11568);
nand U13073 (N_13073,N_11408,N_11455);
and U13074 (N_13074,N_10911,N_10536);
nand U13075 (N_13075,N_11713,N_11581);
and U13076 (N_13076,N_11409,N_11542);
nand U13077 (N_13077,N_10771,N_11297);
nand U13078 (N_13078,N_11435,N_11131);
nand U13079 (N_13079,N_10916,N_11198);
and U13080 (N_13080,N_11445,N_11465);
nor U13081 (N_13081,N_10866,N_11093);
nand U13082 (N_13082,N_11460,N_10999);
xnor U13083 (N_13083,N_11413,N_10809);
nor U13084 (N_13084,N_11997,N_11950);
and U13085 (N_13085,N_11915,N_11799);
nor U13086 (N_13086,N_11305,N_11334);
or U13087 (N_13087,N_11295,N_11071);
and U13088 (N_13088,N_11144,N_11290);
nand U13089 (N_13089,N_10543,N_10698);
or U13090 (N_13090,N_11909,N_10640);
nand U13091 (N_13091,N_11631,N_11750);
nor U13092 (N_13092,N_11195,N_11061);
or U13093 (N_13093,N_11779,N_10556);
nand U13094 (N_13094,N_11345,N_11971);
nand U13095 (N_13095,N_11071,N_10897);
nand U13096 (N_13096,N_11440,N_11368);
nand U13097 (N_13097,N_11177,N_11241);
nand U13098 (N_13098,N_10766,N_11189);
nand U13099 (N_13099,N_10707,N_10678);
nor U13100 (N_13100,N_11442,N_11825);
or U13101 (N_13101,N_11033,N_11329);
and U13102 (N_13102,N_11901,N_10883);
or U13103 (N_13103,N_11423,N_11981);
nor U13104 (N_13104,N_11012,N_11287);
and U13105 (N_13105,N_10608,N_10990);
nand U13106 (N_13106,N_11747,N_11830);
nand U13107 (N_13107,N_10765,N_11548);
or U13108 (N_13108,N_11674,N_11225);
or U13109 (N_13109,N_11197,N_11258);
or U13110 (N_13110,N_10619,N_11195);
nand U13111 (N_13111,N_11555,N_10545);
or U13112 (N_13112,N_11541,N_10787);
or U13113 (N_13113,N_11382,N_11424);
or U13114 (N_13114,N_11632,N_11113);
nand U13115 (N_13115,N_11794,N_11860);
or U13116 (N_13116,N_11522,N_10902);
nand U13117 (N_13117,N_11053,N_10590);
nor U13118 (N_13118,N_10970,N_10652);
nor U13119 (N_13119,N_11742,N_10701);
nor U13120 (N_13120,N_10905,N_11483);
and U13121 (N_13121,N_11528,N_11771);
nand U13122 (N_13122,N_11072,N_11176);
or U13123 (N_13123,N_11908,N_10865);
nor U13124 (N_13124,N_10799,N_11220);
or U13125 (N_13125,N_11121,N_11903);
or U13126 (N_13126,N_10777,N_10959);
or U13127 (N_13127,N_11673,N_11890);
and U13128 (N_13128,N_10836,N_11528);
nand U13129 (N_13129,N_10923,N_11806);
and U13130 (N_13130,N_11204,N_11739);
and U13131 (N_13131,N_11792,N_10720);
or U13132 (N_13132,N_11350,N_11984);
nand U13133 (N_13133,N_11583,N_11035);
nand U13134 (N_13134,N_11418,N_11465);
nand U13135 (N_13135,N_10612,N_11067);
or U13136 (N_13136,N_11682,N_11375);
nand U13137 (N_13137,N_11508,N_10877);
or U13138 (N_13138,N_11617,N_10617);
nor U13139 (N_13139,N_11212,N_11048);
nand U13140 (N_13140,N_11633,N_11988);
xnor U13141 (N_13141,N_10842,N_11340);
or U13142 (N_13142,N_11975,N_10630);
nor U13143 (N_13143,N_11100,N_11586);
or U13144 (N_13144,N_11987,N_11260);
nor U13145 (N_13145,N_11582,N_11545);
and U13146 (N_13146,N_11603,N_11316);
nor U13147 (N_13147,N_11845,N_11071);
or U13148 (N_13148,N_10729,N_11927);
and U13149 (N_13149,N_11720,N_10629);
xnor U13150 (N_13150,N_10781,N_11117);
nand U13151 (N_13151,N_11902,N_10813);
xor U13152 (N_13152,N_11922,N_11189);
nor U13153 (N_13153,N_11959,N_11213);
and U13154 (N_13154,N_11500,N_11980);
and U13155 (N_13155,N_11627,N_10735);
nor U13156 (N_13156,N_11264,N_11299);
and U13157 (N_13157,N_11794,N_11387);
and U13158 (N_13158,N_11630,N_10878);
or U13159 (N_13159,N_11941,N_10705);
and U13160 (N_13160,N_11853,N_11822);
and U13161 (N_13161,N_11013,N_10521);
or U13162 (N_13162,N_11241,N_10595);
nand U13163 (N_13163,N_11416,N_11403);
and U13164 (N_13164,N_11206,N_11357);
nor U13165 (N_13165,N_11003,N_11272);
and U13166 (N_13166,N_11599,N_11910);
and U13167 (N_13167,N_11049,N_11617);
and U13168 (N_13168,N_10895,N_11353);
and U13169 (N_13169,N_11391,N_10900);
nor U13170 (N_13170,N_11568,N_11529);
and U13171 (N_13171,N_10895,N_11359);
and U13172 (N_13172,N_11093,N_11894);
and U13173 (N_13173,N_11158,N_10874);
or U13174 (N_13174,N_11162,N_10663);
and U13175 (N_13175,N_10757,N_10604);
or U13176 (N_13176,N_11400,N_11707);
or U13177 (N_13177,N_11843,N_11308);
nand U13178 (N_13178,N_11557,N_11011);
and U13179 (N_13179,N_11670,N_10949);
or U13180 (N_13180,N_11911,N_11294);
nand U13181 (N_13181,N_11317,N_10924);
or U13182 (N_13182,N_11308,N_11465);
and U13183 (N_13183,N_11750,N_11781);
and U13184 (N_13184,N_10769,N_11891);
nor U13185 (N_13185,N_11304,N_10910);
nor U13186 (N_13186,N_10736,N_11564);
or U13187 (N_13187,N_11292,N_11136);
nand U13188 (N_13188,N_11207,N_11655);
nand U13189 (N_13189,N_10713,N_10850);
or U13190 (N_13190,N_11379,N_11351);
nand U13191 (N_13191,N_10559,N_11559);
nor U13192 (N_13192,N_10797,N_11306);
or U13193 (N_13193,N_10928,N_10936);
or U13194 (N_13194,N_11115,N_11528);
nor U13195 (N_13195,N_10879,N_10728);
or U13196 (N_13196,N_11191,N_11454);
and U13197 (N_13197,N_11100,N_11907);
and U13198 (N_13198,N_10670,N_10891);
and U13199 (N_13199,N_10788,N_10894);
nor U13200 (N_13200,N_10770,N_10745);
nor U13201 (N_13201,N_10559,N_11954);
or U13202 (N_13202,N_10795,N_11431);
or U13203 (N_13203,N_11594,N_11555);
or U13204 (N_13204,N_11947,N_11454);
nand U13205 (N_13205,N_10853,N_11604);
or U13206 (N_13206,N_11683,N_10530);
nor U13207 (N_13207,N_11130,N_10572);
nor U13208 (N_13208,N_10570,N_11823);
nand U13209 (N_13209,N_11242,N_11211);
nand U13210 (N_13210,N_10890,N_10793);
nand U13211 (N_13211,N_11341,N_10617);
and U13212 (N_13212,N_11826,N_11011);
nand U13213 (N_13213,N_11731,N_11934);
nor U13214 (N_13214,N_11800,N_11615);
nand U13215 (N_13215,N_11696,N_11969);
xnor U13216 (N_13216,N_11327,N_11439);
nor U13217 (N_13217,N_10742,N_11109);
or U13218 (N_13218,N_10770,N_11757);
nand U13219 (N_13219,N_11587,N_10882);
or U13220 (N_13220,N_11769,N_11658);
nand U13221 (N_13221,N_10731,N_11038);
nor U13222 (N_13222,N_11153,N_11583);
or U13223 (N_13223,N_11847,N_11148);
and U13224 (N_13224,N_10950,N_11905);
nand U13225 (N_13225,N_11673,N_10975);
nor U13226 (N_13226,N_11471,N_10735);
nand U13227 (N_13227,N_11839,N_10547);
or U13228 (N_13228,N_11944,N_11126);
or U13229 (N_13229,N_10981,N_11374);
or U13230 (N_13230,N_11158,N_11320);
nor U13231 (N_13231,N_10840,N_11854);
or U13232 (N_13232,N_11639,N_10900);
and U13233 (N_13233,N_10839,N_11078);
nor U13234 (N_13234,N_10558,N_11919);
nand U13235 (N_13235,N_11609,N_10801);
and U13236 (N_13236,N_11058,N_10869);
xor U13237 (N_13237,N_10669,N_11253);
or U13238 (N_13238,N_11463,N_11751);
nor U13239 (N_13239,N_11082,N_11266);
nand U13240 (N_13240,N_11316,N_10915);
and U13241 (N_13241,N_11642,N_11471);
and U13242 (N_13242,N_11583,N_10826);
or U13243 (N_13243,N_11074,N_11233);
nand U13244 (N_13244,N_11920,N_10916);
and U13245 (N_13245,N_10547,N_11680);
and U13246 (N_13246,N_11952,N_11142);
nor U13247 (N_13247,N_11245,N_11280);
nor U13248 (N_13248,N_11076,N_11643);
nand U13249 (N_13249,N_11221,N_11860);
nand U13250 (N_13250,N_11010,N_11660);
nor U13251 (N_13251,N_11899,N_11961);
nand U13252 (N_13252,N_11568,N_11388);
and U13253 (N_13253,N_11493,N_11343);
and U13254 (N_13254,N_10529,N_11717);
nand U13255 (N_13255,N_10799,N_10520);
and U13256 (N_13256,N_11891,N_11680);
nor U13257 (N_13257,N_11818,N_11283);
nor U13258 (N_13258,N_11131,N_11712);
and U13259 (N_13259,N_10622,N_11184);
or U13260 (N_13260,N_10896,N_11390);
or U13261 (N_13261,N_11555,N_11518);
and U13262 (N_13262,N_11774,N_10969);
nand U13263 (N_13263,N_11107,N_11632);
or U13264 (N_13264,N_11833,N_10802);
nand U13265 (N_13265,N_11615,N_10518);
or U13266 (N_13266,N_10598,N_11442);
nor U13267 (N_13267,N_11901,N_11219);
nand U13268 (N_13268,N_11235,N_11060);
nor U13269 (N_13269,N_10965,N_10576);
xnor U13270 (N_13270,N_11488,N_10794);
or U13271 (N_13271,N_10609,N_11712);
nor U13272 (N_13272,N_11747,N_11862);
or U13273 (N_13273,N_11564,N_11090);
nand U13274 (N_13274,N_11254,N_10908);
nor U13275 (N_13275,N_11701,N_11412);
xnor U13276 (N_13276,N_10965,N_11703);
or U13277 (N_13277,N_11240,N_10669);
nor U13278 (N_13278,N_11876,N_11047);
nor U13279 (N_13279,N_11412,N_10591);
xor U13280 (N_13280,N_10645,N_11014);
nand U13281 (N_13281,N_11261,N_11094);
nor U13282 (N_13282,N_11548,N_10585);
nand U13283 (N_13283,N_11923,N_11547);
nor U13284 (N_13284,N_11231,N_10900);
or U13285 (N_13285,N_11254,N_10619);
or U13286 (N_13286,N_11041,N_11822);
nand U13287 (N_13287,N_11968,N_11217);
nor U13288 (N_13288,N_10645,N_11314);
or U13289 (N_13289,N_11599,N_10975);
nand U13290 (N_13290,N_11324,N_10980);
nor U13291 (N_13291,N_10829,N_10875);
or U13292 (N_13292,N_11043,N_11736);
or U13293 (N_13293,N_10937,N_10692);
or U13294 (N_13294,N_10653,N_11202);
or U13295 (N_13295,N_11531,N_11190);
and U13296 (N_13296,N_11729,N_10928);
nand U13297 (N_13297,N_10514,N_11826);
and U13298 (N_13298,N_10993,N_11078);
or U13299 (N_13299,N_11327,N_10508);
and U13300 (N_13300,N_11652,N_11347);
nand U13301 (N_13301,N_11622,N_10743);
nor U13302 (N_13302,N_11768,N_11088);
or U13303 (N_13303,N_11158,N_10595);
and U13304 (N_13304,N_11372,N_11429);
or U13305 (N_13305,N_10573,N_11634);
or U13306 (N_13306,N_11061,N_11233);
nor U13307 (N_13307,N_10981,N_11681);
nor U13308 (N_13308,N_10595,N_11849);
nor U13309 (N_13309,N_11452,N_11524);
and U13310 (N_13310,N_11282,N_10584);
nor U13311 (N_13311,N_11133,N_11663);
and U13312 (N_13312,N_11791,N_11561);
nor U13313 (N_13313,N_11086,N_10649);
and U13314 (N_13314,N_11370,N_10500);
nor U13315 (N_13315,N_11629,N_11822);
nor U13316 (N_13316,N_10803,N_10505);
and U13317 (N_13317,N_10873,N_11262);
and U13318 (N_13318,N_11005,N_11820);
and U13319 (N_13319,N_11405,N_11242);
nor U13320 (N_13320,N_10536,N_10865);
and U13321 (N_13321,N_10592,N_11028);
nand U13322 (N_13322,N_11097,N_11055);
nor U13323 (N_13323,N_11259,N_10928);
or U13324 (N_13324,N_11563,N_11742);
and U13325 (N_13325,N_10579,N_10989);
nand U13326 (N_13326,N_11519,N_11907);
nor U13327 (N_13327,N_11129,N_11934);
or U13328 (N_13328,N_10707,N_11296);
xnor U13329 (N_13329,N_11832,N_11959);
nand U13330 (N_13330,N_11154,N_10504);
nor U13331 (N_13331,N_11006,N_10821);
and U13332 (N_13332,N_10615,N_11025);
nor U13333 (N_13333,N_11756,N_10794);
or U13334 (N_13334,N_11824,N_11712);
or U13335 (N_13335,N_10516,N_11757);
nor U13336 (N_13336,N_11040,N_11693);
nor U13337 (N_13337,N_10795,N_11198);
nor U13338 (N_13338,N_10656,N_10653);
nand U13339 (N_13339,N_11692,N_11238);
nor U13340 (N_13340,N_11361,N_10528);
nand U13341 (N_13341,N_11248,N_11074);
and U13342 (N_13342,N_11779,N_11696);
or U13343 (N_13343,N_10797,N_11947);
or U13344 (N_13344,N_10573,N_11342);
or U13345 (N_13345,N_11431,N_11322);
or U13346 (N_13346,N_10825,N_10909);
or U13347 (N_13347,N_10999,N_10920);
nand U13348 (N_13348,N_11896,N_11230);
and U13349 (N_13349,N_11285,N_10763);
nor U13350 (N_13350,N_11959,N_10994);
nor U13351 (N_13351,N_10726,N_11663);
nand U13352 (N_13352,N_11447,N_10591);
nand U13353 (N_13353,N_10842,N_11099);
or U13354 (N_13354,N_11307,N_11119);
nor U13355 (N_13355,N_11506,N_11095);
nand U13356 (N_13356,N_11201,N_11301);
nand U13357 (N_13357,N_10664,N_11901);
and U13358 (N_13358,N_11215,N_10560);
and U13359 (N_13359,N_10682,N_10806);
nand U13360 (N_13360,N_11039,N_11413);
nor U13361 (N_13361,N_11360,N_10786);
or U13362 (N_13362,N_10798,N_11789);
or U13363 (N_13363,N_11731,N_10916);
and U13364 (N_13364,N_10529,N_11804);
nor U13365 (N_13365,N_11606,N_11768);
nand U13366 (N_13366,N_10581,N_11576);
or U13367 (N_13367,N_10963,N_11328);
or U13368 (N_13368,N_10875,N_10968);
or U13369 (N_13369,N_10733,N_10588);
and U13370 (N_13370,N_10680,N_11321);
nand U13371 (N_13371,N_11584,N_10851);
or U13372 (N_13372,N_11077,N_11013);
or U13373 (N_13373,N_11254,N_10667);
and U13374 (N_13374,N_11386,N_10906);
or U13375 (N_13375,N_11988,N_10782);
and U13376 (N_13376,N_11397,N_11646);
nand U13377 (N_13377,N_10509,N_11587);
nand U13378 (N_13378,N_10651,N_11511);
nand U13379 (N_13379,N_11529,N_11282);
or U13380 (N_13380,N_11571,N_10855);
and U13381 (N_13381,N_11001,N_10521);
nor U13382 (N_13382,N_11016,N_11707);
and U13383 (N_13383,N_11717,N_11644);
nor U13384 (N_13384,N_11596,N_10873);
nand U13385 (N_13385,N_10998,N_11768);
nand U13386 (N_13386,N_11389,N_11777);
and U13387 (N_13387,N_11431,N_10966);
or U13388 (N_13388,N_10565,N_10684);
nand U13389 (N_13389,N_11893,N_11316);
nand U13390 (N_13390,N_10991,N_11708);
nor U13391 (N_13391,N_10946,N_10548);
or U13392 (N_13392,N_11655,N_10850);
and U13393 (N_13393,N_11895,N_11722);
nor U13394 (N_13394,N_11097,N_11650);
or U13395 (N_13395,N_11098,N_11673);
and U13396 (N_13396,N_11028,N_11810);
and U13397 (N_13397,N_11225,N_10721);
xor U13398 (N_13398,N_11082,N_10634);
nor U13399 (N_13399,N_11569,N_11118);
nor U13400 (N_13400,N_11897,N_10777);
nor U13401 (N_13401,N_11028,N_10550);
nor U13402 (N_13402,N_11936,N_10772);
and U13403 (N_13403,N_10843,N_10579);
or U13404 (N_13404,N_11504,N_10729);
nor U13405 (N_13405,N_10966,N_11974);
and U13406 (N_13406,N_10640,N_11161);
or U13407 (N_13407,N_11209,N_11655);
and U13408 (N_13408,N_10894,N_10763);
nor U13409 (N_13409,N_11307,N_11447);
nand U13410 (N_13410,N_10712,N_11582);
nand U13411 (N_13411,N_10793,N_11461);
and U13412 (N_13412,N_11495,N_10683);
or U13413 (N_13413,N_11424,N_10818);
and U13414 (N_13414,N_11370,N_11433);
or U13415 (N_13415,N_11017,N_11964);
nand U13416 (N_13416,N_11762,N_10628);
and U13417 (N_13417,N_11187,N_10937);
nor U13418 (N_13418,N_11603,N_10778);
or U13419 (N_13419,N_11399,N_11241);
or U13420 (N_13420,N_11697,N_10732);
or U13421 (N_13421,N_11006,N_11445);
or U13422 (N_13422,N_11685,N_10799);
or U13423 (N_13423,N_10788,N_10646);
or U13424 (N_13424,N_11660,N_11995);
nand U13425 (N_13425,N_11699,N_11074);
and U13426 (N_13426,N_11945,N_10691);
or U13427 (N_13427,N_11421,N_10815);
nor U13428 (N_13428,N_10513,N_10709);
or U13429 (N_13429,N_11882,N_10798);
or U13430 (N_13430,N_11722,N_10805);
nor U13431 (N_13431,N_11514,N_11506);
or U13432 (N_13432,N_11225,N_11398);
nor U13433 (N_13433,N_10935,N_11528);
nand U13434 (N_13434,N_11654,N_11550);
nor U13435 (N_13435,N_11660,N_10738);
nor U13436 (N_13436,N_10764,N_11036);
nand U13437 (N_13437,N_11177,N_11650);
nor U13438 (N_13438,N_11278,N_11353);
nand U13439 (N_13439,N_11807,N_10680);
or U13440 (N_13440,N_10542,N_11987);
nand U13441 (N_13441,N_11641,N_11481);
nand U13442 (N_13442,N_10803,N_11571);
and U13443 (N_13443,N_11788,N_11789);
and U13444 (N_13444,N_11210,N_10999);
nor U13445 (N_13445,N_10915,N_11798);
and U13446 (N_13446,N_10608,N_11734);
nor U13447 (N_13447,N_10718,N_11258);
nand U13448 (N_13448,N_10585,N_11567);
nor U13449 (N_13449,N_11879,N_11959);
or U13450 (N_13450,N_11683,N_10722);
and U13451 (N_13451,N_11097,N_10609);
or U13452 (N_13452,N_10886,N_11961);
nor U13453 (N_13453,N_11703,N_10763);
nor U13454 (N_13454,N_10669,N_11757);
nand U13455 (N_13455,N_11705,N_11027);
and U13456 (N_13456,N_11355,N_11456);
or U13457 (N_13457,N_11416,N_10811);
nand U13458 (N_13458,N_11956,N_10588);
and U13459 (N_13459,N_11658,N_10538);
nand U13460 (N_13460,N_10976,N_10509);
or U13461 (N_13461,N_10554,N_11232);
nand U13462 (N_13462,N_11874,N_11754);
or U13463 (N_13463,N_10595,N_10980);
and U13464 (N_13464,N_11621,N_10952);
or U13465 (N_13465,N_10628,N_11187);
nand U13466 (N_13466,N_11275,N_10996);
or U13467 (N_13467,N_10867,N_10577);
and U13468 (N_13468,N_11030,N_11744);
nor U13469 (N_13469,N_10593,N_11620);
and U13470 (N_13470,N_11766,N_11837);
and U13471 (N_13471,N_11965,N_11984);
nor U13472 (N_13472,N_11913,N_10879);
nand U13473 (N_13473,N_11831,N_11353);
nand U13474 (N_13474,N_11934,N_11369);
or U13475 (N_13475,N_11730,N_11966);
nand U13476 (N_13476,N_10848,N_11729);
nor U13477 (N_13477,N_11509,N_10779);
and U13478 (N_13478,N_11595,N_11660);
nor U13479 (N_13479,N_11940,N_10899);
nor U13480 (N_13480,N_11136,N_11950);
nor U13481 (N_13481,N_11469,N_10901);
nand U13482 (N_13482,N_10922,N_11040);
and U13483 (N_13483,N_11382,N_11408);
nand U13484 (N_13484,N_11861,N_11054);
nor U13485 (N_13485,N_11320,N_11054);
nor U13486 (N_13486,N_11883,N_11202);
nand U13487 (N_13487,N_11261,N_11759);
nand U13488 (N_13488,N_11174,N_10727);
nor U13489 (N_13489,N_11148,N_11612);
nand U13490 (N_13490,N_11059,N_11796);
nor U13491 (N_13491,N_11601,N_11004);
or U13492 (N_13492,N_11439,N_10786);
and U13493 (N_13493,N_11523,N_11020);
and U13494 (N_13494,N_11908,N_10549);
or U13495 (N_13495,N_11151,N_11324);
nor U13496 (N_13496,N_10990,N_10734);
or U13497 (N_13497,N_11994,N_11820);
and U13498 (N_13498,N_11688,N_11176);
or U13499 (N_13499,N_11162,N_11776);
nor U13500 (N_13500,N_12504,N_12660);
or U13501 (N_13501,N_13300,N_13019);
nand U13502 (N_13502,N_12211,N_12711);
or U13503 (N_13503,N_13108,N_12867);
nand U13504 (N_13504,N_12721,N_13177);
or U13505 (N_13505,N_12037,N_12489);
xor U13506 (N_13506,N_12180,N_13048);
or U13507 (N_13507,N_12745,N_13180);
or U13508 (N_13508,N_12222,N_12031);
nor U13509 (N_13509,N_12337,N_12879);
nor U13510 (N_13510,N_12420,N_13020);
and U13511 (N_13511,N_12573,N_12136);
xnor U13512 (N_13512,N_13473,N_12321);
or U13513 (N_13513,N_12816,N_12555);
xor U13514 (N_13514,N_13438,N_13006);
nand U13515 (N_13515,N_13488,N_12778);
nor U13516 (N_13516,N_13160,N_12216);
nand U13517 (N_13517,N_13039,N_12311);
or U13518 (N_13518,N_12923,N_13243);
and U13519 (N_13519,N_12455,N_12052);
nor U13520 (N_13520,N_12678,N_12303);
nand U13521 (N_13521,N_12353,N_13320);
nand U13522 (N_13522,N_12163,N_13178);
nand U13523 (N_13523,N_13443,N_13237);
nand U13524 (N_13524,N_13087,N_13301);
nor U13525 (N_13525,N_12731,N_12483);
or U13526 (N_13526,N_12354,N_12265);
nor U13527 (N_13527,N_12374,N_12545);
nor U13528 (N_13528,N_13088,N_12224);
nor U13529 (N_13529,N_13134,N_13093);
nand U13530 (N_13530,N_12960,N_12677);
nor U13531 (N_13531,N_13421,N_13281);
nor U13532 (N_13532,N_12655,N_12727);
and U13533 (N_13533,N_12911,N_12925);
nand U13534 (N_13534,N_12623,N_13480);
and U13535 (N_13535,N_12498,N_12700);
nand U13536 (N_13536,N_12631,N_13106);
and U13537 (N_13537,N_12949,N_13450);
nand U13538 (N_13538,N_12134,N_12038);
nand U13539 (N_13539,N_12964,N_12282);
nand U13540 (N_13540,N_12517,N_13433);
or U13541 (N_13541,N_12608,N_13241);
and U13542 (N_13542,N_13377,N_12369);
or U13543 (N_13543,N_12034,N_13342);
or U13544 (N_13544,N_13361,N_12690);
nand U13545 (N_13545,N_13169,N_12772);
and U13546 (N_13546,N_12903,N_12006);
nor U13547 (N_13547,N_12326,N_12330);
nand U13548 (N_13548,N_12575,N_13234);
or U13549 (N_13549,N_12680,N_12133);
nand U13550 (N_13550,N_12512,N_13110);
nand U13551 (N_13551,N_12348,N_12790);
nor U13552 (N_13552,N_12984,N_12809);
and U13553 (N_13553,N_12007,N_12782);
or U13554 (N_13554,N_13034,N_13486);
and U13555 (N_13555,N_13332,N_13121);
and U13556 (N_13556,N_12229,N_13145);
nand U13557 (N_13557,N_12565,N_12981);
nor U13558 (N_13558,N_13416,N_12264);
or U13559 (N_13559,N_12233,N_12568);
and U13560 (N_13560,N_12576,N_12689);
nor U13561 (N_13561,N_13076,N_12030);
and U13562 (N_13562,N_12709,N_13477);
xor U13563 (N_13563,N_12556,N_12055);
or U13564 (N_13564,N_12161,N_12705);
nand U13565 (N_13565,N_12550,N_13310);
and U13566 (N_13566,N_13408,N_12827);
nor U13567 (N_13567,N_13347,N_13256);
or U13568 (N_13568,N_13203,N_13367);
or U13569 (N_13569,N_13312,N_12651);
or U13570 (N_13570,N_12848,N_13189);
nand U13571 (N_13571,N_12472,N_12160);
or U13572 (N_13572,N_13061,N_13068);
and U13573 (N_13573,N_12214,N_12875);
or U13574 (N_13574,N_12452,N_13335);
and U13575 (N_13575,N_12273,N_12889);
or U13576 (N_13576,N_12215,N_13456);
nand U13577 (N_13577,N_12488,N_13200);
and U13578 (N_13578,N_12208,N_13182);
or U13579 (N_13579,N_12863,N_13403);
or U13580 (N_13580,N_13454,N_13357);
or U13581 (N_13581,N_12289,N_13100);
and U13582 (N_13582,N_12595,N_13334);
or U13583 (N_13583,N_12364,N_12377);
nor U13584 (N_13584,N_13343,N_12511);
and U13585 (N_13585,N_12694,N_12438);
nand U13586 (N_13586,N_13165,N_12996);
or U13587 (N_13587,N_12917,N_13038);
or U13588 (N_13588,N_13058,N_13043);
or U13589 (N_13589,N_12372,N_12020);
nor U13590 (N_13590,N_12195,N_12248);
nand U13591 (N_13591,N_13054,N_12724);
or U13592 (N_13592,N_13140,N_12450);
nor U13593 (N_13593,N_12636,N_12688);
or U13594 (N_13594,N_12434,N_13468);
and U13595 (N_13595,N_12082,N_12642);
or U13596 (N_13596,N_12999,N_12335);
or U13597 (N_13597,N_12393,N_12704);
and U13598 (N_13598,N_12687,N_12669);
and U13599 (N_13599,N_13164,N_12184);
nand U13600 (N_13600,N_12640,N_12850);
or U13601 (N_13601,N_12402,N_12176);
nand U13602 (N_13602,N_12998,N_12341);
nor U13603 (N_13603,N_12017,N_12625);
nand U13604 (N_13604,N_12773,N_12141);
or U13605 (N_13605,N_12183,N_12127);
nor U13606 (N_13606,N_13149,N_12937);
nor U13607 (N_13607,N_12097,N_13081);
nand U13608 (N_13608,N_12427,N_12532);
or U13609 (N_13609,N_12054,N_13044);
nor U13610 (N_13610,N_12805,N_13172);
or U13611 (N_13611,N_12983,N_12574);
nand U13612 (N_13612,N_12413,N_12632);
or U13613 (N_13613,N_13445,N_12205);
or U13614 (N_13614,N_12293,N_12794);
nand U13615 (N_13615,N_13230,N_13330);
and U13616 (N_13616,N_12061,N_13244);
nor U13617 (N_13617,N_12333,N_13337);
and U13618 (N_13618,N_12280,N_12598);
nor U13619 (N_13619,N_12405,N_12516);
nand U13620 (N_13620,N_12622,N_12548);
nor U13621 (N_13621,N_13092,N_13114);
and U13622 (N_13622,N_12347,N_13078);
and U13623 (N_13623,N_12720,N_12828);
nor U13624 (N_13624,N_12065,N_13295);
nor U13625 (N_13625,N_13036,N_13358);
and U13626 (N_13626,N_12080,N_12649);
or U13627 (N_13627,N_12430,N_12467);
and U13628 (N_13628,N_12398,N_12587);
and U13629 (N_13629,N_12840,N_12066);
and U13630 (N_13630,N_12317,N_12087);
or U13631 (N_13631,N_13344,N_12787);
nand U13632 (N_13632,N_12630,N_12947);
or U13633 (N_13633,N_13063,N_13369);
and U13634 (N_13634,N_12566,N_12744);
nand U13635 (N_13635,N_12880,N_12775);
or U13636 (N_13636,N_12792,N_12712);
and U13637 (N_13637,N_13429,N_12639);
nor U13638 (N_13638,N_12750,N_13419);
nor U13639 (N_13639,N_12121,N_12808);
nor U13640 (N_13640,N_12301,N_13341);
and U13641 (N_13641,N_13207,N_13208);
and U13642 (N_13642,N_12919,N_12883);
nand U13643 (N_13643,N_12841,N_12838);
and U13644 (N_13644,N_12192,N_12886);
or U13645 (N_13645,N_12111,N_12081);
and U13646 (N_13646,N_13352,N_12203);
or U13647 (N_13647,N_12329,N_13440);
nor U13648 (N_13648,N_12915,N_12612);
nor U13649 (N_13649,N_12225,N_12285);
nor U13650 (N_13650,N_12779,N_12118);
nand U13651 (N_13651,N_12601,N_12547);
and U13652 (N_13652,N_13356,N_13015);
xnor U13653 (N_13653,N_12327,N_12737);
nand U13654 (N_13654,N_13292,N_12796);
nor U13655 (N_13655,N_12473,N_12410);
nand U13656 (N_13656,N_12922,N_13112);
or U13657 (N_13657,N_13424,N_12012);
or U13658 (N_13658,N_12159,N_12425);
nand U13659 (N_13659,N_13027,N_13469);
or U13660 (N_13660,N_12124,N_12484);
nand U13661 (N_13661,N_13026,N_12943);
nor U13662 (N_13662,N_12091,N_12619);
nand U13663 (N_13663,N_12200,N_12696);
nand U13664 (N_13664,N_12708,N_12780);
nand U13665 (N_13665,N_13236,N_12461);
nand U13666 (N_13666,N_12620,N_12953);
nor U13667 (N_13667,N_12093,N_13364);
nand U13668 (N_13668,N_12368,N_12380);
or U13669 (N_13669,N_12697,N_13302);
nand U13670 (N_13670,N_13251,N_12256);
nand U13671 (N_13671,N_12637,N_12186);
and U13672 (N_13672,N_12833,N_12825);
xor U13673 (N_13673,N_13472,N_13359);
or U13674 (N_13674,N_12172,N_12339);
nor U13675 (N_13675,N_12157,N_12820);
nor U13676 (N_13676,N_12359,N_12644);
and U13677 (N_13677,N_12344,N_13184);
and U13678 (N_13678,N_12352,N_12583);
nand U13679 (N_13679,N_12907,N_13289);
nor U13680 (N_13680,N_13072,N_12989);
or U13681 (N_13681,N_13288,N_12230);
xor U13682 (N_13682,N_12613,N_12336);
nand U13683 (N_13683,N_12652,N_12785);
and U13684 (N_13684,N_12024,N_13326);
and U13685 (N_13685,N_12499,N_12226);
and U13686 (N_13686,N_12429,N_13309);
or U13687 (N_13687,N_12039,N_13116);
nand U13688 (N_13688,N_13497,N_12509);
nor U13689 (N_13689,N_12490,N_13111);
and U13690 (N_13690,N_12788,N_12323);
nor U13691 (N_13691,N_12977,N_12607);
nor U13692 (N_13692,N_13217,N_12847);
and U13693 (N_13693,N_12213,N_13225);
nand U13694 (N_13694,N_13098,N_12997);
xor U13695 (N_13695,N_12432,N_13004);
nand U13696 (N_13696,N_12870,N_13401);
nand U13697 (N_13697,N_12560,N_12162);
nand U13698 (N_13698,N_13485,N_12518);
nand U13699 (N_13699,N_13386,N_13170);
and U13700 (N_13700,N_12759,N_13482);
nand U13701 (N_13701,N_12234,N_12581);
or U13702 (N_13702,N_12993,N_13452);
and U13703 (N_13703,N_12756,N_13261);
nand U13704 (N_13704,N_12223,N_12714);
nor U13705 (N_13705,N_12171,N_13460);
and U13706 (N_13706,N_13138,N_12921);
nand U13707 (N_13707,N_12807,N_12441);
nor U13708 (N_13708,N_13175,N_13388);
nor U13709 (N_13709,N_13423,N_12202);
nand U13710 (N_13710,N_12757,N_13284);
or U13711 (N_13711,N_12627,N_12194);
nor U13712 (N_13712,N_13147,N_13199);
nor U13713 (N_13713,N_13455,N_13340);
nand U13714 (N_13714,N_13391,N_12699);
nor U13715 (N_13715,N_12853,N_12670);
and U13716 (N_13716,N_12537,N_12324);
nor U13717 (N_13717,N_12113,N_13079);
or U13718 (N_13718,N_13329,N_12218);
nor U13719 (N_13719,N_12249,N_12536);
nor U13720 (N_13720,N_12956,N_12173);
nor U13721 (N_13721,N_12804,N_12274);
or U13722 (N_13722,N_13466,N_13254);
nor U13723 (N_13723,N_12236,N_13339);
and U13724 (N_13724,N_12154,N_12944);
or U13725 (N_13725,N_12514,N_13250);
and U13726 (N_13726,N_12331,N_12412);
or U13727 (N_13727,N_12417,N_13024);
nand U13728 (N_13728,N_12656,N_13205);
or U13729 (N_13729,N_12877,N_12148);
and U13730 (N_13730,N_12507,N_13148);
xnor U13731 (N_13731,N_12104,N_13349);
or U13732 (N_13732,N_12423,N_12152);
xor U13733 (N_13733,N_12358,N_12776);
and U13734 (N_13734,N_12296,N_12752);
or U13735 (N_13735,N_12174,N_12125);
nor U13736 (N_13736,N_12898,N_12023);
and U13737 (N_13737,N_12397,N_12932);
nor U13738 (N_13738,N_13303,N_12271);
nand U13739 (N_13739,N_12421,N_12408);
or U13740 (N_13740,N_12166,N_13018);
nor U13741 (N_13741,N_13035,N_12813);
xor U13742 (N_13742,N_12482,N_12829);
nand U13743 (N_13743,N_13346,N_13161);
or U13744 (N_13744,N_13047,N_12258);
nor U13745 (N_13745,N_12067,N_13327);
nand U13746 (N_13746,N_12307,N_12763);
and U13747 (N_13747,N_13226,N_13298);
nor U13748 (N_13748,N_13484,N_12090);
nor U13749 (N_13749,N_12664,N_12599);
nor U13750 (N_13750,N_12294,N_12422);
nand U13751 (N_13751,N_13458,N_12530);
nand U13752 (N_13752,N_12146,N_12854);
and U13753 (N_13753,N_12367,N_13181);
and U13754 (N_13754,N_12910,N_13461);
nand U13755 (N_13755,N_12147,N_12890);
nand U13756 (N_13756,N_12638,N_12095);
or U13757 (N_13757,N_13381,N_12340);
nand U13758 (N_13758,N_13360,N_12153);
nor U13759 (N_13759,N_12449,N_13496);
nor U13760 (N_13760,N_13224,N_12458);
nor U13761 (N_13761,N_12617,N_12962);
nand U13762 (N_13762,N_12501,N_12447);
nand U13763 (N_13763,N_12798,N_12971);
and U13764 (N_13764,N_12586,N_12199);
nor U13765 (N_13765,N_12343,N_12541);
nor U13766 (N_13766,N_13080,N_13476);
and U13767 (N_13767,N_13065,N_13060);
nor U13768 (N_13768,N_13259,N_12228);
or U13769 (N_13769,N_13030,N_12846);
or U13770 (N_13770,N_12526,N_12382);
or U13771 (N_13771,N_12291,N_12263);
nor U13772 (N_13772,N_12674,N_12279);
and U13773 (N_13773,N_12036,N_13464);
and U13774 (N_13774,N_12391,N_12938);
nor U13775 (N_13775,N_12399,N_12602);
or U13776 (N_13776,N_13307,N_12589);
nor U13777 (N_13777,N_12014,N_13316);
or U13778 (N_13778,N_12675,N_12201);
or U13779 (N_13779,N_13229,N_12857);
or U13780 (N_13780,N_12465,N_12513);
and U13781 (N_13781,N_12777,N_13328);
or U13782 (N_13782,N_13467,N_12924);
and U13783 (N_13783,N_13365,N_12247);
nand U13784 (N_13784,N_13252,N_12569);
nor U13785 (N_13785,N_13426,N_13444);
nand U13786 (N_13786,N_12663,N_13296);
and U13787 (N_13787,N_12156,N_12764);
nor U13788 (N_13788,N_12606,N_12005);
and U13789 (N_13789,N_13264,N_12760);
nor U13790 (N_13790,N_12004,N_13005);
and U13791 (N_13791,N_12206,N_13014);
and U13792 (N_13792,N_12059,N_12819);
and U13793 (N_13793,N_12308,N_12543);
and U13794 (N_13794,N_13071,N_12703);
nor U13795 (N_13795,N_12457,N_13406);
or U13796 (N_13796,N_12831,N_13490);
nand U13797 (N_13797,N_13331,N_13399);
and U13798 (N_13798,N_12320,N_13041);
nor U13799 (N_13799,N_13492,N_13449);
and U13800 (N_13800,N_12822,N_12693);
or U13801 (N_13801,N_12278,N_13413);
and U13802 (N_13802,N_13103,N_13032);
or U13803 (N_13803,N_12978,N_12232);
nand U13804 (N_13804,N_12085,N_12453);
nand U13805 (N_13805,N_13417,N_13314);
or U13806 (N_13806,N_12269,N_12428);
or U13807 (N_13807,N_12715,N_12535);
or U13808 (N_13808,N_12969,N_13168);
or U13809 (N_13809,N_12041,N_12832);
or U13810 (N_13810,N_13099,N_12089);
nand U13811 (N_13811,N_13091,N_12074);
nor U13812 (N_13812,N_12015,N_12237);
nor U13813 (N_13813,N_12316,N_12355);
nand U13814 (N_13814,N_12913,N_12839);
nor U13815 (N_13815,N_13193,N_12585);
and U13816 (N_13816,N_12360,N_12647);
or U13817 (N_13817,N_12468,N_12529);
or U13818 (N_13818,N_12298,N_12987);
nor U13819 (N_13819,N_12920,N_12609);
nand U13820 (N_13820,N_12615,N_13306);
or U13821 (N_13821,N_13368,N_12027);
nand U13822 (N_13822,N_13285,N_12295);
or U13823 (N_13823,N_12029,N_13129);
nand U13824 (N_13824,N_12770,N_12048);
or U13825 (N_13825,N_12844,N_12198);
or U13826 (N_13826,N_12454,N_12893);
nand U13827 (N_13827,N_12527,N_12685);
or U13828 (N_13828,N_12053,N_12753);
and U13829 (N_13829,N_13247,N_12350);
nor U13830 (N_13830,N_12897,N_13031);
nand U13831 (N_13831,N_13318,N_12251);
nor U13832 (N_13832,N_12865,N_12338);
nor U13833 (N_13833,N_13258,N_13475);
and U13834 (N_13834,N_12112,N_12667);
nor U13835 (N_13835,N_12178,N_13104);
nor U13836 (N_13836,N_12751,N_12071);
nand U13837 (N_13837,N_12561,N_12419);
nand U13838 (N_13838,N_13162,N_13394);
or U13839 (N_13839,N_13185,N_12092);
or U13840 (N_13840,N_13190,N_12858);
and U13841 (N_13841,N_12123,N_12105);
and U13842 (N_13842,N_12120,N_13102);
or U13843 (N_13843,N_13187,N_12106);
or U13844 (N_13844,N_12861,N_12765);
nand U13845 (N_13845,N_12456,N_12582);
nand U13846 (N_13846,N_12102,N_13436);
nor U13847 (N_13847,N_12035,N_13223);
nand U13848 (N_13848,N_13389,N_12477);
nand U13849 (N_13849,N_12662,N_12701);
and U13850 (N_13850,N_12723,N_12933);
or U13851 (N_13851,N_12741,N_13249);
and U13852 (N_13852,N_13397,N_12384);
and U13853 (N_13853,N_12390,N_13167);
and U13854 (N_13854,N_12754,N_12431);
or U13855 (N_13855,N_12313,N_12109);
nor U13856 (N_13856,N_12928,N_12657);
or U13857 (N_13857,N_12821,N_13297);
and U13858 (N_13858,N_12144,N_13246);
or U13859 (N_13859,N_12451,N_12876);
nor U13860 (N_13860,N_12003,N_12523);
nor U13861 (N_13861,N_12262,N_12722);
or U13862 (N_13862,N_12626,N_12781);
nor U13863 (N_13863,N_13348,N_13202);
and U13864 (N_13864,N_13253,N_12325);
and U13865 (N_13865,N_12444,N_13214);
nand U13866 (N_13866,N_12332,N_12872);
or U13867 (N_13867,N_12044,N_12869);
and U13868 (N_13868,N_12494,N_12577);
or U13869 (N_13869,N_12672,N_12165);
nand U13870 (N_13870,N_12261,N_12416);
and U13871 (N_13871,N_13291,N_13385);
nor U13872 (N_13872,N_13003,N_12835);
nand U13873 (N_13873,N_12758,N_12395);
xnor U13874 (N_13874,N_12578,N_13231);
or U13875 (N_13875,N_12659,N_12968);
and U13876 (N_13876,N_13268,N_13083);
nor U13877 (N_13877,N_12243,N_13070);
nor U13878 (N_13878,N_13384,N_12021);
and U13879 (N_13879,N_12272,N_12266);
and U13880 (N_13880,N_12736,N_13491);
or U13881 (N_13881,N_12719,N_13023);
and U13882 (N_13882,N_13393,N_13186);
nor U13883 (N_13883,N_12945,N_13299);
and U13884 (N_13884,N_13282,N_12603);
and U13885 (N_13885,N_12167,N_13151);
nor U13886 (N_13886,N_13382,N_12814);
and U13887 (N_13887,N_13028,N_13471);
and U13888 (N_13888,N_13235,N_12967);
nand U13889 (N_13889,N_12480,N_12025);
and U13890 (N_13890,N_12957,N_13267);
and U13891 (N_13891,N_12591,N_13324);
nor U13892 (N_13892,N_12057,N_12929);
nor U13893 (N_13893,N_12975,N_13373);
and U13894 (N_13894,N_12904,N_13355);
nor U13895 (N_13895,N_12558,N_13483);
or U13896 (N_13896,N_13045,N_12695);
xor U13897 (N_13897,N_13451,N_12826);
or U13898 (N_13898,N_12459,N_13398);
nand U13899 (N_13899,N_12096,N_12117);
or U13900 (N_13900,N_12169,N_13383);
and U13901 (N_13901,N_12842,N_12284);
and U13902 (N_13902,N_13412,N_12357);
and U13903 (N_13903,N_13228,N_13407);
nor U13904 (N_13904,N_12855,N_12346);
nor U13905 (N_13905,N_13453,N_12896);
and U13906 (N_13906,N_13010,N_13212);
nor U13907 (N_13907,N_12515,N_12905);
nand U13908 (N_13908,N_12769,N_12959);
and U13909 (N_13909,N_12492,N_12334);
nand U13910 (N_13910,N_12342,N_12707);
nand U13911 (N_13911,N_12318,N_12747);
or U13912 (N_13912,N_13410,N_12140);
nand U13913 (N_13913,N_13096,N_13074);
nand U13914 (N_13914,N_13159,N_12597);
nand U13915 (N_13915,N_13155,N_12995);
or U13916 (N_13916,N_13141,N_13125);
or U13917 (N_13917,N_12963,N_12834);
xor U13918 (N_13918,N_12553,N_13059);
and U13919 (N_13919,N_12376,N_13427);
and U13920 (N_13920,N_13378,N_12137);
and U13921 (N_13921,N_13494,N_12930);
xor U13922 (N_13922,N_13055,N_12463);
nand U13923 (N_13923,N_12524,N_12083);
and U13924 (N_13924,N_12610,N_12939);
or U13925 (N_13925,N_12126,N_12033);
nor U13926 (N_13926,N_12554,N_12802);
or U13927 (N_13927,N_13457,N_12019);
and U13928 (N_13928,N_12493,N_12221);
and U13929 (N_13929,N_12062,N_12666);
nor U13930 (N_13930,N_12155,N_12927);
nand U13931 (N_13931,N_13130,N_12193);
or U13932 (N_13932,N_12815,N_12950);
or U13933 (N_13933,N_13122,N_13422);
xnor U13934 (N_13934,N_12551,N_12860);
nor U13935 (N_13935,N_13150,N_12392);
and U13936 (N_13936,N_12735,N_12411);
nor U13937 (N_13937,N_12580,N_12966);
or U13938 (N_13938,N_12812,N_12179);
xor U13939 (N_13939,N_13489,N_13042);
or U13940 (N_13940,N_12795,N_12799);
or U13941 (N_13941,N_12985,N_12051);
or U13942 (N_13942,N_12309,N_13242);
nand U13943 (N_13943,N_12728,N_12437);
nand U13944 (N_13944,N_12426,N_12611);
and U13945 (N_13945,N_12227,N_13338);
or U13946 (N_13946,N_12182,N_12122);
nor U13947 (N_13947,N_12882,N_13153);
nand U13948 (N_13948,N_13188,N_13317);
nand U13949 (N_13949,N_12098,N_13374);
or U13950 (N_13950,N_12491,N_13211);
nor U13951 (N_13951,N_13126,N_12375);
or U13952 (N_13952,N_12542,N_13051);
and U13953 (N_13953,N_12259,N_13021);
nor U13954 (N_13954,N_12803,N_12668);
nand U13955 (N_13955,N_13294,N_13283);
nor U13956 (N_13956,N_12973,N_12116);
or U13957 (N_13957,N_12418,N_12016);
and U13958 (N_13958,N_12738,N_12972);
nor U13959 (N_13959,N_12557,N_12716);
xor U13960 (N_13960,N_12706,N_12885);
nand U13961 (N_13961,N_13409,N_13215);
or U13962 (N_13962,N_12563,N_12239);
or U13963 (N_13963,N_12594,N_12559);
nor U13964 (N_13964,N_12099,N_12908);
nor U13965 (N_13965,N_13025,N_12824);
or U13966 (N_13966,N_12740,N_12522);
nand U13967 (N_13967,N_12245,N_13481);
nor U13968 (N_13968,N_12531,N_12729);
nand U13969 (N_13969,N_12235,N_12789);
or U13970 (N_13970,N_13273,N_12653);
nor U13971 (N_13971,N_12665,N_12181);
nor U13972 (N_13972,N_12713,N_12864);
nand U13973 (N_13973,N_12887,N_13405);
or U13974 (N_13974,N_13431,N_13430);
or U13975 (N_13975,N_12433,N_12177);
nor U13976 (N_13976,N_12114,N_12884);
and U13977 (N_13977,N_12250,N_12866);
nor U13978 (N_13978,N_13323,N_13255);
nor U13979 (N_13979,N_13050,N_12732);
and U13980 (N_13980,N_12940,N_12648);
nor U13981 (N_13981,N_12242,N_12436);
nor U13982 (N_13982,N_13363,N_13428);
nand U13983 (N_13983,N_12845,N_12040);
nand U13984 (N_13984,N_13272,N_12361);
nor U13985 (N_13985,N_12935,N_12292);
nor U13986 (N_13986,N_13404,N_13442);
or U13987 (N_13987,N_13046,N_12286);
nor U13988 (N_13988,N_12682,N_12139);
xnor U13989 (N_13989,N_12443,N_13201);
xor U13990 (N_13990,N_12328,N_13269);
nand U13991 (N_13991,N_12151,N_13197);
nand U13992 (N_13992,N_12605,N_12698);
nor U13993 (N_13993,N_12733,N_12077);
nand U13994 (N_13994,N_12130,N_13090);
nor U13995 (N_13995,N_12231,N_13319);
or U13996 (N_13996,N_12064,N_12766);
nand U13997 (N_13997,N_12075,N_12414);
nor U13998 (N_13998,N_12614,N_12013);
or U13999 (N_13999,N_12115,N_13209);
or U14000 (N_14000,N_12952,N_13131);
or U14001 (N_14001,N_13013,N_12385);
nor U14002 (N_14002,N_12909,N_12806);
nor U14003 (N_14003,N_12549,N_12868);
or U14004 (N_14004,N_12767,N_13336);
and U14005 (N_14005,N_12439,N_13465);
or U14006 (N_14006,N_12579,N_12389);
nand U14007 (N_14007,N_13133,N_12388);
or U14008 (N_14008,N_13239,N_12002);
or U14009 (N_14009,N_12658,N_12238);
nor U14010 (N_14010,N_13139,N_13086);
nor U14011 (N_14011,N_13195,N_13144);
nor U14012 (N_14012,N_12888,N_13105);
and U14013 (N_14013,N_12260,N_12345);
nand U14014 (N_14014,N_12546,N_12001);
and U14015 (N_14015,N_12086,N_13196);
and U14016 (N_14016,N_13354,N_12894);
or U14017 (N_14017,N_12000,N_12830);
nand U14018 (N_14018,N_12381,N_12288);
nand U14019 (N_14019,N_12955,N_12710);
nor U14020 (N_14020,N_12101,N_13278);
nand U14021 (N_14021,N_12138,N_13400);
nand U14022 (N_14022,N_12299,N_12891);
and U14023 (N_14023,N_12068,N_12060);
nor U14024 (N_14024,N_12084,N_12994);
and U14025 (N_14025,N_12746,N_12976);
or U14026 (N_14026,N_12914,N_12783);
nor U14027 (N_14027,N_13432,N_12275);
nor U14028 (N_14028,N_13007,N_13263);
or U14029 (N_14029,N_12681,N_13115);
nand U14030 (N_14030,N_12045,N_13262);
or U14031 (N_14031,N_13441,N_12009);
or U14032 (N_14032,N_12965,N_12378);
nand U14033 (N_14033,N_13392,N_12982);
nand U14034 (N_14034,N_12257,N_12958);
nand U14035 (N_14035,N_13462,N_12646);
xor U14036 (N_14036,N_12297,N_12590);
and U14037 (N_14037,N_13163,N_12852);
or U14038 (N_14038,N_12533,N_12056);
or U14039 (N_14039,N_12470,N_12244);
and U14040 (N_14040,N_13402,N_12873);
nor U14041 (N_14041,N_12552,N_13265);
or U14042 (N_14042,N_13075,N_12487);
or U14043 (N_14043,N_13420,N_13089);
nand U14044 (N_14044,N_12363,N_13233);
nor U14045 (N_14045,N_12042,N_13128);
nand U14046 (N_14046,N_12592,N_13085);
nor U14047 (N_14047,N_12912,N_12679);
nand U14048 (N_14048,N_13179,N_12050);
and U14049 (N_14049,N_12691,N_13052);
nand U14050 (N_14050,N_12462,N_12508);
nor U14051 (N_14051,N_12209,N_12445);
or U14052 (N_14052,N_13220,N_12371);
and U14053 (N_14053,N_12604,N_12479);
or U14054 (N_14054,N_13311,N_13447);
nand U14055 (N_14055,N_12926,N_12650);
or U14056 (N_14056,N_12784,N_13000);
and U14057 (N_14057,N_13353,N_13062);
nand U14058 (N_14058,N_12768,N_12600);
or U14059 (N_14059,N_12862,N_13304);
and U14060 (N_14060,N_13375,N_12478);
nand U14061 (N_14061,N_12742,N_12175);
and U14062 (N_14062,N_13463,N_12135);
xnor U14063 (N_14063,N_12702,N_12974);
nand U14064 (N_14064,N_12683,N_12481);
nor U14065 (N_14065,N_13434,N_12076);
or U14066 (N_14066,N_12629,N_12145);
and U14067 (N_14067,N_12283,N_12817);
nand U14068 (N_14068,N_13204,N_12871);
nand U14069 (N_14069,N_12748,N_13321);
and U14070 (N_14070,N_12906,N_13439);
and U14071 (N_14071,N_12094,N_13280);
nand U14072 (N_14072,N_12219,N_13351);
nand U14073 (N_14073,N_13143,N_12217);
nand U14074 (N_14074,N_12270,N_12486);
and U14075 (N_14075,N_12310,N_12692);
or U14076 (N_14076,N_12621,N_12892);
nand U14077 (N_14077,N_12851,N_13156);
nand U14078 (N_14078,N_12749,N_13194);
nand U14079 (N_14079,N_13493,N_12899);
nor U14080 (N_14080,N_13276,N_12895);
nor U14081 (N_14081,N_12810,N_12837);
nor U14082 (N_14082,N_12520,N_13192);
or U14083 (N_14083,N_12500,N_12496);
nand U14084 (N_14084,N_13448,N_13056);
or U14085 (N_14085,N_12047,N_12440);
or U14086 (N_14086,N_12485,N_13411);
nand U14087 (N_14087,N_13136,N_13146);
nand U14088 (N_14088,N_13183,N_12349);
nand U14089 (N_14089,N_12633,N_12185);
nor U14090 (N_14090,N_12400,N_12761);
and U14091 (N_14091,N_12356,N_12801);
nor U14092 (N_14092,N_13227,N_12043);
and U14093 (N_14093,N_12103,N_13094);
and U14094 (N_14094,N_12635,N_13009);
and U14095 (N_14095,N_12407,N_13107);
nor U14096 (N_14096,N_13029,N_13124);
nor U14097 (N_14097,N_12132,N_13219);
nand U14098 (N_14098,N_12028,N_13418);
xor U14099 (N_14099,N_13206,N_12916);
nor U14100 (N_14100,N_12931,N_13174);
or U14101 (N_14101,N_12584,N_12951);
nand U14102 (N_14102,N_13037,N_13210);
or U14103 (N_14103,N_12464,N_12878);
or U14104 (N_14104,N_12717,N_12435);
and U14105 (N_14105,N_12220,N_12241);
nor U14106 (N_14106,N_13313,N_12191);
and U14107 (N_14107,N_12150,N_12188);
or U14108 (N_14108,N_13120,N_12197);
nand U14109 (N_14109,N_12918,N_12936);
or U14110 (N_14110,N_13415,N_12634);
and U14111 (N_14111,N_12018,N_12588);
nand U14112 (N_14112,N_12253,N_12624);
or U14113 (N_14113,N_13057,N_12401);
nor U14114 (N_14114,N_13345,N_12366);
nor U14115 (N_14115,N_12128,N_13333);
or U14116 (N_14116,N_12474,N_12394);
and U14117 (N_14117,N_12572,N_12811);
and U14118 (N_14118,N_12793,N_12528);
nor U14119 (N_14119,N_12786,N_12319);
nor U14120 (N_14120,N_13240,N_12628);
and U14121 (N_14121,N_12129,N_13154);
or U14122 (N_14122,N_13064,N_13118);
and U14123 (N_14123,N_12673,N_13371);
nor U14124 (N_14124,N_13101,N_13379);
or U14125 (N_14125,N_13248,N_13257);
and U14126 (N_14126,N_13470,N_12305);
nor U14127 (N_14127,N_12540,N_12149);
nor U14128 (N_14128,N_12990,N_12471);
nor U14129 (N_14129,N_12312,N_13277);
nor U14130 (N_14130,N_12946,N_12306);
or U14131 (N_14131,N_13376,N_12290);
nand U14132 (N_14132,N_13287,N_13171);
and U14133 (N_14133,N_13137,N_12460);
or U14134 (N_14134,N_12255,N_13390);
nor U14135 (N_14135,N_13123,N_13479);
nand U14136 (N_14136,N_12970,N_13366);
and U14137 (N_14137,N_13266,N_12506);
and U14138 (N_14138,N_12902,N_12900);
nor U14139 (N_14139,N_13487,N_12379);
nand U14140 (N_14140,N_13113,N_13437);
or U14141 (N_14141,N_12142,N_12654);
nand U14142 (N_14142,N_13372,N_12387);
nor U14143 (N_14143,N_12570,N_13380);
and U14144 (N_14144,N_12302,N_13222);
or U14145 (N_14145,N_13232,N_12100);
and U14146 (N_14146,N_12362,N_12403);
nand U14147 (N_14147,N_13033,N_13315);
nor U14148 (N_14148,N_12466,N_12158);
and U14149 (N_14149,N_12351,N_12797);
nor U14150 (N_14150,N_13260,N_12986);
or U14151 (N_14151,N_13176,N_12539);
or U14152 (N_14152,N_13077,N_12168);
nor U14153 (N_14153,N_12730,N_12643);
nor U14154 (N_14154,N_13305,N_12836);
or U14155 (N_14155,N_13040,N_13459);
nand U14156 (N_14156,N_12469,N_12934);
or U14157 (N_14157,N_12495,N_13198);
and U14158 (N_14158,N_13293,N_12774);
nor U14159 (N_14159,N_12510,N_12073);
or U14160 (N_14160,N_12645,N_13286);
or U14161 (N_14161,N_12196,N_12268);
and U14162 (N_14162,N_12415,N_13271);
xor U14163 (N_14163,N_13001,N_13308);
nor U14164 (N_14164,N_13218,N_13119);
or U14165 (N_14165,N_12901,N_13084);
and U14166 (N_14166,N_12818,N_12011);
or U14167 (N_14167,N_12596,N_12534);
and U14168 (N_14168,N_12755,N_12383);
nand U14169 (N_14169,N_12204,N_13008);
nand U14170 (N_14170,N_12448,N_13117);
nor U14171 (N_14171,N_13446,N_13082);
nand U14172 (N_14172,N_12277,N_12538);
nor U14173 (N_14173,N_12010,N_13474);
xor U14174 (N_14174,N_12373,N_12739);
nor U14175 (N_14175,N_13270,N_12521);
nand U14176 (N_14176,N_12370,N_13290);
nand U14177 (N_14177,N_13478,N_12386);
nand U14178 (N_14178,N_12856,N_12143);
and U14179 (N_14179,N_12190,N_13370);
and U14180 (N_14180,N_12032,N_12571);
and U14181 (N_14181,N_12254,N_12942);
and U14182 (N_14182,N_13069,N_12948);
and U14183 (N_14183,N_12164,N_12069);
nand U14184 (N_14184,N_13017,N_12503);
or U14185 (N_14185,N_13425,N_12771);
nor U14186 (N_14186,N_12131,N_12843);
nand U14187 (N_14187,N_13109,N_12008);
nor U14188 (N_14188,N_12671,N_12210);
or U14189 (N_14189,N_12276,N_12791);
nand U14190 (N_14190,N_13350,N_12304);
nand U14191 (N_14191,N_12859,N_12941);
or U14192 (N_14192,N_12979,N_12562);
or U14193 (N_14193,N_12980,N_12734);
xnor U14194 (N_14194,N_12564,N_13213);
and U14195 (N_14195,N_12189,N_12287);
nor U14196 (N_14196,N_13142,N_13011);
or U14197 (N_14197,N_13387,N_12525);
nor U14198 (N_14198,N_12988,N_12409);
and U14199 (N_14199,N_13275,N_12315);
and U14200 (N_14200,N_13322,N_13012);
nor U14201 (N_14201,N_12078,N_12406);
nand U14202 (N_14202,N_12475,N_12119);
nand U14203 (N_14203,N_12187,N_12281);
nand U14204 (N_14204,N_13216,N_13499);
and U14205 (N_14205,N_12661,N_13002);
or U14206 (N_14206,N_13362,N_13097);
nor U14207 (N_14207,N_13152,N_13279);
nor U14208 (N_14208,N_12686,N_12365);
xnor U14209 (N_14209,N_12108,N_12881);
nand U14210 (N_14210,N_13067,N_13135);
or U14211 (N_14211,N_13325,N_12641);
or U14212 (N_14212,N_12676,N_13016);
and U14213 (N_14213,N_13053,N_12849);
or U14214 (N_14214,N_13095,N_12743);
and U14215 (N_14215,N_13166,N_12207);
nor U14216 (N_14216,N_12726,N_12404);
or U14217 (N_14217,N_12476,N_12992);
nor U14218 (N_14218,N_12544,N_12107);
nor U14219 (N_14219,N_12424,N_12567);
nor U14220 (N_14220,N_12170,N_12593);
and U14221 (N_14221,N_12072,N_13396);
nor U14222 (N_14222,N_12212,N_13238);
nor U14223 (N_14223,N_12300,N_13191);
and U14224 (N_14224,N_12991,N_12442);
or U14225 (N_14225,N_12088,N_12497);
nand U14226 (N_14226,N_13158,N_13049);
xor U14227 (N_14227,N_12049,N_12618);
and U14228 (N_14228,N_12502,N_12616);
nor U14229 (N_14229,N_13157,N_13221);
nor U14230 (N_14230,N_12322,N_12519);
or U14231 (N_14231,N_12058,N_12800);
nand U14232 (N_14232,N_12063,N_12267);
or U14233 (N_14233,N_13127,N_12110);
and U14234 (N_14234,N_12252,N_12823);
or U14235 (N_14235,N_13132,N_12022);
nor U14236 (N_14236,N_13495,N_12079);
or U14237 (N_14237,N_13245,N_12396);
and U14238 (N_14238,N_12026,N_12874);
or U14239 (N_14239,N_12070,N_12246);
nand U14240 (N_14240,N_12046,N_13066);
and U14241 (N_14241,N_13274,N_12505);
xnor U14242 (N_14242,N_12684,N_13022);
nor U14243 (N_14243,N_12954,N_12240);
and U14244 (N_14244,N_12718,N_12446);
nor U14245 (N_14245,N_13435,N_13073);
xnor U14246 (N_14246,N_12961,N_12314);
or U14247 (N_14247,N_13395,N_12725);
or U14248 (N_14248,N_13498,N_13173);
or U14249 (N_14249,N_13414,N_12762);
and U14250 (N_14250,N_13308,N_12004);
nand U14251 (N_14251,N_12939,N_13409);
nor U14252 (N_14252,N_12480,N_13426);
and U14253 (N_14253,N_12264,N_12439);
nor U14254 (N_14254,N_13119,N_12328);
nand U14255 (N_14255,N_13413,N_13069);
and U14256 (N_14256,N_12478,N_12317);
xnor U14257 (N_14257,N_12335,N_12141);
and U14258 (N_14258,N_13091,N_12577);
nand U14259 (N_14259,N_13243,N_12208);
and U14260 (N_14260,N_12744,N_13292);
nand U14261 (N_14261,N_12694,N_12653);
and U14262 (N_14262,N_13317,N_13484);
and U14263 (N_14263,N_12876,N_12365);
or U14264 (N_14264,N_13293,N_13217);
and U14265 (N_14265,N_13497,N_12529);
or U14266 (N_14266,N_12792,N_12436);
nor U14267 (N_14267,N_12471,N_12951);
and U14268 (N_14268,N_13041,N_12822);
and U14269 (N_14269,N_13322,N_13453);
nor U14270 (N_14270,N_13467,N_12245);
and U14271 (N_14271,N_12546,N_12217);
nor U14272 (N_14272,N_12820,N_12102);
and U14273 (N_14273,N_12967,N_12555);
or U14274 (N_14274,N_13275,N_13217);
and U14275 (N_14275,N_12200,N_13082);
nand U14276 (N_14276,N_12091,N_12252);
nor U14277 (N_14277,N_13485,N_13368);
or U14278 (N_14278,N_12397,N_12799);
and U14279 (N_14279,N_12450,N_12581);
and U14280 (N_14280,N_12119,N_12425);
or U14281 (N_14281,N_12615,N_12901);
nand U14282 (N_14282,N_12428,N_13202);
nand U14283 (N_14283,N_12671,N_12401);
and U14284 (N_14284,N_13210,N_12897);
or U14285 (N_14285,N_12086,N_12654);
or U14286 (N_14286,N_13190,N_12280);
nand U14287 (N_14287,N_12977,N_13191);
nand U14288 (N_14288,N_12943,N_12337);
nand U14289 (N_14289,N_12285,N_12093);
or U14290 (N_14290,N_12707,N_13361);
and U14291 (N_14291,N_12563,N_13484);
or U14292 (N_14292,N_12031,N_12364);
or U14293 (N_14293,N_12870,N_13295);
nand U14294 (N_14294,N_12302,N_12084);
and U14295 (N_14295,N_13012,N_12364);
and U14296 (N_14296,N_12701,N_12600);
nand U14297 (N_14297,N_12344,N_12210);
nand U14298 (N_14298,N_12549,N_12731);
and U14299 (N_14299,N_13205,N_13487);
or U14300 (N_14300,N_12184,N_12912);
and U14301 (N_14301,N_12437,N_12470);
xor U14302 (N_14302,N_13234,N_12078);
or U14303 (N_14303,N_12495,N_13007);
and U14304 (N_14304,N_12023,N_12117);
nand U14305 (N_14305,N_12310,N_13350);
nor U14306 (N_14306,N_12765,N_12320);
nor U14307 (N_14307,N_12898,N_12518);
and U14308 (N_14308,N_12119,N_12464);
nand U14309 (N_14309,N_12701,N_13384);
or U14310 (N_14310,N_12762,N_13322);
nand U14311 (N_14311,N_12585,N_12437);
nand U14312 (N_14312,N_12503,N_12616);
nand U14313 (N_14313,N_12839,N_12344);
nor U14314 (N_14314,N_12025,N_12173);
and U14315 (N_14315,N_12627,N_12026);
nor U14316 (N_14316,N_12495,N_13058);
or U14317 (N_14317,N_12186,N_12599);
and U14318 (N_14318,N_12347,N_13095);
or U14319 (N_14319,N_12458,N_12967);
nor U14320 (N_14320,N_13139,N_12074);
nor U14321 (N_14321,N_12610,N_13106);
nor U14322 (N_14322,N_12379,N_12208);
or U14323 (N_14323,N_12336,N_12722);
nor U14324 (N_14324,N_12615,N_13023);
nor U14325 (N_14325,N_13423,N_12775);
or U14326 (N_14326,N_12134,N_12567);
nand U14327 (N_14327,N_13457,N_13216);
nand U14328 (N_14328,N_12890,N_13267);
and U14329 (N_14329,N_12957,N_13168);
nand U14330 (N_14330,N_12117,N_13356);
nand U14331 (N_14331,N_12845,N_13459);
or U14332 (N_14332,N_13360,N_12098);
nand U14333 (N_14333,N_12908,N_12024);
nand U14334 (N_14334,N_13358,N_12098);
and U14335 (N_14335,N_12219,N_13096);
nand U14336 (N_14336,N_13184,N_12073);
nand U14337 (N_14337,N_12023,N_12920);
or U14338 (N_14338,N_12217,N_12454);
and U14339 (N_14339,N_12665,N_13084);
or U14340 (N_14340,N_13294,N_12346);
nor U14341 (N_14341,N_13166,N_13152);
nor U14342 (N_14342,N_13315,N_12626);
nor U14343 (N_14343,N_12229,N_13075);
or U14344 (N_14344,N_12473,N_12111);
nand U14345 (N_14345,N_12227,N_13268);
or U14346 (N_14346,N_12642,N_12365);
nor U14347 (N_14347,N_13225,N_13396);
nor U14348 (N_14348,N_12475,N_12445);
nor U14349 (N_14349,N_12661,N_13106);
or U14350 (N_14350,N_12841,N_13184);
nor U14351 (N_14351,N_12300,N_12972);
nand U14352 (N_14352,N_12195,N_13079);
nor U14353 (N_14353,N_13390,N_12244);
or U14354 (N_14354,N_12827,N_13141);
nand U14355 (N_14355,N_12583,N_12945);
or U14356 (N_14356,N_12585,N_13176);
and U14357 (N_14357,N_12926,N_13480);
nand U14358 (N_14358,N_12136,N_13084);
nand U14359 (N_14359,N_12265,N_12613);
nand U14360 (N_14360,N_12707,N_12967);
or U14361 (N_14361,N_13152,N_13382);
and U14362 (N_14362,N_13433,N_12575);
nand U14363 (N_14363,N_13237,N_13078);
and U14364 (N_14364,N_13233,N_13037);
nor U14365 (N_14365,N_12609,N_12913);
or U14366 (N_14366,N_13211,N_13266);
nand U14367 (N_14367,N_12802,N_13271);
nor U14368 (N_14368,N_13299,N_12344);
nand U14369 (N_14369,N_13040,N_13224);
or U14370 (N_14370,N_12936,N_12114);
nand U14371 (N_14371,N_13349,N_13445);
and U14372 (N_14372,N_13160,N_13056);
nor U14373 (N_14373,N_13469,N_12212);
or U14374 (N_14374,N_12150,N_12983);
and U14375 (N_14375,N_12446,N_12096);
or U14376 (N_14376,N_12236,N_12612);
or U14377 (N_14377,N_12690,N_12142);
nor U14378 (N_14378,N_12380,N_12944);
nand U14379 (N_14379,N_12024,N_12573);
nand U14380 (N_14380,N_12491,N_13469);
and U14381 (N_14381,N_12561,N_12414);
or U14382 (N_14382,N_12696,N_13341);
nand U14383 (N_14383,N_12304,N_13071);
nor U14384 (N_14384,N_13437,N_12196);
or U14385 (N_14385,N_12499,N_12050);
and U14386 (N_14386,N_12638,N_13046);
and U14387 (N_14387,N_12851,N_12347);
or U14388 (N_14388,N_13063,N_12265);
nor U14389 (N_14389,N_12617,N_13165);
nor U14390 (N_14390,N_12114,N_12032);
or U14391 (N_14391,N_12897,N_12419);
and U14392 (N_14392,N_13136,N_12336);
and U14393 (N_14393,N_12910,N_12345);
and U14394 (N_14394,N_12709,N_12237);
and U14395 (N_14395,N_12153,N_12962);
nand U14396 (N_14396,N_12506,N_13246);
or U14397 (N_14397,N_12640,N_12260);
nor U14398 (N_14398,N_12505,N_12084);
nand U14399 (N_14399,N_12771,N_13325);
nand U14400 (N_14400,N_12594,N_12504);
nand U14401 (N_14401,N_12930,N_13019);
nand U14402 (N_14402,N_12196,N_12762);
nor U14403 (N_14403,N_12067,N_13395);
and U14404 (N_14404,N_13351,N_12955);
or U14405 (N_14405,N_12643,N_12330);
or U14406 (N_14406,N_12798,N_12618);
nor U14407 (N_14407,N_13393,N_12997);
nor U14408 (N_14408,N_12945,N_13058);
and U14409 (N_14409,N_13038,N_13297);
nand U14410 (N_14410,N_13425,N_12777);
or U14411 (N_14411,N_12596,N_13391);
nand U14412 (N_14412,N_12201,N_13427);
and U14413 (N_14413,N_12675,N_12898);
nor U14414 (N_14414,N_12260,N_12576);
nand U14415 (N_14415,N_13205,N_12312);
and U14416 (N_14416,N_12830,N_12036);
nor U14417 (N_14417,N_13057,N_13021);
or U14418 (N_14418,N_12579,N_13252);
and U14419 (N_14419,N_12967,N_12358);
or U14420 (N_14420,N_13215,N_12613);
nor U14421 (N_14421,N_12936,N_13189);
or U14422 (N_14422,N_12889,N_13078);
and U14423 (N_14423,N_12030,N_13050);
and U14424 (N_14424,N_13086,N_12529);
or U14425 (N_14425,N_12925,N_13325);
or U14426 (N_14426,N_12562,N_12364);
nand U14427 (N_14427,N_12304,N_13265);
nor U14428 (N_14428,N_12938,N_13066);
nand U14429 (N_14429,N_12699,N_13342);
xor U14430 (N_14430,N_13490,N_12744);
nand U14431 (N_14431,N_12230,N_13283);
nor U14432 (N_14432,N_13354,N_13246);
nor U14433 (N_14433,N_12006,N_12356);
nand U14434 (N_14434,N_13323,N_12983);
nand U14435 (N_14435,N_13294,N_13369);
or U14436 (N_14436,N_12603,N_12840);
nor U14437 (N_14437,N_12192,N_12234);
nand U14438 (N_14438,N_13093,N_12960);
nand U14439 (N_14439,N_12855,N_13168);
nor U14440 (N_14440,N_13154,N_12088);
nor U14441 (N_14441,N_12324,N_12622);
or U14442 (N_14442,N_13110,N_12703);
nor U14443 (N_14443,N_13073,N_13176);
or U14444 (N_14444,N_13304,N_12086);
nor U14445 (N_14445,N_12628,N_12444);
and U14446 (N_14446,N_12315,N_12604);
nor U14447 (N_14447,N_12417,N_13308);
nand U14448 (N_14448,N_13446,N_12987);
and U14449 (N_14449,N_12021,N_12004);
and U14450 (N_14450,N_12254,N_12507);
and U14451 (N_14451,N_13401,N_12478);
nor U14452 (N_14452,N_13305,N_12763);
nand U14453 (N_14453,N_13148,N_12105);
nand U14454 (N_14454,N_13379,N_12635);
nand U14455 (N_14455,N_13431,N_13203);
nand U14456 (N_14456,N_12895,N_12152);
nand U14457 (N_14457,N_12568,N_13222);
nor U14458 (N_14458,N_12213,N_12729);
nor U14459 (N_14459,N_12543,N_12888);
nor U14460 (N_14460,N_12045,N_13127);
xnor U14461 (N_14461,N_12202,N_13356);
nor U14462 (N_14462,N_12697,N_13113);
nand U14463 (N_14463,N_13299,N_12346);
or U14464 (N_14464,N_12650,N_12102);
or U14465 (N_14465,N_13218,N_12551);
or U14466 (N_14466,N_12508,N_12583);
or U14467 (N_14467,N_13101,N_12521);
nand U14468 (N_14468,N_12126,N_12986);
and U14469 (N_14469,N_12867,N_12468);
xor U14470 (N_14470,N_13374,N_12638);
nor U14471 (N_14471,N_13412,N_12837);
nor U14472 (N_14472,N_12386,N_13093);
nand U14473 (N_14473,N_13279,N_13175);
or U14474 (N_14474,N_12846,N_13025);
and U14475 (N_14475,N_12109,N_12010);
nor U14476 (N_14476,N_12032,N_12179);
or U14477 (N_14477,N_12138,N_12122);
nand U14478 (N_14478,N_12653,N_13087);
or U14479 (N_14479,N_13196,N_12446);
nor U14480 (N_14480,N_12958,N_12679);
or U14481 (N_14481,N_13384,N_13464);
or U14482 (N_14482,N_13344,N_12847);
and U14483 (N_14483,N_12513,N_13480);
and U14484 (N_14484,N_13100,N_12133);
and U14485 (N_14485,N_12053,N_12375);
or U14486 (N_14486,N_12017,N_12209);
or U14487 (N_14487,N_12530,N_12859);
and U14488 (N_14488,N_12894,N_13095);
nor U14489 (N_14489,N_13238,N_13416);
or U14490 (N_14490,N_12579,N_12910);
or U14491 (N_14491,N_12589,N_13085);
and U14492 (N_14492,N_13393,N_13333);
or U14493 (N_14493,N_12948,N_12851);
nor U14494 (N_14494,N_12750,N_12101);
or U14495 (N_14495,N_12350,N_13462);
nand U14496 (N_14496,N_12383,N_13029);
and U14497 (N_14497,N_13145,N_12797);
or U14498 (N_14498,N_12788,N_13071);
and U14499 (N_14499,N_12323,N_13216);
nand U14500 (N_14500,N_12626,N_12479);
nor U14501 (N_14501,N_13059,N_13128);
nand U14502 (N_14502,N_13257,N_12947);
nor U14503 (N_14503,N_12571,N_12972);
nand U14504 (N_14504,N_12884,N_12217);
or U14505 (N_14505,N_13350,N_13021);
nand U14506 (N_14506,N_13259,N_12859);
nand U14507 (N_14507,N_12678,N_12918);
nand U14508 (N_14508,N_13188,N_12023);
nand U14509 (N_14509,N_12654,N_12775);
or U14510 (N_14510,N_12235,N_12398);
nand U14511 (N_14511,N_13299,N_13303);
nand U14512 (N_14512,N_12528,N_12588);
or U14513 (N_14513,N_12927,N_12869);
nand U14514 (N_14514,N_12690,N_12480);
or U14515 (N_14515,N_12289,N_12864);
nand U14516 (N_14516,N_12463,N_12416);
nand U14517 (N_14517,N_13050,N_12446);
nand U14518 (N_14518,N_12005,N_12900);
or U14519 (N_14519,N_12755,N_12171);
nand U14520 (N_14520,N_12771,N_12940);
or U14521 (N_14521,N_13063,N_12824);
nor U14522 (N_14522,N_13239,N_12680);
or U14523 (N_14523,N_12186,N_13018);
nand U14524 (N_14524,N_13058,N_12086);
and U14525 (N_14525,N_12169,N_13385);
nor U14526 (N_14526,N_12469,N_12355);
nand U14527 (N_14527,N_13024,N_12818);
xor U14528 (N_14528,N_12660,N_13242);
or U14529 (N_14529,N_12534,N_12979);
xnor U14530 (N_14530,N_12993,N_12115);
and U14531 (N_14531,N_13109,N_13390);
nand U14532 (N_14532,N_12844,N_12945);
nor U14533 (N_14533,N_12766,N_12552);
or U14534 (N_14534,N_12136,N_13445);
nor U14535 (N_14535,N_13009,N_13344);
nand U14536 (N_14536,N_13104,N_12736);
and U14537 (N_14537,N_12828,N_13015);
and U14538 (N_14538,N_12521,N_13400);
and U14539 (N_14539,N_13445,N_12510);
or U14540 (N_14540,N_13403,N_12153);
nand U14541 (N_14541,N_12897,N_12102);
or U14542 (N_14542,N_13051,N_12682);
and U14543 (N_14543,N_13396,N_12588);
or U14544 (N_14544,N_13070,N_12008);
nand U14545 (N_14545,N_13296,N_13468);
nor U14546 (N_14546,N_12756,N_12404);
and U14547 (N_14547,N_12607,N_12817);
or U14548 (N_14548,N_13103,N_12741);
or U14549 (N_14549,N_13318,N_12846);
nand U14550 (N_14550,N_12223,N_12495);
nand U14551 (N_14551,N_12335,N_13387);
nor U14552 (N_14552,N_13363,N_13206);
nor U14553 (N_14553,N_12009,N_12153);
or U14554 (N_14554,N_12076,N_12486);
or U14555 (N_14555,N_12388,N_12480);
or U14556 (N_14556,N_13030,N_13064);
or U14557 (N_14557,N_13063,N_12286);
and U14558 (N_14558,N_13104,N_12878);
and U14559 (N_14559,N_13349,N_13427);
and U14560 (N_14560,N_13243,N_12857);
and U14561 (N_14561,N_12274,N_13264);
nor U14562 (N_14562,N_12295,N_13138);
and U14563 (N_14563,N_12574,N_12495);
and U14564 (N_14564,N_12681,N_13288);
and U14565 (N_14565,N_12000,N_13105);
and U14566 (N_14566,N_12976,N_12375);
and U14567 (N_14567,N_12205,N_13008);
nor U14568 (N_14568,N_12780,N_12822);
nor U14569 (N_14569,N_12701,N_13051);
and U14570 (N_14570,N_12508,N_13231);
nand U14571 (N_14571,N_13240,N_12398);
nor U14572 (N_14572,N_12451,N_12398);
nor U14573 (N_14573,N_12650,N_12916);
nand U14574 (N_14574,N_12611,N_13493);
nand U14575 (N_14575,N_12118,N_12438);
nand U14576 (N_14576,N_12012,N_12905);
nor U14577 (N_14577,N_12739,N_12142);
or U14578 (N_14578,N_13227,N_12439);
nor U14579 (N_14579,N_13288,N_13198);
nor U14580 (N_14580,N_12204,N_12623);
nand U14581 (N_14581,N_12292,N_13307);
and U14582 (N_14582,N_12019,N_12847);
nand U14583 (N_14583,N_13211,N_13227);
nor U14584 (N_14584,N_13297,N_13315);
nor U14585 (N_14585,N_13290,N_13228);
and U14586 (N_14586,N_12594,N_13392);
or U14587 (N_14587,N_13215,N_12252);
nand U14588 (N_14588,N_12075,N_12988);
nor U14589 (N_14589,N_13286,N_12777);
nand U14590 (N_14590,N_12561,N_12555);
and U14591 (N_14591,N_13459,N_12794);
nor U14592 (N_14592,N_13164,N_12420);
or U14593 (N_14593,N_12309,N_13152);
or U14594 (N_14594,N_12631,N_12310);
xnor U14595 (N_14595,N_13137,N_13479);
nand U14596 (N_14596,N_12662,N_12514);
nor U14597 (N_14597,N_12720,N_12556);
or U14598 (N_14598,N_13112,N_13180);
or U14599 (N_14599,N_12991,N_12773);
and U14600 (N_14600,N_12942,N_12441);
xnor U14601 (N_14601,N_12404,N_13243);
nor U14602 (N_14602,N_12752,N_13049);
and U14603 (N_14603,N_12794,N_13210);
nor U14604 (N_14604,N_13202,N_13406);
nand U14605 (N_14605,N_12729,N_12557);
and U14606 (N_14606,N_12148,N_13343);
nand U14607 (N_14607,N_13427,N_13178);
or U14608 (N_14608,N_12888,N_12280);
or U14609 (N_14609,N_13471,N_12196);
or U14610 (N_14610,N_12684,N_13144);
nor U14611 (N_14611,N_12570,N_12825);
nor U14612 (N_14612,N_12121,N_12475);
or U14613 (N_14613,N_12182,N_13366);
or U14614 (N_14614,N_12198,N_12287);
nand U14615 (N_14615,N_13201,N_12743);
and U14616 (N_14616,N_12498,N_13418);
and U14617 (N_14617,N_12337,N_12920);
xor U14618 (N_14618,N_12256,N_13377);
nand U14619 (N_14619,N_13027,N_13102);
nor U14620 (N_14620,N_12097,N_12670);
or U14621 (N_14621,N_13068,N_12114);
and U14622 (N_14622,N_13391,N_12455);
nor U14623 (N_14623,N_12360,N_12104);
nor U14624 (N_14624,N_13422,N_12464);
nor U14625 (N_14625,N_13430,N_13008);
or U14626 (N_14626,N_12764,N_13474);
nor U14627 (N_14627,N_12860,N_12688);
nand U14628 (N_14628,N_12581,N_12719);
xor U14629 (N_14629,N_12011,N_12670);
or U14630 (N_14630,N_12851,N_12192);
and U14631 (N_14631,N_12811,N_13407);
or U14632 (N_14632,N_13010,N_12970);
nor U14633 (N_14633,N_12426,N_12206);
nand U14634 (N_14634,N_12390,N_12540);
and U14635 (N_14635,N_13353,N_12410);
nor U14636 (N_14636,N_13136,N_12130);
nand U14637 (N_14637,N_13388,N_13002);
nor U14638 (N_14638,N_13393,N_12818);
nand U14639 (N_14639,N_12695,N_12504);
or U14640 (N_14640,N_12048,N_13372);
or U14641 (N_14641,N_12564,N_12874);
and U14642 (N_14642,N_13339,N_12233);
nand U14643 (N_14643,N_13433,N_12771);
nand U14644 (N_14644,N_12573,N_12787);
nand U14645 (N_14645,N_12756,N_12998);
nor U14646 (N_14646,N_12914,N_13314);
nor U14647 (N_14647,N_12028,N_13408);
nand U14648 (N_14648,N_12916,N_13417);
or U14649 (N_14649,N_12679,N_13161);
nor U14650 (N_14650,N_13491,N_13222);
nand U14651 (N_14651,N_13434,N_13327);
or U14652 (N_14652,N_12361,N_12958);
or U14653 (N_14653,N_13059,N_12756);
nand U14654 (N_14654,N_12691,N_12794);
nor U14655 (N_14655,N_12266,N_12581);
nor U14656 (N_14656,N_13311,N_13177);
nor U14657 (N_14657,N_12001,N_13274);
nor U14658 (N_14658,N_12117,N_13209);
nand U14659 (N_14659,N_12724,N_12585);
nor U14660 (N_14660,N_12475,N_13341);
or U14661 (N_14661,N_12941,N_13209);
and U14662 (N_14662,N_12716,N_12031);
or U14663 (N_14663,N_12130,N_13130);
nand U14664 (N_14664,N_12092,N_12425);
or U14665 (N_14665,N_12758,N_12727);
or U14666 (N_14666,N_12689,N_13089);
and U14667 (N_14667,N_13249,N_12883);
nand U14668 (N_14668,N_13255,N_13320);
or U14669 (N_14669,N_13481,N_12626);
nand U14670 (N_14670,N_13121,N_13258);
or U14671 (N_14671,N_12293,N_12486);
and U14672 (N_14672,N_13138,N_12134);
nand U14673 (N_14673,N_12070,N_12988);
and U14674 (N_14674,N_12032,N_12487);
nand U14675 (N_14675,N_12127,N_13305);
and U14676 (N_14676,N_13422,N_12335);
nor U14677 (N_14677,N_13289,N_13372);
nand U14678 (N_14678,N_13349,N_13063);
and U14679 (N_14679,N_12190,N_13231);
nand U14680 (N_14680,N_12519,N_13040);
or U14681 (N_14681,N_12114,N_12376);
and U14682 (N_14682,N_13347,N_13478);
nand U14683 (N_14683,N_13166,N_12137);
and U14684 (N_14684,N_12619,N_12163);
nor U14685 (N_14685,N_12986,N_12904);
nand U14686 (N_14686,N_12266,N_12729);
nor U14687 (N_14687,N_12800,N_13146);
nor U14688 (N_14688,N_13271,N_12601);
and U14689 (N_14689,N_12187,N_12464);
nand U14690 (N_14690,N_12074,N_13354);
nor U14691 (N_14691,N_12318,N_13118);
nand U14692 (N_14692,N_12756,N_13169);
nand U14693 (N_14693,N_12044,N_13245);
nand U14694 (N_14694,N_12619,N_13453);
nor U14695 (N_14695,N_12124,N_13156);
nor U14696 (N_14696,N_12089,N_13370);
xor U14697 (N_14697,N_12082,N_12928);
and U14698 (N_14698,N_12735,N_12902);
or U14699 (N_14699,N_13078,N_12906);
and U14700 (N_14700,N_12546,N_12263);
nand U14701 (N_14701,N_13099,N_13122);
nand U14702 (N_14702,N_12089,N_12581);
nor U14703 (N_14703,N_12496,N_12570);
or U14704 (N_14704,N_12825,N_13232);
and U14705 (N_14705,N_12528,N_12853);
and U14706 (N_14706,N_12513,N_12453);
nor U14707 (N_14707,N_13302,N_12765);
nand U14708 (N_14708,N_12773,N_12587);
xor U14709 (N_14709,N_12531,N_12909);
nand U14710 (N_14710,N_13176,N_12374);
or U14711 (N_14711,N_12875,N_13212);
and U14712 (N_14712,N_12189,N_12416);
or U14713 (N_14713,N_12170,N_13219);
nor U14714 (N_14714,N_12941,N_13244);
or U14715 (N_14715,N_13149,N_13276);
nand U14716 (N_14716,N_13191,N_13061);
nor U14717 (N_14717,N_12419,N_13071);
xnor U14718 (N_14718,N_12377,N_12765);
nand U14719 (N_14719,N_12540,N_12276);
nor U14720 (N_14720,N_12550,N_13359);
nand U14721 (N_14721,N_12651,N_12410);
or U14722 (N_14722,N_12136,N_12085);
or U14723 (N_14723,N_12453,N_12471);
nand U14724 (N_14724,N_13188,N_12470);
nor U14725 (N_14725,N_12186,N_13239);
nor U14726 (N_14726,N_12167,N_12611);
nor U14727 (N_14727,N_13392,N_12958);
and U14728 (N_14728,N_13074,N_12304);
nor U14729 (N_14729,N_12849,N_13430);
or U14730 (N_14730,N_13474,N_12446);
nand U14731 (N_14731,N_13160,N_13320);
xnor U14732 (N_14732,N_12762,N_12708);
or U14733 (N_14733,N_13102,N_13127);
or U14734 (N_14734,N_12989,N_13102);
or U14735 (N_14735,N_13473,N_12092);
xor U14736 (N_14736,N_12136,N_13156);
and U14737 (N_14737,N_12596,N_13114);
nand U14738 (N_14738,N_13031,N_12974);
and U14739 (N_14739,N_12084,N_12938);
and U14740 (N_14740,N_13439,N_13468);
nor U14741 (N_14741,N_12639,N_12396);
nand U14742 (N_14742,N_13005,N_13475);
nand U14743 (N_14743,N_13478,N_12331);
nand U14744 (N_14744,N_13356,N_13321);
or U14745 (N_14745,N_12382,N_12797);
xor U14746 (N_14746,N_12757,N_13308);
and U14747 (N_14747,N_12414,N_13162);
and U14748 (N_14748,N_12767,N_12977);
nor U14749 (N_14749,N_13036,N_13053);
or U14750 (N_14750,N_12589,N_12794);
nand U14751 (N_14751,N_12304,N_12543);
nand U14752 (N_14752,N_12324,N_13124);
nand U14753 (N_14753,N_12653,N_12088);
and U14754 (N_14754,N_13476,N_12157);
or U14755 (N_14755,N_12933,N_13225);
or U14756 (N_14756,N_12238,N_12578);
and U14757 (N_14757,N_13476,N_12059);
nand U14758 (N_14758,N_12397,N_12199);
or U14759 (N_14759,N_12827,N_12662);
nand U14760 (N_14760,N_12917,N_12669);
and U14761 (N_14761,N_12709,N_12316);
nand U14762 (N_14762,N_12606,N_12359);
and U14763 (N_14763,N_13175,N_12492);
nand U14764 (N_14764,N_12358,N_12872);
nor U14765 (N_14765,N_12742,N_13399);
and U14766 (N_14766,N_12851,N_13338);
or U14767 (N_14767,N_12778,N_13020);
and U14768 (N_14768,N_13359,N_12492);
nor U14769 (N_14769,N_13134,N_12980);
nand U14770 (N_14770,N_13369,N_12257);
nand U14771 (N_14771,N_12566,N_12176);
nand U14772 (N_14772,N_12444,N_13319);
and U14773 (N_14773,N_12281,N_12184);
nand U14774 (N_14774,N_12984,N_13274);
nor U14775 (N_14775,N_13145,N_12182);
nand U14776 (N_14776,N_13127,N_12798);
or U14777 (N_14777,N_13288,N_13211);
and U14778 (N_14778,N_13373,N_12420);
or U14779 (N_14779,N_12322,N_13421);
or U14780 (N_14780,N_13209,N_12247);
or U14781 (N_14781,N_12502,N_13233);
nand U14782 (N_14782,N_12757,N_12154);
nand U14783 (N_14783,N_12714,N_12568);
and U14784 (N_14784,N_12191,N_12604);
and U14785 (N_14785,N_12322,N_13065);
nand U14786 (N_14786,N_12537,N_12851);
or U14787 (N_14787,N_12454,N_13111);
and U14788 (N_14788,N_12585,N_12792);
or U14789 (N_14789,N_13368,N_12166);
nand U14790 (N_14790,N_12022,N_12246);
nor U14791 (N_14791,N_12023,N_12482);
and U14792 (N_14792,N_12547,N_12969);
nand U14793 (N_14793,N_12878,N_13463);
nor U14794 (N_14794,N_13104,N_12954);
and U14795 (N_14795,N_13308,N_12551);
nor U14796 (N_14796,N_12932,N_12064);
or U14797 (N_14797,N_13463,N_12125);
nand U14798 (N_14798,N_12085,N_12434);
nor U14799 (N_14799,N_12766,N_12194);
or U14800 (N_14800,N_12947,N_12443);
nor U14801 (N_14801,N_12440,N_12727);
or U14802 (N_14802,N_12774,N_12312);
or U14803 (N_14803,N_12152,N_13346);
or U14804 (N_14804,N_12799,N_12948);
xor U14805 (N_14805,N_13221,N_12728);
and U14806 (N_14806,N_12377,N_12777);
or U14807 (N_14807,N_12140,N_12700);
nor U14808 (N_14808,N_12203,N_12209);
nand U14809 (N_14809,N_12937,N_12243);
and U14810 (N_14810,N_12985,N_12607);
or U14811 (N_14811,N_13353,N_12108);
nand U14812 (N_14812,N_12509,N_12666);
and U14813 (N_14813,N_12606,N_13309);
and U14814 (N_14814,N_13238,N_12508);
and U14815 (N_14815,N_13364,N_12526);
and U14816 (N_14816,N_12290,N_13283);
nor U14817 (N_14817,N_12509,N_12685);
or U14818 (N_14818,N_13155,N_12941);
nand U14819 (N_14819,N_13188,N_13413);
and U14820 (N_14820,N_12776,N_12234);
nor U14821 (N_14821,N_12313,N_12524);
nand U14822 (N_14822,N_12786,N_12665);
and U14823 (N_14823,N_13135,N_12284);
or U14824 (N_14824,N_12478,N_13025);
and U14825 (N_14825,N_13399,N_13485);
or U14826 (N_14826,N_13485,N_13266);
nand U14827 (N_14827,N_12031,N_12238);
or U14828 (N_14828,N_12961,N_13032);
or U14829 (N_14829,N_13454,N_13480);
nor U14830 (N_14830,N_12094,N_12953);
or U14831 (N_14831,N_12377,N_12956);
and U14832 (N_14832,N_13253,N_12749);
nor U14833 (N_14833,N_12618,N_13021);
nand U14834 (N_14834,N_12882,N_12339);
and U14835 (N_14835,N_12015,N_12437);
nor U14836 (N_14836,N_12623,N_13101);
nand U14837 (N_14837,N_13192,N_12801);
nand U14838 (N_14838,N_12049,N_12318);
nor U14839 (N_14839,N_13286,N_13426);
xor U14840 (N_14840,N_13294,N_12712);
nand U14841 (N_14841,N_13112,N_12624);
nor U14842 (N_14842,N_12823,N_12491);
nor U14843 (N_14843,N_12126,N_13351);
nor U14844 (N_14844,N_12864,N_12701);
and U14845 (N_14845,N_12265,N_13174);
nand U14846 (N_14846,N_13023,N_13312);
or U14847 (N_14847,N_12056,N_13006);
and U14848 (N_14848,N_12639,N_13474);
nor U14849 (N_14849,N_12199,N_13008);
nor U14850 (N_14850,N_12320,N_13400);
or U14851 (N_14851,N_13152,N_12040);
nor U14852 (N_14852,N_12999,N_12835);
nand U14853 (N_14853,N_13280,N_13043);
and U14854 (N_14854,N_12986,N_12801);
nor U14855 (N_14855,N_12297,N_13221);
nand U14856 (N_14856,N_13344,N_12201);
or U14857 (N_14857,N_12716,N_12838);
and U14858 (N_14858,N_13030,N_12676);
xnor U14859 (N_14859,N_12325,N_12989);
nor U14860 (N_14860,N_12987,N_13007);
nand U14861 (N_14861,N_12246,N_12593);
nand U14862 (N_14862,N_12036,N_13231);
and U14863 (N_14863,N_13096,N_12493);
or U14864 (N_14864,N_12429,N_13416);
nor U14865 (N_14865,N_12340,N_12405);
nand U14866 (N_14866,N_12286,N_13139);
nor U14867 (N_14867,N_12108,N_13311);
and U14868 (N_14868,N_12229,N_12997);
nand U14869 (N_14869,N_12312,N_12293);
or U14870 (N_14870,N_13378,N_13246);
nor U14871 (N_14871,N_13189,N_13140);
nand U14872 (N_14872,N_12488,N_13132);
nor U14873 (N_14873,N_13167,N_12462);
or U14874 (N_14874,N_12899,N_13003);
and U14875 (N_14875,N_12628,N_12020);
nand U14876 (N_14876,N_12743,N_12580);
or U14877 (N_14877,N_13168,N_12198);
nor U14878 (N_14878,N_12742,N_12810);
nor U14879 (N_14879,N_13236,N_12859);
or U14880 (N_14880,N_13007,N_13328);
nor U14881 (N_14881,N_12440,N_12805);
and U14882 (N_14882,N_13105,N_12980);
or U14883 (N_14883,N_12112,N_13334);
nand U14884 (N_14884,N_13375,N_12065);
nor U14885 (N_14885,N_12296,N_13160);
and U14886 (N_14886,N_12719,N_12301);
or U14887 (N_14887,N_12272,N_13417);
xnor U14888 (N_14888,N_12480,N_13002);
nand U14889 (N_14889,N_13422,N_12680);
and U14890 (N_14890,N_13440,N_13475);
nand U14891 (N_14891,N_12172,N_12237);
nand U14892 (N_14892,N_12651,N_13486);
nand U14893 (N_14893,N_12838,N_12905);
and U14894 (N_14894,N_12482,N_12451);
or U14895 (N_14895,N_13463,N_12943);
nor U14896 (N_14896,N_12939,N_12493);
or U14897 (N_14897,N_12490,N_12310);
and U14898 (N_14898,N_12955,N_13161);
nor U14899 (N_14899,N_13453,N_13256);
or U14900 (N_14900,N_12242,N_12179);
nand U14901 (N_14901,N_12191,N_12714);
xor U14902 (N_14902,N_13125,N_12442);
and U14903 (N_14903,N_12720,N_12565);
nor U14904 (N_14904,N_13149,N_13176);
nand U14905 (N_14905,N_13257,N_13301);
or U14906 (N_14906,N_12302,N_13299);
nand U14907 (N_14907,N_12886,N_12963);
or U14908 (N_14908,N_13280,N_12468);
and U14909 (N_14909,N_12634,N_12921);
and U14910 (N_14910,N_13327,N_12742);
and U14911 (N_14911,N_12644,N_12982);
nor U14912 (N_14912,N_13479,N_12739);
and U14913 (N_14913,N_13277,N_12671);
nand U14914 (N_14914,N_12271,N_12877);
and U14915 (N_14915,N_12476,N_12319);
and U14916 (N_14916,N_13092,N_12739);
or U14917 (N_14917,N_12700,N_13075);
nand U14918 (N_14918,N_12492,N_13035);
nor U14919 (N_14919,N_12153,N_12989);
nor U14920 (N_14920,N_12652,N_13179);
and U14921 (N_14921,N_12657,N_12797);
or U14922 (N_14922,N_13082,N_13114);
nor U14923 (N_14923,N_13221,N_13068);
nand U14924 (N_14924,N_12273,N_13179);
nand U14925 (N_14925,N_12571,N_12451);
and U14926 (N_14926,N_12347,N_12647);
nor U14927 (N_14927,N_13421,N_13080);
xnor U14928 (N_14928,N_12558,N_13220);
nor U14929 (N_14929,N_13453,N_12477);
nand U14930 (N_14930,N_13465,N_13348);
and U14931 (N_14931,N_13478,N_12383);
or U14932 (N_14932,N_12095,N_12700);
or U14933 (N_14933,N_12343,N_12028);
or U14934 (N_14934,N_13137,N_13336);
nand U14935 (N_14935,N_12693,N_12998);
or U14936 (N_14936,N_12765,N_13252);
nor U14937 (N_14937,N_12295,N_12828);
or U14938 (N_14938,N_13116,N_12056);
and U14939 (N_14939,N_12610,N_12693);
or U14940 (N_14940,N_12840,N_12756);
nand U14941 (N_14941,N_13184,N_12361);
and U14942 (N_14942,N_12586,N_13422);
nand U14943 (N_14943,N_13253,N_12609);
or U14944 (N_14944,N_13457,N_12912);
nand U14945 (N_14945,N_13471,N_13026);
nand U14946 (N_14946,N_12957,N_13181);
nor U14947 (N_14947,N_12708,N_12497);
nor U14948 (N_14948,N_13020,N_12139);
and U14949 (N_14949,N_13445,N_12975);
nor U14950 (N_14950,N_12339,N_12773);
nand U14951 (N_14951,N_13072,N_12086);
xor U14952 (N_14952,N_12310,N_13467);
nand U14953 (N_14953,N_12269,N_12478);
nand U14954 (N_14954,N_12692,N_13309);
nor U14955 (N_14955,N_12984,N_12312);
and U14956 (N_14956,N_12851,N_12105);
nor U14957 (N_14957,N_12618,N_12269);
nand U14958 (N_14958,N_13129,N_12038);
xor U14959 (N_14959,N_12465,N_12515);
nor U14960 (N_14960,N_13384,N_12415);
nand U14961 (N_14961,N_13471,N_13496);
nand U14962 (N_14962,N_13463,N_12678);
nor U14963 (N_14963,N_13385,N_13233);
nor U14964 (N_14964,N_12702,N_12368);
or U14965 (N_14965,N_12844,N_13256);
or U14966 (N_14966,N_13291,N_12695);
and U14967 (N_14967,N_12704,N_12197);
or U14968 (N_14968,N_13242,N_12164);
xnor U14969 (N_14969,N_12220,N_13459);
nor U14970 (N_14970,N_12051,N_13281);
nor U14971 (N_14971,N_12446,N_13460);
and U14972 (N_14972,N_12974,N_12200);
nand U14973 (N_14973,N_12879,N_13207);
or U14974 (N_14974,N_12975,N_12633);
and U14975 (N_14975,N_12196,N_12975);
nand U14976 (N_14976,N_12165,N_12434);
nand U14977 (N_14977,N_12015,N_12728);
or U14978 (N_14978,N_13039,N_12602);
or U14979 (N_14979,N_12701,N_12420);
and U14980 (N_14980,N_12376,N_13237);
nand U14981 (N_14981,N_13283,N_13432);
nor U14982 (N_14982,N_12798,N_12975);
or U14983 (N_14983,N_13201,N_12032);
nor U14984 (N_14984,N_12441,N_13004);
nand U14985 (N_14985,N_13078,N_13474);
or U14986 (N_14986,N_12554,N_13250);
nand U14987 (N_14987,N_12428,N_12658);
nor U14988 (N_14988,N_12983,N_13344);
or U14989 (N_14989,N_12450,N_12997);
nor U14990 (N_14990,N_13197,N_12737);
or U14991 (N_14991,N_12560,N_13402);
and U14992 (N_14992,N_13416,N_12605);
nor U14993 (N_14993,N_12874,N_13324);
nand U14994 (N_14994,N_12664,N_12155);
nor U14995 (N_14995,N_12016,N_13332);
and U14996 (N_14996,N_12696,N_12959);
and U14997 (N_14997,N_13357,N_12734);
or U14998 (N_14998,N_12895,N_12784);
and U14999 (N_14999,N_12755,N_12863);
or UO_0 (O_0,N_14234,N_14023);
and UO_1 (O_1,N_14152,N_14143);
nor UO_2 (O_2,N_13793,N_13655);
nor UO_3 (O_3,N_13577,N_14840);
or UO_4 (O_4,N_14775,N_14517);
or UO_5 (O_5,N_14322,N_13689);
nor UO_6 (O_6,N_14557,N_14319);
nand UO_7 (O_7,N_14961,N_14656);
nor UO_8 (O_8,N_13613,N_14107);
or UO_9 (O_9,N_13637,N_13628);
and UO_10 (O_10,N_13982,N_14001);
nor UO_11 (O_11,N_14649,N_14536);
nor UO_12 (O_12,N_13684,N_14175);
or UO_13 (O_13,N_14219,N_14617);
xor UO_14 (O_14,N_13798,N_13851);
nand UO_15 (O_15,N_13873,N_14077);
nor UO_16 (O_16,N_13857,N_14194);
and UO_17 (O_17,N_14661,N_14991);
and UO_18 (O_18,N_13783,N_14804);
nand UO_19 (O_19,N_14109,N_14177);
or UO_20 (O_20,N_14423,N_13975);
and UO_21 (O_21,N_14270,N_13937);
nand UO_22 (O_22,N_14696,N_14101);
nor UO_23 (O_23,N_14193,N_13532);
and UO_24 (O_24,N_13676,N_13965);
nor UO_25 (O_25,N_13558,N_14806);
and UO_26 (O_26,N_14344,N_14292);
nor UO_27 (O_27,N_14660,N_13971);
or UO_28 (O_28,N_14154,N_14890);
and UO_29 (O_29,N_13680,N_14508);
nand UO_30 (O_30,N_13911,N_14261);
and UO_31 (O_31,N_14805,N_14797);
and UO_32 (O_32,N_13967,N_13622);
or UO_33 (O_33,N_14839,N_14418);
xor UO_34 (O_34,N_14711,N_13731);
nor UO_35 (O_35,N_14156,N_14987);
and UO_36 (O_36,N_14305,N_13862);
or UO_37 (O_37,N_13932,N_13512);
nand UO_38 (O_38,N_14010,N_14549);
nor UO_39 (O_39,N_13756,N_14054);
nor UO_40 (O_40,N_13675,N_13682);
nand UO_41 (O_41,N_14932,N_13725);
or UO_42 (O_42,N_13521,N_13536);
nand UO_43 (O_43,N_14600,N_14184);
and UO_44 (O_44,N_14727,N_14901);
xnor UO_45 (O_45,N_14180,N_14581);
nor UO_46 (O_46,N_13698,N_13782);
nand UO_47 (O_47,N_14044,N_13534);
and UO_48 (O_48,N_13823,N_13730);
or UO_49 (O_49,N_14674,N_14560);
nor UO_50 (O_50,N_14274,N_14915);
nor UO_51 (O_51,N_14845,N_13503);
nor UO_52 (O_52,N_14922,N_13580);
or UO_53 (O_53,N_14835,N_14918);
or UO_54 (O_54,N_14823,N_14051);
xor UO_55 (O_55,N_14208,N_13507);
or UO_56 (O_56,N_14937,N_14090);
or UO_57 (O_57,N_14684,N_14138);
and UO_58 (O_58,N_14430,N_13891);
or UO_59 (O_59,N_14119,N_14225);
nand UO_60 (O_60,N_14999,N_14377);
and UO_61 (O_61,N_14167,N_13661);
nand UO_62 (O_62,N_14034,N_13753);
nand UO_63 (O_63,N_13742,N_14139);
or UO_64 (O_64,N_14800,N_13677);
and UO_65 (O_65,N_13665,N_14682);
or UO_66 (O_66,N_14009,N_14692);
or UO_67 (O_67,N_14783,N_14040);
nor UO_68 (O_68,N_13673,N_14151);
nor UO_69 (O_69,N_14820,N_13739);
or UO_70 (O_70,N_14356,N_14616);
and UO_71 (O_71,N_14221,N_14264);
and UO_72 (O_72,N_14770,N_14112);
or UO_73 (O_73,N_14345,N_13687);
nor UO_74 (O_74,N_14150,N_14378);
nor UO_75 (O_75,N_13870,N_14832);
nand UO_76 (O_76,N_13625,N_13566);
nand UO_77 (O_77,N_13883,N_14092);
nand UO_78 (O_78,N_13979,N_13543);
nor UO_79 (O_79,N_14907,N_14947);
nor UO_80 (O_80,N_14240,N_13992);
nor UO_81 (O_81,N_13683,N_14764);
nand UO_82 (O_82,N_14768,N_14538);
nand UO_83 (O_83,N_14332,N_13942);
or UO_84 (O_84,N_13912,N_14945);
or UO_85 (O_85,N_13797,N_14850);
nor UO_86 (O_86,N_13704,N_13824);
nand UO_87 (O_87,N_13618,N_14621);
and UO_88 (O_88,N_14246,N_14210);
nor UO_89 (O_89,N_14665,N_13542);
nand UO_90 (O_90,N_14756,N_14115);
xnor UO_91 (O_91,N_14397,N_14329);
and UO_92 (O_92,N_14169,N_14041);
or UO_93 (O_93,N_14304,N_14867);
or UO_94 (O_94,N_13907,N_14633);
or UO_95 (O_95,N_13744,N_14203);
and UO_96 (O_96,N_14336,N_14342);
nand UO_97 (O_97,N_14120,N_14160);
and UO_98 (O_98,N_14148,N_13959);
nor UO_99 (O_99,N_14874,N_14761);
and UO_100 (O_100,N_14752,N_14352);
and UO_101 (O_101,N_14091,N_13761);
or UO_102 (O_102,N_14291,N_13821);
or UO_103 (O_103,N_13808,N_14364);
and UO_104 (O_104,N_14545,N_14725);
nand UO_105 (O_105,N_14447,N_14944);
and UO_106 (O_106,N_14958,N_14035);
and UO_107 (O_107,N_14533,N_13884);
and UO_108 (O_108,N_14006,N_13656);
and UO_109 (O_109,N_14708,N_14626);
xor UO_110 (O_110,N_14494,N_14717);
or UO_111 (O_111,N_13970,N_14811);
xor UO_112 (O_112,N_13961,N_13602);
or UO_113 (O_113,N_14639,N_14460);
and UO_114 (O_114,N_14644,N_14459);
nand UO_115 (O_115,N_14401,N_13644);
or UO_116 (O_116,N_14297,N_13593);
nor UO_117 (O_117,N_14609,N_14173);
or UO_118 (O_118,N_14384,N_14927);
nor UO_119 (O_119,N_13733,N_14189);
nor UO_120 (O_120,N_13509,N_13991);
xnor UO_121 (O_121,N_14877,N_14339);
and UO_122 (O_122,N_14451,N_13526);
nor UO_123 (O_123,N_14855,N_14940);
and UO_124 (O_124,N_13928,N_14912);
nand UO_125 (O_125,N_13658,N_14552);
or UO_126 (O_126,N_14628,N_14746);
nor UO_127 (O_127,N_13583,N_14469);
nor UO_128 (O_128,N_13943,N_13719);
and UO_129 (O_129,N_14849,N_13803);
or UO_130 (O_130,N_13524,N_14525);
xor UO_131 (O_131,N_14742,N_14938);
or UO_132 (O_132,N_14170,N_14348);
or UO_133 (O_133,N_14518,N_14452);
nand UO_134 (O_134,N_14697,N_13667);
and UO_135 (O_135,N_14934,N_14577);
nor UO_136 (O_136,N_14614,N_13574);
nor UO_137 (O_137,N_14580,N_13799);
nand UO_138 (O_138,N_14710,N_13551);
nor UO_139 (O_139,N_14798,N_14094);
nor UO_140 (O_140,N_13832,N_13576);
nor UO_141 (O_141,N_14427,N_14529);
and UO_142 (O_142,N_13941,N_14970);
or UO_143 (O_143,N_13904,N_13887);
nor UO_144 (O_144,N_14343,N_14540);
and UO_145 (O_145,N_14648,N_14908);
nor UO_146 (O_146,N_14429,N_14113);
xor UO_147 (O_147,N_14905,N_13650);
or UO_148 (O_148,N_14371,N_13915);
nor UO_149 (O_149,N_13867,N_14137);
nor UO_150 (O_150,N_14439,N_14728);
nor UO_151 (O_151,N_13629,N_14869);
and UO_152 (O_152,N_14142,N_13838);
nand UO_153 (O_153,N_14997,N_13517);
and UO_154 (O_154,N_14956,N_14438);
or UO_155 (O_155,N_14388,N_14285);
nand UO_156 (O_156,N_14584,N_13984);
and UO_157 (O_157,N_14543,N_14192);
nor UO_158 (O_158,N_14871,N_14293);
and UO_159 (O_159,N_14755,N_13736);
nand UO_160 (O_160,N_13699,N_13903);
xor UO_161 (O_161,N_14885,N_13901);
or UO_162 (O_162,N_14968,N_13585);
nand UO_163 (O_163,N_14515,N_14008);
nor UO_164 (O_164,N_14812,N_14394);
or UO_165 (O_165,N_14807,N_13711);
and UO_166 (O_166,N_14050,N_13728);
and UO_167 (O_167,N_13801,N_13788);
or UO_168 (O_168,N_13819,N_14262);
nor UO_169 (O_169,N_13952,N_14951);
nor UO_170 (O_170,N_14049,N_14353);
or UO_171 (O_171,N_14444,N_14759);
xnor UO_172 (O_172,N_14410,N_13679);
nor UO_173 (O_173,N_14045,N_14414);
nor UO_174 (O_174,N_13945,N_13501);
and UO_175 (O_175,N_13589,N_14878);
nor UO_176 (O_176,N_13694,N_14317);
or UO_177 (O_177,N_13708,N_14534);
and UO_178 (O_178,N_13748,N_14174);
and UO_179 (O_179,N_14506,N_14406);
and UO_180 (O_180,N_13817,N_14131);
and UO_181 (O_181,N_13999,N_13726);
nor UO_182 (O_182,N_14870,N_13648);
nand UO_183 (O_183,N_14232,N_14749);
or UO_184 (O_184,N_13770,N_14176);
and UO_185 (O_185,N_14729,N_13621);
nor UO_186 (O_186,N_13834,N_14233);
and UO_187 (O_187,N_14791,N_14200);
or UO_188 (O_188,N_13889,N_13617);
nand UO_189 (O_189,N_13606,N_14016);
and UO_190 (O_190,N_13842,N_14315);
or UO_191 (O_191,N_14326,N_14732);
nand UO_192 (O_192,N_13712,N_14790);
nor UO_193 (O_193,N_13569,N_14488);
nor UO_194 (O_194,N_13789,N_14673);
or UO_195 (O_195,N_13519,N_14687);
nand UO_196 (O_196,N_14634,N_14312);
nor UO_197 (O_197,N_14663,N_14162);
or UO_198 (O_198,N_14472,N_14522);
nand UO_199 (O_199,N_13518,N_14570);
nand UO_200 (O_200,N_13765,N_13876);
or UO_201 (O_201,N_14069,N_13856);
or UO_202 (O_202,N_13640,N_14498);
nand UO_203 (O_203,N_14658,N_14409);
and UO_204 (O_204,N_13923,N_13595);
or UO_205 (O_205,N_14482,N_14379);
or UO_206 (O_206,N_14149,N_14751);
nor UO_207 (O_207,N_13780,N_14786);
nor UO_208 (O_208,N_14572,N_13769);
or UO_209 (O_209,N_13531,N_14255);
and UO_210 (O_210,N_13854,N_14209);
and UO_211 (O_211,N_14782,N_14726);
nor UO_212 (O_212,N_14926,N_14579);
and UO_213 (O_213,N_14501,N_13987);
nor UO_214 (O_214,N_14520,N_14398);
nand UO_215 (O_215,N_13603,N_13953);
and UO_216 (O_216,N_13914,N_14833);
nor UO_217 (O_217,N_13816,N_14039);
or UO_218 (O_218,N_14052,N_14257);
nor UO_219 (O_219,N_13643,N_13946);
nor UO_220 (O_220,N_14046,N_14712);
nand UO_221 (O_221,N_13894,N_14033);
and UO_222 (O_222,N_14910,N_13985);
or UO_223 (O_223,N_13792,N_14979);
and UO_224 (O_224,N_14743,N_13590);
nand UO_225 (O_225,N_14415,N_14450);
and UO_226 (O_226,N_14181,N_13795);
nand UO_227 (O_227,N_14683,N_14117);
and UO_228 (O_228,N_14873,N_14638);
or UO_229 (O_229,N_13897,N_14417);
nand UO_230 (O_230,N_14484,N_14948);
and UO_231 (O_231,N_14844,N_14294);
or UO_232 (O_232,N_14590,N_14349);
or UO_233 (O_233,N_14290,N_14437);
nor UO_234 (O_234,N_14239,N_14164);
nand UO_235 (O_235,N_14277,N_13802);
nand UO_236 (O_236,N_13768,N_14686);
and UO_237 (O_237,N_13693,N_13554);
or UO_238 (O_238,N_14188,N_14813);
nand UO_239 (O_239,N_14300,N_14369);
nor UO_240 (O_240,N_14029,N_13721);
or UO_241 (O_241,N_14282,N_13747);
xor UO_242 (O_242,N_14578,N_14363);
and UO_243 (O_243,N_13840,N_14510);
and UO_244 (O_244,N_14493,N_13701);
or UO_245 (O_245,N_13905,N_14923);
and UO_246 (O_246,N_13813,N_14445);
xnor UO_247 (O_247,N_14618,N_13892);
nor UO_248 (O_248,N_14598,N_14168);
or UO_249 (O_249,N_14256,N_14335);
or UO_250 (O_250,N_14036,N_14599);
nor UO_251 (O_251,N_14942,N_13604);
nand UO_252 (O_252,N_14731,N_14744);
and UO_253 (O_253,N_14896,N_14042);
and UO_254 (O_254,N_13716,N_13565);
nor UO_255 (O_255,N_14230,N_14691);
nand UO_256 (O_256,N_14801,N_14704);
and UO_257 (O_257,N_13871,N_14594);
nor UO_258 (O_258,N_14872,N_14121);
nand UO_259 (O_259,N_14243,N_13995);
nor UO_260 (O_260,N_14952,N_13570);
nand UO_261 (O_261,N_14399,N_14486);
nand UO_262 (O_262,N_14466,N_14668);
and UO_263 (O_263,N_14066,N_14434);
nand UO_264 (O_264,N_14985,N_14467);
xnor UO_265 (O_265,N_14136,N_14789);
or UO_266 (O_266,N_13615,N_14100);
nor UO_267 (O_267,N_13776,N_14724);
xor UO_268 (O_268,N_14048,N_14612);
and UO_269 (O_269,N_14116,N_14816);
or UO_270 (O_270,N_14141,N_14003);
or UO_271 (O_271,N_14390,N_14237);
nand UO_272 (O_272,N_14964,N_14808);
xnor UO_273 (O_273,N_13878,N_14779);
or UO_274 (O_274,N_14990,N_13751);
nor UO_275 (O_275,N_14705,N_14604);
nand UO_276 (O_276,N_14569,N_14002);
and UO_277 (O_277,N_14796,N_14993);
nand UO_278 (O_278,N_14657,N_14380);
nor UO_279 (O_279,N_14558,N_14028);
or UO_280 (O_280,N_14500,N_14978);
nor UO_281 (O_281,N_13855,N_14611);
nand UO_282 (O_282,N_13713,N_13852);
nand UO_283 (O_283,N_14974,N_14296);
nand UO_284 (O_284,N_14382,N_13544);
and UO_285 (O_285,N_14794,N_13623);
or UO_286 (O_286,N_13848,N_14868);
nand UO_287 (O_287,N_13822,N_14914);
nand UO_288 (O_288,N_14933,N_13579);
or UO_289 (O_289,N_14053,N_13811);
or UO_290 (O_290,N_14949,N_14433);
nand UO_291 (O_291,N_14354,N_14795);
nand UO_292 (O_292,N_14677,N_14133);
nor UO_293 (O_293,N_14321,N_13796);
nor UO_294 (O_294,N_13685,N_13556);
nand UO_295 (O_295,N_14110,N_14122);
xnor UO_296 (O_296,N_14531,N_14610);
nand UO_297 (O_297,N_13806,N_14513);
or UO_298 (O_298,N_13900,N_13510);
nand UO_299 (O_299,N_13735,N_14280);
or UO_300 (O_300,N_14734,N_14018);
or UO_301 (O_301,N_14242,N_14645);
nor UO_302 (O_302,N_14841,N_14875);
and UO_303 (O_303,N_14685,N_14700);
or UO_304 (O_304,N_14215,N_13869);
xnor UO_305 (O_305,N_14134,N_13934);
and UO_306 (O_306,N_14043,N_14892);
nor UO_307 (O_307,N_14562,N_13664);
and UO_308 (O_308,N_14856,N_13581);
and UO_309 (O_309,N_14089,N_14419);
or UO_310 (O_310,N_14303,N_13921);
or UO_311 (O_311,N_14278,N_14566);
or UO_312 (O_312,N_13791,N_14623);
or UO_313 (O_313,N_13587,N_14007);
nand UO_314 (O_314,N_13881,N_13743);
nand UO_315 (O_315,N_13969,N_13913);
nand UO_316 (O_316,N_14963,N_14055);
and UO_317 (O_317,N_14541,N_14341);
nor UO_318 (O_318,N_14701,N_14375);
nor UO_319 (O_319,N_13691,N_13662);
or UO_320 (O_320,N_14201,N_13927);
or UO_321 (O_321,N_14476,N_14568);
or UO_322 (O_322,N_13764,N_14780);
or UO_323 (O_323,N_13652,N_13841);
nand UO_324 (O_324,N_14252,N_14503);
nor UO_325 (O_325,N_14858,N_14331);
or UO_326 (O_326,N_14882,N_14426);
nand UO_327 (O_327,N_14076,N_14309);
nand UO_328 (O_328,N_14563,N_13763);
nor UO_329 (O_329,N_13778,N_13741);
or UO_330 (O_330,N_14718,N_13988);
xor UO_331 (O_331,N_14367,N_14000);
and UO_332 (O_332,N_13794,N_13948);
nor UO_333 (O_333,N_14980,N_14361);
nand UO_334 (O_334,N_13627,N_14983);
nor UO_335 (O_335,N_14651,N_14766);
or UO_336 (O_336,N_14373,N_14058);
or UO_337 (O_337,N_14251,N_14070);
and UO_338 (O_338,N_14005,N_13962);
and UO_339 (O_339,N_13955,N_13820);
nand UO_340 (O_340,N_14155,N_14227);
and UO_341 (O_341,N_14601,N_14103);
nor UO_342 (O_342,N_13588,N_14479);
nor UO_343 (O_343,N_14477,N_13600);
nand UO_344 (O_344,N_13880,N_14965);
nor UO_345 (O_345,N_14127,N_14575);
or UO_346 (O_346,N_14936,N_13864);
nand UO_347 (O_347,N_14694,N_14098);
nor UO_348 (O_348,N_14553,N_14279);
and UO_349 (O_349,N_14630,N_13674);
nor UO_350 (O_350,N_14818,N_14085);
or UO_351 (O_351,N_14587,N_13703);
nand UO_352 (O_352,N_14996,N_14955);
nor UO_353 (O_353,N_14245,N_13561);
nor UO_354 (O_354,N_14307,N_14462);
nor UO_355 (O_355,N_14573,N_14784);
nor UO_356 (O_356,N_13530,N_13596);
and UO_357 (O_357,N_14720,N_14707);
nand UO_358 (O_358,N_14879,N_14205);
and UO_359 (O_359,N_14846,N_14355);
and UO_360 (O_360,N_13785,N_14071);
xor UO_361 (O_361,N_13516,N_14546);
nor UO_362 (O_362,N_13502,N_13779);
xnor UO_363 (O_363,N_14551,N_13633);
nor UO_364 (O_364,N_14897,N_14523);
and UO_365 (O_365,N_13882,N_13874);
and UO_366 (O_366,N_14235,N_14615);
and UO_367 (O_367,N_14637,N_14214);
or UO_368 (O_368,N_14204,N_14960);
nor UO_369 (O_369,N_14641,N_14586);
nor UO_370 (O_370,N_14223,N_14629);
nand UO_371 (O_371,N_13601,N_13920);
nor UO_372 (O_372,N_13668,N_14592);
nand UO_373 (O_373,N_13700,N_14027);
or UO_374 (O_374,N_14862,N_14900);
nor UO_375 (O_375,N_14843,N_14799);
or UO_376 (O_376,N_14662,N_14253);
nand UO_377 (O_377,N_14715,N_14403);
nor UO_378 (O_378,N_14831,N_14299);
nor UO_379 (O_379,N_14542,N_14198);
and UO_380 (O_380,N_13865,N_14020);
nand UO_381 (O_381,N_14063,N_14888);
nor UO_382 (O_382,N_13972,N_14428);
nor UO_383 (O_383,N_14248,N_14982);
nor UO_384 (O_384,N_14924,N_14387);
or UO_385 (O_385,N_13738,N_14722);
and UO_386 (O_386,N_14883,N_14810);
nor UO_387 (O_387,N_14935,N_14062);
and UO_388 (O_388,N_14745,N_14941);
or UO_389 (O_389,N_13598,N_13760);
and UO_390 (O_390,N_13547,N_14389);
or UO_391 (O_391,N_14516,N_13705);
or UO_392 (O_392,N_13831,N_14654);
and UO_393 (O_393,N_14213,N_14125);
nor UO_394 (O_394,N_14217,N_14202);
or UO_395 (O_395,N_14781,N_14750);
or UO_396 (O_396,N_13599,N_14366);
and UO_397 (O_397,N_14368,N_13790);
and UO_398 (O_398,N_14337,N_14678);
nand UO_399 (O_399,N_14986,N_14605);
nand UO_400 (O_400,N_14258,N_14464);
nor UO_401 (O_401,N_14736,N_13528);
nor UO_402 (O_402,N_14153,N_14454);
nor UO_403 (O_403,N_13895,N_13573);
or UO_404 (O_404,N_14591,N_14381);
or UO_405 (O_405,N_13908,N_14669);
or UO_406 (O_406,N_14973,N_13986);
nor UO_407 (O_407,N_13690,N_14943);
nand UO_408 (O_408,N_14975,N_14431);
nand UO_409 (O_409,N_13688,N_14314);
nor UO_410 (O_410,N_14738,N_14159);
nand UO_411 (O_411,N_14899,N_13755);
nand UO_412 (O_412,N_14411,N_13839);
nand UO_413 (O_413,N_13607,N_14441);
nand UO_414 (O_414,N_14514,N_13678);
or UO_415 (O_415,N_14104,N_14597);
nand UO_416 (O_416,N_14408,N_14440);
nor UO_417 (O_417,N_14474,N_14680);
nor UO_418 (O_418,N_14675,N_14589);
or UO_419 (O_419,N_13750,N_14906);
and UO_420 (O_420,N_13550,N_13879);
and UO_421 (O_421,N_13773,N_14057);
nand UO_422 (O_422,N_14602,N_14402);
nor UO_423 (O_423,N_13944,N_13651);
nand UO_424 (O_424,N_14903,N_14056);
nand UO_425 (O_425,N_14015,N_13641);
nand UO_426 (O_426,N_13616,N_13872);
nand UO_427 (O_427,N_14072,N_14723);
nand UO_428 (O_428,N_14424,N_13560);
nor UO_429 (O_429,N_14446,N_14939);
and UO_430 (O_430,N_14195,N_14929);
nand UO_431 (O_431,N_14509,N_13853);
or UO_432 (O_432,N_14762,N_13863);
nand UO_433 (O_433,N_13568,N_14778);
nor UO_434 (O_434,N_13998,N_13774);
nand UO_435 (O_435,N_14827,N_14088);
nand UO_436 (O_436,N_13947,N_14166);
or UO_437 (O_437,N_13954,N_14754);
nor UO_438 (O_438,N_14084,N_14828);
nand UO_439 (O_439,N_13732,N_13522);
nand UO_440 (O_440,N_14442,N_14060);
nand UO_441 (O_441,N_14880,N_14432);
and UO_442 (O_442,N_14544,N_13775);
nand UO_443 (O_443,N_13663,N_14971);
nand UO_444 (O_444,N_14647,N_13553);
nor UO_445 (O_445,N_14236,N_14537);
or UO_446 (O_446,N_14714,N_14776);
nand UO_447 (O_447,N_14576,N_14393);
nor UO_448 (O_448,N_14695,N_13929);
nor UO_449 (O_449,N_14490,N_13718);
and UO_450 (O_450,N_13898,N_14861);
and UO_451 (O_451,N_14224,N_13612);
or UO_452 (O_452,N_14803,N_13849);
nand UO_453 (O_453,N_14593,N_13868);
and UO_454 (O_454,N_14852,N_13546);
nand UO_455 (O_455,N_14295,N_13592);
and UO_456 (O_456,N_14061,N_13737);
and UO_457 (O_457,N_13837,N_13990);
and UO_458 (O_458,N_13605,N_14333);
nand UO_459 (O_459,N_13537,N_14097);
and UO_460 (O_460,N_14643,N_14817);
nand UO_461 (O_461,N_14025,N_13686);
or UO_462 (O_462,N_14407,N_14187);
and UO_463 (O_463,N_14659,N_13610);
and UO_464 (O_464,N_14310,N_14273);
or UO_465 (O_465,N_14699,N_14895);
nand UO_466 (O_466,N_13636,N_14640);
nand UO_467 (O_467,N_13805,N_14492);
nand UO_468 (O_468,N_14690,N_14535);
and UO_469 (O_469,N_14930,N_14396);
or UO_470 (O_470,N_14249,N_13597);
nor UO_471 (O_471,N_13888,N_13917);
or UO_472 (O_472,N_14238,N_13720);
or UO_473 (O_473,N_13746,N_13766);
nand UO_474 (O_474,N_13787,N_14792);
or UO_475 (O_475,N_13500,N_14124);
nand UO_476 (O_476,N_13541,N_14435);
or UO_477 (O_477,N_13639,N_14567);
nand UO_478 (O_478,N_14838,N_13996);
and UO_479 (O_479,N_14859,N_14913);
nand UO_480 (O_480,N_14969,N_14313);
or UO_481 (O_481,N_14320,N_14916);
nor UO_482 (O_482,N_14383,N_13877);
and UO_483 (O_483,N_14842,N_13723);
nor UO_484 (O_484,N_14526,N_14547);
and UO_485 (O_485,N_14199,N_14241);
nand UO_486 (O_486,N_14739,N_13749);
nor UO_487 (O_487,N_14741,N_13957);
nor UO_488 (O_488,N_13966,N_14866);
or UO_489 (O_489,N_13697,N_14068);
nand UO_490 (O_490,N_14765,N_14802);
nand UO_491 (O_491,N_13666,N_14376);
or UO_492 (O_492,N_13964,N_14911);
and UO_493 (O_493,N_14854,N_14413);
nor UO_494 (O_494,N_14864,N_14338);
nand UO_495 (O_495,N_13631,N_14902);
nor UO_496 (O_496,N_14814,N_14760);
nand UO_497 (O_497,N_13758,N_14716);
nand UO_498 (O_498,N_14093,N_14857);
and UO_499 (O_499,N_14771,N_13994);
or UO_500 (O_500,N_14269,N_13885);
and UO_501 (O_501,N_14702,N_14172);
nor UO_502 (O_502,N_14334,N_14473);
or UO_503 (O_503,N_14962,N_14670);
and UO_504 (O_504,N_14748,N_14197);
nor UO_505 (O_505,N_13654,N_14977);
or UO_506 (O_506,N_13906,N_13714);
nor UO_507 (O_507,N_14650,N_14206);
nor UO_508 (O_508,N_14679,N_14620);
or UO_509 (O_509,N_14998,N_13611);
or UO_510 (O_510,N_13548,N_14370);
and UO_511 (O_511,N_13508,N_13702);
nor UO_512 (O_512,N_13582,N_14012);
and UO_513 (O_513,N_14976,N_13956);
or UO_514 (O_514,N_13835,N_14272);
nor UO_515 (O_515,N_14894,N_14420);
nor UO_516 (O_516,N_14014,N_14860);
nor UO_517 (O_517,N_13624,N_14259);
or UO_518 (O_518,N_14222,N_14220);
nand UO_519 (O_519,N_14953,N_14078);
or UO_520 (O_520,N_14730,N_14228);
nand UO_521 (O_521,N_14735,N_13950);
or UO_522 (O_522,N_13829,N_14276);
and UO_523 (O_523,N_14436,N_13659);
nand UO_524 (O_524,N_14105,N_14688);
nor UO_525 (O_525,N_14283,N_13722);
nand UO_526 (O_526,N_13812,N_14485);
nor UO_527 (O_527,N_14603,N_14848);
or UO_528 (O_528,N_14530,N_14959);
or UO_529 (O_529,N_14323,N_13930);
and UO_530 (O_530,N_14809,N_14889);
nor UO_531 (O_531,N_14499,N_14826);
nor UO_532 (O_532,N_14815,N_13845);
or UO_533 (O_533,N_13653,N_14740);
nor UO_534 (O_534,N_13936,N_14483);
and UO_535 (O_535,N_14308,N_14386);
and UO_536 (O_536,N_14123,N_13539);
or UO_537 (O_537,N_14081,N_13858);
and UO_538 (O_538,N_14465,N_14507);
nor UO_539 (O_539,N_14564,N_14574);
nand UO_540 (O_540,N_14395,N_14984);
or UO_541 (O_541,N_14881,N_13563);
nor UO_542 (O_542,N_13562,N_13657);
or UO_543 (O_543,N_14032,N_13533);
nor UO_544 (O_544,N_13715,N_13771);
nor UO_545 (O_545,N_14561,N_14495);
nand UO_546 (O_546,N_14884,N_14772);
or UO_547 (O_547,N_14019,N_14453);
and UO_548 (O_548,N_14412,N_14359);
and UO_549 (O_549,N_14787,N_14254);
and UO_550 (O_550,N_13632,N_14340);
nor UO_551 (O_551,N_14829,N_13696);
nand UO_552 (O_552,N_14504,N_14497);
or UO_553 (O_553,N_14126,N_14992);
nand UO_554 (O_554,N_14836,N_14921);
and UO_555 (O_555,N_14286,N_14111);
or UO_556 (O_556,N_14636,N_14527);
and UO_557 (O_557,N_13973,N_13935);
nor UO_558 (O_558,N_14229,N_14064);
nand UO_559 (O_559,N_13847,N_13815);
nand UO_560 (O_560,N_13809,N_14559);
nand UO_561 (O_561,N_14102,N_14114);
and UO_562 (O_562,N_14302,N_13859);
xnor UO_563 (O_563,N_13850,N_13578);
or UO_564 (O_564,N_13709,N_13924);
nor UO_565 (O_565,N_14392,N_13968);
or UO_566 (O_566,N_14144,N_13567);
nor UO_567 (O_567,N_13506,N_14622);
nor UO_568 (O_568,N_13983,N_14157);
or UO_569 (O_569,N_14773,N_14405);
nand UO_570 (O_570,N_14519,N_14585);
xnor UO_571 (O_571,N_14822,N_14981);
or UO_572 (O_572,N_14324,N_14819);
or UO_573 (O_573,N_13549,N_13557);
or UO_574 (O_574,N_14737,N_13759);
nand UO_575 (O_575,N_14118,N_14550);
nand UO_576 (O_576,N_14851,N_14385);
or UO_577 (O_577,N_13893,N_14425);
nor UO_578 (O_578,N_14108,N_14186);
or UO_579 (O_579,N_13976,N_14158);
or UO_580 (O_580,N_14244,N_14671);
nand UO_581 (O_581,N_14863,N_14793);
and UO_582 (O_582,N_14306,N_14470);
or UO_583 (O_583,N_13940,N_14834);
and UO_584 (O_584,N_14532,N_14946);
or UO_585 (O_585,N_14478,N_14330);
nor UO_586 (O_586,N_13828,N_13980);
nand UO_587 (O_587,N_13919,N_14207);
or UO_588 (O_588,N_14461,N_14135);
nor UO_589 (O_589,N_14655,N_13670);
or UO_590 (O_590,N_14664,N_13843);
or UO_591 (O_591,N_14231,N_13910);
nand UO_592 (O_592,N_14521,N_14011);
nor UO_593 (O_593,N_14667,N_14404);
nand UO_594 (O_594,N_13710,N_13899);
nor UO_595 (O_595,N_14887,N_13993);
and UO_596 (O_596,N_14165,N_13523);
or UO_597 (O_597,N_14073,N_14769);
nand UO_598 (O_598,N_14505,N_13540);
nand UO_599 (O_599,N_13933,N_13734);
nor UO_600 (O_600,N_13515,N_14179);
and UO_601 (O_601,N_14059,N_14753);
nand UO_602 (O_602,N_14502,N_13672);
and UO_603 (O_603,N_13514,N_14931);
nor UO_604 (O_604,N_13926,N_14281);
and UO_605 (O_605,N_14374,N_14554);
or UO_606 (O_606,N_13978,N_14024);
and UO_607 (O_607,N_13681,N_14693);
or UO_608 (O_608,N_13513,N_13960);
or UO_609 (O_609,N_13909,N_14627);
or UO_610 (O_610,N_14904,N_14950);
nand UO_611 (O_611,N_13772,N_14145);
or UO_612 (O_612,N_13630,N_14013);
or UO_613 (O_613,N_14606,N_14954);
and UO_614 (O_614,N_13767,N_14211);
xnor UO_615 (O_615,N_14065,N_14511);
or UO_616 (O_616,N_14030,N_13706);
and UO_617 (O_617,N_13836,N_14631);
nor UO_618 (O_618,N_14757,N_14837);
nor UO_619 (O_619,N_14555,N_13958);
nor UO_620 (O_620,N_14328,N_13614);
and UO_621 (O_621,N_14457,N_14642);
nand UO_622 (O_622,N_14489,N_13949);
nand UO_623 (O_623,N_13818,N_14909);
or UO_624 (O_624,N_14260,N_13762);
nand UO_625 (O_625,N_14777,N_14372);
nor UO_626 (O_626,N_14972,N_13875);
nand UO_627 (O_627,N_13626,N_14268);
nand UO_628 (O_628,N_14422,N_13825);
or UO_629 (O_629,N_13777,N_14698);
nor UO_630 (O_630,N_13939,N_14635);
nor UO_631 (O_631,N_14391,N_14301);
nand UO_632 (O_632,N_13717,N_14146);
nand UO_633 (O_633,N_13660,N_14613);
or UO_634 (O_634,N_14074,N_14608);
nand UO_635 (O_635,N_13511,N_14891);
nand UO_636 (O_636,N_14925,N_13886);
or UO_637 (O_637,N_14767,N_14672);
or UO_638 (O_638,N_14825,N_14357);
nand UO_639 (O_639,N_13564,N_14082);
or UO_640 (O_640,N_14079,N_13671);
nor UO_641 (O_641,N_13752,N_13638);
nor UO_642 (O_642,N_14416,N_14325);
or UO_643 (O_643,N_13529,N_13981);
nor UO_644 (O_644,N_13757,N_14583);
or UO_645 (O_645,N_14218,N_14216);
or UO_646 (O_646,N_13620,N_13844);
and UO_647 (O_647,N_14524,N_13916);
or UO_648 (O_648,N_13745,N_14080);
and UO_649 (O_649,N_13931,N_13784);
or UO_650 (O_650,N_13535,N_14004);
nand UO_651 (O_651,N_14821,N_14267);
or UO_652 (O_652,N_14703,N_14311);
nor UO_653 (O_653,N_14106,N_14689);
or UO_654 (O_654,N_13545,N_14096);
and UO_655 (O_655,N_13584,N_14463);
xor UO_656 (O_656,N_13833,N_14595);
nor UO_657 (O_657,N_14099,N_14995);
nor UO_658 (O_658,N_14163,N_14265);
or UO_659 (O_659,N_14362,N_13814);
and UO_660 (O_660,N_14646,N_13846);
and UO_661 (O_661,N_14318,N_13608);
nand UO_662 (O_662,N_14266,N_13781);
and UO_663 (O_663,N_13740,N_14596);
or UO_664 (O_664,N_13810,N_14086);
nand UO_665 (O_665,N_14468,N_13669);
nor UO_666 (O_666,N_14571,N_14067);
nor UO_667 (O_667,N_14719,N_14824);
nand UO_668 (O_668,N_14212,N_14458);
and UO_669 (O_669,N_13826,N_13902);
or UO_670 (O_670,N_14548,N_14763);
or UO_671 (O_671,N_14994,N_13727);
and UO_672 (O_672,N_14919,N_14653);
nand UO_673 (O_673,N_14733,N_14190);
and UO_674 (O_674,N_14455,N_13525);
or UO_675 (O_675,N_14443,N_14250);
nand UO_676 (O_676,N_13692,N_14147);
nor UO_677 (O_677,N_13860,N_14400);
or UO_678 (O_678,N_13609,N_14706);
nand UO_679 (O_679,N_14966,N_14847);
nor UO_680 (O_680,N_14539,N_14191);
nor UO_681 (O_681,N_14017,N_14288);
and UO_682 (O_682,N_13575,N_14021);
nor UO_683 (O_683,N_14853,N_13538);
xor UO_684 (O_684,N_14421,N_13586);
nand UO_685 (O_685,N_14196,N_14528);
nand UO_686 (O_686,N_14247,N_13974);
or UO_687 (O_687,N_13552,N_14957);
nand UO_688 (O_688,N_14351,N_13649);
nand UO_689 (O_689,N_14360,N_14487);
nand UO_690 (O_690,N_14652,N_14031);
nor UO_691 (O_691,N_14289,N_13977);
nand UO_692 (O_692,N_13645,N_14182);
xnor UO_693 (O_693,N_13695,N_14676);
and UO_694 (O_694,N_14481,N_14758);
nand UO_695 (O_695,N_14496,N_13925);
nor UO_696 (O_696,N_14666,N_14624);
and UO_697 (O_697,N_14928,N_13647);
and UO_698 (O_698,N_14171,N_13827);
nor UO_699 (O_699,N_14625,N_13571);
nand UO_700 (O_700,N_13572,N_14893);
nor UO_701 (O_701,N_14129,N_13918);
xor UO_702 (O_702,N_14785,N_14747);
nand UO_703 (O_703,N_14298,N_13830);
nand UO_704 (O_704,N_13594,N_14128);
or UO_705 (O_705,N_13804,N_13729);
or UO_706 (O_706,N_14989,N_14026);
xnor UO_707 (O_707,N_14365,N_13997);
or UO_708 (O_708,N_14471,N_13505);
or UO_709 (O_709,N_14161,N_14988);
and UO_710 (O_710,N_14183,N_14917);
nor UO_711 (O_711,N_13520,N_14226);
nand UO_712 (O_712,N_13635,N_13634);
and UO_713 (O_713,N_14491,N_14316);
nand UO_714 (O_714,N_13786,N_13890);
nor UO_715 (O_715,N_14449,N_13807);
or UO_716 (O_716,N_14619,N_14788);
and UO_717 (O_717,N_14075,N_14886);
nand UO_718 (O_718,N_14038,N_14347);
and UO_719 (O_719,N_13619,N_13754);
or UO_720 (O_720,N_13646,N_13504);
or UO_721 (O_721,N_14713,N_13896);
nor UO_722 (O_722,N_14448,N_13707);
or UO_723 (O_723,N_14920,N_14037);
nand UO_724 (O_724,N_14582,N_14632);
or UO_725 (O_725,N_13866,N_13591);
nand UO_726 (O_726,N_14709,N_14876);
nor UO_727 (O_727,N_14607,N_14140);
nor UO_728 (O_728,N_14346,N_13555);
or UO_729 (O_729,N_13724,N_13963);
nor UO_730 (O_730,N_13642,N_14512);
nor UO_731 (O_731,N_14588,N_14327);
or UO_732 (O_732,N_14456,N_14095);
or UO_733 (O_733,N_13989,N_13527);
and UO_734 (O_734,N_14830,N_13559);
and UO_735 (O_735,N_13951,N_14275);
or UO_736 (O_736,N_14263,N_14284);
nor UO_737 (O_737,N_14350,N_14287);
nand UO_738 (O_738,N_13861,N_14178);
and UO_739 (O_739,N_13938,N_14480);
nand UO_740 (O_740,N_14721,N_14087);
nor UO_741 (O_741,N_14967,N_13800);
or UO_742 (O_742,N_14083,N_14556);
and UO_743 (O_743,N_14898,N_14022);
nand UO_744 (O_744,N_14271,N_14130);
nand UO_745 (O_745,N_14774,N_14132);
or UO_746 (O_746,N_14358,N_14865);
or UO_747 (O_747,N_13922,N_14565);
and UO_748 (O_748,N_14681,N_14047);
nor UO_749 (O_749,N_14185,N_14475);
nor UO_750 (O_750,N_14168,N_13548);
or UO_751 (O_751,N_14502,N_13901);
and UO_752 (O_752,N_14974,N_14278);
nor UO_753 (O_753,N_14933,N_14099);
and UO_754 (O_754,N_14685,N_14593);
nand UO_755 (O_755,N_14004,N_14530);
or UO_756 (O_756,N_14539,N_13657);
nand UO_757 (O_757,N_13691,N_13606);
or UO_758 (O_758,N_14735,N_14878);
and UO_759 (O_759,N_14059,N_13606);
and UO_760 (O_760,N_14526,N_13927);
nor UO_761 (O_761,N_13777,N_14278);
nor UO_762 (O_762,N_14658,N_13949);
or UO_763 (O_763,N_14014,N_14536);
or UO_764 (O_764,N_13883,N_13841);
nand UO_765 (O_765,N_14256,N_14348);
and UO_766 (O_766,N_14116,N_13794);
and UO_767 (O_767,N_14337,N_13672);
nor UO_768 (O_768,N_14489,N_14244);
or UO_769 (O_769,N_13629,N_14060);
nor UO_770 (O_770,N_13774,N_14548);
nand UO_771 (O_771,N_14376,N_14433);
nand UO_772 (O_772,N_14061,N_14567);
nor UO_773 (O_773,N_13993,N_14859);
nand UO_774 (O_774,N_14690,N_14391);
nor UO_775 (O_775,N_14075,N_13665);
nor UO_776 (O_776,N_14099,N_14738);
or UO_777 (O_777,N_14847,N_14939);
nand UO_778 (O_778,N_13891,N_13636);
nor UO_779 (O_779,N_13673,N_13671);
nand UO_780 (O_780,N_14942,N_14685);
nor UO_781 (O_781,N_14204,N_13791);
nand UO_782 (O_782,N_14138,N_14354);
nor UO_783 (O_783,N_14186,N_14870);
and UO_784 (O_784,N_14886,N_14339);
or UO_785 (O_785,N_14728,N_14233);
nand UO_786 (O_786,N_14776,N_14500);
and UO_787 (O_787,N_13663,N_14136);
nor UO_788 (O_788,N_13668,N_13671);
or UO_789 (O_789,N_14260,N_14362);
nor UO_790 (O_790,N_14275,N_13775);
nor UO_791 (O_791,N_13684,N_14572);
nand UO_792 (O_792,N_14196,N_14813);
nor UO_793 (O_793,N_14305,N_14170);
nor UO_794 (O_794,N_13896,N_13620);
and UO_795 (O_795,N_14887,N_13955);
and UO_796 (O_796,N_14633,N_14998);
nor UO_797 (O_797,N_14074,N_14131);
nor UO_798 (O_798,N_13567,N_13949);
nor UO_799 (O_799,N_14326,N_13755);
and UO_800 (O_800,N_14437,N_14969);
nand UO_801 (O_801,N_13921,N_14410);
nor UO_802 (O_802,N_14067,N_14033);
nand UO_803 (O_803,N_14515,N_14618);
and UO_804 (O_804,N_13993,N_13683);
and UO_805 (O_805,N_14377,N_14952);
or UO_806 (O_806,N_14472,N_13742);
nor UO_807 (O_807,N_13682,N_14046);
and UO_808 (O_808,N_14743,N_14590);
nand UO_809 (O_809,N_13663,N_14229);
or UO_810 (O_810,N_13566,N_14229);
and UO_811 (O_811,N_14998,N_14114);
and UO_812 (O_812,N_14853,N_14366);
nand UO_813 (O_813,N_13783,N_14355);
nor UO_814 (O_814,N_14335,N_14303);
xor UO_815 (O_815,N_14552,N_14279);
and UO_816 (O_816,N_14179,N_14902);
nand UO_817 (O_817,N_13956,N_13574);
and UO_818 (O_818,N_14950,N_14431);
nor UO_819 (O_819,N_14670,N_14740);
nand UO_820 (O_820,N_13689,N_14096);
nor UO_821 (O_821,N_14443,N_14353);
nor UO_822 (O_822,N_14635,N_13717);
nor UO_823 (O_823,N_14697,N_14677);
and UO_824 (O_824,N_14608,N_13955);
or UO_825 (O_825,N_14259,N_14329);
nand UO_826 (O_826,N_14297,N_13576);
and UO_827 (O_827,N_14162,N_14644);
nor UO_828 (O_828,N_14940,N_14546);
nand UO_829 (O_829,N_13647,N_14646);
and UO_830 (O_830,N_13993,N_13917);
nor UO_831 (O_831,N_14982,N_14501);
nand UO_832 (O_832,N_14581,N_14018);
or UO_833 (O_833,N_13645,N_14089);
nor UO_834 (O_834,N_13804,N_13513);
nor UO_835 (O_835,N_14099,N_14024);
and UO_836 (O_836,N_14284,N_13966);
and UO_837 (O_837,N_14584,N_14763);
nor UO_838 (O_838,N_14876,N_14349);
nor UO_839 (O_839,N_14080,N_14507);
or UO_840 (O_840,N_14888,N_13833);
and UO_841 (O_841,N_14515,N_14436);
nor UO_842 (O_842,N_14475,N_14758);
or UO_843 (O_843,N_13976,N_13723);
nor UO_844 (O_844,N_14340,N_14963);
and UO_845 (O_845,N_14211,N_14336);
nor UO_846 (O_846,N_13831,N_14277);
nand UO_847 (O_847,N_14357,N_14725);
or UO_848 (O_848,N_14935,N_14212);
and UO_849 (O_849,N_14201,N_13991);
nor UO_850 (O_850,N_14813,N_14348);
and UO_851 (O_851,N_14921,N_14712);
or UO_852 (O_852,N_14806,N_14596);
or UO_853 (O_853,N_14922,N_14542);
and UO_854 (O_854,N_14283,N_13509);
nand UO_855 (O_855,N_13711,N_14632);
and UO_856 (O_856,N_13609,N_14525);
nand UO_857 (O_857,N_13550,N_14226);
nand UO_858 (O_858,N_13928,N_14588);
nand UO_859 (O_859,N_14994,N_13668);
or UO_860 (O_860,N_14433,N_13873);
nor UO_861 (O_861,N_13851,N_14976);
or UO_862 (O_862,N_14768,N_14580);
nor UO_863 (O_863,N_13969,N_14583);
nand UO_864 (O_864,N_14920,N_13540);
and UO_865 (O_865,N_13683,N_14894);
nor UO_866 (O_866,N_14281,N_14319);
nor UO_867 (O_867,N_14516,N_14214);
or UO_868 (O_868,N_13953,N_14290);
xnor UO_869 (O_869,N_13762,N_14027);
and UO_870 (O_870,N_14156,N_14901);
or UO_871 (O_871,N_14598,N_13826);
and UO_872 (O_872,N_13836,N_14533);
and UO_873 (O_873,N_14780,N_14042);
and UO_874 (O_874,N_13702,N_14673);
xnor UO_875 (O_875,N_13971,N_14662);
nand UO_876 (O_876,N_13655,N_14952);
and UO_877 (O_877,N_13778,N_14082);
and UO_878 (O_878,N_14379,N_13675);
nand UO_879 (O_879,N_14001,N_14385);
or UO_880 (O_880,N_14563,N_14997);
and UO_881 (O_881,N_14358,N_14036);
and UO_882 (O_882,N_13617,N_14514);
nand UO_883 (O_883,N_14776,N_14453);
nor UO_884 (O_884,N_14626,N_13546);
and UO_885 (O_885,N_14912,N_14132);
nand UO_886 (O_886,N_13761,N_14337);
nor UO_887 (O_887,N_13819,N_14144);
or UO_888 (O_888,N_13935,N_13914);
and UO_889 (O_889,N_14275,N_13600);
or UO_890 (O_890,N_13729,N_14407);
or UO_891 (O_891,N_13968,N_14909);
or UO_892 (O_892,N_13659,N_14887);
xor UO_893 (O_893,N_13681,N_13545);
and UO_894 (O_894,N_14225,N_13680);
nor UO_895 (O_895,N_14161,N_14945);
or UO_896 (O_896,N_13559,N_14016);
nand UO_897 (O_897,N_14772,N_13964);
nand UO_898 (O_898,N_14961,N_14091);
nor UO_899 (O_899,N_14814,N_14968);
and UO_900 (O_900,N_14215,N_14697);
or UO_901 (O_901,N_13681,N_14222);
nand UO_902 (O_902,N_13935,N_14900);
nor UO_903 (O_903,N_14565,N_14534);
nand UO_904 (O_904,N_14431,N_14960);
or UO_905 (O_905,N_14006,N_14080);
xor UO_906 (O_906,N_13520,N_13898);
or UO_907 (O_907,N_14059,N_13552);
nand UO_908 (O_908,N_13672,N_13872);
or UO_909 (O_909,N_13875,N_14323);
nand UO_910 (O_910,N_13812,N_14152);
nand UO_911 (O_911,N_14352,N_13539);
nor UO_912 (O_912,N_13918,N_14641);
nor UO_913 (O_913,N_14778,N_13584);
nand UO_914 (O_914,N_14040,N_13513);
and UO_915 (O_915,N_14218,N_14295);
or UO_916 (O_916,N_14838,N_13801);
and UO_917 (O_917,N_13526,N_13918);
nor UO_918 (O_918,N_14021,N_13569);
or UO_919 (O_919,N_13878,N_14117);
and UO_920 (O_920,N_14458,N_14434);
or UO_921 (O_921,N_14466,N_14078);
nor UO_922 (O_922,N_13567,N_14081);
nor UO_923 (O_923,N_13533,N_14151);
nand UO_924 (O_924,N_14856,N_13959);
nor UO_925 (O_925,N_14526,N_14537);
nand UO_926 (O_926,N_14880,N_14461);
or UO_927 (O_927,N_13936,N_14510);
and UO_928 (O_928,N_14199,N_14679);
nand UO_929 (O_929,N_13825,N_14772);
or UO_930 (O_930,N_13830,N_14993);
or UO_931 (O_931,N_14954,N_13868);
nand UO_932 (O_932,N_14277,N_14607);
nand UO_933 (O_933,N_13597,N_14511);
and UO_934 (O_934,N_14194,N_13904);
and UO_935 (O_935,N_14815,N_13614);
nor UO_936 (O_936,N_13584,N_14440);
or UO_937 (O_937,N_14652,N_13554);
nand UO_938 (O_938,N_14316,N_13897);
and UO_939 (O_939,N_14701,N_14770);
nor UO_940 (O_940,N_14488,N_14996);
and UO_941 (O_941,N_14697,N_13995);
nor UO_942 (O_942,N_13552,N_14398);
nor UO_943 (O_943,N_14334,N_14469);
nand UO_944 (O_944,N_13781,N_14977);
or UO_945 (O_945,N_13952,N_14472);
or UO_946 (O_946,N_13820,N_13855);
nand UO_947 (O_947,N_14244,N_14784);
or UO_948 (O_948,N_14777,N_14570);
or UO_949 (O_949,N_13517,N_14706);
and UO_950 (O_950,N_13663,N_14784);
or UO_951 (O_951,N_14621,N_14216);
nor UO_952 (O_952,N_14186,N_14843);
or UO_953 (O_953,N_14910,N_14755);
nor UO_954 (O_954,N_14281,N_14336);
nor UO_955 (O_955,N_14721,N_14026);
nor UO_956 (O_956,N_14655,N_14900);
or UO_957 (O_957,N_14550,N_14120);
or UO_958 (O_958,N_14181,N_14179);
nor UO_959 (O_959,N_14717,N_13968);
nor UO_960 (O_960,N_14309,N_14749);
nand UO_961 (O_961,N_14403,N_14390);
nor UO_962 (O_962,N_14170,N_13890);
nor UO_963 (O_963,N_13628,N_14081);
or UO_964 (O_964,N_14020,N_14180);
nor UO_965 (O_965,N_14372,N_14838);
nor UO_966 (O_966,N_13662,N_13512);
nand UO_967 (O_967,N_14464,N_13684);
and UO_968 (O_968,N_13630,N_13525);
or UO_969 (O_969,N_14776,N_13929);
and UO_970 (O_970,N_14999,N_13793);
or UO_971 (O_971,N_14891,N_14610);
or UO_972 (O_972,N_14260,N_14412);
nand UO_973 (O_973,N_14091,N_13943);
nand UO_974 (O_974,N_14344,N_13621);
nand UO_975 (O_975,N_13537,N_14259);
or UO_976 (O_976,N_14247,N_14031);
nand UO_977 (O_977,N_14446,N_14135);
or UO_978 (O_978,N_14600,N_14066);
or UO_979 (O_979,N_13758,N_14684);
and UO_980 (O_980,N_13650,N_14620);
or UO_981 (O_981,N_13695,N_14267);
and UO_982 (O_982,N_14720,N_13606);
nor UO_983 (O_983,N_14421,N_14356);
nand UO_984 (O_984,N_14985,N_14144);
and UO_985 (O_985,N_14697,N_13829);
nor UO_986 (O_986,N_14490,N_13532);
nand UO_987 (O_987,N_14149,N_13793);
and UO_988 (O_988,N_13950,N_14986);
nand UO_989 (O_989,N_14189,N_14979);
nand UO_990 (O_990,N_13649,N_14260);
xnor UO_991 (O_991,N_13836,N_14291);
nor UO_992 (O_992,N_14425,N_14451);
or UO_993 (O_993,N_13862,N_14706);
nor UO_994 (O_994,N_14923,N_14944);
and UO_995 (O_995,N_13843,N_14002);
nand UO_996 (O_996,N_14920,N_14990);
and UO_997 (O_997,N_14918,N_14241);
nor UO_998 (O_998,N_14314,N_13770);
and UO_999 (O_999,N_14734,N_14201);
nand UO_1000 (O_1000,N_13643,N_13510);
nor UO_1001 (O_1001,N_13892,N_13902);
or UO_1002 (O_1002,N_14653,N_13707);
nor UO_1003 (O_1003,N_13662,N_14172);
nand UO_1004 (O_1004,N_14361,N_14679);
or UO_1005 (O_1005,N_14636,N_14384);
nor UO_1006 (O_1006,N_14851,N_14946);
or UO_1007 (O_1007,N_14256,N_14798);
nand UO_1008 (O_1008,N_14151,N_14335);
nand UO_1009 (O_1009,N_13771,N_14548);
and UO_1010 (O_1010,N_13853,N_14970);
nor UO_1011 (O_1011,N_13805,N_14695);
or UO_1012 (O_1012,N_13758,N_14116);
or UO_1013 (O_1013,N_14089,N_14138);
nor UO_1014 (O_1014,N_13900,N_14037);
or UO_1015 (O_1015,N_14928,N_13536);
nor UO_1016 (O_1016,N_13809,N_14577);
nor UO_1017 (O_1017,N_14546,N_14218);
nor UO_1018 (O_1018,N_14506,N_13966);
nand UO_1019 (O_1019,N_14530,N_14601);
nor UO_1020 (O_1020,N_13866,N_14932);
nand UO_1021 (O_1021,N_14578,N_14507);
nor UO_1022 (O_1022,N_14171,N_14497);
nand UO_1023 (O_1023,N_14220,N_14493);
nand UO_1024 (O_1024,N_14796,N_14023);
and UO_1025 (O_1025,N_14252,N_14866);
nand UO_1026 (O_1026,N_14672,N_14754);
nor UO_1027 (O_1027,N_13757,N_13656);
nor UO_1028 (O_1028,N_14780,N_14280);
and UO_1029 (O_1029,N_13953,N_14009);
or UO_1030 (O_1030,N_14833,N_13643);
and UO_1031 (O_1031,N_14872,N_14709);
or UO_1032 (O_1032,N_13761,N_14045);
nor UO_1033 (O_1033,N_14859,N_14174);
nand UO_1034 (O_1034,N_14020,N_13575);
or UO_1035 (O_1035,N_13717,N_14600);
nor UO_1036 (O_1036,N_14863,N_14467);
xnor UO_1037 (O_1037,N_14388,N_14434);
nand UO_1038 (O_1038,N_14777,N_14910);
and UO_1039 (O_1039,N_14472,N_14520);
and UO_1040 (O_1040,N_13655,N_14149);
or UO_1041 (O_1041,N_14141,N_13662);
or UO_1042 (O_1042,N_13670,N_14132);
and UO_1043 (O_1043,N_14230,N_14360);
nand UO_1044 (O_1044,N_13798,N_14560);
or UO_1045 (O_1045,N_13615,N_13729);
nand UO_1046 (O_1046,N_14204,N_14116);
nor UO_1047 (O_1047,N_14861,N_13529);
nor UO_1048 (O_1048,N_14921,N_14160);
or UO_1049 (O_1049,N_14903,N_13629);
and UO_1050 (O_1050,N_14760,N_13965);
nor UO_1051 (O_1051,N_13564,N_14282);
nor UO_1052 (O_1052,N_14699,N_14947);
nand UO_1053 (O_1053,N_14660,N_13839);
xnor UO_1054 (O_1054,N_14934,N_14499);
nand UO_1055 (O_1055,N_14634,N_14912);
nand UO_1056 (O_1056,N_14998,N_14506);
or UO_1057 (O_1057,N_14757,N_14124);
nor UO_1058 (O_1058,N_14348,N_14572);
or UO_1059 (O_1059,N_14982,N_13636);
or UO_1060 (O_1060,N_14866,N_14049);
or UO_1061 (O_1061,N_14967,N_14706);
nor UO_1062 (O_1062,N_14373,N_14062);
and UO_1063 (O_1063,N_14410,N_14390);
nor UO_1064 (O_1064,N_13643,N_13507);
nor UO_1065 (O_1065,N_14008,N_14104);
nor UO_1066 (O_1066,N_14452,N_14436);
nand UO_1067 (O_1067,N_14533,N_13732);
nand UO_1068 (O_1068,N_13779,N_14338);
and UO_1069 (O_1069,N_13934,N_14096);
or UO_1070 (O_1070,N_14710,N_13927);
and UO_1071 (O_1071,N_14307,N_13761);
xnor UO_1072 (O_1072,N_14765,N_13659);
and UO_1073 (O_1073,N_14075,N_13903);
or UO_1074 (O_1074,N_14440,N_14969);
or UO_1075 (O_1075,N_14305,N_14703);
and UO_1076 (O_1076,N_13842,N_14729);
nor UO_1077 (O_1077,N_13573,N_14927);
nor UO_1078 (O_1078,N_13779,N_13640);
nor UO_1079 (O_1079,N_14022,N_14121);
nand UO_1080 (O_1080,N_14030,N_14656);
or UO_1081 (O_1081,N_14139,N_14108);
nand UO_1082 (O_1082,N_14300,N_14764);
nand UO_1083 (O_1083,N_14767,N_14987);
and UO_1084 (O_1084,N_13944,N_14746);
nor UO_1085 (O_1085,N_13903,N_13504);
nand UO_1086 (O_1086,N_14852,N_14220);
and UO_1087 (O_1087,N_13613,N_13989);
and UO_1088 (O_1088,N_13616,N_14550);
and UO_1089 (O_1089,N_14237,N_14143);
and UO_1090 (O_1090,N_13614,N_14640);
nand UO_1091 (O_1091,N_14164,N_13705);
nor UO_1092 (O_1092,N_13997,N_14535);
or UO_1093 (O_1093,N_13898,N_14358);
nor UO_1094 (O_1094,N_14516,N_14942);
nor UO_1095 (O_1095,N_13848,N_14516);
nand UO_1096 (O_1096,N_14629,N_14824);
or UO_1097 (O_1097,N_14231,N_13862);
and UO_1098 (O_1098,N_14658,N_13942);
or UO_1099 (O_1099,N_14834,N_13501);
nor UO_1100 (O_1100,N_14509,N_13954);
and UO_1101 (O_1101,N_14102,N_14333);
nor UO_1102 (O_1102,N_13772,N_13918);
nand UO_1103 (O_1103,N_14195,N_14288);
nor UO_1104 (O_1104,N_14969,N_13738);
nor UO_1105 (O_1105,N_14869,N_14763);
nor UO_1106 (O_1106,N_14416,N_14492);
and UO_1107 (O_1107,N_14822,N_13990);
and UO_1108 (O_1108,N_13509,N_13896);
nor UO_1109 (O_1109,N_14131,N_13637);
nand UO_1110 (O_1110,N_14376,N_13832);
nor UO_1111 (O_1111,N_14630,N_14953);
and UO_1112 (O_1112,N_14567,N_14592);
or UO_1113 (O_1113,N_13764,N_14211);
nor UO_1114 (O_1114,N_13946,N_14291);
or UO_1115 (O_1115,N_14961,N_13790);
or UO_1116 (O_1116,N_14510,N_14966);
nand UO_1117 (O_1117,N_14450,N_14876);
nand UO_1118 (O_1118,N_14068,N_14437);
and UO_1119 (O_1119,N_13602,N_14350);
nor UO_1120 (O_1120,N_14857,N_13815);
and UO_1121 (O_1121,N_14277,N_13914);
nor UO_1122 (O_1122,N_14045,N_14332);
nand UO_1123 (O_1123,N_13616,N_14927);
nand UO_1124 (O_1124,N_14409,N_14539);
or UO_1125 (O_1125,N_14556,N_14656);
nor UO_1126 (O_1126,N_13630,N_14101);
or UO_1127 (O_1127,N_14268,N_13646);
nand UO_1128 (O_1128,N_13618,N_13697);
nand UO_1129 (O_1129,N_14013,N_13749);
or UO_1130 (O_1130,N_13916,N_13994);
nand UO_1131 (O_1131,N_14416,N_13970);
or UO_1132 (O_1132,N_14126,N_14176);
or UO_1133 (O_1133,N_14054,N_13907);
and UO_1134 (O_1134,N_13770,N_13743);
or UO_1135 (O_1135,N_14790,N_14124);
nor UO_1136 (O_1136,N_13636,N_14136);
nor UO_1137 (O_1137,N_13575,N_14836);
or UO_1138 (O_1138,N_13750,N_13811);
nor UO_1139 (O_1139,N_13774,N_13970);
nand UO_1140 (O_1140,N_14996,N_14170);
or UO_1141 (O_1141,N_14734,N_14692);
or UO_1142 (O_1142,N_14475,N_14940);
nor UO_1143 (O_1143,N_14231,N_14641);
or UO_1144 (O_1144,N_14638,N_13899);
xnor UO_1145 (O_1145,N_14495,N_13793);
nor UO_1146 (O_1146,N_14276,N_13916);
or UO_1147 (O_1147,N_14893,N_13968);
and UO_1148 (O_1148,N_13773,N_13781);
nor UO_1149 (O_1149,N_13984,N_14680);
and UO_1150 (O_1150,N_14909,N_13775);
nand UO_1151 (O_1151,N_13602,N_14157);
nand UO_1152 (O_1152,N_14941,N_13608);
nor UO_1153 (O_1153,N_14437,N_13518);
xor UO_1154 (O_1154,N_14598,N_14271);
nand UO_1155 (O_1155,N_13575,N_14562);
or UO_1156 (O_1156,N_14184,N_14787);
and UO_1157 (O_1157,N_13837,N_14711);
nor UO_1158 (O_1158,N_14504,N_13684);
nand UO_1159 (O_1159,N_14676,N_13986);
nor UO_1160 (O_1160,N_13648,N_14108);
nand UO_1161 (O_1161,N_13658,N_14484);
nor UO_1162 (O_1162,N_14119,N_14890);
xnor UO_1163 (O_1163,N_14940,N_14172);
nand UO_1164 (O_1164,N_14857,N_14417);
or UO_1165 (O_1165,N_14861,N_14315);
or UO_1166 (O_1166,N_14115,N_14948);
and UO_1167 (O_1167,N_13548,N_14783);
nand UO_1168 (O_1168,N_14682,N_13911);
xor UO_1169 (O_1169,N_14392,N_13548);
nand UO_1170 (O_1170,N_14039,N_14387);
xor UO_1171 (O_1171,N_14012,N_13558);
or UO_1172 (O_1172,N_13505,N_14887);
nor UO_1173 (O_1173,N_14164,N_14676);
nor UO_1174 (O_1174,N_14343,N_14964);
xor UO_1175 (O_1175,N_14115,N_13825);
or UO_1176 (O_1176,N_14450,N_14187);
nor UO_1177 (O_1177,N_14917,N_13637);
and UO_1178 (O_1178,N_14713,N_14319);
or UO_1179 (O_1179,N_14737,N_13544);
nand UO_1180 (O_1180,N_13632,N_14683);
or UO_1181 (O_1181,N_14022,N_14815);
and UO_1182 (O_1182,N_14489,N_14596);
nand UO_1183 (O_1183,N_14869,N_13984);
nand UO_1184 (O_1184,N_14948,N_14802);
or UO_1185 (O_1185,N_14807,N_14898);
nor UO_1186 (O_1186,N_14443,N_14302);
or UO_1187 (O_1187,N_14217,N_13820);
or UO_1188 (O_1188,N_13945,N_14011);
nor UO_1189 (O_1189,N_13782,N_14152);
or UO_1190 (O_1190,N_13590,N_14717);
nor UO_1191 (O_1191,N_14202,N_13994);
nand UO_1192 (O_1192,N_14641,N_14010);
nor UO_1193 (O_1193,N_14135,N_13606);
or UO_1194 (O_1194,N_14081,N_14129);
and UO_1195 (O_1195,N_14163,N_13521);
or UO_1196 (O_1196,N_13789,N_13993);
nor UO_1197 (O_1197,N_14591,N_14518);
or UO_1198 (O_1198,N_13712,N_14173);
nand UO_1199 (O_1199,N_14033,N_14194);
nor UO_1200 (O_1200,N_14866,N_14781);
or UO_1201 (O_1201,N_13627,N_14104);
or UO_1202 (O_1202,N_13731,N_14413);
nand UO_1203 (O_1203,N_14188,N_14542);
nor UO_1204 (O_1204,N_14434,N_13503);
or UO_1205 (O_1205,N_14916,N_14527);
or UO_1206 (O_1206,N_13526,N_14622);
and UO_1207 (O_1207,N_14627,N_14772);
xor UO_1208 (O_1208,N_14744,N_14444);
nand UO_1209 (O_1209,N_13662,N_14523);
nor UO_1210 (O_1210,N_14528,N_14558);
nor UO_1211 (O_1211,N_13993,N_14679);
and UO_1212 (O_1212,N_14567,N_14053);
and UO_1213 (O_1213,N_13538,N_14877);
nand UO_1214 (O_1214,N_13559,N_14992);
nand UO_1215 (O_1215,N_14841,N_14385);
nor UO_1216 (O_1216,N_14735,N_13819);
and UO_1217 (O_1217,N_13928,N_13597);
or UO_1218 (O_1218,N_14303,N_13847);
nand UO_1219 (O_1219,N_14991,N_14212);
or UO_1220 (O_1220,N_14771,N_13927);
nand UO_1221 (O_1221,N_14909,N_14258);
nor UO_1222 (O_1222,N_14296,N_13889);
and UO_1223 (O_1223,N_13573,N_14996);
or UO_1224 (O_1224,N_13504,N_13679);
xor UO_1225 (O_1225,N_13952,N_14243);
nand UO_1226 (O_1226,N_14616,N_14607);
and UO_1227 (O_1227,N_14628,N_14056);
or UO_1228 (O_1228,N_14680,N_13755);
nor UO_1229 (O_1229,N_14183,N_13696);
nand UO_1230 (O_1230,N_13968,N_14074);
nor UO_1231 (O_1231,N_14991,N_13882);
nor UO_1232 (O_1232,N_14782,N_14471);
nand UO_1233 (O_1233,N_13956,N_13775);
or UO_1234 (O_1234,N_14226,N_14040);
nand UO_1235 (O_1235,N_14327,N_13570);
nand UO_1236 (O_1236,N_14404,N_14171);
or UO_1237 (O_1237,N_13842,N_14705);
or UO_1238 (O_1238,N_13535,N_14928);
or UO_1239 (O_1239,N_13576,N_14349);
nand UO_1240 (O_1240,N_14039,N_14043);
nor UO_1241 (O_1241,N_13966,N_14824);
nor UO_1242 (O_1242,N_14537,N_14305);
and UO_1243 (O_1243,N_13903,N_14420);
nor UO_1244 (O_1244,N_14653,N_14089);
or UO_1245 (O_1245,N_14398,N_14694);
or UO_1246 (O_1246,N_14802,N_13694);
nor UO_1247 (O_1247,N_14390,N_14334);
and UO_1248 (O_1248,N_14073,N_13659);
nor UO_1249 (O_1249,N_13546,N_13834);
and UO_1250 (O_1250,N_13853,N_13566);
nor UO_1251 (O_1251,N_14249,N_14977);
or UO_1252 (O_1252,N_14253,N_14784);
or UO_1253 (O_1253,N_14094,N_14888);
and UO_1254 (O_1254,N_13776,N_13564);
and UO_1255 (O_1255,N_14648,N_14636);
or UO_1256 (O_1256,N_14485,N_14389);
nand UO_1257 (O_1257,N_14847,N_14917);
and UO_1258 (O_1258,N_14974,N_13646);
and UO_1259 (O_1259,N_13542,N_13662);
or UO_1260 (O_1260,N_14003,N_13883);
nor UO_1261 (O_1261,N_13738,N_14378);
nor UO_1262 (O_1262,N_13775,N_14285);
nor UO_1263 (O_1263,N_14933,N_14794);
nor UO_1264 (O_1264,N_14702,N_14893);
nor UO_1265 (O_1265,N_13981,N_13556);
or UO_1266 (O_1266,N_14978,N_13684);
or UO_1267 (O_1267,N_14164,N_14031);
and UO_1268 (O_1268,N_14340,N_14559);
or UO_1269 (O_1269,N_13564,N_14045);
and UO_1270 (O_1270,N_14944,N_14592);
and UO_1271 (O_1271,N_14403,N_14888);
or UO_1272 (O_1272,N_14172,N_13954);
xnor UO_1273 (O_1273,N_14952,N_14712);
nand UO_1274 (O_1274,N_14731,N_14912);
or UO_1275 (O_1275,N_13984,N_14884);
nand UO_1276 (O_1276,N_14556,N_14228);
nor UO_1277 (O_1277,N_13695,N_14589);
and UO_1278 (O_1278,N_13704,N_13820);
nor UO_1279 (O_1279,N_13565,N_14284);
nand UO_1280 (O_1280,N_14882,N_14565);
xor UO_1281 (O_1281,N_13870,N_13858);
nor UO_1282 (O_1282,N_14436,N_14636);
or UO_1283 (O_1283,N_13927,N_13712);
nor UO_1284 (O_1284,N_13743,N_14356);
nand UO_1285 (O_1285,N_14584,N_14755);
nand UO_1286 (O_1286,N_13658,N_14179);
and UO_1287 (O_1287,N_14084,N_14519);
and UO_1288 (O_1288,N_14326,N_13610);
nor UO_1289 (O_1289,N_14084,N_13524);
and UO_1290 (O_1290,N_13739,N_14473);
nand UO_1291 (O_1291,N_14644,N_13910);
and UO_1292 (O_1292,N_13664,N_14355);
and UO_1293 (O_1293,N_13740,N_14686);
nand UO_1294 (O_1294,N_13618,N_13693);
nand UO_1295 (O_1295,N_14115,N_14123);
nand UO_1296 (O_1296,N_14911,N_14815);
or UO_1297 (O_1297,N_13606,N_14542);
xor UO_1298 (O_1298,N_14318,N_13994);
and UO_1299 (O_1299,N_14285,N_14997);
nand UO_1300 (O_1300,N_14715,N_13623);
and UO_1301 (O_1301,N_14968,N_13785);
and UO_1302 (O_1302,N_13656,N_14366);
nor UO_1303 (O_1303,N_14381,N_13861);
or UO_1304 (O_1304,N_14875,N_14289);
nand UO_1305 (O_1305,N_13655,N_13772);
nor UO_1306 (O_1306,N_14651,N_14109);
or UO_1307 (O_1307,N_14427,N_14062);
and UO_1308 (O_1308,N_13689,N_14455);
and UO_1309 (O_1309,N_14070,N_14805);
or UO_1310 (O_1310,N_14487,N_14476);
and UO_1311 (O_1311,N_14034,N_14733);
nor UO_1312 (O_1312,N_13873,N_13845);
and UO_1313 (O_1313,N_13621,N_14138);
or UO_1314 (O_1314,N_14058,N_14836);
and UO_1315 (O_1315,N_13614,N_14077);
nor UO_1316 (O_1316,N_14624,N_13733);
xor UO_1317 (O_1317,N_14584,N_14678);
or UO_1318 (O_1318,N_14104,N_13544);
nand UO_1319 (O_1319,N_14651,N_14829);
or UO_1320 (O_1320,N_14829,N_14966);
nand UO_1321 (O_1321,N_13509,N_14791);
and UO_1322 (O_1322,N_14820,N_13741);
or UO_1323 (O_1323,N_14283,N_14654);
or UO_1324 (O_1324,N_14123,N_14473);
or UO_1325 (O_1325,N_14752,N_14419);
and UO_1326 (O_1326,N_14448,N_13897);
and UO_1327 (O_1327,N_14778,N_14613);
nor UO_1328 (O_1328,N_13618,N_14845);
nand UO_1329 (O_1329,N_13580,N_13948);
nand UO_1330 (O_1330,N_14068,N_13717);
or UO_1331 (O_1331,N_14900,N_13934);
nor UO_1332 (O_1332,N_13518,N_14335);
nand UO_1333 (O_1333,N_13996,N_14446);
or UO_1334 (O_1334,N_14826,N_14977);
and UO_1335 (O_1335,N_14984,N_14068);
nor UO_1336 (O_1336,N_14258,N_13895);
and UO_1337 (O_1337,N_13700,N_13550);
xnor UO_1338 (O_1338,N_13571,N_13954);
or UO_1339 (O_1339,N_14950,N_14002);
and UO_1340 (O_1340,N_14933,N_14580);
nand UO_1341 (O_1341,N_14041,N_13943);
and UO_1342 (O_1342,N_14511,N_14489);
or UO_1343 (O_1343,N_13751,N_13524);
nor UO_1344 (O_1344,N_13872,N_14833);
nor UO_1345 (O_1345,N_14012,N_14348);
and UO_1346 (O_1346,N_14773,N_14660);
and UO_1347 (O_1347,N_14707,N_14953);
nor UO_1348 (O_1348,N_14404,N_13799);
or UO_1349 (O_1349,N_14212,N_14533);
nor UO_1350 (O_1350,N_14368,N_13665);
nor UO_1351 (O_1351,N_13960,N_14398);
nand UO_1352 (O_1352,N_13944,N_13532);
and UO_1353 (O_1353,N_14123,N_14251);
nor UO_1354 (O_1354,N_13949,N_14584);
and UO_1355 (O_1355,N_14836,N_13509);
nand UO_1356 (O_1356,N_14277,N_14066);
and UO_1357 (O_1357,N_14258,N_14570);
nor UO_1358 (O_1358,N_13666,N_14526);
or UO_1359 (O_1359,N_14252,N_13646);
or UO_1360 (O_1360,N_14753,N_13893);
nor UO_1361 (O_1361,N_13643,N_14033);
nand UO_1362 (O_1362,N_14173,N_14071);
and UO_1363 (O_1363,N_14839,N_14119);
and UO_1364 (O_1364,N_14860,N_14862);
or UO_1365 (O_1365,N_13902,N_14399);
xnor UO_1366 (O_1366,N_14515,N_14634);
nor UO_1367 (O_1367,N_13720,N_13643);
nor UO_1368 (O_1368,N_13521,N_14829);
xnor UO_1369 (O_1369,N_14737,N_14353);
and UO_1370 (O_1370,N_14275,N_13702);
or UO_1371 (O_1371,N_14469,N_14215);
nand UO_1372 (O_1372,N_13713,N_14449);
nand UO_1373 (O_1373,N_14706,N_13989);
nand UO_1374 (O_1374,N_14514,N_14320);
or UO_1375 (O_1375,N_13790,N_13836);
and UO_1376 (O_1376,N_13540,N_13599);
nand UO_1377 (O_1377,N_14753,N_14280);
and UO_1378 (O_1378,N_13948,N_14536);
and UO_1379 (O_1379,N_13993,N_14375);
and UO_1380 (O_1380,N_13620,N_14706);
and UO_1381 (O_1381,N_13805,N_14735);
or UO_1382 (O_1382,N_13552,N_14766);
and UO_1383 (O_1383,N_13564,N_14646);
nand UO_1384 (O_1384,N_14162,N_14012);
nor UO_1385 (O_1385,N_14850,N_14430);
and UO_1386 (O_1386,N_14369,N_13970);
or UO_1387 (O_1387,N_13552,N_14337);
and UO_1388 (O_1388,N_14251,N_14356);
or UO_1389 (O_1389,N_14320,N_14403);
and UO_1390 (O_1390,N_14904,N_14260);
nor UO_1391 (O_1391,N_14106,N_14914);
or UO_1392 (O_1392,N_14032,N_13783);
and UO_1393 (O_1393,N_14287,N_14005);
nor UO_1394 (O_1394,N_14440,N_14248);
nand UO_1395 (O_1395,N_14486,N_14327);
and UO_1396 (O_1396,N_13563,N_13916);
and UO_1397 (O_1397,N_14968,N_13569);
or UO_1398 (O_1398,N_14683,N_13547);
and UO_1399 (O_1399,N_14478,N_13764);
and UO_1400 (O_1400,N_14879,N_14751);
or UO_1401 (O_1401,N_13781,N_14152);
nand UO_1402 (O_1402,N_14593,N_14296);
and UO_1403 (O_1403,N_13597,N_13839);
and UO_1404 (O_1404,N_14258,N_14844);
nor UO_1405 (O_1405,N_14185,N_14629);
nor UO_1406 (O_1406,N_14790,N_13671);
and UO_1407 (O_1407,N_14730,N_13775);
and UO_1408 (O_1408,N_14164,N_14639);
and UO_1409 (O_1409,N_13613,N_13842);
nor UO_1410 (O_1410,N_13878,N_14226);
nor UO_1411 (O_1411,N_14159,N_14496);
nor UO_1412 (O_1412,N_14310,N_14697);
nor UO_1413 (O_1413,N_14476,N_14389);
and UO_1414 (O_1414,N_13878,N_13627);
and UO_1415 (O_1415,N_14562,N_14695);
nor UO_1416 (O_1416,N_13522,N_14526);
nor UO_1417 (O_1417,N_13668,N_14673);
or UO_1418 (O_1418,N_14554,N_14068);
nand UO_1419 (O_1419,N_14983,N_14610);
nand UO_1420 (O_1420,N_14295,N_14358);
nand UO_1421 (O_1421,N_14585,N_13598);
nand UO_1422 (O_1422,N_13620,N_13829);
nand UO_1423 (O_1423,N_14968,N_14228);
and UO_1424 (O_1424,N_14274,N_14564);
xor UO_1425 (O_1425,N_14997,N_13828);
nor UO_1426 (O_1426,N_14053,N_14320);
nand UO_1427 (O_1427,N_13722,N_14325);
nand UO_1428 (O_1428,N_13761,N_14550);
or UO_1429 (O_1429,N_13905,N_14668);
and UO_1430 (O_1430,N_13504,N_14991);
nor UO_1431 (O_1431,N_14239,N_14110);
or UO_1432 (O_1432,N_14261,N_14118);
nor UO_1433 (O_1433,N_14069,N_14900);
or UO_1434 (O_1434,N_14211,N_14672);
or UO_1435 (O_1435,N_13539,N_14958);
nand UO_1436 (O_1436,N_14533,N_13784);
xnor UO_1437 (O_1437,N_13552,N_14907);
or UO_1438 (O_1438,N_13687,N_13693);
and UO_1439 (O_1439,N_13805,N_14809);
or UO_1440 (O_1440,N_14178,N_14212);
and UO_1441 (O_1441,N_14622,N_14204);
and UO_1442 (O_1442,N_13717,N_14646);
or UO_1443 (O_1443,N_14819,N_13715);
nand UO_1444 (O_1444,N_14520,N_14831);
and UO_1445 (O_1445,N_14147,N_14867);
and UO_1446 (O_1446,N_14704,N_14870);
nand UO_1447 (O_1447,N_14550,N_14088);
nand UO_1448 (O_1448,N_13856,N_13533);
xor UO_1449 (O_1449,N_14873,N_14586);
nor UO_1450 (O_1450,N_14950,N_14418);
and UO_1451 (O_1451,N_14056,N_14599);
and UO_1452 (O_1452,N_14745,N_13568);
nand UO_1453 (O_1453,N_14301,N_14660);
and UO_1454 (O_1454,N_13564,N_13758);
nand UO_1455 (O_1455,N_14471,N_14612);
or UO_1456 (O_1456,N_14535,N_14424);
nand UO_1457 (O_1457,N_14525,N_14163);
or UO_1458 (O_1458,N_14049,N_13819);
nor UO_1459 (O_1459,N_14414,N_14059);
or UO_1460 (O_1460,N_14232,N_13598);
or UO_1461 (O_1461,N_14937,N_13888);
nor UO_1462 (O_1462,N_13569,N_14987);
and UO_1463 (O_1463,N_14614,N_14280);
or UO_1464 (O_1464,N_13882,N_13657);
or UO_1465 (O_1465,N_13875,N_13633);
nand UO_1466 (O_1466,N_14424,N_14862);
nor UO_1467 (O_1467,N_13895,N_13773);
nor UO_1468 (O_1468,N_13774,N_13565);
nand UO_1469 (O_1469,N_14195,N_13995);
and UO_1470 (O_1470,N_14009,N_14177);
or UO_1471 (O_1471,N_14432,N_13867);
and UO_1472 (O_1472,N_14362,N_13516);
nand UO_1473 (O_1473,N_14578,N_13890);
xor UO_1474 (O_1474,N_14056,N_13657);
nor UO_1475 (O_1475,N_14360,N_14696);
nand UO_1476 (O_1476,N_14016,N_13849);
nand UO_1477 (O_1477,N_14244,N_14625);
or UO_1478 (O_1478,N_14187,N_14239);
and UO_1479 (O_1479,N_14220,N_14428);
nand UO_1480 (O_1480,N_14505,N_14080);
nand UO_1481 (O_1481,N_13608,N_13927);
or UO_1482 (O_1482,N_13579,N_14781);
nor UO_1483 (O_1483,N_13934,N_14515);
and UO_1484 (O_1484,N_13586,N_14412);
nand UO_1485 (O_1485,N_14335,N_14620);
nor UO_1486 (O_1486,N_14466,N_14888);
and UO_1487 (O_1487,N_14954,N_14175);
or UO_1488 (O_1488,N_13687,N_13853);
nand UO_1489 (O_1489,N_13705,N_14815);
nand UO_1490 (O_1490,N_14965,N_13554);
nand UO_1491 (O_1491,N_14633,N_14680);
nand UO_1492 (O_1492,N_13603,N_14764);
xor UO_1493 (O_1493,N_14928,N_14891);
nand UO_1494 (O_1494,N_13622,N_14800);
nand UO_1495 (O_1495,N_13969,N_14836);
or UO_1496 (O_1496,N_14108,N_13611);
or UO_1497 (O_1497,N_14834,N_13622);
or UO_1498 (O_1498,N_13600,N_14608);
or UO_1499 (O_1499,N_13826,N_14080);
and UO_1500 (O_1500,N_14561,N_14851);
nand UO_1501 (O_1501,N_14452,N_13598);
or UO_1502 (O_1502,N_14783,N_14057);
nand UO_1503 (O_1503,N_14875,N_13683);
or UO_1504 (O_1504,N_14261,N_14542);
nor UO_1505 (O_1505,N_14231,N_14623);
or UO_1506 (O_1506,N_13525,N_14423);
and UO_1507 (O_1507,N_14223,N_14968);
or UO_1508 (O_1508,N_14033,N_13920);
and UO_1509 (O_1509,N_13556,N_13555);
nor UO_1510 (O_1510,N_14136,N_14879);
nor UO_1511 (O_1511,N_14867,N_14720);
or UO_1512 (O_1512,N_13563,N_13705);
or UO_1513 (O_1513,N_14099,N_14226);
or UO_1514 (O_1514,N_14650,N_13705);
or UO_1515 (O_1515,N_13764,N_13995);
nor UO_1516 (O_1516,N_14135,N_14558);
and UO_1517 (O_1517,N_14805,N_14165);
nand UO_1518 (O_1518,N_14695,N_14541);
nor UO_1519 (O_1519,N_13603,N_14117);
or UO_1520 (O_1520,N_14844,N_13884);
and UO_1521 (O_1521,N_13695,N_13946);
and UO_1522 (O_1522,N_14750,N_14373);
or UO_1523 (O_1523,N_14520,N_14291);
and UO_1524 (O_1524,N_13892,N_14107);
nor UO_1525 (O_1525,N_14254,N_14214);
nand UO_1526 (O_1526,N_14076,N_14754);
nand UO_1527 (O_1527,N_13656,N_14975);
xor UO_1528 (O_1528,N_14127,N_13994);
or UO_1529 (O_1529,N_13864,N_14267);
and UO_1530 (O_1530,N_14292,N_13780);
or UO_1531 (O_1531,N_14182,N_14084);
nand UO_1532 (O_1532,N_14310,N_14408);
nand UO_1533 (O_1533,N_13821,N_13846);
nand UO_1534 (O_1534,N_14630,N_14860);
nor UO_1535 (O_1535,N_14556,N_13558);
and UO_1536 (O_1536,N_14825,N_13704);
nor UO_1537 (O_1537,N_13667,N_14475);
or UO_1538 (O_1538,N_14188,N_14901);
and UO_1539 (O_1539,N_14587,N_14288);
xnor UO_1540 (O_1540,N_13545,N_14545);
and UO_1541 (O_1541,N_14238,N_14109);
or UO_1542 (O_1542,N_13904,N_14367);
and UO_1543 (O_1543,N_14832,N_14459);
nand UO_1544 (O_1544,N_13651,N_14508);
or UO_1545 (O_1545,N_14210,N_13696);
nand UO_1546 (O_1546,N_14967,N_14085);
or UO_1547 (O_1547,N_14927,N_14363);
or UO_1548 (O_1548,N_14823,N_14705);
and UO_1549 (O_1549,N_14366,N_14219);
and UO_1550 (O_1550,N_14208,N_13896);
nor UO_1551 (O_1551,N_13751,N_13929);
or UO_1552 (O_1552,N_14585,N_14064);
or UO_1553 (O_1553,N_14736,N_14947);
nand UO_1554 (O_1554,N_14220,N_14242);
nand UO_1555 (O_1555,N_14275,N_13722);
xnor UO_1556 (O_1556,N_14209,N_13795);
nand UO_1557 (O_1557,N_14844,N_13662);
and UO_1558 (O_1558,N_14272,N_14341);
and UO_1559 (O_1559,N_13674,N_14405);
nor UO_1560 (O_1560,N_14715,N_14104);
nor UO_1561 (O_1561,N_14352,N_14642);
or UO_1562 (O_1562,N_14659,N_13601);
nor UO_1563 (O_1563,N_14192,N_14443);
nor UO_1564 (O_1564,N_14328,N_14344);
nor UO_1565 (O_1565,N_13649,N_14403);
nor UO_1566 (O_1566,N_13637,N_14521);
nand UO_1567 (O_1567,N_13948,N_14913);
or UO_1568 (O_1568,N_14065,N_14246);
nand UO_1569 (O_1569,N_13503,N_14546);
nor UO_1570 (O_1570,N_14392,N_14395);
and UO_1571 (O_1571,N_14818,N_14620);
nand UO_1572 (O_1572,N_14736,N_14087);
nand UO_1573 (O_1573,N_13775,N_14524);
nor UO_1574 (O_1574,N_14346,N_14236);
nor UO_1575 (O_1575,N_14201,N_13645);
nand UO_1576 (O_1576,N_13970,N_13770);
and UO_1577 (O_1577,N_14218,N_14925);
xnor UO_1578 (O_1578,N_13828,N_14954);
or UO_1579 (O_1579,N_14425,N_14919);
nand UO_1580 (O_1580,N_14602,N_13501);
nand UO_1581 (O_1581,N_14786,N_13756);
and UO_1582 (O_1582,N_13973,N_14799);
or UO_1583 (O_1583,N_13551,N_14409);
nand UO_1584 (O_1584,N_13537,N_14519);
nand UO_1585 (O_1585,N_14632,N_14800);
and UO_1586 (O_1586,N_14716,N_14409);
nor UO_1587 (O_1587,N_14309,N_13786);
nand UO_1588 (O_1588,N_14027,N_14414);
nor UO_1589 (O_1589,N_14700,N_14609);
nor UO_1590 (O_1590,N_14806,N_14846);
or UO_1591 (O_1591,N_13604,N_14236);
nor UO_1592 (O_1592,N_14769,N_14060);
and UO_1593 (O_1593,N_14873,N_14842);
nor UO_1594 (O_1594,N_13536,N_14537);
nor UO_1595 (O_1595,N_14260,N_14775);
or UO_1596 (O_1596,N_13752,N_14877);
and UO_1597 (O_1597,N_14190,N_13500);
and UO_1598 (O_1598,N_14140,N_13747);
and UO_1599 (O_1599,N_13975,N_13739);
nand UO_1600 (O_1600,N_14282,N_14201);
nand UO_1601 (O_1601,N_13941,N_14584);
nand UO_1602 (O_1602,N_14690,N_14020);
nand UO_1603 (O_1603,N_14432,N_14044);
or UO_1604 (O_1604,N_13918,N_14443);
or UO_1605 (O_1605,N_14442,N_14603);
nand UO_1606 (O_1606,N_14583,N_14121);
and UO_1607 (O_1607,N_14558,N_13952);
nand UO_1608 (O_1608,N_13606,N_14851);
nor UO_1609 (O_1609,N_14964,N_13668);
and UO_1610 (O_1610,N_14013,N_14267);
or UO_1611 (O_1611,N_13568,N_13736);
and UO_1612 (O_1612,N_14192,N_13520);
or UO_1613 (O_1613,N_14016,N_13868);
nor UO_1614 (O_1614,N_14355,N_14772);
nor UO_1615 (O_1615,N_13744,N_13714);
nand UO_1616 (O_1616,N_14951,N_14115);
and UO_1617 (O_1617,N_14853,N_14852);
or UO_1618 (O_1618,N_13605,N_13889);
nand UO_1619 (O_1619,N_14355,N_13649);
and UO_1620 (O_1620,N_13714,N_14992);
and UO_1621 (O_1621,N_13639,N_13699);
nand UO_1622 (O_1622,N_14252,N_14832);
or UO_1623 (O_1623,N_14496,N_14811);
and UO_1624 (O_1624,N_14444,N_13981);
nor UO_1625 (O_1625,N_14650,N_14051);
nand UO_1626 (O_1626,N_14831,N_14787);
or UO_1627 (O_1627,N_14355,N_14885);
or UO_1628 (O_1628,N_14549,N_14602);
or UO_1629 (O_1629,N_14961,N_13633);
nand UO_1630 (O_1630,N_14183,N_14054);
and UO_1631 (O_1631,N_14053,N_14623);
or UO_1632 (O_1632,N_14394,N_13739);
or UO_1633 (O_1633,N_14201,N_13732);
and UO_1634 (O_1634,N_13631,N_14370);
nor UO_1635 (O_1635,N_14802,N_13501);
nor UO_1636 (O_1636,N_13941,N_13928);
or UO_1637 (O_1637,N_14501,N_14300);
nand UO_1638 (O_1638,N_14687,N_13559);
and UO_1639 (O_1639,N_14849,N_14459);
xor UO_1640 (O_1640,N_14480,N_14548);
nor UO_1641 (O_1641,N_13802,N_13736);
nand UO_1642 (O_1642,N_13898,N_14574);
nor UO_1643 (O_1643,N_14112,N_13882);
and UO_1644 (O_1644,N_14841,N_13561);
and UO_1645 (O_1645,N_13897,N_14687);
nand UO_1646 (O_1646,N_14372,N_14978);
nor UO_1647 (O_1647,N_13933,N_14325);
or UO_1648 (O_1648,N_14129,N_13936);
and UO_1649 (O_1649,N_14335,N_14330);
or UO_1650 (O_1650,N_13555,N_14061);
or UO_1651 (O_1651,N_14596,N_14716);
and UO_1652 (O_1652,N_14961,N_14189);
nor UO_1653 (O_1653,N_14118,N_14793);
nand UO_1654 (O_1654,N_13753,N_14672);
or UO_1655 (O_1655,N_14731,N_14892);
nand UO_1656 (O_1656,N_14823,N_13585);
nor UO_1657 (O_1657,N_14259,N_14688);
or UO_1658 (O_1658,N_14770,N_13751);
nand UO_1659 (O_1659,N_14246,N_14721);
or UO_1660 (O_1660,N_14476,N_14844);
nand UO_1661 (O_1661,N_13823,N_14284);
nor UO_1662 (O_1662,N_14306,N_14847);
and UO_1663 (O_1663,N_14548,N_14406);
nor UO_1664 (O_1664,N_13544,N_14078);
nor UO_1665 (O_1665,N_14829,N_14825);
nor UO_1666 (O_1666,N_14869,N_14358);
or UO_1667 (O_1667,N_14026,N_14384);
and UO_1668 (O_1668,N_13894,N_14446);
xor UO_1669 (O_1669,N_13854,N_14477);
or UO_1670 (O_1670,N_14253,N_14940);
and UO_1671 (O_1671,N_14547,N_14424);
nor UO_1672 (O_1672,N_13651,N_14281);
or UO_1673 (O_1673,N_13754,N_14761);
nor UO_1674 (O_1674,N_14698,N_14766);
nand UO_1675 (O_1675,N_14366,N_14002);
nand UO_1676 (O_1676,N_14136,N_14057);
and UO_1677 (O_1677,N_13652,N_13642);
nor UO_1678 (O_1678,N_14153,N_14730);
nor UO_1679 (O_1679,N_13962,N_14975);
nor UO_1680 (O_1680,N_14305,N_14214);
nor UO_1681 (O_1681,N_14893,N_13935);
and UO_1682 (O_1682,N_13738,N_14567);
or UO_1683 (O_1683,N_13593,N_14623);
nor UO_1684 (O_1684,N_14744,N_14933);
nand UO_1685 (O_1685,N_13860,N_13778);
and UO_1686 (O_1686,N_14720,N_13794);
nand UO_1687 (O_1687,N_13787,N_14516);
or UO_1688 (O_1688,N_14125,N_14283);
and UO_1689 (O_1689,N_14866,N_13617);
nor UO_1690 (O_1690,N_14193,N_14209);
or UO_1691 (O_1691,N_13740,N_14363);
or UO_1692 (O_1692,N_14947,N_14863);
nand UO_1693 (O_1693,N_14065,N_13841);
nor UO_1694 (O_1694,N_14801,N_13996);
nand UO_1695 (O_1695,N_14396,N_14855);
and UO_1696 (O_1696,N_13777,N_13934);
nand UO_1697 (O_1697,N_14567,N_13551);
and UO_1698 (O_1698,N_14989,N_14799);
and UO_1699 (O_1699,N_14419,N_14987);
or UO_1700 (O_1700,N_13980,N_14485);
nand UO_1701 (O_1701,N_14585,N_13654);
nor UO_1702 (O_1702,N_13929,N_13599);
or UO_1703 (O_1703,N_14608,N_14255);
or UO_1704 (O_1704,N_14302,N_13516);
nor UO_1705 (O_1705,N_13868,N_14277);
nor UO_1706 (O_1706,N_14385,N_13568);
nor UO_1707 (O_1707,N_13523,N_14338);
and UO_1708 (O_1708,N_13828,N_14384);
nor UO_1709 (O_1709,N_14795,N_13724);
nor UO_1710 (O_1710,N_14897,N_13906);
nor UO_1711 (O_1711,N_14518,N_14316);
nor UO_1712 (O_1712,N_13887,N_14464);
nand UO_1713 (O_1713,N_13637,N_14635);
and UO_1714 (O_1714,N_14422,N_14960);
or UO_1715 (O_1715,N_14003,N_14316);
or UO_1716 (O_1716,N_13551,N_14443);
or UO_1717 (O_1717,N_14740,N_13820);
nor UO_1718 (O_1718,N_13954,N_13799);
nor UO_1719 (O_1719,N_14334,N_14256);
and UO_1720 (O_1720,N_13755,N_14882);
or UO_1721 (O_1721,N_13772,N_14562);
nor UO_1722 (O_1722,N_14664,N_14331);
or UO_1723 (O_1723,N_14871,N_14335);
nor UO_1724 (O_1724,N_14106,N_13850);
nor UO_1725 (O_1725,N_14230,N_13968);
xor UO_1726 (O_1726,N_14651,N_13561);
nor UO_1727 (O_1727,N_13696,N_13959);
nor UO_1728 (O_1728,N_14370,N_14478);
or UO_1729 (O_1729,N_14236,N_13983);
and UO_1730 (O_1730,N_13961,N_14684);
nor UO_1731 (O_1731,N_13678,N_14950);
or UO_1732 (O_1732,N_13675,N_14305);
nor UO_1733 (O_1733,N_14255,N_13534);
or UO_1734 (O_1734,N_14430,N_13918);
nand UO_1735 (O_1735,N_13578,N_14405);
nand UO_1736 (O_1736,N_13945,N_13910);
or UO_1737 (O_1737,N_13723,N_14376);
and UO_1738 (O_1738,N_13636,N_14481);
and UO_1739 (O_1739,N_14377,N_14387);
nand UO_1740 (O_1740,N_14450,N_14792);
nand UO_1741 (O_1741,N_14044,N_14542);
or UO_1742 (O_1742,N_13619,N_13841);
and UO_1743 (O_1743,N_14520,N_13794);
nand UO_1744 (O_1744,N_14518,N_13866);
nor UO_1745 (O_1745,N_13922,N_13950);
nor UO_1746 (O_1746,N_13612,N_14587);
or UO_1747 (O_1747,N_14287,N_14116);
nand UO_1748 (O_1748,N_14647,N_13963);
nor UO_1749 (O_1749,N_14072,N_13577);
nand UO_1750 (O_1750,N_14770,N_14492);
nand UO_1751 (O_1751,N_14381,N_14984);
nor UO_1752 (O_1752,N_14766,N_14287);
and UO_1753 (O_1753,N_13888,N_14019);
nand UO_1754 (O_1754,N_13566,N_13960);
nand UO_1755 (O_1755,N_14412,N_14651);
nand UO_1756 (O_1756,N_14458,N_13713);
and UO_1757 (O_1757,N_13697,N_14695);
or UO_1758 (O_1758,N_14731,N_13740);
and UO_1759 (O_1759,N_14526,N_14222);
nor UO_1760 (O_1760,N_13587,N_13645);
and UO_1761 (O_1761,N_14575,N_14430);
or UO_1762 (O_1762,N_14137,N_14558);
nor UO_1763 (O_1763,N_13699,N_14786);
and UO_1764 (O_1764,N_14863,N_14563);
or UO_1765 (O_1765,N_14766,N_14433);
nand UO_1766 (O_1766,N_14557,N_14758);
and UO_1767 (O_1767,N_13524,N_13667);
or UO_1768 (O_1768,N_14432,N_14499);
and UO_1769 (O_1769,N_14851,N_14096);
and UO_1770 (O_1770,N_14985,N_13600);
nor UO_1771 (O_1771,N_14062,N_14125);
nor UO_1772 (O_1772,N_14908,N_14918);
or UO_1773 (O_1773,N_13739,N_13659);
xor UO_1774 (O_1774,N_14020,N_13695);
nor UO_1775 (O_1775,N_14451,N_14900);
and UO_1776 (O_1776,N_14029,N_14951);
nand UO_1777 (O_1777,N_13627,N_13921);
or UO_1778 (O_1778,N_14020,N_14672);
and UO_1779 (O_1779,N_14446,N_14356);
or UO_1780 (O_1780,N_13898,N_14912);
nand UO_1781 (O_1781,N_14718,N_14076);
nand UO_1782 (O_1782,N_13596,N_13565);
xor UO_1783 (O_1783,N_14688,N_14701);
nand UO_1784 (O_1784,N_14823,N_14049);
or UO_1785 (O_1785,N_13957,N_14618);
or UO_1786 (O_1786,N_14775,N_13813);
nand UO_1787 (O_1787,N_14119,N_14738);
or UO_1788 (O_1788,N_14336,N_13829);
and UO_1789 (O_1789,N_13805,N_14953);
nand UO_1790 (O_1790,N_13756,N_14599);
nand UO_1791 (O_1791,N_14798,N_13977);
nor UO_1792 (O_1792,N_14541,N_14092);
nor UO_1793 (O_1793,N_14242,N_13782);
nand UO_1794 (O_1794,N_14072,N_13772);
nand UO_1795 (O_1795,N_13762,N_14638);
and UO_1796 (O_1796,N_13683,N_14530);
and UO_1797 (O_1797,N_13542,N_13540);
nor UO_1798 (O_1798,N_14062,N_14635);
and UO_1799 (O_1799,N_14628,N_13944);
or UO_1800 (O_1800,N_13661,N_13755);
or UO_1801 (O_1801,N_14991,N_13764);
and UO_1802 (O_1802,N_14400,N_14893);
nor UO_1803 (O_1803,N_14580,N_13549);
and UO_1804 (O_1804,N_14262,N_14065);
nand UO_1805 (O_1805,N_13507,N_13550);
or UO_1806 (O_1806,N_14004,N_14512);
nor UO_1807 (O_1807,N_14778,N_14283);
and UO_1808 (O_1808,N_13754,N_14545);
nor UO_1809 (O_1809,N_14794,N_14686);
and UO_1810 (O_1810,N_14333,N_14645);
nand UO_1811 (O_1811,N_13628,N_14835);
nor UO_1812 (O_1812,N_14332,N_14598);
or UO_1813 (O_1813,N_14230,N_14582);
nor UO_1814 (O_1814,N_13547,N_13531);
and UO_1815 (O_1815,N_13666,N_14826);
and UO_1816 (O_1816,N_14045,N_14597);
nand UO_1817 (O_1817,N_14448,N_13933);
and UO_1818 (O_1818,N_14625,N_13546);
and UO_1819 (O_1819,N_14435,N_13740);
and UO_1820 (O_1820,N_14301,N_13854);
nor UO_1821 (O_1821,N_14988,N_13574);
nand UO_1822 (O_1822,N_14348,N_14682);
nor UO_1823 (O_1823,N_13798,N_13795);
nor UO_1824 (O_1824,N_14518,N_14310);
nor UO_1825 (O_1825,N_14511,N_13989);
and UO_1826 (O_1826,N_13664,N_13913);
and UO_1827 (O_1827,N_13518,N_14425);
and UO_1828 (O_1828,N_13884,N_13998);
nor UO_1829 (O_1829,N_14866,N_14310);
and UO_1830 (O_1830,N_13516,N_14640);
nor UO_1831 (O_1831,N_13514,N_14112);
nor UO_1832 (O_1832,N_14037,N_13761);
nand UO_1833 (O_1833,N_14287,N_14991);
and UO_1834 (O_1834,N_14898,N_13615);
nand UO_1835 (O_1835,N_13658,N_13703);
and UO_1836 (O_1836,N_13948,N_13927);
and UO_1837 (O_1837,N_14858,N_14563);
nor UO_1838 (O_1838,N_14826,N_13517);
and UO_1839 (O_1839,N_14971,N_13573);
and UO_1840 (O_1840,N_14802,N_14091);
nand UO_1841 (O_1841,N_13956,N_14299);
or UO_1842 (O_1842,N_14450,N_14692);
and UO_1843 (O_1843,N_14247,N_14419);
and UO_1844 (O_1844,N_13951,N_14076);
and UO_1845 (O_1845,N_13550,N_13674);
nand UO_1846 (O_1846,N_13824,N_13649);
nand UO_1847 (O_1847,N_13952,N_13950);
nor UO_1848 (O_1848,N_14872,N_13665);
nand UO_1849 (O_1849,N_14924,N_13606);
nor UO_1850 (O_1850,N_13648,N_14148);
and UO_1851 (O_1851,N_14198,N_13695);
or UO_1852 (O_1852,N_13623,N_14184);
or UO_1853 (O_1853,N_14835,N_13847);
or UO_1854 (O_1854,N_14175,N_14220);
or UO_1855 (O_1855,N_13751,N_13932);
nand UO_1856 (O_1856,N_14340,N_14265);
and UO_1857 (O_1857,N_13837,N_14069);
nor UO_1858 (O_1858,N_14913,N_14841);
nand UO_1859 (O_1859,N_14764,N_14664);
nor UO_1860 (O_1860,N_14482,N_13896);
or UO_1861 (O_1861,N_14925,N_14538);
or UO_1862 (O_1862,N_13798,N_13891);
or UO_1863 (O_1863,N_14183,N_14768);
and UO_1864 (O_1864,N_14756,N_14395);
nor UO_1865 (O_1865,N_13534,N_14058);
and UO_1866 (O_1866,N_13588,N_14403);
or UO_1867 (O_1867,N_14642,N_13982);
nand UO_1868 (O_1868,N_14586,N_14242);
nor UO_1869 (O_1869,N_13809,N_14222);
nor UO_1870 (O_1870,N_14514,N_13578);
and UO_1871 (O_1871,N_13742,N_14470);
nand UO_1872 (O_1872,N_13574,N_14673);
nand UO_1873 (O_1873,N_14284,N_14971);
or UO_1874 (O_1874,N_14606,N_14556);
and UO_1875 (O_1875,N_14635,N_14016);
or UO_1876 (O_1876,N_14564,N_14324);
nor UO_1877 (O_1877,N_14039,N_14795);
nor UO_1878 (O_1878,N_14685,N_13605);
nor UO_1879 (O_1879,N_14710,N_13572);
or UO_1880 (O_1880,N_14118,N_14696);
or UO_1881 (O_1881,N_13630,N_14958);
nand UO_1882 (O_1882,N_13516,N_14335);
and UO_1883 (O_1883,N_13701,N_14458);
nor UO_1884 (O_1884,N_13531,N_14311);
nor UO_1885 (O_1885,N_14893,N_14583);
and UO_1886 (O_1886,N_14527,N_13842);
nand UO_1887 (O_1887,N_14522,N_14688);
and UO_1888 (O_1888,N_13732,N_14334);
and UO_1889 (O_1889,N_13816,N_14259);
and UO_1890 (O_1890,N_14592,N_14175);
nor UO_1891 (O_1891,N_14662,N_14352);
or UO_1892 (O_1892,N_14918,N_14301);
nand UO_1893 (O_1893,N_14820,N_14885);
nand UO_1894 (O_1894,N_14399,N_14734);
or UO_1895 (O_1895,N_14492,N_14521);
and UO_1896 (O_1896,N_14359,N_14190);
or UO_1897 (O_1897,N_13822,N_14502);
or UO_1898 (O_1898,N_14243,N_14489);
nand UO_1899 (O_1899,N_13621,N_13751);
and UO_1900 (O_1900,N_13972,N_14936);
and UO_1901 (O_1901,N_13890,N_13853);
nor UO_1902 (O_1902,N_13876,N_14910);
and UO_1903 (O_1903,N_14695,N_14713);
nor UO_1904 (O_1904,N_14978,N_14737);
or UO_1905 (O_1905,N_14801,N_14009);
and UO_1906 (O_1906,N_14655,N_13734);
nand UO_1907 (O_1907,N_13936,N_13649);
nor UO_1908 (O_1908,N_14666,N_14652);
nand UO_1909 (O_1909,N_14806,N_14761);
nor UO_1910 (O_1910,N_14784,N_14771);
and UO_1911 (O_1911,N_14132,N_14452);
and UO_1912 (O_1912,N_13653,N_14927);
nor UO_1913 (O_1913,N_14322,N_13610);
and UO_1914 (O_1914,N_14795,N_14350);
or UO_1915 (O_1915,N_14411,N_14374);
nor UO_1916 (O_1916,N_14613,N_13944);
and UO_1917 (O_1917,N_14498,N_14836);
or UO_1918 (O_1918,N_14236,N_14722);
or UO_1919 (O_1919,N_14309,N_14620);
or UO_1920 (O_1920,N_14792,N_13627);
nor UO_1921 (O_1921,N_14274,N_13827);
nor UO_1922 (O_1922,N_14080,N_13946);
nand UO_1923 (O_1923,N_14333,N_14452);
nand UO_1924 (O_1924,N_14728,N_13834);
nor UO_1925 (O_1925,N_14820,N_14752);
nand UO_1926 (O_1926,N_13798,N_14825);
nand UO_1927 (O_1927,N_13709,N_13814);
nor UO_1928 (O_1928,N_14718,N_14390);
or UO_1929 (O_1929,N_14257,N_13636);
and UO_1930 (O_1930,N_14759,N_14891);
or UO_1931 (O_1931,N_13780,N_13809);
nor UO_1932 (O_1932,N_14150,N_14166);
nor UO_1933 (O_1933,N_14005,N_13721);
nor UO_1934 (O_1934,N_14218,N_14526);
nor UO_1935 (O_1935,N_14042,N_14296);
nor UO_1936 (O_1936,N_13660,N_13616);
xor UO_1937 (O_1937,N_14832,N_14815);
nand UO_1938 (O_1938,N_14530,N_14116);
or UO_1939 (O_1939,N_14351,N_13760);
or UO_1940 (O_1940,N_14533,N_14443);
nor UO_1941 (O_1941,N_14189,N_13554);
nand UO_1942 (O_1942,N_14317,N_14716);
nand UO_1943 (O_1943,N_14498,N_13501);
nor UO_1944 (O_1944,N_13758,N_14693);
nand UO_1945 (O_1945,N_14655,N_13600);
or UO_1946 (O_1946,N_14418,N_13859);
nand UO_1947 (O_1947,N_14213,N_14228);
and UO_1948 (O_1948,N_13750,N_13685);
and UO_1949 (O_1949,N_14383,N_14781);
nand UO_1950 (O_1950,N_13724,N_14476);
and UO_1951 (O_1951,N_13827,N_14293);
and UO_1952 (O_1952,N_14834,N_14628);
and UO_1953 (O_1953,N_14077,N_13643);
nand UO_1954 (O_1954,N_13537,N_14205);
nand UO_1955 (O_1955,N_13562,N_13643);
and UO_1956 (O_1956,N_14936,N_14955);
or UO_1957 (O_1957,N_14356,N_14083);
or UO_1958 (O_1958,N_14208,N_14397);
or UO_1959 (O_1959,N_14318,N_13942);
and UO_1960 (O_1960,N_13556,N_14995);
nor UO_1961 (O_1961,N_14277,N_14620);
nand UO_1962 (O_1962,N_14292,N_14068);
nand UO_1963 (O_1963,N_13909,N_13579);
or UO_1964 (O_1964,N_14529,N_14181);
nor UO_1965 (O_1965,N_14406,N_14485);
nor UO_1966 (O_1966,N_14700,N_14546);
and UO_1967 (O_1967,N_13878,N_14405);
and UO_1968 (O_1968,N_14367,N_14535);
and UO_1969 (O_1969,N_14947,N_14987);
nand UO_1970 (O_1970,N_13981,N_13670);
nor UO_1971 (O_1971,N_13731,N_14244);
nand UO_1972 (O_1972,N_13706,N_13519);
nand UO_1973 (O_1973,N_13868,N_14645);
or UO_1974 (O_1974,N_13555,N_14269);
nand UO_1975 (O_1975,N_14006,N_13895);
or UO_1976 (O_1976,N_13947,N_13958);
nor UO_1977 (O_1977,N_14448,N_14872);
nand UO_1978 (O_1978,N_14223,N_14419);
and UO_1979 (O_1979,N_13693,N_14796);
nand UO_1980 (O_1980,N_13829,N_14492);
nand UO_1981 (O_1981,N_14829,N_14157);
and UO_1982 (O_1982,N_13939,N_14233);
nand UO_1983 (O_1983,N_13607,N_14169);
or UO_1984 (O_1984,N_13835,N_13504);
and UO_1985 (O_1985,N_14656,N_14319);
and UO_1986 (O_1986,N_14796,N_13934);
nor UO_1987 (O_1987,N_13563,N_14315);
and UO_1988 (O_1988,N_14800,N_13629);
and UO_1989 (O_1989,N_13916,N_14607);
nand UO_1990 (O_1990,N_14054,N_14397);
nand UO_1991 (O_1991,N_14140,N_13749);
nor UO_1992 (O_1992,N_14525,N_14035);
nor UO_1993 (O_1993,N_13592,N_14715);
nand UO_1994 (O_1994,N_14184,N_13990);
or UO_1995 (O_1995,N_14775,N_14515);
nor UO_1996 (O_1996,N_14680,N_14955);
or UO_1997 (O_1997,N_14566,N_14391);
or UO_1998 (O_1998,N_14151,N_13593);
nor UO_1999 (O_1999,N_13810,N_14675);
endmodule