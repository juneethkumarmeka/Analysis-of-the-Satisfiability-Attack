module basic_1000_10000_1500_100_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xnor U0 (N_0,In_547,In_101);
or U1 (N_1,In_628,In_518);
and U2 (N_2,In_617,In_239);
nor U3 (N_3,In_115,In_368);
xor U4 (N_4,In_489,In_873);
xor U5 (N_5,In_701,In_645);
and U6 (N_6,In_844,In_269);
xnor U7 (N_7,In_108,In_236);
or U8 (N_8,In_98,In_987);
or U9 (N_9,In_459,In_960);
and U10 (N_10,In_978,In_143);
nor U11 (N_11,In_800,In_726);
nor U12 (N_12,In_83,In_404);
and U13 (N_13,In_118,In_572);
xor U14 (N_14,In_362,In_832);
nor U15 (N_15,In_158,In_126);
xor U16 (N_16,In_980,In_897);
xor U17 (N_17,In_136,In_743);
xnor U18 (N_18,In_24,In_3);
nand U19 (N_19,In_623,In_846);
or U20 (N_20,In_807,In_263);
nand U21 (N_21,In_984,In_552);
nand U22 (N_22,In_251,In_287);
or U23 (N_23,In_353,In_198);
or U24 (N_24,In_439,In_721);
nand U25 (N_25,In_720,In_478);
nand U26 (N_26,In_218,In_612);
and U27 (N_27,In_438,In_719);
nand U28 (N_28,In_773,In_659);
xnor U29 (N_29,In_190,In_149);
nor U30 (N_30,In_60,In_513);
or U31 (N_31,In_138,In_293);
xor U32 (N_32,In_63,In_970);
or U33 (N_33,In_423,In_44);
nor U34 (N_34,In_7,In_982);
nand U35 (N_35,In_804,In_341);
nor U36 (N_36,In_646,In_966);
nor U37 (N_37,In_21,In_315);
and U38 (N_38,In_576,In_298);
and U39 (N_39,In_699,In_457);
xor U40 (N_40,In_858,In_34);
or U41 (N_41,In_562,In_429);
nand U42 (N_42,In_90,In_245);
nand U43 (N_43,In_910,In_309);
and U44 (N_44,In_6,In_450);
and U45 (N_45,In_510,In_506);
or U46 (N_46,In_401,In_557);
and U47 (N_47,In_172,In_446);
xnor U48 (N_48,In_692,In_884);
or U49 (N_49,In_548,In_267);
or U50 (N_50,In_161,In_246);
and U51 (N_51,In_964,In_345);
nand U52 (N_52,In_586,In_453);
nand U53 (N_53,In_840,In_210);
xnor U54 (N_54,In_393,In_607);
or U55 (N_55,In_878,In_26);
xor U56 (N_56,In_225,In_979);
nand U57 (N_57,In_75,In_913);
nand U58 (N_58,In_31,In_906);
or U59 (N_59,In_886,In_215);
and U60 (N_60,In_93,In_327);
nor U61 (N_61,In_183,In_312);
or U62 (N_62,In_94,In_969);
nor U63 (N_63,In_658,In_512);
nand U64 (N_64,In_498,In_428);
nand U65 (N_65,In_473,In_334);
or U66 (N_66,In_110,In_655);
nand U67 (N_67,In_124,In_823);
xor U68 (N_68,In_988,In_780);
nand U69 (N_69,In_10,In_322);
or U70 (N_70,In_524,In_189);
xor U71 (N_71,In_113,In_733);
or U72 (N_72,In_555,In_741);
nand U73 (N_73,In_575,In_276);
or U74 (N_74,In_656,In_326);
or U75 (N_75,In_717,In_590);
nand U76 (N_76,In_983,In_615);
nor U77 (N_77,In_11,In_782);
and U78 (N_78,In_357,In_783);
nor U79 (N_79,In_205,In_131);
nor U80 (N_80,In_197,In_170);
xor U81 (N_81,In_504,In_471);
nor U82 (N_82,In_916,In_998);
nand U83 (N_83,In_544,In_254);
nor U84 (N_84,In_712,In_523);
and U85 (N_85,In_468,In_714);
xor U86 (N_86,In_372,In_616);
nand U87 (N_87,In_542,In_929);
or U88 (N_88,In_204,In_355);
or U89 (N_89,In_593,In_290);
and U90 (N_90,In_687,In_891);
xor U91 (N_91,In_65,In_601);
nand U92 (N_92,In_705,In_281);
nand U93 (N_93,In_902,In_361);
and U94 (N_94,In_738,In_529);
or U95 (N_95,In_957,In_45);
nand U96 (N_96,In_61,In_303);
nand U97 (N_97,In_127,In_255);
xor U98 (N_98,In_454,In_222);
nor U99 (N_99,In_316,In_793);
nor U100 (N_100,In_975,In_487);
and U101 (N_101,In_639,In_449);
and U102 (N_102,In_962,In_117);
or U103 (N_103,In_624,In_569);
nor U104 (N_104,In_179,In_820);
or U105 (N_105,In_107,In_688);
nor U106 (N_106,In_261,N_40);
or U107 (N_107,In_443,In_648);
or U108 (N_108,In_409,In_839);
xor U109 (N_109,In_981,N_35);
and U110 (N_110,In_908,In_845);
nor U111 (N_111,In_650,In_541);
xor U112 (N_112,In_411,In_427);
and U113 (N_113,In_585,N_66);
nand U114 (N_114,In_20,In_321);
nand U115 (N_115,In_802,In_396);
xor U116 (N_116,In_495,In_715);
nand U117 (N_117,In_491,In_896);
nor U118 (N_118,In_379,In_336);
nor U119 (N_119,N_71,In_208);
xor U120 (N_120,In_815,In_652);
and U121 (N_121,In_14,In_168);
nor U122 (N_122,In_386,In_794);
and U123 (N_123,In_647,In_381);
nand U124 (N_124,In_348,In_243);
nor U125 (N_125,In_852,In_671);
nor U126 (N_126,In_220,In_199);
and U127 (N_127,In_619,In_860);
nand U128 (N_128,In_235,In_458);
and U129 (N_129,In_389,In_344);
xor U130 (N_130,In_193,In_85);
xor U131 (N_131,In_436,In_514);
and U132 (N_132,In_664,In_425);
xnor U133 (N_133,In_856,In_649);
xor U134 (N_134,In_200,In_503);
and U135 (N_135,In_167,In_119);
nor U136 (N_136,In_613,In_812);
xor U137 (N_137,In_776,In_231);
nor U138 (N_138,In_36,In_365);
xor U139 (N_139,In_475,In_260);
or U140 (N_140,In_242,In_638);
nand U141 (N_141,In_564,In_917);
nor U142 (N_142,In_660,N_34);
and U143 (N_143,In_317,In_795);
xnor U144 (N_144,In_227,In_69);
nor U145 (N_145,In_734,In_599);
nand U146 (N_146,In_570,In_670);
and U147 (N_147,In_567,In_892);
nor U148 (N_148,In_736,In_333);
xor U149 (N_149,N_11,In_100);
or U150 (N_150,In_105,In_875);
xnor U151 (N_151,In_967,N_7);
xnor U152 (N_152,In_434,In_870);
nor U153 (N_153,In_855,In_111);
or U154 (N_154,In_497,N_25);
and U155 (N_155,In_191,In_250);
xor U156 (N_156,In_907,N_13);
nor U157 (N_157,In_538,In_256);
nor U158 (N_158,In_784,In_87);
and U159 (N_159,In_696,In_716);
nand U160 (N_160,In_604,In_84);
nand U161 (N_161,In_12,In_201);
nand U162 (N_162,N_6,In_171);
nor U163 (N_163,In_889,In_431);
xnor U164 (N_164,In_597,In_632);
nand U165 (N_165,In_676,N_68);
xnor U166 (N_166,In_626,In_801);
nor U167 (N_167,In_826,In_257);
xnor U168 (N_168,In_850,In_950);
xor U169 (N_169,In_869,In_702);
xor U170 (N_170,In_445,In_730);
xor U171 (N_171,In_943,In_887);
or U172 (N_172,In_834,In_451);
or U173 (N_173,In_992,In_880);
nand U174 (N_174,In_787,In_195);
nand U175 (N_175,In_440,In_781);
xor U176 (N_176,In_744,In_37);
nor U177 (N_177,In_678,In_694);
or U178 (N_178,In_206,In_965);
xnor U179 (N_179,N_21,In_358);
xor U180 (N_180,In_921,In_359);
nand U181 (N_181,In_876,In_686);
nand U182 (N_182,In_857,N_85);
or U183 (N_183,In_92,In_247);
and U184 (N_184,In_419,In_349);
or U185 (N_185,In_866,N_42);
xor U186 (N_186,In_877,N_77);
or U187 (N_187,In_882,In_811);
nor U188 (N_188,In_739,In_174);
xnor U189 (N_189,In_18,In_539);
nor U190 (N_190,In_212,In_278);
or U191 (N_191,N_22,In_282);
xor U192 (N_192,In_797,In_494);
nor U193 (N_193,In_102,In_621);
nor U194 (N_194,In_605,N_46);
or U195 (N_195,In_81,In_872);
and U196 (N_196,N_55,In_972);
or U197 (N_197,In_297,N_1);
nor U198 (N_198,N_9,In_728);
and U199 (N_199,In_849,In_229);
nand U200 (N_200,N_60,In_825);
and U201 (N_201,In_292,In_788);
nand U202 (N_202,In_827,N_123);
and U203 (N_203,In_634,In_582);
nand U204 (N_204,In_153,In_184);
or U205 (N_205,In_633,In_29);
nand U206 (N_206,N_157,N_81);
nand U207 (N_207,N_173,In_620);
xnor U208 (N_208,In_163,In_233);
or U209 (N_209,N_10,N_50);
xor U210 (N_210,In_583,N_105);
xor U211 (N_211,N_30,In_596);
nor U212 (N_212,In_25,N_143);
nor U213 (N_213,N_181,N_197);
and U214 (N_214,In_690,In_435);
nand U215 (N_215,In_155,N_101);
nand U216 (N_216,In_196,In_919);
and U217 (N_217,In_335,N_193);
or U218 (N_218,In_337,In_517);
or U219 (N_219,In_841,In_456);
nor U220 (N_220,In_240,In_40);
nand U221 (N_221,In_611,In_809);
nand U222 (N_222,In_843,In_299);
nor U223 (N_223,In_927,In_133);
and U224 (N_224,In_30,In_38);
and U225 (N_225,N_147,In_816);
nor U226 (N_226,In_937,In_608);
nor U227 (N_227,In_234,In_627);
nor U228 (N_228,In_813,In_684);
xnor U229 (N_229,In_757,N_52);
nor U230 (N_230,N_45,In_618);
or U231 (N_231,In_47,N_114);
nand U232 (N_232,In_22,In_96);
or U233 (N_233,In_178,In_864);
or U234 (N_234,In_779,N_73);
or U235 (N_235,In_4,N_103);
xor U236 (N_236,N_171,In_681);
nand U237 (N_237,N_29,N_169);
nor U238 (N_238,In_519,N_106);
xnor U239 (N_239,In_526,N_5);
nor U240 (N_240,In_437,In_244);
and U241 (N_241,In_534,In_42);
nand U242 (N_242,In_679,In_275);
or U243 (N_243,In_56,N_70);
nor U244 (N_244,In_669,In_977);
xor U245 (N_245,N_18,In_173);
nand U246 (N_246,In_151,In_499);
xor U247 (N_247,In_219,In_66);
and U248 (N_248,In_755,In_375);
or U249 (N_249,In_176,In_675);
nor U250 (N_250,In_477,In_713);
xnor U251 (N_251,In_637,In_367);
nand U252 (N_252,N_140,N_44);
or U253 (N_253,In_595,In_835);
and U254 (N_254,In_46,In_123);
xor U255 (N_255,In_904,N_14);
and U256 (N_256,In_121,N_59);
or U257 (N_257,In_806,In_936);
nand U258 (N_258,In_563,In_141);
or U259 (N_259,N_154,In_848);
or U260 (N_260,In_48,In_180);
nand U261 (N_261,In_695,N_112);
and U262 (N_262,In_948,In_577);
nand U263 (N_263,In_796,In_320);
nor U264 (N_264,In_533,N_74);
nor U265 (N_265,In_328,In_901);
or U266 (N_266,In_528,N_134);
or U267 (N_267,In_640,N_145);
and U268 (N_268,In_752,In_338);
nor U269 (N_269,N_89,In_974);
nand U270 (N_270,N_116,N_167);
nor U271 (N_271,In_600,In_385);
xor U272 (N_272,N_113,N_175);
xor U273 (N_273,N_98,In_828);
nor U274 (N_274,In_397,In_441);
or U275 (N_275,In_481,In_955);
or U276 (N_276,In_631,In_709);
xnor U277 (N_277,N_130,In_516);
or U278 (N_278,N_63,In_76);
xor U279 (N_279,In_708,N_176);
xor U280 (N_280,In_486,In_476);
or U281 (N_281,In_665,In_560);
and U282 (N_282,In_762,In_308);
or U283 (N_283,In_405,In_697);
and U284 (N_284,N_164,In_824);
or U285 (N_285,In_636,In_13);
xor U286 (N_286,In_853,In_408);
xor U287 (N_287,N_24,In_280);
nor U288 (N_288,In_16,N_41);
xor U289 (N_289,In_448,In_112);
nand U290 (N_290,In_579,In_581);
nor U291 (N_291,In_395,In_758);
xnor U292 (N_292,In_963,In_915);
xor U293 (N_293,N_62,In_883);
and U294 (N_294,In_41,In_485);
and U295 (N_295,N_39,In_224);
nor U296 (N_296,In_214,In_894);
or U297 (N_297,N_141,In_403);
xor U298 (N_298,In_422,In_677);
nand U299 (N_299,N_115,In_145);
xor U300 (N_300,N_137,N_295);
and U301 (N_301,In_294,In_706);
and U302 (N_302,In_460,In_890);
and U303 (N_303,In_213,N_159);
or U304 (N_304,In_323,N_102);
or U305 (N_305,N_110,In_469);
nor U306 (N_306,N_174,In_867);
nand U307 (N_307,N_67,In_556);
nand U308 (N_308,In_52,In_27);
nand U309 (N_309,In_767,In_32);
nand U310 (N_310,In_142,In_62);
xor U311 (N_311,N_17,In_945);
nor U312 (N_312,N_119,In_868);
and U313 (N_313,In_470,In_680);
nor U314 (N_314,In_833,N_156);
nor U315 (N_315,In_302,In_914);
or U316 (N_316,N_88,In_685);
nand U317 (N_317,N_87,In_188);
nor U318 (N_318,In_511,N_278);
nand U319 (N_319,In_314,In_594);
nor U320 (N_320,In_509,In_947);
or U321 (N_321,In_573,In_33);
and U322 (N_322,In_759,N_144);
xnor U323 (N_323,In_426,In_953);
nand U324 (N_324,In_58,In_566);
xor U325 (N_325,In_433,N_139);
xnor U326 (N_326,In_424,In_792);
xor U327 (N_327,In_933,In_296);
xor U328 (N_328,N_3,In_985);
nor U329 (N_329,In_159,In_905);
and U330 (N_330,N_75,N_200);
or U331 (N_331,In_331,In_472);
nand U332 (N_332,N_65,In_881);
or U333 (N_333,In_530,In_249);
nor U334 (N_334,In_598,N_244);
and U335 (N_335,In_270,In_641);
and U336 (N_336,In_88,N_268);
and U337 (N_337,N_121,In_392);
and U338 (N_338,In_162,In_462);
xnor U339 (N_339,N_257,In_842);
or U340 (N_340,N_228,In_996);
xnor U341 (N_341,In_775,In_382);
nand U342 (N_342,N_93,In_536);
or U343 (N_343,In_146,N_151);
nand U344 (N_344,N_216,In_653);
nand U345 (N_345,N_31,In_925);
and U346 (N_346,N_72,N_4);
or U347 (N_347,In_939,N_294);
xnor U348 (N_348,In_373,In_324);
or U349 (N_349,In_406,In_148);
and U350 (N_350,N_222,In_588);
nor U351 (N_351,In_991,In_300);
and U352 (N_352,In_537,In_674);
nand U353 (N_353,In_54,In_207);
xor U354 (N_354,In_383,In_387);
nand U355 (N_355,In_463,N_124);
and U356 (N_356,In_415,In_761);
or U357 (N_357,N_56,In_666);
nor U358 (N_358,N_36,In_798);
xor U359 (N_359,In_374,N_108);
xnor U360 (N_360,In_430,In_543);
and U361 (N_361,N_220,N_272);
xnor U362 (N_362,N_275,N_165);
or U363 (N_363,In_942,N_249);
or U364 (N_364,In_932,In_753);
and U365 (N_365,N_43,N_199);
or U366 (N_366,In_305,In_343);
and U367 (N_367,N_210,N_152);
nand U368 (N_368,In_252,N_195);
nand U369 (N_369,In_625,In_642);
and U370 (N_370,In_301,In_727);
nand U371 (N_371,In_663,In_279);
nor U372 (N_372,In_59,In_271);
nor U373 (N_373,In_103,In_703);
or U374 (N_374,N_86,In_522);
and U375 (N_375,N_289,In_754);
nand U376 (N_376,In_230,In_73);
or U377 (N_377,N_276,In_493);
nand U378 (N_378,N_239,In_691);
nand U379 (N_379,In_95,In_574);
nand U380 (N_380,N_162,In_922);
xor U381 (N_381,N_256,In_99);
nand U382 (N_382,In_920,In_421);
nor U383 (N_383,In_893,In_924);
and U384 (N_384,In_187,N_133);
xor U385 (N_385,N_205,N_97);
or U386 (N_386,In_371,In_89);
and U387 (N_387,In_157,N_179);
nor U388 (N_388,In_432,In_8);
or U389 (N_389,In_217,In_186);
and U390 (N_390,In_352,In_474);
or U391 (N_391,N_260,In_558);
nor U392 (N_392,N_263,N_187);
nand U393 (N_393,In_662,In_228);
or U394 (N_394,N_182,In_185);
and U395 (N_395,In_209,In_226);
xnor U396 (N_396,In_837,In_350);
and U397 (N_397,In_53,In_550);
and U398 (N_398,N_279,In_160);
and U399 (N_399,In_750,N_207);
and U400 (N_400,In_49,In_546);
xnor U401 (N_401,In_976,N_325);
nand U402 (N_402,In_938,N_381);
and U403 (N_403,N_226,In_629);
and U404 (N_404,N_300,In_861);
nand U405 (N_405,N_365,In_407);
xor U406 (N_406,In_725,In_283);
nand U407 (N_407,In_805,In_378);
nand U408 (N_408,N_53,N_240);
or U409 (N_409,N_364,In_268);
nor U410 (N_410,In_508,In_584);
xnor U411 (N_411,In_384,In_952);
nor U412 (N_412,N_183,N_32);
nor U413 (N_413,In_64,In_307);
xnor U414 (N_414,In_930,In_748);
and U415 (N_415,N_255,In_718);
xnor U416 (N_416,In_909,N_201);
xor U417 (N_417,N_76,N_211);
and U418 (N_418,In_580,In_635);
nand U419 (N_419,In_956,In_551);
nor U420 (N_420,In_192,In_139);
and U421 (N_421,In_729,N_192);
nor U422 (N_422,In_768,N_8);
and U423 (N_423,In_763,N_221);
nand U424 (N_424,In_990,In_496);
xor U425 (N_425,N_266,N_83);
and U426 (N_426,In_760,N_131);
xor U427 (N_427,In_70,N_315);
xor U428 (N_428,In_223,N_373);
or U429 (N_429,N_196,In_774);
nor U430 (N_430,In_578,In_651);
and U431 (N_431,In_603,In_67);
and U432 (N_432,In_177,N_213);
and U433 (N_433,N_352,N_127);
xnor U434 (N_434,In_821,N_267);
nor U435 (N_435,In_606,In_74);
and U436 (N_436,N_349,N_273);
xnor U437 (N_437,In_91,In_940);
and U438 (N_438,N_377,In_711);
and U439 (N_439,In_722,N_104);
nor U440 (N_440,In_35,N_328);
and U441 (N_441,N_388,N_380);
and U442 (N_442,In_272,In_482);
nand U443 (N_443,N_359,In_756);
and U444 (N_444,N_345,In_479);
xor U445 (N_445,N_391,N_298);
xnor U446 (N_446,In_154,In_789);
and U447 (N_447,In_885,In_899);
nand U448 (N_448,N_218,In_273);
nor U449 (N_449,In_772,In_814);
or U450 (N_450,In_549,N_117);
and U451 (N_451,In_871,In_507);
nand U452 (N_452,In_723,In_654);
xnor U453 (N_453,N_282,N_188);
and U454 (N_454,N_91,In_561);
and U455 (N_455,In_492,In_591);
and U456 (N_456,N_125,N_212);
and U457 (N_457,N_327,N_329);
or U458 (N_458,In_144,In_202);
xnor U459 (N_459,N_259,N_261);
nand U460 (N_460,In_769,In_313);
xor U461 (N_461,In_399,N_281);
and U462 (N_462,In_644,N_198);
nand U463 (N_463,N_204,N_348);
and U464 (N_464,N_190,In_527);
nand U465 (N_465,In_104,N_386);
nor U466 (N_466,N_285,N_107);
nand U467 (N_467,In_515,N_357);
or U468 (N_468,N_37,In_959);
nand U469 (N_469,N_297,N_135);
nand U470 (N_470,In_164,In_152);
nand U471 (N_471,In_829,In_740);
and U472 (N_472,In_175,N_111);
nand U473 (N_473,In_483,N_353);
or U474 (N_474,N_161,N_82);
nor U475 (N_475,In_23,N_232);
nor U476 (N_476,N_229,In_120);
xor U477 (N_477,In_51,In_587);
or U478 (N_478,In_521,In_325);
or U479 (N_479,In_799,In_667);
xor U480 (N_480,N_189,N_334);
or U481 (N_481,N_61,In_288);
or U482 (N_482,In_134,In_946);
and U483 (N_483,N_38,In_785);
xor U484 (N_484,In_80,In_132);
and U485 (N_485,In_262,In_465);
or U486 (N_486,In_50,N_245);
or U487 (N_487,N_155,N_122);
nor U488 (N_488,In_994,In_366);
xnor U489 (N_489,N_356,N_69);
nor U490 (N_490,In_610,N_389);
nor U491 (N_491,In_130,In_765);
nand U492 (N_492,N_337,In_958);
nand U493 (N_493,In_954,In_810);
nand U494 (N_494,In_771,N_0);
and U495 (N_495,In_455,N_224);
or U496 (N_496,In_926,In_39);
and U497 (N_497,N_361,In_928);
and U498 (N_498,In_461,In_808);
xor U499 (N_499,In_707,N_344);
and U500 (N_500,N_435,In_973);
and U501 (N_501,N_311,In_5);
and U502 (N_502,In_888,N_443);
and U503 (N_503,N_404,N_296);
xnor U504 (N_504,N_399,In_746);
or U505 (N_505,N_376,In_169);
or U506 (N_506,In_903,N_303);
nand U507 (N_507,In_912,N_330);
and U508 (N_508,In_79,N_375);
nor U509 (N_509,In_505,In_216);
nand U510 (N_510,N_335,In_614);
and U511 (N_511,N_472,In_764);
nor U512 (N_512,N_417,In_266);
nor U513 (N_513,In_259,In_553);
xor U514 (N_514,N_230,N_340);
xor U515 (N_515,In_291,N_486);
nor U516 (N_516,N_132,N_215);
and U517 (N_517,N_412,N_466);
and U518 (N_518,N_368,N_475);
xnor U519 (N_519,In_836,In_241);
and U520 (N_520,In_668,N_290);
or U521 (N_521,In_277,N_464);
nor U522 (N_522,N_415,N_431);
nor U523 (N_523,In_106,N_202);
xor U524 (N_524,In_704,N_499);
and U525 (N_525,N_471,In_310);
and U526 (N_526,N_149,N_136);
and U527 (N_527,N_405,N_306);
nand U528 (N_528,N_237,N_478);
and U529 (N_529,N_366,N_305);
and U530 (N_530,N_418,N_459);
nor U531 (N_531,In_125,N_54);
nand U532 (N_532,In_329,N_371);
nand U533 (N_533,In_418,In_467);
or U534 (N_534,N_438,In_1);
nand U535 (N_535,N_363,N_318);
nor U536 (N_536,N_444,N_258);
or U537 (N_537,N_497,N_392);
or U538 (N_538,In_464,In_693);
and U539 (N_539,N_128,N_223);
and U540 (N_540,In_400,N_313);
and U541 (N_541,In_819,In_295);
xor U542 (N_542,In_71,In_999);
and U543 (N_543,N_177,In_78);
or U544 (N_544,N_403,In_710);
and U545 (N_545,N_413,In_116);
nor U546 (N_546,N_246,In_790);
and U547 (N_547,N_320,In_554);
nand U548 (N_548,N_476,N_252);
or U549 (N_549,N_274,In_417);
nand U550 (N_550,In_57,In_770);
nor U551 (N_551,N_419,N_441);
nand U552 (N_552,In_416,N_449);
nand U553 (N_553,N_163,In_643);
and U554 (N_554,N_383,N_333);
nand U555 (N_555,N_80,N_414);
nor U556 (N_556,N_468,N_2);
or U557 (N_557,N_146,N_457);
or U558 (N_558,In_854,N_23);
nand U559 (N_559,In_724,N_180);
or U560 (N_560,N_109,N_455);
or U561 (N_561,In_339,In_830);
nor U562 (N_562,In_394,N_423);
nand U563 (N_563,In_995,In_390);
or U564 (N_564,N_450,In_778);
or U565 (N_565,N_452,In_863);
xor U566 (N_566,N_251,N_433);
xnor U567 (N_567,In_140,In_817);
and U568 (N_568,In_444,In_822);
or U569 (N_569,N_225,N_372);
xor U570 (N_570,In_129,In_847);
nor U571 (N_571,In_398,N_203);
nor U572 (N_572,In_971,In_258);
nand U573 (N_573,N_498,In_77);
or U574 (N_574,N_312,In_137);
or U575 (N_575,In_311,N_78);
or U576 (N_576,N_400,N_390);
or U577 (N_577,In_630,N_491);
or U578 (N_578,N_467,N_367);
nor U579 (N_579,In_540,N_217);
and U580 (N_580,In_859,N_489);
nand U581 (N_581,N_321,In_286);
xnor U582 (N_582,In_602,N_385);
nor U583 (N_583,In_737,In_388);
nor U584 (N_584,N_287,N_184);
nand U585 (N_585,N_407,In_156);
nor U586 (N_586,In_380,N_463);
nand U587 (N_587,N_12,N_323);
nor U588 (N_588,N_95,N_422);
and U589 (N_589,N_293,N_186);
and U590 (N_590,N_126,In_238);
and U591 (N_591,N_437,In_274);
nand U592 (N_592,In_264,In_874);
xnor U593 (N_593,N_490,In_831);
nand U594 (N_594,N_484,In_682);
nand U595 (N_595,In_480,N_33);
nand U596 (N_596,N_434,In_900);
or U597 (N_597,In_203,N_317);
xnor U598 (N_598,N_402,In_232);
xor U599 (N_599,N_351,N_447);
nand U600 (N_600,In_525,N_247);
and U601 (N_601,N_474,N_424);
and U602 (N_602,N_522,N_84);
nor U603 (N_603,In_535,N_51);
or U604 (N_604,In_488,In_332);
nor U605 (N_605,N_394,In_531);
nor U606 (N_606,N_508,N_254);
xor U607 (N_607,N_339,N_291);
nand U608 (N_608,N_523,N_342);
nor U609 (N_609,N_597,In_135);
and U610 (N_610,N_527,N_90);
nand U611 (N_611,N_432,N_411);
and U612 (N_612,N_28,In_253);
nor U613 (N_613,In_689,N_592);
or U614 (N_614,N_219,N_559);
xor U615 (N_615,In_318,N_458);
or U616 (N_616,N_545,In_360);
nand U617 (N_617,In_466,In_86);
or U618 (N_618,N_546,In_968);
nor U619 (N_619,In_248,N_421);
and U620 (N_620,In_786,N_429);
and U621 (N_621,In_211,N_487);
and U622 (N_622,N_568,In_565);
or U623 (N_623,N_262,N_331);
nand U624 (N_624,In_997,N_354);
nand U625 (N_625,N_453,In_949);
nand U626 (N_626,N_573,In_993);
xnor U627 (N_627,N_395,N_338);
nand U628 (N_628,N_170,N_555);
nand U629 (N_629,N_94,N_336);
or U630 (N_630,N_288,N_20);
nor U631 (N_631,In_412,In_931);
nor U632 (N_632,N_483,N_553);
nor U633 (N_633,N_519,N_482);
xor U634 (N_634,N_250,N_426);
nor U635 (N_635,N_567,In_319);
or U636 (N_636,In_364,N_578);
nor U637 (N_637,N_410,N_396);
nor U638 (N_638,N_347,N_358);
nand U639 (N_639,In_82,In_377);
xnor U640 (N_640,N_58,In_502);
nor U641 (N_641,N_153,N_590);
nand U642 (N_642,In_109,In_791);
nor U643 (N_643,In_402,N_233);
nor U644 (N_644,In_700,N_589);
nor U645 (N_645,N_283,In_898);
and U646 (N_646,In_951,N_428);
nand U647 (N_647,N_206,In_862);
or U648 (N_648,N_316,In_122);
and U649 (N_649,N_599,N_577);
xor U650 (N_650,N_382,N_515);
nand U651 (N_651,N_284,In_918);
nand U652 (N_652,N_502,In_306);
nand U653 (N_653,N_461,N_15);
and U654 (N_654,N_79,N_534);
and U655 (N_655,N_231,N_280);
nand U656 (N_656,N_408,N_465);
nand U657 (N_657,N_548,N_241);
nor U658 (N_658,In_356,N_234);
xor U659 (N_659,N_319,N_440);
nand U660 (N_660,In_284,In_501);
and U661 (N_661,N_500,N_393);
xnor U662 (N_662,N_120,N_495);
nand U663 (N_663,N_542,N_528);
and U664 (N_664,N_208,In_532);
nor U665 (N_665,N_178,In_520);
nor U666 (N_666,N_593,N_462);
nand U667 (N_667,In_147,N_265);
or U668 (N_668,N_541,N_591);
xor U669 (N_669,N_514,N_596);
xnor U670 (N_670,N_384,In_989);
or U671 (N_671,N_513,In_414);
nand U672 (N_672,In_559,N_374);
nor U673 (N_673,In_265,N_309);
nand U674 (N_674,In_128,N_503);
or U675 (N_675,N_448,N_277);
xor U676 (N_676,In_745,In_672);
and U677 (N_677,N_575,N_533);
nand U678 (N_678,N_526,In_447);
nand U679 (N_679,N_378,N_531);
xnor U680 (N_680,In_330,In_571);
or U681 (N_681,N_166,In_818);
nand U682 (N_682,N_439,N_379);
xnor U683 (N_683,N_511,In_376);
nor U684 (N_684,N_563,N_49);
and U685 (N_685,N_579,In_731);
or U686 (N_686,In_592,In_766);
and U687 (N_687,In_420,N_406);
nor U688 (N_688,N_552,In_97);
and U689 (N_689,N_505,N_158);
or U690 (N_690,N_16,N_350);
xor U691 (N_691,N_539,N_525);
or U692 (N_692,In_944,N_473);
nand U693 (N_693,N_64,N_271);
xnor U694 (N_694,N_301,N_496);
xor U695 (N_695,In_363,N_547);
and U696 (N_696,N_520,N_582);
or U697 (N_697,In_742,In_895);
or U698 (N_698,N_560,In_683);
and U699 (N_699,In_370,N_595);
xnor U700 (N_700,In_72,N_630);
and U701 (N_701,In_369,N_693);
and U702 (N_702,N_92,N_445);
nor U703 (N_703,In_68,N_100);
nor U704 (N_704,N_544,In_181);
nand U705 (N_705,In_622,N_27);
xor U706 (N_706,N_310,N_454);
and U707 (N_707,N_643,In_777);
nand U708 (N_708,N_627,N_676);
xnor U709 (N_709,In_865,N_387);
xor U710 (N_710,N_585,N_427);
nand U711 (N_711,N_536,N_401);
nand U712 (N_712,N_48,N_698);
nor U713 (N_713,In_661,N_646);
and U714 (N_714,N_604,N_614);
xnor U715 (N_715,N_238,N_26);
and U716 (N_716,N_587,N_270);
or U717 (N_717,N_537,N_583);
and U718 (N_718,N_689,N_479);
and U719 (N_719,In_413,N_509);
xnor U720 (N_720,N_138,In_500);
nor U721 (N_721,N_307,In_698);
nor U722 (N_722,N_397,N_645);
nand U723 (N_723,N_686,N_670);
xor U724 (N_724,N_601,N_620);
nand U725 (N_725,N_697,In_285);
nand U726 (N_726,N_602,N_623);
nor U727 (N_727,In_911,N_625);
or U728 (N_728,N_248,In_0);
or U729 (N_729,N_678,N_510);
xnor U730 (N_730,N_616,N_691);
nor U731 (N_731,N_529,N_663);
xnor U732 (N_732,N_362,N_488);
nand U733 (N_733,N_649,N_518);
and U734 (N_734,N_194,N_641);
and U735 (N_735,N_576,In_347);
nor U736 (N_736,In_354,In_19);
xor U737 (N_737,N_690,N_549);
nor U738 (N_738,N_586,In_17);
nand U739 (N_739,N_675,N_214);
or U740 (N_740,N_642,N_558);
xnor U741 (N_741,N_647,N_654);
xnor U742 (N_742,N_343,In_935);
nand U743 (N_743,N_618,N_688);
nor U744 (N_744,N_346,N_469);
nand U745 (N_745,N_598,N_494);
and U746 (N_746,N_600,In_351);
and U747 (N_747,N_129,N_650);
and U748 (N_748,N_299,In_346);
and U749 (N_749,N_610,N_569);
nor U750 (N_750,N_209,N_695);
nor U751 (N_751,N_571,N_653);
xor U752 (N_752,In_150,N_566);
nand U753 (N_753,N_667,N_562);
and U754 (N_754,In_9,In_452);
xnor U755 (N_755,N_621,In_391);
nor U756 (N_756,N_370,N_118);
and U757 (N_757,N_369,N_492);
or U758 (N_758,N_581,N_538);
nor U759 (N_759,N_672,N_637);
nor U760 (N_760,N_485,In_657);
and U761 (N_761,N_292,N_683);
nand U762 (N_762,N_460,In_747);
xnor U763 (N_763,N_150,N_660);
nor U764 (N_764,N_409,N_681);
or U765 (N_765,In_545,N_99);
xnor U766 (N_766,N_477,N_302);
nand U767 (N_767,N_521,N_657);
nand U768 (N_768,N_172,N_550);
or U769 (N_769,N_674,In_55);
nand U770 (N_770,N_556,N_570);
nand U771 (N_771,N_535,N_554);
and U772 (N_772,N_613,N_662);
xnor U773 (N_773,N_286,N_304);
nand U774 (N_774,N_605,N_632);
nand U775 (N_775,N_501,N_607);
or U776 (N_776,N_564,In_28);
nand U777 (N_777,N_651,In_568);
or U778 (N_778,N_360,N_425);
nand U779 (N_779,N_622,N_516);
nand U780 (N_780,In_2,N_631);
nand U781 (N_781,N_687,N_635);
nor U782 (N_782,N_524,N_612);
or U783 (N_783,N_692,In_442);
nor U784 (N_784,N_148,N_696);
nor U785 (N_785,N_451,N_142);
nor U786 (N_786,N_638,In_879);
nor U787 (N_787,N_603,N_442);
and U788 (N_788,N_420,N_504);
nand U789 (N_789,In_749,N_324);
xnor U790 (N_790,In_673,In_221);
or U791 (N_791,N_493,N_543);
and U792 (N_792,N_512,N_636);
xnor U793 (N_793,N_530,In_589);
xnor U794 (N_794,N_574,N_671);
or U795 (N_795,N_588,N_626);
xnor U796 (N_796,In_165,N_430);
nand U797 (N_797,N_235,N_648);
nor U798 (N_798,N_19,N_446);
xor U799 (N_799,N_640,In_15);
nand U800 (N_800,N_791,In_961);
or U801 (N_801,N_685,N_611);
nand U802 (N_802,N_702,N_322);
or U803 (N_803,N_768,N_725);
nand U804 (N_804,N_185,N_713);
and U805 (N_805,N_726,N_666);
and U806 (N_806,N_264,N_754);
or U807 (N_807,N_758,N_769);
and U808 (N_808,N_712,N_710);
and U809 (N_809,N_761,N_795);
nand U810 (N_810,N_699,N_656);
nand U811 (N_811,In_166,N_744);
and U812 (N_812,N_668,N_750);
or U813 (N_813,N_790,N_741);
nand U814 (N_814,N_594,N_480);
and U815 (N_815,N_734,In_851);
or U816 (N_816,N_609,N_694);
nor U817 (N_817,N_416,N_714);
or U818 (N_818,N_737,N_308);
and U819 (N_819,In_732,N_708);
or U820 (N_820,In_941,N_711);
nand U821 (N_821,N_727,N_794);
and U822 (N_822,N_742,N_242);
xnor U823 (N_823,N_762,N_456);
xor U824 (N_824,N_775,N_718);
or U825 (N_825,N_728,In_609);
and U826 (N_826,N_96,N_517);
or U827 (N_827,N_633,N_47);
xor U828 (N_828,N_326,N_717);
and U829 (N_829,N_191,N_168);
xnor U830 (N_830,N_782,N_716);
xor U831 (N_831,N_617,N_557);
xnor U832 (N_832,N_719,N_759);
and U833 (N_833,N_743,N_701);
and U834 (N_834,In_237,N_341);
nand U835 (N_835,N_760,N_755);
or U836 (N_836,In_484,N_731);
nand U837 (N_837,N_724,N_704);
xnor U838 (N_838,N_507,N_540);
xor U839 (N_839,N_160,N_732);
and U840 (N_840,In_986,N_753);
xor U841 (N_841,N_715,N_770);
nor U842 (N_842,N_628,N_780);
nand U843 (N_843,In_194,N_332);
xnor U844 (N_844,N_706,N_655);
and U845 (N_845,N_776,N_729);
and U846 (N_846,N_669,N_740);
and U847 (N_847,N_700,N_766);
nor U848 (N_848,N_767,N_730);
nand U849 (N_849,N_619,In_289);
and U850 (N_850,N_680,N_748);
and U851 (N_851,N_746,N_745);
xor U852 (N_852,N_796,N_756);
or U853 (N_853,N_470,In_803);
or U854 (N_854,In_751,N_707);
nand U855 (N_855,N_634,N_783);
or U856 (N_856,N_749,N_436);
or U857 (N_857,N_639,N_720);
nor U858 (N_858,N_738,N_355);
nor U859 (N_859,N_777,N_793);
nor U860 (N_860,N_786,N_580);
nand U861 (N_861,N_253,N_269);
nand U862 (N_862,N_236,N_227);
or U863 (N_863,N_481,N_736);
nand U864 (N_864,N_679,N_551);
or U865 (N_865,N_792,N_721);
xor U866 (N_866,N_584,In_923);
and U867 (N_867,N_747,N_684);
nand U868 (N_868,N_243,N_779);
or U869 (N_869,In_43,N_774);
or U870 (N_870,N_798,N_398);
nand U871 (N_871,N_739,N_787);
or U872 (N_872,N_797,N_752);
nand U873 (N_873,N_644,N_572);
xor U874 (N_874,N_615,N_789);
or U875 (N_875,N_772,N_771);
or U876 (N_876,N_788,N_733);
nand U877 (N_877,N_703,In_114);
and U878 (N_878,N_314,In_934);
or U879 (N_879,N_764,N_624);
nand U880 (N_880,N_751,N_781);
xnor U881 (N_881,In_182,N_606);
nor U882 (N_882,In_490,N_677);
and U883 (N_883,N_765,In_342);
xnor U884 (N_884,N_659,N_784);
nor U885 (N_885,In_838,N_532);
and U886 (N_886,N_565,N_629);
or U887 (N_887,N_664,N_608);
nor U888 (N_888,N_778,N_773);
or U889 (N_889,N_723,N_722);
xnor U890 (N_890,In_735,N_673);
nor U891 (N_891,N_658,N_665);
xor U892 (N_892,N_57,N_763);
and U893 (N_893,N_561,N_735);
and U894 (N_894,In_410,N_506);
and U895 (N_895,N_757,In_304);
and U896 (N_896,N_652,In_340);
and U897 (N_897,N_661,N_709);
and U898 (N_898,N_799,N_705);
and U899 (N_899,N_682,N_785);
or U900 (N_900,N_854,N_820);
nor U901 (N_901,N_878,N_840);
and U902 (N_902,N_812,N_813);
or U903 (N_903,N_830,N_845);
or U904 (N_904,N_804,N_805);
nor U905 (N_905,N_874,N_891);
xor U906 (N_906,N_859,N_806);
or U907 (N_907,N_871,N_846);
and U908 (N_908,N_897,N_896);
and U909 (N_909,N_832,N_867);
or U910 (N_910,N_866,N_856);
nor U911 (N_911,N_811,N_828);
xor U912 (N_912,N_802,N_863);
or U913 (N_913,N_821,N_849);
and U914 (N_914,N_844,N_868);
xor U915 (N_915,N_899,N_869);
nor U916 (N_916,N_831,N_881);
or U917 (N_917,N_895,N_865);
xor U918 (N_918,N_824,N_885);
nand U919 (N_919,N_816,N_818);
or U920 (N_920,N_884,N_823);
and U921 (N_921,N_839,N_807);
or U922 (N_922,N_882,N_888);
and U923 (N_923,N_826,N_853);
nand U924 (N_924,N_857,N_875);
xnor U925 (N_925,N_836,N_860);
nor U926 (N_926,N_843,N_808);
xnor U927 (N_927,N_879,N_847);
and U928 (N_928,N_814,N_877);
xor U929 (N_929,N_858,N_803);
xnor U930 (N_930,N_815,N_817);
nor U931 (N_931,N_835,N_862);
xnor U932 (N_932,N_870,N_864);
nand U933 (N_933,N_873,N_819);
nand U934 (N_934,N_838,N_898);
nor U935 (N_935,N_887,N_872);
nor U936 (N_936,N_841,N_893);
or U937 (N_937,N_842,N_880);
or U938 (N_938,N_834,N_886);
or U939 (N_939,N_848,N_892);
nor U940 (N_940,N_890,N_825);
and U941 (N_941,N_852,N_883);
or U942 (N_942,N_827,N_800);
xnor U943 (N_943,N_837,N_894);
and U944 (N_944,N_876,N_810);
nand U945 (N_945,N_822,N_851);
nand U946 (N_946,N_801,N_850);
nor U947 (N_947,N_861,N_829);
or U948 (N_948,N_889,N_809);
or U949 (N_949,N_855,N_833);
xor U950 (N_950,N_863,N_865);
nor U951 (N_951,N_885,N_806);
and U952 (N_952,N_889,N_849);
nand U953 (N_953,N_823,N_841);
nor U954 (N_954,N_828,N_841);
or U955 (N_955,N_863,N_893);
xor U956 (N_956,N_851,N_895);
and U957 (N_957,N_851,N_868);
and U958 (N_958,N_886,N_861);
and U959 (N_959,N_881,N_829);
nor U960 (N_960,N_855,N_818);
xor U961 (N_961,N_829,N_810);
nor U962 (N_962,N_827,N_820);
nor U963 (N_963,N_846,N_822);
nand U964 (N_964,N_859,N_844);
or U965 (N_965,N_881,N_859);
nand U966 (N_966,N_838,N_889);
or U967 (N_967,N_810,N_881);
xor U968 (N_968,N_852,N_870);
nor U969 (N_969,N_822,N_857);
nand U970 (N_970,N_865,N_812);
nor U971 (N_971,N_876,N_807);
nor U972 (N_972,N_801,N_809);
nand U973 (N_973,N_866,N_837);
nand U974 (N_974,N_857,N_813);
nand U975 (N_975,N_881,N_893);
and U976 (N_976,N_816,N_895);
and U977 (N_977,N_831,N_871);
nand U978 (N_978,N_842,N_817);
nor U979 (N_979,N_893,N_823);
nor U980 (N_980,N_863,N_800);
and U981 (N_981,N_853,N_851);
or U982 (N_982,N_857,N_847);
nand U983 (N_983,N_888,N_886);
or U984 (N_984,N_818,N_896);
xnor U985 (N_985,N_844,N_866);
nand U986 (N_986,N_873,N_829);
xor U987 (N_987,N_842,N_804);
nand U988 (N_988,N_835,N_887);
and U989 (N_989,N_829,N_821);
nor U990 (N_990,N_845,N_859);
and U991 (N_991,N_847,N_889);
nor U992 (N_992,N_824,N_872);
nand U993 (N_993,N_857,N_843);
nand U994 (N_994,N_844,N_820);
nor U995 (N_995,N_836,N_899);
or U996 (N_996,N_887,N_812);
nand U997 (N_997,N_892,N_891);
nor U998 (N_998,N_859,N_821);
nor U999 (N_999,N_889,N_859);
or U1000 (N_1000,N_949,N_966);
xor U1001 (N_1001,N_974,N_969);
nor U1002 (N_1002,N_963,N_942);
xnor U1003 (N_1003,N_975,N_953);
nand U1004 (N_1004,N_970,N_955);
and U1005 (N_1005,N_951,N_952);
or U1006 (N_1006,N_914,N_948);
xor U1007 (N_1007,N_918,N_985);
or U1008 (N_1008,N_973,N_932);
or U1009 (N_1009,N_938,N_971);
nor U1010 (N_1010,N_965,N_943);
xor U1011 (N_1011,N_989,N_957);
nor U1012 (N_1012,N_978,N_956);
nand U1013 (N_1013,N_913,N_906);
or U1014 (N_1014,N_907,N_977);
xnor U1015 (N_1015,N_944,N_936);
nor U1016 (N_1016,N_926,N_916);
nor U1017 (N_1017,N_911,N_968);
xnor U1018 (N_1018,N_986,N_902);
and U1019 (N_1019,N_903,N_922);
or U1020 (N_1020,N_909,N_950);
and U1021 (N_1021,N_992,N_980);
nand U1022 (N_1022,N_987,N_947);
nand U1023 (N_1023,N_934,N_972);
nand U1024 (N_1024,N_905,N_967);
and U1025 (N_1025,N_983,N_998);
nor U1026 (N_1026,N_994,N_964);
xnor U1027 (N_1027,N_935,N_927);
and U1028 (N_1028,N_958,N_997);
and U1029 (N_1029,N_990,N_924);
or U1030 (N_1030,N_900,N_945);
or U1031 (N_1031,N_954,N_961);
nand U1032 (N_1032,N_920,N_941);
or U1033 (N_1033,N_931,N_940);
xor U1034 (N_1034,N_928,N_996);
or U1035 (N_1035,N_937,N_939);
nor U1036 (N_1036,N_999,N_923);
nor U1037 (N_1037,N_912,N_930);
and U1038 (N_1038,N_960,N_984);
nor U1039 (N_1039,N_929,N_979);
nand U1040 (N_1040,N_933,N_981);
and U1041 (N_1041,N_901,N_919);
nand U1042 (N_1042,N_988,N_921);
and U1043 (N_1043,N_946,N_976);
and U1044 (N_1044,N_908,N_915);
or U1045 (N_1045,N_991,N_993);
xnor U1046 (N_1046,N_910,N_904);
nand U1047 (N_1047,N_925,N_917);
xnor U1048 (N_1048,N_962,N_982);
xor U1049 (N_1049,N_959,N_995);
nand U1050 (N_1050,N_907,N_965);
and U1051 (N_1051,N_939,N_920);
and U1052 (N_1052,N_929,N_981);
xnor U1053 (N_1053,N_970,N_912);
nor U1054 (N_1054,N_912,N_967);
xnor U1055 (N_1055,N_924,N_976);
or U1056 (N_1056,N_987,N_926);
or U1057 (N_1057,N_931,N_962);
xnor U1058 (N_1058,N_973,N_954);
and U1059 (N_1059,N_976,N_963);
xor U1060 (N_1060,N_901,N_952);
and U1061 (N_1061,N_914,N_928);
xnor U1062 (N_1062,N_962,N_973);
and U1063 (N_1063,N_924,N_975);
nor U1064 (N_1064,N_955,N_940);
nor U1065 (N_1065,N_948,N_989);
xor U1066 (N_1066,N_938,N_949);
or U1067 (N_1067,N_903,N_953);
nor U1068 (N_1068,N_917,N_968);
xor U1069 (N_1069,N_946,N_902);
xnor U1070 (N_1070,N_982,N_935);
nand U1071 (N_1071,N_921,N_920);
nand U1072 (N_1072,N_977,N_964);
nand U1073 (N_1073,N_953,N_919);
xnor U1074 (N_1074,N_954,N_916);
xor U1075 (N_1075,N_933,N_935);
xor U1076 (N_1076,N_993,N_983);
or U1077 (N_1077,N_939,N_908);
xnor U1078 (N_1078,N_933,N_912);
and U1079 (N_1079,N_996,N_908);
or U1080 (N_1080,N_958,N_991);
and U1081 (N_1081,N_975,N_907);
xnor U1082 (N_1082,N_944,N_966);
nand U1083 (N_1083,N_933,N_997);
nor U1084 (N_1084,N_994,N_935);
and U1085 (N_1085,N_981,N_965);
or U1086 (N_1086,N_950,N_904);
or U1087 (N_1087,N_964,N_975);
nor U1088 (N_1088,N_990,N_946);
or U1089 (N_1089,N_998,N_942);
xnor U1090 (N_1090,N_956,N_927);
or U1091 (N_1091,N_941,N_911);
nor U1092 (N_1092,N_945,N_966);
or U1093 (N_1093,N_999,N_944);
and U1094 (N_1094,N_907,N_947);
nor U1095 (N_1095,N_902,N_981);
or U1096 (N_1096,N_998,N_961);
or U1097 (N_1097,N_939,N_936);
and U1098 (N_1098,N_913,N_989);
nor U1099 (N_1099,N_954,N_949);
and U1100 (N_1100,N_1063,N_1082);
nor U1101 (N_1101,N_1009,N_1058);
xor U1102 (N_1102,N_1011,N_1042);
nand U1103 (N_1103,N_1007,N_1028);
nor U1104 (N_1104,N_1090,N_1039);
xnor U1105 (N_1105,N_1065,N_1015);
nand U1106 (N_1106,N_1081,N_1077);
or U1107 (N_1107,N_1013,N_1076);
and U1108 (N_1108,N_1008,N_1073);
nor U1109 (N_1109,N_1075,N_1032);
xor U1110 (N_1110,N_1070,N_1014);
nor U1111 (N_1111,N_1020,N_1016);
or U1112 (N_1112,N_1079,N_1094);
and U1113 (N_1113,N_1099,N_1084);
or U1114 (N_1114,N_1071,N_1038);
and U1115 (N_1115,N_1069,N_1006);
nand U1116 (N_1116,N_1098,N_1056);
nor U1117 (N_1117,N_1067,N_1033);
xor U1118 (N_1118,N_1095,N_1001);
nor U1119 (N_1119,N_1017,N_1022);
and U1120 (N_1120,N_1024,N_1036);
and U1121 (N_1121,N_1053,N_1018);
xnor U1122 (N_1122,N_1005,N_1034);
nand U1123 (N_1123,N_1064,N_1061);
xnor U1124 (N_1124,N_1045,N_1055);
and U1125 (N_1125,N_1060,N_1047);
nor U1126 (N_1126,N_1029,N_1031);
and U1127 (N_1127,N_1010,N_1066);
or U1128 (N_1128,N_1041,N_1050);
nand U1129 (N_1129,N_1023,N_1087);
or U1130 (N_1130,N_1059,N_1030);
xnor U1131 (N_1131,N_1091,N_1027);
xor U1132 (N_1132,N_1093,N_1052);
nor U1133 (N_1133,N_1046,N_1083);
nor U1134 (N_1134,N_1062,N_1044);
and U1135 (N_1135,N_1088,N_1012);
and U1136 (N_1136,N_1043,N_1040);
or U1137 (N_1137,N_1025,N_1080);
nor U1138 (N_1138,N_1097,N_1057);
nand U1139 (N_1139,N_1000,N_1026);
nand U1140 (N_1140,N_1004,N_1003);
xnor U1141 (N_1141,N_1072,N_1037);
nor U1142 (N_1142,N_1021,N_1085);
or U1143 (N_1143,N_1092,N_1074);
and U1144 (N_1144,N_1086,N_1078);
xnor U1145 (N_1145,N_1002,N_1068);
nand U1146 (N_1146,N_1035,N_1049);
or U1147 (N_1147,N_1019,N_1089);
or U1148 (N_1148,N_1054,N_1051);
and U1149 (N_1149,N_1096,N_1048);
nand U1150 (N_1150,N_1008,N_1074);
or U1151 (N_1151,N_1056,N_1002);
nor U1152 (N_1152,N_1003,N_1094);
and U1153 (N_1153,N_1023,N_1000);
xnor U1154 (N_1154,N_1015,N_1092);
nor U1155 (N_1155,N_1040,N_1029);
nor U1156 (N_1156,N_1040,N_1061);
or U1157 (N_1157,N_1031,N_1014);
or U1158 (N_1158,N_1046,N_1019);
nor U1159 (N_1159,N_1043,N_1005);
nor U1160 (N_1160,N_1085,N_1090);
nor U1161 (N_1161,N_1003,N_1016);
nor U1162 (N_1162,N_1048,N_1037);
and U1163 (N_1163,N_1052,N_1090);
nand U1164 (N_1164,N_1041,N_1073);
nor U1165 (N_1165,N_1031,N_1022);
nand U1166 (N_1166,N_1040,N_1024);
nand U1167 (N_1167,N_1027,N_1020);
or U1168 (N_1168,N_1004,N_1006);
nand U1169 (N_1169,N_1098,N_1000);
and U1170 (N_1170,N_1010,N_1072);
or U1171 (N_1171,N_1023,N_1075);
xor U1172 (N_1172,N_1070,N_1020);
or U1173 (N_1173,N_1034,N_1004);
and U1174 (N_1174,N_1040,N_1048);
or U1175 (N_1175,N_1065,N_1086);
nor U1176 (N_1176,N_1036,N_1084);
nor U1177 (N_1177,N_1045,N_1033);
xor U1178 (N_1178,N_1025,N_1073);
nand U1179 (N_1179,N_1099,N_1024);
or U1180 (N_1180,N_1039,N_1023);
or U1181 (N_1181,N_1011,N_1017);
and U1182 (N_1182,N_1073,N_1062);
nor U1183 (N_1183,N_1091,N_1055);
nand U1184 (N_1184,N_1098,N_1011);
or U1185 (N_1185,N_1000,N_1087);
or U1186 (N_1186,N_1023,N_1082);
or U1187 (N_1187,N_1066,N_1020);
nand U1188 (N_1188,N_1006,N_1011);
xor U1189 (N_1189,N_1002,N_1088);
nand U1190 (N_1190,N_1018,N_1061);
xnor U1191 (N_1191,N_1036,N_1074);
and U1192 (N_1192,N_1006,N_1005);
xnor U1193 (N_1193,N_1097,N_1065);
and U1194 (N_1194,N_1090,N_1032);
nor U1195 (N_1195,N_1064,N_1066);
nand U1196 (N_1196,N_1081,N_1088);
xnor U1197 (N_1197,N_1068,N_1010);
or U1198 (N_1198,N_1079,N_1049);
xor U1199 (N_1199,N_1005,N_1070);
or U1200 (N_1200,N_1151,N_1105);
and U1201 (N_1201,N_1175,N_1102);
xor U1202 (N_1202,N_1195,N_1180);
and U1203 (N_1203,N_1179,N_1174);
xnor U1204 (N_1204,N_1103,N_1198);
and U1205 (N_1205,N_1156,N_1150);
nor U1206 (N_1206,N_1121,N_1185);
and U1207 (N_1207,N_1160,N_1118);
or U1208 (N_1208,N_1158,N_1119);
nor U1209 (N_1209,N_1173,N_1193);
nand U1210 (N_1210,N_1189,N_1168);
or U1211 (N_1211,N_1167,N_1131);
nor U1212 (N_1212,N_1120,N_1129);
xnor U1213 (N_1213,N_1196,N_1114);
nor U1214 (N_1214,N_1184,N_1100);
nand U1215 (N_1215,N_1177,N_1135);
or U1216 (N_1216,N_1110,N_1142);
xor U1217 (N_1217,N_1133,N_1190);
nor U1218 (N_1218,N_1126,N_1123);
nand U1219 (N_1219,N_1199,N_1182);
nor U1220 (N_1220,N_1161,N_1132);
and U1221 (N_1221,N_1115,N_1163);
nor U1222 (N_1222,N_1176,N_1152);
xor U1223 (N_1223,N_1124,N_1157);
or U1224 (N_1224,N_1186,N_1197);
and U1225 (N_1225,N_1154,N_1138);
or U1226 (N_1226,N_1146,N_1181);
or U1227 (N_1227,N_1183,N_1144);
and U1228 (N_1228,N_1145,N_1139);
nor U1229 (N_1229,N_1178,N_1187);
nand U1230 (N_1230,N_1130,N_1153);
nor U1231 (N_1231,N_1113,N_1171);
or U1232 (N_1232,N_1127,N_1111);
and U1233 (N_1233,N_1134,N_1169);
nor U1234 (N_1234,N_1147,N_1143);
nand U1235 (N_1235,N_1101,N_1116);
nor U1236 (N_1236,N_1164,N_1107);
or U1237 (N_1237,N_1159,N_1106);
nand U1238 (N_1238,N_1109,N_1170);
nor U1239 (N_1239,N_1122,N_1149);
nand U1240 (N_1240,N_1172,N_1194);
xnor U1241 (N_1241,N_1155,N_1117);
nand U1242 (N_1242,N_1125,N_1137);
and U1243 (N_1243,N_1165,N_1191);
and U1244 (N_1244,N_1162,N_1104);
and U1245 (N_1245,N_1108,N_1188);
or U1246 (N_1246,N_1112,N_1128);
or U1247 (N_1247,N_1136,N_1148);
xnor U1248 (N_1248,N_1141,N_1192);
xor U1249 (N_1249,N_1140,N_1166);
nand U1250 (N_1250,N_1194,N_1195);
nand U1251 (N_1251,N_1116,N_1182);
xor U1252 (N_1252,N_1175,N_1165);
nor U1253 (N_1253,N_1185,N_1112);
xnor U1254 (N_1254,N_1119,N_1195);
and U1255 (N_1255,N_1110,N_1155);
or U1256 (N_1256,N_1164,N_1158);
nor U1257 (N_1257,N_1150,N_1147);
xnor U1258 (N_1258,N_1117,N_1165);
nand U1259 (N_1259,N_1141,N_1166);
nand U1260 (N_1260,N_1182,N_1189);
or U1261 (N_1261,N_1137,N_1110);
nand U1262 (N_1262,N_1104,N_1135);
nand U1263 (N_1263,N_1141,N_1170);
or U1264 (N_1264,N_1166,N_1119);
xor U1265 (N_1265,N_1161,N_1100);
xnor U1266 (N_1266,N_1166,N_1146);
xor U1267 (N_1267,N_1159,N_1128);
nor U1268 (N_1268,N_1191,N_1130);
nand U1269 (N_1269,N_1194,N_1170);
or U1270 (N_1270,N_1136,N_1154);
nor U1271 (N_1271,N_1170,N_1112);
nand U1272 (N_1272,N_1104,N_1132);
or U1273 (N_1273,N_1143,N_1171);
and U1274 (N_1274,N_1188,N_1137);
and U1275 (N_1275,N_1136,N_1116);
xnor U1276 (N_1276,N_1130,N_1129);
xnor U1277 (N_1277,N_1140,N_1108);
xnor U1278 (N_1278,N_1174,N_1113);
nand U1279 (N_1279,N_1130,N_1104);
or U1280 (N_1280,N_1133,N_1184);
xor U1281 (N_1281,N_1168,N_1140);
or U1282 (N_1282,N_1162,N_1164);
and U1283 (N_1283,N_1189,N_1161);
nand U1284 (N_1284,N_1193,N_1160);
nor U1285 (N_1285,N_1117,N_1186);
and U1286 (N_1286,N_1153,N_1154);
xor U1287 (N_1287,N_1190,N_1186);
or U1288 (N_1288,N_1158,N_1145);
nor U1289 (N_1289,N_1182,N_1142);
xnor U1290 (N_1290,N_1197,N_1175);
and U1291 (N_1291,N_1190,N_1165);
xnor U1292 (N_1292,N_1159,N_1117);
nor U1293 (N_1293,N_1163,N_1150);
or U1294 (N_1294,N_1190,N_1184);
nand U1295 (N_1295,N_1122,N_1199);
nand U1296 (N_1296,N_1149,N_1143);
and U1297 (N_1297,N_1140,N_1119);
xnor U1298 (N_1298,N_1181,N_1145);
xor U1299 (N_1299,N_1186,N_1174);
and U1300 (N_1300,N_1232,N_1217);
nand U1301 (N_1301,N_1207,N_1229);
and U1302 (N_1302,N_1247,N_1299);
and U1303 (N_1303,N_1271,N_1270);
nor U1304 (N_1304,N_1228,N_1288);
or U1305 (N_1305,N_1235,N_1298);
xnor U1306 (N_1306,N_1280,N_1258);
nor U1307 (N_1307,N_1216,N_1253);
nand U1308 (N_1308,N_1219,N_1226);
nand U1309 (N_1309,N_1295,N_1213);
nand U1310 (N_1310,N_1202,N_1263);
or U1311 (N_1311,N_1294,N_1265);
nor U1312 (N_1312,N_1261,N_1291);
xnor U1313 (N_1313,N_1203,N_1234);
nor U1314 (N_1314,N_1284,N_1208);
or U1315 (N_1315,N_1274,N_1257);
xor U1316 (N_1316,N_1220,N_1225);
nor U1317 (N_1317,N_1243,N_1239);
or U1318 (N_1318,N_1221,N_1268);
nand U1319 (N_1319,N_1215,N_1244);
nand U1320 (N_1320,N_1285,N_1206);
nand U1321 (N_1321,N_1259,N_1240);
xnor U1322 (N_1322,N_1223,N_1266);
and U1323 (N_1323,N_1248,N_1238);
or U1324 (N_1324,N_1245,N_1278);
nand U1325 (N_1325,N_1282,N_1267);
or U1326 (N_1326,N_1200,N_1205);
nand U1327 (N_1327,N_1256,N_1283);
nand U1328 (N_1328,N_1293,N_1255);
nor U1329 (N_1329,N_1264,N_1212);
xor U1330 (N_1330,N_1276,N_1296);
or U1331 (N_1331,N_1252,N_1237);
nand U1332 (N_1332,N_1260,N_1273);
or U1333 (N_1333,N_1236,N_1210);
and U1334 (N_1334,N_1241,N_1281);
or U1335 (N_1335,N_1262,N_1249);
and U1336 (N_1336,N_1275,N_1279);
nand U1337 (N_1337,N_1250,N_1292);
nand U1338 (N_1338,N_1224,N_1242);
nor U1339 (N_1339,N_1227,N_1222);
nand U1340 (N_1340,N_1214,N_1251);
or U1341 (N_1341,N_1289,N_1218);
nand U1342 (N_1342,N_1297,N_1287);
nand U1343 (N_1343,N_1272,N_1277);
nor U1344 (N_1344,N_1211,N_1231);
and U1345 (N_1345,N_1254,N_1209);
or U1346 (N_1346,N_1204,N_1286);
and U1347 (N_1347,N_1233,N_1290);
or U1348 (N_1348,N_1246,N_1269);
and U1349 (N_1349,N_1201,N_1230);
or U1350 (N_1350,N_1293,N_1270);
and U1351 (N_1351,N_1203,N_1278);
nor U1352 (N_1352,N_1249,N_1266);
and U1353 (N_1353,N_1266,N_1230);
xor U1354 (N_1354,N_1212,N_1286);
nor U1355 (N_1355,N_1248,N_1297);
xnor U1356 (N_1356,N_1261,N_1267);
or U1357 (N_1357,N_1295,N_1202);
nor U1358 (N_1358,N_1268,N_1206);
xnor U1359 (N_1359,N_1273,N_1278);
xor U1360 (N_1360,N_1251,N_1280);
xor U1361 (N_1361,N_1287,N_1279);
xnor U1362 (N_1362,N_1252,N_1205);
nand U1363 (N_1363,N_1214,N_1240);
or U1364 (N_1364,N_1286,N_1240);
or U1365 (N_1365,N_1222,N_1213);
or U1366 (N_1366,N_1292,N_1291);
or U1367 (N_1367,N_1276,N_1268);
or U1368 (N_1368,N_1275,N_1214);
nand U1369 (N_1369,N_1221,N_1258);
and U1370 (N_1370,N_1284,N_1281);
nand U1371 (N_1371,N_1266,N_1235);
and U1372 (N_1372,N_1284,N_1288);
and U1373 (N_1373,N_1244,N_1224);
nor U1374 (N_1374,N_1286,N_1282);
nor U1375 (N_1375,N_1213,N_1296);
and U1376 (N_1376,N_1266,N_1274);
nand U1377 (N_1377,N_1233,N_1211);
nand U1378 (N_1378,N_1275,N_1233);
and U1379 (N_1379,N_1239,N_1201);
or U1380 (N_1380,N_1200,N_1299);
and U1381 (N_1381,N_1262,N_1274);
and U1382 (N_1382,N_1261,N_1205);
nand U1383 (N_1383,N_1250,N_1258);
or U1384 (N_1384,N_1297,N_1262);
xor U1385 (N_1385,N_1226,N_1274);
nor U1386 (N_1386,N_1242,N_1231);
xor U1387 (N_1387,N_1203,N_1270);
nor U1388 (N_1388,N_1292,N_1258);
nand U1389 (N_1389,N_1298,N_1208);
and U1390 (N_1390,N_1282,N_1299);
xnor U1391 (N_1391,N_1235,N_1249);
xor U1392 (N_1392,N_1212,N_1276);
nand U1393 (N_1393,N_1273,N_1235);
nor U1394 (N_1394,N_1214,N_1299);
and U1395 (N_1395,N_1209,N_1265);
and U1396 (N_1396,N_1240,N_1278);
nand U1397 (N_1397,N_1241,N_1219);
nand U1398 (N_1398,N_1249,N_1208);
xnor U1399 (N_1399,N_1253,N_1249);
nor U1400 (N_1400,N_1300,N_1316);
or U1401 (N_1401,N_1361,N_1383);
nor U1402 (N_1402,N_1343,N_1393);
nor U1403 (N_1403,N_1375,N_1370);
xor U1404 (N_1404,N_1349,N_1387);
xnor U1405 (N_1405,N_1319,N_1363);
nor U1406 (N_1406,N_1371,N_1323);
or U1407 (N_1407,N_1338,N_1358);
or U1408 (N_1408,N_1345,N_1302);
nor U1409 (N_1409,N_1388,N_1333);
nand U1410 (N_1410,N_1369,N_1307);
and U1411 (N_1411,N_1386,N_1324);
nand U1412 (N_1412,N_1309,N_1365);
nor U1413 (N_1413,N_1303,N_1355);
or U1414 (N_1414,N_1331,N_1325);
or U1415 (N_1415,N_1342,N_1382);
or U1416 (N_1416,N_1310,N_1335);
and U1417 (N_1417,N_1344,N_1337);
and U1418 (N_1418,N_1376,N_1384);
xor U1419 (N_1419,N_1372,N_1351);
nor U1420 (N_1420,N_1392,N_1391);
or U1421 (N_1421,N_1320,N_1341);
and U1422 (N_1422,N_1367,N_1368);
nand U1423 (N_1423,N_1398,N_1348);
xnor U1424 (N_1424,N_1377,N_1336);
nand U1425 (N_1425,N_1389,N_1332);
or U1426 (N_1426,N_1380,N_1327);
and U1427 (N_1427,N_1397,N_1306);
and U1428 (N_1428,N_1340,N_1360);
nand U1429 (N_1429,N_1322,N_1373);
xnor U1430 (N_1430,N_1352,N_1362);
xor U1431 (N_1431,N_1314,N_1366);
nor U1432 (N_1432,N_1379,N_1313);
nand U1433 (N_1433,N_1381,N_1330);
nand U1434 (N_1434,N_1357,N_1394);
nor U1435 (N_1435,N_1308,N_1396);
and U1436 (N_1436,N_1304,N_1390);
or U1437 (N_1437,N_1374,N_1359);
nor U1438 (N_1438,N_1315,N_1328);
or U1439 (N_1439,N_1356,N_1339);
or U1440 (N_1440,N_1321,N_1350);
nand U1441 (N_1441,N_1301,N_1346);
nand U1442 (N_1442,N_1318,N_1354);
xor U1443 (N_1443,N_1334,N_1347);
nor U1444 (N_1444,N_1311,N_1399);
nand U1445 (N_1445,N_1317,N_1378);
or U1446 (N_1446,N_1395,N_1329);
nor U1447 (N_1447,N_1364,N_1385);
and U1448 (N_1448,N_1326,N_1353);
xnor U1449 (N_1449,N_1305,N_1312);
nor U1450 (N_1450,N_1314,N_1362);
and U1451 (N_1451,N_1379,N_1360);
xnor U1452 (N_1452,N_1355,N_1321);
xnor U1453 (N_1453,N_1333,N_1370);
or U1454 (N_1454,N_1360,N_1320);
and U1455 (N_1455,N_1353,N_1331);
nand U1456 (N_1456,N_1358,N_1345);
and U1457 (N_1457,N_1368,N_1358);
xnor U1458 (N_1458,N_1360,N_1396);
nor U1459 (N_1459,N_1383,N_1388);
or U1460 (N_1460,N_1378,N_1323);
xor U1461 (N_1461,N_1349,N_1374);
and U1462 (N_1462,N_1373,N_1307);
nand U1463 (N_1463,N_1373,N_1346);
nand U1464 (N_1464,N_1371,N_1327);
and U1465 (N_1465,N_1388,N_1342);
nand U1466 (N_1466,N_1348,N_1304);
and U1467 (N_1467,N_1382,N_1396);
xor U1468 (N_1468,N_1379,N_1325);
xor U1469 (N_1469,N_1311,N_1379);
nand U1470 (N_1470,N_1370,N_1389);
nand U1471 (N_1471,N_1377,N_1382);
and U1472 (N_1472,N_1343,N_1388);
or U1473 (N_1473,N_1303,N_1351);
or U1474 (N_1474,N_1350,N_1318);
nor U1475 (N_1475,N_1312,N_1386);
and U1476 (N_1476,N_1307,N_1354);
and U1477 (N_1477,N_1359,N_1338);
nand U1478 (N_1478,N_1357,N_1393);
nor U1479 (N_1479,N_1365,N_1360);
nor U1480 (N_1480,N_1302,N_1340);
and U1481 (N_1481,N_1370,N_1346);
or U1482 (N_1482,N_1317,N_1395);
and U1483 (N_1483,N_1324,N_1372);
nor U1484 (N_1484,N_1357,N_1343);
nand U1485 (N_1485,N_1326,N_1376);
nand U1486 (N_1486,N_1365,N_1343);
nand U1487 (N_1487,N_1389,N_1352);
nand U1488 (N_1488,N_1313,N_1348);
and U1489 (N_1489,N_1388,N_1355);
and U1490 (N_1490,N_1354,N_1372);
xnor U1491 (N_1491,N_1371,N_1309);
xnor U1492 (N_1492,N_1392,N_1344);
and U1493 (N_1493,N_1368,N_1306);
or U1494 (N_1494,N_1375,N_1346);
nor U1495 (N_1495,N_1369,N_1365);
or U1496 (N_1496,N_1313,N_1393);
nand U1497 (N_1497,N_1329,N_1386);
and U1498 (N_1498,N_1355,N_1324);
nand U1499 (N_1499,N_1348,N_1374);
nor U1500 (N_1500,N_1468,N_1476);
nor U1501 (N_1501,N_1445,N_1402);
nand U1502 (N_1502,N_1469,N_1431);
nor U1503 (N_1503,N_1411,N_1484);
nor U1504 (N_1504,N_1430,N_1444);
nand U1505 (N_1505,N_1494,N_1435);
xor U1506 (N_1506,N_1475,N_1407);
and U1507 (N_1507,N_1425,N_1499);
or U1508 (N_1508,N_1464,N_1483);
and U1509 (N_1509,N_1486,N_1408);
nor U1510 (N_1510,N_1438,N_1471);
nor U1511 (N_1511,N_1418,N_1472);
and U1512 (N_1512,N_1421,N_1406);
nor U1513 (N_1513,N_1432,N_1450);
or U1514 (N_1514,N_1403,N_1416);
nor U1515 (N_1515,N_1496,N_1451);
and U1516 (N_1516,N_1417,N_1466);
or U1517 (N_1517,N_1457,N_1492);
and U1518 (N_1518,N_1482,N_1401);
xnor U1519 (N_1519,N_1428,N_1488);
nor U1520 (N_1520,N_1420,N_1474);
xnor U1521 (N_1521,N_1405,N_1460);
nand U1522 (N_1522,N_1415,N_1493);
or U1523 (N_1523,N_1429,N_1410);
nand U1524 (N_1524,N_1465,N_1487);
nor U1525 (N_1525,N_1427,N_1443);
and U1526 (N_1526,N_1497,N_1462);
xor U1527 (N_1527,N_1478,N_1490);
nand U1528 (N_1528,N_1433,N_1440);
and U1529 (N_1529,N_1470,N_1455);
xnor U1530 (N_1530,N_1419,N_1413);
nor U1531 (N_1531,N_1426,N_1458);
xor U1532 (N_1532,N_1481,N_1452);
xnor U1533 (N_1533,N_1489,N_1449);
nor U1534 (N_1534,N_1477,N_1434);
nor U1535 (N_1535,N_1439,N_1473);
and U1536 (N_1536,N_1479,N_1404);
and U1537 (N_1537,N_1459,N_1454);
xnor U1538 (N_1538,N_1448,N_1414);
or U1539 (N_1539,N_1409,N_1422);
nor U1540 (N_1540,N_1463,N_1423);
xor U1541 (N_1541,N_1446,N_1495);
and U1542 (N_1542,N_1400,N_1498);
nand U1543 (N_1543,N_1412,N_1436);
or U1544 (N_1544,N_1456,N_1467);
nor U1545 (N_1545,N_1453,N_1424);
and U1546 (N_1546,N_1437,N_1485);
and U1547 (N_1547,N_1447,N_1461);
nor U1548 (N_1548,N_1441,N_1491);
or U1549 (N_1549,N_1480,N_1442);
xnor U1550 (N_1550,N_1435,N_1483);
nand U1551 (N_1551,N_1475,N_1464);
xnor U1552 (N_1552,N_1482,N_1437);
xor U1553 (N_1553,N_1403,N_1451);
xor U1554 (N_1554,N_1413,N_1411);
nor U1555 (N_1555,N_1490,N_1426);
nand U1556 (N_1556,N_1458,N_1403);
nor U1557 (N_1557,N_1466,N_1463);
and U1558 (N_1558,N_1439,N_1459);
nor U1559 (N_1559,N_1464,N_1482);
and U1560 (N_1560,N_1444,N_1427);
nand U1561 (N_1561,N_1472,N_1469);
xor U1562 (N_1562,N_1446,N_1458);
xnor U1563 (N_1563,N_1415,N_1401);
xnor U1564 (N_1564,N_1417,N_1457);
nor U1565 (N_1565,N_1459,N_1403);
and U1566 (N_1566,N_1459,N_1458);
nor U1567 (N_1567,N_1481,N_1415);
or U1568 (N_1568,N_1470,N_1439);
xor U1569 (N_1569,N_1495,N_1494);
and U1570 (N_1570,N_1438,N_1476);
xnor U1571 (N_1571,N_1438,N_1466);
nand U1572 (N_1572,N_1456,N_1499);
nor U1573 (N_1573,N_1484,N_1499);
and U1574 (N_1574,N_1472,N_1481);
xnor U1575 (N_1575,N_1452,N_1497);
xnor U1576 (N_1576,N_1414,N_1498);
nor U1577 (N_1577,N_1438,N_1493);
nor U1578 (N_1578,N_1493,N_1433);
nor U1579 (N_1579,N_1488,N_1441);
and U1580 (N_1580,N_1430,N_1424);
or U1581 (N_1581,N_1479,N_1457);
and U1582 (N_1582,N_1415,N_1459);
nand U1583 (N_1583,N_1480,N_1427);
and U1584 (N_1584,N_1464,N_1477);
xnor U1585 (N_1585,N_1443,N_1451);
or U1586 (N_1586,N_1473,N_1485);
nand U1587 (N_1587,N_1485,N_1474);
or U1588 (N_1588,N_1460,N_1434);
or U1589 (N_1589,N_1434,N_1437);
or U1590 (N_1590,N_1445,N_1449);
nand U1591 (N_1591,N_1440,N_1473);
nor U1592 (N_1592,N_1486,N_1478);
and U1593 (N_1593,N_1431,N_1458);
or U1594 (N_1594,N_1456,N_1452);
and U1595 (N_1595,N_1497,N_1469);
xnor U1596 (N_1596,N_1421,N_1480);
nand U1597 (N_1597,N_1467,N_1441);
nand U1598 (N_1598,N_1476,N_1440);
xnor U1599 (N_1599,N_1465,N_1429);
nand U1600 (N_1600,N_1588,N_1556);
nor U1601 (N_1601,N_1536,N_1502);
nand U1602 (N_1602,N_1565,N_1534);
and U1603 (N_1603,N_1597,N_1577);
or U1604 (N_1604,N_1595,N_1566);
nor U1605 (N_1605,N_1561,N_1562);
and U1606 (N_1606,N_1580,N_1503);
or U1607 (N_1607,N_1560,N_1586);
or U1608 (N_1608,N_1598,N_1547);
and U1609 (N_1609,N_1571,N_1579);
or U1610 (N_1610,N_1576,N_1541);
nand U1611 (N_1611,N_1507,N_1587);
or U1612 (N_1612,N_1501,N_1524);
nand U1613 (N_1613,N_1506,N_1505);
and U1614 (N_1614,N_1578,N_1520);
nand U1615 (N_1615,N_1511,N_1510);
nand U1616 (N_1616,N_1526,N_1546);
nand U1617 (N_1617,N_1529,N_1555);
and U1618 (N_1618,N_1512,N_1599);
or U1619 (N_1619,N_1594,N_1581);
nand U1620 (N_1620,N_1533,N_1523);
nand U1621 (N_1621,N_1527,N_1528);
nor U1622 (N_1622,N_1569,N_1532);
xor U1623 (N_1623,N_1517,N_1574);
nor U1624 (N_1624,N_1531,N_1585);
or U1625 (N_1625,N_1545,N_1596);
and U1626 (N_1626,N_1515,N_1550);
nand U1627 (N_1627,N_1537,N_1573);
and U1628 (N_1628,N_1543,N_1544);
and U1629 (N_1629,N_1508,N_1500);
and U1630 (N_1630,N_1554,N_1519);
or U1631 (N_1631,N_1567,N_1570);
or U1632 (N_1632,N_1584,N_1542);
nand U1633 (N_1633,N_1559,N_1589);
and U1634 (N_1634,N_1553,N_1558);
nor U1635 (N_1635,N_1504,N_1590);
xnor U1636 (N_1636,N_1592,N_1557);
nand U1637 (N_1637,N_1513,N_1548);
xnor U1638 (N_1638,N_1591,N_1540);
nor U1639 (N_1639,N_1552,N_1522);
and U1640 (N_1640,N_1521,N_1525);
xor U1641 (N_1641,N_1593,N_1530);
nand U1642 (N_1642,N_1568,N_1583);
xnor U1643 (N_1643,N_1582,N_1516);
xnor U1644 (N_1644,N_1509,N_1551);
xor U1645 (N_1645,N_1539,N_1563);
nor U1646 (N_1646,N_1564,N_1575);
nand U1647 (N_1647,N_1514,N_1535);
nand U1648 (N_1648,N_1538,N_1518);
or U1649 (N_1649,N_1549,N_1572);
nor U1650 (N_1650,N_1558,N_1567);
nand U1651 (N_1651,N_1510,N_1506);
xnor U1652 (N_1652,N_1528,N_1597);
or U1653 (N_1653,N_1565,N_1523);
or U1654 (N_1654,N_1506,N_1589);
nor U1655 (N_1655,N_1534,N_1519);
nor U1656 (N_1656,N_1520,N_1562);
and U1657 (N_1657,N_1579,N_1582);
nand U1658 (N_1658,N_1508,N_1556);
or U1659 (N_1659,N_1505,N_1515);
nand U1660 (N_1660,N_1567,N_1524);
or U1661 (N_1661,N_1510,N_1515);
nand U1662 (N_1662,N_1572,N_1582);
or U1663 (N_1663,N_1548,N_1586);
or U1664 (N_1664,N_1578,N_1576);
or U1665 (N_1665,N_1510,N_1556);
or U1666 (N_1666,N_1534,N_1594);
nor U1667 (N_1667,N_1581,N_1575);
xnor U1668 (N_1668,N_1547,N_1532);
nand U1669 (N_1669,N_1502,N_1581);
or U1670 (N_1670,N_1570,N_1550);
nand U1671 (N_1671,N_1542,N_1548);
or U1672 (N_1672,N_1597,N_1529);
xnor U1673 (N_1673,N_1504,N_1531);
nand U1674 (N_1674,N_1577,N_1557);
nor U1675 (N_1675,N_1537,N_1584);
or U1676 (N_1676,N_1536,N_1573);
xnor U1677 (N_1677,N_1542,N_1523);
nand U1678 (N_1678,N_1539,N_1528);
nor U1679 (N_1679,N_1544,N_1532);
or U1680 (N_1680,N_1542,N_1517);
or U1681 (N_1681,N_1592,N_1512);
xnor U1682 (N_1682,N_1550,N_1587);
nand U1683 (N_1683,N_1573,N_1515);
and U1684 (N_1684,N_1562,N_1560);
and U1685 (N_1685,N_1587,N_1537);
nor U1686 (N_1686,N_1503,N_1578);
nand U1687 (N_1687,N_1583,N_1535);
nor U1688 (N_1688,N_1590,N_1519);
xnor U1689 (N_1689,N_1542,N_1518);
nand U1690 (N_1690,N_1575,N_1598);
xnor U1691 (N_1691,N_1550,N_1541);
or U1692 (N_1692,N_1508,N_1582);
nor U1693 (N_1693,N_1544,N_1558);
nand U1694 (N_1694,N_1568,N_1537);
nand U1695 (N_1695,N_1512,N_1568);
and U1696 (N_1696,N_1532,N_1545);
and U1697 (N_1697,N_1585,N_1565);
xor U1698 (N_1698,N_1595,N_1544);
or U1699 (N_1699,N_1546,N_1579);
nor U1700 (N_1700,N_1686,N_1608);
and U1701 (N_1701,N_1620,N_1676);
nor U1702 (N_1702,N_1646,N_1654);
xnor U1703 (N_1703,N_1671,N_1662);
xor U1704 (N_1704,N_1634,N_1606);
or U1705 (N_1705,N_1688,N_1651);
nand U1706 (N_1706,N_1682,N_1623);
xor U1707 (N_1707,N_1653,N_1603);
or U1708 (N_1708,N_1655,N_1641);
nand U1709 (N_1709,N_1618,N_1685);
nand U1710 (N_1710,N_1681,N_1638);
or U1711 (N_1711,N_1677,N_1628);
and U1712 (N_1712,N_1664,N_1615);
or U1713 (N_1713,N_1674,N_1666);
nor U1714 (N_1714,N_1683,N_1692);
and U1715 (N_1715,N_1601,N_1696);
and U1716 (N_1716,N_1609,N_1699);
and U1717 (N_1717,N_1652,N_1656);
nand U1718 (N_1718,N_1607,N_1659);
nor U1719 (N_1719,N_1631,N_1643);
nor U1720 (N_1720,N_1629,N_1624);
xor U1721 (N_1721,N_1649,N_1695);
nand U1722 (N_1722,N_1660,N_1689);
nor U1723 (N_1723,N_1658,N_1669);
xnor U1724 (N_1724,N_1622,N_1698);
nor U1725 (N_1725,N_1667,N_1625);
and U1726 (N_1726,N_1627,N_1687);
or U1727 (N_1727,N_1697,N_1665);
nor U1728 (N_1728,N_1680,N_1670);
xnor U1729 (N_1729,N_1675,N_1610);
and U1730 (N_1730,N_1626,N_1645);
xor U1731 (N_1731,N_1668,N_1611);
or U1732 (N_1732,N_1600,N_1690);
or U1733 (N_1733,N_1616,N_1693);
or U1734 (N_1734,N_1642,N_1640);
nor U1735 (N_1735,N_1647,N_1691);
or U1736 (N_1736,N_1614,N_1619);
nand U1737 (N_1737,N_1644,N_1605);
nand U1738 (N_1738,N_1684,N_1657);
nand U1739 (N_1739,N_1679,N_1621);
xor U1740 (N_1740,N_1613,N_1630);
nand U1741 (N_1741,N_1694,N_1636);
and U1742 (N_1742,N_1632,N_1637);
xor U1743 (N_1743,N_1678,N_1639);
nand U1744 (N_1744,N_1673,N_1663);
xor U1745 (N_1745,N_1672,N_1648);
or U1746 (N_1746,N_1635,N_1650);
xor U1747 (N_1747,N_1612,N_1604);
xnor U1748 (N_1748,N_1602,N_1661);
xor U1749 (N_1749,N_1633,N_1617);
and U1750 (N_1750,N_1640,N_1630);
nor U1751 (N_1751,N_1640,N_1641);
nor U1752 (N_1752,N_1606,N_1654);
or U1753 (N_1753,N_1698,N_1626);
nand U1754 (N_1754,N_1620,N_1697);
nand U1755 (N_1755,N_1679,N_1664);
nand U1756 (N_1756,N_1659,N_1617);
nand U1757 (N_1757,N_1661,N_1680);
xor U1758 (N_1758,N_1640,N_1647);
or U1759 (N_1759,N_1625,N_1669);
nand U1760 (N_1760,N_1634,N_1677);
or U1761 (N_1761,N_1631,N_1674);
nand U1762 (N_1762,N_1694,N_1686);
xnor U1763 (N_1763,N_1668,N_1654);
nor U1764 (N_1764,N_1673,N_1660);
xnor U1765 (N_1765,N_1657,N_1661);
nand U1766 (N_1766,N_1687,N_1691);
and U1767 (N_1767,N_1643,N_1615);
or U1768 (N_1768,N_1627,N_1617);
or U1769 (N_1769,N_1675,N_1608);
or U1770 (N_1770,N_1602,N_1684);
xor U1771 (N_1771,N_1615,N_1629);
and U1772 (N_1772,N_1613,N_1611);
xnor U1773 (N_1773,N_1626,N_1667);
or U1774 (N_1774,N_1637,N_1696);
or U1775 (N_1775,N_1688,N_1678);
xor U1776 (N_1776,N_1693,N_1661);
or U1777 (N_1777,N_1688,N_1633);
xnor U1778 (N_1778,N_1645,N_1652);
nor U1779 (N_1779,N_1626,N_1631);
nor U1780 (N_1780,N_1698,N_1660);
or U1781 (N_1781,N_1609,N_1659);
or U1782 (N_1782,N_1646,N_1649);
xor U1783 (N_1783,N_1642,N_1692);
nor U1784 (N_1784,N_1687,N_1666);
xor U1785 (N_1785,N_1659,N_1624);
xnor U1786 (N_1786,N_1631,N_1661);
nand U1787 (N_1787,N_1614,N_1604);
and U1788 (N_1788,N_1618,N_1642);
nor U1789 (N_1789,N_1665,N_1691);
nor U1790 (N_1790,N_1642,N_1622);
nor U1791 (N_1791,N_1647,N_1616);
and U1792 (N_1792,N_1627,N_1690);
and U1793 (N_1793,N_1678,N_1656);
xnor U1794 (N_1794,N_1685,N_1674);
or U1795 (N_1795,N_1653,N_1652);
xor U1796 (N_1796,N_1654,N_1635);
or U1797 (N_1797,N_1678,N_1619);
xor U1798 (N_1798,N_1630,N_1691);
or U1799 (N_1799,N_1649,N_1696);
or U1800 (N_1800,N_1729,N_1744);
xnor U1801 (N_1801,N_1755,N_1715);
or U1802 (N_1802,N_1716,N_1773);
or U1803 (N_1803,N_1775,N_1736);
nand U1804 (N_1804,N_1751,N_1771);
or U1805 (N_1805,N_1790,N_1732);
nand U1806 (N_1806,N_1740,N_1709);
nor U1807 (N_1807,N_1797,N_1798);
or U1808 (N_1808,N_1769,N_1723);
and U1809 (N_1809,N_1741,N_1708);
or U1810 (N_1810,N_1792,N_1737);
nand U1811 (N_1811,N_1784,N_1789);
nor U1812 (N_1812,N_1743,N_1786);
nor U1813 (N_1813,N_1731,N_1712);
nand U1814 (N_1814,N_1787,N_1756);
nand U1815 (N_1815,N_1721,N_1765);
xor U1816 (N_1816,N_1754,N_1714);
nand U1817 (N_1817,N_1794,N_1718);
or U1818 (N_1818,N_1700,N_1703);
nor U1819 (N_1819,N_1702,N_1759);
and U1820 (N_1820,N_1763,N_1725);
or U1821 (N_1821,N_1776,N_1779);
xnor U1822 (N_1822,N_1760,N_1717);
or U1823 (N_1823,N_1758,N_1722);
or U1824 (N_1824,N_1752,N_1706);
or U1825 (N_1825,N_1739,N_1750);
or U1826 (N_1826,N_1753,N_1710);
or U1827 (N_1827,N_1746,N_1757);
xnor U1828 (N_1828,N_1730,N_1796);
and U1829 (N_1829,N_1793,N_1772);
nand U1830 (N_1830,N_1745,N_1747);
xor U1831 (N_1831,N_1768,N_1782);
nand U1832 (N_1832,N_1707,N_1704);
or U1833 (N_1833,N_1781,N_1761);
or U1834 (N_1834,N_1711,N_1701);
xnor U1835 (N_1835,N_1795,N_1735);
nor U1836 (N_1836,N_1766,N_1778);
or U1837 (N_1837,N_1705,N_1713);
nor U1838 (N_1838,N_1726,N_1742);
xnor U1839 (N_1839,N_1749,N_1762);
nand U1840 (N_1840,N_1777,N_1799);
nand U1841 (N_1841,N_1764,N_1767);
nand U1842 (N_1842,N_1727,N_1783);
nand U1843 (N_1843,N_1791,N_1728);
nand U1844 (N_1844,N_1720,N_1774);
or U1845 (N_1845,N_1788,N_1733);
and U1846 (N_1846,N_1738,N_1724);
nand U1847 (N_1847,N_1734,N_1748);
or U1848 (N_1848,N_1780,N_1719);
nor U1849 (N_1849,N_1785,N_1770);
xnor U1850 (N_1850,N_1797,N_1718);
or U1851 (N_1851,N_1781,N_1786);
xnor U1852 (N_1852,N_1755,N_1791);
nand U1853 (N_1853,N_1773,N_1753);
xnor U1854 (N_1854,N_1799,N_1747);
and U1855 (N_1855,N_1783,N_1719);
nor U1856 (N_1856,N_1763,N_1788);
and U1857 (N_1857,N_1737,N_1780);
nor U1858 (N_1858,N_1712,N_1749);
nor U1859 (N_1859,N_1751,N_1704);
xnor U1860 (N_1860,N_1700,N_1763);
xor U1861 (N_1861,N_1741,N_1767);
nand U1862 (N_1862,N_1739,N_1726);
nor U1863 (N_1863,N_1715,N_1772);
nand U1864 (N_1864,N_1709,N_1759);
nand U1865 (N_1865,N_1709,N_1701);
and U1866 (N_1866,N_1719,N_1770);
and U1867 (N_1867,N_1733,N_1705);
and U1868 (N_1868,N_1783,N_1735);
and U1869 (N_1869,N_1797,N_1764);
nand U1870 (N_1870,N_1772,N_1776);
xor U1871 (N_1871,N_1752,N_1789);
and U1872 (N_1872,N_1777,N_1728);
or U1873 (N_1873,N_1780,N_1716);
nand U1874 (N_1874,N_1718,N_1771);
xnor U1875 (N_1875,N_1777,N_1785);
nor U1876 (N_1876,N_1755,N_1770);
and U1877 (N_1877,N_1776,N_1725);
nor U1878 (N_1878,N_1781,N_1762);
or U1879 (N_1879,N_1723,N_1724);
and U1880 (N_1880,N_1795,N_1710);
or U1881 (N_1881,N_1772,N_1741);
nand U1882 (N_1882,N_1765,N_1774);
or U1883 (N_1883,N_1799,N_1733);
and U1884 (N_1884,N_1788,N_1715);
nor U1885 (N_1885,N_1797,N_1714);
xor U1886 (N_1886,N_1716,N_1786);
nand U1887 (N_1887,N_1755,N_1753);
nand U1888 (N_1888,N_1782,N_1773);
or U1889 (N_1889,N_1713,N_1729);
xnor U1890 (N_1890,N_1766,N_1709);
and U1891 (N_1891,N_1730,N_1725);
nand U1892 (N_1892,N_1742,N_1735);
and U1893 (N_1893,N_1717,N_1782);
nor U1894 (N_1894,N_1755,N_1771);
nand U1895 (N_1895,N_1735,N_1731);
nor U1896 (N_1896,N_1704,N_1722);
nand U1897 (N_1897,N_1767,N_1742);
nand U1898 (N_1898,N_1799,N_1794);
and U1899 (N_1899,N_1784,N_1706);
nand U1900 (N_1900,N_1850,N_1854);
and U1901 (N_1901,N_1873,N_1829);
or U1902 (N_1902,N_1853,N_1820);
xor U1903 (N_1903,N_1805,N_1828);
nand U1904 (N_1904,N_1885,N_1832);
nand U1905 (N_1905,N_1830,N_1834);
nor U1906 (N_1906,N_1889,N_1865);
nor U1907 (N_1907,N_1875,N_1899);
nor U1908 (N_1908,N_1874,N_1855);
nand U1909 (N_1909,N_1877,N_1871);
and U1910 (N_1910,N_1821,N_1809);
or U1911 (N_1911,N_1860,N_1851);
and U1912 (N_1912,N_1822,N_1815);
or U1913 (N_1913,N_1879,N_1825);
xor U1914 (N_1914,N_1849,N_1859);
nor U1915 (N_1915,N_1886,N_1861);
nand U1916 (N_1916,N_1883,N_1802);
nand U1917 (N_1917,N_1807,N_1831);
or U1918 (N_1918,N_1887,N_1856);
and U1919 (N_1919,N_1880,N_1840);
nor U1920 (N_1920,N_1866,N_1824);
or U1921 (N_1921,N_1813,N_1898);
nor U1922 (N_1922,N_1836,N_1819);
xor U1923 (N_1923,N_1839,N_1843);
nand U1924 (N_1924,N_1838,N_1846);
xor U1925 (N_1925,N_1882,N_1841);
or U1926 (N_1926,N_1800,N_1893);
nand U1927 (N_1927,N_1801,N_1894);
nand U1928 (N_1928,N_1848,N_1867);
nor U1929 (N_1929,N_1895,N_1896);
or U1930 (N_1930,N_1844,N_1858);
or U1931 (N_1931,N_1810,N_1847);
or U1932 (N_1932,N_1868,N_1876);
or U1933 (N_1933,N_1845,N_1827);
or U1934 (N_1934,N_1857,N_1806);
or U1935 (N_1935,N_1891,N_1814);
and U1936 (N_1936,N_1878,N_1842);
xnor U1937 (N_1937,N_1835,N_1863);
nand U1938 (N_1938,N_1837,N_1888);
or U1939 (N_1939,N_1872,N_1881);
xnor U1940 (N_1940,N_1817,N_1833);
or U1941 (N_1941,N_1816,N_1897);
nand U1942 (N_1942,N_1803,N_1808);
nor U1943 (N_1943,N_1890,N_1862);
nand U1944 (N_1944,N_1892,N_1852);
or U1945 (N_1945,N_1826,N_1812);
xnor U1946 (N_1946,N_1884,N_1818);
nand U1947 (N_1947,N_1823,N_1870);
and U1948 (N_1948,N_1811,N_1864);
or U1949 (N_1949,N_1804,N_1869);
xor U1950 (N_1950,N_1815,N_1890);
xor U1951 (N_1951,N_1857,N_1851);
or U1952 (N_1952,N_1808,N_1894);
xor U1953 (N_1953,N_1836,N_1830);
nand U1954 (N_1954,N_1844,N_1805);
nand U1955 (N_1955,N_1849,N_1891);
xnor U1956 (N_1956,N_1857,N_1821);
xor U1957 (N_1957,N_1813,N_1855);
nand U1958 (N_1958,N_1804,N_1859);
nand U1959 (N_1959,N_1878,N_1829);
nand U1960 (N_1960,N_1869,N_1866);
or U1961 (N_1961,N_1825,N_1841);
and U1962 (N_1962,N_1844,N_1814);
nor U1963 (N_1963,N_1882,N_1815);
nand U1964 (N_1964,N_1845,N_1889);
nor U1965 (N_1965,N_1838,N_1843);
nand U1966 (N_1966,N_1810,N_1835);
nand U1967 (N_1967,N_1845,N_1833);
nand U1968 (N_1968,N_1848,N_1803);
xnor U1969 (N_1969,N_1827,N_1864);
nor U1970 (N_1970,N_1875,N_1807);
and U1971 (N_1971,N_1804,N_1828);
and U1972 (N_1972,N_1811,N_1806);
nor U1973 (N_1973,N_1898,N_1873);
nor U1974 (N_1974,N_1805,N_1872);
nor U1975 (N_1975,N_1891,N_1897);
nor U1976 (N_1976,N_1849,N_1871);
nor U1977 (N_1977,N_1858,N_1834);
or U1978 (N_1978,N_1857,N_1870);
or U1979 (N_1979,N_1851,N_1825);
or U1980 (N_1980,N_1804,N_1857);
xor U1981 (N_1981,N_1882,N_1860);
xor U1982 (N_1982,N_1809,N_1803);
nor U1983 (N_1983,N_1812,N_1810);
nor U1984 (N_1984,N_1866,N_1810);
nor U1985 (N_1985,N_1857,N_1897);
xnor U1986 (N_1986,N_1896,N_1868);
xor U1987 (N_1987,N_1895,N_1838);
or U1988 (N_1988,N_1897,N_1848);
and U1989 (N_1989,N_1878,N_1868);
nor U1990 (N_1990,N_1822,N_1894);
or U1991 (N_1991,N_1841,N_1877);
xor U1992 (N_1992,N_1854,N_1855);
nor U1993 (N_1993,N_1870,N_1893);
and U1994 (N_1994,N_1840,N_1811);
nor U1995 (N_1995,N_1842,N_1873);
and U1996 (N_1996,N_1814,N_1890);
or U1997 (N_1997,N_1812,N_1862);
or U1998 (N_1998,N_1827,N_1892);
nand U1999 (N_1999,N_1820,N_1880);
nor U2000 (N_2000,N_1904,N_1930);
and U2001 (N_2001,N_1979,N_1957);
nand U2002 (N_2002,N_1919,N_1909);
xor U2003 (N_2003,N_1968,N_1991);
and U2004 (N_2004,N_1961,N_1900);
nand U2005 (N_2005,N_1948,N_1976);
nor U2006 (N_2006,N_1972,N_1921);
nand U2007 (N_2007,N_1906,N_1995);
or U2008 (N_2008,N_1944,N_1973);
xnor U2009 (N_2009,N_1999,N_1902);
nand U2010 (N_2010,N_1931,N_1971);
nor U2011 (N_2011,N_1946,N_1916);
or U2012 (N_2012,N_1990,N_1911);
xor U2013 (N_2013,N_1974,N_1914);
and U2014 (N_2014,N_1994,N_1942);
nor U2015 (N_2015,N_1963,N_1955);
nand U2016 (N_2016,N_1927,N_1966);
nand U2017 (N_2017,N_1980,N_1934);
xnor U2018 (N_2018,N_1901,N_1907);
nor U2019 (N_2019,N_1924,N_1981);
nor U2020 (N_2020,N_1967,N_1939);
nor U2021 (N_2021,N_1958,N_1915);
nand U2022 (N_2022,N_1962,N_1970);
or U2023 (N_2023,N_1964,N_1996);
and U2024 (N_2024,N_1985,N_1959);
and U2025 (N_2025,N_1936,N_1913);
or U2026 (N_2026,N_1926,N_1956);
nand U2027 (N_2027,N_1960,N_1943);
nor U2028 (N_2028,N_1953,N_1992);
nand U2029 (N_2029,N_1928,N_1978);
xnor U2030 (N_2030,N_1989,N_1952);
nor U2031 (N_2031,N_1984,N_1938);
nor U2032 (N_2032,N_1940,N_1951);
nand U2033 (N_2033,N_1933,N_1993);
and U2034 (N_2034,N_1923,N_1932);
xor U2035 (N_2035,N_1969,N_1949);
and U2036 (N_2036,N_1950,N_1917);
and U2037 (N_2037,N_1998,N_1997);
nand U2038 (N_2038,N_1941,N_1935);
or U2039 (N_2039,N_1925,N_1920);
or U2040 (N_2040,N_1918,N_1912);
or U2041 (N_2041,N_1905,N_1986);
nand U2042 (N_2042,N_1983,N_1987);
nor U2043 (N_2043,N_1908,N_1947);
nand U2044 (N_2044,N_1937,N_1922);
and U2045 (N_2045,N_1982,N_1975);
nor U2046 (N_2046,N_1954,N_1988);
nor U2047 (N_2047,N_1945,N_1929);
xor U2048 (N_2048,N_1903,N_1910);
and U2049 (N_2049,N_1965,N_1977);
nor U2050 (N_2050,N_1953,N_1982);
nor U2051 (N_2051,N_1917,N_1932);
nand U2052 (N_2052,N_1984,N_1937);
nand U2053 (N_2053,N_1947,N_1997);
xnor U2054 (N_2054,N_1975,N_1909);
or U2055 (N_2055,N_1988,N_1943);
nor U2056 (N_2056,N_1955,N_1958);
nand U2057 (N_2057,N_1966,N_1902);
or U2058 (N_2058,N_1921,N_1951);
nor U2059 (N_2059,N_1936,N_1926);
or U2060 (N_2060,N_1991,N_1951);
and U2061 (N_2061,N_1989,N_1901);
and U2062 (N_2062,N_1972,N_1941);
xor U2063 (N_2063,N_1983,N_1957);
and U2064 (N_2064,N_1903,N_1930);
or U2065 (N_2065,N_1904,N_1952);
nand U2066 (N_2066,N_1977,N_1969);
nand U2067 (N_2067,N_1993,N_1950);
nand U2068 (N_2068,N_1994,N_1991);
and U2069 (N_2069,N_1908,N_1933);
and U2070 (N_2070,N_1981,N_1960);
nand U2071 (N_2071,N_1999,N_1979);
nor U2072 (N_2072,N_1914,N_1949);
nand U2073 (N_2073,N_1977,N_1950);
or U2074 (N_2074,N_1966,N_1951);
xor U2075 (N_2075,N_1902,N_1920);
or U2076 (N_2076,N_1900,N_1903);
xor U2077 (N_2077,N_1956,N_1965);
xnor U2078 (N_2078,N_1902,N_1981);
xnor U2079 (N_2079,N_1925,N_1949);
nand U2080 (N_2080,N_1908,N_1990);
nand U2081 (N_2081,N_1990,N_1920);
or U2082 (N_2082,N_1996,N_1917);
or U2083 (N_2083,N_1937,N_1955);
nor U2084 (N_2084,N_1945,N_1934);
and U2085 (N_2085,N_1971,N_1944);
or U2086 (N_2086,N_1904,N_1911);
nor U2087 (N_2087,N_1947,N_1963);
and U2088 (N_2088,N_1931,N_1973);
xor U2089 (N_2089,N_1958,N_1902);
xnor U2090 (N_2090,N_1955,N_1979);
or U2091 (N_2091,N_1950,N_1945);
nand U2092 (N_2092,N_1904,N_1954);
xor U2093 (N_2093,N_1922,N_1960);
nand U2094 (N_2094,N_1956,N_1981);
nor U2095 (N_2095,N_1918,N_1919);
nor U2096 (N_2096,N_1995,N_1982);
or U2097 (N_2097,N_1915,N_1959);
nor U2098 (N_2098,N_1957,N_1904);
and U2099 (N_2099,N_1979,N_1922);
and U2100 (N_2100,N_2006,N_2091);
nand U2101 (N_2101,N_2004,N_2053);
or U2102 (N_2102,N_2052,N_2084);
nand U2103 (N_2103,N_2062,N_2026);
nor U2104 (N_2104,N_2032,N_2047);
nand U2105 (N_2105,N_2058,N_2021);
and U2106 (N_2106,N_2075,N_2005);
nor U2107 (N_2107,N_2056,N_2033);
xor U2108 (N_2108,N_2028,N_2012);
nand U2109 (N_2109,N_2001,N_2027);
and U2110 (N_2110,N_2083,N_2017);
nor U2111 (N_2111,N_2080,N_2040);
and U2112 (N_2112,N_2081,N_2029);
and U2113 (N_2113,N_2013,N_2000);
xnor U2114 (N_2114,N_2014,N_2009);
nand U2115 (N_2115,N_2041,N_2044);
and U2116 (N_2116,N_2071,N_2036);
and U2117 (N_2117,N_2070,N_2007);
xor U2118 (N_2118,N_2085,N_2097);
or U2119 (N_2119,N_2066,N_2099);
xor U2120 (N_2120,N_2074,N_2020);
xnor U2121 (N_2121,N_2060,N_2077);
or U2122 (N_2122,N_2098,N_2061);
nor U2123 (N_2123,N_2054,N_2087);
xor U2124 (N_2124,N_2031,N_2048);
and U2125 (N_2125,N_2049,N_2023);
nor U2126 (N_2126,N_2016,N_2069);
and U2127 (N_2127,N_2025,N_2059);
nand U2128 (N_2128,N_2008,N_2043);
nand U2129 (N_2129,N_2078,N_2042);
nor U2130 (N_2130,N_2096,N_2055);
nor U2131 (N_2131,N_2022,N_2090);
nand U2132 (N_2132,N_2092,N_2057);
nand U2133 (N_2133,N_2073,N_2038);
nor U2134 (N_2134,N_2045,N_2067);
nand U2135 (N_2135,N_2051,N_2018);
nand U2136 (N_2136,N_2068,N_2037);
and U2137 (N_2137,N_2065,N_2046);
and U2138 (N_2138,N_2072,N_2063);
or U2139 (N_2139,N_2003,N_2019);
and U2140 (N_2140,N_2094,N_2095);
and U2141 (N_2141,N_2082,N_2030);
and U2142 (N_2142,N_2034,N_2050);
or U2143 (N_2143,N_2093,N_2088);
xor U2144 (N_2144,N_2039,N_2010);
nand U2145 (N_2145,N_2079,N_2064);
nand U2146 (N_2146,N_2024,N_2076);
xor U2147 (N_2147,N_2089,N_2002);
nor U2148 (N_2148,N_2035,N_2011);
xor U2149 (N_2149,N_2015,N_2086);
nand U2150 (N_2150,N_2095,N_2049);
xor U2151 (N_2151,N_2016,N_2083);
xor U2152 (N_2152,N_2043,N_2094);
and U2153 (N_2153,N_2064,N_2056);
nor U2154 (N_2154,N_2031,N_2050);
or U2155 (N_2155,N_2022,N_2038);
xor U2156 (N_2156,N_2054,N_2014);
or U2157 (N_2157,N_2072,N_2087);
nand U2158 (N_2158,N_2024,N_2064);
and U2159 (N_2159,N_2067,N_2033);
or U2160 (N_2160,N_2094,N_2028);
nor U2161 (N_2161,N_2068,N_2002);
and U2162 (N_2162,N_2010,N_2052);
nor U2163 (N_2163,N_2082,N_2016);
or U2164 (N_2164,N_2005,N_2089);
or U2165 (N_2165,N_2039,N_2088);
and U2166 (N_2166,N_2076,N_2061);
nand U2167 (N_2167,N_2099,N_2037);
and U2168 (N_2168,N_2021,N_2063);
xnor U2169 (N_2169,N_2029,N_2051);
and U2170 (N_2170,N_2041,N_2052);
nor U2171 (N_2171,N_2084,N_2029);
and U2172 (N_2172,N_2033,N_2093);
xnor U2173 (N_2173,N_2056,N_2024);
and U2174 (N_2174,N_2084,N_2035);
or U2175 (N_2175,N_2074,N_2085);
nand U2176 (N_2176,N_2068,N_2024);
nand U2177 (N_2177,N_2023,N_2017);
nand U2178 (N_2178,N_2085,N_2042);
or U2179 (N_2179,N_2081,N_2049);
or U2180 (N_2180,N_2086,N_2066);
or U2181 (N_2181,N_2074,N_2099);
or U2182 (N_2182,N_2015,N_2069);
xnor U2183 (N_2183,N_2071,N_2091);
and U2184 (N_2184,N_2065,N_2099);
nor U2185 (N_2185,N_2055,N_2004);
or U2186 (N_2186,N_2059,N_2019);
nand U2187 (N_2187,N_2003,N_2064);
nand U2188 (N_2188,N_2056,N_2072);
nor U2189 (N_2189,N_2043,N_2000);
nor U2190 (N_2190,N_2005,N_2088);
or U2191 (N_2191,N_2077,N_2087);
nor U2192 (N_2192,N_2090,N_2086);
nor U2193 (N_2193,N_2060,N_2079);
or U2194 (N_2194,N_2038,N_2059);
xnor U2195 (N_2195,N_2059,N_2032);
and U2196 (N_2196,N_2027,N_2039);
nor U2197 (N_2197,N_2009,N_2079);
nand U2198 (N_2198,N_2028,N_2048);
or U2199 (N_2199,N_2061,N_2009);
nand U2200 (N_2200,N_2167,N_2158);
nor U2201 (N_2201,N_2171,N_2134);
nor U2202 (N_2202,N_2152,N_2156);
nand U2203 (N_2203,N_2194,N_2132);
nand U2204 (N_2204,N_2177,N_2175);
nand U2205 (N_2205,N_2192,N_2127);
nand U2206 (N_2206,N_2115,N_2124);
xnor U2207 (N_2207,N_2197,N_2146);
nor U2208 (N_2208,N_2117,N_2174);
xnor U2209 (N_2209,N_2114,N_2154);
nor U2210 (N_2210,N_2170,N_2136);
and U2211 (N_2211,N_2104,N_2148);
nor U2212 (N_2212,N_2122,N_2107);
or U2213 (N_2213,N_2149,N_2165);
nor U2214 (N_2214,N_2179,N_2160);
or U2215 (N_2215,N_2186,N_2102);
nor U2216 (N_2216,N_2153,N_2187);
or U2217 (N_2217,N_2119,N_2188);
and U2218 (N_2218,N_2144,N_2106);
xnor U2219 (N_2219,N_2181,N_2199);
or U2220 (N_2220,N_2129,N_2176);
and U2221 (N_2221,N_2196,N_2100);
xnor U2222 (N_2222,N_2183,N_2128);
nand U2223 (N_2223,N_2161,N_2121);
nand U2224 (N_2224,N_2111,N_2189);
or U2225 (N_2225,N_2169,N_2178);
and U2226 (N_2226,N_2162,N_2166);
and U2227 (N_2227,N_2101,N_2142);
and U2228 (N_2228,N_2164,N_2140);
and U2229 (N_2229,N_2130,N_2193);
nand U2230 (N_2230,N_2113,N_2123);
xor U2231 (N_2231,N_2185,N_2191);
xnor U2232 (N_2232,N_2184,N_2110);
nand U2233 (N_2233,N_2147,N_2141);
nand U2234 (N_2234,N_2180,N_2112);
and U2235 (N_2235,N_2139,N_2109);
or U2236 (N_2236,N_2120,N_2157);
or U2237 (N_2237,N_2143,N_2135);
or U2238 (N_2238,N_2150,N_2126);
nand U2239 (N_2239,N_2159,N_2105);
nor U2240 (N_2240,N_2137,N_2172);
xor U2241 (N_2241,N_2182,N_2125);
and U2242 (N_2242,N_2168,N_2155);
or U2243 (N_2243,N_2163,N_2151);
xor U2244 (N_2244,N_2198,N_2131);
nand U2245 (N_2245,N_2195,N_2133);
nor U2246 (N_2246,N_2190,N_2118);
xor U2247 (N_2247,N_2103,N_2138);
nor U2248 (N_2248,N_2116,N_2145);
xor U2249 (N_2249,N_2108,N_2173);
nor U2250 (N_2250,N_2172,N_2155);
and U2251 (N_2251,N_2188,N_2169);
nor U2252 (N_2252,N_2137,N_2180);
nor U2253 (N_2253,N_2165,N_2197);
xor U2254 (N_2254,N_2126,N_2155);
xnor U2255 (N_2255,N_2176,N_2107);
nor U2256 (N_2256,N_2175,N_2135);
and U2257 (N_2257,N_2140,N_2117);
nand U2258 (N_2258,N_2134,N_2195);
or U2259 (N_2259,N_2155,N_2141);
and U2260 (N_2260,N_2166,N_2165);
and U2261 (N_2261,N_2145,N_2196);
and U2262 (N_2262,N_2117,N_2199);
nor U2263 (N_2263,N_2138,N_2154);
nand U2264 (N_2264,N_2105,N_2149);
xor U2265 (N_2265,N_2138,N_2130);
and U2266 (N_2266,N_2151,N_2111);
or U2267 (N_2267,N_2125,N_2155);
xor U2268 (N_2268,N_2127,N_2133);
or U2269 (N_2269,N_2102,N_2155);
xor U2270 (N_2270,N_2171,N_2123);
and U2271 (N_2271,N_2149,N_2191);
or U2272 (N_2272,N_2150,N_2154);
nand U2273 (N_2273,N_2192,N_2111);
nand U2274 (N_2274,N_2191,N_2177);
or U2275 (N_2275,N_2110,N_2174);
and U2276 (N_2276,N_2116,N_2187);
nor U2277 (N_2277,N_2138,N_2173);
and U2278 (N_2278,N_2196,N_2112);
nand U2279 (N_2279,N_2171,N_2112);
and U2280 (N_2280,N_2148,N_2183);
and U2281 (N_2281,N_2151,N_2120);
nand U2282 (N_2282,N_2152,N_2145);
or U2283 (N_2283,N_2160,N_2123);
xnor U2284 (N_2284,N_2106,N_2171);
xor U2285 (N_2285,N_2134,N_2196);
and U2286 (N_2286,N_2183,N_2154);
nor U2287 (N_2287,N_2148,N_2154);
nand U2288 (N_2288,N_2169,N_2119);
nand U2289 (N_2289,N_2152,N_2161);
and U2290 (N_2290,N_2136,N_2112);
nand U2291 (N_2291,N_2123,N_2140);
nand U2292 (N_2292,N_2148,N_2121);
and U2293 (N_2293,N_2107,N_2108);
nand U2294 (N_2294,N_2142,N_2199);
or U2295 (N_2295,N_2150,N_2196);
xor U2296 (N_2296,N_2112,N_2146);
nand U2297 (N_2297,N_2168,N_2132);
nor U2298 (N_2298,N_2138,N_2132);
xnor U2299 (N_2299,N_2115,N_2100);
xor U2300 (N_2300,N_2249,N_2259);
or U2301 (N_2301,N_2228,N_2296);
or U2302 (N_2302,N_2251,N_2248);
nand U2303 (N_2303,N_2204,N_2212);
nand U2304 (N_2304,N_2257,N_2292);
or U2305 (N_2305,N_2239,N_2253);
nand U2306 (N_2306,N_2234,N_2269);
nand U2307 (N_2307,N_2207,N_2277);
nand U2308 (N_2308,N_2214,N_2287);
nand U2309 (N_2309,N_2232,N_2201);
or U2310 (N_2310,N_2222,N_2273);
nand U2311 (N_2311,N_2261,N_2299);
nor U2312 (N_2312,N_2235,N_2274);
nor U2313 (N_2313,N_2283,N_2284);
nand U2314 (N_2314,N_2268,N_2293);
nor U2315 (N_2315,N_2267,N_2262);
and U2316 (N_2316,N_2294,N_2245);
or U2317 (N_2317,N_2250,N_2209);
and U2318 (N_2318,N_2221,N_2297);
nor U2319 (N_2319,N_2295,N_2264);
or U2320 (N_2320,N_2219,N_2282);
or U2321 (N_2321,N_2203,N_2237);
nand U2322 (N_2322,N_2243,N_2242);
nor U2323 (N_2323,N_2276,N_2260);
and U2324 (N_2324,N_2210,N_2263);
or U2325 (N_2325,N_2233,N_2240);
or U2326 (N_2326,N_2208,N_2255);
xnor U2327 (N_2327,N_2247,N_2241);
nand U2328 (N_2328,N_2216,N_2224);
xor U2329 (N_2329,N_2225,N_2217);
xor U2330 (N_2330,N_2280,N_2231);
and U2331 (N_2331,N_2200,N_2278);
nor U2332 (N_2332,N_2246,N_2215);
xnor U2333 (N_2333,N_2272,N_2265);
nand U2334 (N_2334,N_2244,N_2206);
and U2335 (N_2335,N_2220,N_2202);
and U2336 (N_2336,N_2298,N_2238);
and U2337 (N_2337,N_2291,N_2211);
nand U2338 (N_2338,N_2229,N_2271);
nand U2339 (N_2339,N_2254,N_2236);
nand U2340 (N_2340,N_2252,N_2285);
and U2341 (N_2341,N_2288,N_2258);
nor U2342 (N_2342,N_2281,N_2290);
or U2343 (N_2343,N_2218,N_2270);
and U2344 (N_2344,N_2266,N_2289);
nand U2345 (N_2345,N_2230,N_2286);
xnor U2346 (N_2346,N_2256,N_2223);
and U2347 (N_2347,N_2205,N_2226);
xnor U2348 (N_2348,N_2279,N_2275);
nand U2349 (N_2349,N_2213,N_2227);
and U2350 (N_2350,N_2215,N_2254);
xnor U2351 (N_2351,N_2216,N_2204);
or U2352 (N_2352,N_2201,N_2297);
xnor U2353 (N_2353,N_2216,N_2254);
nor U2354 (N_2354,N_2253,N_2246);
and U2355 (N_2355,N_2211,N_2228);
nand U2356 (N_2356,N_2206,N_2262);
or U2357 (N_2357,N_2261,N_2250);
xnor U2358 (N_2358,N_2257,N_2251);
nand U2359 (N_2359,N_2263,N_2222);
or U2360 (N_2360,N_2237,N_2223);
nand U2361 (N_2361,N_2261,N_2219);
xor U2362 (N_2362,N_2241,N_2263);
nor U2363 (N_2363,N_2259,N_2267);
and U2364 (N_2364,N_2253,N_2272);
and U2365 (N_2365,N_2224,N_2264);
and U2366 (N_2366,N_2220,N_2273);
and U2367 (N_2367,N_2285,N_2216);
xor U2368 (N_2368,N_2266,N_2293);
xor U2369 (N_2369,N_2299,N_2244);
nor U2370 (N_2370,N_2227,N_2255);
or U2371 (N_2371,N_2262,N_2292);
and U2372 (N_2372,N_2213,N_2249);
and U2373 (N_2373,N_2216,N_2203);
xor U2374 (N_2374,N_2278,N_2296);
nor U2375 (N_2375,N_2285,N_2273);
and U2376 (N_2376,N_2292,N_2221);
and U2377 (N_2377,N_2258,N_2203);
and U2378 (N_2378,N_2273,N_2206);
and U2379 (N_2379,N_2218,N_2206);
xnor U2380 (N_2380,N_2206,N_2249);
xor U2381 (N_2381,N_2227,N_2295);
or U2382 (N_2382,N_2201,N_2241);
and U2383 (N_2383,N_2283,N_2227);
nand U2384 (N_2384,N_2287,N_2286);
or U2385 (N_2385,N_2299,N_2286);
nand U2386 (N_2386,N_2288,N_2272);
or U2387 (N_2387,N_2215,N_2243);
xnor U2388 (N_2388,N_2245,N_2275);
and U2389 (N_2389,N_2215,N_2258);
nand U2390 (N_2390,N_2265,N_2209);
and U2391 (N_2391,N_2247,N_2243);
or U2392 (N_2392,N_2298,N_2276);
and U2393 (N_2393,N_2269,N_2288);
nor U2394 (N_2394,N_2235,N_2213);
xor U2395 (N_2395,N_2254,N_2211);
nor U2396 (N_2396,N_2270,N_2217);
xor U2397 (N_2397,N_2201,N_2280);
and U2398 (N_2398,N_2213,N_2240);
nand U2399 (N_2399,N_2208,N_2206);
or U2400 (N_2400,N_2388,N_2375);
and U2401 (N_2401,N_2374,N_2372);
or U2402 (N_2402,N_2393,N_2300);
nor U2403 (N_2403,N_2352,N_2395);
nand U2404 (N_2404,N_2362,N_2376);
nand U2405 (N_2405,N_2327,N_2398);
xnor U2406 (N_2406,N_2384,N_2335);
and U2407 (N_2407,N_2339,N_2309);
and U2408 (N_2408,N_2340,N_2351);
and U2409 (N_2409,N_2337,N_2330);
and U2410 (N_2410,N_2353,N_2358);
nand U2411 (N_2411,N_2383,N_2360);
xor U2412 (N_2412,N_2336,N_2302);
nor U2413 (N_2413,N_2348,N_2318);
xnor U2414 (N_2414,N_2370,N_2354);
xnor U2415 (N_2415,N_2361,N_2303);
xor U2416 (N_2416,N_2317,N_2341);
nand U2417 (N_2417,N_2310,N_2347);
or U2418 (N_2418,N_2390,N_2319);
xor U2419 (N_2419,N_2369,N_2389);
nand U2420 (N_2420,N_2396,N_2394);
or U2421 (N_2421,N_2343,N_2326);
xor U2422 (N_2422,N_2315,N_2344);
and U2423 (N_2423,N_2380,N_2377);
or U2424 (N_2424,N_2322,N_2356);
and U2425 (N_2425,N_2329,N_2381);
xor U2426 (N_2426,N_2349,N_2332);
nand U2427 (N_2427,N_2364,N_2368);
or U2428 (N_2428,N_2314,N_2365);
xor U2429 (N_2429,N_2399,N_2387);
or U2430 (N_2430,N_2392,N_2308);
or U2431 (N_2431,N_2366,N_2323);
xor U2432 (N_2432,N_2304,N_2307);
or U2433 (N_2433,N_2378,N_2345);
xor U2434 (N_2434,N_2311,N_2331);
nor U2435 (N_2435,N_2338,N_2324);
and U2436 (N_2436,N_2371,N_2386);
nor U2437 (N_2437,N_2301,N_2346);
and U2438 (N_2438,N_2379,N_2312);
nand U2439 (N_2439,N_2385,N_2359);
or U2440 (N_2440,N_2316,N_2320);
xor U2441 (N_2441,N_2373,N_2328);
nor U2442 (N_2442,N_2363,N_2334);
or U2443 (N_2443,N_2382,N_2325);
and U2444 (N_2444,N_2342,N_2321);
or U2445 (N_2445,N_2355,N_2367);
and U2446 (N_2446,N_2357,N_2391);
and U2447 (N_2447,N_2397,N_2305);
nor U2448 (N_2448,N_2333,N_2350);
nand U2449 (N_2449,N_2306,N_2313);
xor U2450 (N_2450,N_2334,N_2362);
or U2451 (N_2451,N_2333,N_2355);
nor U2452 (N_2452,N_2336,N_2311);
and U2453 (N_2453,N_2341,N_2383);
and U2454 (N_2454,N_2390,N_2326);
and U2455 (N_2455,N_2326,N_2393);
xnor U2456 (N_2456,N_2383,N_2338);
nor U2457 (N_2457,N_2369,N_2319);
or U2458 (N_2458,N_2370,N_2387);
and U2459 (N_2459,N_2357,N_2348);
nand U2460 (N_2460,N_2393,N_2382);
nand U2461 (N_2461,N_2310,N_2319);
or U2462 (N_2462,N_2369,N_2300);
nor U2463 (N_2463,N_2372,N_2341);
nor U2464 (N_2464,N_2326,N_2300);
or U2465 (N_2465,N_2389,N_2352);
or U2466 (N_2466,N_2376,N_2349);
or U2467 (N_2467,N_2397,N_2334);
nor U2468 (N_2468,N_2365,N_2323);
nand U2469 (N_2469,N_2327,N_2358);
xnor U2470 (N_2470,N_2354,N_2314);
xnor U2471 (N_2471,N_2312,N_2390);
or U2472 (N_2472,N_2367,N_2314);
nand U2473 (N_2473,N_2306,N_2395);
nor U2474 (N_2474,N_2387,N_2333);
nand U2475 (N_2475,N_2388,N_2354);
and U2476 (N_2476,N_2321,N_2325);
and U2477 (N_2477,N_2344,N_2383);
xnor U2478 (N_2478,N_2364,N_2385);
and U2479 (N_2479,N_2349,N_2347);
and U2480 (N_2480,N_2365,N_2312);
or U2481 (N_2481,N_2387,N_2345);
nand U2482 (N_2482,N_2397,N_2354);
nand U2483 (N_2483,N_2317,N_2308);
or U2484 (N_2484,N_2387,N_2395);
nor U2485 (N_2485,N_2316,N_2391);
nand U2486 (N_2486,N_2335,N_2391);
or U2487 (N_2487,N_2341,N_2376);
nor U2488 (N_2488,N_2319,N_2328);
and U2489 (N_2489,N_2384,N_2309);
or U2490 (N_2490,N_2367,N_2326);
nand U2491 (N_2491,N_2342,N_2337);
xor U2492 (N_2492,N_2388,N_2330);
xor U2493 (N_2493,N_2364,N_2333);
nor U2494 (N_2494,N_2389,N_2340);
nand U2495 (N_2495,N_2324,N_2391);
and U2496 (N_2496,N_2331,N_2382);
nand U2497 (N_2497,N_2397,N_2308);
nand U2498 (N_2498,N_2355,N_2305);
nand U2499 (N_2499,N_2337,N_2399);
nor U2500 (N_2500,N_2416,N_2430);
and U2501 (N_2501,N_2415,N_2480);
and U2502 (N_2502,N_2411,N_2467);
or U2503 (N_2503,N_2439,N_2454);
nand U2504 (N_2504,N_2479,N_2421);
xnor U2505 (N_2505,N_2493,N_2466);
xor U2506 (N_2506,N_2431,N_2484);
xnor U2507 (N_2507,N_2478,N_2403);
nand U2508 (N_2508,N_2444,N_2455);
xnor U2509 (N_2509,N_2488,N_2458);
and U2510 (N_2510,N_2463,N_2440);
xnor U2511 (N_2511,N_2494,N_2401);
xor U2512 (N_2512,N_2472,N_2498);
nor U2513 (N_2513,N_2400,N_2434);
xnor U2514 (N_2514,N_2420,N_2468);
xnor U2515 (N_2515,N_2437,N_2435);
nand U2516 (N_2516,N_2412,N_2442);
xnor U2517 (N_2517,N_2427,N_2465);
or U2518 (N_2518,N_2404,N_2489);
nand U2519 (N_2519,N_2426,N_2485);
nand U2520 (N_2520,N_2473,N_2441);
nand U2521 (N_2521,N_2410,N_2486);
xor U2522 (N_2522,N_2422,N_2428);
and U2523 (N_2523,N_2496,N_2438);
xnor U2524 (N_2524,N_2490,N_2417);
and U2525 (N_2525,N_2495,N_2456);
nor U2526 (N_2526,N_2406,N_2475);
or U2527 (N_2527,N_2457,N_2470);
and U2528 (N_2528,N_2405,N_2419);
and U2529 (N_2529,N_2446,N_2459);
nor U2530 (N_2530,N_2451,N_2448);
xnor U2531 (N_2531,N_2477,N_2432);
xnor U2532 (N_2532,N_2452,N_2481);
xor U2533 (N_2533,N_2429,N_2424);
xnor U2534 (N_2534,N_2482,N_2425);
xnor U2535 (N_2535,N_2436,N_2474);
xnor U2536 (N_2536,N_2491,N_2464);
nor U2537 (N_2537,N_2450,N_2487);
and U2538 (N_2538,N_2445,N_2499);
and U2539 (N_2539,N_2449,N_2460);
and U2540 (N_2540,N_2483,N_2407);
nor U2541 (N_2541,N_2447,N_2433);
or U2542 (N_2542,N_2418,N_2409);
nand U2543 (N_2543,N_2469,N_2471);
xnor U2544 (N_2544,N_2423,N_2402);
xor U2545 (N_2545,N_2408,N_2453);
xnor U2546 (N_2546,N_2413,N_2414);
nand U2547 (N_2547,N_2461,N_2476);
xor U2548 (N_2548,N_2462,N_2497);
or U2549 (N_2549,N_2443,N_2492);
xnor U2550 (N_2550,N_2453,N_2492);
or U2551 (N_2551,N_2495,N_2499);
and U2552 (N_2552,N_2474,N_2460);
or U2553 (N_2553,N_2487,N_2417);
and U2554 (N_2554,N_2480,N_2473);
or U2555 (N_2555,N_2431,N_2467);
or U2556 (N_2556,N_2401,N_2464);
or U2557 (N_2557,N_2433,N_2440);
nor U2558 (N_2558,N_2417,N_2435);
or U2559 (N_2559,N_2465,N_2443);
or U2560 (N_2560,N_2419,N_2448);
and U2561 (N_2561,N_2470,N_2402);
nor U2562 (N_2562,N_2419,N_2474);
or U2563 (N_2563,N_2480,N_2499);
xor U2564 (N_2564,N_2481,N_2497);
or U2565 (N_2565,N_2439,N_2403);
and U2566 (N_2566,N_2458,N_2472);
and U2567 (N_2567,N_2430,N_2463);
and U2568 (N_2568,N_2482,N_2435);
and U2569 (N_2569,N_2431,N_2495);
or U2570 (N_2570,N_2495,N_2420);
nand U2571 (N_2571,N_2480,N_2417);
and U2572 (N_2572,N_2418,N_2485);
and U2573 (N_2573,N_2469,N_2448);
or U2574 (N_2574,N_2459,N_2429);
nor U2575 (N_2575,N_2453,N_2478);
xor U2576 (N_2576,N_2419,N_2453);
or U2577 (N_2577,N_2425,N_2456);
and U2578 (N_2578,N_2424,N_2454);
xor U2579 (N_2579,N_2425,N_2450);
and U2580 (N_2580,N_2461,N_2436);
or U2581 (N_2581,N_2494,N_2491);
xnor U2582 (N_2582,N_2454,N_2425);
nor U2583 (N_2583,N_2408,N_2467);
nand U2584 (N_2584,N_2459,N_2491);
xor U2585 (N_2585,N_2462,N_2472);
or U2586 (N_2586,N_2418,N_2404);
nor U2587 (N_2587,N_2461,N_2415);
and U2588 (N_2588,N_2471,N_2459);
xnor U2589 (N_2589,N_2437,N_2436);
nor U2590 (N_2590,N_2446,N_2453);
and U2591 (N_2591,N_2495,N_2494);
nand U2592 (N_2592,N_2436,N_2416);
nand U2593 (N_2593,N_2471,N_2466);
or U2594 (N_2594,N_2430,N_2460);
or U2595 (N_2595,N_2425,N_2499);
xor U2596 (N_2596,N_2433,N_2495);
or U2597 (N_2597,N_2464,N_2439);
and U2598 (N_2598,N_2447,N_2457);
and U2599 (N_2599,N_2497,N_2431);
and U2600 (N_2600,N_2575,N_2566);
nor U2601 (N_2601,N_2501,N_2544);
or U2602 (N_2602,N_2525,N_2598);
nand U2603 (N_2603,N_2554,N_2534);
or U2604 (N_2604,N_2578,N_2568);
nand U2605 (N_2605,N_2547,N_2527);
or U2606 (N_2606,N_2530,N_2514);
and U2607 (N_2607,N_2549,N_2545);
nor U2608 (N_2608,N_2588,N_2529);
nand U2609 (N_2609,N_2586,N_2587);
nand U2610 (N_2610,N_2502,N_2582);
xnor U2611 (N_2611,N_2546,N_2551);
and U2612 (N_2612,N_2571,N_2550);
and U2613 (N_2613,N_2507,N_2572);
xor U2614 (N_2614,N_2509,N_2533);
nand U2615 (N_2615,N_2532,N_2556);
or U2616 (N_2616,N_2512,N_2506);
nand U2617 (N_2617,N_2517,N_2513);
nor U2618 (N_2618,N_2538,N_2521);
xnor U2619 (N_2619,N_2516,N_2595);
and U2620 (N_2620,N_2524,N_2540);
xnor U2621 (N_2621,N_2577,N_2536);
nand U2622 (N_2622,N_2593,N_2585);
and U2623 (N_2623,N_2564,N_2569);
nor U2624 (N_2624,N_2579,N_2508);
or U2625 (N_2625,N_2528,N_2570);
nand U2626 (N_2626,N_2592,N_2574);
and U2627 (N_2627,N_2555,N_2596);
nand U2628 (N_2628,N_2580,N_2510);
nand U2629 (N_2629,N_2511,N_2523);
xor U2630 (N_2630,N_2561,N_2504);
nor U2631 (N_2631,N_2597,N_2552);
nor U2632 (N_2632,N_2560,N_2565);
nand U2633 (N_2633,N_2594,N_2557);
or U2634 (N_2634,N_2505,N_2584);
and U2635 (N_2635,N_2518,N_2519);
nand U2636 (N_2636,N_2590,N_2581);
nand U2637 (N_2637,N_2503,N_2522);
and U2638 (N_2638,N_2535,N_2589);
xor U2639 (N_2639,N_2567,N_2553);
and U2640 (N_2640,N_2573,N_2541);
or U2641 (N_2641,N_2542,N_2526);
or U2642 (N_2642,N_2562,N_2599);
nor U2643 (N_2643,N_2559,N_2531);
and U2644 (N_2644,N_2543,N_2520);
or U2645 (N_2645,N_2515,N_2537);
or U2646 (N_2646,N_2548,N_2583);
or U2647 (N_2647,N_2500,N_2558);
and U2648 (N_2648,N_2539,N_2563);
xnor U2649 (N_2649,N_2576,N_2591);
nand U2650 (N_2650,N_2569,N_2538);
xnor U2651 (N_2651,N_2590,N_2510);
xnor U2652 (N_2652,N_2545,N_2502);
xnor U2653 (N_2653,N_2507,N_2561);
nand U2654 (N_2654,N_2512,N_2544);
xnor U2655 (N_2655,N_2510,N_2518);
and U2656 (N_2656,N_2577,N_2570);
and U2657 (N_2657,N_2505,N_2523);
xnor U2658 (N_2658,N_2523,N_2518);
nand U2659 (N_2659,N_2513,N_2551);
xor U2660 (N_2660,N_2574,N_2539);
nand U2661 (N_2661,N_2583,N_2527);
or U2662 (N_2662,N_2560,N_2569);
nor U2663 (N_2663,N_2532,N_2518);
or U2664 (N_2664,N_2544,N_2530);
and U2665 (N_2665,N_2517,N_2594);
nand U2666 (N_2666,N_2578,N_2534);
nor U2667 (N_2667,N_2563,N_2582);
and U2668 (N_2668,N_2545,N_2536);
or U2669 (N_2669,N_2522,N_2557);
xor U2670 (N_2670,N_2560,N_2566);
xor U2671 (N_2671,N_2590,N_2543);
nor U2672 (N_2672,N_2546,N_2539);
xor U2673 (N_2673,N_2570,N_2512);
or U2674 (N_2674,N_2560,N_2567);
nand U2675 (N_2675,N_2565,N_2563);
and U2676 (N_2676,N_2589,N_2531);
or U2677 (N_2677,N_2577,N_2590);
nand U2678 (N_2678,N_2580,N_2500);
or U2679 (N_2679,N_2555,N_2542);
or U2680 (N_2680,N_2520,N_2568);
and U2681 (N_2681,N_2502,N_2520);
nor U2682 (N_2682,N_2520,N_2546);
or U2683 (N_2683,N_2515,N_2518);
xor U2684 (N_2684,N_2594,N_2532);
xor U2685 (N_2685,N_2500,N_2552);
nand U2686 (N_2686,N_2555,N_2524);
nor U2687 (N_2687,N_2502,N_2570);
nor U2688 (N_2688,N_2544,N_2592);
or U2689 (N_2689,N_2544,N_2511);
nor U2690 (N_2690,N_2503,N_2508);
xor U2691 (N_2691,N_2529,N_2559);
xnor U2692 (N_2692,N_2525,N_2546);
nor U2693 (N_2693,N_2587,N_2508);
and U2694 (N_2694,N_2593,N_2584);
nor U2695 (N_2695,N_2547,N_2545);
nand U2696 (N_2696,N_2567,N_2561);
nand U2697 (N_2697,N_2535,N_2548);
or U2698 (N_2698,N_2588,N_2502);
and U2699 (N_2699,N_2504,N_2599);
and U2700 (N_2700,N_2647,N_2659);
or U2701 (N_2701,N_2658,N_2618);
nor U2702 (N_2702,N_2606,N_2675);
nor U2703 (N_2703,N_2676,N_2692);
xor U2704 (N_2704,N_2607,N_2663);
nor U2705 (N_2705,N_2627,N_2610);
nor U2706 (N_2706,N_2615,N_2665);
or U2707 (N_2707,N_2608,N_2678);
nand U2708 (N_2708,N_2666,N_2650);
and U2709 (N_2709,N_2686,N_2633);
or U2710 (N_2710,N_2611,N_2698);
and U2711 (N_2711,N_2694,N_2643);
or U2712 (N_2712,N_2653,N_2677);
xnor U2713 (N_2713,N_2684,N_2644);
or U2714 (N_2714,N_2648,N_2626);
and U2715 (N_2715,N_2681,N_2697);
or U2716 (N_2716,N_2661,N_2628);
and U2717 (N_2717,N_2652,N_2619);
xor U2718 (N_2718,N_2693,N_2673);
xor U2719 (N_2719,N_2635,N_2632);
nand U2720 (N_2720,N_2646,N_2613);
nand U2721 (N_2721,N_2639,N_2683);
nand U2722 (N_2722,N_2642,N_2671);
nand U2723 (N_2723,N_2654,N_2656);
xnor U2724 (N_2724,N_2690,N_2664);
or U2725 (N_2725,N_2699,N_2601);
nor U2726 (N_2726,N_2651,N_2670);
nor U2727 (N_2727,N_2623,N_2616);
or U2728 (N_2728,N_2668,N_2630);
nor U2729 (N_2729,N_2624,N_2617);
and U2730 (N_2730,N_2691,N_2669);
nor U2731 (N_2731,N_2680,N_2645);
nand U2732 (N_2732,N_2672,N_2604);
nor U2733 (N_2733,N_2625,N_2603);
xnor U2734 (N_2734,N_2696,N_2688);
and U2735 (N_2735,N_2682,N_2689);
and U2736 (N_2736,N_2621,N_2657);
nor U2737 (N_2737,N_2614,N_2600);
nand U2738 (N_2738,N_2602,N_2660);
nand U2739 (N_2739,N_2629,N_2662);
or U2740 (N_2740,N_2695,N_2679);
and U2741 (N_2741,N_2612,N_2620);
xnor U2742 (N_2742,N_2655,N_2641);
nand U2743 (N_2743,N_2622,N_2609);
and U2744 (N_2744,N_2636,N_2685);
nor U2745 (N_2745,N_2631,N_2640);
nand U2746 (N_2746,N_2649,N_2667);
xnor U2747 (N_2747,N_2605,N_2687);
nand U2748 (N_2748,N_2634,N_2637);
nand U2749 (N_2749,N_2674,N_2638);
or U2750 (N_2750,N_2678,N_2674);
nor U2751 (N_2751,N_2626,N_2611);
and U2752 (N_2752,N_2679,N_2634);
and U2753 (N_2753,N_2699,N_2654);
or U2754 (N_2754,N_2640,N_2663);
xor U2755 (N_2755,N_2662,N_2674);
nor U2756 (N_2756,N_2649,N_2661);
or U2757 (N_2757,N_2699,N_2637);
nor U2758 (N_2758,N_2688,N_2602);
nor U2759 (N_2759,N_2600,N_2699);
and U2760 (N_2760,N_2660,N_2616);
xor U2761 (N_2761,N_2693,N_2609);
or U2762 (N_2762,N_2642,N_2699);
and U2763 (N_2763,N_2635,N_2640);
nand U2764 (N_2764,N_2625,N_2693);
or U2765 (N_2765,N_2661,N_2637);
and U2766 (N_2766,N_2652,N_2663);
xnor U2767 (N_2767,N_2659,N_2698);
nand U2768 (N_2768,N_2671,N_2650);
nand U2769 (N_2769,N_2651,N_2681);
nand U2770 (N_2770,N_2629,N_2650);
and U2771 (N_2771,N_2681,N_2603);
and U2772 (N_2772,N_2660,N_2656);
or U2773 (N_2773,N_2646,N_2683);
nand U2774 (N_2774,N_2665,N_2623);
or U2775 (N_2775,N_2614,N_2685);
or U2776 (N_2776,N_2602,N_2635);
or U2777 (N_2777,N_2641,N_2622);
or U2778 (N_2778,N_2607,N_2637);
or U2779 (N_2779,N_2645,N_2610);
and U2780 (N_2780,N_2685,N_2604);
xor U2781 (N_2781,N_2655,N_2616);
or U2782 (N_2782,N_2637,N_2665);
or U2783 (N_2783,N_2685,N_2690);
nor U2784 (N_2784,N_2618,N_2695);
and U2785 (N_2785,N_2610,N_2641);
nor U2786 (N_2786,N_2602,N_2613);
or U2787 (N_2787,N_2694,N_2693);
xor U2788 (N_2788,N_2629,N_2675);
nor U2789 (N_2789,N_2646,N_2602);
nor U2790 (N_2790,N_2694,N_2648);
nor U2791 (N_2791,N_2616,N_2601);
xnor U2792 (N_2792,N_2611,N_2639);
xor U2793 (N_2793,N_2682,N_2658);
nand U2794 (N_2794,N_2648,N_2686);
nor U2795 (N_2795,N_2639,N_2672);
nand U2796 (N_2796,N_2669,N_2614);
nand U2797 (N_2797,N_2653,N_2642);
and U2798 (N_2798,N_2626,N_2645);
or U2799 (N_2799,N_2669,N_2615);
xor U2800 (N_2800,N_2721,N_2793);
and U2801 (N_2801,N_2720,N_2754);
nor U2802 (N_2802,N_2784,N_2757);
xnor U2803 (N_2803,N_2769,N_2733);
or U2804 (N_2804,N_2728,N_2729);
nand U2805 (N_2805,N_2744,N_2761);
nand U2806 (N_2806,N_2701,N_2752);
or U2807 (N_2807,N_2775,N_2700);
xor U2808 (N_2808,N_2758,N_2713);
or U2809 (N_2809,N_2703,N_2773);
or U2810 (N_2810,N_2786,N_2798);
xnor U2811 (N_2811,N_2704,N_2759);
xor U2812 (N_2812,N_2779,N_2756);
xnor U2813 (N_2813,N_2727,N_2723);
nor U2814 (N_2814,N_2764,N_2787);
nand U2815 (N_2815,N_2783,N_2770);
or U2816 (N_2816,N_2738,N_2748);
and U2817 (N_2817,N_2755,N_2780);
nand U2818 (N_2818,N_2711,N_2795);
and U2819 (N_2819,N_2739,N_2785);
xor U2820 (N_2820,N_2753,N_2705);
or U2821 (N_2821,N_2725,N_2708);
or U2822 (N_2822,N_2726,N_2763);
xor U2823 (N_2823,N_2766,N_2776);
and U2824 (N_2824,N_2782,N_2707);
nand U2825 (N_2825,N_2745,N_2797);
or U2826 (N_2826,N_2771,N_2778);
nor U2827 (N_2827,N_2750,N_2706);
or U2828 (N_2828,N_2772,N_2790);
or U2829 (N_2829,N_2715,N_2719);
or U2830 (N_2830,N_2762,N_2735);
nor U2831 (N_2831,N_2718,N_2792);
xnor U2832 (N_2832,N_2747,N_2774);
nand U2833 (N_2833,N_2736,N_2768);
and U2834 (N_2834,N_2760,N_2741);
or U2835 (N_2835,N_2749,N_2781);
nor U2836 (N_2836,N_2724,N_2777);
xor U2837 (N_2837,N_2743,N_2722);
nand U2838 (N_2838,N_2737,N_2796);
nand U2839 (N_2839,N_2788,N_2767);
nor U2840 (N_2840,N_2751,N_2765);
and U2841 (N_2841,N_2730,N_2732);
and U2842 (N_2842,N_2712,N_2746);
or U2843 (N_2843,N_2716,N_2709);
and U2844 (N_2844,N_2794,N_2731);
xor U2845 (N_2845,N_2799,N_2791);
or U2846 (N_2846,N_2702,N_2789);
or U2847 (N_2847,N_2734,N_2710);
and U2848 (N_2848,N_2742,N_2717);
or U2849 (N_2849,N_2740,N_2714);
nor U2850 (N_2850,N_2753,N_2770);
xor U2851 (N_2851,N_2719,N_2740);
or U2852 (N_2852,N_2720,N_2711);
xnor U2853 (N_2853,N_2726,N_2733);
or U2854 (N_2854,N_2746,N_2725);
or U2855 (N_2855,N_2750,N_2702);
nor U2856 (N_2856,N_2768,N_2742);
nor U2857 (N_2857,N_2706,N_2775);
nor U2858 (N_2858,N_2721,N_2706);
nor U2859 (N_2859,N_2753,N_2771);
xnor U2860 (N_2860,N_2795,N_2757);
xnor U2861 (N_2861,N_2715,N_2731);
and U2862 (N_2862,N_2735,N_2715);
xor U2863 (N_2863,N_2755,N_2796);
nand U2864 (N_2864,N_2774,N_2789);
and U2865 (N_2865,N_2757,N_2748);
and U2866 (N_2866,N_2797,N_2734);
nor U2867 (N_2867,N_2717,N_2785);
nor U2868 (N_2868,N_2761,N_2783);
xor U2869 (N_2869,N_2707,N_2752);
nand U2870 (N_2870,N_2708,N_2789);
and U2871 (N_2871,N_2729,N_2793);
nand U2872 (N_2872,N_2765,N_2757);
and U2873 (N_2873,N_2777,N_2720);
nor U2874 (N_2874,N_2763,N_2737);
nand U2875 (N_2875,N_2771,N_2767);
nor U2876 (N_2876,N_2747,N_2788);
xnor U2877 (N_2877,N_2715,N_2754);
nand U2878 (N_2878,N_2771,N_2715);
or U2879 (N_2879,N_2764,N_2775);
nor U2880 (N_2880,N_2758,N_2749);
xor U2881 (N_2881,N_2710,N_2753);
or U2882 (N_2882,N_2735,N_2727);
or U2883 (N_2883,N_2748,N_2742);
nor U2884 (N_2884,N_2732,N_2714);
and U2885 (N_2885,N_2765,N_2789);
xnor U2886 (N_2886,N_2758,N_2764);
and U2887 (N_2887,N_2730,N_2741);
or U2888 (N_2888,N_2792,N_2796);
nand U2889 (N_2889,N_2717,N_2799);
nand U2890 (N_2890,N_2741,N_2725);
nand U2891 (N_2891,N_2738,N_2776);
or U2892 (N_2892,N_2745,N_2732);
nand U2893 (N_2893,N_2753,N_2755);
nand U2894 (N_2894,N_2757,N_2727);
nor U2895 (N_2895,N_2785,N_2767);
xor U2896 (N_2896,N_2741,N_2790);
xor U2897 (N_2897,N_2769,N_2703);
nor U2898 (N_2898,N_2783,N_2710);
xor U2899 (N_2899,N_2768,N_2741);
and U2900 (N_2900,N_2801,N_2861);
and U2901 (N_2901,N_2880,N_2843);
nor U2902 (N_2902,N_2828,N_2808);
nor U2903 (N_2903,N_2856,N_2862);
and U2904 (N_2904,N_2807,N_2896);
nor U2905 (N_2905,N_2872,N_2827);
nand U2906 (N_2906,N_2826,N_2893);
xor U2907 (N_2907,N_2811,N_2819);
or U2908 (N_2908,N_2838,N_2863);
nor U2909 (N_2909,N_2854,N_2844);
nand U2910 (N_2910,N_2886,N_2852);
and U2911 (N_2911,N_2858,N_2846);
and U2912 (N_2912,N_2832,N_2816);
nor U2913 (N_2913,N_2885,N_2806);
nor U2914 (N_2914,N_2897,N_2820);
or U2915 (N_2915,N_2878,N_2853);
or U2916 (N_2916,N_2870,N_2867);
or U2917 (N_2917,N_2873,N_2814);
nor U2918 (N_2918,N_2898,N_2892);
nand U2919 (N_2919,N_2857,N_2849);
nor U2920 (N_2920,N_2802,N_2882);
xnor U2921 (N_2921,N_2850,N_2881);
xnor U2922 (N_2922,N_2818,N_2891);
and U2923 (N_2923,N_2804,N_2879);
nor U2924 (N_2924,N_2836,N_2884);
or U2925 (N_2925,N_2855,N_2869);
and U2926 (N_2926,N_2829,N_2876);
and U2927 (N_2927,N_2847,N_2851);
or U2928 (N_2928,N_2888,N_2813);
nor U2929 (N_2929,N_2871,N_2866);
xnor U2930 (N_2930,N_2824,N_2810);
nor U2931 (N_2931,N_2859,N_2834);
and U2932 (N_2932,N_2815,N_2874);
xnor U2933 (N_2933,N_2817,N_2833);
nor U2934 (N_2934,N_2845,N_2860);
or U2935 (N_2935,N_2887,N_2894);
or U2936 (N_2936,N_2864,N_2875);
and U2937 (N_2937,N_2848,N_2877);
or U2938 (N_2938,N_2865,N_2899);
nor U2939 (N_2939,N_2895,N_2839);
nand U2940 (N_2940,N_2868,N_2841);
nor U2941 (N_2941,N_2800,N_2821);
xnor U2942 (N_2942,N_2835,N_2822);
and U2943 (N_2943,N_2812,N_2837);
xnor U2944 (N_2944,N_2889,N_2803);
nor U2945 (N_2945,N_2809,N_2840);
or U2946 (N_2946,N_2883,N_2823);
nand U2947 (N_2947,N_2825,N_2831);
nand U2948 (N_2948,N_2890,N_2830);
xnor U2949 (N_2949,N_2805,N_2842);
nand U2950 (N_2950,N_2850,N_2846);
xor U2951 (N_2951,N_2828,N_2871);
and U2952 (N_2952,N_2881,N_2849);
nand U2953 (N_2953,N_2885,N_2879);
or U2954 (N_2954,N_2874,N_2821);
or U2955 (N_2955,N_2828,N_2825);
and U2956 (N_2956,N_2876,N_2852);
or U2957 (N_2957,N_2843,N_2801);
and U2958 (N_2958,N_2808,N_2848);
and U2959 (N_2959,N_2892,N_2879);
nor U2960 (N_2960,N_2846,N_2863);
and U2961 (N_2961,N_2846,N_2880);
and U2962 (N_2962,N_2883,N_2898);
xor U2963 (N_2963,N_2834,N_2838);
and U2964 (N_2964,N_2810,N_2857);
nand U2965 (N_2965,N_2881,N_2835);
and U2966 (N_2966,N_2849,N_2842);
and U2967 (N_2967,N_2841,N_2895);
xnor U2968 (N_2968,N_2819,N_2803);
and U2969 (N_2969,N_2849,N_2854);
or U2970 (N_2970,N_2810,N_2819);
or U2971 (N_2971,N_2890,N_2873);
nand U2972 (N_2972,N_2879,N_2899);
nor U2973 (N_2973,N_2811,N_2849);
and U2974 (N_2974,N_2833,N_2898);
nand U2975 (N_2975,N_2808,N_2898);
nand U2976 (N_2976,N_2895,N_2866);
xor U2977 (N_2977,N_2857,N_2879);
xnor U2978 (N_2978,N_2855,N_2817);
xor U2979 (N_2979,N_2836,N_2808);
xor U2980 (N_2980,N_2823,N_2841);
xor U2981 (N_2981,N_2809,N_2854);
xor U2982 (N_2982,N_2889,N_2859);
xor U2983 (N_2983,N_2892,N_2834);
xnor U2984 (N_2984,N_2882,N_2825);
nor U2985 (N_2985,N_2859,N_2830);
nor U2986 (N_2986,N_2857,N_2830);
xnor U2987 (N_2987,N_2880,N_2800);
and U2988 (N_2988,N_2830,N_2838);
or U2989 (N_2989,N_2810,N_2811);
or U2990 (N_2990,N_2830,N_2860);
xnor U2991 (N_2991,N_2814,N_2864);
or U2992 (N_2992,N_2853,N_2801);
xor U2993 (N_2993,N_2876,N_2838);
nor U2994 (N_2994,N_2869,N_2818);
and U2995 (N_2995,N_2839,N_2814);
or U2996 (N_2996,N_2839,N_2835);
nand U2997 (N_2997,N_2845,N_2848);
nand U2998 (N_2998,N_2894,N_2881);
nand U2999 (N_2999,N_2831,N_2842);
nor U3000 (N_3000,N_2963,N_2905);
nor U3001 (N_3001,N_2922,N_2950);
and U3002 (N_3002,N_2976,N_2901);
nand U3003 (N_3003,N_2986,N_2921);
nor U3004 (N_3004,N_2933,N_2907);
nand U3005 (N_3005,N_2982,N_2940);
xnor U3006 (N_3006,N_2975,N_2910);
xor U3007 (N_3007,N_2946,N_2974);
nand U3008 (N_3008,N_2959,N_2951);
xnor U3009 (N_3009,N_2965,N_2929);
or U3010 (N_3010,N_2914,N_2989);
or U3011 (N_3011,N_2988,N_2912);
and U3012 (N_3012,N_2985,N_2941);
or U3013 (N_3013,N_2939,N_2916);
or U3014 (N_3014,N_2926,N_2978);
nor U3015 (N_3015,N_2971,N_2972);
nor U3016 (N_3016,N_2983,N_2958);
nor U3017 (N_3017,N_2932,N_2995);
xor U3018 (N_3018,N_2994,N_2952);
nor U3019 (N_3019,N_2984,N_2920);
nand U3020 (N_3020,N_2973,N_2993);
or U3021 (N_3021,N_2966,N_2934);
xor U3022 (N_3022,N_2999,N_2998);
and U3023 (N_3023,N_2962,N_2935);
xor U3024 (N_3024,N_2991,N_2903);
nor U3025 (N_3025,N_2915,N_2992);
and U3026 (N_3026,N_2913,N_2964);
and U3027 (N_3027,N_2980,N_2954);
nor U3028 (N_3028,N_2931,N_2956);
or U3029 (N_3029,N_2981,N_2908);
nor U3030 (N_3030,N_2996,N_2948);
nor U3031 (N_3031,N_2967,N_2970);
nor U3032 (N_3032,N_2987,N_2927);
and U3033 (N_3033,N_2953,N_2911);
nand U3034 (N_3034,N_2955,N_2969);
nor U3035 (N_3035,N_2947,N_2904);
or U3036 (N_3036,N_2990,N_2949);
or U3037 (N_3037,N_2968,N_2937);
or U3038 (N_3038,N_2960,N_2943);
and U3039 (N_3039,N_2900,N_2925);
and U3040 (N_3040,N_2957,N_2906);
nor U3041 (N_3041,N_2917,N_2942);
or U3042 (N_3042,N_2909,N_2930);
nand U3043 (N_3043,N_2928,N_2944);
xnor U3044 (N_3044,N_2945,N_2961);
nor U3045 (N_3045,N_2938,N_2997);
and U3046 (N_3046,N_2923,N_2979);
and U3047 (N_3047,N_2902,N_2924);
nand U3048 (N_3048,N_2936,N_2977);
nand U3049 (N_3049,N_2918,N_2919);
xor U3050 (N_3050,N_2985,N_2936);
or U3051 (N_3051,N_2971,N_2908);
nor U3052 (N_3052,N_2956,N_2966);
nor U3053 (N_3053,N_2973,N_2990);
xor U3054 (N_3054,N_2944,N_2992);
nand U3055 (N_3055,N_2903,N_2972);
or U3056 (N_3056,N_2965,N_2940);
nor U3057 (N_3057,N_2917,N_2941);
or U3058 (N_3058,N_2962,N_2932);
nand U3059 (N_3059,N_2972,N_2958);
xor U3060 (N_3060,N_2975,N_2940);
nand U3061 (N_3061,N_2964,N_2931);
nand U3062 (N_3062,N_2933,N_2965);
or U3063 (N_3063,N_2973,N_2951);
and U3064 (N_3064,N_2953,N_2957);
nand U3065 (N_3065,N_2998,N_2969);
nand U3066 (N_3066,N_2970,N_2990);
or U3067 (N_3067,N_2973,N_2987);
or U3068 (N_3068,N_2937,N_2957);
and U3069 (N_3069,N_2949,N_2961);
and U3070 (N_3070,N_2923,N_2929);
nor U3071 (N_3071,N_2998,N_2982);
nand U3072 (N_3072,N_2941,N_2907);
xor U3073 (N_3073,N_2963,N_2928);
or U3074 (N_3074,N_2901,N_2944);
or U3075 (N_3075,N_2948,N_2949);
or U3076 (N_3076,N_2912,N_2934);
and U3077 (N_3077,N_2966,N_2965);
nand U3078 (N_3078,N_2944,N_2971);
or U3079 (N_3079,N_2978,N_2986);
nor U3080 (N_3080,N_2942,N_2980);
nor U3081 (N_3081,N_2979,N_2960);
or U3082 (N_3082,N_2940,N_2989);
nand U3083 (N_3083,N_2989,N_2916);
xnor U3084 (N_3084,N_2969,N_2959);
or U3085 (N_3085,N_2948,N_2955);
nor U3086 (N_3086,N_2977,N_2999);
nand U3087 (N_3087,N_2923,N_2994);
nand U3088 (N_3088,N_2965,N_2962);
and U3089 (N_3089,N_2929,N_2985);
or U3090 (N_3090,N_2909,N_2979);
or U3091 (N_3091,N_2935,N_2993);
xnor U3092 (N_3092,N_2943,N_2955);
xor U3093 (N_3093,N_2909,N_2980);
nand U3094 (N_3094,N_2964,N_2949);
and U3095 (N_3095,N_2940,N_2984);
and U3096 (N_3096,N_2933,N_2914);
nor U3097 (N_3097,N_2950,N_2944);
or U3098 (N_3098,N_2912,N_2915);
xor U3099 (N_3099,N_2951,N_2950);
nor U3100 (N_3100,N_3026,N_3002);
and U3101 (N_3101,N_3043,N_3088);
or U3102 (N_3102,N_3045,N_3031);
xnor U3103 (N_3103,N_3078,N_3052);
xnor U3104 (N_3104,N_3018,N_3064);
xnor U3105 (N_3105,N_3068,N_3080);
and U3106 (N_3106,N_3087,N_3099);
nand U3107 (N_3107,N_3057,N_3077);
and U3108 (N_3108,N_3038,N_3054);
and U3109 (N_3109,N_3016,N_3062);
xor U3110 (N_3110,N_3059,N_3034);
or U3111 (N_3111,N_3001,N_3019);
nand U3112 (N_3112,N_3037,N_3071);
nand U3113 (N_3113,N_3056,N_3061);
nor U3114 (N_3114,N_3007,N_3044);
nand U3115 (N_3115,N_3082,N_3063);
xor U3116 (N_3116,N_3015,N_3060);
nor U3117 (N_3117,N_3072,N_3055);
nand U3118 (N_3118,N_3020,N_3004);
or U3119 (N_3119,N_3024,N_3095);
and U3120 (N_3120,N_3008,N_3074);
xnor U3121 (N_3121,N_3076,N_3075);
xnor U3122 (N_3122,N_3029,N_3050);
or U3123 (N_3123,N_3046,N_3097);
nand U3124 (N_3124,N_3048,N_3047);
and U3125 (N_3125,N_3017,N_3005);
xnor U3126 (N_3126,N_3092,N_3032);
nand U3127 (N_3127,N_3022,N_3023);
or U3128 (N_3128,N_3042,N_3083);
nand U3129 (N_3129,N_3028,N_3051);
nand U3130 (N_3130,N_3039,N_3014);
and U3131 (N_3131,N_3027,N_3011);
nor U3132 (N_3132,N_3073,N_3091);
nor U3133 (N_3133,N_3067,N_3070);
or U3134 (N_3134,N_3041,N_3090);
nand U3135 (N_3135,N_3086,N_3006);
xnor U3136 (N_3136,N_3000,N_3033);
nor U3137 (N_3137,N_3065,N_3013);
or U3138 (N_3138,N_3085,N_3053);
xor U3139 (N_3139,N_3040,N_3058);
and U3140 (N_3140,N_3035,N_3093);
nor U3141 (N_3141,N_3021,N_3030);
nor U3142 (N_3142,N_3069,N_3003);
or U3143 (N_3143,N_3049,N_3084);
nand U3144 (N_3144,N_3066,N_3098);
nor U3145 (N_3145,N_3025,N_3089);
or U3146 (N_3146,N_3010,N_3081);
nand U3147 (N_3147,N_3096,N_3036);
and U3148 (N_3148,N_3012,N_3079);
or U3149 (N_3149,N_3094,N_3009);
or U3150 (N_3150,N_3091,N_3081);
or U3151 (N_3151,N_3001,N_3092);
nand U3152 (N_3152,N_3066,N_3086);
and U3153 (N_3153,N_3091,N_3007);
xnor U3154 (N_3154,N_3050,N_3075);
and U3155 (N_3155,N_3029,N_3000);
nor U3156 (N_3156,N_3044,N_3098);
and U3157 (N_3157,N_3025,N_3073);
nand U3158 (N_3158,N_3044,N_3096);
and U3159 (N_3159,N_3051,N_3032);
or U3160 (N_3160,N_3014,N_3085);
nor U3161 (N_3161,N_3020,N_3038);
xor U3162 (N_3162,N_3022,N_3010);
nor U3163 (N_3163,N_3045,N_3076);
xnor U3164 (N_3164,N_3001,N_3077);
nand U3165 (N_3165,N_3042,N_3008);
nor U3166 (N_3166,N_3000,N_3085);
xnor U3167 (N_3167,N_3069,N_3068);
xor U3168 (N_3168,N_3076,N_3091);
nor U3169 (N_3169,N_3086,N_3056);
or U3170 (N_3170,N_3056,N_3032);
nor U3171 (N_3171,N_3007,N_3024);
nor U3172 (N_3172,N_3003,N_3042);
or U3173 (N_3173,N_3052,N_3041);
nor U3174 (N_3174,N_3079,N_3009);
xor U3175 (N_3175,N_3005,N_3022);
xor U3176 (N_3176,N_3000,N_3050);
nor U3177 (N_3177,N_3035,N_3059);
xnor U3178 (N_3178,N_3086,N_3083);
nand U3179 (N_3179,N_3087,N_3040);
nand U3180 (N_3180,N_3088,N_3069);
xnor U3181 (N_3181,N_3042,N_3013);
or U3182 (N_3182,N_3022,N_3099);
nand U3183 (N_3183,N_3015,N_3041);
xor U3184 (N_3184,N_3054,N_3066);
or U3185 (N_3185,N_3055,N_3070);
and U3186 (N_3186,N_3067,N_3000);
xnor U3187 (N_3187,N_3086,N_3005);
nor U3188 (N_3188,N_3099,N_3098);
xnor U3189 (N_3189,N_3047,N_3083);
and U3190 (N_3190,N_3049,N_3036);
or U3191 (N_3191,N_3081,N_3012);
nor U3192 (N_3192,N_3045,N_3063);
xor U3193 (N_3193,N_3042,N_3066);
nor U3194 (N_3194,N_3005,N_3048);
nor U3195 (N_3195,N_3066,N_3093);
nand U3196 (N_3196,N_3073,N_3057);
nand U3197 (N_3197,N_3068,N_3025);
and U3198 (N_3198,N_3015,N_3098);
xor U3199 (N_3199,N_3082,N_3060);
or U3200 (N_3200,N_3198,N_3144);
nor U3201 (N_3201,N_3197,N_3164);
nand U3202 (N_3202,N_3128,N_3140);
or U3203 (N_3203,N_3168,N_3113);
nand U3204 (N_3204,N_3105,N_3123);
nand U3205 (N_3205,N_3184,N_3112);
nor U3206 (N_3206,N_3139,N_3151);
nor U3207 (N_3207,N_3114,N_3191);
and U3208 (N_3208,N_3138,N_3143);
xnor U3209 (N_3209,N_3166,N_3133);
xnor U3210 (N_3210,N_3187,N_3160);
or U3211 (N_3211,N_3122,N_3111);
and U3212 (N_3212,N_3141,N_3131);
and U3213 (N_3213,N_3174,N_3107);
and U3214 (N_3214,N_3193,N_3189);
and U3215 (N_3215,N_3118,N_3155);
nor U3216 (N_3216,N_3161,N_3181);
nor U3217 (N_3217,N_3115,N_3154);
xnor U3218 (N_3218,N_3108,N_3132);
or U3219 (N_3219,N_3183,N_3101);
or U3220 (N_3220,N_3180,N_3150);
and U3221 (N_3221,N_3188,N_3173);
xnor U3222 (N_3222,N_3170,N_3106);
or U3223 (N_3223,N_3117,N_3102);
nand U3224 (N_3224,N_3165,N_3190);
and U3225 (N_3225,N_3120,N_3135);
nand U3226 (N_3226,N_3142,N_3152);
or U3227 (N_3227,N_3195,N_3137);
nor U3228 (N_3228,N_3179,N_3196);
or U3229 (N_3229,N_3163,N_3126);
nand U3230 (N_3230,N_3153,N_3124);
or U3231 (N_3231,N_3127,N_3159);
nand U3232 (N_3232,N_3110,N_3199);
nor U3233 (N_3233,N_3129,N_3116);
xor U3234 (N_3234,N_3146,N_3192);
nand U3235 (N_3235,N_3177,N_3121);
nor U3236 (N_3236,N_3109,N_3104);
nand U3237 (N_3237,N_3172,N_3194);
xor U3238 (N_3238,N_3176,N_3182);
nor U3239 (N_3239,N_3103,N_3156);
nand U3240 (N_3240,N_3167,N_3125);
and U3241 (N_3241,N_3147,N_3134);
nand U3242 (N_3242,N_3145,N_3178);
xnor U3243 (N_3243,N_3186,N_3130);
nand U3244 (N_3244,N_3175,N_3100);
nand U3245 (N_3245,N_3136,N_3149);
and U3246 (N_3246,N_3148,N_3171);
xor U3247 (N_3247,N_3185,N_3119);
xnor U3248 (N_3248,N_3162,N_3169);
nand U3249 (N_3249,N_3157,N_3158);
and U3250 (N_3250,N_3103,N_3172);
xor U3251 (N_3251,N_3109,N_3185);
nor U3252 (N_3252,N_3166,N_3198);
or U3253 (N_3253,N_3122,N_3127);
nand U3254 (N_3254,N_3198,N_3146);
xnor U3255 (N_3255,N_3175,N_3147);
nor U3256 (N_3256,N_3191,N_3178);
xor U3257 (N_3257,N_3125,N_3188);
xnor U3258 (N_3258,N_3100,N_3158);
or U3259 (N_3259,N_3116,N_3103);
and U3260 (N_3260,N_3142,N_3165);
xor U3261 (N_3261,N_3191,N_3125);
xnor U3262 (N_3262,N_3159,N_3107);
or U3263 (N_3263,N_3156,N_3173);
xnor U3264 (N_3264,N_3188,N_3144);
and U3265 (N_3265,N_3139,N_3172);
nand U3266 (N_3266,N_3198,N_3173);
nand U3267 (N_3267,N_3104,N_3143);
nor U3268 (N_3268,N_3139,N_3121);
nor U3269 (N_3269,N_3189,N_3187);
or U3270 (N_3270,N_3179,N_3160);
nand U3271 (N_3271,N_3190,N_3103);
nor U3272 (N_3272,N_3140,N_3129);
nor U3273 (N_3273,N_3196,N_3151);
or U3274 (N_3274,N_3176,N_3123);
or U3275 (N_3275,N_3129,N_3191);
xnor U3276 (N_3276,N_3160,N_3147);
or U3277 (N_3277,N_3193,N_3192);
and U3278 (N_3278,N_3153,N_3198);
nand U3279 (N_3279,N_3112,N_3146);
nor U3280 (N_3280,N_3157,N_3111);
xor U3281 (N_3281,N_3194,N_3113);
nor U3282 (N_3282,N_3170,N_3157);
nand U3283 (N_3283,N_3121,N_3165);
nor U3284 (N_3284,N_3119,N_3127);
nand U3285 (N_3285,N_3140,N_3160);
nand U3286 (N_3286,N_3183,N_3182);
xnor U3287 (N_3287,N_3186,N_3176);
xnor U3288 (N_3288,N_3136,N_3193);
xor U3289 (N_3289,N_3142,N_3156);
xnor U3290 (N_3290,N_3185,N_3164);
or U3291 (N_3291,N_3145,N_3189);
xor U3292 (N_3292,N_3135,N_3149);
or U3293 (N_3293,N_3160,N_3162);
or U3294 (N_3294,N_3138,N_3165);
and U3295 (N_3295,N_3174,N_3188);
xnor U3296 (N_3296,N_3137,N_3162);
nor U3297 (N_3297,N_3183,N_3160);
nand U3298 (N_3298,N_3113,N_3150);
nor U3299 (N_3299,N_3123,N_3163);
nand U3300 (N_3300,N_3266,N_3238);
nand U3301 (N_3301,N_3227,N_3233);
nor U3302 (N_3302,N_3251,N_3255);
nand U3303 (N_3303,N_3219,N_3229);
and U3304 (N_3304,N_3221,N_3286);
and U3305 (N_3305,N_3291,N_3216);
or U3306 (N_3306,N_3282,N_3294);
or U3307 (N_3307,N_3268,N_3273);
and U3308 (N_3308,N_3265,N_3240);
nand U3309 (N_3309,N_3247,N_3204);
or U3310 (N_3310,N_3217,N_3208);
or U3311 (N_3311,N_3234,N_3235);
and U3312 (N_3312,N_3253,N_3296);
xnor U3313 (N_3313,N_3281,N_3298);
and U3314 (N_3314,N_3210,N_3241);
or U3315 (N_3315,N_3299,N_3249);
nor U3316 (N_3316,N_3228,N_3239);
or U3317 (N_3317,N_3260,N_3209);
or U3318 (N_3318,N_3205,N_3248);
nand U3319 (N_3319,N_3293,N_3201);
or U3320 (N_3320,N_3250,N_3297);
nor U3321 (N_3321,N_3200,N_3223);
and U3322 (N_3322,N_3222,N_3256);
or U3323 (N_3323,N_3245,N_3252);
and U3324 (N_3324,N_3206,N_3231);
and U3325 (N_3325,N_3292,N_3254);
xnor U3326 (N_3326,N_3230,N_3279);
xor U3327 (N_3327,N_3276,N_3271);
xnor U3328 (N_3328,N_3280,N_3288);
xnor U3329 (N_3329,N_3202,N_3224);
or U3330 (N_3330,N_3243,N_3218);
nand U3331 (N_3331,N_3214,N_3272);
or U3332 (N_3332,N_3270,N_3285);
nand U3333 (N_3333,N_3278,N_3295);
or U3334 (N_3334,N_3236,N_3203);
and U3335 (N_3335,N_3242,N_3225);
xnor U3336 (N_3336,N_3283,N_3259);
xnor U3337 (N_3337,N_3261,N_3262);
xnor U3338 (N_3338,N_3290,N_3287);
or U3339 (N_3339,N_3207,N_3246);
and U3340 (N_3340,N_3232,N_3263);
nand U3341 (N_3341,N_3258,N_3244);
or U3342 (N_3342,N_3257,N_3267);
and U3343 (N_3343,N_3213,N_3211);
nand U3344 (N_3344,N_3284,N_3212);
nand U3345 (N_3345,N_3275,N_3264);
nand U3346 (N_3346,N_3277,N_3274);
or U3347 (N_3347,N_3215,N_3237);
and U3348 (N_3348,N_3220,N_3269);
or U3349 (N_3349,N_3226,N_3289);
nand U3350 (N_3350,N_3293,N_3269);
nor U3351 (N_3351,N_3225,N_3244);
or U3352 (N_3352,N_3256,N_3234);
xnor U3353 (N_3353,N_3248,N_3225);
or U3354 (N_3354,N_3209,N_3250);
nand U3355 (N_3355,N_3215,N_3265);
nor U3356 (N_3356,N_3269,N_3248);
and U3357 (N_3357,N_3273,N_3236);
xor U3358 (N_3358,N_3241,N_3277);
nor U3359 (N_3359,N_3259,N_3211);
xnor U3360 (N_3360,N_3246,N_3260);
xor U3361 (N_3361,N_3219,N_3242);
xnor U3362 (N_3362,N_3249,N_3245);
xnor U3363 (N_3363,N_3292,N_3240);
nor U3364 (N_3364,N_3214,N_3249);
nor U3365 (N_3365,N_3296,N_3212);
nor U3366 (N_3366,N_3250,N_3274);
nor U3367 (N_3367,N_3224,N_3231);
and U3368 (N_3368,N_3230,N_3211);
nor U3369 (N_3369,N_3219,N_3283);
xnor U3370 (N_3370,N_3229,N_3279);
and U3371 (N_3371,N_3288,N_3283);
nand U3372 (N_3372,N_3222,N_3214);
nor U3373 (N_3373,N_3261,N_3293);
and U3374 (N_3374,N_3216,N_3221);
and U3375 (N_3375,N_3235,N_3204);
xor U3376 (N_3376,N_3212,N_3228);
and U3377 (N_3377,N_3237,N_3233);
nand U3378 (N_3378,N_3205,N_3271);
nand U3379 (N_3379,N_3241,N_3225);
nand U3380 (N_3380,N_3279,N_3292);
or U3381 (N_3381,N_3244,N_3259);
nand U3382 (N_3382,N_3207,N_3288);
xor U3383 (N_3383,N_3238,N_3253);
nand U3384 (N_3384,N_3282,N_3264);
nor U3385 (N_3385,N_3224,N_3281);
or U3386 (N_3386,N_3203,N_3205);
nor U3387 (N_3387,N_3256,N_3294);
or U3388 (N_3388,N_3209,N_3296);
or U3389 (N_3389,N_3285,N_3235);
nand U3390 (N_3390,N_3231,N_3222);
nand U3391 (N_3391,N_3282,N_3216);
xnor U3392 (N_3392,N_3264,N_3206);
and U3393 (N_3393,N_3207,N_3271);
nand U3394 (N_3394,N_3288,N_3213);
nand U3395 (N_3395,N_3266,N_3279);
and U3396 (N_3396,N_3234,N_3287);
xnor U3397 (N_3397,N_3289,N_3216);
or U3398 (N_3398,N_3204,N_3209);
nor U3399 (N_3399,N_3260,N_3234);
nor U3400 (N_3400,N_3333,N_3380);
xor U3401 (N_3401,N_3370,N_3308);
nor U3402 (N_3402,N_3394,N_3302);
nand U3403 (N_3403,N_3320,N_3397);
nor U3404 (N_3404,N_3372,N_3387);
nand U3405 (N_3405,N_3356,N_3311);
and U3406 (N_3406,N_3393,N_3352);
xor U3407 (N_3407,N_3385,N_3382);
nor U3408 (N_3408,N_3378,N_3319);
nor U3409 (N_3409,N_3339,N_3326);
nand U3410 (N_3410,N_3371,N_3399);
nand U3411 (N_3411,N_3316,N_3310);
and U3412 (N_3412,N_3373,N_3367);
or U3413 (N_3413,N_3301,N_3366);
nand U3414 (N_3414,N_3318,N_3345);
nand U3415 (N_3415,N_3328,N_3369);
and U3416 (N_3416,N_3355,N_3358);
nor U3417 (N_3417,N_3376,N_3312);
or U3418 (N_3418,N_3331,N_3325);
nand U3419 (N_3419,N_3306,N_3364);
and U3420 (N_3420,N_3315,N_3353);
nand U3421 (N_3421,N_3354,N_3321);
and U3422 (N_3422,N_3349,N_3343);
xor U3423 (N_3423,N_3392,N_3322);
or U3424 (N_3424,N_3346,N_3340);
nand U3425 (N_3425,N_3383,N_3335);
and U3426 (N_3426,N_3361,N_3327);
or U3427 (N_3427,N_3300,N_3307);
nand U3428 (N_3428,N_3304,N_3388);
and U3429 (N_3429,N_3374,N_3332);
and U3430 (N_3430,N_3330,N_3395);
nor U3431 (N_3431,N_3363,N_3303);
xor U3432 (N_3432,N_3379,N_3350);
xor U3433 (N_3433,N_3381,N_3375);
and U3434 (N_3434,N_3314,N_3398);
nor U3435 (N_3435,N_3309,N_3323);
or U3436 (N_3436,N_3337,N_3386);
nor U3437 (N_3437,N_3351,N_3359);
nand U3438 (N_3438,N_3344,N_3317);
xnor U3439 (N_3439,N_3342,N_3324);
nor U3440 (N_3440,N_3384,N_3390);
nand U3441 (N_3441,N_3334,N_3305);
nor U3442 (N_3442,N_3329,N_3336);
nand U3443 (N_3443,N_3347,N_3389);
nor U3444 (N_3444,N_3341,N_3338);
nand U3445 (N_3445,N_3348,N_3396);
nor U3446 (N_3446,N_3368,N_3362);
and U3447 (N_3447,N_3391,N_3357);
nor U3448 (N_3448,N_3313,N_3377);
nor U3449 (N_3449,N_3360,N_3365);
or U3450 (N_3450,N_3326,N_3394);
nor U3451 (N_3451,N_3379,N_3388);
nand U3452 (N_3452,N_3355,N_3330);
xnor U3453 (N_3453,N_3374,N_3397);
and U3454 (N_3454,N_3376,N_3383);
nand U3455 (N_3455,N_3340,N_3377);
and U3456 (N_3456,N_3350,N_3317);
xor U3457 (N_3457,N_3394,N_3337);
nand U3458 (N_3458,N_3386,N_3369);
nand U3459 (N_3459,N_3353,N_3326);
nand U3460 (N_3460,N_3366,N_3300);
nand U3461 (N_3461,N_3384,N_3323);
xor U3462 (N_3462,N_3361,N_3351);
xnor U3463 (N_3463,N_3359,N_3395);
nand U3464 (N_3464,N_3348,N_3371);
nand U3465 (N_3465,N_3346,N_3373);
or U3466 (N_3466,N_3305,N_3324);
or U3467 (N_3467,N_3375,N_3301);
and U3468 (N_3468,N_3385,N_3323);
nor U3469 (N_3469,N_3302,N_3386);
xnor U3470 (N_3470,N_3363,N_3349);
or U3471 (N_3471,N_3397,N_3353);
or U3472 (N_3472,N_3361,N_3374);
and U3473 (N_3473,N_3343,N_3389);
nor U3474 (N_3474,N_3357,N_3336);
and U3475 (N_3475,N_3347,N_3357);
and U3476 (N_3476,N_3312,N_3346);
nor U3477 (N_3477,N_3331,N_3393);
or U3478 (N_3478,N_3396,N_3398);
nand U3479 (N_3479,N_3367,N_3300);
nor U3480 (N_3480,N_3319,N_3333);
nor U3481 (N_3481,N_3334,N_3364);
and U3482 (N_3482,N_3380,N_3312);
nand U3483 (N_3483,N_3322,N_3367);
and U3484 (N_3484,N_3373,N_3321);
nand U3485 (N_3485,N_3371,N_3327);
xnor U3486 (N_3486,N_3367,N_3311);
nand U3487 (N_3487,N_3329,N_3370);
nand U3488 (N_3488,N_3384,N_3321);
nor U3489 (N_3489,N_3377,N_3353);
and U3490 (N_3490,N_3342,N_3362);
xnor U3491 (N_3491,N_3362,N_3366);
xor U3492 (N_3492,N_3364,N_3303);
or U3493 (N_3493,N_3366,N_3394);
nor U3494 (N_3494,N_3399,N_3300);
xor U3495 (N_3495,N_3308,N_3346);
nand U3496 (N_3496,N_3399,N_3396);
xor U3497 (N_3497,N_3363,N_3393);
or U3498 (N_3498,N_3305,N_3329);
and U3499 (N_3499,N_3388,N_3375);
or U3500 (N_3500,N_3491,N_3472);
and U3501 (N_3501,N_3441,N_3422);
and U3502 (N_3502,N_3405,N_3487);
nor U3503 (N_3503,N_3461,N_3476);
and U3504 (N_3504,N_3482,N_3462);
xor U3505 (N_3505,N_3447,N_3416);
or U3506 (N_3506,N_3481,N_3449);
nor U3507 (N_3507,N_3408,N_3429);
and U3508 (N_3508,N_3460,N_3415);
or U3509 (N_3509,N_3485,N_3411);
or U3510 (N_3510,N_3403,N_3438);
nand U3511 (N_3511,N_3423,N_3496);
nand U3512 (N_3512,N_3488,N_3486);
and U3513 (N_3513,N_3459,N_3465);
or U3514 (N_3514,N_3432,N_3484);
or U3515 (N_3515,N_3418,N_3477);
and U3516 (N_3516,N_3412,N_3499);
xor U3517 (N_3517,N_3444,N_3446);
xor U3518 (N_3518,N_3448,N_3410);
and U3519 (N_3519,N_3435,N_3419);
xor U3520 (N_3520,N_3421,N_3494);
nor U3521 (N_3521,N_3427,N_3458);
nand U3522 (N_3522,N_3467,N_3468);
and U3523 (N_3523,N_3436,N_3406);
nand U3524 (N_3524,N_3475,N_3439);
nand U3525 (N_3525,N_3431,N_3466);
nor U3526 (N_3526,N_3450,N_3464);
and U3527 (N_3527,N_3492,N_3433);
nand U3528 (N_3528,N_3471,N_3497);
and U3529 (N_3529,N_3453,N_3498);
nand U3530 (N_3530,N_3440,N_3489);
nand U3531 (N_3531,N_3474,N_3455);
nand U3532 (N_3532,N_3493,N_3457);
nor U3533 (N_3533,N_3400,N_3420);
nor U3534 (N_3534,N_3495,N_3437);
xor U3535 (N_3535,N_3480,N_3434);
nand U3536 (N_3536,N_3479,N_3451);
and U3537 (N_3537,N_3407,N_3401);
nor U3538 (N_3538,N_3424,N_3456);
nand U3539 (N_3539,N_3470,N_3490);
nor U3540 (N_3540,N_3430,N_3409);
xor U3541 (N_3541,N_3452,N_3454);
nand U3542 (N_3542,N_3413,N_3414);
nand U3543 (N_3543,N_3483,N_3442);
xnor U3544 (N_3544,N_3417,N_3463);
and U3545 (N_3545,N_3469,N_3473);
nand U3546 (N_3546,N_3425,N_3478);
or U3547 (N_3547,N_3426,N_3443);
xnor U3548 (N_3548,N_3402,N_3445);
nand U3549 (N_3549,N_3404,N_3428);
xnor U3550 (N_3550,N_3454,N_3468);
and U3551 (N_3551,N_3472,N_3445);
xor U3552 (N_3552,N_3418,N_3423);
nor U3553 (N_3553,N_3417,N_3427);
nor U3554 (N_3554,N_3401,N_3455);
xor U3555 (N_3555,N_3499,N_3492);
xnor U3556 (N_3556,N_3478,N_3451);
nand U3557 (N_3557,N_3493,N_3427);
xor U3558 (N_3558,N_3465,N_3480);
and U3559 (N_3559,N_3430,N_3416);
or U3560 (N_3560,N_3404,N_3477);
nand U3561 (N_3561,N_3425,N_3436);
nor U3562 (N_3562,N_3496,N_3499);
nor U3563 (N_3563,N_3487,N_3447);
nor U3564 (N_3564,N_3456,N_3455);
and U3565 (N_3565,N_3474,N_3435);
or U3566 (N_3566,N_3412,N_3402);
nor U3567 (N_3567,N_3426,N_3415);
xnor U3568 (N_3568,N_3416,N_3491);
or U3569 (N_3569,N_3456,N_3436);
and U3570 (N_3570,N_3441,N_3434);
nor U3571 (N_3571,N_3489,N_3441);
nor U3572 (N_3572,N_3464,N_3466);
or U3573 (N_3573,N_3462,N_3451);
xnor U3574 (N_3574,N_3431,N_3493);
nand U3575 (N_3575,N_3468,N_3461);
nand U3576 (N_3576,N_3410,N_3490);
nand U3577 (N_3577,N_3406,N_3469);
or U3578 (N_3578,N_3431,N_3467);
xnor U3579 (N_3579,N_3431,N_3492);
nand U3580 (N_3580,N_3439,N_3472);
nand U3581 (N_3581,N_3477,N_3478);
nor U3582 (N_3582,N_3450,N_3484);
or U3583 (N_3583,N_3403,N_3457);
xor U3584 (N_3584,N_3477,N_3466);
xor U3585 (N_3585,N_3496,N_3489);
nand U3586 (N_3586,N_3422,N_3427);
and U3587 (N_3587,N_3481,N_3489);
nand U3588 (N_3588,N_3477,N_3407);
or U3589 (N_3589,N_3427,N_3434);
and U3590 (N_3590,N_3425,N_3442);
xnor U3591 (N_3591,N_3471,N_3492);
nor U3592 (N_3592,N_3464,N_3446);
and U3593 (N_3593,N_3481,N_3445);
xor U3594 (N_3594,N_3414,N_3476);
nand U3595 (N_3595,N_3429,N_3495);
xor U3596 (N_3596,N_3471,N_3425);
and U3597 (N_3597,N_3424,N_3468);
xnor U3598 (N_3598,N_3490,N_3408);
and U3599 (N_3599,N_3490,N_3458);
or U3600 (N_3600,N_3576,N_3517);
xnor U3601 (N_3601,N_3572,N_3563);
nor U3602 (N_3602,N_3593,N_3552);
nor U3603 (N_3603,N_3573,N_3529);
nand U3604 (N_3604,N_3500,N_3519);
and U3605 (N_3605,N_3559,N_3532);
nand U3606 (N_3606,N_3558,N_3579);
xnor U3607 (N_3607,N_3536,N_3587);
and U3608 (N_3608,N_3585,N_3537);
nor U3609 (N_3609,N_3538,N_3518);
nand U3610 (N_3610,N_3592,N_3509);
and U3611 (N_3611,N_3578,N_3597);
and U3612 (N_3612,N_3503,N_3551);
nor U3613 (N_3613,N_3542,N_3520);
nand U3614 (N_3614,N_3553,N_3535);
nor U3615 (N_3615,N_3512,N_3511);
or U3616 (N_3616,N_3556,N_3504);
nor U3617 (N_3617,N_3505,N_3568);
nor U3618 (N_3618,N_3575,N_3571);
xor U3619 (N_3619,N_3540,N_3595);
and U3620 (N_3620,N_3560,N_3521);
xnor U3621 (N_3621,N_3580,N_3510);
or U3622 (N_3622,N_3530,N_3533);
nand U3623 (N_3623,N_3539,N_3544);
or U3624 (N_3624,N_3590,N_3557);
or U3625 (N_3625,N_3531,N_3589);
and U3626 (N_3626,N_3569,N_3583);
or U3627 (N_3627,N_3507,N_3513);
and U3628 (N_3628,N_3577,N_3574);
or U3629 (N_3629,N_3526,N_3516);
or U3630 (N_3630,N_3514,N_3570);
or U3631 (N_3631,N_3525,N_3528);
nand U3632 (N_3632,N_3588,N_3502);
nor U3633 (N_3633,N_3554,N_3566);
or U3634 (N_3634,N_3501,N_3506);
xnor U3635 (N_3635,N_3548,N_3594);
nor U3636 (N_3636,N_3543,N_3586);
or U3637 (N_3637,N_3534,N_3567);
or U3638 (N_3638,N_3522,N_3584);
nand U3639 (N_3639,N_3565,N_3527);
nor U3640 (N_3640,N_3598,N_3541);
xnor U3641 (N_3641,N_3596,N_3523);
nand U3642 (N_3642,N_3550,N_3545);
nand U3643 (N_3643,N_3599,N_3515);
nand U3644 (N_3644,N_3591,N_3582);
or U3645 (N_3645,N_3561,N_3546);
nand U3646 (N_3646,N_3547,N_3524);
and U3647 (N_3647,N_3549,N_3581);
or U3648 (N_3648,N_3564,N_3555);
or U3649 (N_3649,N_3562,N_3508);
xnor U3650 (N_3650,N_3545,N_3515);
xor U3651 (N_3651,N_3513,N_3527);
and U3652 (N_3652,N_3551,N_3528);
xnor U3653 (N_3653,N_3552,N_3548);
or U3654 (N_3654,N_3587,N_3557);
nor U3655 (N_3655,N_3559,N_3561);
nand U3656 (N_3656,N_3583,N_3595);
and U3657 (N_3657,N_3586,N_3578);
xor U3658 (N_3658,N_3589,N_3587);
xnor U3659 (N_3659,N_3541,N_3553);
and U3660 (N_3660,N_3590,N_3506);
nand U3661 (N_3661,N_3529,N_3596);
xnor U3662 (N_3662,N_3567,N_3574);
xnor U3663 (N_3663,N_3530,N_3573);
xnor U3664 (N_3664,N_3532,N_3544);
and U3665 (N_3665,N_3508,N_3560);
xnor U3666 (N_3666,N_3514,N_3521);
xnor U3667 (N_3667,N_3545,N_3551);
nand U3668 (N_3668,N_3580,N_3503);
xnor U3669 (N_3669,N_3577,N_3504);
nor U3670 (N_3670,N_3504,N_3598);
nand U3671 (N_3671,N_3579,N_3546);
or U3672 (N_3672,N_3566,N_3502);
xor U3673 (N_3673,N_3517,N_3508);
nand U3674 (N_3674,N_3590,N_3565);
nor U3675 (N_3675,N_3557,N_3516);
and U3676 (N_3676,N_3596,N_3586);
nor U3677 (N_3677,N_3532,N_3553);
nor U3678 (N_3678,N_3597,N_3516);
xnor U3679 (N_3679,N_3519,N_3576);
and U3680 (N_3680,N_3517,N_3512);
or U3681 (N_3681,N_3508,N_3575);
or U3682 (N_3682,N_3593,N_3555);
nand U3683 (N_3683,N_3584,N_3573);
nor U3684 (N_3684,N_3571,N_3599);
nand U3685 (N_3685,N_3554,N_3523);
nand U3686 (N_3686,N_3514,N_3584);
and U3687 (N_3687,N_3510,N_3597);
or U3688 (N_3688,N_3524,N_3515);
or U3689 (N_3689,N_3512,N_3553);
or U3690 (N_3690,N_3536,N_3598);
and U3691 (N_3691,N_3595,N_3596);
and U3692 (N_3692,N_3578,N_3528);
and U3693 (N_3693,N_3550,N_3573);
and U3694 (N_3694,N_3528,N_3529);
xor U3695 (N_3695,N_3519,N_3545);
and U3696 (N_3696,N_3523,N_3565);
or U3697 (N_3697,N_3522,N_3582);
and U3698 (N_3698,N_3515,N_3587);
nor U3699 (N_3699,N_3544,N_3540);
nand U3700 (N_3700,N_3679,N_3663);
and U3701 (N_3701,N_3642,N_3631);
or U3702 (N_3702,N_3659,N_3625);
or U3703 (N_3703,N_3657,N_3675);
and U3704 (N_3704,N_3695,N_3619);
nand U3705 (N_3705,N_3614,N_3684);
nor U3706 (N_3706,N_3694,N_3674);
xor U3707 (N_3707,N_3683,N_3600);
nor U3708 (N_3708,N_3639,N_3635);
nand U3709 (N_3709,N_3611,N_3665);
and U3710 (N_3710,N_3612,N_3686);
or U3711 (N_3711,N_3664,N_3670);
nand U3712 (N_3712,N_3698,N_3681);
or U3713 (N_3713,N_3638,N_3602);
or U3714 (N_3714,N_3653,N_3692);
nand U3715 (N_3715,N_3610,N_3699);
or U3716 (N_3716,N_3615,N_3633);
xor U3717 (N_3717,N_3676,N_3624);
or U3718 (N_3718,N_3666,N_3628);
nor U3719 (N_3719,N_3691,N_3608);
or U3720 (N_3720,N_3667,N_3649);
xnor U3721 (N_3721,N_3603,N_3644);
xnor U3722 (N_3722,N_3605,N_3641);
nand U3723 (N_3723,N_3623,N_3671);
and U3724 (N_3724,N_3688,N_3616);
or U3725 (N_3725,N_3622,N_3689);
nor U3726 (N_3726,N_3647,N_3621);
nand U3727 (N_3727,N_3696,N_3673);
xor U3728 (N_3728,N_3636,N_3620);
nand U3729 (N_3729,N_3643,N_3651);
nand U3730 (N_3730,N_3661,N_3656);
xnor U3731 (N_3731,N_3654,N_3680);
nand U3732 (N_3732,N_3618,N_3662);
or U3733 (N_3733,N_3630,N_3645);
nand U3734 (N_3734,N_3617,N_3668);
nor U3735 (N_3735,N_3601,N_3660);
and U3736 (N_3736,N_3658,N_3646);
and U3737 (N_3737,N_3613,N_3693);
nor U3738 (N_3738,N_3652,N_3690);
nand U3739 (N_3739,N_3607,N_3678);
nor U3740 (N_3740,N_3648,N_3626);
nor U3741 (N_3741,N_3669,N_3627);
nand U3742 (N_3742,N_3697,N_3629);
and U3743 (N_3743,N_3634,N_3606);
xor U3744 (N_3744,N_3609,N_3672);
xnor U3745 (N_3745,N_3685,N_3637);
nor U3746 (N_3746,N_3655,N_3640);
and U3747 (N_3747,N_3682,N_3604);
or U3748 (N_3748,N_3650,N_3632);
and U3749 (N_3749,N_3677,N_3687);
nand U3750 (N_3750,N_3635,N_3656);
nand U3751 (N_3751,N_3673,N_3677);
xnor U3752 (N_3752,N_3641,N_3669);
xnor U3753 (N_3753,N_3630,N_3620);
or U3754 (N_3754,N_3675,N_3635);
nand U3755 (N_3755,N_3645,N_3694);
nor U3756 (N_3756,N_3614,N_3612);
or U3757 (N_3757,N_3670,N_3656);
xnor U3758 (N_3758,N_3683,N_3623);
nor U3759 (N_3759,N_3604,N_3678);
nor U3760 (N_3760,N_3620,N_3617);
nand U3761 (N_3761,N_3667,N_3697);
or U3762 (N_3762,N_3631,N_3675);
xnor U3763 (N_3763,N_3651,N_3668);
nor U3764 (N_3764,N_3610,N_3623);
and U3765 (N_3765,N_3636,N_3691);
nand U3766 (N_3766,N_3657,N_3685);
xor U3767 (N_3767,N_3612,N_3645);
nor U3768 (N_3768,N_3630,N_3665);
nor U3769 (N_3769,N_3615,N_3602);
or U3770 (N_3770,N_3626,N_3692);
xor U3771 (N_3771,N_3685,N_3676);
or U3772 (N_3772,N_3614,N_3601);
and U3773 (N_3773,N_3668,N_3665);
nor U3774 (N_3774,N_3694,N_3644);
nor U3775 (N_3775,N_3618,N_3670);
or U3776 (N_3776,N_3659,N_3651);
nor U3777 (N_3777,N_3692,N_3674);
and U3778 (N_3778,N_3698,N_3696);
nor U3779 (N_3779,N_3685,N_3631);
or U3780 (N_3780,N_3636,N_3607);
or U3781 (N_3781,N_3640,N_3692);
nor U3782 (N_3782,N_3694,N_3613);
nor U3783 (N_3783,N_3679,N_3677);
nand U3784 (N_3784,N_3673,N_3688);
or U3785 (N_3785,N_3680,N_3699);
xnor U3786 (N_3786,N_3668,N_3611);
and U3787 (N_3787,N_3635,N_3633);
and U3788 (N_3788,N_3673,N_3641);
and U3789 (N_3789,N_3633,N_3668);
xor U3790 (N_3790,N_3645,N_3693);
or U3791 (N_3791,N_3609,N_3602);
nand U3792 (N_3792,N_3699,N_3692);
and U3793 (N_3793,N_3693,N_3617);
or U3794 (N_3794,N_3617,N_3600);
nor U3795 (N_3795,N_3662,N_3610);
nor U3796 (N_3796,N_3604,N_3676);
and U3797 (N_3797,N_3695,N_3667);
nor U3798 (N_3798,N_3697,N_3646);
nor U3799 (N_3799,N_3631,N_3643);
xor U3800 (N_3800,N_3789,N_3737);
nor U3801 (N_3801,N_3746,N_3743);
nand U3802 (N_3802,N_3723,N_3780);
or U3803 (N_3803,N_3742,N_3795);
or U3804 (N_3804,N_3768,N_3765);
or U3805 (N_3805,N_3711,N_3745);
xor U3806 (N_3806,N_3747,N_3721);
nor U3807 (N_3807,N_3770,N_3740);
nor U3808 (N_3808,N_3709,N_3787);
or U3809 (N_3809,N_3718,N_3762);
or U3810 (N_3810,N_3728,N_3794);
nand U3811 (N_3811,N_3790,N_3705);
xnor U3812 (N_3812,N_3776,N_3782);
or U3813 (N_3813,N_3727,N_3793);
xnor U3814 (N_3814,N_3708,N_3753);
xor U3815 (N_3815,N_3706,N_3710);
xnor U3816 (N_3816,N_3717,N_3730);
or U3817 (N_3817,N_3757,N_3763);
nand U3818 (N_3818,N_3777,N_3749);
and U3819 (N_3819,N_3760,N_3702);
nand U3820 (N_3820,N_3736,N_3720);
nor U3821 (N_3821,N_3738,N_3771);
nand U3822 (N_3822,N_3761,N_3755);
and U3823 (N_3823,N_3759,N_3739);
nand U3824 (N_3824,N_3734,N_3773);
nand U3825 (N_3825,N_3722,N_3781);
or U3826 (N_3826,N_3733,N_3701);
nand U3827 (N_3827,N_3791,N_3798);
and U3828 (N_3828,N_3792,N_3741);
nor U3829 (N_3829,N_3783,N_3724);
nand U3830 (N_3830,N_3750,N_3799);
or U3831 (N_3831,N_3796,N_3744);
nor U3832 (N_3832,N_3731,N_3719);
nand U3833 (N_3833,N_3713,N_3729);
nand U3834 (N_3834,N_3788,N_3779);
and U3835 (N_3835,N_3700,N_3707);
nand U3836 (N_3836,N_3774,N_3758);
or U3837 (N_3837,N_3732,N_3769);
nor U3838 (N_3838,N_3797,N_3764);
or U3839 (N_3839,N_3784,N_3712);
xor U3840 (N_3840,N_3766,N_3714);
nand U3841 (N_3841,N_3751,N_3726);
or U3842 (N_3842,N_3775,N_3785);
nor U3843 (N_3843,N_3703,N_3756);
nand U3844 (N_3844,N_3704,N_3778);
nand U3845 (N_3845,N_3754,N_3725);
nand U3846 (N_3846,N_3772,N_3735);
xor U3847 (N_3847,N_3716,N_3715);
and U3848 (N_3848,N_3752,N_3767);
nor U3849 (N_3849,N_3786,N_3748);
nor U3850 (N_3850,N_3749,N_3757);
xor U3851 (N_3851,N_3715,N_3705);
nor U3852 (N_3852,N_3736,N_3755);
xor U3853 (N_3853,N_3712,N_3754);
nand U3854 (N_3854,N_3770,N_3705);
nand U3855 (N_3855,N_3750,N_3715);
xor U3856 (N_3856,N_3729,N_3749);
xnor U3857 (N_3857,N_3764,N_3777);
nor U3858 (N_3858,N_3734,N_3794);
nor U3859 (N_3859,N_3717,N_3721);
nand U3860 (N_3860,N_3747,N_3780);
or U3861 (N_3861,N_3740,N_3730);
nand U3862 (N_3862,N_3737,N_3776);
nor U3863 (N_3863,N_3719,N_3770);
and U3864 (N_3864,N_3718,N_3730);
nand U3865 (N_3865,N_3782,N_3727);
nor U3866 (N_3866,N_3731,N_3770);
xor U3867 (N_3867,N_3773,N_3700);
and U3868 (N_3868,N_3759,N_3790);
nand U3869 (N_3869,N_3726,N_3717);
nor U3870 (N_3870,N_3754,N_3756);
nor U3871 (N_3871,N_3795,N_3707);
or U3872 (N_3872,N_3730,N_3709);
xnor U3873 (N_3873,N_3708,N_3792);
xor U3874 (N_3874,N_3776,N_3733);
nor U3875 (N_3875,N_3740,N_3783);
xor U3876 (N_3876,N_3789,N_3778);
nor U3877 (N_3877,N_3736,N_3794);
nor U3878 (N_3878,N_3781,N_3773);
or U3879 (N_3879,N_3789,N_3747);
xnor U3880 (N_3880,N_3702,N_3741);
nor U3881 (N_3881,N_3728,N_3702);
xnor U3882 (N_3882,N_3724,N_3742);
nor U3883 (N_3883,N_3726,N_3747);
or U3884 (N_3884,N_3712,N_3729);
nor U3885 (N_3885,N_3777,N_3714);
xnor U3886 (N_3886,N_3755,N_3708);
and U3887 (N_3887,N_3776,N_3730);
xnor U3888 (N_3888,N_3754,N_3731);
and U3889 (N_3889,N_3746,N_3786);
nand U3890 (N_3890,N_3788,N_3765);
or U3891 (N_3891,N_3748,N_3708);
and U3892 (N_3892,N_3774,N_3711);
or U3893 (N_3893,N_3774,N_3755);
nor U3894 (N_3894,N_3788,N_3738);
nand U3895 (N_3895,N_3719,N_3796);
and U3896 (N_3896,N_3782,N_3752);
and U3897 (N_3897,N_3743,N_3793);
xor U3898 (N_3898,N_3739,N_3744);
and U3899 (N_3899,N_3712,N_3795);
or U3900 (N_3900,N_3814,N_3859);
xor U3901 (N_3901,N_3832,N_3892);
nor U3902 (N_3902,N_3851,N_3835);
or U3903 (N_3903,N_3850,N_3816);
nor U3904 (N_3904,N_3868,N_3883);
nand U3905 (N_3905,N_3808,N_3857);
nand U3906 (N_3906,N_3800,N_3824);
xnor U3907 (N_3907,N_3890,N_3811);
or U3908 (N_3908,N_3879,N_3878);
nand U3909 (N_3909,N_3858,N_3867);
or U3910 (N_3910,N_3821,N_3887);
nand U3911 (N_3911,N_3802,N_3813);
or U3912 (N_3912,N_3809,N_3864);
or U3913 (N_3913,N_3803,N_3815);
xnor U3914 (N_3914,N_3860,N_3880);
xor U3915 (N_3915,N_3836,N_3854);
and U3916 (N_3916,N_3898,N_3889);
and U3917 (N_3917,N_3845,N_3818);
nor U3918 (N_3918,N_3899,N_3897);
nor U3919 (N_3919,N_3846,N_3877);
nor U3920 (N_3920,N_3825,N_3822);
or U3921 (N_3921,N_3812,N_3861);
nor U3922 (N_3922,N_3831,N_3820);
xnor U3923 (N_3923,N_3838,N_3801);
or U3924 (N_3924,N_3847,N_3894);
or U3925 (N_3925,N_3893,N_3834);
nand U3926 (N_3926,N_3870,N_3823);
nand U3927 (N_3927,N_3863,N_3827);
and U3928 (N_3928,N_3848,N_3826);
and U3929 (N_3929,N_3895,N_3817);
nand U3930 (N_3930,N_3866,N_3853);
or U3931 (N_3931,N_3852,N_3830);
or U3932 (N_3932,N_3807,N_3841);
nand U3933 (N_3933,N_3882,N_3873);
nor U3934 (N_3934,N_3810,N_3885);
and U3935 (N_3935,N_3855,N_3856);
xor U3936 (N_3936,N_3839,N_3872);
nand U3937 (N_3937,N_3819,N_3828);
xor U3938 (N_3938,N_3875,N_3804);
nand U3939 (N_3939,N_3874,N_3806);
and U3940 (N_3940,N_3884,N_3849);
and U3941 (N_3941,N_3876,N_3842);
and U3942 (N_3942,N_3840,N_3886);
nand U3943 (N_3943,N_3871,N_3869);
nand U3944 (N_3944,N_3891,N_3805);
nand U3945 (N_3945,N_3862,N_3888);
nor U3946 (N_3946,N_3829,N_3865);
nor U3947 (N_3947,N_3837,N_3896);
or U3948 (N_3948,N_3833,N_3844);
and U3949 (N_3949,N_3843,N_3881);
nor U3950 (N_3950,N_3892,N_3808);
nor U3951 (N_3951,N_3810,N_3804);
or U3952 (N_3952,N_3862,N_3859);
nor U3953 (N_3953,N_3844,N_3867);
xnor U3954 (N_3954,N_3865,N_3888);
nor U3955 (N_3955,N_3878,N_3895);
and U3956 (N_3956,N_3868,N_3896);
or U3957 (N_3957,N_3865,N_3852);
nor U3958 (N_3958,N_3803,N_3822);
or U3959 (N_3959,N_3801,N_3873);
and U3960 (N_3960,N_3832,N_3899);
nand U3961 (N_3961,N_3862,N_3820);
or U3962 (N_3962,N_3898,N_3873);
xor U3963 (N_3963,N_3883,N_3839);
nor U3964 (N_3964,N_3818,N_3811);
and U3965 (N_3965,N_3827,N_3871);
nand U3966 (N_3966,N_3865,N_3858);
nand U3967 (N_3967,N_3897,N_3839);
xnor U3968 (N_3968,N_3824,N_3876);
xor U3969 (N_3969,N_3807,N_3852);
nor U3970 (N_3970,N_3888,N_3831);
nor U3971 (N_3971,N_3842,N_3884);
and U3972 (N_3972,N_3801,N_3889);
nand U3973 (N_3973,N_3833,N_3875);
nor U3974 (N_3974,N_3829,N_3828);
nor U3975 (N_3975,N_3831,N_3893);
xor U3976 (N_3976,N_3898,N_3883);
nand U3977 (N_3977,N_3884,N_3809);
and U3978 (N_3978,N_3848,N_3859);
nand U3979 (N_3979,N_3876,N_3840);
nand U3980 (N_3980,N_3889,N_3827);
xor U3981 (N_3981,N_3875,N_3892);
or U3982 (N_3982,N_3837,N_3848);
nand U3983 (N_3983,N_3875,N_3885);
nand U3984 (N_3984,N_3863,N_3831);
nand U3985 (N_3985,N_3801,N_3824);
nor U3986 (N_3986,N_3822,N_3846);
nand U3987 (N_3987,N_3827,N_3855);
or U3988 (N_3988,N_3862,N_3864);
or U3989 (N_3989,N_3888,N_3833);
xnor U3990 (N_3990,N_3803,N_3841);
nand U3991 (N_3991,N_3895,N_3807);
nand U3992 (N_3992,N_3801,N_3814);
or U3993 (N_3993,N_3847,N_3827);
or U3994 (N_3994,N_3836,N_3824);
xor U3995 (N_3995,N_3850,N_3822);
nand U3996 (N_3996,N_3831,N_3825);
and U3997 (N_3997,N_3883,N_3842);
nor U3998 (N_3998,N_3827,N_3803);
nor U3999 (N_3999,N_3892,N_3807);
and U4000 (N_4000,N_3980,N_3959);
and U4001 (N_4001,N_3939,N_3988);
nor U4002 (N_4002,N_3943,N_3905);
nand U4003 (N_4003,N_3985,N_3964);
nor U4004 (N_4004,N_3933,N_3950);
or U4005 (N_4005,N_3912,N_3999);
xor U4006 (N_4006,N_3962,N_3955);
and U4007 (N_4007,N_3983,N_3917);
nor U4008 (N_4008,N_3976,N_3995);
or U4009 (N_4009,N_3913,N_3963);
or U4010 (N_4010,N_3987,N_3931);
and U4011 (N_4011,N_3982,N_3970);
nor U4012 (N_4012,N_3938,N_3945);
nand U4013 (N_4013,N_3903,N_3975);
nand U4014 (N_4014,N_3919,N_3902);
or U4015 (N_4015,N_3918,N_3952);
and U4016 (N_4016,N_3986,N_3991);
and U4017 (N_4017,N_3923,N_3935);
nor U4018 (N_4018,N_3993,N_3990);
and U4019 (N_4019,N_3930,N_3900);
nand U4020 (N_4020,N_3984,N_3911);
or U4021 (N_4021,N_3989,N_3994);
nor U4022 (N_4022,N_3960,N_3910);
or U4023 (N_4023,N_3973,N_3916);
or U4024 (N_4024,N_3937,N_3998);
nor U4025 (N_4025,N_3957,N_3934);
or U4026 (N_4026,N_3924,N_3958);
nor U4027 (N_4027,N_3954,N_3941);
or U4028 (N_4028,N_3904,N_3949);
nand U4029 (N_4029,N_3921,N_3974);
xnor U4030 (N_4030,N_3915,N_3926);
nand U4031 (N_4031,N_3997,N_3914);
nand U4032 (N_4032,N_3901,N_3925);
nand U4033 (N_4033,N_3981,N_3927);
nor U4034 (N_4034,N_3944,N_3996);
or U4035 (N_4035,N_3992,N_3920);
nand U4036 (N_4036,N_3946,N_3907);
xor U4037 (N_4037,N_3942,N_3951);
and U4038 (N_4038,N_3947,N_3948);
and U4039 (N_4039,N_3967,N_3906);
nor U4040 (N_4040,N_3953,N_3922);
or U4041 (N_4041,N_3940,N_3965);
nand U4042 (N_4042,N_3908,N_3979);
and U4043 (N_4043,N_3966,N_3968);
nand U4044 (N_4044,N_3936,N_3909);
nand U4045 (N_4045,N_3969,N_3977);
nor U4046 (N_4046,N_3972,N_3932);
nand U4047 (N_4047,N_3978,N_3929);
or U4048 (N_4048,N_3928,N_3971);
or U4049 (N_4049,N_3961,N_3956);
or U4050 (N_4050,N_3902,N_3922);
xor U4051 (N_4051,N_3941,N_3931);
or U4052 (N_4052,N_3987,N_3960);
nor U4053 (N_4053,N_3911,N_3927);
nand U4054 (N_4054,N_3932,N_3968);
or U4055 (N_4055,N_3968,N_3920);
nor U4056 (N_4056,N_3928,N_3974);
or U4057 (N_4057,N_3913,N_3938);
nand U4058 (N_4058,N_3912,N_3974);
nor U4059 (N_4059,N_3931,N_3962);
nor U4060 (N_4060,N_3974,N_3917);
xnor U4061 (N_4061,N_3911,N_3989);
nand U4062 (N_4062,N_3987,N_3923);
xnor U4063 (N_4063,N_3955,N_3945);
xnor U4064 (N_4064,N_3941,N_3952);
nand U4065 (N_4065,N_3974,N_3934);
or U4066 (N_4066,N_3934,N_3977);
nand U4067 (N_4067,N_3914,N_3915);
and U4068 (N_4068,N_3994,N_3930);
and U4069 (N_4069,N_3965,N_3941);
and U4070 (N_4070,N_3916,N_3987);
nand U4071 (N_4071,N_3985,N_3931);
and U4072 (N_4072,N_3927,N_3935);
or U4073 (N_4073,N_3946,N_3913);
nand U4074 (N_4074,N_3903,N_3950);
or U4075 (N_4075,N_3955,N_3926);
or U4076 (N_4076,N_3992,N_3934);
or U4077 (N_4077,N_3981,N_3989);
nor U4078 (N_4078,N_3927,N_3931);
and U4079 (N_4079,N_3996,N_3986);
and U4080 (N_4080,N_3937,N_3974);
xnor U4081 (N_4081,N_3953,N_3995);
nor U4082 (N_4082,N_3947,N_3995);
and U4083 (N_4083,N_3914,N_3924);
nor U4084 (N_4084,N_3958,N_3965);
nor U4085 (N_4085,N_3987,N_3915);
or U4086 (N_4086,N_3955,N_3917);
nand U4087 (N_4087,N_3912,N_3910);
nand U4088 (N_4088,N_3963,N_3960);
xnor U4089 (N_4089,N_3970,N_3904);
nand U4090 (N_4090,N_3975,N_3999);
and U4091 (N_4091,N_3967,N_3997);
nand U4092 (N_4092,N_3967,N_3976);
xnor U4093 (N_4093,N_3925,N_3960);
xnor U4094 (N_4094,N_3928,N_3998);
or U4095 (N_4095,N_3952,N_3989);
xor U4096 (N_4096,N_3905,N_3985);
xnor U4097 (N_4097,N_3969,N_3991);
nor U4098 (N_4098,N_3901,N_3966);
nor U4099 (N_4099,N_3923,N_3948);
and U4100 (N_4100,N_4022,N_4015);
xor U4101 (N_4101,N_4029,N_4007);
and U4102 (N_4102,N_4039,N_4071);
and U4103 (N_4103,N_4088,N_4092);
and U4104 (N_4104,N_4072,N_4035);
and U4105 (N_4105,N_4017,N_4012);
nor U4106 (N_4106,N_4043,N_4011);
and U4107 (N_4107,N_4079,N_4001);
nand U4108 (N_4108,N_4098,N_4009);
or U4109 (N_4109,N_4040,N_4060);
or U4110 (N_4110,N_4047,N_4036);
and U4111 (N_4111,N_4077,N_4010);
or U4112 (N_4112,N_4099,N_4055);
nor U4113 (N_4113,N_4090,N_4032);
or U4114 (N_4114,N_4059,N_4038);
nand U4115 (N_4115,N_4004,N_4034);
nor U4116 (N_4116,N_4084,N_4057);
and U4117 (N_4117,N_4003,N_4093);
and U4118 (N_4118,N_4014,N_4024);
nand U4119 (N_4119,N_4050,N_4086);
nor U4120 (N_4120,N_4065,N_4096);
nor U4121 (N_4121,N_4054,N_4042);
nor U4122 (N_4122,N_4094,N_4033);
nand U4123 (N_4123,N_4074,N_4051);
nand U4124 (N_4124,N_4095,N_4073);
nand U4125 (N_4125,N_4023,N_4026);
and U4126 (N_4126,N_4000,N_4052);
xnor U4127 (N_4127,N_4076,N_4031);
nand U4128 (N_4128,N_4068,N_4025);
or U4129 (N_4129,N_4030,N_4063);
or U4130 (N_4130,N_4082,N_4056);
nor U4131 (N_4131,N_4089,N_4002);
nand U4132 (N_4132,N_4006,N_4078);
and U4133 (N_4133,N_4048,N_4005);
nor U4134 (N_4134,N_4061,N_4021);
or U4135 (N_4135,N_4085,N_4027);
or U4136 (N_4136,N_4041,N_4067);
and U4137 (N_4137,N_4044,N_4062);
xnor U4138 (N_4138,N_4020,N_4070);
nor U4139 (N_4139,N_4087,N_4097);
nor U4140 (N_4140,N_4083,N_4075);
nor U4141 (N_4141,N_4046,N_4016);
nand U4142 (N_4142,N_4081,N_4028);
nor U4143 (N_4143,N_4018,N_4080);
xor U4144 (N_4144,N_4019,N_4045);
nor U4145 (N_4145,N_4069,N_4013);
and U4146 (N_4146,N_4049,N_4058);
xnor U4147 (N_4147,N_4066,N_4064);
or U4148 (N_4148,N_4091,N_4037);
nand U4149 (N_4149,N_4053,N_4008);
nor U4150 (N_4150,N_4065,N_4080);
nand U4151 (N_4151,N_4004,N_4078);
nor U4152 (N_4152,N_4039,N_4048);
xor U4153 (N_4153,N_4040,N_4049);
nand U4154 (N_4154,N_4056,N_4026);
nand U4155 (N_4155,N_4013,N_4017);
nor U4156 (N_4156,N_4030,N_4075);
nand U4157 (N_4157,N_4086,N_4003);
or U4158 (N_4158,N_4056,N_4071);
or U4159 (N_4159,N_4066,N_4003);
nor U4160 (N_4160,N_4058,N_4008);
and U4161 (N_4161,N_4094,N_4051);
nor U4162 (N_4162,N_4016,N_4035);
xor U4163 (N_4163,N_4088,N_4001);
xnor U4164 (N_4164,N_4083,N_4062);
xnor U4165 (N_4165,N_4006,N_4069);
and U4166 (N_4166,N_4031,N_4069);
or U4167 (N_4167,N_4046,N_4070);
xnor U4168 (N_4168,N_4001,N_4034);
nor U4169 (N_4169,N_4094,N_4016);
and U4170 (N_4170,N_4077,N_4012);
nor U4171 (N_4171,N_4010,N_4041);
or U4172 (N_4172,N_4011,N_4077);
and U4173 (N_4173,N_4065,N_4010);
or U4174 (N_4174,N_4032,N_4018);
nand U4175 (N_4175,N_4018,N_4020);
and U4176 (N_4176,N_4084,N_4082);
xnor U4177 (N_4177,N_4074,N_4093);
nand U4178 (N_4178,N_4089,N_4007);
or U4179 (N_4179,N_4033,N_4005);
nor U4180 (N_4180,N_4090,N_4089);
or U4181 (N_4181,N_4036,N_4003);
xnor U4182 (N_4182,N_4008,N_4044);
nor U4183 (N_4183,N_4052,N_4027);
and U4184 (N_4184,N_4082,N_4035);
xor U4185 (N_4185,N_4076,N_4074);
and U4186 (N_4186,N_4043,N_4072);
nor U4187 (N_4187,N_4082,N_4085);
nor U4188 (N_4188,N_4074,N_4033);
and U4189 (N_4189,N_4004,N_4056);
and U4190 (N_4190,N_4019,N_4088);
and U4191 (N_4191,N_4019,N_4014);
or U4192 (N_4192,N_4065,N_4013);
xor U4193 (N_4193,N_4029,N_4076);
or U4194 (N_4194,N_4009,N_4075);
or U4195 (N_4195,N_4076,N_4014);
nand U4196 (N_4196,N_4024,N_4015);
nor U4197 (N_4197,N_4094,N_4018);
nor U4198 (N_4198,N_4013,N_4049);
nor U4199 (N_4199,N_4056,N_4040);
nor U4200 (N_4200,N_4196,N_4153);
nor U4201 (N_4201,N_4195,N_4174);
nand U4202 (N_4202,N_4125,N_4118);
nor U4203 (N_4203,N_4127,N_4130);
nor U4204 (N_4204,N_4112,N_4168);
nand U4205 (N_4205,N_4110,N_4104);
nor U4206 (N_4206,N_4178,N_4117);
nor U4207 (N_4207,N_4140,N_4184);
nor U4208 (N_4208,N_4170,N_4129);
and U4209 (N_4209,N_4106,N_4144);
nor U4210 (N_4210,N_4142,N_4143);
or U4211 (N_4211,N_4182,N_4133);
nor U4212 (N_4212,N_4179,N_4165);
nor U4213 (N_4213,N_4186,N_4113);
xnor U4214 (N_4214,N_4134,N_4173);
nor U4215 (N_4215,N_4120,N_4157);
or U4216 (N_4216,N_4148,N_4149);
nor U4217 (N_4217,N_4183,N_4105);
xnor U4218 (N_4218,N_4181,N_4193);
xnor U4219 (N_4219,N_4187,N_4131);
xor U4220 (N_4220,N_4111,N_4145);
and U4221 (N_4221,N_4108,N_4188);
nor U4222 (N_4222,N_4156,N_4159);
or U4223 (N_4223,N_4139,N_4138);
xnor U4224 (N_4224,N_4198,N_4176);
or U4225 (N_4225,N_4132,N_4152);
and U4226 (N_4226,N_4147,N_4160);
and U4227 (N_4227,N_4162,N_4124);
nor U4228 (N_4228,N_4194,N_4128);
and U4229 (N_4229,N_4167,N_4126);
nor U4230 (N_4230,N_4123,N_4100);
nand U4231 (N_4231,N_4171,N_4172);
nor U4232 (N_4232,N_4150,N_4190);
xor U4233 (N_4233,N_4136,N_4169);
xnor U4234 (N_4234,N_4166,N_4175);
nand U4235 (N_4235,N_4191,N_4180);
and U4236 (N_4236,N_4102,N_4101);
or U4237 (N_4237,N_4107,N_4137);
nand U4238 (N_4238,N_4116,N_4121);
and U4239 (N_4239,N_4185,N_4158);
nand U4240 (N_4240,N_4177,N_4154);
xnor U4241 (N_4241,N_4103,N_4192);
nor U4242 (N_4242,N_4189,N_4114);
or U4243 (N_4243,N_4155,N_4122);
xor U4244 (N_4244,N_4119,N_4141);
xor U4245 (N_4245,N_4146,N_4151);
nor U4246 (N_4246,N_4135,N_4199);
or U4247 (N_4247,N_4164,N_4163);
xnor U4248 (N_4248,N_4115,N_4161);
xnor U4249 (N_4249,N_4109,N_4197);
nor U4250 (N_4250,N_4185,N_4165);
nor U4251 (N_4251,N_4173,N_4182);
nand U4252 (N_4252,N_4176,N_4150);
nand U4253 (N_4253,N_4186,N_4127);
xnor U4254 (N_4254,N_4141,N_4126);
nor U4255 (N_4255,N_4103,N_4146);
nand U4256 (N_4256,N_4195,N_4131);
and U4257 (N_4257,N_4166,N_4174);
nand U4258 (N_4258,N_4135,N_4198);
xor U4259 (N_4259,N_4196,N_4132);
nor U4260 (N_4260,N_4105,N_4157);
nand U4261 (N_4261,N_4102,N_4154);
nor U4262 (N_4262,N_4139,N_4152);
nor U4263 (N_4263,N_4123,N_4181);
xor U4264 (N_4264,N_4188,N_4118);
or U4265 (N_4265,N_4137,N_4171);
or U4266 (N_4266,N_4136,N_4177);
nand U4267 (N_4267,N_4112,N_4121);
or U4268 (N_4268,N_4171,N_4133);
or U4269 (N_4269,N_4195,N_4177);
nand U4270 (N_4270,N_4130,N_4171);
or U4271 (N_4271,N_4165,N_4105);
xor U4272 (N_4272,N_4157,N_4196);
nand U4273 (N_4273,N_4161,N_4126);
or U4274 (N_4274,N_4129,N_4156);
and U4275 (N_4275,N_4137,N_4160);
xnor U4276 (N_4276,N_4162,N_4174);
xor U4277 (N_4277,N_4153,N_4143);
xnor U4278 (N_4278,N_4119,N_4153);
and U4279 (N_4279,N_4122,N_4182);
or U4280 (N_4280,N_4149,N_4126);
or U4281 (N_4281,N_4176,N_4177);
and U4282 (N_4282,N_4177,N_4167);
xor U4283 (N_4283,N_4195,N_4157);
nor U4284 (N_4284,N_4100,N_4101);
nand U4285 (N_4285,N_4134,N_4114);
and U4286 (N_4286,N_4140,N_4145);
nand U4287 (N_4287,N_4109,N_4120);
nor U4288 (N_4288,N_4110,N_4151);
xor U4289 (N_4289,N_4114,N_4111);
or U4290 (N_4290,N_4129,N_4193);
or U4291 (N_4291,N_4124,N_4137);
xor U4292 (N_4292,N_4114,N_4183);
and U4293 (N_4293,N_4162,N_4131);
nor U4294 (N_4294,N_4164,N_4148);
nand U4295 (N_4295,N_4123,N_4116);
nand U4296 (N_4296,N_4132,N_4192);
nor U4297 (N_4297,N_4163,N_4147);
nand U4298 (N_4298,N_4138,N_4193);
nand U4299 (N_4299,N_4106,N_4105);
and U4300 (N_4300,N_4242,N_4289);
and U4301 (N_4301,N_4277,N_4232);
or U4302 (N_4302,N_4203,N_4260);
xor U4303 (N_4303,N_4273,N_4298);
and U4304 (N_4304,N_4264,N_4229);
nand U4305 (N_4305,N_4251,N_4243);
nand U4306 (N_4306,N_4200,N_4255);
and U4307 (N_4307,N_4217,N_4220);
and U4308 (N_4308,N_4223,N_4271);
or U4309 (N_4309,N_4299,N_4250);
or U4310 (N_4310,N_4270,N_4214);
nor U4311 (N_4311,N_4240,N_4288);
nor U4312 (N_4312,N_4235,N_4252);
or U4313 (N_4313,N_4227,N_4230);
or U4314 (N_4314,N_4253,N_4207);
or U4315 (N_4315,N_4258,N_4205);
or U4316 (N_4316,N_4249,N_4286);
nor U4317 (N_4317,N_4237,N_4226);
xor U4318 (N_4318,N_4266,N_4246);
nand U4319 (N_4319,N_4295,N_4211);
nand U4320 (N_4320,N_4228,N_4231);
xor U4321 (N_4321,N_4290,N_4234);
nand U4322 (N_4322,N_4281,N_4291);
nand U4323 (N_4323,N_4265,N_4221);
or U4324 (N_4324,N_4222,N_4218);
or U4325 (N_4325,N_4272,N_4241);
nor U4326 (N_4326,N_4287,N_4276);
or U4327 (N_4327,N_4208,N_4219);
or U4328 (N_4328,N_4268,N_4275);
nor U4329 (N_4329,N_4210,N_4233);
and U4330 (N_4330,N_4274,N_4239);
xor U4331 (N_4331,N_4263,N_4238);
xnor U4332 (N_4332,N_4215,N_4257);
or U4333 (N_4333,N_4278,N_4285);
and U4334 (N_4334,N_4261,N_4296);
xnor U4335 (N_4335,N_4212,N_4225);
or U4336 (N_4336,N_4224,N_4280);
and U4337 (N_4337,N_4256,N_4216);
and U4338 (N_4338,N_4262,N_4294);
nand U4339 (N_4339,N_4244,N_4293);
and U4340 (N_4340,N_4282,N_4247);
nand U4341 (N_4341,N_4297,N_4292);
or U4342 (N_4342,N_4279,N_4213);
nand U4343 (N_4343,N_4209,N_4201);
nor U4344 (N_4344,N_4206,N_4284);
and U4345 (N_4345,N_4204,N_4245);
or U4346 (N_4346,N_4248,N_4254);
nor U4347 (N_4347,N_4236,N_4202);
or U4348 (N_4348,N_4283,N_4259);
nor U4349 (N_4349,N_4267,N_4269);
nor U4350 (N_4350,N_4226,N_4236);
xor U4351 (N_4351,N_4226,N_4207);
nand U4352 (N_4352,N_4232,N_4211);
nand U4353 (N_4353,N_4216,N_4233);
xor U4354 (N_4354,N_4204,N_4282);
or U4355 (N_4355,N_4273,N_4206);
nand U4356 (N_4356,N_4213,N_4206);
nor U4357 (N_4357,N_4202,N_4243);
nor U4358 (N_4358,N_4231,N_4222);
nor U4359 (N_4359,N_4228,N_4256);
xnor U4360 (N_4360,N_4278,N_4226);
and U4361 (N_4361,N_4289,N_4287);
xor U4362 (N_4362,N_4280,N_4299);
xnor U4363 (N_4363,N_4241,N_4237);
nor U4364 (N_4364,N_4248,N_4258);
nand U4365 (N_4365,N_4258,N_4260);
or U4366 (N_4366,N_4203,N_4220);
xor U4367 (N_4367,N_4255,N_4245);
or U4368 (N_4368,N_4223,N_4297);
xnor U4369 (N_4369,N_4215,N_4219);
nor U4370 (N_4370,N_4259,N_4263);
nand U4371 (N_4371,N_4279,N_4295);
xor U4372 (N_4372,N_4272,N_4284);
and U4373 (N_4373,N_4284,N_4224);
nand U4374 (N_4374,N_4257,N_4229);
or U4375 (N_4375,N_4261,N_4205);
or U4376 (N_4376,N_4263,N_4203);
xnor U4377 (N_4377,N_4289,N_4219);
or U4378 (N_4378,N_4260,N_4246);
nor U4379 (N_4379,N_4278,N_4262);
xor U4380 (N_4380,N_4285,N_4245);
or U4381 (N_4381,N_4216,N_4259);
nand U4382 (N_4382,N_4207,N_4236);
nand U4383 (N_4383,N_4271,N_4222);
and U4384 (N_4384,N_4280,N_4234);
nand U4385 (N_4385,N_4287,N_4246);
or U4386 (N_4386,N_4233,N_4299);
and U4387 (N_4387,N_4254,N_4296);
and U4388 (N_4388,N_4236,N_4265);
or U4389 (N_4389,N_4214,N_4212);
xor U4390 (N_4390,N_4213,N_4266);
or U4391 (N_4391,N_4277,N_4225);
nor U4392 (N_4392,N_4219,N_4288);
or U4393 (N_4393,N_4276,N_4218);
nand U4394 (N_4394,N_4215,N_4282);
xnor U4395 (N_4395,N_4231,N_4244);
and U4396 (N_4396,N_4216,N_4205);
xnor U4397 (N_4397,N_4226,N_4290);
nand U4398 (N_4398,N_4217,N_4287);
or U4399 (N_4399,N_4255,N_4269);
or U4400 (N_4400,N_4346,N_4339);
and U4401 (N_4401,N_4374,N_4396);
xnor U4402 (N_4402,N_4334,N_4320);
or U4403 (N_4403,N_4304,N_4364);
xnor U4404 (N_4404,N_4347,N_4380);
nand U4405 (N_4405,N_4350,N_4302);
nor U4406 (N_4406,N_4391,N_4366);
nand U4407 (N_4407,N_4344,N_4317);
nand U4408 (N_4408,N_4316,N_4300);
xor U4409 (N_4409,N_4341,N_4362);
nor U4410 (N_4410,N_4377,N_4324);
or U4411 (N_4411,N_4398,N_4322);
nand U4412 (N_4412,N_4399,N_4338);
xor U4413 (N_4413,N_4389,N_4309);
nand U4414 (N_4414,N_4326,N_4360);
xor U4415 (N_4415,N_4305,N_4359);
nand U4416 (N_4416,N_4306,N_4384);
xor U4417 (N_4417,N_4327,N_4315);
or U4418 (N_4418,N_4336,N_4375);
nand U4419 (N_4419,N_4357,N_4373);
or U4420 (N_4420,N_4307,N_4308);
nor U4421 (N_4421,N_4361,N_4343);
xor U4422 (N_4422,N_4397,N_4369);
nand U4423 (N_4423,N_4332,N_4378);
or U4424 (N_4424,N_4312,N_4355);
nand U4425 (N_4425,N_4382,N_4331);
and U4426 (N_4426,N_4352,N_4386);
or U4427 (N_4427,N_4348,N_4321);
nand U4428 (N_4428,N_4319,N_4314);
and U4429 (N_4429,N_4388,N_4367);
nor U4430 (N_4430,N_4390,N_4381);
or U4431 (N_4431,N_4311,N_4376);
nor U4432 (N_4432,N_4349,N_4353);
or U4433 (N_4433,N_4371,N_4310);
and U4434 (N_4434,N_4313,N_4393);
xnor U4435 (N_4435,N_4323,N_4387);
or U4436 (N_4436,N_4379,N_4368);
nor U4437 (N_4437,N_4351,N_4337);
nand U4438 (N_4438,N_4370,N_4358);
nand U4439 (N_4439,N_4372,N_4363);
nor U4440 (N_4440,N_4328,N_4325);
and U4441 (N_4441,N_4385,N_4342);
or U4442 (N_4442,N_4395,N_4303);
nand U4443 (N_4443,N_4356,N_4345);
or U4444 (N_4444,N_4392,N_4318);
and U4445 (N_4445,N_4301,N_4394);
xnor U4446 (N_4446,N_4335,N_4365);
nand U4447 (N_4447,N_4330,N_4340);
nor U4448 (N_4448,N_4329,N_4333);
xnor U4449 (N_4449,N_4354,N_4383);
xnor U4450 (N_4450,N_4317,N_4398);
or U4451 (N_4451,N_4318,N_4350);
nor U4452 (N_4452,N_4388,N_4331);
and U4453 (N_4453,N_4365,N_4302);
and U4454 (N_4454,N_4303,N_4350);
nor U4455 (N_4455,N_4301,N_4393);
nor U4456 (N_4456,N_4321,N_4334);
nor U4457 (N_4457,N_4351,N_4366);
or U4458 (N_4458,N_4302,N_4362);
or U4459 (N_4459,N_4317,N_4351);
and U4460 (N_4460,N_4360,N_4378);
nor U4461 (N_4461,N_4317,N_4339);
xnor U4462 (N_4462,N_4336,N_4349);
xnor U4463 (N_4463,N_4378,N_4389);
nor U4464 (N_4464,N_4391,N_4393);
xor U4465 (N_4465,N_4390,N_4319);
and U4466 (N_4466,N_4307,N_4320);
or U4467 (N_4467,N_4371,N_4320);
and U4468 (N_4468,N_4379,N_4386);
nor U4469 (N_4469,N_4323,N_4386);
or U4470 (N_4470,N_4346,N_4331);
nand U4471 (N_4471,N_4316,N_4311);
or U4472 (N_4472,N_4388,N_4345);
nor U4473 (N_4473,N_4312,N_4369);
or U4474 (N_4474,N_4372,N_4321);
and U4475 (N_4475,N_4336,N_4343);
or U4476 (N_4476,N_4309,N_4339);
and U4477 (N_4477,N_4357,N_4397);
or U4478 (N_4478,N_4381,N_4315);
nor U4479 (N_4479,N_4397,N_4323);
nor U4480 (N_4480,N_4375,N_4301);
and U4481 (N_4481,N_4332,N_4373);
xor U4482 (N_4482,N_4389,N_4337);
nor U4483 (N_4483,N_4328,N_4357);
and U4484 (N_4484,N_4333,N_4357);
nor U4485 (N_4485,N_4310,N_4382);
xor U4486 (N_4486,N_4328,N_4329);
or U4487 (N_4487,N_4327,N_4321);
and U4488 (N_4488,N_4341,N_4354);
and U4489 (N_4489,N_4311,N_4355);
and U4490 (N_4490,N_4379,N_4304);
nand U4491 (N_4491,N_4338,N_4302);
or U4492 (N_4492,N_4393,N_4352);
nand U4493 (N_4493,N_4339,N_4312);
and U4494 (N_4494,N_4365,N_4333);
xnor U4495 (N_4495,N_4305,N_4371);
or U4496 (N_4496,N_4319,N_4324);
and U4497 (N_4497,N_4320,N_4351);
xor U4498 (N_4498,N_4363,N_4343);
xor U4499 (N_4499,N_4393,N_4339);
nor U4500 (N_4500,N_4438,N_4447);
nand U4501 (N_4501,N_4496,N_4407);
or U4502 (N_4502,N_4463,N_4483);
xnor U4503 (N_4503,N_4430,N_4421);
nor U4504 (N_4504,N_4459,N_4476);
and U4505 (N_4505,N_4498,N_4450);
nand U4506 (N_4506,N_4409,N_4448);
xnor U4507 (N_4507,N_4479,N_4484);
nand U4508 (N_4508,N_4403,N_4420);
nand U4509 (N_4509,N_4470,N_4415);
nor U4510 (N_4510,N_4426,N_4491);
nand U4511 (N_4511,N_4445,N_4406);
nand U4512 (N_4512,N_4472,N_4412);
nand U4513 (N_4513,N_4469,N_4458);
and U4514 (N_4514,N_4480,N_4442);
xor U4515 (N_4515,N_4418,N_4446);
xor U4516 (N_4516,N_4401,N_4486);
xor U4517 (N_4517,N_4489,N_4492);
and U4518 (N_4518,N_4499,N_4465);
or U4519 (N_4519,N_4449,N_4461);
nand U4520 (N_4520,N_4490,N_4423);
nor U4521 (N_4521,N_4404,N_4468);
nor U4522 (N_4522,N_4460,N_4481);
nand U4523 (N_4523,N_4402,N_4466);
nand U4524 (N_4524,N_4437,N_4441);
nand U4525 (N_4525,N_4414,N_4432);
nor U4526 (N_4526,N_4435,N_4413);
xnor U4527 (N_4527,N_4454,N_4425);
and U4528 (N_4528,N_4451,N_4416);
or U4529 (N_4529,N_4429,N_4473);
or U4530 (N_4530,N_4410,N_4422);
or U4531 (N_4531,N_4474,N_4427);
and U4532 (N_4532,N_4443,N_4495);
or U4533 (N_4533,N_4467,N_4436);
or U4534 (N_4534,N_4431,N_4444);
and U4535 (N_4535,N_4417,N_4493);
xor U4536 (N_4536,N_4455,N_4494);
nor U4537 (N_4537,N_4456,N_4433);
or U4538 (N_4538,N_4497,N_4462);
xnor U4539 (N_4539,N_4485,N_4482);
nor U4540 (N_4540,N_4411,N_4419);
nor U4541 (N_4541,N_4453,N_4440);
nand U4542 (N_4542,N_4477,N_4475);
or U4543 (N_4543,N_4471,N_4428);
nand U4544 (N_4544,N_4405,N_4400);
and U4545 (N_4545,N_4452,N_4488);
nor U4546 (N_4546,N_4434,N_4478);
nor U4547 (N_4547,N_4439,N_4457);
or U4548 (N_4548,N_4487,N_4464);
or U4549 (N_4549,N_4424,N_4408);
and U4550 (N_4550,N_4497,N_4417);
and U4551 (N_4551,N_4448,N_4480);
nor U4552 (N_4552,N_4459,N_4485);
xor U4553 (N_4553,N_4418,N_4410);
nor U4554 (N_4554,N_4430,N_4463);
nand U4555 (N_4555,N_4408,N_4401);
and U4556 (N_4556,N_4454,N_4493);
nand U4557 (N_4557,N_4429,N_4476);
and U4558 (N_4558,N_4482,N_4431);
nand U4559 (N_4559,N_4449,N_4488);
nand U4560 (N_4560,N_4458,N_4413);
and U4561 (N_4561,N_4400,N_4404);
xnor U4562 (N_4562,N_4420,N_4415);
nand U4563 (N_4563,N_4439,N_4499);
nand U4564 (N_4564,N_4444,N_4473);
nor U4565 (N_4565,N_4408,N_4426);
nor U4566 (N_4566,N_4448,N_4467);
nor U4567 (N_4567,N_4449,N_4446);
and U4568 (N_4568,N_4418,N_4492);
and U4569 (N_4569,N_4482,N_4494);
or U4570 (N_4570,N_4475,N_4471);
xor U4571 (N_4571,N_4494,N_4489);
or U4572 (N_4572,N_4466,N_4441);
or U4573 (N_4573,N_4431,N_4470);
xor U4574 (N_4574,N_4404,N_4466);
nor U4575 (N_4575,N_4428,N_4467);
or U4576 (N_4576,N_4475,N_4487);
and U4577 (N_4577,N_4484,N_4402);
nor U4578 (N_4578,N_4471,N_4408);
and U4579 (N_4579,N_4401,N_4475);
nor U4580 (N_4580,N_4473,N_4492);
xnor U4581 (N_4581,N_4417,N_4462);
nor U4582 (N_4582,N_4464,N_4495);
xnor U4583 (N_4583,N_4490,N_4447);
nor U4584 (N_4584,N_4422,N_4474);
nand U4585 (N_4585,N_4422,N_4487);
nor U4586 (N_4586,N_4424,N_4403);
xnor U4587 (N_4587,N_4471,N_4485);
and U4588 (N_4588,N_4489,N_4459);
nor U4589 (N_4589,N_4421,N_4422);
and U4590 (N_4590,N_4451,N_4457);
nand U4591 (N_4591,N_4418,N_4400);
and U4592 (N_4592,N_4419,N_4425);
and U4593 (N_4593,N_4419,N_4446);
nor U4594 (N_4594,N_4428,N_4483);
xor U4595 (N_4595,N_4481,N_4492);
or U4596 (N_4596,N_4451,N_4488);
nand U4597 (N_4597,N_4461,N_4457);
or U4598 (N_4598,N_4457,N_4449);
nand U4599 (N_4599,N_4431,N_4490);
or U4600 (N_4600,N_4561,N_4564);
or U4601 (N_4601,N_4585,N_4568);
and U4602 (N_4602,N_4594,N_4572);
and U4603 (N_4603,N_4586,N_4595);
nand U4604 (N_4604,N_4549,N_4559);
nand U4605 (N_4605,N_4541,N_4562);
xnor U4606 (N_4606,N_4502,N_4516);
nand U4607 (N_4607,N_4552,N_4542);
and U4608 (N_4608,N_4548,N_4500);
or U4609 (N_4609,N_4599,N_4588);
nor U4610 (N_4610,N_4579,N_4535);
or U4611 (N_4611,N_4581,N_4574);
and U4612 (N_4612,N_4577,N_4587);
nand U4613 (N_4613,N_4512,N_4523);
or U4614 (N_4614,N_4593,N_4554);
or U4615 (N_4615,N_4551,N_4598);
xor U4616 (N_4616,N_4547,N_4524);
nor U4617 (N_4617,N_4550,N_4544);
or U4618 (N_4618,N_4575,N_4576);
or U4619 (N_4619,N_4530,N_4515);
and U4620 (N_4620,N_4528,N_4596);
or U4621 (N_4621,N_4545,N_4506);
nor U4622 (N_4622,N_4563,N_4558);
nor U4623 (N_4623,N_4521,N_4527);
or U4624 (N_4624,N_4538,N_4517);
nand U4625 (N_4625,N_4583,N_4536);
nand U4626 (N_4626,N_4522,N_4589);
or U4627 (N_4627,N_4509,N_4519);
and U4628 (N_4628,N_4501,N_4511);
xnor U4629 (N_4629,N_4533,N_4580);
or U4630 (N_4630,N_4510,N_4571);
nor U4631 (N_4631,N_4592,N_4513);
and U4632 (N_4632,N_4584,N_4520);
and U4633 (N_4633,N_4505,N_4507);
nor U4634 (N_4634,N_4566,N_4518);
nor U4635 (N_4635,N_4567,N_4553);
nand U4636 (N_4636,N_4504,N_4540);
and U4637 (N_4637,N_4534,N_4597);
nand U4638 (N_4638,N_4508,N_4573);
and U4639 (N_4639,N_4532,N_4531);
nor U4640 (N_4640,N_4529,N_4543);
xor U4641 (N_4641,N_4556,N_4539);
nor U4642 (N_4642,N_4569,N_4557);
xnor U4643 (N_4643,N_4555,N_4526);
xor U4644 (N_4644,N_4560,N_4570);
and U4645 (N_4645,N_4537,N_4514);
or U4646 (N_4646,N_4546,N_4590);
or U4647 (N_4647,N_4591,N_4582);
and U4648 (N_4648,N_4565,N_4503);
nand U4649 (N_4649,N_4525,N_4578);
or U4650 (N_4650,N_4558,N_4597);
nand U4651 (N_4651,N_4524,N_4539);
nand U4652 (N_4652,N_4567,N_4541);
nand U4653 (N_4653,N_4510,N_4548);
nand U4654 (N_4654,N_4554,N_4592);
xnor U4655 (N_4655,N_4587,N_4596);
and U4656 (N_4656,N_4569,N_4505);
nand U4657 (N_4657,N_4506,N_4543);
and U4658 (N_4658,N_4521,N_4524);
or U4659 (N_4659,N_4506,N_4550);
and U4660 (N_4660,N_4534,N_4566);
xor U4661 (N_4661,N_4549,N_4535);
nor U4662 (N_4662,N_4574,N_4562);
nand U4663 (N_4663,N_4551,N_4526);
xnor U4664 (N_4664,N_4593,N_4574);
nand U4665 (N_4665,N_4526,N_4520);
nand U4666 (N_4666,N_4525,N_4572);
or U4667 (N_4667,N_4558,N_4524);
xor U4668 (N_4668,N_4560,N_4586);
xor U4669 (N_4669,N_4586,N_4537);
nand U4670 (N_4670,N_4512,N_4521);
and U4671 (N_4671,N_4558,N_4507);
xnor U4672 (N_4672,N_4592,N_4541);
and U4673 (N_4673,N_4556,N_4575);
nand U4674 (N_4674,N_4560,N_4531);
and U4675 (N_4675,N_4527,N_4552);
and U4676 (N_4676,N_4558,N_4542);
nor U4677 (N_4677,N_4518,N_4531);
and U4678 (N_4678,N_4506,N_4595);
nand U4679 (N_4679,N_4513,N_4575);
or U4680 (N_4680,N_4534,N_4538);
nand U4681 (N_4681,N_4575,N_4509);
xor U4682 (N_4682,N_4540,N_4557);
nand U4683 (N_4683,N_4536,N_4543);
and U4684 (N_4684,N_4534,N_4530);
nand U4685 (N_4685,N_4586,N_4541);
or U4686 (N_4686,N_4570,N_4526);
or U4687 (N_4687,N_4539,N_4531);
and U4688 (N_4688,N_4546,N_4520);
xnor U4689 (N_4689,N_4584,N_4546);
nor U4690 (N_4690,N_4596,N_4506);
nor U4691 (N_4691,N_4593,N_4584);
or U4692 (N_4692,N_4564,N_4596);
or U4693 (N_4693,N_4582,N_4519);
nor U4694 (N_4694,N_4555,N_4508);
xnor U4695 (N_4695,N_4520,N_4514);
or U4696 (N_4696,N_4567,N_4562);
nand U4697 (N_4697,N_4551,N_4544);
and U4698 (N_4698,N_4506,N_4508);
nor U4699 (N_4699,N_4568,N_4594);
and U4700 (N_4700,N_4679,N_4665);
or U4701 (N_4701,N_4618,N_4637);
and U4702 (N_4702,N_4688,N_4634);
and U4703 (N_4703,N_4643,N_4677);
and U4704 (N_4704,N_4671,N_4656);
and U4705 (N_4705,N_4696,N_4623);
nand U4706 (N_4706,N_4640,N_4672);
nand U4707 (N_4707,N_4645,N_4608);
xnor U4708 (N_4708,N_4628,N_4600);
or U4709 (N_4709,N_4668,N_4693);
nor U4710 (N_4710,N_4605,N_4658);
and U4711 (N_4711,N_4607,N_4622);
nor U4712 (N_4712,N_4675,N_4633);
or U4713 (N_4713,N_4692,N_4619);
xor U4714 (N_4714,N_4651,N_4683);
and U4715 (N_4715,N_4631,N_4630);
nor U4716 (N_4716,N_4690,N_4616);
xor U4717 (N_4717,N_4652,N_4662);
nand U4718 (N_4718,N_4655,N_4614);
or U4719 (N_4719,N_4602,N_4621);
or U4720 (N_4720,N_4601,N_4609);
or U4721 (N_4721,N_4627,N_4629);
or U4722 (N_4722,N_4639,N_4654);
nand U4723 (N_4723,N_4620,N_4689);
xor U4724 (N_4724,N_4680,N_4625);
or U4725 (N_4725,N_4660,N_4657);
and U4726 (N_4726,N_4681,N_4642);
or U4727 (N_4727,N_4698,N_4699);
xnor U4728 (N_4728,N_4666,N_4626);
and U4729 (N_4729,N_4676,N_4669);
xor U4730 (N_4730,N_4685,N_4649);
and U4731 (N_4731,N_4653,N_4678);
xnor U4732 (N_4732,N_4617,N_4673);
nand U4733 (N_4733,N_4659,N_4687);
and U4734 (N_4734,N_4686,N_4684);
or U4735 (N_4735,N_4691,N_4638);
nand U4736 (N_4736,N_4606,N_4644);
xor U4737 (N_4737,N_4682,N_4646);
and U4738 (N_4738,N_4615,N_4670);
and U4739 (N_4739,N_4661,N_4650);
xor U4740 (N_4740,N_4636,N_4648);
nor U4741 (N_4741,N_4603,N_4635);
nand U4742 (N_4742,N_4632,N_4604);
and U4743 (N_4743,N_4647,N_4613);
nor U4744 (N_4744,N_4610,N_4697);
xor U4745 (N_4745,N_4695,N_4611);
xor U4746 (N_4746,N_4663,N_4694);
or U4747 (N_4747,N_4612,N_4641);
nor U4748 (N_4748,N_4624,N_4674);
nor U4749 (N_4749,N_4667,N_4664);
nand U4750 (N_4750,N_4649,N_4639);
xnor U4751 (N_4751,N_4632,N_4602);
xnor U4752 (N_4752,N_4610,N_4603);
xnor U4753 (N_4753,N_4674,N_4617);
xnor U4754 (N_4754,N_4640,N_4654);
nor U4755 (N_4755,N_4632,N_4608);
or U4756 (N_4756,N_4673,N_4600);
nand U4757 (N_4757,N_4697,N_4673);
or U4758 (N_4758,N_4627,N_4658);
nand U4759 (N_4759,N_4699,N_4666);
xor U4760 (N_4760,N_4673,N_4615);
and U4761 (N_4761,N_4618,N_4638);
nor U4762 (N_4762,N_4621,N_4624);
and U4763 (N_4763,N_4629,N_4611);
or U4764 (N_4764,N_4697,N_4601);
xor U4765 (N_4765,N_4657,N_4651);
nor U4766 (N_4766,N_4634,N_4655);
nand U4767 (N_4767,N_4680,N_4636);
or U4768 (N_4768,N_4624,N_4698);
or U4769 (N_4769,N_4697,N_4660);
nor U4770 (N_4770,N_4654,N_4665);
or U4771 (N_4771,N_4683,N_4647);
nand U4772 (N_4772,N_4649,N_4684);
or U4773 (N_4773,N_4660,N_4612);
or U4774 (N_4774,N_4617,N_4622);
and U4775 (N_4775,N_4634,N_4696);
nand U4776 (N_4776,N_4663,N_4646);
and U4777 (N_4777,N_4690,N_4681);
or U4778 (N_4778,N_4683,N_4678);
nor U4779 (N_4779,N_4687,N_4617);
or U4780 (N_4780,N_4688,N_4626);
nand U4781 (N_4781,N_4682,N_4670);
and U4782 (N_4782,N_4603,N_4683);
and U4783 (N_4783,N_4661,N_4607);
nor U4784 (N_4784,N_4618,N_4687);
xor U4785 (N_4785,N_4625,N_4685);
and U4786 (N_4786,N_4649,N_4636);
xnor U4787 (N_4787,N_4645,N_4624);
nand U4788 (N_4788,N_4693,N_4652);
or U4789 (N_4789,N_4638,N_4610);
nand U4790 (N_4790,N_4604,N_4624);
or U4791 (N_4791,N_4662,N_4658);
nand U4792 (N_4792,N_4619,N_4624);
or U4793 (N_4793,N_4603,N_4646);
and U4794 (N_4794,N_4679,N_4634);
or U4795 (N_4795,N_4675,N_4640);
and U4796 (N_4796,N_4621,N_4625);
or U4797 (N_4797,N_4622,N_4633);
and U4798 (N_4798,N_4681,N_4618);
xnor U4799 (N_4799,N_4603,N_4609);
and U4800 (N_4800,N_4748,N_4701);
and U4801 (N_4801,N_4706,N_4789);
xor U4802 (N_4802,N_4778,N_4720);
xnor U4803 (N_4803,N_4712,N_4747);
and U4804 (N_4804,N_4734,N_4793);
and U4805 (N_4805,N_4752,N_4770);
nand U4806 (N_4806,N_4717,N_4791);
xnor U4807 (N_4807,N_4786,N_4722);
nor U4808 (N_4808,N_4728,N_4733);
or U4809 (N_4809,N_4702,N_4783);
nand U4810 (N_4810,N_4709,N_4779);
and U4811 (N_4811,N_4755,N_4719);
or U4812 (N_4812,N_4716,N_4727);
and U4813 (N_4813,N_4724,N_4740);
xor U4814 (N_4814,N_4797,N_4718);
and U4815 (N_4815,N_4767,N_4781);
nand U4816 (N_4816,N_4758,N_4761);
xnor U4817 (N_4817,N_4730,N_4790);
nand U4818 (N_4818,N_4775,N_4798);
or U4819 (N_4819,N_4773,N_4787);
nand U4820 (N_4820,N_4723,N_4796);
nand U4821 (N_4821,N_4714,N_4750);
nor U4822 (N_4822,N_4785,N_4782);
nand U4823 (N_4823,N_4737,N_4799);
and U4824 (N_4824,N_4765,N_4772);
and U4825 (N_4825,N_4721,N_4792);
or U4826 (N_4826,N_4711,N_4700);
or U4827 (N_4827,N_4713,N_4731);
and U4828 (N_4828,N_4774,N_4703);
nor U4829 (N_4829,N_4795,N_4746);
nor U4830 (N_4830,N_4766,N_4777);
nand U4831 (N_4831,N_4756,N_4739);
and U4832 (N_4832,N_4736,N_4749);
xnor U4833 (N_4833,N_4704,N_4751);
xor U4834 (N_4834,N_4732,N_4745);
and U4835 (N_4835,N_4768,N_4763);
or U4836 (N_4836,N_4776,N_4764);
nor U4837 (N_4837,N_4753,N_4794);
and U4838 (N_4838,N_4726,N_4735);
or U4839 (N_4839,N_4741,N_4759);
or U4840 (N_4840,N_4744,N_4710);
nor U4841 (N_4841,N_4780,N_4784);
nor U4842 (N_4842,N_4742,N_4754);
xor U4843 (N_4843,N_4769,N_4771);
and U4844 (N_4844,N_4715,N_4743);
or U4845 (N_4845,N_4725,N_4707);
nand U4846 (N_4846,N_4762,N_4788);
nor U4847 (N_4847,N_4708,N_4729);
and U4848 (N_4848,N_4705,N_4760);
and U4849 (N_4849,N_4738,N_4757);
and U4850 (N_4850,N_4740,N_4738);
nor U4851 (N_4851,N_4760,N_4741);
nand U4852 (N_4852,N_4714,N_4791);
nor U4853 (N_4853,N_4774,N_4719);
or U4854 (N_4854,N_4778,N_4715);
and U4855 (N_4855,N_4752,N_4799);
nand U4856 (N_4856,N_4749,N_4765);
xnor U4857 (N_4857,N_4773,N_4714);
xor U4858 (N_4858,N_4742,N_4783);
or U4859 (N_4859,N_4796,N_4777);
nand U4860 (N_4860,N_4790,N_4788);
or U4861 (N_4861,N_4753,N_4725);
or U4862 (N_4862,N_4756,N_4762);
nor U4863 (N_4863,N_4750,N_4742);
nor U4864 (N_4864,N_4748,N_4704);
xor U4865 (N_4865,N_4731,N_4761);
xor U4866 (N_4866,N_4764,N_4773);
or U4867 (N_4867,N_4739,N_4764);
or U4868 (N_4868,N_4746,N_4747);
xnor U4869 (N_4869,N_4766,N_4743);
nor U4870 (N_4870,N_4708,N_4782);
or U4871 (N_4871,N_4794,N_4707);
and U4872 (N_4872,N_4752,N_4791);
nor U4873 (N_4873,N_4794,N_4748);
and U4874 (N_4874,N_4761,N_4788);
and U4875 (N_4875,N_4742,N_4734);
nand U4876 (N_4876,N_4758,N_4781);
nor U4877 (N_4877,N_4761,N_4767);
nor U4878 (N_4878,N_4772,N_4702);
nand U4879 (N_4879,N_4778,N_4759);
or U4880 (N_4880,N_4791,N_4740);
nor U4881 (N_4881,N_4751,N_4735);
or U4882 (N_4882,N_4767,N_4703);
and U4883 (N_4883,N_4786,N_4742);
nor U4884 (N_4884,N_4716,N_4750);
or U4885 (N_4885,N_4797,N_4769);
nand U4886 (N_4886,N_4765,N_4766);
nand U4887 (N_4887,N_4766,N_4726);
and U4888 (N_4888,N_4732,N_4759);
xnor U4889 (N_4889,N_4786,N_4762);
nor U4890 (N_4890,N_4772,N_4705);
nor U4891 (N_4891,N_4762,N_4715);
or U4892 (N_4892,N_4782,N_4759);
and U4893 (N_4893,N_4792,N_4715);
or U4894 (N_4894,N_4794,N_4790);
xor U4895 (N_4895,N_4777,N_4788);
nand U4896 (N_4896,N_4769,N_4781);
nor U4897 (N_4897,N_4772,N_4770);
xor U4898 (N_4898,N_4756,N_4731);
nor U4899 (N_4899,N_4761,N_4700);
nand U4900 (N_4900,N_4867,N_4821);
nand U4901 (N_4901,N_4882,N_4802);
or U4902 (N_4902,N_4805,N_4854);
nor U4903 (N_4903,N_4873,N_4839);
xor U4904 (N_4904,N_4857,N_4816);
nor U4905 (N_4905,N_4851,N_4888);
and U4906 (N_4906,N_4860,N_4846);
and U4907 (N_4907,N_4875,N_4809);
nor U4908 (N_4908,N_4861,N_4810);
nand U4909 (N_4909,N_4841,N_4830);
xnor U4910 (N_4910,N_4817,N_4832);
nor U4911 (N_4911,N_4894,N_4835);
nand U4912 (N_4912,N_4868,N_4881);
and U4913 (N_4913,N_4878,N_4853);
nand U4914 (N_4914,N_4865,N_4814);
nor U4915 (N_4915,N_4806,N_4897);
or U4916 (N_4916,N_4826,N_4880);
and U4917 (N_4917,N_4859,N_4812);
nor U4918 (N_4918,N_4811,N_4847);
nand U4919 (N_4919,N_4808,N_4819);
nor U4920 (N_4920,N_4845,N_4801);
nand U4921 (N_4921,N_4813,N_4884);
xor U4922 (N_4922,N_4879,N_4824);
and U4923 (N_4923,N_4872,N_4886);
xnor U4924 (N_4924,N_4843,N_4823);
and U4925 (N_4925,N_4893,N_4895);
or U4926 (N_4926,N_4833,N_4883);
xnor U4927 (N_4927,N_4822,N_4862);
nand U4928 (N_4928,N_4838,N_4874);
or U4929 (N_4929,N_4891,N_4842);
xnor U4930 (N_4930,N_4890,N_4800);
nand U4931 (N_4931,N_4887,N_4855);
xor U4932 (N_4932,N_4829,N_4836);
nand U4933 (N_4933,N_4892,N_4863);
and U4934 (N_4934,N_4896,N_4899);
nor U4935 (N_4935,N_4831,N_4885);
nand U4936 (N_4936,N_4828,N_4852);
xor U4937 (N_4937,N_4825,N_4864);
nor U4938 (N_4938,N_4850,N_4844);
and U4939 (N_4939,N_4804,N_4889);
and U4940 (N_4940,N_4820,N_4803);
and U4941 (N_4941,N_4866,N_4834);
or U4942 (N_4942,N_4871,N_4877);
xnor U4943 (N_4943,N_4869,N_4898);
or U4944 (N_4944,N_4856,N_4827);
nor U4945 (N_4945,N_4815,N_4849);
xnor U4946 (N_4946,N_4858,N_4837);
xor U4947 (N_4947,N_4840,N_4848);
nor U4948 (N_4948,N_4818,N_4870);
nor U4949 (N_4949,N_4807,N_4876);
nor U4950 (N_4950,N_4892,N_4857);
xnor U4951 (N_4951,N_4824,N_4821);
or U4952 (N_4952,N_4824,N_4855);
or U4953 (N_4953,N_4822,N_4852);
and U4954 (N_4954,N_4817,N_4855);
or U4955 (N_4955,N_4844,N_4812);
nand U4956 (N_4956,N_4854,N_4860);
xnor U4957 (N_4957,N_4859,N_4838);
xor U4958 (N_4958,N_4875,N_4842);
xnor U4959 (N_4959,N_4838,N_4886);
xor U4960 (N_4960,N_4801,N_4809);
or U4961 (N_4961,N_4807,N_4800);
nand U4962 (N_4962,N_4827,N_4874);
or U4963 (N_4963,N_4849,N_4850);
or U4964 (N_4964,N_4816,N_4850);
or U4965 (N_4965,N_4876,N_4830);
nand U4966 (N_4966,N_4815,N_4837);
and U4967 (N_4967,N_4833,N_4849);
nand U4968 (N_4968,N_4809,N_4882);
and U4969 (N_4969,N_4830,N_4829);
nand U4970 (N_4970,N_4857,N_4843);
or U4971 (N_4971,N_4864,N_4815);
and U4972 (N_4972,N_4892,N_4825);
nand U4973 (N_4973,N_4808,N_4848);
xnor U4974 (N_4974,N_4813,N_4893);
nor U4975 (N_4975,N_4809,N_4860);
and U4976 (N_4976,N_4871,N_4804);
and U4977 (N_4977,N_4884,N_4843);
xor U4978 (N_4978,N_4824,N_4853);
nor U4979 (N_4979,N_4882,N_4866);
nor U4980 (N_4980,N_4845,N_4804);
and U4981 (N_4981,N_4885,N_4816);
nand U4982 (N_4982,N_4853,N_4889);
or U4983 (N_4983,N_4814,N_4897);
xor U4984 (N_4984,N_4856,N_4821);
and U4985 (N_4985,N_4880,N_4894);
and U4986 (N_4986,N_4848,N_4825);
nand U4987 (N_4987,N_4899,N_4874);
nand U4988 (N_4988,N_4820,N_4860);
xor U4989 (N_4989,N_4863,N_4803);
and U4990 (N_4990,N_4831,N_4887);
xnor U4991 (N_4991,N_4841,N_4804);
and U4992 (N_4992,N_4822,N_4872);
xnor U4993 (N_4993,N_4840,N_4895);
and U4994 (N_4994,N_4835,N_4823);
or U4995 (N_4995,N_4861,N_4885);
or U4996 (N_4996,N_4815,N_4816);
or U4997 (N_4997,N_4866,N_4805);
or U4998 (N_4998,N_4838,N_4801);
and U4999 (N_4999,N_4863,N_4842);
xnor U5000 (N_5000,N_4961,N_4990);
nand U5001 (N_5001,N_4991,N_4916);
or U5002 (N_5002,N_4949,N_4966);
or U5003 (N_5003,N_4973,N_4931);
nor U5004 (N_5004,N_4935,N_4950);
xor U5005 (N_5005,N_4929,N_4946);
and U5006 (N_5006,N_4902,N_4928);
or U5007 (N_5007,N_4923,N_4945);
nand U5008 (N_5008,N_4909,N_4942);
nand U5009 (N_5009,N_4925,N_4954);
nand U5010 (N_5010,N_4940,N_4926);
or U5011 (N_5011,N_4974,N_4911);
nand U5012 (N_5012,N_4962,N_4972);
and U5013 (N_5013,N_4984,N_4971);
xor U5014 (N_5014,N_4913,N_4921);
and U5015 (N_5015,N_4993,N_4968);
nor U5016 (N_5016,N_4953,N_4917);
xnor U5017 (N_5017,N_4934,N_4979);
nor U5018 (N_5018,N_4977,N_4936);
nor U5019 (N_5019,N_4907,N_4918);
nor U5020 (N_5020,N_4914,N_4969);
or U5021 (N_5021,N_4952,N_4919);
nor U5022 (N_5022,N_4956,N_4905);
nor U5023 (N_5023,N_4999,N_4983);
xnor U5024 (N_5024,N_4965,N_4951);
or U5025 (N_5025,N_4967,N_4985);
and U5026 (N_5026,N_4975,N_4932);
nor U5027 (N_5027,N_4948,N_4908);
and U5028 (N_5028,N_4900,N_4998);
nor U5029 (N_5029,N_4995,N_4904);
or U5030 (N_5030,N_4903,N_4912);
nor U5031 (N_5031,N_4997,N_4959);
nand U5032 (N_5032,N_4982,N_4944);
xnor U5033 (N_5033,N_4922,N_4976);
or U5034 (N_5034,N_4980,N_4930);
xor U5035 (N_5035,N_4915,N_4978);
or U5036 (N_5036,N_4964,N_4988);
nor U5037 (N_5037,N_4992,N_4955);
or U5038 (N_5038,N_4924,N_4958);
or U5039 (N_5039,N_4957,N_4963);
nand U5040 (N_5040,N_4994,N_4960);
nor U5041 (N_5041,N_4989,N_4939);
xnor U5042 (N_5042,N_4920,N_4947);
nor U5043 (N_5043,N_4937,N_4938);
and U5044 (N_5044,N_4943,N_4927);
and U5045 (N_5045,N_4910,N_4987);
and U5046 (N_5046,N_4901,N_4970);
nand U5047 (N_5047,N_4933,N_4986);
and U5048 (N_5048,N_4941,N_4906);
and U5049 (N_5049,N_4996,N_4981);
or U5050 (N_5050,N_4996,N_4924);
nor U5051 (N_5051,N_4911,N_4917);
or U5052 (N_5052,N_4944,N_4956);
xor U5053 (N_5053,N_4998,N_4941);
and U5054 (N_5054,N_4925,N_4984);
nor U5055 (N_5055,N_4932,N_4908);
nor U5056 (N_5056,N_4998,N_4907);
or U5057 (N_5057,N_4915,N_4986);
xnor U5058 (N_5058,N_4921,N_4907);
or U5059 (N_5059,N_4990,N_4960);
nor U5060 (N_5060,N_4966,N_4970);
nor U5061 (N_5061,N_4962,N_4994);
and U5062 (N_5062,N_4924,N_4915);
or U5063 (N_5063,N_4980,N_4940);
xor U5064 (N_5064,N_4926,N_4917);
nand U5065 (N_5065,N_4987,N_4977);
xnor U5066 (N_5066,N_4928,N_4916);
and U5067 (N_5067,N_4962,N_4907);
or U5068 (N_5068,N_4965,N_4919);
and U5069 (N_5069,N_4949,N_4953);
or U5070 (N_5070,N_4903,N_4952);
nor U5071 (N_5071,N_4991,N_4983);
and U5072 (N_5072,N_4906,N_4904);
nand U5073 (N_5073,N_4986,N_4973);
and U5074 (N_5074,N_4945,N_4909);
xnor U5075 (N_5075,N_4978,N_4941);
or U5076 (N_5076,N_4975,N_4961);
and U5077 (N_5077,N_4943,N_4987);
and U5078 (N_5078,N_4947,N_4939);
or U5079 (N_5079,N_4992,N_4917);
and U5080 (N_5080,N_4957,N_4987);
nor U5081 (N_5081,N_4976,N_4902);
nor U5082 (N_5082,N_4910,N_4996);
nand U5083 (N_5083,N_4901,N_4983);
or U5084 (N_5084,N_4965,N_4912);
nand U5085 (N_5085,N_4952,N_4943);
xnor U5086 (N_5086,N_4946,N_4911);
or U5087 (N_5087,N_4917,N_4907);
and U5088 (N_5088,N_4994,N_4958);
xnor U5089 (N_5089,N_4914,N_4976);
nor U5090 (N_5090,N_4998,N_4935);
and U5091 (N_5091,N_4986,N_4945);
nand U5092 (N_5092,N_4915,N_4947);
xor U5093 (N_5093,N_4997,N_4922);
and U5094 (N_5094,N_4983,N_4919);
and U5095 (N_5095,N_4976,N_4905);
and U5096 (N_5096,N_4900,N_4972);
or U5097 (N_5097,N_4901,N_4979);
nand U5098 (N_5098,N_4959,N_4943);
nor U5099 (N_5099,N_4984,N_4926);
or U5100 (N_5100,N_5020,N_5075);
nand U5101 (N_5101,N_5053,N_5081);
and U5102 (N_5102,N_5001,N_5062);
nand U5103 (N_5103,N_5054,N_5017);
or U5104 (N_5104,N_5091,N_5027);
nor U5105 (N_5105,N_5096,N_5066);
xnor U5106 (N_5106,N_5069,N_5049);
and U5107 (N_5107,N_5064,N_5013);
nor U5108 (N_5108,N_5021,N_5014);
or U5109 (N_5109,N_5037,N_5070);
xor U5110 (N_5110,N_5047,N_5057);
nand U5111 (N_5111,N_5028,N_5098);
nand U5112 (N_5112,N_5026,N_5042);
and U5113 (N_5113,N_5085,N_5055);
xor U5114 (N_5114,N_5073,N_5024);
nor U5115 (N_5115,N_5031,N_5063);
and U5116 (N_5116,N_5032,N_5079);
or U5117 (N_5117,N_5025,N_5061);
nor U5118 (N_5118,N_5059,N_5009);
xnor U5119 (N_5119,N_5071,N_5043);
nor U5120 (N_5120,N_5097,N_5086);
and U5121 (N_5121,N_5019,N_5030);
and U5122 (N_5122,N_5000,N_5094);
nor U5123 (N_5123,N_5093,N_5050);
xnor U5124 (N_5124,N_5015,N_5029);
nand U5125 (N_5125,N_5058,N_5056);
and U5126 (N_5126,N_5078,N_5041);
xnor U5127 (N_5127,N_5035,N_5065);
xnor U5128 (N_5128,N_5003,N_5068);
and U5129 (N_5129,N_5005,N_5051);
xor U5130 (N_5130,N_5004,N_5090);
xnor U5131 (N_5131,N_5006,N_5052);
or U5132 (N_5132,N_5040,N_5011);
xnor U5133 (N_5133,N_5023,N_5036);
or U5134 (N_5134,N_5088,N_5099);
nand U5135 (N_5135,N_5089,N_5002);
and U5136 (N_5136,N_5045,N_5072);
or U5137 (N_5137,N_5048,N_5087);
xor U5138 (N_5138,N_5033,N_5076);
and U5139 (N_5139,N_5092,N_5044);
xor U5140 (N_5140,N_5082,N_5080);
nand U5141 (N_5141,N_5060,N_5038);
or U5142 (N_5142,N_5022,N_5008);
xnor U5143 (N_5143,N_5007,N_5039);
nand U5144 (N_5144,N_5077,N_5083);
or U5145 (N_5145,N_5046,N_5016);
or U5146 (N_5146,N_5084,N_5067);
nor U5147 (N_5147,N_5074,N_5012);
and U5148 (N_5148,N_5095,N_5018);
or U5149 (N_5149,N_5010,N_5034);
nand U5150 (N_5150,N_5043,N_5066);
and U5151 (N_5151,N_5009,N_5074);
nor U5152 (N_5152,N_5020,N_5049);
and U5153 (N_5153,N_5077,N_5072);
or U5154 (N_5154,N_5043,N_5070);
nand U5155 (N_5155,N_5033,N_5016);
and U5156 (N_5156,N_5014,N_5098);
nand U5157 (N_5157,N_5024,N_5049);
nor U5158 (N_5158,N_5058,N_5051);
nor U5159 (N_5159,N_5045,N_5092);
xor U5160 (N_5160,N_5012,N_5035);
nor U5161 (N_5161,N_5037,N_5060);
or U5162 (N_5162,N_5084,N_5030);
and U5163 (N_5163,N_5078,N_5021);
and U5164 (N_5164,N_5068,N_5026);
nor U5165 (N_5165,N_5008,N_5093);
nand U5166 (N_5166,N_5011,N_5002);
and U5167 (N_5167,N_5000,N_5084);
nand U5168 (N_5168,N_5050,N_5006);
nand U5169 (N_5169,N_5031,N_5064);
or U5170 (N_5170,N_5039,N_5022);
nor U5171 (N_5171,N_5075,N_5086);
nor U5172 (N_5172,N_5072,N_5046);
nand U5173 (N_5173,N_5085,N_5030);
nand U5174 (N_5174,N_5029,N_5043);
xor U5175 (N_5175,N_5063,N_5098);
nor U5176 (N_5176,N_5012,N_5026);
nor U5177 (N_5177,N_5028,N_5072);
nand U5178 (N_5178,N_5019,N_5017);
and U5179 (N_5179,N_5024,N_5085);
or U5180 (N_5180,N_5064,N_5001);
nor U5181 (N_5181,N_5062,N_5045);
xnor U5182 (N_5182,N_5081,N_5025);
nand U5183 (N_5183,N_5035,N_5017);
nand U5184 (N_5184,N_5053,N_5068);
or U5185 (N_5185,N_5034,N_5056);
xor U5186 (N_5186,N_5039,N_5086);
or U5187 (N_5187,N_5008,N_5057);
or U5188 (N_5188,N_5088,N_5075);
nor U5189 (N_5189,N_5016,N_5018);
and U5190 (N_5190,N_5015,N_5049);
or U5191 (N_5191,N_5008,N_5074);
xnor U5192 (N_5192,N_5014,N_5058);
nand U5193 (N_5193,N_5081,N_5065);
xor U5194 (N_5194,N_5095,N_5008);
and U5195 (N_5195,N_5011,N_5067);
nor U5196 (N_5196,N_5000,N_5070);
or U5197 (N_5197,N_5051,N_5047);
nand U5198 (N_5198,N_5082,N_5025);
and U5199 (N_5199,N_5067,N_5074);
nand U5200 (N_5200,N_5176,N_5124);
xor U5201 (N_5201,N_5177,N_5130);
or U5202 (N_5202,N_5114,N_5189);
and U5203 (N_5203,N_5117,N_5141);
xor U5204 (N_5204,N_5153,N_5138);
or U5205 (N_5205,N_5158,N_5162);
or U5206 (N_5206,N_5109,N_5103);
nand U5207 (N_5207,N_5188,N_5128);
and U5208 (N_5208,N_5101,N_5159);
or U5209 (N_5209,N_5145,N_5132);
nor U5210 (N_5210,N_5156,N_5104);
nor U5211 (N_5211,N_5161,N_5102);
xnor U5212 (N_5212,N_5186,N_5160);
nor U5213 (N_5213,N_5123,N_5185);
xnor U5214 (N_5214,N_5142,N_5164);
nor U5215 (N_5215,N_5173,N_5137);
xnor U5216 (N_5216,N_5171,N_5167);
and U5217 (N_5217,N_5144,N_5199);
and U5218 (N_5218,N_5155,N_5193);
or U5219 (N_5219,N_5146,N_5182);
xnor U5220 (N_5220,N_5113,N_5190);
nor U5221 (N_5221,N_5163,N_5127);
or U5222 (N_5222,N_5174,N_5118);
and U5223 (N_5223,N_5131,N_5154);
xnor U5224 (N_5224,N_5181,N_5116);
xnor U5225 (N_5225,N_5122,N_5194);
nand U5226 (N_5226,N_5150,N_5121);
nand U5227 (N_5227,N_5106,N_5115);
or U5228 (N_5228,N_5149,N_5126);
and U5229 (N_5229,N_5168,N_5129);
nand U5230 (N_5230,N_5107,N_5184);
nor U5231 (N_5231,N_5125,N_5192);
nor U5232 (N_5232,N_5178,N_5134);
or U5233 (N_5233,N_5136,N_5183);
nand U5234 (N_5234,N_5180,N_5147);
xnor U5235 (N_5235,N_5179,N_5170);
nand U5236 (N_5236,N_5139,N_5108);
xnor U5237 (N_5237,N_5135,N_5187);
nand U5238 (N_5238,N_5143,N_5169);
or U5239 (N_5239,N_5191,N_5110);
nand U5240 (N_5240,N_5157,N_5140);
nand U5241 (N_5241,N_5196,N_5148);
xnor U5242 (N_5242,N_5151,N_5166);
or U5243 (N_5243,N_5198,N_5112);
and U5244 (N_5244,N_5172,N_5111);
nand U5245 (N_5245,N_5105,N_5119);
or U5246 (N_5246,N_5165,N_5152);
nor U5247 (N_5247,N_5175,N_5100);
or U5248 (N_5248,N_5133,N_5120);
or U5249 (N_5249,N_5195,N_5197);
nand U5250 (N_5250,N_5188,N_5123);
or U5251 (N_5251,N_5144,N_5102);
nor U5252 (N_5252,N_5186,N_5106);
nand U5253 (N_5253,N_5123,N_5149);
xor U5254 (N_5254,N_5148,N_5189);
xnor U5255 (N_5255,N_5181,N_5173);
nor U5256 (N_5256,N_5141,N_5154);
nand U5257 (N_5257,N_5143,N_5122);
nor U5258 (N_5258,N_5172,N_5157);
nor U5259 (N_5259,N_5103,N_5114);
or U5260 (N_5260,N_5147,N_5159);
or U5261 (N_5261,N_5123,N_5127);
and U5262 (N_5262,N_5132,N_5144);
nand U5263 (N_5263,N_5198,N_5185);
xor U5264 (N_5264,N_5144,N_5160);
nor U5265 (N_5265,N_5124,N_5160);
xor U5266 (N_5266,N_5158,N_5123);
or U5267 (N_5267,N_5173,N_5107);
nor U5268 (N_5268,N_5106,N_5112);
and U5269 (N_5269,N_5146,N_5189);
and U5270 (N_5270,N_5165,N_5162);
nor U5271 (N_5271,N_5143,N_5167);
nand U5272 (N_5272,N_5100,N_5119);
nor U5273 (N_5273,N_5195,N_5143);
nand U5274 (N_5274,N_5128,N_5178);
nand U5275 (N_5275,N_5118,N_5148);
nor U5276 (N_5276,N_5178,N_5190);
and U5277 (N_5277,N_5179,N_5121);
nor U5278 (N_5278,N_5198,N_5170);
or U5279 (N_5279,N_5147,N_5177);
or U5280 (N_5280,N_5150,N_5136);
xor U5281 (N_5281,N_5197,N_5122);
nand U5282 (N_5282,N_5136,N_5193);
and U5283 (N_5283,N_5120,N_5110);
nor U5284 (N_5284,N_5144,N_5133);
nand U5285 (N_5285,N_5105,N_5159);
xnor U5286 (N_5286,N_5167,N_5196);
or U5287 (N_5287,N_5117,N_5156);
xor U5288 (N_5288,N_5147,N_5144);
nand U5289 (N_5289,N_5168,N_5141);
and U5290 (N_5290,N_5153,N_5164);
xor U5291 (N_5291,N_5139,N_5143);
and U5292 (N_5292,N_5159,N_5109);
and U5293 (N_5293,N_5188,N_5157);
xnor U5294 (N_5294,N_5197,N_5124);
and U5295 (N_5295,N_5115,N_5122);
and U5296 (N_5296,N_5199,N_5121);
or U5297 (N_5297,N_5155,N_5105);
and U5298 (N_5298,N_5192,N_5156);
and U5299 (N_5299,N_5147,N_5135);
and U5300 (N_5300,N_5235,N_5278);
xor U5301 (N_5301,N_5226,N_5266);
and U5302 (N_5302,N_5246,N_5209);
xnor U5303 (N_5303,N_5265,N_5267);
nor U5304 (N_5304,N_5262,N_5269);
or U5305 (N_5305,N_5297,N_5245);
or U5306 (N_5306,N_5260,N_5281);
or U5307 (N_5307,N_5249,N_5210);
nor U5308 (N_5308,N_5200,N_5254);
and U5309 (N_5309,N_5273,N_5224);
or U5310 (N_5310,N_5268,N_5244);
or U5311 (N_5311,N_5258,N_5274);
or U5312 (N_5312,N_5271,N_5221);
nor U5313 (N_5313,N_5299,N_5223);
xor U5314 (N_5314,N_5292,N_5204);
xnor U5315 (N_5315,N_5264,N_5298);
nand U5316 (N_5316,N_5257,N_5287);
xor U5317 (N_5317,N_5283,N_5296);
and U5318 (N_5318,N_5220,N_5205);
nor U5319 (N_5319,N_5232,N_5242);
and U5320 (N_5320,N_5247,N_5212);
nor U5321 (N_5321,N_5241,N_5222);
nand U5322 (N_5322,N_5206,N_5236);
and U5323 (N_5323,N_5207,N_5295);
nand U5324 (N_5324,N_5202,N_5216);
or U5325 (N_5325,N_5284,N_5285);
xor U5326 (N_5326,N_5227,N_5293);
or U5327 (N_5327,N_5231,N_5276);
nor U5328 (N_5328,N_5256,N_5229);
nand U5329 (N_5329,N_5291,N_5261);
nor U5330 (N_5330,N_5294,N_5243);
or U5331 (N_5331,N_5230,N_5286);
or U5332 (N_5332,N_5208,N_5225);
nand U5333 (N_5333,N_5214,N_5237);
nand U5334 (N_5334,N_5234,N_5280);
xor U5335 (N_5335,N_5213,N_5255);
nand U5336 (N_5336,N_5272,N_5289);
xnor U5337 (N_5337,N_5288,N_5275);
nor U5338 (N_5338,N_5251,N_5203);
nor U5339 (N_5339,N_5218,N_5240);
and U5340 (N_5340,N_5277,N_5239);
nand U5341 (N_5341,N_5259,N_5228);
nand U5342 (N_5342,N_5290,N_5201);
or U5343 (N_5343,N_5270,N_5253);
or U5344 (N_5344,N_5215,N_5211);
and U5345 (N_5345,N_5238,N_5282);
or U5346 (N_5346,N_5248,N_5252);
nor U5347 (N_5347,N_5279,N_5219);
xor U5348 (N_5348,N_5233,N_5263);
xnor U5349 (N_5349,N_5217,N_5250);
xnor U5350 (N_5350,N_5215,N_5234);
nor U5351 (N_5351,N_5236,N_5231);
xor U5352 (N_5352,N_5235,N_5262);
or U5353 (N_5353,N_5275,N_5270);
xor U5354 (N_5354,N_5225,N_5257);
nor U5355 (N_5355,N_5264,N_5216);
or U5356 (N_5356,N_5281,N_5235);
and U5357 (N_5357,N_5280,N_5230);
nor U5358 (N_5358,N_5231,N_5266);
nand U5359 (N_5359,N_5234,N_5249);
xnor U5360 (N_5360,N_5226,N_5236);
nand U5361 (N_5361,N_5255,N_5280);
and U5362 (N_5362,N_5292,N_5299);
nor U5363 (N_5363,N_5215,N_5238);
nand U5364 (N_5364,N_5283,N_5295);
and U5365 (N_5365,N_5211,N_5222);
and U5366 (N_5366,N_5212,N_5264);
nand U5367 (N_5367,N_5297,N_5239);
nand U5368 (N_5368,N_5256,N_5226);
xor U5369 (N_5369,N_5233,N_5219);
xor U5370 (N_5370,N_5226,N_5244);
nor U5371 (N_5371,N_5282,N_5283);
nand U5372 (N_5372,N_5268,N_5271);
nand U5373 (N_5373,N_5214,N_5233);
and U5374 (N_5374,N_5259,N_5207);
and U5375 (N_5375,N_5274,N_5254);
nand U5376 (N_5376,N_5266,N_5267);
and U5377 (N_5377,N_5224,N_5265);
xor U5378 (N_5378,N_5217,N_5236);
nor U5379 (N_5379,N_5206,N_5289);
nor U5380 (N_5380,N_5214,N_5241);
nor U5381 (N_5381,N_5212,N_5295);
or U5382 (N_5382,N_5241,N_5230);
and U5383 (N_5383,N_5271,N_5202);
or U5384 (N_5384,N_5271,N_5211);
and U5385 (N_5385,N_5265,N_5230);
or U5386 (N_5386,N_5200,N_5264);
or U5387 (N_5387,N_5251,N_5243);
xnor U5388 (N_5388,N_5264,N_5267);
xnor U5389 (N_5389,N_5251,N_5278);
nor U5390 (N_5390,N_5286,N_5223);
xor U5391 (N_5391,N_5259,N_5235);
or U5392 (N_5392,N_5262,N_5230);
xor U5393 (N_5393,N_5256,N_5237);
or U5394 (N_5394,N_5262,N_5241);
and U5395 (N_5395,N_5242,N_5241);
nand U5396 (N_5396,N_5239,N_5264);
nor U5397 (N_5397,N_5202,N_5269);
xnor U5398 (N_5398,N_5237,N_5212);
xnor U5399 (N_5399,N_5226,N_5291);
xnor U5400 (N_5400,N_5314,N_5351);
xor U5401 (N_5401,N_5371,N_5326);
and U5402 (N_5402,N_5313,N_5308);
nand U5403 (N_5403,N_5360,N_5303);
or U5404 (N_5404,N_5387,N_5370);
or U5405 (N_5405,N_5358,N_5365);
or U5406 (N_5406,N_5354,N_5372);
nor U5407 (N_5407,N_5361,N_5383);
nor U5408 (N_5408,N_5338,N_5304);
nand U5409 (N_5409,N_5368,N_5390);
and U5410 (N_5410,N_5355,N_5386);
nand U5411 (N_5411,N_5311,N_5300);
xor U5412 (N_5412,N_5369,N_5391);
nor U5413 (N_5413,N_5366,N_5328);
nor U5414 (N_5414,N_5348,N_5394);
and U5415 (N_5415,N_5317,N_5339);
and U5416 (N_5416,N_5335,N_5321);
nor U5417 (N_5417,N_5357,N_5374);
and U5418 (N_5418,N_5309,N_5333);
nor U5419 (N_5419,N_5334,N_5380);
nand U5420 (N_5420,N_5340,N_5392);
nand U5421 (N_5421,N_5346,N_5316);
nor U5422 (N_5422,N_5345,N_5343);
xor U5423 (N_5423,N_5322,N_5336);
xnor U5424 (N_5424,N_5363,N_5337);
and U5425 (N_5425,N_5344,N_5381);
or U5426 (N_5426,N_5350,N_5356);
nand U5427 (N_5427,N_5396,N_5325);
nor U5428 (N_5428,N_5301,N_5306);
nor U5429 (N_5429,N_5305,N_5302);
and U5430 (N_5430,N_5331,N_5324);
nand U5431 (N_5431,N_5393,N_5342);
nand U5432 (N_5432,N_5330,N_5362);
or U5433 (N_5433,N_5332,N_5349);
nor U5434 (N_5434,N_5319,N_5323);
or U5435 (N_5435,N_5373,N_5389);
xor U5436 (N_5436,N_5359,N_5364);
and U5437 (N_5437,N_5399,N_5375);
or U5438 (N_5438,N_5329,N_5327);
nor U5439 (N_5439,N_5397,N_5382);
or U5440 (N_5440,N_5312,N_5398);
and U5441 (N_5441,N_5320,N_5307);
nor U5442 (N_5442,N_5395,N_5367);
or U5443 (N_5443,N_5384,N_5377);
xnor U5444 (N_5444,N_5385,N_5379);
xnor U5445 (N_5445,N_5341,N_5347);
and U5446 (N_5446,N_5310,N_5352);
nand U5447 (N_5447,N_5378,N_5318);
or U5448 (N_5448,N_5376,N_5315);
nor U5449 (N_5449,N_5388,N_5353);
nand U5450 (N_5450,N_5316,N_5337);
xor U5451 (N_5451,N_5386,N_5311);
xnor U5452 (N_5452,N_5333,N_5384);
nand U5453 (N_5453,N_5344,N_5356);
nor U5454 (N_5454,N_5330,N_5347);
nand U5455 (N_5455,N_5360,N_5371);
nand U5456 (N_5456,N_5302,N_5328);
xor U5457 (N_5457,N_5329,N_5353);
or U5458 (N_5458,N_5389,N_5301);
and U5459 (N_5459,N_5388,N_5368);
nand U5460 (N_5460,N_5354,N_5332);
nor U5461 (N_5461,N_5364,N_5320);
and U5462 (N_5462,N_5371,N_5372);
nand U5463 (N_5463,N_5345,N_5321);
xor U5464 (N_5464,N_5311,N_5376);
nand U5465 (N_5465,N_5328,N_5343);
nor U5466 (N_5466,N_5351,N_5304);
nor U5467 (N_5467,N_5315,N_5325);
and U5468 (N_5468,N_5372,N_5386);
nor U5469 (N_5469,N_5352,N_5379);
xnor U5470 (N_5470,N_5396,N_5359);
nor U5471 (N_5471,N_5312,N_5353);
and U5472 (N_5472,N_5312,N_5380);
nand U5473 (N_5473,N_5301,N_5377);
or U5474 (N_5474,N_5341,N_5349);
or U5475 (N_5475,N_5343,N_5301);
and U5476 (N_5476,N_5350,N_5398);
or U5477 (N_5477,N_5300,N_5354);
nor U5478 (N_5478,N_5364,N_5345);
nor U5479 (N_5479,N_5368,N_5341);
nand U5480 (N_5480,N_5396,N_5320);
nor U5481 (N_5481,N_5360,N_5357);
or U5482 (N_5482,N_5336,N_5301);
and U5483 (N_5483,N_5396,N_5339);
xor U5484 (N_5484,N_5353,N_5350);
and U5485 (N_5485,N_5301,N_5370);
or U5486 (N_5486,N_5359,N_5356);
nand U5487 (N_5487,N_5310,N_5354);
and U5488 (N_5488,N_5360,N_5351);
and U5489 (N_5489,N_5313,N_5312);
and U5490 (N_5490,N_5385,N_5314);
and U5491 (N_5491,N_5369,N_5330);
nor U5492 (N_5492,N_5337,N_5391);
and U5493 (N_5493,N_5377,N_5333);
or U5494 (N_5494,N_5327,N_5354);
nand U5495 (N_5495,N_5388,N_5326);
nand U5496 (N_5496,N_5398,N_5397);
and U5497 (N_5497,N_5330,N_5385);
nand U5498 (N_5498,N_5327,N_5395);
or U5499 (N_5499,N_5325,N_5399);
or U5500 (N_5500,N_5410,N_5453);
nand U5501 (N_5501,N_5477,N_5495);
xor U5502 (N_5502,N_5485,N_5467);
xor U5503 (N_5503,N_5438,N_5419);
nor U5504 (N_5504,N_5466,N_5423);
nor U5505 (N_5505,N_5431,N_5425);
nor U5506 (N_5506,N_5439,N_5430);
and U5507 (N_5507,N_5475,N_5448);
and U5508 (N_5508,N_5456,N_5421);
xnor U5509 (N_5509,N_5457,N_5460);
nand U5510 (N_5510,N_5446,N_5464);
or U5511 (N_5511,N_5496,N_5433);
or U5512 (N_5512,N_5418,N_5406);
nor U5513 (N_5513,N_5426,N_5444);
nor U5514 (N_5514,N_5494,N_5440);
nand U5515 (N_5515,N_5478,N_5443);
and U5516 (N_5516,N_5452,N_5432);
xnor U5517 (N_5517,N_5458,N_5490);
xnor U5518 (N_5518,N_5486,N_5427);
nand U5519 (N_5519,N_5445,N_5493);
nand U5520 (N_5520,N_5498,N_5488);
nand U5521 (N_5521,N_5465,N_5411);
or U5522 (N_5522,N_5408,N_5437);
and U5523 (N_5523,N_5499,N_5487);
nand U5524 (N_5524,N_5462,N_5407);
and U5525 (N_5525,N_5449,N_5429);
and U5526 (N_5526,N_5435,N_5482);
or U5527 (N_5527,N_5441,N_5491);
or U5528 (N_5528,N_5455,N_5417);
nand U5529 (N_5529,N_5472,N_5424);
and U5530 (N_5530,N_5442,N_5402);
nand U5531 (N_5531,N_5412,N_5483);
and U5532 (N_5532,N_5459,N_5473);
and U5533 (N_5533,N_5409,N_5479);
or U5534 (N_5534,N_5484,N_5415);
or U5535 (N_5535,N_5471,N_5403);
or U5536 (N_5536,N_5428,N_5416);
and U5537 (N_5537,N_5400,N_5434);
or U5538 (N_5538,N_5492,N_5468);
xnor U5539 (N_5539,N_5476,N_5414);
nand U5540 (N_5540,N_5454,N_5469);
xnor U5541 (N_5541,N_5401,N_5420);
or U5542 (N_5542,N_5404,N_5470);
nand U5543 (N_5543,N_5450,N_5480);
nand U5544 (N_5544,N_5436,N_5422);
xnor U5545 (N_5545,N_5413,N_5447);
xnor U5546 (N_5546,N_5451,N_5497);
nand U5547 (N_5547,N_5481,N_5489);
or U5548 (N_5548,N_5461,N_5463);
or U5549 (N_5549,N_5405,N_5474);
nand U5550 (N_5550,N_5405,N_5471);
nand U5551 (N_5551,N_5451,N_5403);
nor U5552 (N_5552,N_5469,N_5442);
nand U5553 (N_5553,N_5417,N_5454);
nor U5554 (N_5554,N_5460,N_5463);
xnor U5555 (N_5555,N_5497,N_5411);
nand U5556 (N_5556,N_5424,N_5425);
nand U5557 (N_5557,N_5456,N_5402);
xor U5558 (N_5558,N_5456,N_5484);
nand U5559 (N_5559,N_5417,N_5483);
xor U5560 (N_5560,N_5482,N_5431);
nand U5561 (N_5561,N_5416,N_5450);
and U5562 (N_5562,N_5438,N_5499);
xnor U5563 (N_5563,N_5448,N_5480);
nand U5564 (N_5564,N_5467,N_5432);
nor U5565 (N_5565,N_5432,N_5457);
or U5566 (N_5566,N_5439,N_5483);
nand U5567 (N_5567,N_5489,N_5433);
nor U5568 (N_5568,N_5444,N_5464);
or U5569 (N_5569,N_5459,N_5406);
and U5570 (N_5570,N_5467,N_5402);
or U5571 (N_5571,N_5437,N_5494);
xnor U5572 (N_5572,N_5465,N_5440);
nor U5573 (N_5573,N_5407,N_5418);
and U5574 (N_5574,N_5405,N_5463);
nand U5575 (N_5575,N_5440,N_5426);
and U5576 (N_5576,N_5485,N_5446);
nand U5577 (N_5577,N_5431,N_5434);
nand U5578 (N_5578,N_5434,N_5462);
nor U5579 (N_5579,N_5467,N_5421);
nor U5580 (N_5580,N_5476,N_5404);
nand U5581 (N_5581,N_5402,N_5408);
xor U5582 (N_5582,N_5449,N_5497);
nor U5583 (N_5583,N_5487,N_5452);
nand U5584 (N_5584,N_5497,N_5432);
xor U5585 (N_5585,N_5499,N_5497);
nor U5586 (N_5586,N_5451,N_5481);
and U5587 (N_5587,N_5479,N_5451);
xor U5588 (N_5588,N_5468,N_5417);
or U5589 (N_5589,N_5426,N_5498);
xnor U5590 (N_5590,N_5402,N_5424);
xor U5591 (N_5591,N_5462,N_5438);
xnor U5592 (N_5592,N_5496,N_5434);
and U5593 (N_5593,N_5467,N_5469);
or U5594 (N_5594,N_5464,N_5427);
nand U5595 (N_5595,N_5423,N_5406);
or U5596 (N_5596,N_5495,N_5409);
or U5597 (N_5597,N_5402,N_5410);
and U5598 (N_5598,N_5417,N_5443);
or U5599 (N_5599,N_5404,N_5490);
or U5600 (N_5600,N_5588,N_5595);
xnor U5601 (N_5601,N_5534,N_5584);
nand U5602 (N_5602,N_5549,N_5589);
xor U5603 (N_5603,N_5597,N_5567);
or U5604 (N_5604,N_5508,N_5545);
xor U5605 (N_5605,N_5590,N_5509);
or U5606 (N_5606,N_5537,N_5511);
and U5607 (N_5607,N_5503,N_5539);
and U5608 (N_5608,N_5535,N_5552);
nor U5609 (N_5609,N_5596,N_5524);
nand U5610 (N_5610,N_5517,N_5502);
nor U5611 (N_5611,N_5566,N_5591);
xor U5612 (N_5612,N_5506,N_5565);
and U5613 (N_5613,N_5547,N_5516);
and U5614 (N_5614,N_5572,N_5510);
nand U5615 (N_5615,N_5518,N_5582);
xnor U5616 (N_5616,N_5512,N_5513);
nor U5617 (N_5617,N_5561,N_5548);
nand U5618 (N_5618,N_5521,N_5520);
nor U5619 (N_5619,N_5526,N_5528);
nor U5620 (N_5620,N_5569,N_5541);
and U5621 (N_5621,N_5557,N_5599);
or U5622 (N_5622,N_5536,N_5556);
nand U5623 (N_5623,N_5515,N_5587);
xor U5624 (N_5624,N_5573,N_5500);
nor U5625 (N_5625,N_5504,N_5581);
nor U5626 (N_5626,N_5533,N_5571);
nand U5627 (N_5627,N_5532,N_5576);
nand U5628 (N_5628,N_5519,N_5583);
xor U5629 (N_5629,N_5594,N_5574);
or U5630 (N_5630,N_5586,N_5577);
or U5631 (N_5631,N_5538,N_5501);
nand U5632 (N_5632,N_5514,N_5507);
and U5633 (N_5633,N_5563,N_5522);
nor U5634 (N_5634,N_5505,N_5542);
nand U5635 (N_5635,N_5568,N_5564);
or U5636 (N_5636,N_5540,N_5529);
xor U5637 (N_5637,N_5575,N_5525);
and U5638 (N_5638,N_5530,N_5598);
xnor U5639 (N_5639,N_5551,N_5527);
nand U5640 (N_5640,N_5544,N_5554);
nand U5641 (N_5641,N_5570,N_5558);
and U5642 (N_5642,N_5562,N_5553);
nand U5643 (N_5643,N_5531,N_5592);
nand U5644 (N_5644,N_5546,N_5585);
or U5645 (N_5645,N_5559,N_5593);
or U5646 (N_5646,N_5543,N_5580);
nand U5647 (N_5647,N_5550,N_5579);
nor U5648 (N_5648,N_5578,N_5560);
nor U5649 (N_5649,N_5555,N_5523);
xnor U5650 (N_5650,N_5570,N_5598);
and U5651 (N_5651,N_5592,N_5573);
xor U5652 (N_5652,N_5593,N_5569);
nor U5653 (N_5653,N_5555,N_5578);
nor U5654 (N_5654,N_5590,N_5516);
nor U5655 (N_5655,N_5534,N_5539);
nor U5656 (N_5656,N_5581,N_5552);
nor U5657 (N_5657,N_5500,N_5507);
nand U5658 (N_5658,N_5516,N_5579);
xnor U5659 (N_5659,N_5506,N_5599);
nand U5660 (N_5660,N_5540,N_5542);
and U5661 (N_5661,N_5553,N_5501);
or U5662 (N_5662,N_5540,N_5593);
nor U5663 (N_5663,N_5507,N_5563);
xor U5664 (N_5664,N_5543,N_5517);
or U5665 (N_5665,N_5548,N_5542);
or U5666 (N_5666,N_5517,N_5507);
xnor U5667 (N_5667,N_5508,N_5528);
nand U5668 (N_5668,N_5550,N_5544);
or U5669 (N_5669,N_5525,N_5517);
nand U5670 (N_5670,N_5585,N_5562);
nand U5671 (N_5671,N_5532,N_5526);
and U5672 (N_5672,N_5598,N_5568);
or U5673 (N_5673,N_5553,N_5549);
nand U5674 (N_5674,N_5578,N_5515);
or U5675 (N_5675,N_5582,N_5530);
or U5676 (N_5676,N_5554,N_5518);
and U5677 (N_5677,N_5537,N_5516);
xnor U5678 (N_5678,N_5516,N_5571);
or U5679 (N_5679,N_5572,N_5543);
nor U5680 (N_5680,N_5565,N_5572);
nor U5681 (N_5681,N_5564,N_5525);
nand U5682 (N_5682,N_5553,N_5561);
nor U5683 (N_5683,N_5533,N_5518);
xor U5684 (N_5684,N_5526,N_5511);
nand U5685 (N_5685,N_5527,N_5560);
nor U5686 (N_5686,N_5550,N_5508);
nor U5687 (N_5687,N_5589,N_5542);
and U5688 (N_5688,N_5534,N_5567);
xnor U5689 (N_5689,N_5544,N_5540);
and U5690 (N_5690,N_5545,N_5595);
and U5691 (N_5691,N_5504,N_5585);
xor U5692 (N_5692,N_5547,N_5513);
and U5693 (N_5693,N_5560,N_5516);
or U5694 (N_5694,N_5580,N_5560);
or U5695 (N_5695,N_5581,N_5573);
or U5696 (N_5696,N_5536,N_5591);
xnor U5697 (N_5697,N_5505,N_5573);
and U5698 (N_5698,N_5598,N_5582);
xor U5699 (N_5699,N_5564,N_5594);
nand U5700 (N_5700,N_5669,N_5685);
xnor U5701 (N_5701,N_5615,N_5667);
nand U5702 (N_5702,N_5664,N_5631);
nand U5703 (N_5703,N_5693,N_5601);
xnor U5704 (N_5704,N_5679,N_5675);
or U5705 (N_5705,N_5613,N_5659);
nor U5706 (N_5706,N_5655,N_5682);
nand U5707 (N_5707,N_5690,N_5673);
and U5708 (N_5708,N_5683,N_5658);
xnor U5709 (N_5709,N_5686,N_5698);
or U5710 (N_5710,N_5648,N_5614);
xor U5711 (N_5711,N_5610,N_5623);
nand U5712 (N_5712,N_5695,N_5634);
nand U5713 (N_5713,N_5652,N_5653);
nand U5714 (N_5714,N_5661,N_5629);
xnor U5715 (N_5715,N_5619,N_5666);
nand U5716 (N_5716,N_5684,N_5642);
nand U5717 (N_5717,N_5628,N_5608);
nand U5718 (N_5718,N_5645,N_5691);
or U5719 (N_5719,N_5689,N_5627);
xor U5720 (N_5720,N_5605,N_5600);
or U5721 (N_5721,N_5654,N_5604);
xnor U5722 (N_5722,N_5650,N_5696);
xnor U5723 (N_5723,N_5636,N_5688);
nor U5724 (N_5724,N_5622,N_5672);
nor U5725 (N_5725,N_5633,N_5609);
nor U5726 (N_5726,N_5616,N_5647);
nor U5727 (N_5727,N_5671,N_5643);
nor U5728 (N_5728,N_5687,N_5692);
xor U5729 (N_5729,N_5699,N_5677);
or U5730 (N_5730,N_5611,N_5632);
nand U5731 (N_5731,N_5626,N_5665);
nor U5732 (N_5732,N_5625,N_5617);
nand U5733 (N_5733,N_5670,N_5602);
or U5734 (N_5734,N_5641,N_5680);
and U5735 (N_5735,N_5621,N_5674);
or U5736 (N_5736,N_5638,N_5668);
nor U5737 (N_5737,N_5637,N_5656);
or U5738 (N_5738,N_5663,N_5651);
nand U5739 (N_5739,N_5620,N_5660);
xor U5740 (N_5740,N_5618,N_5639);
nor U5741 (N_5741,N_5635,N_5649);
nand U5742 (N_5742,N_5603,N_5640);
nand U5743 (N_5743,N_5612,N_5644);
and U5744 (N_5744,N_5697,N_5657);
xor U5745 (N_5745,N_5678,N_5607);
and U5746 (N_5746,N_5646,N_5694);
xor U5747 (N_5747,N_5676,N_5606);
nand U5748 (N_5748,N_5681,N_5662);
and U5749 (N_5749,N_5630,N_5624);
xor U5750 (N_5750,N_5696,N_5675);
or U5751 (N_5751,N_5693,N_5694);
and U5752 (N_5752,N_5667,N_5628);
nor U5753 (N_5753,N_5676,N_5699);
and U5754 (N_5754,N_5635,N_5678);
xnor U5755 (N_5755,N_5657,N_5615);
nand U5756 (N_5756,N_5678,N_5681);
nor U5757 (N_5757,N_5673,N_5661);
nor U5758 (N_5758,N_5642,N_5637);
and U5759 (N_5759,N_5630,N_5693);
and U5760 (N_5760,N_5653,N_5672);
nor U5761 (N_5761,N_5663,N_5660);
nand U5762 (N_5762,N_5661,N_5646);
xnor U5763 (N_5763,N_5628,N_5619);
or U5764 (N_5764,N_5698,N_5682);
and U5765 (N_5765,N_5609,N_5608);
nor U5766 (N_5766,N_5615,N_5620);
xor U5767 (N_5767,N_5616,N_5643);
nor U5768 (N_5768,N_5673,N_5624);
and U5769 (N_5769,N_5638,N_5650);
xnor U5770 (N_5770,N_5667,N_5644);
and U5771 (N_5771,N_5635,N_5604);
nand U5772 (N_5772,N_5643,N_5636);
nor U5773 (N_5773,N_5604,N_5686);
xnor U5774 (N_5774,N_5605,N_5635);
nand U5775 (N_5775,N_5639,N_5697);
and U5776 (N_5776,N_5668,N_5608);
or U5777 (N_5777,N_5661,N_5618);
nand U5778 (N_5778,N_5671,N_5653);
nand U5779 (N_5779,N_5659,N_5606);
xnor U5780 (N_5780,N_5696,N_5626);
nand U5781 (N_5781,N_5699,N_5673);
and U5782 (N_5782,N_5693,N_5644);
xor U5783 (N_5783,N_5602,N_5622);
nand U5784 (N_5784,N_5631,N_5639);
nor U5785 (N_5785,N_5646,N_5699);
and U5786 (N_5786,N_5634,N_5630);
nor U5787 (N_5787,N_5616,N_5636);
nand U5788 (N_5788,N_5615,N_5641);
or U5789 (N_5789,N_5611,N_5693);
nand U5790 (N_5790,N_5675,N_5650);
xor U5791 (N_5791,N_5610,N_5673);
or U5792 (N_5792,N_5606,N_5670);
and U5793 (N_5793,N_5670,N_5667);
xnor U5794 (N_5794,N_5641,N_5674);
xor U5795 (N_5795,N_5606,N_5665);
and U5796 (N_5796,N_5623,N_5601);
and U5797 (N_5797,N_5671,N_5638);
nand U5798 (N_5798,N_5654,N_5699);
xor U5799 (N_5799,N_5633,N_5669);
xnor U5800 (N_5800,N_5772,N_5749);
or U5801 (N_5801,N_5720,N_5758);
and U5802 (N_5802,N_5733,N_5713);
or U5803 (N_5803,N_5711,N_5712);
nand U5804 (N_5804,N_5761,N_5770);
nand U5805 (N_5805,N_5737,N_5729);
or U5806 (N_5806,N_5722,N_5750);
nand U5807 (N_5807,N_5746,N_5784);
or U5808 (N_5808,N_5765,N_5718);
nor U5809 (N_5809,N_5743,N_5783);
xnor U5810 (N_5810,N_5710,N_5779);
or U5811 (N_5811,N_5700,N_5752);
and U5812 (N_5812,N_5794,N_5725);
nor U5813 (N_5813,N_5782,N_5742);
nor U5814 (N_5814,N_5787,N_5745);
and U5815 (N_5815,N_5766,N_5780);
nand U5816 (N_5816,N_5756,N_5786);
and U5817 (N_5817,N_5768,N_5791);
nand U5818 (N_5818,N_5776,N_5785);
xor U5819 (N_5819,N_5714,N_5735);
or U5820 (N_5820,N_5740,N_5738);
or U5821 (N_5821,N_5739,N_5796);
and U5822 (N_5822,N_5767,N_5763);
nand U5823 (N_5823,N_5706,N_5719);
or U5824 (N_5824,N_5790,N_5734);
and U5825 (N_5825,N_5797,N_5753);
xnor U5826 (N_5826,N_5721,N_5774);
or U5827 (N_5827,N_5731,N_5705);
nor U5828 (N_5828,N_5773,N_5762);
nand U5829 (N_5829,N_5723,N_5741);
nand U5830 (N_5830,N_5795,N_5728);
nor U5831 (N_5831,N_5709,N_5792);
nor U5832 (N_5832,N_5788,N_5760);
or U5833 (N_5833,N_5736,N_5730);
nor U5834 (N_5834,N_5769,N_5757);
nand U5835 (N_5835,N_5755,N_5777);
or U5836 (N_5836,N_5771,N_5775);
nor U5837 (N_5837,N_5793,N_5799);
xnor U5838 (N_5838,N_5726,N_5715);
xnor U5839 (N_5839,N_5717,N_5744);
nor U5840 (N_5840,N_5727,N_5704);
or U5841 (N_5841,N_5708,N_5778);
and U5842 (N_5842,N_5759,N_5707);
nand U5843 (N_5843,N_5747,N_5702);
and U5844 (N_5844,N_5732,N_5716);
xnor U5845 (N_5845,N_5703,N_5798);
or U5846 (N_5846,N_5751,N_5781);
nor U5847 (N_5847,N_5724,N_5748);
and U5848 (N_5848,N_5764,N_5754);
nor U5849 (N_5849,N_5701,N_5789);
nand U5850 (N_5850,N_5767,N_5704);
and U5851 (N_5851,N_5763,N_5789);
nand U5852 (N_5852,N_5787,N_5737);
nand U5853 (N_5853,N_5733,N_5761);
nor U5854 (N_5854,N_5724,N_5784);
nand U5855 (N_5855,N_5775,N_5770);
nand U5856 (N_5856,N_5729,N_5763);
or U5857 (N_5857,N_5793,N_5718);
xor U5858 (N_5858,N_5726,N_5747);
xnor U5859 (N_5859,N_5796,N_5720);
or U5860 (N_5860,N_5720,N_5726);
xnor U5861 (N_5861,N_5787,N_5799);
and U5862 (N_5862,N_5773,N_5756);
nor U5863 (N_5863,N_5719,N_5776);
xor U5864 (N_5864,N_5750,N_5794);
nor U5865 (N_5865,N_5706,N_5712);
and U5866 (N_5866,N_5749,N_5771);
or U5867 (N_5867,N_5737,N_5712);
nand U5868 (N_5868,N_5736,N_5702);
xnor U5869 (N_5869,N_5718,N_5731);
nor U5870 (N_5870,N_5760,N_5729);
nand U5871 (N_5871,N_5780,N_5767);
and U5872 (N_5872,N_5714,N_5713);
xor U5873 (N_5873,N_5753,N_5764);
and U5874 (N_5874,N_5724,N_5732);
and U5875 (N_5875,N_5753,N_5720);
xnor U5876 (N_5876,N_5745,N_5763);
nand U5877 (N_5877,N_5795,N_5718);
or U5878 (N_5878,N_5727,N_5787);
nor U5879 (N_5879,N_5757,N_5713);
xnor U5880 (N_5880,N_5745,N_5736);
nor U5881 (N_5881,N_5750,N_5704);
or U5882 (N_5882,N_5766,N_5707);
and U5883 (N_5883,N_5766,N_5772);
and U5884 (N_5884,N_5712,N_5739);
and U5885 (N_5885,N_5730,N_5764);
nor U5886 (N_5886,N_5754,N_5773);
nand U5887 (N_5887,N_5798,N_5717);
xnor U5888 (N_5888,N_5713,N_5704);
and U5889 (N_5889,N_5787,N_5768);
nor U5890 (N_5890,N_5755,N_5748);
nor U5891 (N_5891,N_5735,N_5708);
nand U5892 (N_5892,N_5751,N_5777);
nand U5893 (N_5893,N_5763,N_5784);
xnor U5894 (N_5894,N_5768,N_5756);
xnor U5895 (N_5895,N_5792,N_5791);
nand U5896 (N_5896,N_5723,N_5730);
xor U5897 (N_5897,N_5784,N_5764);
xnor U5898 (N_5898,N_5702,N_5769);
nor U5899 (N_5899,N_5771,N_5739);
nand U5900 (N_5900,N_5822,N_5873);
xnor U5901 (N_5901,N_5831,N_5847);
nand U5902 (N_5902,N_5800,N_5844);
xnor U5903 (N_5903,N_5869,N_5889);
nor U5904 (N_5904,N_5893,N_5802);
xnor U5905 (N_5905,N_5811,N_5857);
or U5906 (N_5906,N_5826,N_5878);
nor U5907 (N_5907,N_5875,N_5818);
nor U5908 (N_5908,N_5841,N_5892);
xor U5909 (N_5909,N_5804,N_5836);
nand U5910 (N_5910,N_5866,N_5828);
nor U5911 (N_5911,N_5840,N_5852);
nor U5912 (N_5912,N_5890,N_5813);
and U5913 (N_5913,N_5882,N_5829);
and U5914 (N_5914,N_5868,N_5881);
and U5915 (N_5915,N_5850,N_5839);
nand U5916 (N_5916,N_5848,N_5805);
xor U5917 (N_5917,N_5842,N_5887);
nor U5918 (N_5918,N_5801,N_5814);
xnor U5919 (N_5919,N_5895,N_5870);
and U5920 (N_5920,N_5825,N_5867);
nor U5921 (N_5921,N_5880,N_5812);
nor U5922 (N_5922,N_5886,N_5810);
xor U5923 (N_5923,N_5858,N_5894);
or U5924 (N_5924,N_5856,N_5860);
xor U5925 (N_5925,N_5806,N_5834);
or U5926 (N_5926,N_5807,N_5888);
nand U5927 (N_5927,N_5820,N_5874);
nor U5928 (N_5928,N_5872,N_5862);
nand U5929 (N_5929,N_5808,N_5821);
or U5930 (N_5930,N_5876,N_5864);
or U5931 (N_5931,N_5837,N_5845);
xnor U5932 (N_5932,N_5803,N_5863);
and U5933 (N_5933,N_5897,N_5824);
nor U5934 (N_5934,N_5883,N_5859);
or U5935 (N_5935,N_5865,N_5817);
or U5936 (N_5936,N_5815,N_5891);
nand U5937 (N_5937,N_5853,N_5899);
nor U5938 (N_5938,N_5843,N_5854);
xnor U5939 (N_5939,N_5846,N_5849);
nand U5940 (N_5940,N_5835,N_5809);
xnor U5941 (N_5941,N_5896,N_5819);
nand U5942 (N_5942,N_5885,N_5861);
or U5943 (N_5943,N_5827,N_5823);
nor U5944 (N_5944,N_5879,N_5833);
nor U5945 (N_5945,N_5816,N_5855);
or U5946 (N_5946,N_5877,N_5830);
xnor U5947 (N_5947,N_5871,N_5838);
or U5948 (N_5948,N_5832,N_5898);
xnor U5949 (N_5949,N_5884,N_5851);
nand U5950 (N_5950,N_5831,N_5881);
and U5951 (N_5951,N_5816,N_5803);
nand U5952 (N_5952,N_5835,N_5825);
nand U5953 (N_5953,N_5876,N_5878);
or U5954 (N_5954,N_5862,N_5861);
nand U5955 (N_5955,N_5870,N_5843);
or U5956 (N_5956,N_5882,N_5846);
nor U5957 (N_5957,N_5897,N_5826);
nor U5958 (N_5958,N_5807,N_5853);
nor U5959 (N_5959,N_5879,N_5878);
and U5960 (N_5960,N_5819,N_5804);
xnor U5961 (N_5961,N_5868,N_5822);
or U5962 (N_5962,N_5801,N_5894);
or U5963 (N_5963,N_5802,N_5816);
nand U5964 (N_5964,N_5816,N_5856);
nand U5965 (N_5965,N_5891,N_5805);
nor U5966 (N_5966,N_5898,N_5860);
and U5967 (N_5967,N_5874,N_5881);
or U5968 (N_5968,N_5874,N_5844);
or U5969 (N_5969,N_5875,N_5850);
nor U5970 (N_5970,N_5834,N_5853);
nand U5971 (N_5971,N_5812,N_5851);
or U5972 (N_5972,N_5834,N_5885);
nor U5973 (N_5973,N_5804,N_5851);
or U5974 (N_5974,N_5835,N_5866);
or U5975 (N_5975,N_5864,N_5873);
and U5976 (N_5976,N_5821,N_5865);
xnor U5977 (N_5977,N_5894,N_5802);
and U5978 (N_5978,N_5815,N_5871);
nand U5979 (N_5979,N_5896,N_5855);
or U5980 (N_5980,N_5840,N_5889);
or U5981 (N_5981,N_5851,N_5853);
nor U5982 (N_5982,N_5848,N_5839);
xnor U5983 (N_5983,N_5837,N_5883);
xor U5984 (N_5984,N_5836,N_5860);
nor U5985 (N_5985,N_5831,N_5855);
nor U5986 (N_5986,N_5859,N_5837);
or U5987 (N_5987,N_5862,N_5844);
xor U5988 (N_5988,N_5890,N_5829);
xnor U5989 (N_5989,N_5810,N_5813);
or U5990 (N_5990,N_5841,N_5829);
nand U5991 (N_5991,N_5856,N_5834);
xnor U5992 (N_5992,N_5815,N_5822);
or U5993 (N_5993,N_5834,N_5855);
nand U5994 (N_5994,N_5804,N_5880);
nand U5995 (N_5995,N_5859,N_5882);
and U5996 (N_5996,N_5812,N_5810);
and U5997 (N_5997,N_5847,N_5860);
nor U5998 (N_5998,N_5820,N_5883);
nand U5999 (N_5999,N_5843,N_5822);
and U6000 (N_6000,N_5964,N_5937);
or U6001 (N_6001,N_5952,N_5951);
nor U6002 (N_6002,N_5911,N_5947);
and U6003 (N_6003,N_5933,N_5912);
and U6004 (N_6004,N_5981,N_5924);
and U6005 (N_6005,N_5980,N_5903);
xnor U6006 (N_6006,N_5996,N_5945);
nand U6007 (N_6007,N_5907,N_5977);
nand U6008 (N_6008,N_5992,N_5969);
or U6009 (N_6009,N_5915,N_5906);
nor U6010 (N_6010,N_5923,N_5913);
nor U6011 (N_6011,N_5901,N_5987);
xor U6012 (N_6012,N_5925,N_5998);
and U6013 (N_6013,N_5978,N_5918);
nand U6014 (N_6014,N_5982,N_5914);
or U6015 (N_6015,N_5928,N_5979);
nand U6016 (N_6016,N_5950,N_5986);
xor U6017 (N_6017,N_5968,N_5963);
or U6018 (N_6018,N_5984,N_5946);
and U6019 (N_6019,N_5935,N_5938);
and U6020 (N_6020,N_5993,N_5932);
xnor U6021 (N_6021,N_5941,N_5919);
nand U6022 (N_6022,N_5967,N_5959);
nand U6023 (N_6023,N_5957,N_5965);
nand U6024 (N_6024,N_5955,N_5910);
nor U6025 (N_6025,N_5962,N_5900);
nor U6026 (N_6026,N_5976,N_5917);
nand U6027 (N_6027,N_5940,N_5909);
or U6028 (N_6028,N_5989,N_5995);
nand U6029 (N_6029,N_5948,N_5970);
nor U6030 (N_6030,N_5922,N_5997);
and U6031 (N_6031,N_5973,N_5966);
nor U6032 (N_6032,N_5931,N_5944);
or U6033 (N_6033,N_5916,N_5942);
xnor U6034 (N_6034,N_5983,N_5988);
nor U6035 (N_6035,N_5960,N_5902);
or U6036 (N_6036,N_5930,N_5905);
or U6037 (N_6037,N_5920,N_5934);
xor U6038 (N_6038,N_5974,N_5904);
nand U6039 (N_6039,N_5943,N_5971);
or U6040 (N_6040,N_5990,N_5958);
nor U6041 (N_6041,N_5949,N_5954);
nor U6042 (N_6042,N_5927,N_5908);
xnor U6043 (N_6043,N_5961,N_5994);
and U6044 (N_6044,N_5929,N_5999);
or U6045 (N_6045,N_5972,N_5953);
nor U6046 (N_6046,N_5921,N_5985);
nand U6047 (N_6047,N_5975,N_5936);
xnor U6048 (N_6048,N_5939,N_5956);
or U6049 (N_6049,N_5926,N_5991);
nand U6050 (N_6050,N_5907,N_5904);
nor U6051 (N_6051,N_5935,N_5930);
and U6052 (N_6052,N_5970,N_5975);
nor U6053 (N_6053,N_5965,N_5934);
nand U6054 (N_6054,N_5956,N_5921);
or U6055 (N_6055,N_5915,N_5932);
and U6056 (N_6056,N_5908,N_5994);
or U6057 (N_6057,N_5953,N_5926);
nor U6058 (N_6058,N_5970,N_5947);
or U6059 (N_6059,N_5980,N_5913);
and U6060 (N_6060,N_5984,N_5953);
or U6061 (N_6061,N_5951,N_5928);
nor U6062 (N_6062,N_5921,N_5952);
xnor U6063 (N_6063,N_5927,N_5996);
and U6064 (N_6064,N_5993,N_5940);
xor U6065 (N_6065,N_5982,N_5999);
xor U6066 (N_6066,N_5992,N_5966);
nand U6067 (N_6067,N_5964,N_5994);
and U6068 (N_6068,N_5945,N_5993);
or U6069 (N_6069,N_5956,N_5995);
nand U6070 (N_6070,N_5903,N_5955);
nor U6071 (N_6071,N_5968,N_5908);
nor U6072 (N_6072,N_5916,N_5971);
or U6073 (N_6073,N_5941,N_5900);
xor U6074 (N_6074,N_5962,N_5944);
nand U6075 (N_6075,N_5998,N_5915);
or U6076 (N_6076,N_5956,N_5986);
nor U6077 (N_6077,N_5963,N_5914);
nand U6078 (N_6078,N_5950,N_5914);
and U6079 (N_6079,N_5958,N_5943);
nand U6080 (N_6080,N_5952,N_5917);
nor U6081 (N_6081,N_5979,N_5915);
or U6082 (N_6082,N_5912,N_5944);
xnor U6083 (N_6083,N_5927,N_5960);
nand U6084 (N_6084,N_5946,N_5912);
and U6085 (N_6085,N_5983,N_5952);
xor U6086 (N_6086,N_5925,N_5937);
and U6087 (N_6087,N_5925,N_5901);
and U6088 (N_6088,N_5936,N_5910);
nor U6089 (N_6089,N_5983,N_5972);
xnor U6090 (N_6090,N_5961,N_5942);
nand U6091 (N_6091,N_5949,N_5938);
and U6092 (N_6092,N_5976,N_5934);
xnor U6093 (N_6093,N_5962,N_5902);
nand U6094 (N_6094,N_5948,N_5954);
nand U6095 (N_6095,N_5958,N_5946);
and U6096 (N_6096,N_5940,N_5925);
and U6097 (N_6097,N_5922,N_5994);
or U6098 (N_6098,N_5989,N_5918);
nor U6099 (N_6099,N_5994,N_5937);
nand U6100 (N_6100,N_6065,N_6031);
nand U6101 (N_6101,N_6076,N_6020);
nand U6102 (N_6102,N_6048,N_6028);
and U6103 (N_6103,N_6066,N_6030);
nand U6104 (N_6104,N_6087,N_6091);
nor U6105 (N_6105,N_6069,N_6059);
and U6106 (N_6106,N_6094,N_6061);
or U6107 (N_6107,N_6085,N_6018);
nor U6108 (N_6108,N_6003,N_6058);
xnor U6109 (N_6109,N_6027,N_6055);
nand U6110 (N_6110,N_6036,N_6074);
nand U6111 (N_6111,N_6013,N_6099);
nor U6112 (N_6112,N_6090,N_6071);
and U6113 (N_6113,N_6043,N_6038);
xor U6114 (N_6114,N_6054,N_6029);
nand U6115 (N_6115,N_6008,N_6060);
or U6116 (N_6116,N_6052,N_6002);
nand U6117 (N_6117,N_6077,N_6072);
nand U6118 (N_6118,N_6005,N_6096);
xnor U6119 (N_6119,N_6047,N_6082);
nand U6120 (N_6120,N_6022,N_6001);
and U6121 (N_6121,N_6068,N_6088);
nor U6122 (N_6122,N_6093,N_6024);
and U6123 (N_6123,N_6017,N_6000);
xor U6124 (N_6124,N_6034,N_6070);
xnor U6125 (N_6125,N_6039,N_6051);
xor U6126 (N_6126,N_6086,N_6041);
or U6127 (N_6127,N_6062,N_6019);
xor U6128 (N_6128,N_6011,N_6092);
and U6129 (N_6129,N_6035,N_6015);
xnor U6130 (N_6130,N_6089,N_6042);
xor U6131 (N_6131,N_6073,N_6084);
nor U6132 (N_6132,N_6050,N_6046);
nor U6133 (N_6133,N_6007,N_6095);
or U6134 (N_6134,N_6032,N_6023);
nand U6135 (N_6135,N_6012,N_6040);
nor U6136 (N_6136,N_6057,N_6080);
or U6137 (N_6137,N_6021,N_6098);
or U6138 (N_6138,N_6033,N_6025);
or U6139 (N_6139,N_6078,N_6045);
xor U6140 (N_6140,N_6075,N_6083);
and U6141 (N_6141,N_6010,N_6097);
nand U6142 (N_6142,N_6053,N_6009);
xor U6143 (N_6143,N_6081,N_6067);
or U6144 (N_6144,N_6044,N_6063);
nand U6145 (N_6145,N_6064,N_6049);
and U6146 (N_6146,N_6006,N_6037);
or U6147 (N_6147,N_6004,N_6016);
nor U6148 (N_6148,N_6014,N_6079);
xnor U6149 (N_6149,N_6056,N_6026);
nand U6150 (N_6150,N_6007,N_6088);
xor U6151 (N_6151,N_6018,N_6043);
or U6152 (N_6152,N_6059,N_6020);
nand U6153 (N_6153,N_6052,N_6003);
nand U6154 (N_6154,N_6084,N_6091);
nor U6155 (N_6155,N_6041,N_6020);
or U6156 (N_6156,N_6018,N_6052);
or U6157 (N_6157,N_6045,N_6080);
nor U6158 (N_6158,N_6061,N_6018);
nor U6159 (N_6159,N_6055,N_6002);
nand U6160 (N_6160,N_6063,N_6091);
nand U6161 (N_6161,N_6070,N_6018);
nor U6162 (N_6162,N_6057,N_6069);
and U6163 (N_6163,N_6004,N_6050);
xor U6164 (N_6164,N_6071,N_6038);
nand U6165 (N_6165,N_6078,N_6060);
xnor U6166 (N_6166,N_6085,N_6021);
or U6167 (N_6167,N_6041,N_6094);
or U6168 (N_6168,N_6080,N_6099);
xnor U6169 (N_6169,N_6072,N_6031);
and U6170 (N_6170,N_6063,N_6071);
nor U6171 (N_6171,N_6034,N_6062);
and U6172 (N_6172,N_6023,N_6034);
nor U6173 (N_6173,N_6003,N_6096);
and U6174 (N_6174,N_6040,N_6048);
or U6175 (N_6175,N_6053,N_6080);
xor U6176 (N_6176,N_6081,N_6066);
or U6177 (N_6177,N_6019,N_6027);
xor U6178 (N_6178,N_6058,N_6063);
or U6179 (N_6179,N_6067,N_6020);
and U6180 (N_6180,N_6003,N_6062);
and U6181 (N_6181,N_6061,N_6072);
or U6182 (N_6182,N_6043,N_6081);
nand U6183 (N_6183,N_6086,N_6025);
and U6184 (N_6184,N_6021,N_6046);
nor U6185 (N_6185,N_6012,N_6026);
xor U6186 (N_6186,N_6023,N_6022);
or U6187 (N_6187,N_6066,N_6035);
nand U6188 (N_6188,N_6016,N_6073);
or U6189 (N_6189,N_6013,N_6052);
or U6190 (N_6190,N_6011,N_6021);
and U6191 (N_6191,N_6048,N_6038);
and U6192 (N_6192,N_6013,N_6094);
or U6193 (N_6193,N_6086,N_6032);
xnor U6194 (N_6194,N_6082,N_6058);
xnor U6195 (N_6195,N_6025,N_6037);
and U6196 (N_6196,N_6089,N_6050);
or U6197 (N_6197,N_6090,N_6005);
nor U6198 (N_6198,N_6092,N_6050);
and U6199 (N_6199,N_6022,N_6039);
and U6200 (N_6200,N_6116,N_6128);
nand U6201 (N_6201,N_6193,N_6162);
or U6202 (N_6202,N_6117,N_6187);
and U6203 (N_6203,N_6124,N_6134);
nor U6204 (N_6204,N_6111,N_6107);
or U6205 (N_6205,N_6100,N_6196);
and U6206 (N_6206,N_6147,N_6177);
xor U6207 (N_6207,N_6131,N_6120);
and U6208 (N_6208,N_6118,N_6161);
nand U6209 (N_6209,N_6188,N_6185);
xnor U6210 (N_6210,N_6165,N_6127);
and U6211 (N_6211,N_6126,N_6137);
or U6212 (N_6212,N_6155,N_6144);
and U6213 (N_6213,N_6167,N_6191);
nand U6214 (N_6214,N_6141,N_6108);
nand U6215 (N_6215,N_6146,N_6143);
xor U6216 (N_6216,N_6184,N_6179);
or U6217 (N_6217,N_6168,N_6174);
nand U6218 (N_6218,N_6106,N_6152);
nor U6219 (N_6219,N_6145,N_6139);
nor U6220 (N_6220,N_6156,N_6151);
or U6221 (N_6221,N_6110,N_6136);
xor U6222 (N_6222,N_6138,N_6190);
xor U6223 (N_6223,N_6103,N_6173);
nand U6224 (N_6224,N_6142,N_6166);
xnor U6225 (N_6225,N_6172,N_6169);
nor U6226 (N_6226,N_6122,N_6153);
nor U6227 (N_6227,N_6158,N_6102);
or U6228 (N_6228,N_6170,N_6197);
and U6229 (N_6229,N_6189,N_6135);
nand U6230 (N_6230,N_6140,N_6104);
nand U6231 (N_6231,N_6171,N_6178);
or U6232 (N_6232,N_6183,N_6194);
xor U6233 (N_6233,N_6105,N_6149);
nor U6234 (N_6234,N_6130,N_6133);
or U6235 (N_6235,N_6199,N_6129);
nor U6236 (N_6236,N_6181,N_6157);
nand U6237 (N_6237,N_6182,N_6125);
and U6238 (N_6238,N_6195,N_6115);
or U6239 (N_6239,N_6113,N_6198);
nand U6240 (N_6240,N_6154,N_6132);
and U6241 (N_6241,N_6112,N_6121);
or U6242 (N_6242,N_6101,N_6176);
nor U6243 (N_6243,N_6192,N_6186);
xor U6244 (N_6244,N_6180,N_6159);
xor U6245 (N_6245,N_6114,N_6163);
nand U6246 (N_6246,N_6119,N_6109);
xor U6247 (N_6247,N_6123,N_6148);
xnor U6248 (N_6248,N_6175,N_6150);
and U6249 (N_6249,N_6164,N_6160);
nand U6250 (N_6250,N_6109,N_6118);
xnor U6251 (N_6251,N_6138,N_6122);
xnor U6252 (N_6252,N_6108,N_6110);
nand U6253 (N_6253,N_6190,N_6117);
xor U6254 (N_6254,N_6173,N_6162);
nor U6255 (N_6255,N_6162,N_6159);
or U6256 (N_6256,N_6196,N_6122);
nand U6257 (N_6257,N_6189,N_6187);
xor U6258 (N_6258,N_6140,N_6174);
xor U6259 (N_6259,N_6174,N_6153);
nand U6260 (N_6260,N_6190,N_6187);
and U6261 (N_6261,N_6132,N_6129);
and U6262 (N_6262,N_6133,N_6173);
nand U6263 (N_6263,N_6102,N_6141);
nand U6264 (N_6264,N_6133,N_6140);
and U6265 (N_6265,N_6149,N_6154);
nor U6266 (N_6266,N_6163,N_6117);
and U6267 (N_6267,N_6163,N_6190);
and U6268 (N_6268,N_6155,N_6196);
xor U6269 (N_6269,N_6103,N_6162);
and U6270 (N_6270,N_6157,N_6164);
xor U6271 (N_6271,N_6135,N_6142);
nand U6272 (N_6272,N_6187,N_6103);
nor U6273 (N_6273,N_6177,N_6183);
nor U6274 (N_6274,N_6198,N_6133);
or U6275 (N_6275,N_6169,N_6163);
nand U6276 (N_6276,N_6148,N_6115);
nor U6277 (N_6277,N_6135,N_6131);
nor U6278 (N_6278,N_6170,N_6196);
nor U6279 (N_6279,N_6181,N_6114);
or U6280 (N_6280,N_6152,N_6160);
xnor U6281 (N_6281,N_6169,N_6199);
and U6282 (N_6282,N_6156,N_6146);
or U6283 (N_6283,N_6163,N_6115);
nor U6284 (N_6284,N_6111,N_6170);
or U6285 (N_6285,N_6111,N_6186);
xnor U6286 (N_6286,N_6194,N_6172);
nor U6287 (N_6287,N_6177,N_6123);
or U6288 (N_6288,N_6175,N_6181);
nand U6289 (N_6289,N_6106,N_6145);
xor U6290 (N_6290,N_6179,N_6133);
and U6291 (N_6291,N_6178,N_6197);
xnor U6292 (N_6292,N_6106,N_6142);
or U6293 (N_6293,N_6175,N_6184);
and U6294 (N_6294,N_6103,N_6116);
nor U6295 (N_6295,N_6129,N_6135);
xnor U6296 (N_6296,N_6110,N_6169);
xnor U6297 (N_6297,N_6192,N_6110);
or U6298 (N_6298,N_6146,N_6124);
and U6299 (N_6299,N_6149,N_6129);
and U6300 (N_6300,N_6290,N_6270);
nand U6301 (N_6301,N_6216,N_6208);
xnor U6302 (N_6302,N_6202,N_6264);
nand U6303 (N_6303,N_6228,N_6284);
nand U6304 (N_6304,N_6260,N_6278);
xnor U6305 (N_6305,N_6224,N_6223);
or U6306 (N_6306,N_6220,N_6239);
or U6307 (N_6307,N_6222,N_6229);
xnor U6308 (N_6308,N_6214,N_6247);
nand U6309 (N_6309,N_6227,N_6217);
and U6310 (N_6310,N_6253,N_6203);
nand U6311 (N_6311,N_6241,N_6206);
nand U6312 (N_6312,N_6271,N_6280);
and U6313 (N_6313,N_6221,N_6200);
and U6314 (N_6314,N_6275,N_6295);
nand U6315 (N_6315,N_6233,N_6276);
and U6316 (N_6316,N_6263,N_6245);
nand U6317 (N_6317,N_6244,N_6225);
or U6318 (N_6318,N_6257,N_6268);
xnor U6319 (N_6319,N_6265,N_6234);
nand U6320 (N_6320,N_6219,N_6266);
nand U6321 (N_6321,N_6248,N_6287);
nand U6322 (N_6322,N_6289,N_6205);
nor U6323 (N_6323,N_6237,N_6249);
nor U6324 (N_6324,N_6281,N_6273);
nor U6325 (N_6325,N_6279,N_6232);
xor U6326 (N_6326,N_6293,N_6294);
xor U6327 (N_6327,N_6211,N_6242);
nand U6328 (N_6328,N_6209,N_6252);
and U6329 (N_6329,N_6296,N_6207);
or U6330 (N_6330,N_6261,N_6201);
nand U6331 (N_6331,N_6298,N_6297);
nand U6332 (N_6332,N_6274,N_6277);
and U6333 (N_6333,N_6286,N_6259);
or U6334 (N_6334,N_6210,N_6240);
and U6335 (N_6335,N_6262,N_6291);
or U6336 (N_6336,N_6256,N_6299);
or U6337 (N_6337,N_6254,N_6218);
nor U6338 (N_6338,N_6283,N_6272);
or U6339 (N_6339,N_6226,N_6238);
or U6340 (N_6340,N_6255,N_6215);
and U6341 (N_6341,N_6251,N_6204);
and U6342 (N_6342,N_6269,N_6288);
and U6343 (N_6343,N_6292,N_6246);
nand U6344 (N_6344,N_6212,N_6235);
nor U6345 (N_6345,N_6250,N_6231);
xnor U6346 (N_6346,N_6267,N_6236);
nand U6347 (N_6347,N_6243,N_6282);
xor U6348 (N_6348,N_6213,N_6285);
and U6349 (N_6349,N_6258,N_6230);
xor U6350 (N_6350,N_6279,N_6200);
xnor U6351 (N_6351,N_6251,N_6267);
nor U6352 (N_6352,N_6268,N_6273);
nand U6353 (N_6353,N_6252,N_6262);
nor U6354 (N_6354,N_6294,N_6213);
and U6355 (N_6355,N_6218,N_6225);
nor U6356 (N_6356,N_6257,N_6283);
and U6357 (N_6357,N_6266,N_6298);
xor U6358 (N_6358,N_6217,N_6226);
nand U6359 (N_6359,N_6242,N_6205);
or U6360 (N_6360,N_6269,N_6290);
nand U6361 (N_6361,N_6257,N_6249);
nor U6362 (N_6362,N_6272,N_6233);
xnor U6363 (N_6363,N_6207,N_6203);
or U6364 (N_6364,N_6253,N_6249);
and U6365 (N_6365,N_6232,N_6255);
nor U6366 (N_6366,N_6247,N_6287);
and U6367 (N_6367,N_6227,N_6287);
and U6368 (N_6368,N_6220,N_6213);
nor U6369 (N_6369,N_6250,N_6249);
nor U6370 (N_6370,N_6225,N_6279);
nand U6371 (N_6371,N_6248,N_6257);
nor U6372 (N_6372,N_6259,N_6267);
and U6373 (N_6373,N_6290,N_6229);
and U6374 (N_6374,N_6298,N_6263);
xor U6375 (N_6375,N_6225,N_6215);
or U6376 (N_6376,N_6228,N_6238);
nor U6377 (N_6377,N_6292,N_6242);
nor U6378 (N_6378,N_6212,N_6298);
or U6379 (N_6379,N_6265,N_6225);
nand U6380 (N_6380,N_6228,N_6264);
xnor U6381 (N_6381,N_6278,N_6292);
and U6382 (N_6382,N_6294,N_6278);
xnor U6383 (N_6383,N_6270,N_6293);
xor U6384 (N_6384,N_6294,N_6267);
xnor U6385 (N_6385,N_6270,N_6272);
and U6386 (N_6386,N_6218,N_6273);
nor U6387 (N_6387,N_6234,N_6244);
and U6388 (N_6388,N_6257,N_6286);
nor U6389 (N_6389,N_6206,N_6259);
nor U6390 (N_6390,N_6299,N_6208);
nand U6391 (N_6391,N_6241,N_6242);
nor U6392 (N_6392,N_6223,N_6277);
and U6393 (N_6393,N_6202,N_6284);
and U6394 (N_6394,N_6281,N_6236);
and U6395 (N_6395,N_6285,N_6274);
xnor U6396 (N_6396,N_6265,N_6202);
xor U6397 (N_6397,N_6235,N_6222);
nor U6398 (N_6398,N_6257,N_6297);
or U6399 (N_6399,N_6200,N_6257);
xnor U6400 (N_6400,N_6335,N_6352);
nor U6401 (N_6401,N_6303,N_6355);
and U6402 (N_6402,N_6343,N_6320);
xor U6403 (N_6403,N_6319,N_6308);
nor U6404 (N_6404,N_6385,N_6377);
xor U6405 (N_6405,N_6324,N_6382);
nor U6406 (N_6406,N_6334,N_6338);
and U6407 (N_6407,N_6375,N_6371);
nand U6408 (N_6408,N_6394,N_6353);
nor U6409 (N_6409,N_6364,N_6345);
nand U6410 (N_6410,N_6384,N_6391);
or U6411 (N_6411,N_6350,N_6347);
xnor U6412 (N_6412,N_6331,N_6387);
nor U6413 (N_6413,N_6348,N_6367);
or U6414 (N_6414,N_6392,N_6346);
and U6415 (N_6415,N_6369,N_6380);
and U6416 (N_6416,N_6313,N_6310);
nor U6417 (N_6417,N_6368,N_6378);
and U6418 (N_6418,N_6399,N_6314);
and U6419 (N_6419,N_6351,N_6366);
or U6420 (N_6420,N_6396,N_6316);
and U6421 (N_6421,N_6341,N_6306);
nand U6422 (N_6422,N_6357,N_6361);
nand U6423 (N_6423,N_6373,N_6311);
or U6424 (N_6424,N_6342,N_6356);
nand U6425 (N_6425,N_6300,N_6302);
or U6426 (N_6426,N_6325,N_6390);
xnor U6427 (N_6427,N_6318,N_6379);
nand U6428 (N_6428,N_6388,N_6363);
nand U6429 (N_6429,N_6395,N_6307);
nand U6430 (N_6430,N_6327,N_6365);
nand U6431 (N_6431,N_6315,N_6386);
nor U6432 (N_6432,N_6322,N_6389);
and U6433 (N_6433,N_6344,N_6332);
and U6434 (N_6434,N_6362,N_6323);
and U6435 (N_6435,N_6333,N_6370);
nand U6436 (N_6436,N_6337,N_6340);
nor U6437 (N_6437,N_6312,N_6398);
or U6438 (N_6438,N_6358,N_6383);
xor U6439 (N_6439,N_6317,N_6330);
nor U6440 (N_6440,N_6336,N_6393);
xor U6441 (N_6441,N_6329,N_6360);
nand U6442 (N_6442,N_6339,N_6397);
and U6443 (N_6443,N_6328,N_6374);
nand U6444 (N_6444,N_6326,N_6376);
nor U6445 (N_6445,N_6309,N_6349);
nor U6446 (N_6446,N_6354,N_6301);
or U6447 (N_6447,N_6304,N_6372);
nor U6448 (N_6448,N_6321,N_6305);
or U6449 (N_6449,N_6359,N_6381);
nor U6450 (N_6450,N_6306,N_6325);
nor U6451 (N_6451,N_6338,N_6324);
nand U6452 (N_6452,N_6378,N_6329);
and U6453 (N_6453,N_6321,N_6355);
and U6454 (N_6454,N_6345,N_6355);
xnor U6455 (N_6455,N_6318,N_6381);
and U6456 (N_6456,N_6364,N_6334);
xnor U6457 (N_6457,N_6319,N_6352);
nand U6458 (N_6458,N_6324,N_6329);
xnor U6459 (N_6459,N_6352,N_6348);
and U6460 (N_6460,N_6343,N_6370);
nand U6461 (N_6461,N_6306,N_6329);
and U6462 (N_6462,N_6328,N_6315);
nor U6463 (N_6463,N_6357,N_6315);
or U6464 (N_6464,N_6320,N_6331);
nand U6465 (N_6465,N_6362,N_6373);
nor U6466 (N_6466,N_6341,N_6395);
xor U6467 (N_6467,N_6390,N_6328);
and U6468 (N_6468,N_6318,N_6355);
or U6469 (N_6469,N_6319,N_6345);
nor U6470 (N_6470,N_6313,N_6360);
nor U6471 (N_6471,N_6381,N_6337);
or U6472 (N_6472,N_6309,N_6356);
nor U6473 (N_6473,N_6383,N_6395);
nand U6474 (N_6474,N_6313,N_6355);
and U6475 (N_6475,N_6320,N_6338);
nand U6476 (N_6476,N_6370,N_6392);
or U6477 (N_6477,N_6322,N_6364);
and U6478 (N_6478,N_6399,N_6308);
nand U6479 (N_6479,N_6323,N_6383);
nor U6480 (N_6480,N_6397,N_6346);
or U6481 (N_6481,N_6368,N_6321);
xor U6482 (N_6482,N_6314,N_6343);
nand U6483 (N_6483,N_6304,N_6353);
xnor U6484 (N_6484,N_6358,N_6371);
nor U6485 (N_6485,N_6395,N_6354);
and U6486 (N_6486,N_6388,N_6385);
xor U6487 (N_6487,N_6320,N_6321);
xor U6488 (N_6488,N_6309,N_6345);
nor U6489 (N_6489,N_6306,N_6379);
nand U6490 (N_6490,N_6353,N_6307);
nand U6491 (N_6491,N_6320,N_6350);
xor U6492 (N_6492,N_6387,N_6341);
nor U6493 (N_6493,N_6372,N_6342);
or U6494 (N_6494,N_6318,N_6376);
and U6495 (N_6495,N_6324,N_6388);
xor U6496 (N_6496,N_6344,N_6327);
xnor U6497 (N_6497,N_6358,N_6347);
or U6498 (N_6498,N_6342,N_6312);
and U6499 (N_6499,N_6394,N_6318);
and U6500 (N_6500,N_6441,N_6452);
xnor U6501 (N_6501,N_6420,N_6470);
xor U6502 (N_6502,N_6438,N_6424);
or U6503 (N_6503,N_6484,N_6499);
xor U6504 (N_6504,N_6475,N_6479);
or U6505 (N_6505,N_6423,N_6461);
xor U6506 (N_6506,N_6442,N_6422);
nor U6507 (N_6507,N_6413,N_6495);
nor U6508 (N_6508,N_6444,N_6410);
nor U6509 (N_6509,N_6476,N_6489);
or U6510 (N_6510,N_6460,N_6412);
nand U6511 (N_6511,N_6404,N_6436);
xor U6512 (N_6512,N_6473,N_6482);
or U6513 (N_6513,N_6431,N_6414);
xnor U6514 (N_6514,N_6439,N_6491);
and U6515 (N_6515,N_6400,N_6402);
nor U6516 (N_6516,N_6401,N_6490);
nor U6517 (N_6517,N_6497,N_6468);
and U6518 (N_6518,N_6471,N_6433);
xor U6519 (N_6519,N_6455,N_6411);
xor U6520 (N_6520,N_6406,N_6437);
or U6521 (N_6521,N_6492,N_6483);
nand U6522 (N_6522,N_6458,N_6427);
and U6523 (N_6523,N_6477,N_6498);
xnor U6524 (N_6524,N_6496,N_6403);
nor U6525 (N_6525,N_6421,N_6449);
xor U6526 (N_6526,N_6487,N_6426);
or U6527 (N_6527,N_6472,N_6453);
nor U6528 (N_6528,N_6417,N_6480);
xnor U6529 (N_6529,N_6469,N_6459);
and U6530 (N_6530,N_6457,N_6409);
xnor U6531 (N_6531,N_6467,N_6446);
and U6532 (N_6532,N_6407,N_6447);
and U6533 (N_6533,N_6408,N_6456);
nor U6534 (N_6534,N_6454,N_6464);
or U6535 (N_6535,N_6430,N_6494);
nand U6536 (N_6536,N_6440,N_6465);
or U6537 (N_6537,N_6462,N_6478);
nand U6538 (N_6538,N_6466,N_6415);
nand U6539 (N_6539,N_6448,N_6493);
nor U6540 (N_6540,N_6432,N_6450);
or U6541 (N_6541,N_6418,N_6425);
xnor U6542 (N_6542,N_6451,N_6445);
nand U6543 (N_6543,N_6486,N_6434);
nor U6544 (N_6544,N_6481,N_6419);
xor U6545 (N_6545,N_6435,N_6443);
nand U6546 (N_6546,N_6474,N_6429);
and U6547 (N_6547,N_6416,N_6463);
and U6548 (N_6548,N_6485,N_6488);
nand U6549 (N_6549,N_6405,N_6428);
and U6550 (N_6550,N_6433,N_6481);
nand U6551 (N_6551,N_6425,N_6451);
nand U6552 (N_6552,N_6454,N_6414);
and U6553 (N_6553,N_6489,N_6477);
nor U6554 (N_6554,N_6454,N_6478);
and U6555 (N_6555,N_6472,N_6459);
xor U6556 (N_6556,N_6492,N_6426);
xor U6557 (N_6557,N_6439,N_6425);
and U6558 (N_6558,N_6446,N_6404);
nand U6559 (N_6559,N_6496,N_6432);
nand U6560 (N_6560,N_6487,N_6498);
xnor U6561 (N_6561,N_6485,N_6441);
and U6562 (N_6562,N_6405,N_6421);
nand U6563 (N_6563,N_6495,N_6402);
nand U6564 (N_6564,N_6481,N_6415);
nand U6565 (N_6565,N_6442,N_6464);
nand U6566 (N_6566,N_6476,N_6486);
and U6567 (N_6567,N_6453,N_6460);
and U6568 (N_6568,N_6492,N_6433);
nand U6569 (N_6569,N_6427,N_6499);
xor U6570 (N_6570,N_6416,N_6449);
nor U6571 (N_6571,N_6447,N_6403);
and U6572 (N_6572,N_6403,N_6469);
and U6573 (N_6573,N_6484,N_6451);
xnor U6574 (N_6574,N_6479,N_6413);
nand U6575 (N_6575,N_6411,N_6433);
and U6576 (N_6576,N_6456,N_6420);
or U6577 (N_6577,N_6413,N_6468);
xnor U6578 (N_6578,N_6494,N_6478);
nand U6579 (N_6579,N_6466,N_6427);
and U6580 (N_6580,N_6473,N_6494);
nor U6581 (N_6581,N_6424,N_6419);
nand U6582 (N_6582,N_6402,N_6411);
xor U6583 (N_6583,N_6464,N_6470);
nor U6584 (N_6584,N_6403,N_6401);
and U6585 (N_6585,N_6470,N_6433);
and U6586 (N_6586,N_6497,N_6481);
xor U6587 (N_6587,N_6441,N_6491);
or U6588 (N_6588,N_6407,N_6423);
nor U6589 (N_6589,N_6421,N_6419);
xor U6590 (N_6590,N_6469,N_6479);
and U6591 (N_6591,N_6442,N_6421);
nand U6592 (N_6592,N_6434,N_6453);
and U6593 (N_6593,N_6454,N_6498);
nand U6594 (N_6594,N_6437,N_6455);
or U6595 (N_6595,N_6486,N_6443);
nand U6596 (N_6596,N_6440,N_6479);
xor U6597 (N_6597,N_6469,N_6423);
or U6598 (N_6598,N_6485,N_6429);
and U6599 (N_6599,N_6483,N_6411);
and U6600 (N_6600,N_6559,N_6583);
xnor U6601 (N_6601,N_6584,N_6575);
xor U6602 (N_6602,N_6573,N_6545);
or U6603 (N_6603,N_6553,N_6547);
and U6604 (N_6604,N_6591,N_6518);
or U6605 (N_6605,N_6576,N_6512);
xnor U6606 (N_6606,N_6571,N_6552);
nor U6607 (N_6607,N_6505,N_6580);
or U6608 (N_6608,N_6517,N_6569);
or U6609 (N_6609,N_6581,N_6509);
or U6610 (N_6610,N_6550,N_6599);
and U6611 (N_6611,N_6589,N_6506);
and U6612 (N_6612,N_6527,N_6524);
nor U6613 (N_6613,N_6577,N_6574);
nor U6614 (N_6614,N_6536,N_6537);
nor U6615 (N_6615,N_6541,N_6525);
or U6616 (N_6616,N_6504,N_6508);
or U6617 (N_6617,N_6542,N_6500);
and U6618 (N_6618,N_6592,N_6523);
nor U6619 (N_6619,N_6521,N_6567);
nand U6620 (N_6620,N_6579,N_6554);
and U6621 (N_6621,N_6572,N_6560);
nor U6622 (N_6622,N_6526,N_6549);
nor U6623 (N_6623,N_6501,N_6532);
nand U6624 (N_6624,N_6558,N_6566);
nor U6625 (N_6625,N_6582,N_6511);
xnor U6626 (N_6626,N_6561,N_6551);
and U6627 (N_6627,N_6530,N_6503);
xor U6628 (N_6628,N_6516,N_6528);
nand U6629 (N_6629,N_6533,N_6564);
and U6630 (N_6630,N_6594,N_6548);
xor U6631 (N_6631,N_6529,N_6515);
and U6632 (N_6632,N_6543,N_6570);
nand U6633 (N_6633,N_6546,N_6502);
nand U6634 (N_6634,N_6520,N_6544);
and U6635 (N_6635,N_6519,N_6595);
nor U6636 (N_6636,N_6597,N_6565);
or U6637 (N_6637,N_6562,N_6510);
or U6638 (N_6638,N_6555,N_6540);
and U6639 (N_6639,N_6557,N_6507);
and U6640 (N_6640,N_6556,N_6522);
xor U6641 (N_6641,N_6538,N_6531);
xnor U6642 (N_6642,N_6590,N_6534);
nand U6643 (N_6643,N_6585,N_6568);
or U6644 (N_6644,N_6539,N_6587);
and U6645 (N_6645,N_6598,N_6588);
xor U6646 (N_6646,N_6578,N_6535);
xor U6647 (N_6647,N_6586,N_6514);
or U6648 (N_6648,N_6563,N_6593);
nand U6649 (N_6649,N_6596,N_6513);
nand U6650 (N_6650,N_6531,N_6584);
and U6651 (N_6651,N_6599,N_6597);
or U6652 (N_6652,N_6587,N_6542);
xor U6653 (N_6653,N_6520,N_6592);
and U6654 (N_6654,N_6590,N_6573);
nand U6655 (N_6655,N_6578,N_6528);
and U6656 (N_6656,N_6594,N_6561);
and U6657 (N_6657,N_6588,N_6572);
nor U6658 (N_6658,N_6514,N_6538);
or U6659 (N_6659,N_6543,N_6541);
nand U6660 (N_6660,N_6575,N_6567);
and U6661 (N_6661,N_6552,N_6516);
nor U6662 (N_6662,N_6543,N_6585);
xor U6663 (N_6663,N_6575,N_6553);
or U6664 (N_6664,N_6560,N_6507);
nor U6665 (N_6665,N_6534,N_6515);
or U6666 (N_6666,N_6572,N_6585);
and U6667 (N_6667,N_6584,N_6583);
and U6668 (N_6668,N_6550,N_6565);
nand U6669 (N_6669,N_6546,N_6515);
nor U6670 (N_6670,N_6565,N_6559);
xnor U6671 (N_6671,N_6595,N_6524);
nand U6672 (N_6672,N_6502,N_6590);
or U6673 (N_6673,N_6517,N_6589);
xor U6674 (N_6674,N_6592,N_6514);
nor U6675 (N_6675,N_6592,N_6509);
nand U6676 (N_6676,N_6546,N_6540);
nor U6677 (N_6677,N_6574,N_6554);
or U6678 (N_6678,N_6515,N_6590);
xor U6679 (N_6679,N_6564,N_6585);
nor U6680 (N_6680,N_6530,N_6555);
or U6681 (N_6681,N_6546,N_6590);
xor U6682 (N_6682,N_6592,N_6591);
nor U6683 (N_6683,N_6536,N_6598);
and U6684 (N_6684,N_6524,N_6522);
nor U6685 (N_6685,N_6598,N_6502);
and U6686 (N_6686,N_6534,N_6577);
nand U6687 (N_6687,N_6551,N_6515);
or U6688 (N_6688,N_6502,N_6531);
or U6689 (N_6689,N_6540,N_6598);
or U6690 (N_6690,N_6546,N_6533);
nand U6691 (N_6691,N_6509,N_6575);
or U6692 (N_6692,N_6537,N_6565);
xor U6693 (N_6693,N_6500,N_6560);
xor U6694 (N_6694,N_6589,N_6557);
nand U6695 (N_6695,N_6568,N_6583);
nor U6696 (N_6696,N_6559,N_6543);
nor U6697 (N_6697,N_6586,N_6504);
xor U6698 (N_6698,N_6542,N_6595);
nor U6699 (N_6699,N_6581,N_6560);
xor U6700 (N_6700,N_6672,N_6617);
or U6701 (N_6701,N_6698,N_6686);
xor U6702 (N_6702,N_6687,N_6625);
nor U6703 (N_6703,N_6654,N_6679);
xnor U6704 (N_6704,N_6604,N_6664);
and U6705 (N_6705,N_6606,N_6660);
nand U6706 (N_6706,N_6650,N_6661);
or U6707 (N_6707,N_6638,N_6683);
xor U6708 (N_6708,N_6697,N_6692);
xor U6709 (N_6709,N_6636,N_6674);
xnor U6710 (N_6710,N_6602,N_6612);
nand U6711 (N_6711,N_6631,N_6655);
nand U6712 (N_6712,N_6668,N_6622);
nor U6713 (N_6713,N_6643,N_6644);
nand U6714 (N_6714,N_6649,N_6680);
nor U6715 (N_6715,N_6632,N_6685);
or U6716 (N_6716,N_6699,N_6623);
nand U6717 (N_6717,N_6693,N_6663);
and U6718 (N_6718,N_6656,N_6611);
and U6719 (N_6719,N_6691,N_6616);
or U6720 (N_6720,N_6669,N_6653);
xor U6721 (N_6721,N_6648,N_6675);
or U6722 (N_6722,N_6629,N_6614);
nand U6723 (N_6723,N_6639,N_6609);
xnor U6724 (N_6724,N_6695,N_6677);
or U6725 (N_6725,N_6613,N_6601);
or U6726 (N_6726,N_6633,N_6682);
nand U6727 (N_6727,N_6667,N_6665);
nor U6728 (N_6728,N_6694,N_6630);
nor U6729 (N_6729,N_6626,N_6651);
and U6730 (N_6730,N_6657,N_6689);
or U6731 (N_6731,N_6607,N_6615);
or U6732 (N_6732,N_6658,N_6647);
or U6733 (N_6733,N_6659,N_6628);
nor U6734 (N_6734,N_6690,N_6642);
xor U6735 (N_6735,N_6635,N_6666);
or U6736 (N_6736,N_6671,N_6662);
and U6737 (N_6737,N_6641,N_6637);
nor U6738 (N_6738,N_6645,N_6646);
xnor U6739 (N_6739,N_6681,N_6673);
nor U6740 (N_6740,N_6608,N_6684);
or U6741 (N_6741,N_6605,N_6621);
or U6742 (N_6742,N_6634,N_6676);
nand U6743 (N_6743,N_6696,N_6610);
xor U6744 (N_6744,N_6688,N_6603);
xnor U6745 (N_6745,N_6600,N_6620);
xor U6746 (N_6746,N_6678,N_6670);
nand U6747 (N_6747,N_6619,N_6618);
and U6748 (N_6748,N_6624,N_6627);
or U6749 (N_6749,N_6652,N_6640);
xnor U6750 (N_6750,N_6678,N_6699);
nor U6751 (N_6751,N_6620,N_6606);
and U6752 (N_6752,N_6648,N_6606);
or U6753 (N_6753,N_6680,N_6671);
nand U6754 (N_6754,N_6600,N_6698);
nand U6755 (N_6755,N_6636,N_6618);
nand U6756 (N_6756,N_6686,N_6687);
and U6757 (N_6757,N_6645,N_6696);
or U6758 (N_6758,N_6602,N_6619);
or U6759 (N_6759,N_6617,N_6616);
nand U6760 (N_6760,N_6689,N_6646);
nor U6761 (N_6761,N_6677,N_6681);
and U6762 (N_6762,N_6619,N_6654);
nand U6763 (N_6763,N_6636,N_6689);
or U6764 (N_6764,N_6687,N_6601);
nor U6765 (N_6765,N_6634,N_6623);
xor U6766 (N_6766,N_6654,N_6637);
nor U6767 (N_6767,N_6667,N_6636);
or U6768 (N_6768,N_6647,N_6690);
nor U6769 (N_6769,N_6626,N_6658);
or U6770 (N_6770,N_6699,N_6690);
xnor U6771 (N_6771,N_6612,N_6643);
xnor U6772 (N_6772,N_6697,N_6631);
or U6773 (N_6773,N_6686,N_6616);
and U6774 (N_6774,N_6699,N_6650);
nand U6775 (N_6775,N_6682,N_6613);
or U6776 (N_6776,N_6649,N_6639);
nand U6777 (N_6777,N_6657,N_6605);
nor U6778 (N_6778,N_6661,N_6617);
nand U6779 (N_6779,N_6678,N_6689);
and U6780 (N_6780,N_6616,N_6645);
nand U6781 (N_6781,N_6671,N_6640);
nor U6782 (N_6782,N_6640,N_6661);
or U6783 (N_6783,N_6648,N_6626);
or U6784 (N_6784,N_6660,N_6699);
nor U6785 (N_6785,N_6655,N_6629);
nand U6786 (N_6786,N_6692,N_6684);
nand U6787 (N_6787,N_6615,N_6659);
xor U6788 (N_6788,N_6654,N_6625);
or U6789 (N_6789,N_6666,N_6680);
nand U6790 (N_6790,N_6612,N_6630);
xnor U6791 (N_6791,N_6613,N_6656);
xor U6792 (N_6792,N_6641,N_6638);
or U6793 (N_6793,N_6648,N_6678);
nand U6794 (N_6794,N_6696,N_6671);
and U6795 (N_6795,N_6668,N_6660);
nor U6796 (N_6796,N_6619,N_6622);
or U6797 (N_6797,N_6691,N_6600);
or U6798 (N_6798,N_6676,N_6604);
nor U6799 (N_6799,N_6649,N_6662);
nand U6800 (N_6800,N_6770,N_6799);
nand U6801 (N_6801,N_6793,N_6754);
nor U6802 (N_6802,N_6741,N_6796);
and U6803 (N_6803,N_6700,N_6753);
or U6804 (N_6804,N_6757,N_6731);
nor U6805 (N_6805,N_6751,N_6756);
nand U6806 (N_6806,N_6784,N_6727);
nand U6807 (N_6807,N_6742,N_6704);
and U6808 (N_6808,N_6766,N_6724);
nand U6809 (N_6809,N_6772,N_6735);
nor U6810 (N_6810,N_6738,N_6785);
and U6811 (N_6811,N_6733,N_6791);
or U6812 (N_6812,N_6759,N_6760);
xor U6813 (N_6813,N_6715,N_6712);
xnor U6814 (N_6814,N_6778,N_6774);
nor U6815 (N_6815,N_6737,N_6794);
and U6816 (N_6816,N_6714,N_6787);
nand U6817 (N_6817,N_6716,N_6747);
or U6818 (N_6818,N_6729,N_6706);
or U6819 (N_6819,N_6736,N_6788);
nor U6820 (N_6820,N_6797,N_6718);
xor U6821 (N_6821,N_6773,N_6728);
nand U6822 (N_6822,N_6744,N_6782);
nor U6823 (N_6823,N_6771,N_6775);
nor U6824 (N_6824,N_6798,N_6789);
xor U6825 (N_6825,N_6758,N_6732);
or U6826 (N_6826,N_6763,N_6764);
and U6827 (N_6827,N_6739,N_6786);
xnor U6828 (N_6828,N_6769,N_6730);
or U6829 (N_6829,N_6740,N_6709);
and U6830 (N_6830,N_6777,N_6795);
xnor U6831 (N_6831,N_6749,N_6767);
nor U6832 (N_6832,N_6721,N_6783);
xor U6833 (N_6833,N_6711,N_6743);
nor U6834 (N_6834,N_6726,N_6762);
xnor U6835 (N_6835,N_6768,N_6790);
nor U6836 (N_6836,N_6707,N_6710);
nand U6837 (N_6837,N_6713,N_6701);
nor U6838 (N_6838,N_6702,N_6746);
and U6839 (N_6839,N_6779,N_6780);
or U6840 (N_6840,N_6719,N_6705);
xor U6841 (N_6841,N_6750,N_6765);
or U6842 (N_6842,N_6755,N_6748);
xnor U6843 (N_6843,N_6734,N_6722);
xor U6844 (N_6844,N_6703,N_6781);
nor U6845 (N_6845,N_6720,N_6776);
xnor U6846 (N_6846,N_6708,N_6717);
nor U6847 (N_6847,N_6792,N_6761);
nand U6848 (N_6848,N_6752,N_6723);
nor U6849 (N_6849,N_6725,N_6745);
or U6850 (N_6850,N_6793,N_6700);
nor U6851 (N_6851,N_6744,N_6772);
or U6852 (N_6852,N_6712,N_6782);
nor U6853 (N_6853,N_6798,N_6724);
or U6854 (N_6854,N_6707,N_6768);
nor U6855 (N_6855,N_6776,N_6768);
nor U6856 (N_6856,N_6786,N_6776);
and U6857 (N_6857,N_6710,N_6726);
xnor U6858 (N_6858,N_6757,N_6780);
nor U6859 (N_6859,N_6731,N_6736);
xnor U6860 (N_6860,N_6744,N_6755);
and U6861 (N_6861,N_6762,N_6754);
or U6862 (N_6862,N_6764,N_6756);
or U6863 (N_6863,N_6721,N_6798);
or U6864 (N_6864,N_6778,N_6713);
nand U6865 (N_6865,N_6755,N_6751);
or U6866 (N_6866,N_6711,N_6768);
nand U6867 (N_6867,N_6775,N_6784);
and U6868 (N_6868,N_6752,N_6796);
or U6869 (N_6869,N_6752,N_6717);
nor U6870 (N_6870,N_6793,N_6798);
or U6871 (N_6871,N_6726,N_6711);
nand U6872 (N_6872,N_6744,N_6768);
xor U6873 (N_6873,N_6771,N_6702);
nand U6874 (N_6874,N_6733,N_6724);
nand U6875 (N_6875,N_6769,N_6786);
or U6876 (N_6876,N_6718,N_6757);
nor U6877 (N_6877,N_6748,N_6741);
xor U6878 (N_6878,N_6750,N_6712);
nor U6879 (N_6879,N_6761,N_6724);
or U6880 (N_6880,N_6718,N_6722);
nand U6881 (N_6881,N_6766,N_6733);
xnor U6882 (N_6882,N_6708,N_6726);
nor U6883 (N_6883,N_6724,N_6730);
and U6884 (N_6884,N_6772,N_6756);
xor U6885 (N_6885,N_6701,N_6789);
nand U6886 (N_6886,N_6777,N_6722);
nand U6887 (N_6887,N_6758,N_6708);
and U6888 (N_6888,N_6719,N_6763);
xnor U6889 (N_6889,N_6750,N_6786);
and U6890 (N_6890,N_6741,N_6782);
nor U6891 (N_6891,N_6733,N_6770);
and U6892 (N_6892,N_6712,N_6792);
or U6893 (N_6893,N_6782,N_6702);
or U6894 (N_6894,N_6750,N_6742);
nand U6895 (N_6895,N_6799,N_6773);
and U6896 (N_6896,N_6728,N_6789);
and U6897 (N_6897,N_6782,N_6750);
and U6898 (N_6898,N_6770,N_6786);
nand U6899 (N_6899,N_6713,N_6709);
xnor U6900 (N_6900,N_6872,N_6874);
or U6901 (N_6901,N_6811,N_6845);
xnor U6902 (N_6902,N_6856,N_6816);
nor U6903 (N_6903,N_6873,N_6863);
nand U6904 (N_6904,N_6878,N_6834);
or U6905 (N_6905,N_6896,N_6837);
nor U6906 (N_6906,N_6830,N_6846);
nand U6907 (N_6907,N_6836,N_6889);
or U6908 (N_6908,N_6871,N_6815);
nor U6909 (N_6909,N_6851,N_6875);
xor U6910 (N_6910,N_6849,N_6800);
nand U6911 (N_6911,N_6857,N_6805);
and U6912 (N_6912,N_6802,N_6801);
and U6913 (N_6913,N_6893,N_6828);
xnor U6914 (N_6914,N_6864,N_6854);
or U6915 (N_6915,N_6898,N_6861);
nor U6916 (N_6916,N_6825,N_6877);
nand U6917 (N_6917,N_6844,N_6819);
and U6918 (N_6918,N_6879,N_6897);
and U6919 (N_6919,N_6848,N_6804);
nor U6920 (N_6920,N_6894,N_6809);
and U6921 (N_6921,N_6826,N_6886);
and U6922 (N_6922,N_6899,N_6833);
xnor U6923 (N_6923,N_6890,N_6866);
nand U6924 (N_6924,N_6884,N_6852);
and U6925 (N_6925,N_6829,N_6859);
or U6926 (N_6926,N_6850,N_6827);
nand U6927 (N_6927,N_6832,N_6842);
nor U6928 (N_6928,N_6853,N_6862);
or U6929 (N_6929,N_6882,N_6812);
nor U6930 (N_6930,N_6835,N_6821);
xor U6931 (N_6931,N_6839,N_6888);
nand U6932 (N_6932,N_6808,N_6867);
and U6933 (N_6933,N_6807,N_6803);
and U6934 (N_6934,N_6814,N_6820);
and U6935 (N_6935,N_6869,N_6860);
nor U6936 (N_6936,N_6806,N_6865);
xor U6937 (N_6937,N_6881,N_6824);
or U6938 (N_6938,N_6847,N_6876);
nor U6939 (N_6939,N_6838,N_6831);
or U6940 (N_6940,N_6892,N_6841);
or U6941 (N_6941,N_6887,N_6883);
xor U6942 (N_6942,N_6810,N_6813);
xor U6943 (N_6943,N_6880,N_6843);
nor U6944 (N_6944,N_6870,N_6895);
or U6945 (N_6945,N_6891,N_6818);
and U6946 (N_6946,N_6885,N_6858);
nor U6947 (N_6947,N_6868,N_6855);
or U6948 (N_6948,N_6823,N_6822);
and U6949 (N_6949,N_6817,N_6840);
and U6950 (N_6950,N_6824,N_6879);
nor U6951 (N_6951,N_6836,N_6824);
and U6952 (N_6952,N_6839,N_6884);
nand U6953 (N_6953,N_6836,N_6821);
or U6954 (N_6954,N_6845,N_6820);
nor U6955 (N_6955,N_6898,N_6852);
xnor U6956 (N_6956,N_6811,N_6836);
and U6957 (N_6957,N_6895,N_6862);
and U6958 (N_6958,N_6846,N_6894);
xor U6959 (N_6959,N_6860,N_6884);
xnor U6960 (N_6960,N_6899,N_6883);
nor U6961 (N_6961,N_6861,N_6820);
or U6962 (N_6962,N_6852,N_6862);
nand U6963 (N_6963,N_6875,N_6822);
nor U6964 (N_6964,N_6844,N_6837);
and U6965 (N_6965,N_6811,N_6871);
nand U6966 (N_6966,N_6867,N_6804);
nor U6967 (N_6967,N_6896,N_6878);
and U6968 (N_6968,N_6884,N_6875);
xor U6969 (N_6969,N_6889,N_6878);
or U6970 (N_6970,N_6854,N_6891);
xor U6971 (N_6971,N_6865,N_6895);
and U6972 (N_6972,N_6826,N_6845);
and U6973 (N_6973,N_6833,N_6871);
nand U6974 (N_6974,N_6821,N_6873);
and U6975 (N_6975,N_6891,N_6805);
xnor U6976 (N_6976,N_6869,N_6833);
nand U6977 (N_6977,N_6868,N_6894);
nand U6978 (N_6978,N_6803,N_6827);
nand U6979 (N_6979,N_6815,N_6867);
and U6980 (N_6980,N_6896,N_6841);
nand U6981 (N_6981,N_6838,N_6858);
or U6982 (N_6982,N_6817,N_6823);
nor U6983 (N_6983,N_6808,N_6860);
nand U6984 (N_6984,N_6827,N_6805);
nor U6985 (N_6985,N_6815,N_6879);
nand U6986 (N_6986,N_6826,N_6857);
and U6987 (N_6987,N_6840,N_6898);
nor U6988 (N_6988,N_6896,N_6848);
and U6989 (N_6989,N_6847,N_6871);
or U6990 (N_6990,N_6818,N_6885);
or U6991 (N_6991,N_6847,N_6866);
and U6992 (N_6992,N_6807,N_6833);
nor U6993 (N_6993,N_6817,N_6837);
and U6994 (N_6994,N_6882,N_6820);
and U6995 (N_6995,N_6832,N_6874);
nor U6996 (N_6996,N_6833,N_6835);
nand U6997 (N_6997,N_6861,N_6816);
xor U6998 (N_6998,N_6857,N_6804);
or U6999 (N_6999,N_6899,N_6842);
xor U7000 (N_7000,N_6939,N_6931);
and U7001 (N_7001,N_6992,N_6907);
nand U7002 (N_7002,N_6984,N_6924);
or U7003 (N_7003,N_6941,N_6910);
xor U7004 (N_7004,N_6962,N_6999);
xnor U7005 (N_7005,N_6914,N_6912);
nand U7006 (N_7006,N_6927,N_6944);
or U7007 (N_7007,N_6951,N_6919);
or U7008 (N_7008,N_6903,N_6994);
and U7009 (N_7009,N_6916,N_6997);
xor U7010 (N_7010,N_6909,N_6996);
nand U7011 (N_7011,N_6929,N_6906);
or U7012 (N_7012,N_6982,N_6920);
nand U7013 (N_7013,N_6928,N_6945);
xor U7014 (N_7014,N_6993,N_6976);
nand U7015 (N_7015,N_6970,N_6926);
or U7016 (N_7016,N_6932,N_6900);
nand U7017 (N_7017,N_6956,N_6952);
xor U7018 (N_7018,N_6968,N_6987);
nor U7019 (N_7019,N_6953,N_6983);
or U7020 (N_7020,N_6960,N_6988);
nand U7021 (N_7021,N_6913,N_6985);
nor U7022 (N_7022,N_6957,N_6955);
or U7023 (N_7023,N_6973,N_6930);
nand U7024 (N_7024,N_6961,N_6998);
and U7025 (N_7025,N_6974,N_6989);
and U7026 (N_7026,N_6921,N_6978);
or U7027 (N_7027,N_6938,N_6971);
nand U7028 (N_7028,N_6925,N_6948);
and U7029 (N_7029,N_6943,N_6991);
nand U7030 (N_7030,N_6986,N_6964);
or U7031 (N_7031,N_6990,N_6947);
and U7032 (N_7032,N_6915,N_6908);
and U7033 (N_7033,N_6933,N_6922);
nand U7034 (N_7034,N_6901,N_6979);
xor U7035 (N_7035,N_6936,N_6965);
or U7036 (N_7036,N_6966,N_6977);
or U7037 (N_7037,N_6950,N_6911);
xor U7038 (N_7038,N_6963,N_6942);
nand U7039 (N_7039,N_6904,N_6967);
xor U7040 (N_7040,N_6917,N_6969);
and U7041 (N_7041,N_6958,N_6980);
xnor U7042 (N_7042,N_6923,N_6972);
or U7043 (N_7043,N_6905,N_6902);
nand U7044 (N_7044,N_6918,N_6934);
nand U7045 (N_7045,N_6940,N_6981);
or U7046 (N_7046,N_6949,N_6946);
or U7047 (N_7047,N_6995,N_6954);
nand U7048 (N_7048,N_6937,N_6959);
xor U7049 (N_7049,N_6935,N_6975);
and U7050 (N_7050,N_6951,N_6916);
and U7051 (N_7051,N_6901,N_6933);
and U7052 (N_7052,N_6942,N_6971);
and U7053 (N_7053,N_6944,N_6921);
nor U7054 (N_7054,N_6995,N_6918);
and U7055 (N_7055,N_6924,N_6918);
or U7056 (N_7056,N_6968,N_6925);
or U7057 (N_7057,N_6998,N_6965);
nor U7058 (N_7058,N_6997,N_6975);
or U7059 (N_7059,N_6915,N_6927);
or U7060 (N_7060,N_6905,N_6955);
nand U7061 (N_7061,N_6900,N_6950);
and U7062 (N_7062,N_6904,N_6978);
or U7063 (N_7063,N_6974,N_6930);
nand U7064 (N_7064,N_6944,N_6916);
xor U7065 (N_7065,N_6917,N_6993);
nor U7066 (N_7066,N_6957,N_6968);
xor U7067 (N_7067,N_6966,N_6950);
and U7068 (N_7068,N_6964,N_6925);
nor U7069 (N_7069,N_6936,N_6979);
and U7070 (N_7070,N_6943,N_6997);
and U7071 (N_7071,N_6989,N_6924);
and U7072 (N_7072,N_6969,N_6939);
nand U7073 (N_7073,N_6975,N_6926);
nand U7074 (N_7074,N_6966,N_6984);
nor U7075 (N_7075,N_6948,N_6994);
nand U7076 (N_7076,N_6956,N_6969);
and U7077 (N_7077,N_6976,N_6943);
or U7078 (N_7078,N_6998,N_6912);
and U7079 (N_7079,N_6902,N_6985);
and U7080 (N_7080,N_6997,N_6955);
nand U7081 (N_7081,N_6913,N_6924);
nand U7082 (N_7082,N_6961,N_6952);
xnor U7083 (N_7083,N_6902,N_6934);
and U7084 (N_7084,N_6938,N_6939);
nor U7085 (N_7085,N_6966,N_6988);
and U7086 (N_7086,N_6921,N_6949);
xor U7087 (N_7087,N_6935,N_6998);
nor U7088 (N_7088,N_6976,N_6961);
and U7089 (N_7089,N_6963,N_6955);
and U7090 (N_7090,N_6959,N_6970);
nand U7091 (N_7091,N_6972,N_6909);
xnor U7092 (N_7092,N_6938,N_6950);
or U7093 (N_7093,N_6955,N_6983);
nor U7094 (N_7094,N_6946,N_6980);
xnor U7095 (N_7095,N_6906,N_6984);
nor U7096 (N_7096,N_6981,N_6915);
nand U7097 (N_7097,N_6989,N_6949);
nor U7098 (N_7098,N_6984,N_6990);
or U7099 (N_7099,N_6924,N_6917);
nor U7100 (N_7100,N_7095,N_7007);
xnor U7101 (N_7101,N_7070,N_7049);
nor U7102 (N_7102,N_7023,N_7067);
xor U7103 (N_7103,N_7056,N_7071);
nor U7104 (N_7104,N_7047,N_7036);
nor U7105 (N_7105,N_7074,N_7064);
nor U7106 (N_7106,N_7082,N_7024);
or U7107 (N_7107,N_7030,N_7093);
nand U7108 (N_7108,N_7099,N_7014);
xor U7109 (N_7109,N_7018,N_7044);
or U7110 (N_7110,N_7065,N_7001);
nor U7111 (N_7111,N_7059,N_7045);
nand U7112 (N_7112,N_7084,N_7069);
nand U7113 (N_7113,N_7000,N_7010);
and U7114 (N_7114,N_7090,N_7072);
nand U7115 (N_7115,N_7083,N_7080);
nor U7116 (N_7116,N_7038,N_7012);
and U7117 (N_7117,N_7068,N_7089);
or U7118 (N_7118,N_7011,N_7091);
nor U7119 (N_7119,N_7022,N_7031);
xnor U7120 (N_7120,N_7061,N_7042);
and U7121 (N_7121,N_7027,N_7035);
nand U7122 (N_7122,N_7092,N_7097);
xnor U7123 (N_7123,N_7015,N_7087);
nor U7124 (N_7124,N_7094,N_7078);
nand U7125 (N_7125,N_7017,N_7004);
nand U7126 (N_7126,N_7002,N_7021);
nor U7127 (N_7127,N_7073,N_7009);
nand U7128 (N_7128,N_7052,N_7066);
nor U7129 (N_7129,N_7062,N_7028);
nand U7130 (N_7130,N_7060,N_7050);
or U7131 (N_7131,N_7046,N_7075);
nor U7132 (N_7132,N_7088,N_7016);
nor U7133 (N_7133,N_7039,N_7057);
nand U7134 (N_7134,N_7013,N_7077);
nand U7135 (N_7135,N_7041,N_7008);
nor U7136 (N_7136,N_7076,N_7033);
and U7137 (N_7137,N_7081,N_7006);
nor U7138 (N_7138,N_7040,N_7096);
nor U7139 (N_7139,N_7051,N_7058);
and U7140 (N_7140,N_7098,N_7005);
xor U7141 (N_7141,N_7020,N_7037);
xnor U7142 (N_7142,N_7025,N_7053);
or U7143 (N_7143,N_7034,N_7055);
xnor U7144 (N_7144,N_7086,N_7026);
nor U7145 (N_7145,N_7048,N_7079);
xor U7146 (N_7146,N_7054,N_7032);
and U7147 (N_7147,N_7003,N_7029);
or U7148 (N_7148,N_7063,N_7043);
xnor U7149 (N_7149,N_7085,N_7019);
or U7150 (N_7150,N_7069,N_7037);
nand U7151 (N_7151,N_7092,N_7096);
or U7152 (N_7152,N_7010,N_7089);
nor U7153 (N_7153,N_7016,N_7004);
and U7154 (N_7154,N_7070,N_7089);
and U7155 (N_7155,N_7004,N_7001);
and U7156 (N_7156,N_7048,N_7002);
or U7157 (N_7157,N_7048,N_7052);
or U7158 (N_7158,N_7068,N_7012);
nand U7159 (N_7159,N_7089,N_7074);
and U7160 (N_7160,N_7084,N_7055);
nand U7161 (N_7161,N_7070,N_7011);
or U7162 (N_7162,N_7020,N_7048);
nor U7163 (N_7163,N_7077,N_7072);
or U7164 (N_7164,N_7004,N_7064);
nand U7165 (N_7165,N_7078,N_7004);
or U7166 (N_7166,N_7036,N_7081);
or U7167 (N_7167,N_7048,N_7005);
nand U7168 (N_7168,N_7050,N_7089);
and U7169 (N_7169,N_7039,N_7066);
and U7170 (N_7170,N_7086,N_7083);
and U7171 (N_7171,N_7049,N_7050);
nand U7172 (N_7172,N_7060,N_7057);
nor U7173 (N_7173,N_7061,N_7063);
and U7174 (N_7174,N_7088,N_7023);
and U7175 (N_7175,N_7091,N_7075);
xnor U7176 (N_7176,N_7039,N_7016);
nand U7177 (N_7177,N_7056,N_7085);
xor U7178 (N_7178,N_7084,N_7001);
nand U7179 (N_7179,N_7032,N_7089);
and U7180 (N_7180,N_7035,N_7029);
xnor U7181 (N_7181,N_7057,N_7070);
nor U7182 (N_7182,N_7089,N_7062);
nand U7183 (N_7183,N_7086,N_7016);
xor U7184 (N_7184,N_7037,N_7084);
and U7185 (N_7185,N_7070,N_7027);
nor U7186 (N_7186,N_7095,N_7046);
nor U7187 (N_7187,N_7091,N_7085);
or U7188 (N_7188,N_7053,N_7073);
nand U7189 (N_7189,N_7052,N_7091);
nor U7190 (N_7190,N_7026,N_7074);
nor U7191 (N_7191,N_7047,N_7066);
and U7192 (N_7192,N_7083,N_7091);
xor U7193 (N_7193,N_7041,N_7020);
and U7194 (N_7194,N_7074,N_7044);
nor U7195 (N_7195,N_7057,N_7028);
nand U7196 (N_7196,N_7051,N_7048);
nand U7197 (N_7197,N_7081,N_7039);
nor U7198 (N_7198,N_7090,N_7045);
or U7199 (N_7199,N_7015,N_7059);
nor U7200 (N_7200,N_7114,N_7185);
xnor U7201 (N_7201,N_7130,N_7165);
nor U7202 (N_7202,N_7134,N_7148);
xnor U7203 (N_7203,N_7124,N_7162);
nand U7204 (N_7204,N_7167,N_7146);
and U7205 (N_7205,N_7166,N_7192);
nor U7206 (N_7206,N_7173,N_7110);
nand U7207 (N_7207,N_7193,N_7199);
and U7208 (N_7208,N_7106,N_7109);
xor U7209 (N_7209,N_7133,N_7153);
and U7210 (N_7210,N_7126,N_7170);
xor U7211 (N_7211,N_7150,N_7151);
xnor U7212 (N_7212,N_7178,N_7122);
and U7213 (N_7213,N_7132,N_7147);
nor U7214 (N_7214,N_7190,N_7188);
or U7215 (N_7215,N_7176,N_7136);
nand U7216 (N_7216,N_7100,N_7197);
xnor U7217 (N_7217,N_7112,N_7142);
or U7218 (N_7218,N_7120,N_7108);
xor U7219 (N_7219,N_7118,N_7160);
or U7220 (N_7220,N_7154,N_7104);
and U7221 (N_7221,N_7117,N_7129);
nand U7222 (N_7222,N_7181,N_7179);
nor U7223 (N_7223,N_7182,N_7135);
or U7224 (N_7224,N_7116,N_7159);
xor U7225 (N_7225,N_7164,N_7198);
nor U7226 (N_7226,N_7140,N_7158);
xor U7227 (N_7227,N_7113,N_7189);
xnor U7228 (N_7228,N_7177,N_7152);
nand U7229 (N_7229,N_7161,N_7128);
nor U7230 (N_7230,N_7107,N_7111);
nor U7231 (N_7231,N_7169,N_7195);
nor U7232 (N_7232,N_7105,N_7157);
and U7233 (N_7233,N_7174,N_7180);
nand U7234 (N_7234,N_7143,N_7187);
nor U7235 (N_7235,N_7115,N_7123);
or U7236 (N_7236,N_7141,N_7145);
and U7237 (N_7237,N_7101,N_7137);
xor U7238 (N_7238,N_7144,N_7184);
xor U7239 (N_7239,N_7125,N_7172);
and U7240 (N_7240,N_7156,N_7102);
nor U7241 (N_7241,N_7163,N_7196);
nand U7242 (N_7242,N_7119,N_7121);
and U7243 (N_7243,N_7194,N_7103);
or U7244 (N_7244,N_7168,N_7149);
and U7245 (N_7245,N_7127,N_7139);
or U7246 (N_7246,N_7131,N_7191);
nand U7247 (N_7247,N_7155,N_7138);
or U7248 (N_7248,N_7186,N_7183);
or U7249 (N_7249,N_7171,N_7175);
nor U7250 (N_7250,N_7120,N_7173);
nor U7251 (N_7251,N_7120,N_7100);
or U7252 (N_7252,N_7176,N_7134);
nor U7253 (N_7253,N_7152,N_7119);
and U7254 (N_7254,N_7103,N_7187);
nand U7255 (N_7255,N_7130,N_7173);
xnor U7256 (N_7256,N_7153,N_7170);
nor U7257 (N_7257,N_7118,N_7152);
or U7258 (N_7258,N_7176,N_7123);
nor U7259 (N_7259,N_7186,N_7120);
and U7260 (N_7260,N_7100,N_7135);
nand U7261 (N_7261,N_7156,N_7152);
and U7262 (N_7262,N_7126,N_7148);
or U7263 (N_7263,N_7171,N_7141);
and U7264 (N_7264,N_7195,N_7138);
or U7265 (N_7265,N_7181,N_7161);
nand U7266 (N_7266,N_7107,N_7199);
nand U7267 (N_7267,N_7174,N_7168);
nor U7268 (N_7268,N_7103,N_7126);
and U7269 (N_7269,N_7109,N_7185);
and U7270 (N_7270,N_7165,N_7171);
and U7271 (N_7271,N_7195,N_7187);
nand U7272 (N_7272,N_7193,N_7147);
xor U7273 (N_7273,N_7138,N_7110);
and U7274 (N_7274,N_7149,N_7104);
nor U7275 (N_7275,N_7187,N_7138);
or U7276 (N_7276,N_7114,N_7174);
nand U7277 (N_7277,N_7154,N_7153);
xor U7278 (N_7278,N_7116,N_7161);
or U7279 (N_7279,N_7113,N_7174);
and U7280 (N_7280,N_7199,N_7164);
or U7281 (N_7281,N_7196,N_7110);
nor U7282 (N_7282,N_7129,N_7180);
xor U7283 (N_7283,N_7150,N_7189);
nand U7284 (N_7284,N_7107,N_7106);
or U7285 (N_7285,N_7159,N_7131);
xor U7286 (N_7286,N_7110,N_7163);
and U7287 (N_7287,N_7125,N_7164);
nand U7288 (N_7288,N_7167,N_7114);
or U7289 (N_7289,N_7146,N_7147);
nor U7290 (N_7290,N_7186,N_7194);
nor U7291 (N_7291,N_7191,N_7144);
nand U7292 (N_7292,N_7198,N_7192);
or U7293 (N_7293,N_7194,N_7174);
and U7294 (N_7294,N_7106,N_7168);
or U7295 (N_7295,N_7154,N_7174);
and U7296 (N_7296,N_7167,N_7126);
nand U7297 (N_7297,N_7102,N_7186);
xor U7298 (N_7298,N_7167,N_7137);
or U7299 (N_7299,N_7157,N_7148);
nor U7300 (N_7300,N_7247,N_7222);
xnor U7301 (N_7301,N_7233,N_7254);
or U7302 (N_7302,N_7266,N_7231);
nand U7303 (N_7303,N_7273,N_7215);
xor U7304 (N_7304,N_7223,N_7229);
or U7305 (N_7305,N_7232,N_7253);
nor U7306 (N_7306,N_7256,N_7275);
nand U7307 (N_7307,N_7200,N_7262);
and U7308 (N_7308,N_7226,N_7267);
nor U7309 (N_7309,N_7241,N_7201);
xnor U7310 (N_7310,N_7276,N_7290);
nor U7311 (N_7311,N_7249,N_7242);
nor U7312 (N_7312,N_7280,N_7292);
nand U7313 (N_7313,N_7296,N_7207);
nor U7314 (N_7314,N_7206,N_7295);
nor U7315 (N_7315,N_7228,N_7208);
or U7316 (N_7316,N_7244,N_7205);
nor U7317 (N_7317,N_7283,N_7211);
and U7318 (N_7318,N_7219,N_7218);
nand U7319 (N_7319,N_7216,N_7245);
nor U7320 (N_7320,N_7214,N_7261);
xnor U7321 (N_7321,N_7237,N_7299);
xor U7322 (N_7322,N_7271,N_7264);
or U7323 (N_7323,N_7250,N_7285);
nor U7324 (N_7324,N_7236,N_7281);
xor U7325 (N_7325,N_7204,N_7212);
or U7326 (N_7326,N_7202,N_7243);
nand U7327 (N_7327,N_7210,N_7260);
xnor U7328 (N_7328,N_7230,N_7217);
nor U7329 (N_7329,N_7203,N_7272);
nand U7330 (N_7330,N_7259,N_7252);
nor U7331 (N_7331,N_7297,N_7224);
nand U7332 (N_7332,N_7277,N_7234);
nor U7333 (N_7333,N_7289,N_7221);
and U7334 (N_7334,N_7287,N_7258);
xnor U7335 (N_7335,N_7298,N_7269);
xnor U7336 (N_7336,N_7220,N_7238);
xnor U7337 (N_7337,N_7240,N_7278);
nand U7338 (N_7338,N_7257,N_7291);
xor U7339 (N_7339,N_7265,N_7282);
or U7340 (N_7340,N_7209,N_7246);
nand U7341 (N_7341,N_7274,N_7255);
nor U7342 (N_7342,N_7263,N_7286);
nand U7343 (N_7343,N_7225,N_7288);
nand U7344 (N_7344,N_7270,N_7279);
nor U7345 (N_7345,N_7293,N_7268);
or U7346 (N_7346,N_7284,N_7251);
and U7347 (N_7347,N_7227,N_7248);
or U7348 (N_7348,N_7294,N_7235);
xnor U7349 (N_7349,N_7239,N_7213);
nand U7350 (N_7350,N_7265,N_7217);
and U7351 (N_7351,N_7249,N_7209);
and U7352 (N_7352,N_7202,N_7236);
xor U7353 (N_7353,N_7234,N_7250);
xnor U7354 (N_7354,N_7238,N_7208);
and U7355 (N_7355,N_7218,N_7210);
and U7356 (N_7356,N_7241,N_7291);
or U7357 (N_7357,N_7274,N_7258);
or U7358 (N_7358,N_7217,N_7251);
xor U7359 (N_7359,N_7216,N_7249);
and U7360 (N_7360,N_7296,N_7271);
and U7361 (N_7361,N_7234,N_7214);
nand U7362 (N_7362,N_7267,N_7229);
or U7363 (N_7363,N_7259,N_7219);
nand U7364 (N_7364,N_7230,N_7297);
and U7365 (N_7365,N_7292,N_7278);
xor U7366 (N_7366,N_7251,N_7287);
nor U7367 (N_7367,N_7222,N_7289);
xor U7368 (N_7368,N_7294,N_7216);
nor U7369 (N_7369,N_7288,N_7264);
nand U7370 (N_7370,N_7209,N_7289);
nand U7371 (N_7371,N_7282,N_7286);
xor U7372 (N_7372,N_7217,N_7209);
or U7373 (N_7373,N_7221,N_7252);
and U7374 (N_7374,N_7207,N_7225);
and U7375 (N_7375,N_7255,N_7209);
xnor U7376 (N_7376,N_7278,N_7296);
xor U7377 (N_7377,N_7231,N_7285);
xnor U7378 (N_7378,N_7242,N_7227);
nand U7379 (N_7379,N_7206,N_7220);
xor U7380 (N_7380,N_7201,N_7295);
xor U7381 (N_7381,N_7240,N_7230);
nand U7382 (N_7382,N_7287,N_7220);
or U7383 (N_7383,N_7263,N_7230);
nand U7384 (N_7384,N_7290,N_7273);
xnor U7385 (N_7385,N_7234,N_7289);
and U7386 (N_7386,N_7293,N_7275);
xnor U7387 (N_7387,N_7283,N_7247);
nand U7388 (N_7388,N_7279,N_7268);
or U7389 (N_7389,N_7218,N_7299);
and U7390 (N_7390,N_7259,N_7285);
or U7391 (N_7391,N_7218,N_7221);
nor U7392 (N_7392,N_7277,N_7263);
nand U7393 (N_7393,N_7284,N_7224);
nor U7394 (N_7394,N_7244,N_7255);
xor U7395 (N_7395,N_7253,N_7261);
nor U7396 (N_7396,N_7201,N_7217);
nor U7397 (N_7397,N_7252,N_7287);
and U7398 (N_7398,N_7290,N_7244);
or U7399 (N_7399,N_7258,N_7296);
xor U7400 (N_7400,N_7314,N_7323);
xnor U7401 (N_7401,N_7343,N_7380);
nand U7402 (N_7402,N_7344,N_7307);
nand U7403 (N_7403,N_7389,N_7337);
nor U7404 (N_7404,N_7356,N_7348);
nor U7405 (N_7405,N_7368,N_7341);
or U7406 (N_7406,N_7321,N_7396);
nor U7407 (N_7407,N_7340,N_7386);
nor U7408 (N_7408,N_7339,N_7399);
nor U7409 (N_7409,N_7303,N_7319);
and U7410 (N_7410,N_7375,N_7354);
nand U7411 (N_7411,N_7349,N_7304);
or U7412 (N_7412,N_7373,N_7350);
or U7413 (N_7413,N_7359,N_7301);
nor U7414 (N_7414,N_7391,N_7338);
and U7415 (N_7415,N_7342,N_7312);
or U7416 (N_7416,N_7327,N_7300);
and U7417 (N_7417,N_7315,N_7384);
xor U7418 (N_7418,N_7346,N_7385);
or U7419 (N_7419,N_7362,N_7328);
and U7420 (N_7420,N_7325,N_7320);
and U7421 (N_7421,N_7397,N_7372);
and U7422 (N_7422,N_7318,N_7376);
xor U7423 (N_7423,N_7379,N_7365);
and U7424 (N_7424,N_7398,N_7329);
and U7425 (N_7425,N_7322,N_7358);
nor U7426 (N_7426,N_7351,N_7324);
nor U7427 (N_7427,N_7311,N_7367);
or U7428 (N_7428,N_7394,N_7305);
and U7429 (N_7429,N_7395,N_7302);
or U7430 (N_7430,N_7333,N_7313);
and U7431 (N_7431,N_7317,N_7352);
nand U7432 (N_7432,N_7371,N_7355);
nand U7433 (N_7433,N_7336,N_7363);
and U7434 (N_7434,N_7374,N_7332);
and U7435 (N_7435,N_7387,N_7326);
xor U7436 (N_7436,N_7383,N_7364);
and U7437 (N_7437,N_7309,N_7330);
xnor U7438 (N_7438,N_7382,N_7360);
nand U7439 (N_7439,N_7357,N_7366);
xnor U7440 (N_7440,N_7310,N_7369);
nor U7441 (N_7441,N_7347,N_7361);
or U7442 (N_7442,N_7331,N_7392);
or U7443 (N_7443,N_7353,N_7377);
nor U7444 (N_7444,N_7381,N_7370);
nand U7445 (N_7445,N_7316,N_7306);
and U7446 (N_7446,N_7388,N_7308);
or U7447 (N_7447,N_7334,N_7378);
or U7448 (N_7448,N_7345,N_7393);
and U7449 (N_7449,N_7335,N_7390);
nand U7450 (N_7450,N_7329,N_7380);
or U7451 (N_7451,N_7342,N_7330);
or U7452 (N_7452,N_7324,N_7393);
xor U7453 (N_7453,N_7302,N_7370);
nand U7454 (N_7454,N_7327,N_7372);
or U7455 (N_7455,N_7303,N_7378);
nand U7456 (N_7456,N_7396,N_7365);
or U7457 (N_7457,N_7334,N_7370);
xnor U7458 (N_7458,N_7316,N_7395);
or U7459 (N_7459,N_7387,N_7300);
nand U7460 (N_7460,N_7367,N_7307);
nor U7461 (N_7461,N_7335,N_7333);
nand U7462 (N_7462,N_7314,N_7328);
and U7463 (N_7463,N_7375,N_7370);
nor U7464 (N_7464,N_7320,N_7313);
xor U7465 (N_7465,N_7384,N_7391);
nor U7466 (N_7466,N_7391,N_7399);
nor U7467 (N_7467,N_7395,N_7338);
nor U7468 (N_7468,N_7395,N_7375);
xnor U7469 (N_7469,N_7321,N_7337);
xor U7470 (N_7470,N_7312,N_7375);
or U7471 (N_7471,N_7326,N_7360);
nor U7472 (N_7472,N_7387,N_7310);
nand U7473 (N_7473,N_7358,N_7372);
xor U7474 (N_7474,N_7336,N_7323);
nand U7475 (N_7475,N_7383,N_7389);
and U7476 (N_7476,N_7376,N_7378);
xor U7477 (N_7477,N_7302,N_7371);
nor U7478 (N_7478,N_7344,N_7354);
nand U7479 (N_7479,N_7308,N_7306);
or U7480 (N_7480,N_7341,N_7303);
nor U7481 (N_7481,N_7307,N_7334);
nand U7482 (N_7482,N_7369,N_7359);
and U7483 (N_7483,N_7371,N_7368);
and U7484 (N_7484,N_7366,N_7396);
and U7485 (N_7485,N_7383,N_7395);
and U7486 (N_7486,N_7386,N_7351);
nor U7487 (N_7487,N_7334,N_7396);
or U7488 (N_7488,N_7303,N_7323);
nor U7489 (N_7489,N_7342,N_7313);
xor U7490 (N_7490,N_7362,N_7342);
nor U7491 (N_7491,N_7381,N_7391);
nor U7492 (N_7492,N_7364,N_7303);
nor U7493 (N_7493,N_7325,N_7336);
or U7494 (N_7494,N_7312,N_7346);
and U7495 (N_7495,N_7351,N_7335);
xor U7496 (N_7496,N_7324,N_7348);
nor U7497 (N_7497,N_7369,N_7306);
nor U7498 (N_7498,N_7359,N_7339);
and U7499 (N_7499,N_7372,N_7342);
nor U7500 (N_7500,N_7495,N_7403);
nand U7501 (N_7501,N_7446,N_7427);
nor U7502 (N_7502,N_7431,N_7473);
nand U7503 (N_7503,N_7496,N_7406);
or U7504 (N_7504,N_7490,N_7408);
xor U7505 (N_7505,N_7443,N_7488);
or U7506 (N_7506,N_7428,N_7438);
nand U7507 (N_7507,N_7480,N_7441);
nand U7508 (N_7508,N_7453,N_7445);
and U7509 (N_7509,N_7412,N_7461);
and U7510 (N_7510,N_7489,N_7484);
and U7511 (N_7511,N_7414,N_7458);
nand U7512 (N_7512,N_7454,N_7474);
nor U7513 (N_7513,N_7486,N_7432);
xnor U7514 (N_7514,N_7404,N_7485);
and U7515 (N_7515,N_7491,N_7426);
xor U7516 (N_7516,N_7421,N_7457);
nand U7517 (N_7517,N_7465,N_7482);
nor U7518 (N_7518,N_7471,N_7402);
and U7519 (N_7519,N_7459,N_7440);
xor U7520 (N_7520,N_7475,N_7429);
or U7521 (N_7521,N_7472,N_7477);
nor U7522 (N_7522,N_7407,N_7444);
or U7523 (N_7523,N_7411,N_7483);
xnor U7524 (N_7524,N_7456,N_7478);
nand U7525 (N_7525,N_7499,N_7467);
or U7526 (N_7526,N_7413,N_7436);
or U7527 (N_7527,N_7423,N_7410);
xor U7528 (N_7528,N_7401,N_7425);
nor U7529 (N_7529,N_7400,N_7447);
and U7530 (N_7530,N_7435,N_7434);
and U7531 (N_7531,N_7498,N_7466);
nor U7532 (N_7532,N_7417,N_7437);
and U7533 (N_7533,N_7430,N_7415);
nor U7534 (N_7534,N_7424,N_7468);
nand U7535 (N_7535,N_7476,N_7481);
and U7536 (N_7536,N_7492,N_7442);
nor U7537 (N_7537,N_7420,N_7452);
or U7538 (N_7538,N_7455,N_7463);
or U7539 (N_7539,N_7493,N_7462);
nand U7540 (N_7540,N_7419,N_7494);
nand U7541 (N_7541,N_7422,N_7409);
or U7542 (N_7542,N_7464,N_7450);
and U7543 (N_7543,N_7418,N_7470);
or U7544 (N_7544,N_7487,N_7416);
or U7545 (N_7545,N_7451,N_7449);
xor U7546 (N_7546,N_7448,N_7479);
nor U7547 (N_7547,N_7469,N_7460);
nand U7548 (N_7548,N_7497,N_7405);
and U7549 (N_7549,N_7433,N_7439);
nor U7550 (N_7550,N_7490,N_7471);
nand U7551 (N_7551,N_7494,N_7468);
nand U7552 (N_7552,N_7431,N_7459);
nor U7553 (N_7553,N_7474,N_7477);
nand U7554 (N_7554,N_7488,N_7440);
and U7555 (N_7555,N_7492,N_7403);
and U7556 (N_7556,N_7429,N_7419);
nand U7557 (N_7557,N_7470,N_7456);
xor U7558 (N_7558,N_7495,N_7438);
nand U7559 (N_7559,N_7400,N_7418);
nor U7560 (N_7560,N_7416,N_7452);
and U7561 (N_7561,N_7463,N_7415);
nand U7562 (N_7562,N_7445,N_7479);
nand U7563 (N_7563,N_7436,N_7469);
or U7564 (N_7564,N_7432,N_7489);
or U7565 (N_7565,N_7499,N_7466);
nand U7566 (N_7566,N_7411,N_7432);
nor U7567 (N_7567,N_7463,N_7468);
and U7568 (N_7568,N_7442,N_7458);
xor U7569 (N_7569,N_7463,N_7459);
or U7570 (N_7570,N_7485,N_7442);
or U7571 (N_7571,N_7453,N_7446);
and U7572 (N_7572,N_7486,N_7488);
and U7573 (N_7573,N_7493,N_7451);
nor U7574 (N_7574,N_7464,N_7493);
nor U7575 (N_7575,N_7498,N_7449);
nand U7576 (N_7576,N_7468,N_7420);
xnor U7577 (N_7577,N_7435,N_7466);
xnor U7578 (N_7578,N_7467,N_7423);
and U7579 (N_7579,N_7412,N_7411);
nor U7580 (N_7580,N_7473,N_7466);
xnor U7581 (N_7581,N_7495,N_7428);
and U7582 (N_7582,N_7472,N_7440);
xnor U7583 (N_7583,N_7420,N_7427);
or U7584 (N_7584,N_7425,N_7448);
nand U7585 (N_7585,N_7431,N_7464);
nand U7586 (N_7586,N_7408,N_7412);
nor U7587 (N_7587,N_7484,N_7459);
xnor U7588 (N_7588,N_7453,N_7431);
nand U7589 (N_7589,N_7436,N_7404);
and U7590 (N_7590,N_7499,N_7427);
and U7591 (N_7591,N_7456,N_7458);
nand U7592 (N_7592,N_7464,N_7496);
and U7593 (N_7593,N_7418,N_7413);
or U7594 (N_7594,N_7409,N_7489);
xnor U7595 (N_7595,N_7424,N_7498);
nor U7596 (N_7596,N_7442,N_7403);
or U7597 (N_7597,N_7429,N_7476);
nor U7598 (N_7598,N_7496,N_7417);
nor U7599 (N_7599,N_7451,N_7413);
xnor U7600 (N_7600,N_7522,N_7592);
nand U7601 (N_7601,N_7562,N_7558);
nor U7602 (N_7602,N_7550,N_7552);
nand U7603 (N_7603,N_7544,N_7517);
nor U7604 (N_7604,N_7593,N_7508);
xnor U7605 (N_7605,N_7513,N_7501);
or U7606 (N_7606,N_7524,N_7541);
nor U7607 (N_7607,N_7526,N_7539);
xor U7608 (N_7608,N_7565,N_7520);
xor U7609 (N_7609,N_7530,N_7540);
or U7610 (N_7610,N_7590,N_7597);
and U7611 (N_7611,N_7563,N_7545);
nor U7612 (N_7612,N_7532,N_7512);
or U7613 (N_7613,N_7560,N_7571);
nand U7614 (N_7614,N_7500,N_7583);
nand U7615 (N_7615,N_7591,N_7564);
and U7616 (N_7616,N_7510,N_7575);
nor U7617 (N_7617,N_7599,N_7503);
and U7618 (N_7618,N_7548,N_7594);
xor U7619 (N_7619,N_7523,N_7557);
xor U7620 (N_7620,N_7506,N_7574);
and U7621 (N_7621,N_7515,N_7525);
xnor U7622 (N_7622,N_7509,N_7598);
and U7623 (N_7623,N_7568,N_7578);
xnor U7624 (N_7624,N_7569,N_7549);
and U7625 (N_7625,N_7561,N_7519);
and U7626 (N_7626,N_7596,N_7589);
xnor U7627 (N_7627,N_7538,N_7582);
or U7628 (N_7628,N_7547,N_7585);
nor U7629 (N_7629,N_7531,N_7554);
and U7630 (N_7630,N_7505,N_7546);
and U7631 (N_7631,N_7559,N_7588);
xnor U7632 (N_7632,N_7536,N_7521);
xnor U7633 (N_7633,N_7504,N_7543);
and U7634 (N_7634,N_7518,N_7586);
and U7635 (N_7635,N_7553,N_7570);
and U7636 (N_7636,N_7584,N_7551);
nor U7637 (N_7637,N_7537,N_7577);
xor U7638 (N_7638,N_7587,N_7555);
or U7639 (N_7639,N_7573,N_7527);
nand U7640 (N_7640,N_7511,N_7528);
and U7641 (N_7641,N_7534,N_7581);
nand U7642 (N_7642,N_7556,N_7576);
nor U7643 (N_7643,N_7516,N_7566);
and U7644 (N_7644,N_7529,N_7567);
xor U7645 (N_7645,N_7514,N_7579);
nand U7646 (N_7646,N_7535,N_7542);
xnor U7647 (N_7647,N_7502,N_7507);
and U7648 (N_7648,N_7572,N_7595);
or U7649 (N_7649,N_7580,N_7533);
xor U7650 (N_7650,N_7597,N_7578);
nand U7651 (N_7651,N_7575,N_7552);
nor U7652 (N_7652,N_7531,N_7507);
nand U7653 (N_7653,N_7572,N_7551);
xnor U7654 (N_7654,N_7587,N_7542);
nor U7655 (N_7655,N_7505,N_7538);
or U7656 (N_7656,N_7579,N_7558);
xor U7657 (N_7657,N_7505,N_7586);
nor U7658 (N_7658,N_7580,N_7515);
nor U7659 (N_7659,N_7583,N_7548);
nor U7660 (N_7660,N_7514,N_7517);
nor U7661 (N_7661,N_7502,N_7542);
nor U7662 (N_7662,N_7531,N_7562);
nor U7663 (N_7663,N_7535,N_7503);
nand U7664 (N_7664,N_7553,N_7593);
nand U7665 (N_7665,N_7578,N_7585);
or U7666 (N_7666,N_7513,N_7527);
or U7667 (N_7667,N_7582,N_7527);
nand U7668 (N_7668,N_7551,N_7570);
or U7669 (N_7669,N_7539,N_7541);
and U7670 (N_7670,N_7510,N_7514);
nor U7671 (N_7671,N_7520,N_7573);
nand U7672 (N_7672,N_7549,N_7527);
xnor U7673 (N_7673,N_7523,N_7538);
and U7674 (N_7674,N_7520,N_7511);
nor U7675 (N_7675,N_7552,N_7596);
or U7676 (N_7676,N_7548,N_7572);
and U7677 (N_7677,N_7594,N_7525);
nand U7678 (N_7678,N_7562,N_7593);
nor U7679 (N_7679,N_7591,N_7510);
nand U7680 (N_7680,N_7512,N_7585);
nor U7681 (N_7681,N_7517,N_7587);
xor U7682 (N_7682,N_7587,N_7506);
nor U7683 (N_7683,N_7546,N_7524);
and U7684 (N_7684,N_7552,N_7597);
or U7685 (N_7685,N_7545,N_7547);
nor U7686 (N_7686,N_7554,N_7557);
nand U7687 (N_7687,N_7566,N_7552);
and U7688 (N_7688,N_7527,N_7522);
nor U7689 (N_7689,N_7575,N_7564);
nor U7690 (N_7690,N_7569,N_7593);
nand U7691 (N_7691,N_7599,N_7530);
nor U7692 (N_7692,N_7545,N_7581);
nand U7693 (N_7693,N_7597,N_7537);
xor U7694 (N_7694,N_7593,N_7523);
nor U7695 (N_7695,N_7577,N_7590);
xor U7696 (N_7696,N_7573,N_7561);
and U7697 (N_7697,N_7594,N_7591);
or U7698 (N_7698,N_7508,N_7585);
nor U7699 (N_7699,N_7598,N_7508);
xnor U7700 (N_7700,N_7669,N_7666);
nor U7701 (N_7701,N_7650,N_7611);
nor U7702 (N_7702,N_7635,N_7648);
and U7703 (N_7703,N_7626,N_7677);
or U7704 (N_7704,N_7667,N_7646);
nor U7705 (N_7705,N_7682,N_7691);
or U7706 (N_7706,N_7636,N_7639);
and U7707 (N_7707,N_7622,N_7652);
or U7708 (N_7708,N_7675,N_7656);
nand U7709 (N_7709,N_7610,N_7687);
and U7710 (N_7710,N_7600,N_7695);
nand U7711 (N_7711,N_7643,N_7674);
xnor U7712 (N_7712,N_7629,N_7608);
xnor U7713 (N_7713,N_7657,N_7697);
nand U7714 (N_7714,N_7678,N_7612);
nor U7715 (N_7715,N_7661,N_7606);
nor U7716 (N_7716,N_7623,N_7655);
or U7717 (N_7717,N_7658,N_7663);
nor U7718 (N_7718,N_7653,N_7644);
nor U7719 (N_7719,N_7603,N_7640);
nor U7720 (N_7720,N_7694,N_7698);
and U7721 (N_7721,N_7638,N_7679);
nor U7722 (N_7722,N_7634,N_7625);
or U7723 (N_7723,N_7602,N_7615);
xnor U7724 (N_7724,N_7683,N_7628);
and U7725 (N_7725,N_7627,N_7685);
nand U7726 (N_7726,N_7673,N_7680);
nor U7727 (N_7727,N_7684,N_7604);
xnor U7728 (N_7728,N_7671,N_7613);
xor U7729 (N_7729,N_7654,N_7631);
and U7730 (N_7730,N_7637,N_7616);
nand U7731 (N_7731,N_7621,N_7660);
and U7732 (N_7732,N_7670,N_7693);
nor U7733 (N_7733,N_7642,N_7692);
xor U7734 (N_7734,N_7617,N_7665);
or U7735 (N_7735,N_7633,N_7614);
nand U7736 (N_7736,N_7668,N_7641);
nor U7737 (N_7737,N_7618,N_7647);
or U7738 (N_7738,N_7630,N_7609);
nor U7739 (N_7739,N_7605,N_7620);
nor U7740 (N_7740,N_7607,N_7696);
xor U7741 (N_7741,N_7681,N_7676);
xor U7742 (N_7742,N_7662,N_7689);
xor U7743 (N_7743,N_7688,N_7664);
or U7744 (N_7744,N_7632,N_7601);
nor U7745 (N_7745,N_7699,N_7690);
or U7746 (N_7746,N_7672,N_7659);
or U7747 (N_7747,N_7651,N_7686);
xor U7748 (N_7748,N_7649,N_7624);
xor U7749 (N_7749,N_7645,N_7619);
nor U7750 (N_7750,N_7632,N_7602);
and U7751 (N_7751,N_7678,N_7675);
nand U7752 (N_7752,N_7602,N_7638);
nor U7753 (N_7753,N_7639,N_7693);
xnor U7754 (N_7754,N_7678,N_7650);
or U7755 (N_7755,N_7690,N_7632);
xnor U7756 (N_7756,N_7620,N_7640);
and U7757 (N_7757,N_7645,N_7687);
xnor U7758 (N_7758,N_7672,N_7640);
and U7759 (N_7759,N_7657,N_7642);
xor U7760 (N_7760,N_7639,N_7697);
nand U7761 (N_7761,N_7600,N_7646);
or U7762 (N_7762,N_7611,N_7612);
nand U7763 (N_7763,N_7699,N_7684);
nand U7764 (N_7764,N_7620,N_7600);
nand U7765 (N_7765,N_7635,N_7671);
xnor U7766 (N_7766,N_7656,N_7660);
nor U7767 (N_7767,N_7694,N_7613);
and U7768 (N_7768,N_7653,N_7684);
and U7769 (N_7769,N_7632,N_7609);
xnor U7770 (N_7770,N_7616,N_7623);
nand U7771 (N_7771,N_7666,N_7626);
nand U7772 (N_7772,N_7632,N_7680);
or U7773 (N_7773,N_7676,N_7603);
nand U7774 (N_7774,N_7686,N_7681);
or U7775 (N_7775,N_7692,N_7651);
and U7776 (N_7776,N_7629,N_7691);
or U7777 (N_7777,N_7646,N_7678);
xnor U7778 (N_7778,N_7611,N_7681);
or U7779 (N_7779,N_7622,N_7607);
nand U7780 (N_7780,N_7693,N_7687);
nand U7781 (N_7781,N_7632,N_7646);
or U7782 (N_7782,N_7641,N_7604);
or U7783 (N_7783,N_7664,N_7619);
nand U7784 (N_7784,N_7630,N_7626);
nor U7785 (N_7785,N_7687,N_7621);
xnor U7786 (N_7786,N_7603,N_7656);
or U7787 (N_7787,N_7623,N_7683);
nor U7788 (N_7788,N_7613,N_7607);
and U7789 (N_7789,N_7603,N_7624);
and U7790 (N_7790,N_7658,N_7653);
xor U7791 (N_7791,N_7623,N_7610);
or U7792 (N_7792,N_7643,N_7696);
nand U7793 (N_7793,N_7662,N_7622);
nand U7794 (N_7794,N_7602,N_7624);
nand U7795 (N_7795,N_7643,N_7695);
nor U7796 (N_7796,N_7604,N_7674);
nand U7797 (N_7797,N_7623,N_7635);
and U7798 (N_7798,N_7679,N_7646);
nand U7799 (N_7799,N_7604,N_7603);
xor U7800 (N_7800,N_7764,N_7717);
and U7801 (N_7801,N_7707,N_7705);
nand U7802 (N_7802,N_7748,N_7773);
nand U7803 (N_7803,N_7713,N_7703);
xnor U7804 (N_7804,N_7777,N_7706);
nor U7805 (N_7805,N_7729,N_7718);
nor U7806 (N_7806,N_7712,N_7702);
or U7807 (N_7807,N_7765,N_7725);
nand U7808 (N_7808,N_7797,N_7700);
and U7809 (N_7809,N_7791,N_7723);
nand U7810 (N_7810,N_7770,N_7739);
nand U7811 (N_7811,N_7751,N_7731);
xnor U7812 (N_7812,N_7732,N_7761);
or U7813 (N_7813,N_7752,N_7743);
or U7814 (N_7814,N_7708,N_7744);
nand U7815 (N_7815,N_7728,N_7720);
or U7816 (N_7816,N_7749,N_7716);
or U7817 (N_7817,N_7710,N_7715);
and U7818 (N_7818,N_7741,N_7726);
nand U7819 (N_7819,N_7709,N_7795);
nor U7820 (N_7820,N_7745,N_7794);
and U7821 (N_7821,N_7776,N_7783);
nor U7822 (N_7822,N_7780,N_7734);
and U7823 (N_7823,N_7767,N_7787);
and U7824 (N_7824,N_7754,N_7721);
xor U7825 (N_7825,N_7793,N_7742);
or U7826 (N_7826,N_7769,N_7727);
nor U7827 (N_7827,N_7768,N_7730);
and U7828 (N_7828,N_7762,N_7740);
or U7829 (N_7829,N_7750,N_7753);
nand U7830 (N_7830,N_7798,N_7774);
or U7831 (N_7831,N_7771,N_7738);
or U7832 (N_7832,N_7737,N_7756);
or U7833 (N_7833,N_7724,N_7746);
or U7834 (N_7834,N_7766,N_7772);
or U7835 (N_7835,N_7735,N_7704);
nor U7836 (N_7836,N_7719,N_7790);
nor U7837 (N_7837,N_7714,N_7781);
and U7838 (N_7838,N_7784,N_7711);
xor U7839 (N_7839,N_7757,N_7788);
xnor U7840 (N_7840,N_7759,N_7747);
and U7841 (N_7841,N_7792,N_7701);
nand U7842 (N_7842,N_7785,N_7760);
xor U7843 (N_7843,N_7736,N_7778);
nand U7844 (N_7844,N_7775,N_7722);
or U7845 (N_7845,N_7789,N_7758);
xor U7846 (N_7846,N_7733,N_7782);
or U7847 (N_7847,N_7796,N_7799);
nand U7848 (N_7848,N_7786,N_7755);
nand U7849 (N_7849,N_7779,N_7763);
nor U7850 (N_7850,N_7750,N_7762);
or U7851 (N_7851,N_7777,N_7731);
nand U7852 (N_7852,N_7782,N_7764);
and U7853 (N_7853,N_7765,N_7738);
xnor U7854 (N_7854,N_7747,N_7722);
and U7855 (N_7855,N_7722,N_7761);
nand U7856 (N_7856,N_7780,N_7709);
nor U7857 (N_7857,N_7789,N_7727);
or U7858 (N_7858,N_7794,N_7722);
nor U7859 (N_7859,N_7770,N_7768);
nor U7860 (N_7860,N_7755,N_7757);
and U7861 (N_7861,N_7734,N_7793);
nor U7862 (N_7862,N_7760,N_7758);
xnor U7863 (N_7863,N_7714,N_7710);
and U7864 (N_7864,N_7759,N_7723);
nor U7865 (N_7865,N_7772,N_7765);
or U7866 (N_7866,N_7723,N_7763);
and U7867 (N_7867,N_7770,N_7776);
nor U7868 (N_7868,N_7743,N_7742);
and U7869 (N_7869,N_7780,N_7738);
nor U7870 (N_7870,N_7746,N_7710);
nor U7871 (N_7871,N_7795,N_7738);
or U7872 (N_7872,N_7767,N_7712);
xnor U7873 (N_7873,N_7740,N_7766);
or U7874 (N_7874,N_7743,N_7794);
xnor U7875 (N_7875,N_7727,N_7706);
and U7876 (N_7876,N_7739,N_7763);
xnor U7877 (N_7877,N_7716,N_7748);
nor U7878 (N_7878,N_7723,N_7748);
and U7879 (N_7879,N_7707,N_7766);
nor U7880 (N_7880,N_7717,N_7719);
xnor U7881 (N_7881,N_7772,N_7713);
or U7882 (N_7882,N_7787,N_7757);
nand U7883 (N_7883,N_7785,N_7754);
xnor U7884 (N_7884,N_7790,N_7773);
nor U7885 (N_7885,N_7707,N_7715);
and U7886 (N_7886,N_7715,N_7756);
nand U7887 (N_7887,N_7765,N_7784);
nor U7888 (N_7888,N_7778,N_7704);
or U7889 (N_7889,N_7799,N_7724);
or U7890 (N_7890,N_7743,N_7736);
xnor U7891 (N_7891,N_7706,N_7733);
nand U7892 (N_7892,N_7758,N_7743);
nand U7893 (N_7893,N_7722,N_7718);
nor U7894 (N_7894,N_7790,N_7734);
xor U7895 (N_7895,N_7766,N_7749);
and U7896 (N_7896,N_7755,N_7744);
nand U7897 (N_7897,N_7709,N_7726);
nor U7898 (N_7898,N_7737,N_7762);
nand U7899 (N_7899,N_7773,N_7774);
xnor U7900 (N_7900,N_7838,N_7862);
or U7901 (N_7901,N_7841,N_7804);
and U7902 (N_7902,N_7861,N_7871);
xnor U7903 (N_7903,N_7873,N_7868);
xor U7904 (N_7904,N_7856,N_7848);
xnor U7905 (N_7905,N_7809,N_7822);
and U7906 (N_7906,N_7814,N_7888);
nor U7907 (N_7907,N_7876,N_7870);
or U7908 (N_7908,N_7824,N_7859);
or U7909 (N_7909,N_7815,N_7816);
nor U7910 (N_7910,N_7890,N_7892);
nor U7911 (N_7911,N_7878,N_7872);
nor U7912 (N_7912,N_7821,N_7826);
nand U7913 (N_7913,N_7857,N_7885);
nand U7914 (N_7914,N_7800,N_7865);
nand U7915 (N_7915,N_7864,N_7886);
or U7916 (N_7916,N_7858,N_7811);
nor U7917 (N_7917,N_7837,N_7884);
nor U7918 (N_7918,N_7833,N_7839);
and U7919 (N_7919,N_7808,N_7801);
or U7920 (N_7920,N_7832,N_7883);
or U7921 (N_7921,N_7812,N_7897);
or U7922 (N_7922,N_7898,N_7863);
nor U7923 (N_7923,N_7855,N_7891);
nor U7924 (N_7924,N_7810,N_7813);
or U7925 (N_7925,N_7807,N_7803);
nand U7926 (N_7926,N_7843,N_7893);
nand U7927 (N_7927,N_7825,N_7823);
nor U7928 (N_7928,N_7887,N_7818);
and U7929 (N_7929,N_7852,N_7875);
xor U7930 (N_7930,N_7831,N_7879);
nand U7931 (N_7931,N_7819,N_7827);
nor U7932 (N_7932,N_7844,N_7853);
or U7933 (N_7933,N_7845,N_7851);
and U7934 (N_7934,N_7836,N_7849);
xor U7935 (N_7935,N_7805,N_7881);
nand U7936 (N_7936,N_7806,N_7829);
or U7937 (N_7937,N_7817,N_7850);
nand U7938 (N_7938,N_7866,N_7874);
or U7939 (N_7939,N_7882,N_7830);
xnor U7940 (N_7940,N_7847,N_7899);
or U7941 (N_7941,N_7869,N_7842);
nand U7942 (N_7942,N_7835,N_7834);
xor U7943 (N_7943,N_7820,N_7802);
or U7944 (N_7944,N_7889,N_7877);
and U7945 (N_7945,N_7860,N_7880);
nand U7946 (N_7946,N_7867,N_7896);
nor U7947 (N_7947,N_7895,N_7828);
xnor U7948 (N_7948,N_7846,N_7894);
nor U7949 (N_7949,N_7840,N_7854);
and U7950 (N_7950,N_7875,N_7843);
or U7951 (N_7951,N_7811,N_7887);
or U7952 (N_7952,N_7883,N_7805);
nor U7953 (N_7953,N_7844,N_7893);
and U7954 (N_7954,N_7884,N_7822);
nor U7955 (N_7955,N_7855,N_7877);
nor U7956 (N_7956,N_7817,N_7879);
or U7957 (N_7957,N_7890,N_7820);
nor U7958 (N_7958,N_7801,N_7876);
and U7959 (N_7959,N_7864,N_7896);
xor U7960 (N_7960,N_7828,N_7859);
and U7961 (N_7961,N_7839,N_7858);
xor U7962 (N_7962,N_7840,N_7882);
nand U7963 (N_7963,N_7820,N_7868);
xor U7964 (N_7964,N_7877,N_7811);
or U7965 (N_7965,N_7883,N_7874);
and U7966 (N_7966,N_7854,N_7869);
or U7967 (N_7967,N_7851,N_7848);
and U7968 (N_7968,N_7810,N_7800);
and U7969 (N_7969,N_7861,N_7859);
and U7970 (N_7970,N_7872,N_7804);
nand U7971 (N_7971,N_7819,N_7848);
nor U7972 (N_7972,N_7819,N_7883);
nand U7973 (N_7973,N_7809,N_7868);
xor U7974 (N_7974,N_7857,N_7845);
or U7975 (N_7975,N_7866,N_7871);
nor U7976 (N_7976,N_7839,N_7830);
xnor U7977 (N_7977,N_7863,N_7852);
nand U7978 (N_7978,N_7830,N_7885);
nor U7979 (N_7979,N_7876,N_7804);
or U7980 (N_7980,N_7853,N_7894);
xnor U7981 (N_7981,N_7881,N_7815);
nand U7982 (N_7982,N_7807,N_7818);
and U7983 (N_7983,N_7824,N_7806);
nand U7984 (N_7984,N_7885,N_7849);
nand U7985 (N_7985,N_7883,N_7856);
nand U7986 (N_7986,N_7801,N_7822);
or U7987 (N_7987,N_7863,N_7832);
and U7988 (N_7988,N_7816,N_7824);
and U7989 (N_7989,N_7873,N_7834);
and U7990 (N_7990,N_7850,N_7801);
xor U7991 (N_7991,N_7893,N_7804);
nor U7992 (N_7992,N_7868,N_7850);
xor U7993 (N_7993,N_7879,N_7888);
xor U7994 (N_7994,N_7856,N_7892);
nor U7995 (N_7995,N_7883,N_7871);
and U7996 (N_7996,N_7851,N_7817);
or U7997 (N_7997,N_7842,N_7881);
nand U7998 (N_7998,N_7899,N_7835);
and U7999 (N_7999,N_7899,N_7855);
nand U8000 (N_8000,N_7950,N_7949);
nand U8001 (N_8001,N_7972,N_7981);
and U8002 (N_8002,N_7982,N_7961);
and U8003 (N_8003,N_7921,N_7912);
nand U8004 (N_8004,N_7976,N_7969);
xnor U8005 (N_8005,N_7959,N_7908);
and U8006 (N_8006,N_7989,N_7971);
nand U8007 (N_8007,N_7902,N_7918);
and U8008 (N_8008,N_7963,N_7916);
nor U8009 (N_8009,N_7964,N_7948);
nand U8010 (N_8010,N_7910,N_7978);
nand U8011 (N_8011,N_7945,N_7924);
nor U8012 (N_8012,N_7998,N_7986);
xnor U8013 (N_8013,N_7925,N_7951);
nand U8014 (N_8014,N_7974,N_7952);
nand U8015 (N_8015,N_7984,N_7953);
nor U8016 (N_8016,N_7929,N_7970);
nor U8017 (N_8017,N_7928,N_7943);
nor U8018 (N_8018,N_7991,N_7988);
and U8019 (N_8019,N_7913,N_7994);
nor U8020 (N_8020,N_7983,N_7939);
nor U8021 (N_8021,N_7936,N_7940);
xnor U8022 (N_8022,N_7979,N_7968);
xor U8023 (N_8023,N_7934,N_7966);
and U8024 (N_8024,N_7957,N_7997);
or U8025 (N_8025,N_7958,N_7941);
or U8026 (N_8026,N_7917,N_7922);
or U8027 (N_8027,N_7973,N_7926);
nand U8028 (N_8028,N_7975,N_7992);
and U8029 (N_8029,N_7919,N_7956);
xor U8030 (N_8030,N_7901,N_7938);
and U8031 (N_8031,N_7937,N_7980);
or U8032 (N_8032,N_7960,N_7947);
nand U8033 (N_8033,N_7909,N_7932);
nand U8034 (N_8034,N_7906,N_7933);
xor U8035 (N_8035,N_7967,N_7903);
nand U8036 (N_8036,N_7930,N_7944);
or U8037 (N_8037,N_7905,N_7977);
and U8038 (N_8038,N_7962,N_7914);
nand U8039 (N_8039,N_7955,N_7999);
and U8040 (N_8040,N_7942,N_7911);
and U8041 (N_8041,N_7965,N_7993);
nor U8042 (N_8042,N_7990,N_7900);
or U8043 (N_8043,N_7923,N_7904);
and U8044 (N_8044,N_7985,N_7931);
nand U8045 (N_8045,N_7987,N_7946);
or U8046 (N_8046,N_7954,N_7907);
nor U8047 (N_8047,N_7915,N_7995);
xnor U8048 (N_8048,N_7996,N_7920);
nor U8049 (N_8049,N_7935,N_7927);
and U8050 (N_8050,N_7967,N_7999);
nor U8051 (N_8051,N_7943,N_7965);
nor U8052 (N_8052,N_7996,N_7955);
nor U8053 (N_8053,N_7996,N_7999);
nand U8054 (N_8054,N_7930,N_7977);
or U8055 (N_8055,N_7950,N_7948);
and U8056 (N_8056,N_7947,N_7988);
xnor U8057 (N_8057,N_7910,N_7986);
xor U8058 (N_8058,N_7989,N_7968);
or U8059 (N_8059,N_7948,N_7953);
or U8060 (N_8060,N_7921,N_7998);
xnor U8061 (N_8061,N_7931,N_7923);
nand U8062 (N_8062,N_7913,N_7927);
and U8063 (N_8063,N_7974,N_7992);
or U8064 (N_8064,N_7938,N_7913);
nor U8065 (N_8065,N_7916,N_7932);
nand U8066 (N_8066,N_7935,N_7943);
and U8067 (N_8067,N_7941,N_7930);
nor U8068 (N_8068,N_7919,N_7992);
and U8069 (N_8069,N_7971,N_7951);
or U8070 (N_8070,N_7974,N_7993);
xnor U8071 (N_8071,N_7951,N_7992);
nor U8072 (N_8072,N_7956,N_7960);
and U8073 (N_8073,N_7940,N_7969);
xnor U8074 (N_8074,N_7947,N_7974);
or U8075 (N_8075,N_7957,N_7919);
and U8076 (N_8076,N_7906,N_7902);
or U8077 (N_8077,N_7932,N_7969);
or U8078 (N_8078,N_7969,N_7960);
or U8079 (N_8079,N_7906,N_7970);
or U8080 (N_8080,N_7994,N_7985);
nor U8081 (N_8081,N_7935,N_7925);
nand U8082 (N_8082,N_7915,N_7945);
or U8083 (N_8083,N_7980,N_7971);
xnor U8084 (N_8084,N_7923,N_7999);
and U8085 (N_8085,N_7902,N_7955);
or U8086 (N_8086,N_7977,N_7999);
nand U8087 (N_8087,N_7922,N_7968);
and U8088 (N_8088,N_7960,N_7946);
nor U8089 (N_8089,N_7994,N_7991);
and U8090 (N_8090,N_7957,N_7950);
nor U8091 (N_8091,N_7966,N_7958);
nand U8092 (N_8092,N_7950,N_7965);
and U8093 (N_8093,N_7919,N_7974);
and U8094 (N_8094,N_7906,N_7909);
and U8095 (N_8095,N_7903,N_7975);
and U8096 (N_8096,N_7976,N_7955);
or U8097 (N_8097,N_7903,N_7959);
and U8098 (N_8098,N_7990,N_7961);
nand U8099 (N_8099,N_7934,N_7960);
xor U8100 (N_8100,N_8022,N_8082);
nand U8101 (N_8101,N_8032,N_8076);
xor U8102 (N_8102,N_8015,N_8000);
xor U8103 (N_8103,N_8096,N_8047);
or U8104 (N_8104,N_8091,N_8062);
xor U8105 (N_8105,N_8030,N_8013);
or U8106 (N_8106,N_8090,N_8009);
or U8107 (N_8107,N_8018,N_8017);
and U8108 (N_8108,N_8002,N_8039);
xnor U8109 (N_8109,N_8095,N_8099);
and U8110 (N_8110,N_8086,N_8004);
or U8111 (N_8111,N_8024,N_8041);
and U8112 (N_8112,N_8025,N_8038);
xor U8113 (N_8113,N_8027,N_8011);
xor U8114 (N_8114,N_8097,N_8057);
xor U8115 (N_8115,N_8059,N_8003);
and U8116 (N_8116,N_8026,N_8056);
and U8117 (N_8117,N_8020,N_8021);
nor U8118 (N_8118,N_8065,N_8034);
and U8119 (N_8119,N_8014,N_8079);
nor U8120 (N_8120,N_8052,N_8092);
xnor U8121 (N_8121,N_8046,N_8078);
nor U8122 (N_8122,N_8074,N_8054);
or U8123 (N_8123,N_8043,N_8042);
or U8124 (N_8124,N_8067,N_8066);
nand U8125 (N_8125,N_8016,N_8036);
nor U8126 (N_8126,N_8005,N_8058);
or U8127 (N_8127,N_8028,N_8094);
or U8128 (N_8128,N_8080,N_8055);
and U8129 (N_8129,N_8083,N_8069);
xnor U8130 (N_8130,N_8051,N_8098);
or U8131 (N_8131,N_8072,N_8048);
or U8132 (N_8132,N_8019,N_8070);
and U8133 (N_8133,N_8064,N_8089);
xnor U8134 (N_8134,N_8037,N_8081);
nor U8135 (N_8135,N_8075,N_8063);
nand U8136 (N_8136,N_8077,N_8001);
or U8137 (N_8137,N_8031,N_8087);
nand U8138 (N_8138,N_8010,N_8007);
nor U8139 (N_8139,N_8088,N_8093);
and U8140 (N_8140,N_8035,N_8033);
or U8141 (N_8141,N_8071,N_8053);
xor U8142 (N_8142,N_8049,N_8045);
nor U8143 (N_8143,N_8073,N_8006);
nand U8144 (N_8144,N_8068,N_8050);
xor U8145 (N_8145,N_8085,N_8012);
nor U8146 (N_8146,N_8029,N_8023);
nand U8147 (N_8147,N_8084,N_8008);
and U8148 (N_8148,N_8060,N_8040);
or U8149 (N_8149,N_8044,N_8061);
and U8150 (N_8150,N_8017,N_8046);
or U8151 (N_8151,N_8020,N_8061);
and U8152 (N_8152,N_8085,N_8069);
nor U8153 (N_8153,N_8006,N_8077);
or U8154 (N_8154,N_8019,N_8074);
nor U8155 (N_8155,N_8097,N_8053);
or U8156 (N_8156,N_8015,N_8067);
nand U8157 (N_8157,N_8026,N_8096);
and U8158 (N_8158,N_8076,N_8007);
xor U8159 (N_8159,N_8037,N_8083);
or U8160 (N_8160,N_8014,N_8058);
or U8161 (N_8161,N_8006,N_8002);
xor U8162 (N_8162,N_8003,N_8011);
or U8163 (N_8163,N_8022,N_8010);
and U8164 (N_8164,N_8048,N_8000);
xor U8165 (N_8165,N_8076,N_8094);
or U8166 (N_8166,N_8023,N_8034);
nor U8167 (N_8167,N_8024,N_8048);
nor U8168 (N_8168,N_8009,N_8052);
nand U8169 (N_8169,N_8057,N_8061);
xor U8170 (N_8170,N_8040,N_8019);
xor U8171 (N_8171,N_8022,N_8074);
nor U8172 (N_8172,N_8005,N_8046);
or U8173 (N_8173,N_8003,N_8027);
and U8174 (N_8174,N_8055,N_8083);
and U8175 (N_8175,N_8011,N_8062);
and U8176 (N_8176,N_8041,N_8067);
nor U8177 (N_8177,N_8030,N_8000);
nand U8178 (N_8178,N_8023,N_8015);
xnor U8179 (N_8179,N_8079,N_8011);
and U8180 (N_8180,N_8034,N_8039);
and U8181 (N_8181,N_8098,N_8060);
nand U8182 (N_8182,N_8062,N_8069);
nor U8183 (N_8183,N_8042,N_8069);
and U8184 (N_8184,N_8072,N_8037);
nor U8185 (N_8185,N_8040,N_8057);
xor U8186 (N_8186,N_8022,N_8057);
nand U8187 (N_8187,N_8080,N_8033);
nand U8188 (N_8188,N_8085,N_8017);
nor U8189 (N_8189,N_8073,N_8059);
or U8190 (N_8190,N_8098,N_8018);
nor U8191 (N_8191,N_8013,N_8021);
and U8192 (N_8192,N_8039,N_8038);
nand U8193 (N_8193,N_8046,N_8007);
nand U8194 (N_8194,N_8089,N_8007);
nand U8195 (N_8195,N_8064,N_8010);
and U8196 (N_8196,N_8045,N_8032);
or U8197 (N_8197,N_8074,N_8041);
or U8198 (N_8198,N_8028,N_8041);
and U8199 (N_8199,N_8049,N_8086);
nor U8200 (N_8200,N_8184,N_8183);
xor U8201 (N_8201,N_8143,N_8159);
xnor U8202 (N_8202,N_8155,N_8195);
or U8203 (N_8203,N_8113,N_8165);
and U8204 (N_8204,N_8118,N_8147);
nand U8205 (N_8205,N_8131,N_8198);
or U8206 (N_8206,N_8173,N_8175);
nand U8207 (N_8207,N_8116,N_8144);
or U8208 (N_8208,N_8127,N_8190);
and U8209 (N_8209,N_8167,N_8174);
nor U8210 (N_8210,N_8139,N_8109);
nand U8211 (N_8211,N_8141,N_8142);
nand U8212 (N_8212,N_8106,N_8120);
nand U8213 (N_8213,N_8150,N_8104);
nand U8214 (N_8214,N_8172,N_8191);
xnor U8215 (N_8215,N_8140,N_8138);
and U8216 (N_8216,N_8164,N_8178);
nor U8217 (N_8217,N_8179,N_8161);
nor U8218 (N_8218,N_8130,N_8137);
or U8219 (N_8219,N_8133,N_8124);
xnor U8220 (N_8220,N_8129,N_8192);
or U8221 (N_8221,N_8169,N_8122);
and U8222 (N_8222,N_8193,N_8170);
and U8223 (N_8223,N_8171,N_8105);
nor U8224 (N_8224,N_8189,N_8185);
and U8225 (N_8225,N_8153,N_8110);
nand U8226 (N_8226,N_8114,N_8160);
xnor U8227 (N_8227,N_8119,N_8107);
nand U8228 (N_8228,N_8135,N_8100);
xnor U8229 (N_8229,N_8126,N_8115);
xnor U8230 (N_8230,N_8136,N_8134);
xor U8231 (N_8231,N_8180,N_8168);
or U8232 (N_8232,N_8187,N_8157);
xnor U8233 (N_8233,N_8125,N_8182);
or U8234 (N_8234,N_8112,N_8149);
nor U8235 (N_8235,N_8108,N_8162);
xnor U8236 (N_8236,N_8145,N_8123);
nand U8237 (N_8237,N_8146,N_8152);
nand U8238 (N_8238,N_8194,N_8111);
and U8239 (N_8239,N_8163,N_8132);
xor U8240 (N_8240,N_8102,N_8196);
and U8241 (N_8241,N_8121,N_8181);
nand U8242 (N_8242,N_8176,N_8186);
xnor U8243 (N_8243,N_8199,N_8188);
nor U8244 (N_8244,N_8156,N_8154);
nand U8245 (N_8245,N_8151,N_8166);
nand U8246 (N_8246,N_8197,N_8101);
and U8247 (N_8247,N_8128,N_8117);
and U8248 (N_8248,N_8177,N_8148);
and U8249 (N_8249,N_8158,N_8103);
nand U8250 (N_8250,N_8167,N_8138);
or U8251 (N_8251,N_8109,N_8162);
nor U8252 (N_8252,N_8186,N_8175);
xor U8253 (N_8253,N_8105,N_8115);
nand U8254 (N_8254,N_8188,N_8133);
xor U8255 (N_8255,N_8180,N_8171);
or U8256 (N_8256,N_8100,N_8114);
and U8257 (N_8257,N_8175,N_8142);
or U8258 (N_8258,N_8182,N_8193);
or U8259 (N_8259,N_8158,N_8161);
and U8260 (N_8260,N_8177,N_8110);
or U8261 (N_8261,N_8144,N_8163);
nand U8262 (N_8262,N_8138,N_8166);
nand U8263 (N_8263,N_8192,N_8190);
nor U8264 (N_8264,N_8183,N_8104);
nor U8265 (N_8265,N_8160,N_8106);
nor U8266 (N_8266,N_8195,N_8150);
and U8267 (N_8267,N_8193,N_8104);
xor U8268 (N_8268,N_8178,N_8157);
nor U8269 (N_8269,N_8196,N_8194);
nor U8270 (N_8270,N_8161,N_8188);
xnor U8271 (N_8271,N_8148,N_8153);
or U8272 (N_8272,N_8143,N_8140);
xor U8273 (N_8273,N_8150,N_8165);
or U8274 (N_8274,N_8198,N_8125);
or U8275 (N_8275,N_8131,N_8105);
nand U8276 (N_8276,N_8129,N_8189);
and U8277 (N_8277,N_8129,N_8149);
and U8278 (N_8278,N_8156,N_8114);
xor U8279 (N_8279,N_8115,N_8162);
xnor U8280 (N_8280,N_8114,N_8158);
or U8281 (N_8281,N_8149,N_8120);
nor U8282 (N_8282,N_8196,N_8120);
xor U8283 (N_8283,N_8173,N_8116);
nand U8284 (N_8284,N_8119,N_8199);
nand U8285 (N_8285,N_8195,N_8136);
or U8286 (N_8286,N_8187,N_8124);
or U8287 (N_8287,N_8196,N_8158);
and U8288 (N_8288,N_8174,N_8187);
nor U8289 (N_8289,N_8110,N_8135);
or U8290 (N_8290,N_8106,N_8113);
and U8291 (N_8291,N_8173,N_8192);
nor U8292 (N_8292,N_8150,N_8109);
nand U8293 (N_8293,N_8154,N_8108);
nor U8294 (N_8294,N_8110,N_8178);
or U8295 (N_8295,N_8129,N_8145);
nand U8296 (N_8296,N_8125,N_8110);
nor U8297 (N_8297,N_8181,N_8190);
nor U8298 (N_8298,N_8155,N_8144);
xnor U8299 (N_8299,N_8143,N_8171);
nor U8300 (N_8300,N_8258,N_8210);
or U8301 (N_8301,N_8215,N_8266);
nor U8302 (N_8302,N_8270,N_8232);
or U8303 (N_8303,N_8254,N_8255);
and U8304 (N_8304,N_8236,N_8245);
nand U8305 (N_8305,N_8260,N_8208);
nand U8306 (N_8306,N_8278,N_8277);
xor U8307 (N_8307,N_8204,N_8225);
or U8308 (N_8308,N_8276,N_8252);
nand U8309 (N_8309,N_8257,N_8226);
nor U8310 (N_8310,N_8296,N_8200);
nor U8311 (N_8311,N_8205,N_8286);
and U8312 (N_8312,N_8207,N_8287);
nand U8313 (N_8313,N_8263,N_8271);
or U8314 (N_8314,N_8242,N_8291);
or U8315 (N_8315,N_8220,N_8221);
and U8316 (N_8316,N_8217,N_8202);
nor U8317 (N_8317,N_8280,N_8283);
and U8318 (N_8318,N_8227,N_8253);
nor U8319 (N_8319,N_8269,N_8275);
or U8320 (N_8320,N_8211,N_8292);
nor U8321 (N_8321,N_8234,N_8214);
or U8322 (N_8322,N_8241,N_8203);
or U8323 (N_8323,N_8251,N_8218);
xnor U8324 (N_8324,N_8239,N_8209);
and U8325 (N_8325,N_8299,N_8238);
xnor U8326 (N_8326,N_8279,N_8224);
nor U8327 (N_8327,N_8228,N_8240);
nor U8328 (N_8328,N_8259,N_8256);
nand U8329 (N_8329,N_8294,N_8284);
or U8330 (N_8330,N_8216,N_8248);
nand U8331 (N_8331,N_8272,N_8281);
xor U8332 (N_8332,N_8206,N_8244);
or U8333 (N_8333,N_8290,N_8268);
xor U8334 (N_8334,N_8298,N_8273);
xnor U8335 (N_8335,N_8274,N_8243);
or U8336 (N_8336,N_8262,N_8246);
or U8337 (N_8337,N_8293,N_8285);
and U8338 (N_8338,N_8213,N_8230);
or U8339 (N_8339,N_8235,N_8282);
nand U8340 (N_8340,N_8288,N_8212);
and U8341 (N_8341,N_8267,N_8222);
or U8342 (N_8342,N_8295,N_8261);
and U8343 (N_8343,N_8297,N_8237);
nand U8344 (N_8344,N_8289,N_8223);
nor U8345 (N_8345,N_8201,N_8233);
and U8346 (N_8346,N_8219,N_8247);
nor U8347 (N_8347,N_8264,N_8229);
or U8348 (N_8348,N_8265,N_8231);
nor U8349 (N_8349,N_8249,N_8250);
or U8350 (N_8350,N_8288,N_8254);
nand U8351 (N_8351,N_8276,N_8266);
nor U8352 (N_8352,N_8209,N_8282);
or U8353 (N_8353,N_8276,N_8299);
and U8354 (N_8354,N_8264,N_8254);
xor U8355 (N_8355,N_8220,N_8260);
nand U8356 (N_8356,N_8259,N_8249);
or U8357 (N_8357,N_8292,N_8222);
or U8358 (N_8358,N_8271,N_8216);
xor U8359 (N_8359,N_8244,N_8283);
nand U8360 (N_8360,N_8245,N_8289);
nand U8361 (N_8361,N_8296,N_8277);
nor U8362 (N_8362,N_8291,N_8254);
and U8363 (N_8363,N_8215,N_8271);
or U8364 (N_8364,N_8274,N_8267);
xnor U8365 (N_8365,N_8243,N_8226);
and U8366 (N_8366,N_8232,N_8277);
nor U8367 (N_8367,N_8234,N_8201);
nand U8368 (N_8368,N_8277,N_8247);
or U8369 (N_8369,N_8264,N_8216);
nor U8370 (N_8370,N_8226,N_8278);
xnor U8371 (N_8371,N_8256,N_8223);
or U8372 (N_8372,N_8269,N_8210);
and U8373 (N_8373,N_8242,N_8283);
nand U8374 (N_8374,N_8283,N_8252);
nand U8375 (N_8375,N_8267,N_8290);
nor U8376 (N_8376,N_8205,N_8254);
nor U8377 (N_8377,N_8209,N_8295);
nor U8378 (N_8378,N_8231,N_8251);
or U8379 (N_8379,N_8265,N_8252);
nor U8380 (N_8380,N_8255,N_8219);
or U8381 (N_8381,N_8224,N_8285);
nor U8382 (N_8382,N_8286,N_8269);
and U8383 (N_8383,N_8209,N_8279);
xor U8384 (N_8384,N_8234,N_8287);
xnor U8385 (N_8385,N_8205,N_8202);
and U8386 (N_8386,N_8212,N_8231);
and U8387 (N_8387,N_8265,N_8214);
xor U8388 (N_8388,N_8257,N_8290);
nand U8389 (N_8389,N_8295,N_8203);
and U8390 (N_8390,N_8262,N_8240);
or U8391 (N_8391,N_8223,N_8216);
nand U8392 (N_8392,N_8232,N_8287);
and U8393 (N_8393,N_8232,N_8281);
and U8394 (N_8394,N_8245,N_8233);
or U8395 (N_8395,N_8229,N_8206);
nor U8396 (N_8396,N_8232,N_8203);
nand U8397 (N_8397,N_8281,N_8226);
xnor U8398 (N_8398,N_8242,N_8223);
and U8399 (N_8399,N_8228,N_8269);
nor U8400 (N_8400,N_8378,N_8324);
nor U8401 (N_8401,N_8396,N_8364);
nor U8402 (N_8402,N_8370,N_8387);
and U8403 (N_8403,N_8313,N_8347);
and U8404 (N_8404,N_8379,N_8343);
nand U8405 (N_8405,N_8377,N_8349);
xnor U8406 (N_8406,N_8382,N_8311);
and U8407 (N_8407,N_8328,N_8395);
or U8408 (N_8408,N_8389,N_8331);
xor U8409 (N_8409,N_8304,N_8373);
or U8410 (N_8410,N_8302,N_8333);
nor U8411 (N_8411,N_8307,N_8335);
or U8412 (N_8412,N_8393,N_8325);
or U8413 (N_8413,N_8319,N_8309);
nor U8414 (N_8414,N_8330,N_8355);
nor U8415 (N_8415,N_8323,N_8342);
or U8416 (N_8416,N_8344,N_8352);
xor U8417 (N_8417,N_8332,N_8300);
nand U8418 (N_8418,N_8341,N_8354);
xnor U8419 (N_8419,N_8346,N_8318);
or U8420 (N_8420,N_8350,N_8391);
xor U8421 (N_8421,N_8336,N_8356);
xor U8422 (N_8422,N_8338,N_8372);
and U8423 (N_8423,N_8326,N_8366);
or U8424 (N_8424,N_8315,N_8316);
nor U8425 (N_8425,N_8303,N_8380);
nand U8426 (N_8426,N_8374,N_8322);
xor U8427 (N_8427,N_8399,N_8312);
xnor U8428 (N_8428,N_8385,N_8345);
and U8429 (N_8429,N_8376,N_8388);
xnor U8430 (N_8430,N_8305,N_8321);
or U8431 (N_8431,N_8353,N_8348);
and U8432 (N_8432,N_8363,N_8365);
or U8433 (N_8433,N_8317,N_8397);
and U8434 (N_8434,N_8381,N_8308);
or U8435 (N_8435,N_8367,N_8357);
nand U8436 (N_8436,N_8383,N_8384);
xnor U8437 (N_8437,N_8329,N_8301);
nor U8438 (N_8438,N_8310,N_8334);
xor U8439 (N_8439,N_8327,N_8340);
nand U8440 (N_8440,N_8390,N_8320);
nor U8441 (N_8441,N_8398,N_8351);
and U8442 (N_8442,N_8394,N_8337);
nand U8443 (N_8443,N_8306,N_8339);
xor U8444 (N_8444,N_8360,N_8358);
xor U8445 (N_8445,N_8371,N_8368);
and U8446 (N_8446,N_8392,N_8386);
and U8447 (N_8447,N_8369,N_8362);
or U8448 (N_8448,N_8375,N_8361);
and U8449 (N_8449,N_8314,N_8359);
nand U8450 (N_8450,N_8323,N_8349);
nor U8451 (N_8451,N_8344,N_8311);
xnor U8452 (N_8452,N_8328,N_8303);
or U8453 (N_8453,N_8357,N_8382);
and U8454 (N_8454,N_8384,N_8319);
and U8455 (N_8455,N_8329,N_8396);
xnor U8456 (N_8456,N_8383,N_8361);
xor U8457 (N_8457,N_8305,N_8324);
nor U8458 (N_8458,N_8362,N_8352);
nand U8459 (N_8459,N_8330,N_8306);
and U8460 (N_8460,N_8361,N_8369);
and U8461 (N_8461,N_8374,N_8362);
nand U8462 (N_8462,N_8315,N_8379);
and U8463 (N_8463,N_8329,N_8395);
or U8464 (N_8464,N_8320,N_8363);
and U8465 (N_8465,N_8312,N_8311);
or U8466 (N_8466,N_8306,N_8392);
xor U8467 (N_8467,N_8370,N_8396);
nor U8468 (N_8468,N_8369,N_8357);
xor U8469 (N_8469,N_8362,N_8377);
nand U8470 (N_8470,N_8399,N_8369);
xnor U8471 (N_8471,N_8339,N_8399);
or U8472 (N_8472,N_8394,N_8348);
and U8473 (N_8473,N_8320,N_8306);
and U8474 (N_8474,N_8357,N_8388);
nor U8475 (N_8475,N_8354,N_8386);
nand U8476 (N_8476,N_8336,N_8379);
nand U8477 (N_8477,N_8395,N_8305);
or U8478 (N_8478,N_8309,N_8373);
or U8479 (N_8479,N_8302,N_8320);
xnor U8480 (N_8480,N_8306,N_8384);
or U8481 (N_8481,N_8370,N_8382);
xnor U8482 (N_8482,N_8375,N_8319);
and U8483 (N_8483,N_8301,N_8309);
xor U8484 (N_8484,N_8326,N_8353);
nor U8485 (N_8485,N_8309,N_8348);
nor U8486 (N_8486,N_8332,N_8356);
nand U8487 (N_8487,N_8366,N_8397);
or U8488 (N_8488,N_8320,N_8367);
and U8489 (N_8489,N_8370,N_8373);
and U8490 (N_8490,N_8324,N_8307);
xor U8491 (N_8491,N_8392,N_8335);
xor U8492 (N_8492,N_8301,N_8320);
or U8493 (N_8493,N_8372,N_8306);
or U8494 (N_8494,N_8379,N_8309);
nor U8495 (N_8495,N_8372,N_8359);
and U8496 (N_8496,N_8388,N_8319);
xnor U8497 (N_8497,N_8396,N_8302);
nand U8498 (N_8498,N_8360,N_8306);
xnor U8499 (N_8499,N_8312,N_8372);
nor U8500 (N_8500,N_8471,N_8414);
nand U8501 (N_8501,N_8437,N_8492);
nor U8502 (N_8502,N_8445,N_8451);
nand U8503 (N_8503,N_8409,N_8487);
or U8504 (N_8504,N_8431,N_8490);
and U8505 (N_8505,N_8491,N_8461);
or U8506 (N_8506,N_8436,N_8438);
nor U8507 (N_8507,N_8469,N_8433);
and U8508 (N_8508,N_8428,N_8413);
or U8509 (N_8509,N_8483,N_8486);
nand U8510 (N_8510,N_8476,N_8410);
xor U8511 (N_8511,N_8408,N_8411);
and U8512 (N_8512,N_8432,N_8426);
or U8513 (N_8513,N_8478,N_8412);
and U8514 (N_8514,N_8488,N_8425);
or U8515 (N_8515,N_8463,N_8480);
and U8516 (N_8516,N_8498,N_8443);
or U8517 (N_8517,N_8423,N_8434);
nor U8518 (N_8518,N_8406,N_8401);
xnor U8519 (N_8519,N_8446,N_8450);
and U8520 (N_8520,N_8477,N_8493);
or U8521 (N_8521,N_8427,N_8462);
nor U8522 (N_8522,N_8489,N_8472);
xor U8523 (N_8523,N_8466,N_8497);
nand U8524 (N_8524,N_8459,N_8465);
or U8525 (N_8525,N_8407,N_8415);
xnor U8526 (N_8526,N_8479,N_8424);
or U8527 (N_8527,N_8468,N_8481);
nand U8528 (N_8528,N_8447,N_8470);
nand U8529 (N_8529,N_8499,N_8454);
xor U8530 (N_8530,N_8473,N_8441);
xor U8531 (N_8531,N_8418,N_8405);
nand U8532 (N_8532,N_8458,N_8484);
nor U8533 (N_8533,N_8435,N_8402);
and U8534 (N_8534,N_8467,N_8482);
xnor U8535 (N_8535,N_8457,N_8456);
or U8536 (N_8536,N_8494,N_8430);
or U8537 (N_8537,N_8448,N_8460);
xor U8538 (N_8538,N_8485,N_8421);
and U8539 (N_8539,N_8439,N_8419);
or U8540 (N_8540,N_8403,N_8420);
nand U8541 (N_8541,N_8400,N_8442);
nor U8542 (N_8542,N_8464,N_8404);
xor U8543 (N_8543,N_8455,N_8449);
and U8544 (N_8544,N_8474,N_8496);
xnor U8545 (N_8545,N_8453,N_8495);
xor U8546 (N_8546,N_8440,N_8422);
xnor U8547 (N_8547,N_8444,N_8417);
nand U8548 (N_8548,N_8429,N_8475);
or U8549 (N_8549,N_8452,N_8416);
nor U8550 (N_8550,N_8481,N_8466);
or U8551 (N_8551,N_8407,N_8483);
and U8552 (N_8552,N_8431,N_8478);
nor U8553 (N_8553,N_8424,N_8469);
and U8554 (N_8554,N_8408,N_8487);
nor U8555 (N_8555,N_8474,N_8411);
xnor U8556 (N_8556,N_8493,N_8481);
xor U8557 (N_8557,N_8454,N_8444);
and U8558 (N_8558,N_8416,N_8489);
xnor U8559 (N_8559,N_8486,N_8484);
or U8560 (N_8560,N_8443,N_8442);
nor U8561 (N_8561,N_8435,N_8410);
xnor U8562 (N_8562,N_8465,N_8454);
nand U8563 (N_8563,N_8459,N_8411);
and U8564 (N_8564,N_8474,N_8448);
and U8565 (N_8565,N_8465,N_8495);
nand U8566 (N_8566,N_8447,N_8417);
xnor U8567 (N_8567,N_8421,N_8481);
nand U8568 (N_8568,N_8460,N_8485);
nor U8569 (N_8569,N_8426,N_8456);
and U8570 (N_8570,N_8423,N_8478);
nand U8571 (N_8571,N_8493,N_8471);
nor U8572 (N_8572,N_8440,N_8408);
or U8573 (N_8573,N_8481,N_8458);
or U8574 (N_8574,N_8490,N_8459);
and U8575 (N_8575,N_8422,N_8478);
xor U8576 (N_8576,N_8491,N_8453);
nand U8577 (N_8577,N_8494,N_8438);
nand U8578 (N_8578,N_8460,N_8447);
and U8579 (N_8579,N_8418,N_8491);
xnor U8580 (N_8580,N_8489,N_8490);
nand U8581 (N_8581,N_8400,N_8495);
nor U8582 (N_8582,N_8498,N_8442);
xor U8583 (N_8583,N_8469,N_8458);
nand U8584 (N_8584,N_8481,N_8492);
or U8585 (N_8585,N_8460,N_8438);
nand U8586 (N_8586,N_8470,N_8401);
nand U8587 (N_8587,N_8416,N_8426);
xnor U8588 (N_8588,N_8407,N_8464);
xnor U8589 (N_8589,N_8408,N_8416);
and U8590 (N_8590,N_8437,N_8425);
and U8591 (N_8591,N_8402,N_8424);
and U8592 (N_8592,N_8489,N_8469);
xnor U8593 (N_8593,N_8437,N_8403);
or U8594 (N_8594,N_8457,N_8492);
or U8595 (N_8595,N_8461,N_8410);
xnor U8596 (N_8596,N_8476,N_8470);
and U8597 (N_8597,N_8492,N_8488);
and U8598 (N_8598,N_8448,N_8445);
nor U8599 (N_8599,N_8406,N_8430);
xor U8600 (N_8600,N_8581,N_8515);
nand U8601 (N_8601,N_8502,N_8565);
nor U8602 (N_8602,N_8504,N_8591);
nand U8603 (N_8603,N_8508,N_8523);
xnor U8604 (N_8604,N_8528,N_8570);
xnor U8605 (N_8605,N_8595,N_8536);
and U8606 (N_8606,N_8586,N_8519);
xor U8607 (N_8607,N_8525,N_8532);
xor U8608 (N_8608,N_8563,N_8544);
nand U8609 (N_8609,N_8553,N_8548);
and U8610 (N_8610,N_8514,N_8557);
xnor U8611 (N_8611,N_8538,N_8590);
and U8612 (N_8612,N_8535,N_8543);
and U8613 (N_8613,N_8594,N_8583);
nor U8614 (N_8614,N_8593,N_8509);
and U8615 (N_8615,N_8556,N_8559);
xor U8616 (N_8616,N_8571,N_8524);
and U8617 (N_8617,N_8577,N_8513);
xor U8618 (N_8618,N_8546,N_8561);
or U8619 (N_8619,N_8578,N_8575);
or U8620 (N_8620,N_8501,N_8547);
nor U8621 (N_8621,N_8511,N_8506);
or U8622 (N_8622,N_8589,N_8555);
nand U8623 (N_8623,N_8566,N_8564);
xor U8624 (N_8624,N_8598,N_8584);
or U8625 (N_8625,N_8526,N_8579);
and U8626 (N_8626,N_8517,N_8510);
nor U8627 (N_8627,N_8596,N_8542);
and U8628 (N_8628,N_8537,N_8560);
xnor U8629 (N_8629,N_8568,N_8585);
nor U8630 (N_8630,N_8530,N_8567);
nand U8631 (N_8631,N_8522,N_8539);
nor U8632 (N_8632,N_8533,N_8576);
or U8633 (N_8633,N_8588,N_8554);
nand U8634 (N_8634,N_8500,N_8580);
xnor U8635 (N_8635,N_8541,N_8512);
and U8636 (N_8636,N_8540,N_8550);
and U8637 (N_8637,N_8572,N_8587);
xor U8638 (N_8638,N_8549,N_8520);
or U8639 (N_8639,N_8599,N_8582);
nand U8640 (N_8640,N_8531,N_8558);
nor U8641 (N_8641,N_8527,N_8518);
or U8642 (N_8642,N_8562,N_8503);
nand U8643 (N_8643,N_8534,N_8574);
and U8644 (N_8644,N_8545,N_8573);
and U8645 (N_8645,N_8505,N_8507);
nor U8646 (N_8646,N_8516,N_8597);
xnor U8647 (N_8647,N_8529,N_8552);
and U8648 (N_8648,N_8521,N_8551);
nor U8649 (N_8649,N_8569,N_8592);
nand U8650 (N_8650,N_8511,N_8554);
or U8651 (N_8651,N_8578,N_8501);
or U8652 (N_8652,N_8571,N_8539);
and U8653 (N_8653,N_8541,N_8579);
xor U8654 (N_8654,N_8599,N_8500);
nor U8655 (N_8655,N_8562,N_8533);
and U8656 (N_8656,N_8569,N_8541);
nand U8657 (N_8657,N_8539,N_8565);
or U8658 (N_8658,N_8572,N_8563);
and U8659 (N_8659,N_8586,N_8553);
or U8660 (N_8660,N_8525,N_8502);
and U8661 (N_8661,N_8540,N_8560);
nor U8662 (N_8662,N_8530,N_8598);
or U8663 (N_8663,N_8534,N_8568);
nand U8664 (N_8664,N_8597,N_8566);
and U8665 (N_8665,N_8510,N_8593);
xor U8666 (N_8666,N_8501,N_8572);
nor U8667 (N_8667,N_8550,N_8530);
and U8668 (N_8668,N_8582,N_8529);
or U8669 (N_8669,N_8568,N_8513);
xor U8670 (N_8670,N_8591,N_8553);
xor U8671 (N_8671,N_8580,N_8573);
nand U8672 (N_8672,N_8555,N_8502);
and U8673 (N_8673,N_8523,N_8558);
xnor U8674 (N_8674,N_8526,N_8587);
nor U8675 (N_8675,N_8561,N_8566);
nor U8676 (N_8676,N_8551,N_8505);
nor U8677 (N_8677,N_8538,N_8518);
xor U8678 (N_8678,N_8501,N_8545);
and U8679 (N_8679,N_8517,N_8508);
and U8680 (N_8680,N_8531,N_8552);
and U8681 (N_8681,N_8566,N_8565);
nor U8682 (N_8682,N_8588,N_8575);
nor U8683 (N_8683,N_8502,N_8505);
xor U8684 (N_8684,N_8505,N_8511);
nand U8685 (N_8685,N_8591,N_8561);
nor U8686 (N_8686,N_8552,N_8585);
nand U8687 (N_8687,N_8575,N_8590);
and U8688 (N_8688,N_8584,N_8560);
xor U8689 (N_8689,N_8502,N_8526);
xor U8690 (N_8690,N_8597,N_8537);
nor U8691 (N_8691,N_8516,N_8590);
nor U8692 (N_8692,N_8505,N_8574);
nand U8693 (N_8693,N_8563,N_8587);
and U8694 (N_8694,N_8516,N_8545);
nand U8695 (N_8695,N_8582,N_8507);
and U8696 (N_8696,N_8546,N_8596);
or U8697 (N_8697,N_8581,N_8500);
xor U8698 (N_8698,N_8539,N_8579);
xnor U8699 (N_8699,N_8583,N_8518);
xor U8700 (N_8700,N_8685,N_8661);
or U8701 (N_8701,N_8645,N_8682);
xor U8702 (N_8702,N_8670,N_8694);
nor U8703 (N_8703,N_8633,N_8699);
xnor U8704 (N_8704,N_8695,N_8627);
xor U8705 (N_8705,N_8696,N_8632);
nand U8706 (N_8706,N_8642,N_8604);
nor U8707 (N_8707,N_8610,N_8637);
and U8708 (N_8708,N_8629,N_8617);
nor U8709 (N_8709,N_8673,N_8601);
and U8710 (N_8710,N_8666,N_8687);
xor U8711 (N_8711,N_8644,N_8691);
xnor U8712 (N_8712,N_8609,N_8669);
or U8713 (N_8713,N_8663,N_8603);
and U8714 (N_8714,N_8650,N_8636);
or U8715 (N_8715,N_8635,N_8657);
nor U8716 (N_8716,N_8693,N_8697);
or U8717 (N_8717,N_8660,N_8647);
and U8718 (N_8718,N_8656,N_8643);
nor U8719 (N_8719,N_8634,N_8622);
nor U8720 (N_8720,N_8676,N_8698);
nor U8721 (N_8721,N_8654,N_8607);
and U8722 (N_8722,N_8619,N_8688);
or U8723 (N_8723,N_8648,N_8625);
xor U8724 (N_8724,N_8628,N_8683);
nand U8725 (N_8725,N_8600,N_8606);
nor U8726 (N_8726,N_8659,N_8630);
xor U8727 (N_8727,N_8689,N_8646);
and U8728 (N_8728,N_8658,N_8655);
and U8729 (N_8729,N_8616,N_8678);
xor U8730 (N_8730,N_8608,N_8690);
nor U8731 (N_8731,N_8671,N_8624);
nor U8732 (N_8732,N_8612,N_8649);
nor U8733 (N_8733,N_8602,N_8684);
nand U8734 (N_8734,N_8653,N_8651);
or U8735 (N_8735,N_8640,N_8638);
and U8736 (N_8736,N_8611,N_8639);
nand U8737 (N_8737,N_8686,N_8621);
or U8738 (N_8738,N_8613,N_8680);
nand U8739 (N_8739,N_8641,N_8674);
or U8740 (N_8740,N_8677,N_8620);
nand U8741 (N_8741,N_8662,N_8615);
or U8742 (N_8742,N_8631,N_8614);
xnor U8743 (N_8743,N_8679,N_8692);
and U8744 (N_8744,N_8665,N_8626);
and U8745 (N_8745,N_8664,N_8672);
xor U8746 (N_8746,N_8618,N_8667);
and U8747 (N_8747,N_8681,N_8675);
or U8748 (N_8748,N_8668,N_8605);
nand U8749 (N_8749,N_8623,N_8652);
or U8750 (N_8750,N_8626,N_8612);
and U8751 (N_8751,N_8641,N_8684);
nand U8752 (N_8752,N_8698,N_8680);
nor U8753 (N_8753,N_8621,N_8600);
nor U8754 (N_8754,N_8655,N_8605);
and U8755 (N_8755,N_8617,N_8690);
and U8756 (N_8756,N_8638,N_8641);
or U8757 (N_8757,N_8692,N_8652);
or U8758 (N_8758,N_8656,N_8606);
nand U8759 (N_8759,N_8625,N_8619);
nand U8760 (N_8760,N_8680,N_8604);
nor U8761 (N_8761,N_8641,N_8647);
nor U8762 (N_8762,N_8622,N_8656);
xor U8763 (N_8763,N_8642,N_8618);
or U8764 (N_8764,N_8665,N_8623);
and U8765 (N_8765,N_8653,N_8698);
xnor U8766 (N_8766,N_8635,N_8656);
nor U8767 (N_8767,N_8661,N_8656);
or U8768 (N_8768,N_8634,N_8658);
and U8769 (N_8769,N_8612,N_8608);
xor U8770 (N_8770,N_8623,N_8609);
and U8771 (N_8771,N_8613,N_8630);
or U8772 (N_8772,N_8631,N_8630);
xor U8773 (N_8773,N_8606,N_8636);
nand U8774 (N_8774,N_8646,N_8694);
nor U8775 (N_8775,N_8697,N_8694);
nand U8776 (N_8776,N_8680,N_8656);
and U8777 (N_8777,N_8688,N_8604);
nand U8778 (N_8778,N_8689,N_8628);
or U8779 (N_8779,N_8601,N_8694);
or U8780 (N_8780,N_8637,N_8626);
or U8781 (N_8781,N_8640,N_8657);
nand U8782 (N_8782,N_8600,N_8693);
xor U8783 (N_8783,N_8670,N_8696);
nand U8784 (N_8784,N_8625,N_8642);
or U8785 (N_8785,N_8666,N_8649);
nand U8786 (N_8786,N_8602,N_8607);
nor U8787 (N_8787,N_8627,N_8681);
xor U8788 (N_8788,N_8621,N_8604);
or U8789 (N_8789,N_8616,N_8636);
nand U8790 (N_8790,N_8626,N_8643);
or U8791 (N_8791,N_8620,N_8696);
nand U8792 (N_8792,N_8687,N_8608);
nor U8793 (N_8793,N_8685,N_8624);
nand U8794 (N_8794,N_8605,N_8645);
and U8795 (N_8795,N_8636,N_8691);
and U8796 (N_8796,N_8642,N_8689);
xnor U8797 (N_8797,N_8680,N_8692);
xor U8798 (N_8798,N_8618,N_8698);
or U8799 (N_8799,N_8664,N_8681);
nor U8800 (N_8800,N_8717,N_8765);
nand U8801 (N_8801,N_8787,N_8785);
and U8802 (N_8802,N_8732,N_8792);
nand U8803 (N_8803,N_8788,N_8790);
and U8804 (N_8804,N_8754,N_8796);
nand U8805 (N_8805,N_8798,N_8704);
nand U8806 (N_8806,N_8728,N_8745);
nor U8807 (N_8807,N_8784,N_8725);
and U8808 (N_8808,N_8703,N_8752);
nand U8809 (N_8809,N_8780,N_8778);
nor U8810 (N_8810,N_8773,N_8701);
and U8811 (N_8811,N_8768,N_8791);
xor U8812 (N_8812,N_8781,N_8709);
or U8813 (N_8813,N_8748,N_8715);
xor U8814 (N_8814,N_8731,N_8736);
nor U8815 (N_8815,N_8740,N_8708);
xor U8816 (N_8816,N_8705,N_8774);
nand U8817 (N_8817,N_8751,N_8795);
nor U8818 (N_8818,N_8770,N_8720);
or U8819 (N_8819,N_8783,N_8702);
and U8820 (N_8820,N_8775,N_8743);
xor U8821 (N_8821,N_8746,N_8713);
and U8822 (N_8822,N_8757,N_8733);
nand U8823 (N_8823,N_8742,N_8706);
nor U8824 (N_8824,N_8716,N_8749);
nand U8825 (N_8825,N_8750,N_8777);
or U8826 (N_8826,N_8799,N_8739);
nor U8827 (N_8827,N_8729,N_8797);
xor U8828 (N_8828,N_8734,N_8714);
nor U8829 (N_8829,N_8730,N_8789);
xor U8830 (N_8830,N_8772,N_8753);
and U8831 (N_8831,N_8737,N_8744);
and U8832 (N_8832,N_8759,N_8710);
xor U8833 (N_8833,N_8779,N_8794);
and U8834 (N_8834,N_8700,N_8776);
nand U8835 (N_8835,N_8763,N_8723);
or U8836 (N_8836,N_8711,N_8726);
nor U8837 (N_8837,N_8762,N_8719);
and U8838 (N_8838,N_8755,N_8712);
xor U8839 (N_8839,N_8760,N_8756);
or U8840 (N_8840,N_8741,N_8782);
nand U8841 (N_8841,N_8724,N_8718);
nand U8842 (N_8842,N_8707,N_8764);
nand U8843 (N_8843,N_8769,N_8761);
xor U8844 (N_8844,N_8735,N_8758);
xnor U8845 (N_8845,N_8793,N_8722);
xnor U8846 (N_8846,N_8786,N_8766);
nand U8847 (N_8847,N_8767,N_8721);
nand U8848 (N_8848,N_8771,N_8738);
or U8849 (N_8849,N_8747,N_8727);
nand U8850 (N_8850,N_8763,N_8796);
xnor U8851 (N_8851,N_8747,N_8760);
nor U8852 (N_8852,N_8724,N_8748);
and U8853 (N_8853,N_8796,N_8732);
nand U8854 (N_8854,N_8773,N_8765);
nand U8855 (N_8855,N_8745,N_8789);
nor U8856 (N_8856,N_8785,N_8741);
xnor U8857 (N_8857,N_8759,N_8729);
nand U8858 (N_8858,N_8762,N_8723);
and U8859 (N_8859,N_8740,N_8722);
and U8860 (N_8860,N_8736,N_8799);
xor U8861 (N_8861,N_8772,N_8729);
and U8862 (N_8862,N_8747,N_8768);
nand U8863 (N_8863,N_8785,N_8798);
and U8864 (N_8864,N_8798,N_8730);
or U8865 (N_8865,N_8719,N_8771);
or U8866 (N_8866,N_8722,N_8732);
nor U8867 (N_8867,N_8791,N_8728);
nand U8868 (N_8868,N_8722,N_8748);
nand U8869 (N_8869,N_8756,N_8714);
nor U8870 (N_8870,N_8719,N_8736);
nand U8871 (N_8871,N_8757,N_8735);
and U8872 (N_8872,N_8739,N_8743);
nand U8873 (N_8873,N_8775,N_8732);
or U8874 (N_8874,N_8737,N_8712);
and U8875 (N_8875,N_8775,N_8741);
nand U8876 (N_8876,N_8796,N_8722);
and U8877 (N_8877,N_8701,N_8793);
and U8878 (N_8878,N_8735,N_8766);
xnor U8879 (N_8879,N_8759,N_8742);
nor U8880 (N_8880,N_8732,N_8728);
xor U8881 (N_8881,N_8748,N_8735);
or U8882 (N_8882,N_8762,N_8737);
or U8883 (N_8883,N_8757,N_8722);
nand U8884 (N_8884,N_8724,N_8791);
or U8885 (N_8885,N_8746,N_8719);
and U8886 (N_8886,N_8728,N_8797);
xnor U8887 (N_8887,N_8750,N_8760);
xor U8888 (N_8888,N_8708,N_8763);
and U8889 (N_8889,N_8704,N_8719);
or U8890 (N_8890,N_8738,N_8725);
and U8891 (N_8891,N_8752,N_8778);
nor U8892 (N_8892,N_8754,N_8767);
xor U8893 (N_8893,N_8799,N_8704);
nor U8894 (N_8894,N_8753,N_8782);
xnor U8895 (N_8895,N_8704,N_8740);
nand U8896 (N_8896,N_8716,N_8725);
and U8897 (N_8897,N_8728,N_8741);
nor U8898 (N_8898,N_8715,N_8757);
nor U8899 (N_8899,N_8797,N_8710);
xor U8900 (N_8900,N_8832,N_8882);
nand U8901 (N_8901,N_8828,N_8874);
nor U8902 (N_8902,N_8897,N_8857);
nor U8903 (N_8903,N_8837,N_8886);
and U8904 (N_8904,N_8804,N_8896);
nand U8905 (N_8905,N_8800,N_8820);
xor U8906 (N_8906,N_8872,N_8818);
and U8907 (N_8907,N_8878,N_8834);
xor U8908 (N_8908,N_8885,N_8843);
xnor U8909 (N_8909,N_8825,N_8803);
or U8910 (N_8910,N_8892,N_8809);
nor U8911 (N_8911,N_8869,N_8893);
or U8912 (N_8912,N_8889,N_8830);
xor U8913 (N_8913,N_8819,N_8852);
and U8914 (N_8914,N_8823,N_8840);
nand U8915 (N_8915,N_8833,N_8801);
and U8916 (N_8916,N_8890,N_8812);
nand U8917 (N_8917,N_8854,N_8887);
and U8918 (N_8918,N_8868,N_8891);
and U8919 (N_8919,N_8899,N_8876);
nand U8920 (N_8920,N_8814,N_8849);
or U8921 (N_8921,N_8846,N_8850);
and U8922 (N_8922,N_8895,N_8806);
or U8923 (N_8923,N_8827,N_8802);
or U8924 (N_8924,N_8861,N_8863);
nand U8925 (N_8925,N_8829,N_8859);
nand U8926 (N_8926,N_8821,N_8848);
nand U8927 (N_8927,N_8805,N_8844);
xor U8928 (N_8928,N_8815,N_8879);
and U8929 (N_8929,N_8888,N_8842);
nor U8930 (N_8930,N_8894,N_8813);
and U8931 (N_8931,N_8875,N_8867);
and U8932 (N_8932,N_8826,N_8880);
xor U8933 (N_8933,N_8847,N_8871);
and U8934 (N_8934,N_8831,N_8810);
nand U8935 (N_8935,N_8862,N_8811);
nor U8936 (N_8936,N_8864,N_8838);
nor U8937 (N_8937,N_8881,N_8877);
and U8938 (N_8938,N_8855,N_8858);
xor U8939 (N_8939,N_8873,N_8808);
or U8940 (N_8940,N_8884,N_8839);
or U8941 (N_8941,N_8865,N_8807);
nand U8942 (N_8942,N_8845,N_8824);
nor U8943 (N_8943,N_8841,N_8817);
or U8944 (N_8944,N_8835,N_8822);
nand U8945 (N_8945,N_8860,N_8816);
or U8946 (N_8946,N_8836,N_8856);
nor U8947 (N_8947,N_8870,N_8853);
nand U8948 (N_8948,N_8866,N_8898);
or U8949 (N_8949,N_8851,N_8883);
xor U8950 (N_8950,N_8832,N_8855);
nand U8951 (N_8951,N_8870,N_8866);
and U8952 (N_8952,N_8890,N_8813);
and U8953 (N_8953,N_8878,N_8856);
xnor U8954 (N_8954,N_8875,N_8876);
nor U8955 (N_8955,N_8829,N_8804);
nor U8956 (N_8956,N_8895,N_8844);
or U8957 (N_8957,N_8828,N_8803);
nand U8958 (N_8958,N_8878,N_8861);
or U8959 (N_8959,N_8824,N_8855);
or U8960 (N_8960,N_8856,N_8825);
nand U8961 (N_8961,N_8871,N_8876);
or U8962 (N_8962,N_8814,N_8853);
or U8963 (N_8963,N_8846,N_8829);
and U8964 (N_8964,N_8859,N_8848);
nor U8965 (N_8965,N_8846,N_8852);
and U8966 (N_8966,N_8870,N_8832);
nand U8967 (N_8967,N_8818,N_8866);
nand U8968 (N_8968,N_8850,N_8874);
and U8969 (N_8969,N_8800,N_8877);
nand U8970 (N_8970,N_8870,N_8883);
nand U8971 (N_8971,N_8807,N_8846);
or U8972 (N_8972,N_8853,N_8806);
xor U8973 (N_8973,N_8887,N_8823);
nor U8974 (N_8974,N_8820,N_8819);
and U8975 (N_8975,N_8864,N_8861);
or U8976 (N_8976,N_8850,N_8849);
and U8977 (N_8977,N_8846,N_8819);
xnor U8978 (N_8978,N_8876,N_8854);
or U8979 (N_8979,N_8800,N_8810);
and U8980 (N_8980,N_8875,N_8807);
xnor U8981 (N_8981,N_8843,N_8897);
nor U8982 (N_8982,N_8838,N_8827);
nand U8983 (N_8983,N_8874,N_8882);
nor U8984 (N_8984,N_8898,N_8805);
or U8985 (N_8985,N_8821,N_8891);
or U8986 (N_8986,N_8838,N_8839);
or U8987 (N_8987,N_8867,N_8804);
xor U8988 (N_8988,N_8805,N_8861);
or U8989 (N_8989,N_8882,N_8875);
or U8990 (N_8990,N_8855,N_8867);
nor U8991 (N_8991,N_8886,N_8883);
xor U8992 (N_8992,N_8896,N_8868);
nand U8993 (N_8993,N_8856,N_8847);
or U8994 (N_8994,N_8805,N_8813);
xnor U8995 (N_8995,N_8832,N_8878);
or U8996 (N_8996,N_8853,N_8871);
xnor U8997 (N_8997,N_8851,N_8849);
xnor U8998 (N_8998,N_8881,N_8899);
or U8999 (N_8999,N_8832,N_8816);
xor U9000 (N_9000,N_8982,N_8922);
xnor U9001 (N_9001,N_8985,N_8908);
nand U9002 (N_9002,N_8954,N_8980);
and U9003 (N_9003,N_8920,N_8935);
xor U9004 (N_9004,N_8939,N_8961);
xnor U9005 (N_9005,N_8928,N_8962);
nand U9006 (N_9006,N_8904,N_8917);
nand U9007 (N_9007,N_8931,N_8909);
nor U9008 (N_9008,N_8990,N_8944);
or U9009 (N_9009,N_8941,N_8978);
or U9010 (N_9010,N_8993,N_8923);
nand U9011 (N_9011,N_8948,N_8988);
and U9012 (N_9012,N_8996,N_8919);
and U9013 (N_9013,N_8946,N_8938);
and U9014 (N_9014,N_8976,N_8975);
nor U9015 (N_9015,N_8950,N_8907);
and U9016 (N_9016,N_8927,N_8963);
or U9017 (N_9017,N_8957,N_8958);
nand U9018 (N_9018,N_8971,N_8966);
nor U9019 (N_9019,N_8910,N_8952);
xor U9020 (N_9020,N_8979,N_8949);
nand U9021 (N_9021,N_8986,N_8967);
and U9022 (N_9022,N_8959,N_8900);
and U9023 (N_9023,N_8921,N_8987);
xor U9024 (N_9024,N_8911,N_8955);
nand U9025 (N_9025,N_8997,N_8947);
xor U9026 (N_9026,N_8960,N_8972);
and U9027 (N_9027,N_8964,N_8951);
nor U9028 (N_9028,N_8969,N_8973);
xnor U9029 (N_9029,N_8977,N_8906);
xnor U9030 (N_9030,N_8995,N_8940);
or U9031 (N_9031,N_8924,N_8915);
or U9032 (N_9032,N_8981,N_8933);
and U9033 (N_9033,N_8998,N_8991);
and U9034 (N_9034,N_8932,N_8925);
or U9035 (N_9035,N_8914,N_8970);
nand U9036 (N_9036,N_8930,N_8994);
nand U9037 (N_9037,N_8984,N_8934);
xnor U9038 (N_9038,N_8983,N_8903);
or U9039 (N_9039,N_8956,N_8901);
nor U9040 (N_9040,N_8936,N_8943);
and U9041 (N_9041,N_8965,N_8945);
and U9042 (N_9042,N_8989,N_8918);
nand U9043 (N_9043,N_8916,N_8926);
or U9044 (N_9044,N_8953,N_8999);
or U9045 (N_9045,N_8942,N_8992);
xnor U9046 (N_9046,N_8937,N_8905);
or U9047 (N_9047,N_8974,N_8929);
or U9048 (N_9048,N_8912,N_8913);
and U9049 (N_9049,N_8902,N_8968);
xor U9050 (N_9050,N_8920,N_8931);
nand U9051 (N_9051,N_8912,N_8931);
xor U9052 (N_9052,N_8950,N_8981);
and U9053 (N_9053,N_8931,N_8918);
nand U9054 (N_9054,N_8986,N_8952);
and U9055 (N_9055,N_8975,N_8905);
or U9056 (N_9056,N_8954,N_8984);
or U9057 (N_9057,N_8916,N_8994);
or U9058 (N_9058,N_8909,N_8925);
xnor U9059 (N_9059,N_8946,N_8931);
xnor U9060 (N_9060,N_8948,N_8981);
or U9061 (N_9061,N_8990,N_8930);
xnor U9062 (N_9062,N_8916,N_8935);
xor U9063 (N_9063,N_8917,N_8910);
nor U9064 (N_9064,N_8965,N_8914);
nor U9065 (N_9065,N_8906,N_8920);
xnor U9066 (N_9066,N_8960,N_8967);
xnor U9067 (N_9067,N_8995,N_8941);
xor U9068 (N_9068,N_8981,N_8991);
nand U9069 (N_9069,N_8975,N_8938);
nor U9070 (N_9070,N_8944,N_8983);
and U9071 (N_9071,N_8969,N_8941);
nor U9072 (N_9072,N_8997,N_8998);
or U9073 (N_9073,N_8982,N_8930);
nor U9074 (N_9074,N_8995,N_8930);
xor U9075 (N_9075,N_8938,N_8912);
nand U9076 (N_9076,N_8933,N_8965);
nor U9077 (N_9077,N_8980,N_8957);
xor U9078 (N_9078,N_8954,N_8995);
and U9079 (N_9079,N_8925,N_8934);
and U9080 (N_9080,N_8902,N_8907);
nand U9081 (N_9081,N_8977,N_8995);
nand U9082 (N_9082,N_8919,N_8907);
or U9083 (N_9083,N_8979,N_8917);
nand U9084 (N_9084,N_8953,N_8933);
nand U9085 (N_9085,N_8982,N_8960);
or U9086 (N_9086,N_8939,N_8959);
nor U9087 (N_9087,N_8901,N_8974);
nand U9088 (N_9088,N_8966,N_8997);
and U9089 (N_9089,N_8975,N_8969);
xor U9090 (N_9090,N_8988,N_8946);
and U9091 (N_9091,N_8932,N_8965);
xor U9092 (N_9092,N_8922,N_8949);
xnor U9093 (N_9093,N_8963,N_8991);
or U9094 (N_9094,N_8935,N_8989);
xor U9095 (N_9095,N_8949,N_8997);
nor U9096 (N_9096,N_8942,N_8964);
xnor U9097 (N_9097,N_8984,N_8959);
xnor U9098 (N_9098,N_8902,N_8998);
nand U9099 (N_9099,N_8963,N_8956);
nor U9100 (N_9100,N_9098,N_9064);
and U9101 (N_9101,N_9099,N_9044);
or U9102 (N_9102,N_9032,N_9034);
nor U9103 (N_9103,N_9095,N_9008);
and U9104 (N_9104,N_9009,N_9058);
or U9105 (N_9105,N_9025,N_9083);
or U9106 (N_9106,N_9087,N_9074);
xor U9107 (N_9107,N_9049,N_9068);
nand U9108 (N_9108,N_9026,N_9002);
xor U9109 (N_9109,N_9051,N_9062);
or U9110 (N_9110,N_9045,N_9091);
nor U9111 (N_9111,N_9006,N_9080);
xnor U9112 (N_9112,N_9007,N_9043);
or U9113 (N_9113,N_9097,N_9057);
nor U9114 (N_9114,N_9081,N_9016);
and U9115 (N_9115,N_9076,N_9060);
and U9116 (N_9116,N_9048,N_9023);
xnor U9117 (N_9117,N_9029,N_9077);
xor U9118 (N_9118,N_9031,N_9092);
or U9119 (N_9119,N_9052,N_9038);
nor U9120 (N_9120,N_9072,N_9088);
nor U9121 (N_9121,N_9030,N_9078);
and U9122 (N_9122,N_9020,N_9035);
nand U9123 (N_9123,N_9096,N_9073);
or U9124 (N_9124,N_9066,N_9012);
and U9125 (N_9125,N_9063,N_9089);
and U9126 (N_9126,N_9090,N_9069);
or U9127 (N_9127,N_9005,N_9041);
or U9128 (N_9128,N_9071,N_9014);
or U9129 (N_9129,N_9011,N_9028);
nor U9130 (N_9130,N_9070,N_9003);
or U9131 (N_9131,N_9067,N_9054);
or U9132 (N_9132,N_9065,N_9018);
xor U9133 (N_9133,N_9017,N_9053);
nor U9134 (N_9134,N_9010,N_9050);
xor U9135 (N_9135,N_9042,N_9093);
or U9136 (N_9136,N_9013,N_9039);
nor U9137 (N_9137,N_9004,N_9040);
or U9138 (N_9138,N_9046,N_9047);
and U9139 (N_9139,N_9033,N_9015);
nand U9140 (N_9140,N_9022,N_9082);
and U9141 (N_9141,N_9027,N_9055);
or U9142 (N_9142,N_9086,N_9036);
and U9143 (N_9143,N_9037,N_9075);
and U9144 (N_9144,N_9084,N_9059);
nand U9145 (N_9145,N_9085,N_9061);
nand U9146 (N_9146,N_9001,N_9000);
nor U9147 (N_9147,N_9024,N_9019);
or U9148 (N_9148,N_9021,N_9056);
and U9149 (N_9149,N_9079,N_9094);
or U9150 (N_9150,N_9009,N_9096);
and U9151 (N_9151,N_9089,N_9064);
or U9152 (N_9152,N_9095,N_9028);
nand U9153 (N_9153,N_9024,N_9039);
nor U9154 (N_9154,N_9082,N_9071);
and U9155 (N_9155,N_9046,N_9048);
xnor U9156 (N_9156,N_9052,N_9089);
nor U9157 (N_9157,N_9077,N_9000);
and U9158 (N_9158,N_9092,N_9023);
and U9159 (N_9159,N_9031,N_9089);
xnor U9160 (N_9160,N_9046,N_9043);
nor U9161 (N_9161,N_9063,N_9008);
xnor U9162 (N_9162,N_9083,N_9064);
xnor U9163 (N_9163,N_9091,N_9028);
nand U9164 (N_9164,N_9057,N_9042);
and U9165 (N_9165,N_9070,N_9018);
xor U9166 (N_9166,N_9081,N_9023);
and U9167 (N_9167,N_9094,N_9046);
or U9168 (N_9168,N_9011,N_9051);
nand U9169 (N_9169,N_9017,N_9034);
or U9170 (N_9170,N_9041,N_9010);
or U9171 (N_9171,N_9075,N_9033);
or U9172 (N_9172,N_9069,N_9077);
nand U9173 (N_9173,N_9071,N_9024);
and U9174 (N_9174,N_9027,N_9059);
nand U9175 (N_9175,N_9056,N_9034);
nor U9176 (N_9176,N_9021,N_9009);
and U9177 (N_9177,N_9006,N_9093);
nor U9178 (N_9178,N_9064,N_9010);
xnor U9179 (N_9179,N_9098,N_9042);
and U9180 (N_9180,N_9002,N_9030);
xor U9181 (N_9181,N_9089,N_9086);
or U9182 (N_9182,N_9043,N_9010);
or U9183 (N_9183,N_9019,N_9074);
nor U9184 (N_9184,N_9006,N_9091);
or U9185 (N_9185,N_9047,N_9056);
or U9186 (N_9186,N_9053,N_9014);
nor U9187 (N_9187,N_9068,N_9073);
nor U9188 (N_9188,N_9082,N_9006);
and U9189 (N_9189,N_9050,N_9060);
nand U9190 (N_9190,N_9094,N_9032);
xnor U9191 (N_9191,N_9087,N_9000);
xnor U9192 (N_9192,N_9091,N_9087);
nand U9193 (N_9193,N_9057,N_9015);
xnor U9194 (N_9194,N_9089,N_9005);
nand U9195 (N_9195,N_9004,N_9010);
or U9196 (N_9196,N_9033,N_9035);
nor U9197 (N_9197,N_9059,N_9039);
nor U9198 (N_9198,N_9004,N_9053);
nor U9199 (N_9199,N_9096,N_9061);
xnor U9200 (N_9200,N_9148,N_9181);
nand U9201 (N_9201,N_9143,N_9167);
and U9202 (N_9202,N_9191,N_9119);
nand U9203 (N_9203,N_9117,N_9190);
and U9204 (N_9204,N_9128,N_9171);
or U9205 (N_9205,N_9149,N_9194);
and U9206 (N_9206,N_9184,N_9193);
nand U9207 (N_9207,N_9140,N_9113);
nor U9208 (N_9208,N_9124,N_9129);
or U9209 (N_9209,N_9134,N_9125);
xor U9210 (N_9210,N_9195,N_9133);
or U9211 (N_9211,N_9139,N_9127);
and U9212 (N_9212,N_9155,N_9138);
xor U9213 (N_9213,N_9187,N_9110);
and U9214 (N_9214,N_9199,N_9192);
nand U9215 (N_9215,N_9183,N_9156);
and U9216 (N_9216,N_9111,N_9182);
and U9217 (N_9217,N_9176,N_9160);
nor U9218 (N_9218,N_9108,N_9109);
nor U9219 (N_9219,N_9141,N_9135);
nand U9220 (N_9220,N_9198,N_9137);
nand U9221 (N_9221,N_9112,N_9163);
and U9222 (N_9222,N_9179,N_9122);
and U9223 (N_9223,N_9115,N_9116);
xnor U9224 (N_9224,N_9150,N_9131);
xnor U9225 (N_9225,N_9174,N_9121);
nor U9226 (N_9226,N_9189,N_9114);
and U9227 (N_9227,N_9177,N_9132);
or U9228 (N_9228,N_9107,N_9197);
and U9229 (N_9229,N_9158,N_9180);
xnor U9230 (N_9230,N_9152,N_9142);
nand U9231 (N_9231,N_9157,N_9106);
or U9232 (N_9232,N_9168,N_9100);
and U9233 (N_9233,N_9162,N_9147);
and U9234 (N_9234,N_9105,N_9175);
xor U9235 (N_9235,N_9159,N_9136);
or U9236 (N_9236,N_9118,N_9169);
or U9237 (N_9237,N_9120,N_9186);
or U9238 (N_9238,N_9166,N_9102);
nor U9239 (N_9239,N_9161,N_9145);
or U9240 (N_9240,N_9123,N_9104);
xnor U9241 (N_9241,N_9173,N_9103);
nor U9242 (N_9242,N_9165,N_9188);
xor U9243 (N_9243,N_9178,N_9101);
nor U9244 (N_9244,N_9164,N_9170);
xor U9245 (N_9245,N_9185,N_9126);
xor U9246 (N_9246,N_9196,N_9130);
xnor U9247 (N_9247,N_9144,N_9151);
nand U9248 (N_9248,N_9172,N_9153);
nor U9249 (N_9249,N_9146,N_9154);
xnor U9250 (N_9250,N_9139,N_9142);
nand U9251 (N_9251,N_9130,N_9117);
and U9252 (N_9252,N_9179,N_9190);
and U9253 (N_9253,N_9195,N_9183);
and U9254 (N_9254,N_9196,N_9170);
or U9255 (N_9255,N_9122,N_9196);
xor U9256 (N_9256,N_9100,N_9125);
or U9257 (N_9257,N_9146,N_9128);
nor U9258 (N_9258,N_9152,N_9196);
xnor U9259 (N_9259,N_9136,N_9149);
xor U9260 (N_9260,N_9194,N_9161);
xnor U9261 (N_9261,N_9185,N_9109);
nor U9262 (N_9262,N_9107,N_9175);
or U9263 (N_9263,N_9103,N_9191);
xnor U9264 (N_9264,N_9156,N_9198);
nor U9265 (N_9265,N_9192,N_9182);
nor U9266 (N_9266,N_9142,N_9172);
and U9267 (N_9267,N_9174,N_9114);
xnor U9268 (N_9268,N_9167,N_9131);
nor U9269 (N_9269,N_9151,N_9108);
nor U9270 (N_9270,N_9177,N_9199);
xor U9271 (N_9271,N_9129,N_9149);
or U9272 (N_9272,N_9134,N_9174);
nor U9273 (N_9273,N_9161,N_9175);
xnor U9274 (N_9274,N_9167,N_9176);
or U9275 (N_9275,N_9104,N_9137);
or U9276 (N_9276,N_9104,N_9145);
and U9277 (N_9277,N_9118,N_9197);
xor U9278 (N_9278,N_9112,N_9171);
and U9279 (N_9279,N_9154,N_9162);
nor U9280 (N_9280,N_9148,N_9158);
nand U9281 (N_9281,N_9126,N_9168);
nand U9282 (N_9282,N_9173,N_9197);
and U9283 (N_9283,N_9131,N_9132);
nor U9284 (N_9284,N_9159,N_9199);
nor U9285 (N_9285,N_9155,N_9150);
nand U9286 (N_9286,N_9117,N_9178);
or U9287 (N_9287,N_9190,N_9121);
xnor U9288 (N_9288,N_9164,N_9184);
nor U9289 (N_9289,N_9132,N_9199);
or U9290 (N_9290,N_9177,N_9193);
or U9291 (N_9291,N_9165,N_9127);
nand U9292 (N_9292,N_9144,N_9189);
xnor U9293 (N_9293,N_9174,N_9188);
or U9294 (N_9294,N_9146,N_9193);
and U9295 (N_9295,N_9154,N_9176);
and U9296 (N_9296,N_9130,N_9167);
or U9297 (N_9297,N_9181,N_9141);
xnor U9298 (N_9298,N_9163,N_9140);
nor U9299 (N_9299,N_9157,N_9117);
and U9300 (N_9300,N_9237,N_9260);
nand U9301 (N_9301,N_9256,N_9243);
nor U9302 (N_9302,N_9239,N_9225);
nand U9303 (N_9303,N_9292,N_9207);
xor U9304 (N_9304,N_9214,N_9245);
xnor U9305 (N_9305,N_9252,N_9273);
and U9306 (N_9306,N_9262,N_9229);
and U9307 (N_9307,N_9209,N_9271);
and U9308 (N_9308,N_9253,N_9294);
or U9309 (N_9309,N_9238,N_9234);
or U9310 (N_9310,N_9230,N_9215);
nand U9311 (N_9311,N_9297,N_9200);
or U9312 (N_9312,N_9295,N_9250);
xor U9313 (N_9313,N_9290,N_9287);
nor U9314 (N_9314,N_9216,N_9274);
nand U9315 (N_9315,N_9280,N_9246);
xor U9316 (N_9316,N_9233,N_9220);
or U9317 (N_9317,N_9289,N_9281);
xor U9318 (N_9318,N_9244,N_9212);
and U9319 (N_9319,N_9240,N_9242);
nand U9320 (N_9320,N_9231,N_9276);
and U9321 (N_9321,N_9277,N_9226);
nand U9322 (N_9322,N_9232,N_9275);
xnor U9323 (N_9323,N_9266,N_9270);
nor U9324 (N_9324,N_9236,N_9223);
nor U9325 (N_9325,N_9286,N_9211);
nand U9326 (N_9326,N_9265,N_9248);
xnor U9327 (N_9327,N_9282,N_9278);
nand U9328 (N_9328,N_9217,N_9213);
or U9329 (N_9329,N_9247,N_9222);
nand U9330 (N_9330,N_9293,N_9299);
xor U9331 (N_9331,N_9206,N_9283);
nand U9332 (N_9332,N_9205,N_9259);
or U9333 (N_9333,N_9284,N_9224);
and U9334 (N_9334,N_9210,N_9269);
xor U9335 (N_9335,N_9208,N_9227);
or U9336 (N_9336,N_9267,N_9204);
nand U9337 (N_9337,N_9249,N_9298);
nor U9338 (N_9338,N_9218,N_9264);
or U9339 (N_9339,N_9268,N_9288);
nor U9340 (N_9340,N_9258,N_9285);
nor U9341 (N_9341,N_9251,N_9296);
xnor U9342 (N_9342,N_9272,N_9261);
or U9343 (N_9343,N_9202,N_9221);
xor U9344 (N_9344,N_9263,N_9279);
xnor U9345 (N_9345,N_9241,N_9228);
xor U9346 (N_9346,N_9219,N_9257);
nand U9347 (N_9347,N_9201,N_9291);
nor U9348 (N_9348,N_9235,N_9254);
nor U9349 (N_9349,N_9255,N_9203);
and U9350 (N_9350,N_9243,N_9228);
and U9351 (N_9351,N_9258,N_9273);
and U9352 (N_9352,N_9261,N_9244);
and U9353 (N_9353,N_9270,N_9222);
xor U9354 (N_9354,N_9200,N_9222);
xor U9355 (N_9355,N_9299,N_9241);
nor U9356 (N_9356,N_9242,N_9229);
and U9357 (N_9357,N_9276,N_9250);
and U9358 (N_9358,N_9210,N_9214);
and U9359 (N_9359,N_9209,N_9256);
and U9360 (N_9360,N_9244,N_9218);
or U9361 (N_9361,N_9294,N_9276);
or U9362 (N_9362,N_9260,N_9289);
and U9363 (N_9363,N_9209,N_9225);
xnor U9364 (N_9364,N_9231,N_9211);
xor U9365 (N_9365,N_9248,N_9256);
nor U9366 (N_9366,N_9272,N_9264);
nand U9367 (N_9367,N_9286,N_9202);
xor U9368 (N_9368,N_9214,N_9217);
nand U9369 (N_9369,N_9256,N_9278);
nand U9370 (N_9370,N_9296,N_9273);
nand U9371 (N_9371,N_9247,N_9210);
and U9372 (N_9372,N_9229,N_9249);
xnor U9373 (N_9373,N_9202,N_9287);
nand U9374 (N_9374,N_9283,N_9240);
nor U9375 (N_9375,N_9201,N_9298);
nand U9376 (N_9376,N_9245,N_9264);
or U9377 (N_9377,N_9287,N_9212);
and U9378 (N_9378,N_9244,N_9245);
xnor U9379 (N_9379,N_9258,N_9228);
nor U9380 (N_9380,N_9209,N_9215);
and U9381 (N_9381,N_9260,N_9231);
xnor U9382 (N_9382,N_9206,N_9233);
nand U9383 (N_9383,N_9209,N_9243);
or U9384 (N_9384,N_9210,N_9255);
nor U9385 (N_9385,N_9255,N_9276);
or U9386 (N_9386,N_9254,N_9237);
xor U9387 (N_9387,N_9215,N_9268);
nand U9388 (N_9388,N_9216,N_9298);
or U9389 (N_9389,N_9215,N_9241);
nor U9390 (N_9390,N_9292,N_9245);
or U9391 (N_9391,N_9286,N_9239);
xnor U9392 (N_9392,N_9292,N_9289);
nor U9393 (N_9393,N_9242,N_9232);
nand U9394 (N_9394,N_9207,N_9268);
nor U9395 (N_9395,N_9234,N_9231);
xnor U9396 (N_9396,N_9253,N_9224);
and U9397 (N_9397,N_9289,N_9218);
or U9398 (N_9398,N_9247,N_9224);
nor U9399 (N_9399,N_9232,N_9239);
xnor U9400 (N_9400,N_9388,N_9392);
nand U9401 (N_9401,N_9342,N_9318);
or U9402 (N_9402,N_9323,N_9390);
nand U9403 (N_9403,N_9383,N_9357);
and U9404 (N_9404,N_9393,N_9380);
nor U9405 (N_9405,N_9320,N_9302);
nor U9406 (N_9406,N_9365,N_9341);
nor U9407 (N_9407,N_9373,N_9321);
nor U9408 (N_9408,N_9315,N_9371);
and U9409 (N_9409,N_9361,N_9378);
xor U9410 (N_9410,N_9376,N_9329);
xor U9411 (N_9411,N_9384,N_9300);
or U9412 (N_9412,N_9386,N_9350);
or U9413 (N_9413,N_9353,N_9327);
nor U9414 (N_9414,N_9395,N_9344);
xor U9415 (N_9415,N_9348,N_9326);
and U9416 (N_9416,N_9338,N_9370);
xnor U9417 (N_9417,N_9312,N_9382);
or U9418 (N_9418,N_9359,N_9314);
xnor U9419 (N_9419,N_9304,N_9354);
nor U9420 (N_9420,N_9387,N_9328);
xor U9421 (N_9421,N_9345,N_9339);
or U9422 (N_9422,N_9319,N_9309);
and U9423 (N_9423,N_9349,N_9313);
or U9424 (N_9424,N_9351,N_9389);
nand U9425 (N_9425,N_9305,N_9301);
xnor U9426 (N_9426,N_9347,N_9363);
nand U9427 (N_9427,N_9358,N_9364);
and U9428 (N_9428,N_9385,N_9362);
nand U9429 (N_9429,N_9372,N_9391);
or U9430 (N_9430,N_9308,N_9346);
and U9431 (N_9431,N_9340,N_9332);
and U9432 (N_9432,N_9379,N_9306);
and U9433 (N_9433,N_9367,N_9375);
nand U9434 (N_9434,N_9352,N_9397);
and U9435 (N_9435,N_9355,N_9311);
and U9436 (N_9436,N_9398,N_9394);
nand U9437 (N_9437,N_9316,N_9356);
or U9438 (N_9438,N_9368,N_9374);
nor U9439 (N_9439,N_9399,N_9381);
and U9440 (N_9440,N_9334,N_9343);
and U9441 (N_9441,N_9366,N_9336);
xor U9442 (N_9442,N_9360,N_9303);
or U9443 (N_9443,N_9330,N_9322);
xnor U9444 (N_9444,N_9317,N_9310);
xnor U9445 (N_9445,N_9333,N_9337);
nand U9446 (N_9446,N_9377,N_9369);
nor U9447 (N_9447,N_9335,N_9396);
and U9448 (N_9448,N_9324,N_9307);
or U9449 (N_9449,N_9325,N_9331);
xnor U9450 (N_9450,N_9393,N_9342);
xnor U9451 (N_9451,N_9394,N_9316);
xor U9452 (N_9452,N_9364,N_9368);
nor U9453 (N_9453,N_9353,N_9348);
nor U9454 (N_9454,N_9344,N_9398);
nor U9455 (N_9455,N_9345,N_9350);
nand U9456 (N_9456,N_9365,N_9376);
and U9457 (N_9457,N_9390,N_9330);
or U9458 (N_9458,N_9381,N_9325);
or U9459 (N_9459,N_9346,N_9351);
xor U9460 (N_9460,N_9388,N_9394);
and U9461 (N_9461,N_9352,N_9362);
or U9462 (N_9462,N_9304,N_9367);
or U9463 (N_9463,N_9393,N_9324);
and U9464 (N_9464,N_9360,N_9367);
or U9465 (N_9465,N_9381,N_9320);
or U9466 (N_9466,N_9396,N_9334);
xnor U9467 (N_9467,N_9385,N_9306);
or U9468 (N_9468,N_9360,N_9371);
nand U9469 (N_9469,N_9300,N_9379);
nor U9470 (N_9470,N_9312,N_9399);
xor U9471 (N_9471,N_9398,N_9331);
nor U9472 (N_9472,N_9396,N_9364);
xnor U9473 (N_9473,N_9396,N_9357);
or U9474 (N_9474,N_9347,N_9301);
and U9475 (N_9475,N_9399,N_9340);
or U9476 (N_9476,N_9334,N_9344);
nand U9477 (N_9477,N_9387,N_9356);
nor U9478 (N_9478,N_9350,N_9357);
xor U9479 (N_9479,N_9336,N_9375);
nor U9480 (N_9480,N_9349,N_9386);
nand U9481 (N_9481,N_9353,N_9370);
or U9482 (N_9482,N_9344,N_9368);
nand U9483 (N_9483,N_9351,N_9334);
and U9484 (N_9484,N_9384,N_9373);
and U9485 (N_9485,N_9340,N_9387);
or U9486 (N_9486,N_9315,N_9387);
xnor U9487 (N_9487,N_9386,N_9363);
nand U9488 (N_9488,N_9387,N_9397);
and U9489 (N_9489,N_9394,N_9320);
xor U9490 (N_9490,N_9380,N_9315);
nor U9491 (N_9491,N_9359,N_9332);
or U9492 (N_9492,N_9319,N_9307);
xnor U9493 (N_9493,N_9372,N_9370);
and U9494 (N_9494,N_9390,N_9357);
xor U9495 (N_9495,N_9373,N_9374);
nand U9496 (N_9496,N_9390,N_9342);
nor U9497 (N_9497,N_9342,N_9394);
xnor U9498 (N_9498,N_9306,N_9344);
nand U9499 (N_9499,N_9342,N_9367);
nor U9500 (N_9500,N_9456,N_9426);
xor U9501 (N_9501,N_9417,N_9450);
xor U9502 (N_9502,N_9497,N_9428);
or U9503 (N_9503,N_9434,N_9469);
and U9504 (N_9504,N_9453,N_9429);
or U9505 (N_9505,N_9464,N_9423);
and U9506 (N_9506,N_9474,N_9409);
and U9507 (N_9507,N_9479,N_9451);
and U9508 (N_9508,N_9406,N_9407);
nor U9509 (N_9509,N_9472,N_9483);
xor U9510 (N_9510,N_9466,N_9489);
xor U9511 (N_9511,N_9415,N_9444);
or U9512 (N_9512,N_9413,N_9427);
nor U9513 (N_9513,N_9400,N_9460);
nand U9514 (N_9514,N_9403,N_9414);
xor U9515 (N_9515,N_9473,N_9425);
xnor U9516 (N_9516,N_9477,N_9435);
nor U9517 (N_9517,N_9499,N_9441);
xor U9518 (N_9518,N_9438,N_9495);
xor U9519 (N_9519,N_9411,N_9418);
nand U9520 (N_9520,N_9484,N_9454);
and U9521 (N_9521,N_9476,N_9459);
xor U9522 (N_9522,N_9458,N_9452);
nand U9523 (N_9523,N_9449,N_9470);
nand U9524 (N_9524,N_9439,N_9475);
or U9525 (N_9525,N_9487,N_9455);
or U9526 (N_9526,N_9492,N_9433);
nor U9527 (N_9527,N_9457,N_9416);
nor U9528 (N_9528,N_9448,N_9401);
xor U9529 (N_9529,N_9471,N_9462);
nor U9530 (N_9530,N_9486,N_9421);
nand U9531 (N_9531,N_9436,N_9490);
nor U9532 (N_9532,N_9431,N_9422);
or U9533 (N_9533,N_9481,N_9493);
or U9534 (N_9534,N_9430,N_9494);
nor U9535 (N_9535,N_9478,N_9410);
and U9536 (N_9536,N_9461,N_9463);
nor U9537 (N_9537,N_9465,N_9402);
xor U9538 (N_9538,N_9442,N_9424);
nor U9539 (N_9539,N_9496,N_9412);
nand U9540 (N_9540,N_9408,N_9440);
xnor U9541 (N_9541,N_9447,N_9445);
nor U9542 (N_9542,N_9405,N_9480);
xor U9543 (N_9543,N_9485,N_9491);
nand U9544 (N_9544,N_9404,N_9432);
nor U9545 (N_9545,N_9437,N_9420);
nor U9546 (N_9546,N_9467,N_9443);
or U9547 (N_9547,N_9488,N_9419);
nand U9548 (N_9548,N_9482,N_9446);
and U9549 (N_9549,N_9468,N_9498);
and U9550 (N_9550,N_9424,N_9416);
nor U9551 (N_9551,N_9447,N_9411);
and U9552 (N_9552,N_9450,N_9406);
or U9553 (N_9553,N_9499,N_9495);
and U9554 (N_9554,N_9401,N_9478);
xor U9555 (N_9555,N_9458,N_9461);
or U9556 (N_9556,N_9463,N_9417);
xnor U9557 (N_9557,N_9409,N_9486);
and U9558 (N_9558,N_9429,N_9409);
nand U9559 (N_9559,N_9492,N_9429);
and U9560 (N_9560,N_9440,N_9430);
xnor U9561 (N_9561,N_9424,N_9455);
nand U9562 (N_9562,N_9495,N_9450);
or U9563 (N_9563,N_9416,N_9408);
nor U9564 (N_9564,N_9489,N_9497);
and U9565 (N_9565,N_9425,N_9439);
or U9566 (N_9566,N_9448,N_9475);
nand U9567 (N_9567,N_9479,N_9470);
and U9568 (N_9568,N_9487,N_9459);
xnor U9569 (N_9569,N_9423,N_9459);
and U9570 (N_9570,N_9439,N_9468);
nor U9571 (N_9571,N_9412,N_9424);
nor U9572 (N_9572,N_9474,N_9421);
nand U9573 (N_9573,N_9405,N_9404);
and U9574 (N_9574,N_9477,N_9498);
xnor U9575 (N_9575,N_9447,N_9443);
and U9576 (N_9576,N_9434,N_9464);
and U9577 (N_9577,N_9460,N_9483);
or U9578 (N_9578,N_9438,N_9416);
and U9579 (N_9579,N_9434,N_9432);
nor U9580 (N_9580,N_9473,N_9474);
xor U9581 (N_9581,N_9498,N_9430);
and U9582 (N_9582,N_9463,N_9408);
and U9583 (N_9583,N_9408,N_9465);
nand U9584 (N_9584,N_9447,N_9467);
xor U9585 (N_9585,N_9424,N_9463);
or U9586 (N_9586,N_9404,N_9493);
and U9587 (N_9587,N_9449,N_9409);
and U9588 (N_9588,N_9493,N_9412);
and U9589 (N_9589,N_9455,N_9404);
or U9590 (N_9590,N_9482,N_9474);
xor U9591 (N_9591,N_9449,N_9414);
or U9592 (N_9592,N_9468,N_9452);
nand U9593 (N_9593,N_9472,N_9427);
nand U9594 (N_9594,N_9455,N_9401);
nor U9595 (N_9595,N_9470,N_9488);
nand U9596 (N_9596,N_9405,N_9452);
and U9597 (N_9597,N_9492,N_9479);
nand U9598 (N_9598,N_9402,N_9417);
xnor U9599 (N_9599,N_9458,N_9447);
nor U9600 (N_9600,N_9582,N_9511);
nand U9601 (N_9601,N_9514,N_9558);
nor U9602 (N_9602,N_9549,N_9542);
nor U9603 (N_9603,N_9523,N_9596);
nand U9604 (N_9604,N_9528,N_9559);
nor U9605 (N_9605,N_9576,N_9554);
xnor U9606 (N_9606,N_9574,N_9543);
nor U9607 (N_9607,N_9590,N_9525);
and U9608 (N_9608,N_9592,N_9553);
nand U9609 (N_9609,N_9568,N_9598);
or U9610 (N_9610,N_9547,N_9597);
and U9611 (N_9611,N_9524,N_9571);
and U9612 (N_9612,N_9580,N_9503);
and U9613 (N_9613,N_9504,N_9516);
nand U9614 (N_9614,N_9535,N_9569);
or U9615 (N_9615,N_9536,N_9577);
nor U9616 (N_9616,N_9527,N_9564);
xnor U9617 (N_9617,N_9591,N_9501);
nand U9618 (N_9618,N_9588,N_9561);
xnor U9619 (N_9619,N_9586,N_9552);
and U9620 (N_9620,N_9594,N_9565);
and U9621 (N_9621,N_9533,N_9541);
nor U9622 (N_9622,N_9573,N_9539);
xor U9623 (N_9623,N_9507,N_9595);
nor U9624 (N_9624,N_9509,N_9587);
xor U9625 (N_9625,N_9505,N_9515);
or U9626 (N_9626,N_9544,N_9556);
or U9627 (N_9627,N_9517,N_9537);
and U9628 (N_9628,N_9532,N_9585);
xor U9629 (N_9629,N_9545,N_9546);
and U9630 (N_9630,N_9538,N_9551);
nand U9631 (N_9631,N_9584,N_9506);
and U9632 (N_9632,N_9508,N_9510);
nor U9633 (N_9633,N_9502,N_9513);
or U9634 (N_9634,N_9531,N_9560);
nand U9635 (N_9635,N_9581,N_9518);
nor U9636 (N_9636,N_9599,N_9575);
and U9637 (N_9637,N_9579,N_9512);
xnor U9638 (N_9638,N_9540,N_9548);
nor U9639 (N_9639,N_9570,N_9529);
xnor U9640 (N_9640,N_9534,N_9562);
nand U9641 (N_9641,N_9578,N_9567);
and U9642 (N_9642,N_9583,N_9500);
xnor U9643 (N_9643,N_9572,N_9526);
xnor U9644 (N_9644,N_9550,N_9563);
or U9645 (N_9645,N_9589,N_9520);
or U9646 (N_9646,N_9555,N_9522);
or U9647 (N_9647,N_9566,N_9530);
or U9648 (N_9648,N_9593,N_9557);
or U9649 (N_9649,N_9521,N_9519);
or U9650 (N_9650,N_9560,N_9573);
and U9651 (N_9651,N_9573,N_9549);
xnor U9652 (N_9652,N_9593,N_9576);
nand U9653 (N_9653,N_9500,N_9598);
and U9654 (N_9654,N_9535,N_9546);
nor U9655 (N_9655,N_9598,N_9503);
or U9656 (N_9656,N_9523,N_9575);
nand U9657 (N_9657,N_9591,N_9587);
xor U9658 (N_9658,N_9598,N_9591);
and U9659 (N_9659,N_9534,N_9514);
and U9660 (N_9660,N_9509,N_9522);
and U9661 (N_9661,N_9592,N_9573);
nand U9662 (N_9662,N_9557,N_9598);
nor U9663 (N_9663,N_9573,N_9546);
nand U9664 (N_9664,N_9536,N_9590);
xor U9665 (N_9665,N_9561,N_9530);
xnor U9666 (N_9666,N_9512,N_9508);
nand U9667 (N_9667,N_9534,N_9532);
and U9668 (N_9668,N_9580,N_9545);
nand U9669 (N_9669,N_9514,N_9582);
or U9670 (N_9670,N_9513,N_9577);
xor U9671 (N_9671,N_9529,N_9580);
and U9672 (N_9672,N_9572,N_9557);
nand U9673 (N_9673,N_9516,N_9518);
and U9674 (N_9674,N_9522,N_9544);
xor U9675 (N_9675,N_9516,N_9525);
nand U9676 (N_9676,N_9535,N_9506);
and U9677 (N_9677,N_9519,N_9576);
nor U9678 (N_9678,N_9532,N_9560);
and U9679 (N_9679,N_9550,N_9561);
nand U9680 (N_9680,N_9599,N_9591);
nor U9681 (N_9681,N_9552,N_9557);
nand U9682 (N_9682,N_9514,N_9597);
or U9683 (N_9683,N_9569,N_9552);
xor U9684 (N_9684,N_9577,N_9575);
xor U9685 (N_9685,N_9527,N_9507);
and U9686 (N_9686,N_9517,N_9562);
nor U9687 (N_9687,N_9504,N_9585);
nand U9688 (N_9688,N_9525,N_9537);
and U9689 (N_9689,N_9592,N_9539);
and U9690 (N_9690,N_9557,N_9568);
nor U9691 (N_9691,N_9576,N_9550);
nor U9692 (N_9692,N_9569,N_9566);
or U9693 (N_9693,N_9567,N_9576);
and U9694 (N_9694,N_9528,N_9548);
xnor U9695 (N_9695,N_9573,N_9534);
or U9696 (N_9696,N_9540,N_9521);
and U9697 (N_9697,N_9557,N_9589);
and U9698 (N_9698,N_9561,N_9501);
nand U9699 (N_9699,N_9555,N_9510);
or U9700 (N_9700,N_9628,N_9642);
or U9701 (N_9701,N_9681,N_9600);
xor U9702 (N_9702,N_9661,N_9643);
nand U9703 (N_9703,N_9676,N_9696);
nor U9704 (N_9704,N_9607,N_9660);
or U9705 (N_9705,N_9680,N_9608);
nand U9706 (N_9706,N_9666,N_9654);
xor U9707 (N_9707,N_9687,N_9684);
or U9708 (N_9708,N_9617,N_9678);
nor U9709 (N_9709,N_9612,N_9698);
and U9710 (N_9710,N_9640,N_9634);
and U9711 (N_9711,N_9625,N_9663);
and U9712 (N_9712,N_9606,N_9620);
nor U9713 (N_9713,N_9648,N_9615);
nand U9714 (N_9714,N_9621,N_9673);
nor U9715 (N_9715,N_9638,N_9644);
xnor U9716 (N_9716,N_9667,N_9633);
nor U9717 (N_9717,N_9669,N_9675);
and U9718 (N_9718,N_9604,N_9636);
or U9719 (N_9719,N_9647,N_9679);
xnor U9720 (N_9720,N_9602,N_9651);
or U9721 (N_9721,N_9686,N_9627);
and U9722 (N_9722,N_9695,N_9629);
or U9723 (N_9723,N_9671,N_9692);
and U9724 (N_9724,N_9637,N_9685);
and U9725 (N_9725,N_9674,N_9672);
xnor U9726 (N_9726,N_9650,N_9605);
and U9727 (N_9727,N_9641,N_9652);
or U9728 (N_9728,N_9649,N_9631);
or U9729 (N_9729,N_9645,N_9682);
xnor U9730 (N_9730,N_9616,N_9699);
nor U9731 (N_9731,N_9691,N_9653);
and U9732 (N_9732,N_9614,N_9658);
xor U9733 (N_9733,N_9656,N_9618);
or U9734 (N_9734,N_9662,N_9694);
nor U9735 (N_9735,N_9611,N_9630);
or U9736 (N_9736,N_9622,N_9610);
or U9737 (N_9737,N_9623,N_9609);
nand U9738 (N_9738,N_9668,N_9619);
and U9739 (N_9739,N_9689,N_9657);
nand U9740 (N_9740,N_9655,N_9639);
or U9741 (N_9741,N_9601,N_9693);
xor U9742 (N_9742,N_9635,N_9613);
and U9743 (N_9743,N_9664,N_9697);
nor U9744 (N_9744,N_9603,N_9677);
nand U9745 (N_9745,N_9665,N_9683);
nor U9746 (N_9746,N_9670,N_9624);
nand U9747 (N_9747,N_9690,N_9688);
nor U9748 (N_9748,N_9632,N_9646);
and U9749 (N_9749,N_9626,N_9659);
xor U9750 (N_9750,N_9679,N_9655);
nor U9751 (N_9751,N_9620,N_9633);
nor U9752 (N_9752,N_9614,N_9684);
and U9753 (N_9753,N_9630,N_9603);
and U9754 (N_9754,N_9682,N_9632);
and U9755 (N_9755,N_9680,N_9656);
or U9756 (N_9756,N_9624,N_9697);
nor U9757 (N_9757,N_9635,N_9657);
and U9758 (N_9758,N_9655,N_9651);
xor U9759 (N_9759,N_9606,N_9699);
xnor U9760 (N_9760,N_9603,N_9660);
and U9761 (N_9761,N_9687,N_9608);
nor U9762 (N_9762,N_9644,N_9664);
and U9763 (N_9763,N_9639,N_9653);
nand U9764 (N_9764,N_9629,N_9699);
nand U9765 (N_9765,N_9696,N_9684);
and U9766 (N_9766,N_9686,N_9616);
and U9767 (N_9767,N_9672,N_9689);
nor U9768 (N_9768,N_9694,N_9671);
xor U9769 (N_9769,N_9640,N_9693);
nor U9770 (N_9770,N_9647,N_9698);
and U9771 (N_9771,N_9686,N_9617);
and U9772 (N_9772,N_9667,N_9639);
xnor U9773 (N_9773,N_9605,N_9612);
or U9774 (N_9774,N_9629,N_9615);
nand U9775 (N_9775,N_9637,N_9678);
xnor U9776 (N_9776,N_9643,N_9695);
and U9777 (N_9777,N_9698,N_9616);
xnor U9778 (N_9778,N_9656,N_9695);
or U9779 (N_9779,N_9611,N_9608);
nand U9780 (N_9780,N_9687,N_9625);
nand U9781 (N_9781,N_9649,N_9662);
xor U9782 (N_9782,N_9634,N_9695);
or U9783 (N_9783,N_9625,N_9608);
and U9784 (N_9784,N_9667,N_9660);
and U9785 (N_9785,N_9676,N_9678);
and U9786 (N_9786,N_9628,N_9637);
and U9787 (N_9787,N_9662,N_9698);
nand U9788 (N_9788,N_9677,N_9682);
xnor U9789 (N_9789,N_9685,N_9625);
and U9790 (N_9790,N_9662,N_9603);
nor U9791 (N_9791,N_9608,N_9655);
or U9792 (N_9792,N_9620,N_9619);
and U9793 (N_9793,N_9648,N_9661);
nand U9794 (N_9794,N_9631,N_9673);
nand U9795 (N_9795,N_9697,N_9610);
nor U9796 (N_9796,N_9633,N_9641);
and U9797 (N_9797,N_9676,N_9607);
nand U9798 (N_9798,N_9610,N_9625);
nor U9799 (N_9799,N_9624,N_9603);
and U9800 (N_9800,N_9759,N_9741);
and U9801 (N_9801,N_9764,N_9707);
xnor U9802 (N_9802,N_9729,N_9709);
nand U9803 (N_9803,N_9748,N_9785);
nor U9804 (N_9804,N_9706,N_9750);
and U9805 (N_9805,N_9782,N_9711);
and U9806 (N_9806,N_9758,N_9756);
or U9807 (N_9807,N_9797,N_9736);
and U9808 (N_9808,N_9704,N_9788);
nor U9809 (N_9809,N_9715,N_9752);
nand U9810 (N_9810,N_9793,N_9720);
nand U9811 (N_9811,N_9718,N_9733);
nor U9812 (N_9812,N_9738,N_9717);
xnor U9813 (N_9813,N_9784,N_9755);
xor U9814 (N_9814,N_9713,N_9778);
and U9815 (N_9815,N_9701,N_9745);
or U9816 (N_9816,N_9774,N_9771);
and U9817 (N_9817,N_9795,N_9792);
nand U9818 (N_9818,N_9767,N_9772);
xor U9819 (N_9819,N_9735,N_9742);
xor U9820 (N_9820,N_9779,N_9702);
or U9821 (N_9821,N_9716,N_9790);
and U9822 (N_9822,N_9747,N_9773);
and U9823 (N_9823,N_9799,N_9757);
and U9824 (N_9824,N_9719,N_9777);
and U9825 (N_9825,N_9714,N_9769);
nor U9826 (N_9826,N_9765,N_9781);
and U9827 (N_9827,N_9783,N_9740);
and U9828 (N_9828,N_9722,N_9789);
or U9829 (N_9829,N_9700,N_9734);
and U9830 (N_9830,N_9787,N_9739);
and U9831 (N_9831,N_9737,N_9705);
xor U9832 (N_9832,N_9743,N_9766);
and U9833 (N_9833,N_9730,N_9725);
or U9834 (N_9834,N_9763,N_9744);
xnor U9835 (N_9835,N_9794,N_9710);
and U9836 (N_9836,N_9712,N_9727);
xor U9837 (N_9837,N_9732,N_9780);
or U9838 (N_9838,N_9723,N_9761);
nand U9839 (N_9839,N_9775,N_9703);
nor U9840 (N_9840,N_9796,N_9791);
xor U9841 (N_9841,N_9776,N_9786);
nor U9842 (N_9842,N_9762,N_9746);
nand U9843 (N_9843,N_9708,N_9754);
and U9844 (N_9844,N_9760,N_9728);
or U9845 (N_9845,N_9753,N_9770);
xnor U9846 (N_9846,N_9724,N_9726);
and U9847 (N_9847,N_9721,N_9749);
or U9848 (N_9848,N_9731,N_9798);
or U9849 (N_9849,N_9768,N_9751);
xor U9850 (N_9850,N_9769,N_9781);
xnor U9851 (N_9851,N_9793,N_9726);
nor U9852 (N_9852,N_9766,N_9705);
xnor U9853 (N_9853,N_9781,N_9785);
and U9854 (N_9854,N_9759,N_9799);
nor U9855 (N_9855,N_9731,N_9721);
or U9856 (N_9856,N_9709,N_9750);
or U9857 (N_9857,N_9769,N_9721);
nand U9858 (N_9858,N_9725,N_9711);
and U9859 (N_9859,N_9702,N_9747);
and U9860 (N_9860,N_9756,N_9720);
and U9861 (N_9861,N_9723,N_9797);
xor U9862 (N_9862,N_9702,N_9748);
or U9863 (N_9863,N_9736,N_9733);
nor U9864 (N_9864,N_9706,N_9742);
xor U9865 (N_9865,N_9700,N_9763);
nor U9866 (N_9866,N_9765,N_9701);
or U9867 (N_9867,N_9770,N_9734);
or U9868 (N_9868,N_9791,N_9711);
xor U9869 (N_9869,N_9765,N_9782);
nor U9870 (N_9870,N_9794,N_9764);
or U9871 (N_9871,N_9747,N_9778);
nand U9872 (N_9872,N_9703,N_9768);
or U9873 (N_9873,N_9762,N_9744);
xnor U9874 (N_9874,N_9735,N_9788);
nor U9875 (N_9875,N_9722,N_9700);
nor U9876 (N_9876,N_9734,N_9714);
xnor U9877 (N_9877,N_9720,N_9773);
or U9878 (N_9878,N_9796,N_9792);
nor U9879 (N_9879,N_9782,N_9738);
nand U9880 (N_9880,N_9775,N_9787);
or U9881 (N_9881,N_9703,N_9756);
nand U9882 (N_9882,N_9761,N_9789);
nand U9883 (N_9883,N_9733,N_9717);
nor U9884 (N_9884,N_9720,N_9740);
and U9885 (N_9885,N_9707,N_9728);
nor U9886 (N_9886,N_9766,N_9729);
or U9887 (N_9887,N_9745,N_9734);
xnor U9888 (N_9888,N_9777,N_9756);
and U9889 (N_9889,N_9722,N_9787);
xnor U9890 (N_9890,N_9787,N_9726);
nor U9891 (N_9891,N_9710,N_9792);
nand U9892 (N_9892,N_9758,N_9791);
and U9893 (N_9893,N_9728,N_9720);
and U9894 (N_9894,N_9735,N_9757);
nand U9895 (N_9895,N_9750,N_9724);
xor U9896 (N_9896,N_9741,N_9783);
or U9897 (N_9897,N_9745,N_9792);
nor U9898 (N_9898,N_9769,N_9762);
or U9899 (N_9899,N_9753,N_9784);
or U9900 (N_9900,N_9820,N_9854);
and U9901 (N_9901,N_9882,N_9889);
or U9902 (N_9902,N_9830,N_9849);
and U9903 (N_9903,N_9887,N_9856);
xnor U9904 (N_9904,N_9814,N_9801);
nand U9905 (N_9905,N_9817,N_9867);
nand U9906 (N_9906,N_9899,N_9865);
or U9907 (N_9907,N_9855,N_9842);
nand U9908 (N_9908,N_9831,N_9876);
xnor U9909 (N_9909,N_9839,N_9880);
xnor U9910 (N_9910,N_9862,N_9895);
or U9911 (N_9911,N_9828,N_9836);
and U9912 (N_9912,N_9848,N_9809);
nand U9913 (N_9913,N_9838,N_9872);
xor U9914 (N_9914,N_9802,N_9834);
xor U9915 (N_9915,N_9851,N_9835);
and U9916 (N_9916,N_9861,N_9870);
or U9917 (N_9917,N_9868,N_9888);
and U9918 (N_9918,N_9819,N_9890);
xor U9919 (N_9919,N_9881,N_9827);
nand U9920 (N_9920,N_9847,N_9823);
xnor U9921 (N_9921,N_9853,N_9806);
xor U9922 (N_9922,N_9812,N_9808);
nand U9923 (N_9923,N_9800,N_9883);
nand U9924 (N_9924,N_9816,N_9873);
nor U9925 (N_9925,N_9803,N_9884);
or U9926 (N_9926,N_9892,N_9860);
nand U9927 (N_9927,N_9826,N_9822);
and U9928 (N_9928,N_9825,N_9878);
nor U9929 (N_9929,N_9829,N_9858);
xor U9930 (N_9930,N_9843,N_9804);
nand U9931 (N_9931,N_9811,N_9893);
or U9932 (N_9932,N_9894,N_9850);
xnor U9933 (N_9933,N_9898,N_9869);
nor U9934 (N_9934,N_9845,N_9852);
nand U9935 (N_9935,N_9875,N_9813);
nor U9936 (N_9936,N_9885,N_9815);
xnor U9937 (N_9937,N_9821,N_9896);
nand U9938 (N_9938,N_9844,N_9824);
nor U9939 (N_9939,N_9857,N_9863);
nor U9940 (N_9940,N_9891,N_9833);
nor U9941 (N_9941,N_9846,N_9840);
nand U9942 (N_9942,N_9874,N_9841);
and U9943 (N_9943,N_9871,N_9879);
or U9944 (N_9944,N_9837,N_9832);
xor U9945 (N_9945,N_9807,N_9877);
nand U9946 (N_9946,N_9866,N_9886);
nor U9947 (N_9947,N_9864,N_9859);
nand U9948 (N_9948,N_9897,N_9805);
nand U9949 (N_9949,N_9810,N_9818);
and U9950 (N_9950,N_9859,N_9813);
nand U9951 (N_9951,N_9865,N_9843);
nor U9952 (N_9952,N_9819,N_9814);
or U9953 (N_9953,N_9898,N_9863);
xor U9954 (N_9954,N_9812,N_9871);
or U9955 (N_9955,N_9820,N_9894);
or U9956 (N_9956,N_9818,N_9805);
nor U9957 (N_9957,N_9876,N_9865);
or U9958 (N_9958,N_9855,N_9858);
or U9959 (N_9959,N_9823,N_9861);
and U9960 (N_9960,N_9831,N_9832);
nor U9961 (N_9961,N_9810,N_9870);
nor U9962 (N_9962,N_9888,N_9806);
xnor U9963 (N_9963,N_9875,N_9844);
nand U9964 (N_9964,N_9869,N_9857);
xor U9965 (N_9965,N_9803,N_9867);
xnor U9966 (N_9966,N_9834,N_9858);
nor U9967 (N_9967,N_9800,N_9824);
xor U9968 (N_9968,N_9801,N_9848);
xnor U9969 (N_9969,N_9861,N_9802);
and U9970 (N_9970,N_9814,N_9837);
and U9971 (N_9971,N_9846,N_9847);
and U9972 (N_9972,N_9884,N_9852);
or U9973 (N_9973,N_9894,N_9832);
and U9974 (N_9974,N_9892,N_9841);
xnor U9975 (N_9975,N_9890,N_9841);
nor U9976 (N_9976,N_9824,N_9811);
xor U9977 (N_9977,N_9842,N_9810);
nor U9978 (N_9978,N_9820,N_9887);
or U9979 (N_9979,N_9878,N_9897);
nor U9980 (N_9980,N_9808,N_9892);
nor U9981 (N_9981,N_9857,N_9845);
xnor U9982 (N_9982,N_9862,N_9884);
or U9983 (N_9983,N_9862,N_9806);
and U9984 (N_9984,N_9882,N_9868);
or U9985 (N_9985,N_9826,N_9874);
xor U9986 (N_9986,N_9854,N_9877);
or U9987 (N_9987,N_9897,N_9888);
xnor U9988 (N_9988,N_9839,N_9892);
or U9989 (N_9989,N_9848,N_9850);
or U9990 (N_9990,N_9861,N_9884);
xnor U9991 (N_9991,N_9881,N_9875);
and U9992 (N_9992,N_9838,N_9894);
and U9993 (N_9993,N_9844,N_9881);
nor U9994 (N_9994,N_9872,N_9821);
nor U9995 (N_9995,N_9816,N_9844);
nor U9996 (N_9996,N_9845,N_9805);
xnor U9997 (N_9997,N_9835,N_9841);
and U9998 (N_9998,N_9842,N_9836);
or U9999 (N_9999,N_9863,N_9884);
xnor UO_0 (O_0,N_9903,N_9926);
and UO_1 (O_1,N_9948,N_9988);
and UO_2 (O_2,N_9982,N_9915);
or UO_3 (O_3,N_9966,N_9905);
nor UO_4 (O_4,N_9958,N_9963);
xor UO_5 (O_5,N_9999,N_9932);
nand UO_6 (O_6,N_9987,N_9937);
xnor UO_7 (O_7,N_9906,N_9941);
nand UO_8 (O_8,N_9957,N_9985);
or UO_9 (O_9,N_9959,N_9981);
nand UO_10 (O_10,N_9994,N_9935);
nand UO_11 (O_11,N_9919,N_9950);
nand UO_12 (O_12,N_9964,N_9940);
nor UO_13 (O_13,N_9952,N_9992);
nand UO_14 (O_14,N_9996,N_9929);
and UO_15 (O_15,N_9908,N_9990);
nand UO_16 (O_16,N_9942,N_9930);
and UO_17 (O_17,N_9911,N_9924);
and UO_18 (O_18,N_9914,N_9928);
nand UO_19 (O_19,N_9976,N_9910);
xor UO_20 (O_20,N_9989,N_9995);
nand UO_21 (O_21,N_9923,N_9931);
xor UO_22 (O_22,N_9978,N_9962);
or UO_23 (O_23,N_9947,N_9968);
nor UO_24 (O_24,N_9933,N_9974);
nand UO_25 (O_25,N_9961,N_9993);
or UO_26 (O_26,N_9907,N_9983);
and UO_27 (O_27,N_9918,N_9945);
and UO_28 (O_28,N_9922,N_9969);
xnor UO_29 (O_29,N_9913,N_9943);
nand UO_30 (O_30,N_9953,N_9920);
and UO_31 (O_31,N_9944,N_9902);
or UO_32 (O_32,N_9939,N_9917);
and UO_33 (O_33,N_9970,N_9927);
and UO_34 (O_34,N_9904,N_9901);
or UO_35 (O_35,N_9925,N_9977);
and UO_36 (O_36,N_9998,N_9912);
nor UO_37 (O_37,N_9921,N_9971);
nor UO_38 (O_38,N_9938,N_9954);
xnor UO_39 (O_39,N_9991,N_9916);
nand UO_40 (O_40,N_9972,N_9955);
nand UO_41 (O_41,N_9951,N_9986);
and UO_42 (O_42,N_9975,N_9934);
nand UO_43 (O_43,N_9980,N_9909);
and UO_44 (O_44,N_9936,N_9967);
or UO_45 (O_45,N_9956,N_9984);
nand UO_46 (O_46,N_9973,N_9900);
xor UO_47 (O_47,N_9979,N_9946);
or UO_48 (O_48,N_9949,N_9965);
and UO_49 (O_49,N_9997,N_9960);
and UO_50 (O_50,N_9912,N_9910);
nor UO_51 (O_51,N_9953,N_9975);
and UO_52 (O_52,N_9947,N_9979);
xor UO_53 (O_53,N_9958,N_9983);
and UO_54 (O_54,N_9953,N_9930);
nand UO_55 (O_55,N_9910,N_9934);
nor UO_56 (O_56,N_9913,N_9932);
nor UO_57 (O_57,N_9958,N_9913);
and UO_58 (O_58,N_9969,N_9931);
nand UO_59 (O_59,N_9996,N_9944);
xnor UO_60 (O_60,N_9901,N_9956);
xnor UO_61 (O_61,N_9977,N_9979);
and UO_62 (O_62,N_9908,N_9947);
and UO_63 (O_63,N_9958,N_9942);
or UO_64 (O_64,N_9959,N_9979);
nor UO_65 (O_65,N_9976,N_9903);
nor UO_66 (O_66,N_9925,N_9969);
xnor UO_67 (O_67,N_9955,N_9941);
or UO_68 (O_68,N_9943,N_9912);
xnor UO_69 (O_69,N_9962,N_9976);
nand UO_70 (O_70,N_9921,N_9958);
xnor UO_71 (O_71,N_9969,N_9989);
and UO_72 (O_72,N_9912,N_9926);
or UO_73 (O_73,N_9910,N_9974);
xor UO_74 (O_74,N_9932,N_9995);
nor UO_75 (O_75,N_9946,N_9981);
nand UO_76 (O_76,N_9904,N_9929);
and UO_77 (O_77,N_9985,N_9943);
xor UO_78 (O_78,N_9987,N_9998);
nand UO_79 (O_79,N_9922,N_9957);
nor UO_80 (O_80,N_9943,N_9990);
or UO_81 (O_81,N_9912,N_9984);
nand UO_82 (O_82,N_9995,N_9999);
nand UO_83 (O_83,N_9976,N_9938);
or UO_84 (O_84,N_9996,N_9915);
nand UO_85 (O_85,N_9988,N_9951);
and UO_86 (O_86,N_9968,N_9940);
nand UO_87 (O_87,N_9920,N_9999);
xor UO_88 (O_88,N_9908,N_9983);
nand UO_89 (O_89,N_9917,N_9910);
xor UO_90 (O_90,N_9914,N_9979);
nor UO_91 (O_91,N_9916,N_9953);
or UO_92 (O_92,N_9908,N_9944);
or UO_93 (O_93,N_9907,N_9945);
nor UO_94 (O_94,N_9937,N_9933);
xnor UO_95 (O_95,N_9963,N_9912);
nand UO_96 (O_96,N_9934,N_9938);
nor UO_97 (O_97,N_9982,N_9914);
or UO_98 (O_98,N_9983,N_9903);
and UO_99 (O_99,N_9987,N_9957);
nor UO_100 (O_100,N_9909,N_9975);
xor UO_101 (O_101,N_9945,N_9927);
nor UO_102 (O_102,N_9999,N_9994);
nand UO_103 (O_103,N_9952,N_9973);
or UO_104 (O_104,N_9914,N_9961);
and UO_105 (O_105,N_9900,N_9933);
nor UO_106 (O_106,N_9946,N_9974);
nand UO_107 (O_107,N_9987,N_9977);
nor UO_108 (O_108,N_9989,N_9919);
and UO_109 (O_109,N_9970,N_9990);
nor UO_110 (O_110,N_9921,N_9924);
and UO_111 (O_111,N_9987,N_9925);
xor UO_112 (O_112,N_9980,N_9900);
and UO_113 (O_113,N_9926,N_9937);
or UO_114 (O_114,N_9941,N_9945);
or UO_115 (O_115,N_9992,N_9993);
or UO_116 (O_116,N_9904,N_9903);
nor UO_117 (O_117,N_9943,N_9980);
nor UO_118 (O_118,N_9945,N_9975);
nor UO_119 (O_119,N_9958,N_9922);
xnor UO_120 (O_120,N_9986,N_9967);
and UO_121 (O_121,N_9970,N_9969);
nor UO_122 (O_122,N_9918,N_9917);
and UO_123 (O_123,N_9984,N_9955);
or UO_124 (O_124,N_9978,N_9985);
or UO_125 (O_125,N_9928,N_9993);
or UO_126 (O_126,N_9911,N_9900);
or UO_127 (O_127,N_9928,N_9967);
nand UO_128 (O_128,N_9977,N_9910);
nor UO_129 (O_129,N_9955,N_9997);
and UO_130 (O_130,N_9914,N_9900);
xnor UO_131 (O_131,N_9925,N_9918);
or UO_132 (O_132,N_9947,N_9981);
nand UO_133 (O_133,N_9940,N_9920);
xor UO_134 (O_134,N_9903,N_9941);
or UO_135 (O_135,N_9990,N_9947);
xnor UO_136 (O_136,N_9922,N_9918);
nor UO_137 (O_137,N_9912,N_9990);
or UO_138 (O_138,N_9972,N_9942);
nor UO_139 (O_139,N_9971,N_9960);
nand UO_140 (O_140,N_9936,N_9961);
nor UO_141 (O_141,N_9935,N_9950);
nand UO_142 (O_142,N_9935,N_9930);
and UO_143 (O_143,N_9910,N_9951);
nor UO_144 (O_144,N_9921,N_9957);
and UO_145 (O_145,N_9910,N_9954);
nor UO_146 (O_146,N_9978,N_9911);
or UO_147 (O_147,N_9994,N_9914);
or UO_148 (O_148,N_9940,N_9950);
nor UO_149 (O_149,N_9945,N_9989);
and UO_150 (O_150,N_9943,N_9928);
xor UO_151 (O_151,N_9994,N_9916);
xor UO_152 (O_152,N_9925,N_9910);
nand UO_153 (O_153,N_9910,N_9981);
and UO_154 (O_154,N_9921,N_9904);
nor UO_155 (O_155,N_9912,N_9913);
and UO_156 (O_156,N_9974,N_9978);
and UO_157 (O_157,N_9936,N_9981);
and UO_158 (O_158,N_9972,N_9956);
and UO_159 (O_159,N_9907,N_9991);
or UO_160 (O_160,N_9921,N_9951);
nand UO_161 (O_161,N_9915,N_9938);
or UO_162 (O_162,N_9900,N_9921);
xnor UO_163 (O_163,N_9999,N_9981);
or UO_164 (O_164,N_9936,N_9946);
nand UO_165 (O_165,N_9994,N_9925);
or UO_166 (O_166,N_9969,N_9905);
or UO_167 (O_167,N_9941,N_9939);
xor UO_168 (O_168,N_9909,N_9945);
and UO_169 (O_169,N_9910,N_9938);
xor UO_170 (O_170,N_9984,N_9900);
nand UO_171 (O_171,N_9929,N_9973);
and UO_172 (O_172,N_9906,N_9938);
xnor UO_173 (O_173,N_9913,N_9938);
nor UO_174 (O_174,N_9971,N_9976);
and UO_175 (O_175,N_9957,N_9927);
nor UO_176 (O_176,N_9937,N_9917);
or UO_177 (O_177,N_9927,N_9993);
nand UO_178 (O_178,N_9932,N_9966);
nor UO_179 (O_179,N_9959,N_9945);
or UO_180 (O_180,N_9971,N_9991);
nor UO_181 (O_181,N_9922,N_9979);
nor UO_182 (O_182,N_9995,N_9959);
nand UO_183 (O_183,N_9940,N_9980);
or UO_184 (O_184,N_9965,N_9991);
or UO_185 (O_185,N_9953,N_9940);
nand UO_186 (O_186,N_9989,N_9926);
nor UO_187 (O_187,N_9991,N_9950);
nor UO_188 (O_188,N_9997,N_9967);
or UO_189 (O_189,N_9960,N_9985);
nor UO_190 (O_190,N_9950,N_9931);
nand UO_191 (O_191,N_9985,N_9951);
xor UO_192 (O_192,N_9961,N_9944);
nand UO_193 (O_193,N_9930,N_9988);
nor UO_194 (O_194,N_9925,N_9953);
and UO_195 (O_195,N_9911,N_9930);
xor UO_196 (O_196,N_9945,N_9961);
nand UO_197 (O_197,N_9956,N_9946);
nand UO_198 (O_198,N_9938,N_9901);
xor UO_199 (O_199,N_9945,N_9971);
nand UO_200 (O_200,N_9989,N_9981);
and UO_201 (O_201,N_9954,N_9997);
nand UO_202 (O_202,N_9932,N_9942);
xnor UO_203 (O_203,N_9922,N_9925);
and UO_204 (O_204,N_9937,N_9920);
xnor UO_205 (O_205,N_9925,N_9924);
and UO_206 (O_206,N_9978,N_9966);
or UO_207 (O_207,N_9993,N_9931);
or UO_208 (O_208,N_9921,N_9915);
or UO_209 (O_209,N_9993,N_9964);
nand UO_210 (O_210,N_9920,N_9970);
or UO_211 (O_211,N_9946,N_9920);
xor UO_212 (O_212,N_9937,N_9909);
nand UO_213 (O_213,N_9973,N_9935);
nand UO_214 (O_214,N_9985,N_9994);
and UO_215 (O_215,N_9926,N_9962);
and UO_216 (O_216,N_9962,N_9985);
xnor UO_217 (O_217,N_9969,N_9985);
xor UO_218 (O_218,N_9948,N_9955);
nor UO_219 (O_219,N_9929,N_9946);
xor UO_220 (O_220,N_9954,N_9982);
nand UO_221 (O_221,N_9934,N_9997);
nor UO_222 (O_222,N_9951,N_9944);
and UO_223 (O_223,N_9998,N_9949);
or UO_224 (O_224,N_9902,N_9957);
nor UO_225 (O_225,N_9918,N_9940);
xor UO_226 (O_226,N_9945,N_9982);
nand UO_227 (O_227,N_9920,N_9988);
nor UO_228 (O_228,N_9910,N_9933);
and UO_229 (O_229,N_9967,N_9931);
xnor UO_230 (O_230,N_9965,N_9947);
nor UO_231 (O_231,N_9933,N_9954);
nand UO_232 (O_232,N_9972,N_9981);
nor UO_233 (O_233,N_9932,N_9949);
and UO_234 (O_234,N_9951,N_9942);
or UO_235 (O_235,N_9905,N_9959);
and UO_236 (O_236,N_9971,N_9961);
nor UO_237 (O_237,N_9960,N_9925);
xnor UO_238 (O_238,N_9990,N_9989);
nor UO_239 (O_239,N_9968,N_9910);
and UO_240 (O_240,N_9978,N_9991);
xnor UO_241 (O_241,N_9970,N_9936);
nor UO_242 (O_242,N_9918,N_9919);
and UO_243 (O_243,N_9964,N_9984);
or UO_244 (O_244,N_9970,N_9933);
xnor UO_245 (O_245,N_9936,N_9901);
nor UO_246 (O_246,N_9998,N_9948);
nor UO_247 (O_247,N_9910,N_9913);
nor UO_248 (O_248,N_9934,N_9971);
and UO_249 (O_249,N_9932,N_9915);
or UO_250 (O_250,N_9994,N_9921);
and UO_251 (O_251,N_9927,N_9923);
or UO_252 (O_252,N_9992,N_9901);
nor UO_253 (O_253,N_9910,N_9958);
and UO_254 (O_254,N_9956,N_9939);
and UO_255 (O_255,N_9966,N_9934);
nand UO_256 (O_256,N_9928,N_9912);
or UO_257 (O_257,N_9953,N_9904);
nor UO_258 (O_258,N_9974,N_9967);
nand UO_259 (O_259,N_9974,N_9945);
nor UO_260 (O_260,N_9902,N_9971);
xnor UO_261 (O_261,N_9964,N_9999);
xor UO_262 (O_262,N_9946,N_9977);
nor UO_263 (O_263,N_9939,N_9964);
or UO_264 (O_264,N_9942,N_9940);
or UO_265 (O_265,N_9908,N_9971);
or UO_266 (O_266,N_9972,N_9931);
xnor UO_267 (O_267,N_9969,N_9938);
nand UO_268 (O_268,N_9938,N_9950);
nand UO_269 (O_269,N_9914,N_9965);
nand UO_270 (O_270,N_9964,N_9908);
nor UO_271 (O_271,N_9970,N_9917);
and UO_272 (O_272,N_9927,N_9980);
or UO_273 (O_273,N_9972,N_9908);
xnor UO_274 (O_274,N_9959,N_9941);
and UO_275 (O_275,N_9999,N_9998);
nand UO_276 (O_276,N_9907,N_9986);
or UO_277 (O_277,N_9944,N_9905);
or UO_278 (O_278,N_9932,N_9998);
and UO_279 (O_279,N_9952,N_9971);
or UO_280 (O_280,N_9984,N_9949);
nand UO_281 (O_281,N_9972,N_9969);
xor UO_282 (O_282,N_9920,N_9991);
nand UO_283 (O_283,N_9974,N_9905);
xor UO_284 (O_284,N_9928,N_9909);
nor UO_285 (O_285,N_9901,N_9952);
nor UO_286 (O_286,N_9913,N_9988);
or UO_287 (O_287,N_9934,N_9944);
or UO_288 (O_288,N_9944,N_9921);
or UO_289 (O_289,N_9990,N_9928);
nand UO_290 (O_290,N_9980,N_9920);
nor UO_291 (O_291,N_9912,N_9902);
and UO_292 (O_292,N_9986,N_9957);
and UO_293 (O_293,N_9980,N_9977);
nor UO_294 (O_294,N_9917,N_9980);
and UO_295 (O_295,N_9957,N_9990);
nand UO_296 (O_296,N_9940,N_9965);
or UO_297 (O_297,N_9919,N_9988);
and UO_298 (O_298,N_9933,N_9990);
xnor UO_299 (O_299,N_9946,N_9906);
xnor UO_300 (O_300,N_9930,N_9920);
and UO_301 (O_301,N_9961,N_9923);
or UO_302 (O_302,N_9985,N_9968);
nand UO_303 (O_303,N_9926,N_9992);
nand UO_304 (O_304,N_9909,N_9956);
and UO_305 (O_305,N_9954,N_9960);
nand UO_306 (O_306,N_9902,N_9941);
nand UO_307 (O_307,N_9985,N_9923);
nor UO_308 (O_308,N_9900,N_9990);
nand UO_309 (O_309,N_9935,N_9915);
nand UO_310 (O_310,N_9992,N_9983);
or UO_311 (O_311,N_9905,N_9963);
nand UO_312 (O_312,N_9972,N_9996);
nor UO_313 (O_313,N_9990,N_9902);
or UO_314 (O_314,N_9949,N_9907);
nor UO_315 (O_315,N_9930,N_9934);
nor UO_316 (O_316,N_9924,N_9978);
nand UO_317 (O_317,N_9956,N_9917);
nand UO_318 (O_318,N_9984,N_9981);
nor UO_319 (O_319,N_9915,N_9901);
and UO_320 (O_320,N_9930,N_9980);
nor UO_321 (O_321,N_9902,N_9938);
or UO_322 (O_322,N_9939,N_9993);
or UO_323 (O_323,N_9973,N_9907);
and UO_324 (O_324,N_9944,N_9950);
nand UO_325 (O_325,N_9942,N_9983);
nand UO_326 (O_326,N_9916,N_9949);
nand UO_327 (O_327,N_9925,N_9920);
or UO_328 (O_328,N_9913,N_9982);
nor UO_329 (O_329,N_9935,N_9947);
or UO_330 (O_330,N_9939,N_9982);
nor UO_331 (O_331,N_9946,N_9944);
and UO_332 (O_332,N_9916,N_9921);
nand UO_333 (O_333,N_9951,N_9938);
xor UO_334 (O_334,N_9967,N_9906);
or UO_335 (O_335,N_9940,N_9984);
and UO_336 (O_336,N_9927,N_9971);
nor UO_337 (O_337,N_9925,N_9975);
and UO_338 (O_338,N_9989,N_9975);
xnor UO_339 (O_339,N_9997,N_9959);
and UO_340 (O_340,N_9933,N_9999);
xnor UO_341 (O_341,N_9990,N_9996);
nor UO_342 (O_342,N_9936,N_9919);
nor UO_343 (O_343,N_9984,N_9939);
xor UO_344 (O_344,N_9973,N_9970);
and UO_345 (O_345,N_9953,N_9935);
or UO_346 (O_346,N_9924,N_9975);
nand UO_347 (O_347,N_9969,N_9933);
nor UO_348 (O_348,N_9988,N_9973);
nand UO_349 (O_349,N_9958,N_9924);
nand UO_350 (O_350,N_9909,N_9935);
nor UO_351 (O_351,N_9908,N_9979);
xnor UO_352 (O_352,N_9911,N_9945);
nand UO_353 (O_353,N_9943,N_9907);
or UO_354 (O_354,N_9962,N_9968);
nand UO_355 (O_355,N_9980,N_9955);
or UO_356 (O_356,N_9900,N_9947);
and UO_357 (O_357,N_9949,N_9995);
nand UO_358 (O_358,N_9930,N_9976);
nor UO_359 (O_359,N_9960,N_9946);
nor UO_360 (O_360,N_9959,N_9978);
nor UO_361 (O_361,N_9942,N_9905);
xnor UO_362 (O_362,N_9992,N_9985);
and UO_363 (O_363,N_9931,N_9994);
xnor UO_364 (O_364,N_9998,N_9968);
nand UO_365 (O_365,N_9925,N_9911);
nor UO_366 (O_366,N_9916,N_9965);
nand UO_367 (O_367,N_9967,N_9919);
nor UO_368 (O_368,N_9989,N_9904);
nor UO_369 (O_369,N_9972,N_9960);
nand UO_370 (O_370,N_9966,N_9926);
nor UO_371 (O_371,N_9969,N_9956);
and UO_372 (O_372,N_9974,N_9952);
and UO_373 (O_373,N_9967,N_9957);
or UO_374 (O_374,N_9933,N_9961);
nor UO_375 (O_375,N_9924,N_9939);
xor UO_376 (O_376,N_9949,N_9904);
nor UO_377 (O_377,N_9940,N_9944);
or UO_378 (O_378,N_9944,N_9988);
nor UO_379 (O_379,N_9939,N_9905);
nor UO_380 (O_380,N_9915,N_9972);
and UO_381 (O_381,N_9982,N_9902);
nand UO_382 (O_382,N_9911,N_9990);
nand UO_383 (O_383,N_9950,N_9951);
or UO_384 (O_384,N_9979,N_9952);
nand UO_385 (O_385,N_9911,N_9947);
nand UO_386 (O_386,N_9952,N_9966);
xnor UO_387 (O_387,N_9902,N_9999);
or UO_388 (O_388,N_9989,N_9930);
nor UO_389 (O_389,N_9963,N_9931);
nand UO_390 (O_390,N_9984,N_9945);
or UO_391 (O_391,N_9959,N_9940);
or UO_392 (O_392,N_9971,N_9956);
or UO_393 (O_393,N_9986,N_9964);
or UO_394 (O_394,N_9967,N_9933);
nor UO_395 (O_395,N_9945,N_9913);
nand UO_396 (O_396,N_9907,N_9939);
xor UO_397 (O_397,N_9911,N_9984);
nand UO_398 (O_398,N_9914,N_9971);
xor UO_399 (O_399,N_9916,N_9913);
nor UO_400 (O_400,N_9916,N_9967);
xnor UO_401 (O_401,N_9975,N_9903);
xor UO_402 (O_402,N_9962,N_9992);
xor UO_403 (O_403,N_9971,N_9946);
nor UO_404 (O_404,N_9947,N_9999);
nand UO_405 (O_405,N_9993,N_9953);
and UO_406 (O_406,N_9912,N_9970);
xor UO_407 (O_407,N_9944,N_9928);
and UO_408 (O_408,N_9953,N_9913);
and UO_409 (O_409,N_9915,N_9904);
and UO_410 (O_410,N_9929,N_9928);
and UO_411 (O_411,N_9969,N_9919);
or UO_412 (O_412,N_9984,N_9919);
xor UO_413 (O_413,N_9993,N_9965);
nand UO_414 (O_414,N_9920,N_9948);
and UO_415 (O_415,N_9996,N_9907);
or UO_416 (O_416,N_9979,N_9981);
nand UO_417 (O_417,N_9987,N_9960);
and UO_418 (O_418,N_9982,N_9905);
nand UO_419 (O_419,N_9906,N_9939);
or UO_420 (O_420,N_9939,N_9902);
and UO_421 (O_421,N_9952,N_9968);
nor UO_422 (O_422,N_9924,N_9988);
or UO_423 (O_423,N_9992,N_9903);
and UO_424 (O_424,N_9992,N_9991);
xor UO_425 (O_425,N_9999,N_9984);
nand UO_426 (O_426,N_9924,N_9906);
nor UO_427 (O_427,N_9935,N_9966);
nor UO_428 (O_428,N_9943,N_9948);
or UO_429 (O_429,N_9943,N_9977);
nand UO_430 (O_430,N_9927,N_9989);
or UO_431 (O_431,N_9994,N_9923);
or UO_432 (O_432,N_9952,N_9955);
and UO_433 (O_433,N_9991,N_9903);
or UO_434 (O_434,N_9987,N_9969);
nand UO_435 (O_435,N_9905,N_9920);
nor UO_436 (O_436,N_9922,N_9977);
or UO_437 (O_437,N_9959,N_9984);
and UO_438 (O_438,N_9907,N_9994);
and UO_439 (O_439,N_9955,N_9906);
nor UO_440 (O_440,N_9937,N_9914);
nand UO_441 (O_441,N_9981,N_9941);
nand UO_442 (O_442,N_9953,N_9964);
nor UO_443 (O_443,N_9932,N_9990);
nor UO_444 (O_444,N_9922,N_9917);
nor UO_445 (O_445,N_9985,N_9945);
nand UO_446 (O_446,N_9964,N_9982);
or UO_447 (O_447,N_9933,N_9925);
xnor UO_448 (O_448,N_9982,N_9933);
nand UO_449 (O_449,N_9932,N_9982);
xor UO_450 (O_450,N_9996,N_9964);
or UO_451 (O_451,N_9969,N_9975);
or UO_452 (O_452,N_9978,N_9947);
xnor UO_453 (O_453,N_9968,N_9964);
and UO_454 (O_454,N_9955,N_9959);
nand UO_455 (O_455,N_9918,N_9974);
xnor UO_456 (O_456,N_9976,N_9974);
and UO_457 (O_457,N_9962,N_9974);
nor UO_458 (O_458,N_9965,N_9977);
and UO_459 (O_459,N_9992,N_9904);
xor UO_460 (O_460,N_9932,N_9921);
or UO_461 (O_461,N_9913,N_9991);
and UO_462 (O_462,N_9923,N_9954);
xnor UO_463 (O_463,N_9979,N_9957);
nor UO_464 (O_464,N_9966,N_9913);
nand UO_465 (O_465,N_9910,N_9994);
xnor UO_466 (O_466,N_9988,N_9950);
and UO_467 (O_467,N_9919,N_9968);
nor UO_468 (O_468,N_9918,N_9976);
xnor UO_469 (O_469,N_9967,N_9972);
nand UO_470 (O_470,N_9946,N_9951);
nand UO_471 (O_471,N_9924,N_9969);
nor UO_472 (O_472,N_9906,N_9988);
and UO_473 (O_473,N_9930,N_9912);
nand UO_474 (O_474,N_9946,N_9904);
xnor UO_475 (O_475,N_9972,N_9946);
or UO_476 (O_476,N_9979,N_9963);
nor UO_477 (O_477,N_9900,N_9904);
and UO_478 (O_478,N_9944,N_9987);
xor UO_479 (O_479,N_9962,N_9923);
and UO_480 (O_480,N_9952,N_9964);
xor UO_481 (O_481,N_9966,N_9909);
and UO_482 (O_482,N_9972,N_9948);
nor UO_483 (O_483,N_9991,N_9969);
or UO_484 (O_484,N_9986,N_9993);
and UO_485 (O_485,N_9976,N_9906);
nor UO_486 (O_486,N_9963,N_9984);
and UO_487 (O_487,N_9945,N_9994);
xor UO_488 (O_488,N_9917,N_9945);
nand UO_489 (O_489,N_9986,N_9997);
and UO_490 (O_490,N_9949,N_9996);
nand UO_491 (O_491,N_9976,N_9965);
xor UO_492 (O_492,N_9992,N_9988);
xor UO_493 (O_493,N_9931,N_9986);
and UO_494 (O_494,N_9938,N_9917);
xnor UO_495 (O_495,N_9962,N_9979);
nor UO_496 (O_496,N_9960,N_9921);
and UO_497 (O_497,N_9988,N_9908);
nand UO_498 (O_498,N_9947,N_9986);
and UO_499 (O_499,N_9975,N_9984);
xnor UO_500 (O_500,N_9982,N_9944);
xor UO_501 (O_501,N_9965,N_9909);
and UO_502 (O_502,N_9975,N_9943);
nor UO_503 (O_503,N_9917,N_9997);
or UO_504 (O_504,N_9953,N_9989);
xnor UO_505 (O_505,N_9960,N_9907);
nor UO_506 (O_506,N_9929,N_9951);
or UO_507 (O_507,N_9984,N_9989);
and UO_508 (O_508,N_9900,N_9943);
nor UO_509 (O_509,N_9945,N_9929);
and UO_510 (O_510,N_9996,N_9958);
nor UO_511 (O_511,N_9968,N_9915);
nor UO_512 (O_512,N_9968,N_9984);
and UO_513 (O_513,N_9956,N_9914);
nor UO_514 (O_514,N_9971,N_9953);
and UO_515 (O_515,N_9918,N_9943);
nor UO_516 (O_516,N_9967,N_9930);
or UO_517 (O_517,N_9993,N_9925);
nand UO_518 (O_518,N_9963,N_9951);
nand UO_519 (O_519,N_9950,N_9928);
and UO_520 (O_520,N_9969,N_9901);
nand UO_521 (O_521,N_9927,N_9931);
or UO_522 (O_522,N_9956,N_9996);
xnor UO_523 (O_523,N_9984,N_9901);
nand UO_524 (O_524,N_9956,N_9903);
or UO_525 (O_525,N_9984,N_9922);
or UO_526 (O_526,N_9966,N_9971);
or UO_527 (O_527,N_9975,N_9957);
or UO_528 (O_528,N_9900,N_9910);
nand UO_529 (O_529,N_9931,N_9914);
nand UO_530 (O_530,N_9963,N_9921);
nand UO_531 (O_531,N_9938,N_9991);
nor UO_532 (O_532,N_9924,N_9955);
nand UO_533 (O_533,N_9940,N_9989);
xor UO_534 (O_534,N_9998,N_9995);
or UO_535 (O_535,N_9989,N_9928);
and UO_536 (O_536,N_9991,N_9931);
or UO_537 (O_537,N_9983,N_9916);
xnor UO_538 (O_538,N_9926,N_9957);
nand UO_539 (O_539,N_9946,N_9965);
and UO_540 (O_540,N_9998,N_9906);
nand UO_541 (O_541,N_9976,N_9908);
nor UO_542 (O_542,N_9929,N_9947);
nand UO_543 (O_543,N_9999,N_9931);
xnor UO_544 (O_544,N_9977,N_9950);
xnor UO_545 (O_545,N_9966,N_9998);
and UO_546 (O_546,N_9971,N_9916);
or UO_547 (O_547,N_9985,N_9980);
nor UO_548 (O_548,N_9953,N_9906);
nor UO_549 (O_549,N_9904,N_9969);
or UO_550 (O_550,N_9952,N_9940);
xnor UO_551 (O_551,N_9961,N_9918);
xnor UO_552 (O_552,N_9933,N_9909);
and UO_553 (O_553,N_9915,N_9992);
or UO_554 (O_554,N_9944,N_9964);
nand UO_555 (O_555,N_9979,N_9907);
and UO_556 (O_556,N_9993,N_9942);
and UO_557 (O_557,N_9952,N_9980);
and UO_558 (O_558,N_9979,N_9915);
xor UO_559 (O_559,N_9964,N_9948);
nor UO_560 (O_560,N_9920,N_9938);
nand UO_561 (O_561,N_9942,N_9944);
or UO_562 (O_562,N_9992,N_9998);
and UO_563 (O_563,N_9935,N_9914);
xor UO_564 (O_564,N_9946,N_9964);
nand UO_565 (O_565,N_9931,N_9906);
nand UO_566 (O_566,N_9998,N_9971);
nand UO_567 (O_567,N_9949,N_9973);
or UO_568 (O_568,N_9907,N_9909);
xnor UO_569 (O_569,N_9963,N_9960);
or UO_570 (O_570,N_9976,N_9915);
and UO_571 (O_571,N_9934,N_9906);
nor UO_572 (O_572,N_9985,N_9914);
xor UO_573 (O_573,N_9918,N_9932);
and UO_574 (O_574,N_9918,N_9981);
or UO_575 (O_575,N_9945,N_9938);
and UO_576 (O_576,N_9913,N_9906);
and UO_577 (O_577,N_9986,N_9971);
nor UO_578 (O_578,N_9947,N_9904);
nor UO_579 (O_579,N_9965,N_9989);
xnor UO_580 (O_580,N_9983,N_9981);
or UO_581 (O_581,N_9930,N_9960);
or UO_582 (O_582,N_9928,N_9971);
and UO_583 (O_583,N_9938,N_9995);
nand UO_584 (O_584,N_9902,N_9916);
nand UO_585 (O_585,N_9992,N_9920);
and UO_586 (O_586,N_9955,N_9925);
and UO_587 (O_587,N_9938,N_9970);
xnor UO_588 (O_588,N_9902,N_9952);
nand UO_589 (O_589,N_9960,N_9966);
or UO_590 (O_590,N_9997,N_9969);
and UO_591 (O_591,N_9955,N_9939);
or UO_592 (O_592,N_9923,N_9973);
or UO_593 (O_593,N_9990,N_9917);
or UO_594 (O_594,N_9966,N_9941);
xnor UO_595 (O_595,N_9950,N_9969);
xnor UO_596 (O_596,N_9985,N_9932);
or UO_597 (O_597,N_9915,N_9940);
and UO_598 (O_598,N_9909,N_9923);
and UO_599 (O_599,N_9989,N_9960);
nand UO_600 (O_600,N_9937,N_9932);
xnor UO_601 (O_601,N_9902,N_9917);
nand UO_602 (O_602,N_9940,N_9926);
nand UO_603 (O_603,N_9901,N_9932);
and UO_604 (O_604,N_9938,N_9962);
nor UO_605 (O_605,N_9944,N_9907);
xor UO_606 (O_606,N_9979,N_9910);
and UO_607 (O_607,N_9961,N_9952);
or UO_608 (O_608,N_9940,N_9976);
or UO_609 (O_609,N_9932,N_9908);
xor UO_610 (O_610,N_9901,N_9980);
or UO_611 (O_611,N_9905,N_9999);
nor UO_612 (O_612,N_9917,N_9906);
or UO_613 (O_613,N_9922,N_9952);
and UO_614 (O_614,N_9929,N_9988);
nand UO_615 (O_615,N_9925,N_9988);
nand UO_616 (O_616,N_9933,N_9927);
and UO_617 (O_617,N_9987,N_9912);
xor UO_618 (O_618,N_9977,N_9901);
nand UO_619 (O_619,N_9981,N_9970);
and UO_620 (O_620,N_9958,N_9915);
or UO_621 (O_621,N_9954,N_9922);
or UO_622 (O_622,N_9925,N_9981);
xnor UO_623 (O_623,N_9988,N_9954);
nor UO_624 (O_624,N_9980,N_9981);
nand UO_625 (O_625,N_9982,N_9984);
or UO_626 (O_626,N_9906,N_9979);
nand UO_627 (O_627,N_9995,N_9903);
nand UO_628 (O_628,N_9917,N_9908);
and UO_629 (O_629,N_9907,N_9936);
nand UO_630 (O_630,N_9964,N_9905);
or UO_631 (O_631,N_9906,N_9989);
nand UO_632 (O_632,N_9980,N_9910);
nor UO_633 (O_633,N_9940,N_9943);
xor UO_634 (O_634,N_9972,N_9989);
xnor UO_635 (O_635,N_9903,N_9945);
and UO_636 (O_636,N_9907,N_9923);
nor UO_637 (O_637,N_9929,N_9983);
nor UO_638 (O_638,N_9983,N_9940);
and UO_639 (O_639,N_9998,N_9974);
or UO_640 (O_640,N_9927,N_9916);
and UO_641 (O_641,N_9986,N_9905);
nand UO_642 (O_642,N_9907,N_9989);
xor UO_643 (O_643,N_9906,N_9950);
nand UO_644 (O_644,N_9968,N_9976);
or UO_645 (O_645,N_9994,N_9977);
xnor UO_646 (O_646,N_9964,N_9991);
xnor UO_647 (O_647,N_9970,N_9987);
or UO_648 (O_648,N_9955,N_9914);
or UO_649 (O_649,N_9975,N_9902);
or UO_650 (O_650,N_9971,N_9904);
xor UO_651 (O_651,N_9974,N_9980);
nand UO_652 (O_652,N_9964,N_9966);
xor UO_653 (O_653,N_9976,N_9941);
nor UO_654 (O_654,N_9939,N_9962);
xnor UO_655 (O_655,N_9916,N_9918);
nand UO_656 (O_656,N_9986,N_9995);
or UO_657 (O_657,N_9901,N_9931);
and UO_658 (O_658,N_9936,N_9988);
or UO_659 (O_659,N_9972,N_9923);
xnor UO_660 (O_660,N_9964,N_9931);
nor UO_661 (O_661,N_9930,N_9929);
nand UO_662 (O_662,N_9959,N_9964);
nor UO_663 (O_663,N_9988,N_9963);
nand UO_664 (O_664,N_9910,N_9926);
xnor UO_665 (O_665,N_9908,N_9977);
or UO_666 (O_666,N_9941,N_9924);
xnor UO_667 (O_667,N_9979,N_9958);
and UO_668 (O_668,N_9996,N_9981);
and UO_669 (O_669,N_9927,N_9956);
nand UO_670 (O_670,N_9931,N_9996);
nand UO_671 (O_671,N_9936,N_9913);
nand UO_672 (O_672,N_9997,N_9925);
nand UO_673 (O_673,N_9970,N_9955);
nor UO_674 (O_674,N_9963,N_9900);
nor UO_675 (O_675,N_9990,N_9968);
or UO_676 (O_676,N_9961,N_9940);
and UO_677 (O_677,N_9942,N_9946);
or UO_678 (O_678,N_9948,N_9926);
nand UO_679 (O_679,N_9900,N_9962);
nand UO_680 (O_680,N_9929,N_9998);
and UO_681 (O_681,N_9909,N_9924);
and UO_682 (O_682,N_9941,N_9992);
or UO_683 (O_683,N_9929,N_9957);
and UO_684 (O_684,N_9911,N_9929);
and UO_685 (O_685,N_9979,N_9938);
and UO_686 (O_686,N_9932,N_9943);
or UO_687 (O_687,N_9982,N_9903);
nor UO_688 (O_688,N_9978,N_9960);
xor UO_689 (O_689,N_9963,N_9909);
xor UO_690 (O_690,N_9989,N_9901);
nand UO_691 (O_691,N_9938,N_9952);
nand UO_692 (O_692,N_9986,N_9980);
xor UO_693 (O_693,N_9925,N_9978);
nand UO_694 (O_694,N_9944,N_9970);
nand UO_695 (O_695,N_9965,N_9941);
and UO_696 (O_696,N_9915,N_9957);
and UO_697 (O_697,N_9946,N_9913);
and UO_698 (O_698,N_9969,N_9916);
xnor UO_699 (O_699,N_9903,N_9943);
nand UO_700 (O_700,N_9991,N_9944);
and UO_701 (O_701,N_9950,N_9964);
nand UO_702 (O_702,N_9965,N_9918);
nor UO_703 (O_703,N_9978,N_9912);
nor UO_704 (O_704,N_9945,N_9921);
and UO_705 (O_705,N_9911,N_9999);
or UO_706 (O_706,N_9923,N_9903);
or UO_707 (O_707,N_9905,N_9921);
and UO_708 (O_708,N_9952,N_9918);
or UO_709 (O_709,N_9999,N_9924);
xor UO_710 (O_710,N_9986,N_9989);
or UO_711 (O_711,N_9912,N_9985);
xnor UO_712 (O_712,N_9936,N_9900);
xor UO_713 (O_713,N_9978,N_9936);
or UO_714 (O_714,N_9977,N_9920);
xnor UO_715 (O_715,N_9958,N_9931);
xnor UO_716 (O_716,N_9951,N_9924);
nand UO_717 (O_717,N_9909,N_9950);
and UO_718 (O_718,N_9902,N_9908);
nor UO_719 (O_719,N_9931,N_9909);
nor UO_720 (O_720,N_9930,N_9919);
nand UO_721 (O_721,N_9941,N_9988);
and UO_722 (O_722,N_9963,N_9991);
and UO_723 (O_723,N_9947,N_9966);
and UO_724 (O_724,N_9985,N_9996);
nand UO_725 (O_725,N_9944,N_9900);
nand UO_726 (O_726,N_9943,N_9992);
xnor UO_727 (O_727,N_9963,N_9999);
or UO_728 (O_728,N_9909,N_9948);
and UO_729 (O_729,N_9941,N_9915);
or UO_730 (O_730,N_9999,N_9977);
nand UO_731 (O_731,N_9918,N_9987);
nand UO_732 (O_732,N_9977,N_9924);
and UO_733 (O_733,N_9921,N_9977);
or UO_734 (O_734,N_9948,N_9960);
xor UO_735 (O_735,N_9974,N_9995);
and UO_736 (O_736,N_9925,N_9945);
nor UO_737 (O_737,N_9968,N_9981);
xnor UO_738 (O_738,N_9946,N_9985);
or UO_739 (O_739,N_9903,N_9910);
and UO_740 (O_740,N_9965,N_9930);
nand UO_741 (O_741,N_9965,N_9944);
xor UO_742 (O_742,N_9933,N_9947);
nand UO_743 (O_743,N_9970,N_9991);
or UO_744 (O_744,N_9947,N_9943);
nor UO_745 (O_745,N_9960,N_9915);
and UO_746 (O_746,N_9905,N_9951);
xnor UO_747 (O_747,N_9959,N_9966);
nor UO_748 (O_748,N_9978,N_9926);
nand UO_749 (O_749,N_9993,N_9938);
and UO_750 (O_750,N_9902,N_9972);
and UO_751 (O_751,N_9997,N_9950);
or UO_752 (O_752,N_9956,N_9962);
nand UO_753 (O_753,N_9918,N_9930);
and UO_754 (O_754,N_9978,N_9976);
nor UO_755 (O_755,N_9987,N_9986);
or UO_756 (O_756,N_9939,N_9958);
nand UO_757 (O_757,N_9925,N_9938);
nor UO_758 (O_758,N_9953,N_9938);
nand UO_759 (O_759,N_9903,N_9929);
or UO_760 (O_760,N_9970,N_9965);
or UO_761 (O_761,N_9995,N_9934);
nand UO_762 (O_762,N_9943,N_9981);
and UO_763 (O_763,N_9914,N_9923);
and UO_764 (O_764,N_9938,N_9971);
xnor UO_765 (O_765,N_9949,N_9909);
and UO_766 (O_766,N_9900,N_9912);
nand UO_767 (O_767,N_9958,N_9902);
xor UO_768 (O_768,N_9918,N_9912);
nand UO_769 (O_769,N_9991,N_9975);
nand UO_770 (O_770,N_9988,N_9905);
nand UO_771 (O_771,N_9986,N_9991);
nor UO_772 (O_772,N_9927,N_9951);
nor UO_773 (O_773,N_9916,N_9950);
nor UO_774 (O_774,N_9911,N_9981);
nand UO_775 (O_775,N_9900,N_9923);
nor UO_776 (O_776,N_9967,N_9945);
xor UO_777 (O_777,N_9904,N_9960);
nor UO_778 (O_778,N_9941,N_9949);
nor UO_779 (O_779,N_9930,N_9907);
nor UO_780 (O_780,N_9921,N_9911);
nor UO_781 (O_781,N_9948,N_9989);
or UO_782 (O_782,N_9994,N_9902);
nand UO_783 (O_783,N_9921,N_9939);
or UO_784 (O_784,N_9912,N_9923);
nor UO_785 (O_785,N_9992,N_9990);
nand UO_786 (O_786,N_9937,N_9955);
nand UO_787 (O_787,N_9991,N_9919);
xnor UO_788 (O_788,N_9921,N_9946);
xnor UO_789 (O_789,N_9923,N_9939);
and UO_790 (O_790,N_9979,N_9934);
nand UO_791 (O_791,N_9964,N_9995);
or UO_792 (O_792,N_9943,N_9915);
xnor UO_793 (O_793,N_9980,N_9956);
or UO_794 (O_794,N_9940,N_9988);
and UO_795 (O_795,N_9942,N_9999);
and UO_796 (O_796,N_9984,N_9910);
xnor UO_797 (O_797,N_9955,N_9933);
nand UO_798 (O_798,N_9907,N_9931);
nor UO_799 (O_799,N_9929,N_9940);
and UO_800 (O_800,N_9904,N_9961);
nand UO_801 (O_801,N_9991,N_9921);
xnor UO_802 (O_802,N_9900,N_9915);
or UO_803 (O_803,N_9923,N_9935);
and UO_804 (O_804,N_9992,N_9959);
nand UO_805 (O_805,N_9923,N_9942);
nand UO_806 (O_806,N_9904,N_9999);
xor UO_807 (O_807,N_9977,N_9917);
nor UO_808 (O_808,N_9906,N_9900);
nor UO_809 (O_809,N_9994,N_9912);
and UO_810 (O_810,N_9965,N_9982);
nand UO_811 (O_811,N_9967,N_9982);
nor UO_812 (O_812,N_9910,N_9924);
nand UO_813 (O_813,N_9951,N_9965);
or UO_814 (O_814,N_9934,N_9987);
and UO_815 (O_815,N_9949,N_9951);
xor UO_816 (O_816,N_9905,N_9949);
xor UO_817 (O_817,N_9902,N_9978);
nand UO_818 (O_818,N_9937,N_9947);
nand UO_819 (O_819,N_9907,N_9948);
nor UO_820 (O_820,N_9905,N_9973);
and UO_821 (O_821,N_9965,N_9966);
or UO_822 (O_822,N_9944,N_9968);
or UO_823 (O_823,N_9923,N_9925);
nand UO_824 (O_824,N_9937,N_9940);
nor UO_825 (O_825,N_9950,N_9960);
nand UO_826 (O_826,N_9958,N_9992);
or UO_827 (O_827,N_9938,N_9965);
nand UO_828 (O_828,N_9923,N_9992);
nor UO_829 (O_829,N_9979,N_9901);
or UO_830 (O_830,N_9967,N_9990);
nand UO_831 (O_831,N_9992,N_9939);
or UO_832 (O_832,N_9902,N_9913);
nor UO_833 (O_833,N_9986,N_9946);
or UO_834 (O_834,N_9942,N_9990);
xnor UO_835 (O_835,N_9937,N_9974);
xor UO_836 (O_836,N_9982,N_9998);
and UO_837 (O_837,N_9942,N_9994);
nor UO_838 (O_838,N_9940,N_9966);
or UO_839 (O_839,N_9946,N_9937);
nand UO_840 (O_840,N_9924,N_9997);
and UO_841 (O_841,N_9901,N_9981);
and UO_842 (O_842,N_9906,N_9973);
nand UO_843 (O_843,N_9926,N_9932);
nand UO_844 (O_844,N_9988,N_9927);
nand UO_845 (O_845,N_9995,N_9978);
xnor UO_846 (O_846,N_9999,N_9908);
xnor UO_847 (O_847,N_9952,N_9995);
nand UO_848 (O_848,N_9949,N_9993);
or UO_849 (O_849,N_9961,N_9967);
xnor UO_850 (O_850,N_9969,N_9996);
nand UO_851 (O_851,N_9945,N_9928);
or UO_852 (O_852,N_9937,N_9942);
xnor UO_853 (O_853,N_9921,N_9933);
or UO_854 (O_854,N_9908,N_9916);
or UO_855 (O_855,N_9984,N_9996);
xor UO_856 (O_856,N_9965,N_9979);
and UO_857 (O_857,N_9967,N_9988);
nor UO_858 (O_858,N_9983,N_9900);
nor UO_859 (O_859,N_9922,N_9945);
xor UO_860 (O_860,N_9955,N_9950);
xnor UO_861 (O_861,N_9914,N_9969);
nand UO_862 (O_862,N_9984,N_9972);
nor UO_863 (O_863,N_9937,N_9973);
nor UO_864 (O_864,N_9927,N_9964);
xor UO_865 (O_865,N_9993,N_9935);
nand UO_866 (O_866,N_9992,N_9961);
nand UO_867 (O_867,N_9998,N_9935);
nand UO_868 (O_868,N_9914,N_9960);
nand UO_869 (O_869,N_9903,N_9902);
and UO_870 (O_870,N_9914,N_9997);
and UO_871 (O_871,N_9946,N_9900);
nand UO_872 (O_872,N_9982,N_9958);
xor UO_873 (O_873,N_9961,N_9951);
nor UO_874 (O_874,N_9980,N_9944);
xnor UO_875 (O_875,N_9929,N_9920);
and UO_876 (O_876,N_9932,N_9930);
or UO_877 (O_877,N_9967,N_9968);
nor UO_878 (O_878,N_9931,N_9928);
and UO_879 (O_879,N_9975,N_9994);
nor UO_880 (O_880,N_9949,N_9983);
nand UO_881 (O_881,N_9903,N_9907);
or UO_882 (O_882,N_9901,N_9909);
xor UO_883 (O_883,N_9921,N_9903);
nand UO_884 (O_884,N_9926,N_9930);
xor UO_885 (O_885,N_9972,N_9990);
and UO_886 (O_886,N_9925,N_9976);
and UO_887 (O_887,N_9936,N_9968);
nand UO_888 (O_888,N_9936,N_9930);
nand UO_889 (O_889,N_9983,N_9915);
xnor UO_890 (O_890,N_9974,N_9916);
and UO_891 (O_891,N_9988,N_9960);
and UO_892 (O_892,N_9995,N_9922);
nor UO_893 (O_893,N_9958,N_9905);
xor UO_894 (O_894,N_9971,N_9979);
or UO_895 (O_895,N_9957,N_9942);
nand UO_896 (O_896,N_9901,N_9991);
xnor UO_897 (O_897,N_9984,N_9946);
xnor UO_898 (O_898,N_9995,N_9925);
xor UO_899 (O_899,N_9967,N_9924);
nor UO_900 (O_900,N_9950,N_9986);
nand UO_901 (O_901,N_9978,N_9954);
or UO_902 (O_902,N_9935,N_9983);
or UO_903 (O_903,N_9992,N_9934);
or UO_904 (O_904,N_9977,N_9962);
nor UO_905 (O_905,N_9957,N_9900);
xnor UO_906 (O_906,N_9912,N_9953);
and UO_907 (O_907,N_9968,N_9953);
xor UO_908 (O_908,N_9943,N_9910);
and UO_909 (O_909,N_9973,N_9908);
nand UO_910 (O_910,N_9931,N_9992);
nand UO_911 (O_911,N_9975,N_9981);
nand UO_912 (O_912,N_9965,N_9985);
xnor UO_913 (O_913,N_9978,N_9904);
and UO_914 (O_914,N_9993,N_9909);
nand UO_915 (O_915,N_9968,N_9973);
nand UO_916 (O_916,N_9957,N_9906);
or UO_917 (O_917,N_9988,N_9986);
xor UO_918 (O_918,N_9900,N_9932);
nand UO_919 (O_919,N_9965,N_9917);
nor UO_920 (O_920,N_9941,N_9977);
xnor UO_921 (O_921,N_9954,N_9907);
nand UO_922 (O_922,N_9997,N_9900);
and UO_923 (O_923,N_9941,N_9986);
nand UO_924 (O_924,N_9929,N_9963);
or UO_925 (O_925,N_9966,N_9991);
nand UO_926 (O_926,N_9903,N_9994);
and UO_927 (O_927,N_9929,N_9935);
or UO_928 (O_928,N_9954,N_9986);
or UO_929 (O_929,N_9910,N_9988);
and UO_930 (O_930,N_9993,N_9998);
xnor UO_931 (O_931,N_9941,N_9970);
xnor UO_932 (O_932,N_9971,N_9929);
xnor UO_933 (O_933,N_9988,N_9958);
nand UO_934 (O_934,N_9964,N_9997);
and UO_935 (O_935,N_9992,N_9974);
nor UO_936 (O_936,N_9967,N_9913);
and UO_937 (O_937,N_9917,N_9935);
and UO_938 (O_938,N_9945,N_9933);
nand UO_939 (O_939,N_9928,N_9980);
and UO_940 (O_940,N_9917,N_9928);
and UO_941 (O_941,N_9964,N_9914);
nand UO_942 (O_942,N_9992,N_9933);
nand UO_943 (O_943,N_9941,N_9908);
and UO_944 (O_944,N_9986,N_9984);
xor UO_945 (O_945,N_9991,N_9928);
nand UO_946 (O_946,N_9989,N_9929);
and UO_947 (O_947,N_9937,N_9984);
or UO_948 (O_948,N_9939,N_9977);
nor UO_949 (O_949,N_9955,N_9988);
xnor UO_950 (O_950,N_9909,N_9982);
or UO_951 (O_951,N_9910,N_9955);
xor UO_952 (O_952,N_9969,N_9953);
and UO_953 (O_953,N_9974,N_9913);
nor UO_954 (O_954,N_9952,N_9946);
and UO_955 (O_955,N_9987,N_9956);
and UO_956 (O_956,N_9928,N_9920);
nand UO_957 (O_957,N_9911,N_9955);
nand UO_958 (O_958,N_9932,N_9963);
xnor UO_959 (O_959,N_9983,N_9921);
nor UO_960 (O_960,N_9972,N_9929);
nor UO_961 (O_961,N_9930,N_9945);
and UO_962 (O_962,N_9984,N_9935);
nand UO_963 (O_963,N_9955,N_9971);
or UO_964 (O_964,N_9929,N_9902);
or UO_965 (O_965,N_9923,N_9975);
nor UO_966 (O_966,N_9976,N_9981);
xnor UO_967 (O_967,N_9916,N_9959);
xnor UO_968 (O_968,N_9991,N_9951);
and UO_969 (O_969,N_9924,N_9930);
or UO_970 (O_970,N_9958,N_9999);
nand UO_971 (O_971,N_9923,N_9916);
or UO_972 (O_972,N_9977,N_9938);
nor UO_973 (O_973,N_9902,N_9911);
xnor UO_974 (O_974,N_9941,N_9904);
xnor UO_975 (O_975,N_9979,N_9956);
xnor UO_976 (O_976,N_9907,N_9966);
xor UO_977 (O_977,N_9961,N_9949);
xor UO_978 (O_978,N_9923,N_9968);
xor UO_979 (O_979,N_9946,N_9949);
xnor UO_980 (O_980,N_9909,N_9976);
xnor UO_981 (O_981,N_9999,N_9959);
nor UO_982 (O_982,N_9944,N_9912);
and UO_983 (O_983,N_9953,N_9946);
xnor UO_984 (O_984,N_9977,N_9978);
xor UO_985 (O_985,N_9921,N_9978);
or UO_986 (O_986,N_9911,N_9967);
nand UO_987 (O_987,N_9919,N_9935);
xnor UO_988 (O_988,N_9965,N_9939);
xnor UO_989 (O_989,N_9927,N_9990);
or UO_990 (O_990,N_9934,N_9921);
nand UO_991 (O_991,N_9904,N_9998);
nor UO_992 (O_992,N_9954,N_9959);
nor UO_993 (O_993,N_9903,N_9916);
nand UO_994 (O_994,N_9917,N_9943);
nand UO_995 (O_995,N_9910,N_9920);
xnor UO_996 (O_996,N_9937,N_9950);
or UO_997 (O_997,N_9956,N_9915);
or UO_998 (O_998,N_9909,N_9990);
nand UO_999 (O_999,N_9982,N_9929);
and UO_1000 (O_1000,N_9916,N_9989);
and UO_1001 (O_1001,N_9909,N_9953);
nor UO_1002 (O_1002,N_9987,N_9917);
nor UO_1003 (O_1003,N_9974,N_9972);
or UO_1004 (O_1004,N_9917,N_9985);
nor UO_1005 (O_1005,N_9950,N_9992);
or UO_1006 (O_1006,N_9963,N_9942);
nor UO_1007 (O_1007,N_9970,N_9959);
nand UO_1008 (O_1008,N_9950,N_9973);
nand UO_1009 (O_1009,N_9916,N_9944);
nand UO_1010 (O_1010,N_9943,N_9905);
or UO_1011 (O_1011,N_9921,N_9992);
nor UO_1012 (O_1012,N_9931,N_9933);
nand UO_1013 (O_1013,N_9967,N_9981);
and UO_1014 (O_1014,N_9959,N_9967);
nand UO_1015 (O_1015,N_9923,N_9977);
or UO_1016 (O_1016,N_9929,N_9913);
and UO_1017 (O_1017,N_9934,N_9945);
nor UO_1018 (O_1018,N_9963,N_9943);
nand UO_1019 (O_1019,N_9954,N_9930);
nand UO_1020 (O_1020,N_9998,N_9980);
xnor UO_1021 (O_1021,N_9945,N_9948);
nor UO_1022 (O_1022,N_9942,N_9960);
nor UO_1023 (O_1023,N_9979,N_9903);
nand UO_1024 (O_1024,N_9935,N_9927);
or UO_1025 (O_1025,N_9981,N_9923);
xor UO_1026 (O_1026,N_9920,N_9906);
xor UO_1027 (O_1027,N_9928,N_9900);
nand UO_1028 (O_1028,N_9954,N_9965);
nor UO_1029 (O_1029,N_9902,N_9942);
nand UO_1030 (O_1030,N_9977,N_9947);
or UO_1031 (O_1031,N_9909,N_9955);
and UO_1032 (O_1032,N_9970,N_9982);
nand UO_1033 (O_1033,N_9925,N_9986);
xor UO_1034 (O_1034,N_9960,N_9938);
xnor UO_1035 (O_1035,N_9909,N_9941);
xor UO_1036 (O_1036,N_9975,N_9906);
nor UO_1037 (O_1037,N_9918,N_9998);
and UO_1038 (O_1038,N_9945,N_9936);
xor UO_1039 (O_1039,N_9965,N_9948);
nor UO_1040 (O_1040,N_9914,N_9921);
nor UO_1041 (O_1041,N_9963,N_9989);
and UO_1042 (O_1042,N_9962,N_9972);
nand UO_1043 (O_1043,N_9945,N_9976);
nor UO_1044 (O_1044,N_9991,N_9984);
or UO_1045 (O_1045,N_9959,N_9939);
and UO_1046 (O_1046,N_9984,N_9936);
xor UO_1047 (O_1047,N_9998,N_9910);
and UO_1048 (O_1048,N_9988,N_9915);
and UO_1049 (O_1049,N_9906,N_9945);
xor UO_1050 (O_1050,N_9928,N_9918);
xor UO_1051 (O_1051,N_9998,N_9903);
nand UO_1052 (O_1052,N_9934,N_9962);
nand UO_1053 (O_1053,N_9929,N_9942);
nor UO_1054 (O_1054,N_9942,N_9916);
xor UO_1055 (O_1055,N_9960,N_9992);
or UO_1056 (O_1056,N_9938,N_9989);
xor UO_1057 (O_1057,N_9911,N_9968);
nand UO_1058 (O_1058,N_9980,N_9958);
and UO_1059 (O_1059,N_9953,N_9922);
or UO_1060 (O_1060,N_9967,N_9953);
or UO_1061 (O_1061,N_9941,N_9990);
xor UO_1062 (O_1062,N_9956,N_9978);
xnor UO_1063 (O_1063,N_9977,N_9982);
nor UO_1064 (O_1064,N_9978,N_9941);
and UO_1065 (O_1065,N_9951,N_9941);
xor UO_1066 (O_1066,N_9919,N_9993);
nand UO_1067 (O_1067,N_9988,N_9926);
and UO_1068 (O_1068,N_9941,N_9961);
nand UO_1069 (O_1069,N_9924,N_9995);
nand UO_1070 (O_1070,N_9910,N_9936);
nand UO_1071 (O_1071,N_9996,N_9948);
nand UO_1072 (O_1072,N_9940,N_9921);
or UO_1073 (O_1073,N_9945,N_9997);
xor UO_1074 (O_1074,N_9964,N_9965);
nor UO_1075 (O_1075,N_9908,N_9975);
xnor UO_1076 (O_1076,N_9924,N_9989);
or UO_1077 (O_1077,N_9966,N_9979);
and UO_1078 (O_1078,N_9988,N_9938);
and UO_1079 (O_1079,N_9920,N_9984);
xor UO_1080 (O_1080,N_9953,N_9985);
xnor UO_1081 (O_1081,N_9930,N_9979);
nand UO_1082 (O_1082,N_9984,N_9921);
nor UO_1083 (O_1083,N_9913,N_9990);
and UO_1084 (O_1084,N_9996,N_9910);
nor UO_1085 (O_1085,N_9966,N_9902);
nand UO_1086 (O_1086,N_9913,N_9973);
or UO_1087 (O_1087,N_9995,N_9983);
nor UO_1088 (O_1088,N_9972,N_9994);
nor UO_1089 (O_1089,N_9979,N_9980);
or UO_1090 (O_1090,N_9956,N_9968);
or UO_1091 (O_1091,N_9924,N_9901);
nand UO_1092 (O_1092,N_9901,N_9942);
nand UO_1093 (O_1093,N_9913,N_9933);
nand UO_1094 (O_1094,N_9915,N_9970);
xnor UO_1095 (O_1095,N_9932,N_9940);
or UO_1096 (O_1096,N_9970,N_9926);
or UO_1097 (O_1097,N_9912,N_9981);
nor UO_1098 (O_1098,N_9959,N_9988);
nand UO_1099 (O_1099,N_9948,N_9973);
xor UO_1100 (O_1100,N_9939,N_9913);
nand UO_1101 (O_1101,N_9941,N_9950);
nand UO_1102 (O_1102,N_9928,N_9907);
and UO_1103 (O_1103,N_9967,N_9958);
or UO_1104 (O_1104,N_9911,N_9983);
and UO_1105 (O_1105,N_9970,N_9972);
nor UO_1106 (O_1106,N_9960,N_9975);
and UO_1107 (O_1107,N_9998,N_9979);
nand UO_1108 (O_1108,N_9979,N_9986);
nor UO_1109 (O_1109,N_9930,N_9940);
nand UO_1110 (O_1110,N_9957,N_9983);
or UO_1111 (O_1111,N_9961,N_9954);
or UO_1112 (O_1112,N_9926,N_9908);
xor UO_1113 (O_1113,N_9901,N_9995);
and UO_1114 (O_1114,N_9934,N_9982);
nor UO_1115 (O_1115,N_9996,N_9905);
nand UO_1116 (O_1116,N_9981,N_9937);
or UO_1117 (O_1117,N_9955,N_9981);
nand UO_1118 (O_1118,N_9969,N_9921);
and UO_1119 (O_1119,N_9962,N_9980);
nand UO_1120 (O_1120,N_9904,N_9925);
or UO_1121 (O_1121,N_9930,N_9923);
or UO_1122 (O_1122,N_9969,N_9995);
and UO_1123 (O_1123,N_9932,N_9945);
xor UO_1124 (O_1124,N_9908,N_9919);
nor UO_1125 (O_1125,N_9993,N_9999);
or UO_1126 (O_1126,N_9965,N_9926);
and UO_1127 (O_1127,N_9923,N_9948);
and UO_1128 (O_1128,N_9924,N_9994);
or UO_1129 (O_1129,N_9927,N_9938);
nand UO_1130 (O_1130,N_9978,N_9988);
or UO_1131 (O_1131,N_9928,N_9901);
nand UO_1132 (O_1132,N_9902,N_9900);
xnor UO_1133 (O_1133,N_9993,N_9947);
nand UO_1134 (O_1134,N_9982,N_9920);
or UO_1135 (O_1135,N_9909,N_9906);
xnor UO_1136 (O_1136,N_9928,N_9983);
xor UO_1137 (O_1137,N_9971,N_9923);
or UO_1138 (O_1138,N_9986,N_9927);
and UO_1139 (O_1139,N_9997,N_9907);
and UO_1140 (O_1140,N_9971,N_9906);
or UO_1141 (O_1141,N_9970,N_9928);
or UO_1142 (O_1142,N_9912,N_9931);
nand UO_1143 (O_1143,N_9922,N_9902);
or UO_1144 (O_1144,N_9949,N_9943);
nand UO_1145 (O_1145,N_9934,N_9968);
or UO_1146 (O_1146,N_9994,N_9943);
nand UO_1147 (O_1147,N_9916,N_9972);
or UO_1148 (O_1148,N_9930,N_9961);
nand UO_1149 (O_1149,N_9989,N_9967);
or UO_1150 (O_1150,N_9955,N_9998);
or UO_1151 (O_1151,N_9960,N_9901);
xnor UO_1152 (O_1152,N_9929,N_9969);
nand UO_1153 (O_1153,N_9905,N_9904);
xnor UO_1154 (O_1154,N_9952,N_9935);
nand UO_1155 (O_1155,N_9919,N_9980);
or UO_1156 (O_1156,N_9904,N_9976);
xnor UO_1157 (O_1157,N_9994,N_9906);
nor UO_1158 (O_1158,N_9958,N_9941);
or UO_1159 (O_1159,N_9997,N_9901);
nand UO_1160 (O_1160,N_9931,N_9934);
and UO_1161 (O_1161,N_9995,N_9904);
xor UO_1162 (O_1162,N_9928,N_9955);
and UO_1163 (O_1163,N_9941,N_9932);
and UO_1164 (O_1164,N_9915,N_9934);
and UO_1165 (O_1165,N_9910,N_9967);
xnor UO_1166 (O_1166,N_9933,N_9924);
nand UO_1167 (O_1167,N_9949,N_9942);
xnor UO_1168 (O_1168,N_9930,N_9975);
nor UO_1169 (O_1169,N_9942,N_9931);
nor UO_1170 (O_1170,N_9914,N_9901);
nor UO_1171 (O_1171,N_9955,N_9932);
nor UO_1172 (O_1172,N_9963,N_9910);
nor UO_1173 (O_1173,N_9922,N_9999);
nand UO_1174 (O_1174,N_9909,N_9916);
nor UO_1175 (O_1175,N_9909,N_9985);
or UO_1176 (O_1176,N_9980,N_9982);
nor UO_1177 (O_1177,N_9973,N_9957);
or UO_1178 (O_1178,N_9954,N_9949);
or UO_1179 (O_1179,N_9992,N_9979);
nand UO_1180 (O_1180,N_9979,N_9929);
nor UO_1181 (O_1181,N_9945,N_9957);
xnor UO_1182 (O_1182,N_9991,N_9968);
nor UO_1183 (O_1183,N_9947,N_9971);
or UO_1184 (O_1184,N_9904,N_9967);
xor UO_1185 (O_1185,N_9974,N_9928);
xnor UO_1186 (O_1186,N_9921,N_9938);
nand UO_1187 (O_1187,N_9969,N_9988);
xor UO_1188 (O_1188,N_9973,N_9909);
nor UO_1189 (O_1189,N_9902,N_9927);
xor UO_1190 (O_1190,N_9962,N_9994);
or UO_1191 (O_1191,N_9971,N_9995);
nor UO_1192 (O_1192,N_9903,N_9958);
xor UO_1193 (O_1193,N_9953,N_9988);
or UO_1194 (O_1194,N_9948,N_9982);
nand UO_1195 (O_1195,N_9941,N_9954);
or UO_1196 (O_1196,N_9971,N_9975);
nor UO_1197 (O_1197,N_9933,N_9914);
xor UO_1198 (O_1198,N_9914,N_9953);
and UO_1199 (O_1199,N_9905,N_9981);
xnor UO_1200 (O_1200,N_9925,N_9930);
or UO_1201 (O_1201,N_9959,N_9994);
and UO_1202 (O_1202,N_9905,N_9927);
nand UO_1203 (O_1203,N_9924,N_9959);
nor UO_1204 (O_1204,N_9989,N_9905);
xor UO_1205 (O_1205,N_9958,N_9952);
and UO_1206 (O_1206,N_9974,N_9961);
nand UO_1207 (O_1207,N_9952,N_9941);
nand UO_1208 (O_1208,N_9903,N_9947);
nand UO_1209 (O_1209,N_9995,N_9930);
nand UO_1210 (O_1210,N_9947,N_9944);
xnor UO_1211 (O_1211,N_9972,N_9998);
or UO_1212 (O_1212,N_9968,N_9971);
xnor UO_1213 (O_1213,N_9939,N_9972);
xor UO_1214 (O_1214,N_9974,N_9907);
and UO_1215 (O_1215,N_9993,N_9917);
nand UO_1216 (O_1216,N_9922,N_9940);
or UO_1217 (O_1217,N_9968,N_9974);
and UO_1218 (O_1218,N_9914,N_9957);
xor UO_1219 (O_1219,N_9919,N_9926);
and UO_1220 (O_1220,N_9992,N_9925);
nor UO_1221 (O_1221,N_9952,N_9984);
or UO_1222 (O_1222,N_9971,N_9957);
xnor UO_1223 (O_1223,N_9980,N_9964);
nor UO_1224 (O_1224,N_9994,N_9928);
or UO_1225 (O_1225,N_9916,N_9992);
and UO_1226 (O_1226,N_9927,N_9904);
nor UO_1227 (O_1227,N_9996,N_9913);
nand UO_1228 (O_1228,N_9913,N_9952);
xor UO_1229 (O_1229,N_9966,N_9986);
nor UO_1230 (O_1230,N_9948,N_9956);
and UO_1231 (O_1231,N_9937,N_9990);
or UO_1232 (O_1232,N_9994,N_9900);
xnor UO_1233 (O_1233,N_9938,N_9936);
nand UO_1234 (O_1234,N_9970,N_9913);
xnor UO_1235 (O_1235,N_9941,N_9933);
nor UO_1236 (O_1236,N_9913,N_9919);
and UO_1237 (O_1237,N_9957,N_9984);
xor UO_1238 (O_1238,N_9909,N_9984);
xor UO_1239 (O_1239,N_9907,N_9902);
nand UO_1240 (O_1240,N_9944,N_9903);
nor UO_1241 (O_1241,N_9922,N_9973);
and UO_1242 (O_1242,N_9908,N_9978);
or UO_1243 (O_1243,N_9958,N_9966);
xor UO_1244 (O_1244,N_9920,N_9995);
or UO_1245 (O_1245,N_9915,N_9931);
xor UO_1246 (O_1246,N_9964,N_9949);
xnor UO_1247 (O_1247,N_9991,N_9979);
and UO_1248 (O_1248,N_9981,N_9934);
nand UO_1249 (O_1249,N_9994,N_9919);
xnor UO_1250 (O_1250,N_9975,N_9970);
nor UO_1251 (O_1251,N_9974,N_9954);
nor UO_1252 (O_1252,N_9979,N_9944);
nor UO_1253 (O_1253,N_9910,N_9919);
or UO_1254 (O_1254,N_9970,N_9999);
xor UO_1255 (O_1255,N_9997,N_9999);
nor UO_1256 (O_1256,N_9958,N_9944);
and UO_1257 (O_1257,N_9920,N_9900);
nand UO_1258 (O_1258,N_9919,N_9927);
nand UO_1259 (O_1259,N_9972,N_9988);
nor UO_1260 (O_1260,N_9993,N_9995);
nor UO_1261 (O_1261,N_9939,N_9948);
nor UO_1262 (O_1262,N_9945,N_9991);
nor UO_1263 (O_1263,N_9995,N_9941);
nand UO_1264 (O_1264,N_9946,N_9931);
xnor UO_1265 (O_1265,N_9934,N_9901);
nand UO_1266 (O_1266,N_9945,N_9954);
nand UO_1267 (O_1267,N_9903,N_9912);
nor UO_1268 (O_1268,N_9986,N_9918);
and UO_1269 (O_1269,N_9959,N_9974);
nand UO_1270 (O_1270,N_9985,N_9973);
xor UO_1271 (O_1271,N_9939,N_9942);
xnor UO_1272 (O_1272,N_9938,N_9940);
and UO_1273 (O_1273,N_9913,N_9960);
nor UO_1274 (O_1274,N_9982,N_9943);
or UO_1275 (O_1275,N_9948,N_9924);
nand UO_1276 (O_1276,N_9912,N_9968);
nor UO_1277 (O_1277,N_9992,N_9910);
nand UO_1278 (O_1278,N_9953,N_9972);
nor UO_1279 (O_1279,N_9921,N_9952);
or UO_1280 (O_1280,N_9915,N_9978);
and UO_1281 (O_1281,N_9967,N_9998);
nor UO_1282 (O_1282,N_9976,N_9934);
nor UO_1283 (O_1283,N_9970,N_9945);
and UO_1284 (O_1284,N_9952,N_9942);
nand UO_1285 (O_1285,N_9913,N_9920);
and UO_1286 (O_1286,N_9953,N_9994);
xnor UO_1287 (O_1287,N_9912,N_9939);
nand UO_1288 (O_1288,N_9986,N_9933);
or UO_1289 (O_1289,N_9920,N_9941);
nand UO_1290 (O_1290,N_9987,N_9976);
xnor UO_1291 (O_1291,N_9942,N_9971);
or UO_1292 (O_1292,N_9978,N_9999);
or UO_1293 (O_1293,N_9929,N_9955);
nand UO_1294 (O_1294,N_9995,N_9966);
nor UO_1295 (O_1295,N_9959,N_9948);
xnor UO_1296 (O_1296,N_9940,N_9946);
nor UO_1297 (O_1297,N_9946,N_9993);
nand UO_1298 (O_1298,N_9973,N_9930);
xnor UO_1299 (O_1299,N_9921,N_9961);
or UO_1300 (O_1300,N_9937,N_9931);
nor UO_1301 (O_1301,N_9914,N_9977);
nand UO_1302 (O_1302,N_9930,N_9955);
or UO_1303 (O_1303,N_9995,N_9942);
or UO_1304 (O_1304,N_9951,N_9926);
nand UO_1305 (O_1305,N_9915,N_9990);
nand UO_1306 (O_1306,N_9953,N_9927);
and UO_1307 (O_1307,N_9968,N_9972);
or UO_1308 (O_1308,N_9925,N_9951);
or UO_1309 (O_1309,N_9992,N_9963);
and UO_1310 (O_1310,N_9928,N_9962);
or UO_1311 (O_1311,N_9982,N_9901);
nand UO_1312 (O_1312,N_9952,N_9947);
nand UO_1313 (O_1313,N_9951,N_9973);
xnor UO_1314 (O_1314,N_9905,N_9912);
nor UO_1315 (O_1315,N_9946,N_9939);
xnor UO_1316 (O_1316,N_9995,N_9912);
nor UO_1317 (O_1317,N_9958,N_9923);
xor UO_1318 (O_1318,N_9968,N_9932);
or UO_1319 (O_1319,N_9986,N_9926);
xor UO_1320 (O_1320,N_9910,N_9950);
xnor UO_1321 (O_1321,N_9925,N_9912);
xor UO_1322 (O_1322,N_9956,N_9995);
and UO_1323 (O_1323,N_9910,N_9995);
and UO_1324 (O_1324,N_9984,N_9965);
nand UO_1325 (O_1325,N_9938,N_9984);
or UO_1326 (O_1326,N_9915,N_9929);
nor UO_1327 (O_1327,N_9918,N_9921);
nor UO_1328 (O_1328,N_9974,N_9983);
nand UO_1329 (O_1329,N_9924,N_9990);
nor UO_1330 (O_1330,N_9975,N_9926);
xor UO_1331 (O_1331,N_9978,N_9906);
nor UO_1332 (O_1332,N_9906,N_9982);
or UO_1333 (O_1333,N_9998,N_9962);
or UO_1334 (O_1334,N_9932,N_9962);
or UO_1335 (O_1335,N_9967,N_9969);
or UO_1336 (O_1336,N_9928,N_9985);
nor UO_1337 (O_1337,N_9905,N_9947);
or UO_1338 (O_1338,N_9956,N_9941);
nand UO_1339 (O_1339,N_9983,N_9948);
nor UO_1340 (O_1340,N_9914,N_9978);
nand UO_1341 (O_1341,N_9997,N_9923);
nor UO_1342 (O_1342,N_9907,N_9905);
and UO_1343 (O_1343,N_9965,N_9908);
or UO_1344 (O_1344,N_9921,N_9974);
xnor UO_1345 (O_1345,N_9960,N_9979);
or UO_1346 (O_1346,N_9989,N_9935);
nor UO_1347 (O_1347,N_9940,N_9993);
or UO_1348 (O_1348,N_9930,N_9957);
nand UO_1349 (O_1349,N_9962,N_9983);
xnor UO_1350 (O_1350,N_9911,N_9948);
xnor UO_1351 (O_1351,N_9910,N_9941);
or UO_1352 (O_1352,N_9926,N_9906);
or UO_1353 (O_1353,N_9934,N_9965);
nor UO_1354 (O_1354,N_9925,N_9983);
and UO_1355 (O_1355,N_9900,N_9934);
nand UO_1356 (O_1356,N_9975,N_9973);
and UO_1357 (O_1357,N_9960,N_9973);
nand UO_1358 (O_1358,N_9938,N_9982);
nor UO_1359 (O_1359,N_9937,N_9941);
xnor UO_1360 (O_1360,N_9988,N_9991);
nor UO_1361 (O_1361,N_9941,N_9982);
nand UO_1362 (O_1362,N_9906,N_9916);
and UO_1363 (O_1363,N_9965,N_9942);
xor UO_1364 (O_1364,N_9935,N_9908);
or UO_1365 (O_1365,N_9912,N_9927);
and UO_1366 (O_1366,N_9912,N_9962);
nor UO_1367 (O_1367,N_9937,N_9907);
or UO_1368 (O_1368,N_9960,N_9955);
or UO_1369 (O_1369,N_9918,N_9993);
or UO_1370 (O_1370,N_9947,N_9924);
nor UO_1371 (O_1371,N_9923,N_9915);
and UO_1372 (O_1372,N_9912,N_9961);
nor UO_1373 (O_1373,N_9974,N_9957);
and UO_1374 (O_1374,N_9931,N_9911);
and UO_1375 (O_1375,N_9927,N_9949);
xnor UO_1376 (O_1376,N_9956,N_9921);
nor UO_1377 (O_1377,N_9927,N_9994);
and UO_1378 (O_1378,N_9952,N_9900);
and UO_1379 (O_1379,N_9934,N_9905);
or UO_1380 (O_1380,N_9914,N_9948);
or UO_1381 (O_1381,N_9972,N_9919);
or UO_1382 (O_1382,N_9974,N_9917);
and UO_1383 (O_1383,N_9958,N_9987);
and UO_1384 (O_1384,N_9983,N_9970);
nand UO_1385 (O_1385,N_9938,N_9992);
or UO_1386 (O_1386,N_9939,N_9931);
or UO_1387 (O_1387,N_9976,N_9914);
and UO_1388 (O_1388,N_9954,N_9905);
nor UO_1389 (O_1389,N_9933,N_9966);
nor UO_1390 (O_1390,N_9980,N_9999);
xnor UO_1391 (O_1391,N_9944,N_9924);
nor UO_1392 (O_1392,N_9938,N_9918);
xnor UO_1393 (O_1393,N_9955,N_9990);
and UO_1394 (O_1394,N_9921,N_9965);
and UO_1395 (O_1395,N_9975,N_9920);
or UO_1396 (O_1396,N_9962,N_9964);
xor UO_1397 (O_1397,N_9973,N_9946);
nor UO_1398 (O_1398,N_9950,N_9907);
and UO_1399 (O_1399,N_9950,N_9989);
nor UO_1400 (O_1400,N_9974,N_9996);
xor UO_1401 (O_1401,N_9932,N_9923);
or UO_1402 (O_1402,N_9925,N_9902);
nor UO_1403 (O_1403,N_9915,N_9961);
nand UO_1404 (O_1404,N_9941,N_9980);
nor UO_1405 (O_1405,N_9916,N_9920);
or UO_1406 (O_1406,N_9914,N_9973);
or UO_1407 (O_1407,N_9906,N_9986);
nand UO_1408 (O_1408,N_9978,N_9928);
nor UO_1409 (O_1409,N_9933,N_9946);
and UO_1410 (O_1410,N_9947,N_9959);
and UO_1411 (O_1411,N_9983,N_9951);
xnor UO_1412 (O_1412,N_9915,N_9974);
nand UO_1413 (O_1413,N_9949,N_9970);
xnor UO_1414 (O_1414,N_9942,N_9956);
xor UO_1415 (O_1415,N_9981,N_9945);
or UO_1416 (O_1416,N_9932,N_9927);
xor UO_1417 (O_1417,N_9974,N_9986);
nand UO_1418 (O_1418,N_9969,N_9936);
nand UO_1419 (O_1419,N_9929,N_9965);
nor UO_1420 (O_1420,N_9960,N_9996);
nor UO_1421 (O_1421,N_9928,N_9932);
nor UO_1422 (O_1422,N_9995,N_9951);
nand UO_1423 (O_1423,N_9990,N_9974);
or UO_1424 (O_1424,N_9954,N_9939);
nand UO_1425 (O_1425,N_9909,N_9998);
nand UO_1426 (O_1426,N_9960,N_9994);
xnor UO_1427 (O_1427,N_9998,N_9956);
or UO_1428 (O_1428,N_9957,N_9981);
and UO_1429 (O_1429,N_9924,N_9927);
xnor UO_1430 (O_1430,N_9935,N_9971);
nand UO_1431 (O_1431,N_9935,N_9906);
nor UO_1432 (O_1432,N_9977,N_9988);
xor UO_1433 (O_1433,N_9966,N_9989);
or UO_1434 (O_1434,N_9996,N_9936);
nor UO_1435 (O_1435,N_9943,N_9971);
xnor UO_1436 (O_1436,N_9934,N_9913);
xnor UO_1437 (O_1437,N_9975,N_9907);
or UO_1438 (O_1438,N_9988,N_9946);
nor UO_1439 (O_1439,N_9978,N_9942);
nand UO_1440 (O_1440,N_9913,N_9914);
xnor UO_1441 (O_1441,N_9905,N_9923);
or UO_1442 (O_1442,N_9917,N_9946);
nand UO_1443 (O_1443,N_9939,N_9929);
xnor UO_1444 (O_1444,N_9983,N_9950);
and UO_1445 (O_1445,N_9994,N_9963);
nand UO_1446 (O_1446,N_9987,N_9929);
or UO_1447 (O_1447,N_9979,N_9932);
nand UO_1448 (O_1448,N_9955,N_9922);
xnor UO_1449 (O_1449,N_9988,N_9916);
or UO_1450 (O_1450,N_9971,N_9909);
and UO_1451 (O_1451,N_9999,N_9937);
or UO_1452 (O_1452,N_9949,N_9974);
nor UO_1453 (O_1453,N_9985,N_9906);
nor UO_1454 (O_1454,N_9966,N_9963);
nor UO_1455 (O_1455,N_9919,N_9922);
nand UO_1456 (O_1456,N_9983,N_9947);
and UO_1457 (O_1457,N_9958,N_9909);
or UO_1458 (O_1458,N_9974,N_9940);
xnor UO_1459 (O_1459,N_9971,N_9903);
xnor UO_1460 (O_1460,N_9930,N_9950);
nand UO_1461 (O_1461,N_9901,N_9999);
nand UO_1462 (O_1462,N_9985,N_9999);
nor UO_1463 (O_1463,N_9926,N_9900);
xor UO_1464 (O_1464,N_9995,N_9906);
nor UO_1465 (O_1465,N_9909,N_9991);
and UO_1466 (O_1466,N_9949,N_9903);
and UO_1467 (O_1467,N_9967,N_9991);
or UO_1468 (O_1468,N_9948,N_9952);
or UO_1469 (O_1469,N_9906,N_9949);
and UO_1470 (O_1470,N_9974,N_9989);
or UO_1471 (O_1471,N_9992,N_9965);
or UO_1472 (O_1472,N_9966,N_9931);
xor UO_1473 (O_1473,N_9985,N_9902);
nor UO_1474 (O_1474,N_9928,N_9926);
or UO_1475 (O_1475,N_9911,N_9913);
or UO_1476 (O_1476,N_9908,N_9913);
nand UO_1477 (O_1477,N_9918,N_9982);
or UO_1478 (O_1478,N_9926,N_9985);
nand UO_1479 (O_1479,N_9976,N_9936);
or UO_1480 (O_1480,N_9985,N_9997);
nand UO_1481 (O_1481,N_9932,N_9944);
nor UO_1482 (O_1482,N_9953,N_9911);
or UO_1483 (O_1483,N_9941,N_9901);
nand UO_1484 (O_1484,N_9908,N_9907);
nor UO_1485 (O_1485,N_9907,N_9982);
nor UO_1486 (O_1486,N_9989,N_9998);
nor UO_1487 (O_1487,N_9914,N_9927);
nor UO_1488 (O_1488,N_9901,N_9958);
nand UO_1489 (O_1489,N_9927,N_9911);
nor UO_1490 (O_1490,N_9980,N_9961);
and UO_1491 (O_1491,N_9940,N_9987);
and UO_1492 (O_1492,N_9975,N_9996);
nor UO_1493 (O_1493,N_9937,N_9913);
and UO_1494 (O_1494,N_9919,N_9923);
and UO_1495 (O_1495,N_9949,N_9921);
nor UO_1496 (O_1496,N_9928,N_9940);
and UO_1497 (O_1497,N_9904,N_9966);
nand UO_1498 (O_1498,N_9960,N_9968);
nand UO_1499 (O_1499,N_9940,N_9904);
endmodule