module basic_2000_20000_2500_125_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_878,In_820);
nor U1 (N_1,In_1257,In_1623);
nand U2 (N_2,In_1084,In_286);
nand U3 (N_3,In_297,In_755);
and U4 (N_4,In_553,In_1289);
nor U5 (N_5,In_737,In_638);
or U6 (N_6,In_1189,In_70);
nor U7 (N_7,In_8,In_852);
xor U8 (N_8,In_748,In_1833);
and U9 (N_9,In_199,In_200);
nor U10 (N_10,In_1192,In_1901);
nand U11 (N_11,In_881,In_356);
nor U12 (N_12,In_1430,In_1755);
nor U13 (N_13,In_1645,In_29);
xnor U14 (N_14,In_1991,In_54);
nor U15 (N_15,In_1500,In_1984);
and U16 (N_16,In_583,In_656);
nand U17 (N_17,In_1043,In_1550);
nor U18 (N_18,In_733,In_438);
xor U19 (N_19,In_260,In_636);
xnor U20 (N_20,In_699,In_1770);
nor U21 (N_21,In_845,In_252);
and U22 (N_22,In_538,In_1543);
or U23 (N_23,In_1752,In_360);
nor U24 (N_24,In_370,In_138);
xor U25 (N_25,In_729,In_1126);
or U26 (N_26,In_9,In_402);
or U27 (N_27,In_1506,In_713);
nor U28 (N_28,In_279,In_1869);
xnor U29 (N_29,In_509,In_110);
or U30 (N_30,In_1951,In_1692);
nand U31 (N_31,In_162,In_1916);
nand U32 (N_32,In_940,In_1021);
and U33 (N_33,In_854,In_452);
nand U34 (N_34,In_744,In_1022);
nand U35 (N_35,In_962,In_652);
and U36 (N_36,In_475,In_43);
xnor U37 (N_37,In_499,In_1166);
and U38 (N_38,In_909,In_479);
xor U39 (N_39,In_1883,In_1710);
nand U40 (N_40,In_856,In_1317);
and U41 (N_41,In_1024,In_145);
xor U42 (N_42,In_1779,In_253);
nor U43 (N_43,In_451,In_1254);
and U44 (N_44,In_290,In_417);
nand U45 (N_45,In_1130,In_365);
or U46 (N_46,In_1591,In_597);
nor U47 (N_47,In_1854,In_1820);
xor U48 (N_48,In_1015,In_798);
or U49 (N_49,In_1338,In_1025);
nand U50 (N_50,In_1844,In_24);
nor U51 (N_51,In_968,In_1896);
xnor U52 (N_52,In_1594,In_93);
nor U53 (N_53,In_492,In_1846);
or U54 (N_54,In_1640,In_600);
nand U55 (N_55,In_503,In_1754);
nor U56 (N_56,In_179,In_735);
nand U57 (N_57,In_1475,In_423);
xor U58 (N_58,In_1644,In_1147);
xor U59 (N_59,In_1913,In_953);
or U60 (N_60,In_1787,In_1476);
nor U61 (N_61,In_604,In_855);
and U62 (N_62,In_27,In_231);
or U63 (N_63,In_922,In_689);
nor U64 (N_64,In_1961,In_1701);
xor U65 (N_65,In_1059,In_1208);
nand U66 (N_66,In_1628,In_892);
or U67 (N_67,In_1228,In_1784);
nor U68 (N_68,In_530,In_413);
and U69 (N_69,In_578,In_384);
and U70 (N_70,In_811,In_944);
xor U71 (N_71,In_342,In_774);
nand U72 (N_72,In_1538,In_895);
xor U73 (N_73,In_1344,In_1255);
nor U74 (N_74,In_144,In_428);
or U75 (N_75,In_400,In_1705);
and U76 (N_76,In_1541,In_1213);
nand U77 (N_77,In_1034,In_1658);
and U78 (N_78,In_640,In_1797);
nor U79 (N_79,In_866,In_63);
xor U80 (N_80,In_694,In_222);
or U81 (N_81,In_603,In_294);
xnor U82 (N_82,In_26,In_230);
or U83 (N_83,In_842,In_1112);
xor U84 (N_84,In_91,In_1146);
nor U85 (N_85,In_1005,In_605);
or U86 (N_86,In_1927,In_679);
and U87 (N_87,In_1220,In_1125);
nor U88 (N_88,In_1935,In_1567);
and U89 (N_89,In_4,In_317);
xnor U90 (N_90,In_1118,In_1686);
nor U91 (N_91,In_271,In_427);
nor U92 (N_92,In_1744,In_1008);
xor U93 (N_93,In_965,In_1378);
nand U94 (N_94,In_513,In_708);
or U95 (N_95,In_1574,In_1109);
nor U96 (N_96,In_1900,In_1994);
nor U97 (N_97,In_1948,In_1096);
nor U98 (N_98,In_305,In_1424);
nor U99 (N_99,In_128,In_1877);
nand U100 (N_100,In_998,In_268);
nor U101 (N_101,In_1922,In_1072);
nand U102 (N_102,In_206,In_169);
nor U103 (N_103,In_1173,In_1428);
nor U104 (N_104,In_1942,In_921);
or U105 (N_105,In_1646,In_1694);
nor U106 (N_106,In_1577,In_1753);
nor U107 (N_107,In_308,In_867);
or U108 (N_108,In_1825,In_812);
and U109 (N_109,In_361,In_363);
nand U110 (N_110,In_900,In_450);
nand U111 (N_111,In_767,In_1078);
or U112 (N_112,In_1389,In_550);
nand U113 (N_113,In_1725,In_107);
or U114 (N_114,In_1308,In_0);
nand U115 (N_115,In_1136,In_569);
nand U116 (N_116,In_1265,In_1131);
and U117 (N_117,In_254,In_1669);
and U118 (N_118,In_701,In_505);
and U119 (N_119,In_81,In_1803);
and U120 (N_120,In_1572,In_267);
xnor U121 (N_121,In_1127,In_341);
xor U122 (N_122,In_557,In_512);
nand U123 (N_123,In_1480,In_1938);
or U124 (N_124,In_1724,In_506);
and U125 (N_125,In_25,In_1741);
nor U126 (N_126,In_34,In_580);
or U127 (N_127,In_776,In_1287);
nor U128 (N_128,In_1397,In_1926);
or U129 (N_129,In_468,In_1680);
and U130 (N_130,In_44,In_1761);
nand U131 (N_131,In_657,In_1183);
nor U132 (N_132,In_1246,In_1674);
nor U133 (N_133,In_1821,In_1046);
or U134 (N_134,In_1798,In_502);
nor U135 (N_135,In_534,In_1056);
xnor U136 (N_136,In_1226,In_695);
or U137 (N_137,In_1533,In_1108);
or U138 (N_138,In_644,In_234);
nor U139 (N_139,In_1531,In_788);
and U140 (N_140,In_1740,In_564);
nand U141 (N_141,In_609,In_2);
and U142 (N_142,In_164,In_667);
and U143 (N_143,In_326,In_1930);
nor U144 (N_144,In_1429,In_1720);
nand U145 (N_145,In_936,In_122);
nor U146 (N_146,In_1449,In_1241);
nand U147 (N_147,In_1,In_507);
nor U148 (N_148,In_582,In_800);
nor U149 (N_149,In_1876,In_1081);
nand U150 (N_150,In_519,In_246);
xor U151 (N_151,In_727,In_533);
and U152 (N_152,In_1000,In_374);
nand U153 (N_153,In_276,In_1564);
nand U154 (N_154,In_781,In_1573);
and U155 (N_155,In_621,In_875);
or U156 (N_156,In_1988,In_586);
xor U157 (N_157,In_1184,In_1718);
nor U158 (N_158,In_1302,In_17);
or U159 (N_159,In_1617,In_315);
or U160 (N_160,N_24,In_763);
xor U161 (N_161,In_802,In_1408);
nand U162 (N_162,In_823,In_1012);
nor U163 (N_163,In_1945,In_1041);
nand U164 (N_164,In_1151,In_990);
nor U165 (N_165,In_1283,In_1132);
xnor U166 (N_166,In_435,In_1641);
and U167 (N_167,In_379,In_217);
or U168 (N_168,In_345,In_1160);
nand U169 (N_169,In_381,In_929);
and U170 (N_170,In_1479,In_1445);
xnor U171 (N_171,In_1978,In_284);
xor U172 (N_172,In_1831,In_573);
xnor U173 (N_173,In_899,In_483);
and U174 (N_174,In_157,In_1726);
or U175 (N_175,In_399,In_177);
or U176 (N_176,In_1643,In_992);
xor U177 (N_177,In_1441,In_426);
and U178 (N_178,In_1898,In_1561);
and U179 (N_179,In_184,In_790);
and U180 (N_180,N_43,In_1092);
nand U181 (N_181,In_1366,In_1974);
or U182 (N_182,In_1636,In_602);
and U183 (N_183,In_386,In_1304);
and U184 (N_184,In_1786,In_196);
xor U185 (N_185,In_1460,In_841);
or U186 (N_186,In_1847,In_1235);
xnor U187 (N_187,In_522,In_1867);
nor U188 (N_188,In_510,In_385);
and U189 (N_189,In_433,In_1165);
xor U190 (N_190,In_48,In_406);
and U191 (N_191,In_1764,In_625);
nand U192 (N_192,In_1027,In_1377);
nand U193 (N_193,In_816,In_916);
nand U194 (N_194,In_1952,In_837);
or U195 (N_195,In_1273,N_23);
or U196 (N_196,In_1331,In_526);
nand U197 (N_197,N_2,In_1719);
nor U198 (N_198,In_544,In_313);
nor U199 (N_199,In_293,In_1285);
and U200 (N_200,In_612,In_309);
nor U201 (N_201,In_1153,In_1157);
nor U202 (N_202,In_931,In_1219);
or U203 (N_203,In_686,In_1452);
nor U204 (N_204,In_587,In_1765);
nand U205 (N_205,In_1492,N_0);
nand U206 (N_206,In_1294,In_1487);
nor U207 (N_207,In_847,In_250);
xnor U208 (N_208,In_1070,In_1100);
nor U209 (N_209,N_28,In_444);
nand U210 (N_210,In_559,In_1504);
nand U211 (N_211,In_938,In_38);
nor U212 (N_212,In_1884,In_947);
xnor U213 (N_213,In_1601,In_1528);
or U214 (N_214,In_1722,In_1274);
and U215 (N_215,In_1544,In_996);
nand U216 (N_216,In_988,In_1392);
and U217 (N_217,In_78,N_58);
nand U218 (N_218,In_72,In_683);
nand U219 (N_219,N_106,In_752);
xor U220 (N_220,In_810,In_1734);
nand U221 (N_221,N_66,In_191);
nand U222 (N_222,In_1456,In_1375);
xnor U223 (N_223,In_1608,N_83);
or U224 (N_224,N_50,In_189);
xnor U225 (N_225,In_53,In_368);
nor U226 (N_226,In_1532,In_1879);
nor U227 (N_227,In_1700,In_818);
or U228 (N_228,In_1431,In_760);
nand U229 (N_229,In_887,In_1767);
nand U230 (N_230,In_941,In_1300);
nand U231 (N_231,In_39,N_35);
or U232 (N_232,In_865,In_117);
or U233 (N_233,In_741,In_19);
nor U234 (N_234,In_743,In_487);
nor U235 (N_235,In_80,In_894);
and U236 (N_236,In_1060,In_1966);
or U237 (N_237,In_1447,In_1275);
nor U238 (N_238,N_82,In_1748);
nor U239 (N_239,In_1416,In_1950);
nor U240 (N_240,In_1800,In_1399);
or U241 (N_241,In_1400,In_458);
and U242 (N_242,In_1494,In_1483);
and U243 (N_243,In_407,In_1737);
and U244 (N_244,In_976,In_1298);
nand U245 (N_245,In_1864,In_886);
xor U246 (N_246,In_822,In_1872);
and U247 (N_247,In_1536,In_1326);
nand U248 (N_248,In_872,In_1835);
xnor U249 (N_249,In_396,N_80);
or U250 (N_250,In_615,In_684);
and U251 (N_251,In_651,In_1040);
xnor U252 (N_252,In_724,In_1135);
nor U253 (N_253,In_1816,In_1290);
nor U254 (N_254,In_494,In_1619);
nand U255 (N_255,In_457,In_1868);
and U256 (N_256,In_490,In_1804);
nor U257 (N_257,In_991,In_459);
xor U258 (N_258,In_296,In_1620);
and U259 (N_259,In_1307,In_601);
and U260 (N_260,In_190,In_1064);
nand U261 (N_261,In_1518,N_119);
nor U262 (N_262,In_1314,In_766);
or U263 (N_263,In_570,In_288);
nand U264 (N_264,In_1547,In_868);
xor U265 (N_265,In_1267,In_925);
xnor U266 (N_266,In_397,In_77);
nand U267 (N_267,In_671,In_498);
and U268 (N_268,In_1380,In_257);
and U269 (N_269,In_273,In_1612);
or U270 (N_270,In_86,In_208);
nand U271 (N_271,N_140,In_1079);
nand U272 (N_272,In_1230,In_101);
nor U273 (N_273,In_1286,In_1863);
and U274 (N_274,In_1364,In_1683);
nor U275 (N_275,In_460,In_1899);
xnor U276 (N_276,In_1458,In_1932);
xnor U277 (N_277,In_994,In_514);
nor U278 (N_278,In_1962,In_283);
xor U279 (N_279,In_907,In_1266);
nand U280 (N_280,In_995,In_1203);
nor U281 (N_281,In_136,In_1090);
xor U282 (N_282,In_431,N_60);
nand U283 (N_283,In_1461,N_72);
nand U284 (N_284,In_1919,In_1340);
nor U285 (N_285,In_261,N_44);
xnor U286 (N_286,In_1023,In_504);
nand U287 (N_287,In_799,In_1053);
xnor U288 (N_288,N_77,In_338);
and U289 (N_289,In_410,In_480);
or U290 (N_290,In_1848,N_53);
nand U291 (N_291,In_687,In_849);
nor U292 (N_292,In_376,In_1515);
nor U293 (N_293,In_1468,In_723);
nand U294 (N_294,In_148,In_1401);
nor U295 (N_295,In_1665,In_861);
nor U296 (N_296,In_325,In_1063);
or U297 (N_297,In_243,N_47);
or U298 (N_298,In_839,In_1769);
nand U299 (N_299,N_158,In_387);
xor U300 (N_300,In_1336,In_1339);
or U301 (N_301,In_1174,In_1579);
nor U302 (N_302,In_420,In_449);
nand U303 (N_303,In_119,In_1355);
or U304 (N_304,N_102,In_1604);
nand U305 (N_305,In_1976,In_1634);
nor U306 (N_306,In_1361,In_591);
nor U307 (N_307,In_1170,In_803);
and U308 (N_308,In_1996,In_862);
and U309 (N_309,In_496,In_454);
xnor U310 (N_310,In_1971,In_531);
nor U311 (N_311,N_149,In_106);
xnor U312 (N_312,In_1693,In_408);
or U313 (N_313,In_131,In_1677);
and U314 (N_314,In_306,In_1394);
nor U315 (N_315,In_1215,In_579);
xor U316 (N_316,In_1346,In_568);
nand U317 (N_317,In_113,In_108);
nor U318 (N_318,In_1123,In_782);
or U319 (N_319,In_1055,In_1805);
nand U320 (N_320,In_547,N_69);
nor U321 (N_321,In_1337,In_1373);
nand U322 (N_322,In_1918,In_501);
nor U323 (N_323,In_1663,N_180);
nor U324 (N_324,In_1312,In_731);
nand U325 (N_325,In_495,In_198);
and U326 (N_326,In_1268,In_404);
or U327 (N_327,N_33,In_1472);
xnor U328 (N_328,In_1478,N_281);
nor U329 (N_329,In_430,In_18);
and U330 (N_330,N_75,In_1537);
xnor U331 (N_331,In_147,In_263);
nand U332 (N_332,In_97,N_252);
and U333 (N_333,In_517,In_1849);
nand U334 (N_334,In_676,In_977);
nor U335 (N_335,In_1507,N_20);
or U336 (N_336,In_1358,N_95);
and U337 (N_337,In_1360,In_20);
or U338 (N_338,N_233,In_132);
nand U339 (N_339,In_1703,In_1288);
and U340 (N_340,In_1353,In_919);
nand U341 (N_341,In_824,N_273);
xor U342 (N_342,In_1202,N_112);
nand U343 (N_343,In_718,N_279);
and U344 (N_344,In_14,In_1093);
or U345 (N_345,In_1795,In_275);
nor U346 (N_346,In_634,In_967);
or U347 (N_347,In_1892,In_660);
nand U348 (N_348,In_369,In_906);
and U349 (N_349,In_1581,In_1354);
and U350 (N_350,In_792,In_1037);
nor U351 (N_351,In_937,In_935);
xor U352 (N_352,In_801,In_1178);
and U353 (N_353,In_1749,In_1614);
and U354 (N_354,In_1842,In_508);
xnor U355 (N_355,In_1292,In_1785);
or U356 (N_356,In_1033,N_295);
xnor U357 (N_357,In_1965,In_1672);
nor U358 (N_358,N_64,In_1655);
nand U359 (N_359,In_562,N_203);
and U360 (N_360,In_158,In_1327);
or U361 (N_361,In_806,In_446);
and U362 (N_362,In_624,In_1776);
and U363 (N_363,N_280,In_1809);
nor U364 (N_364,In_928,In_425);
or U365 (N_365,In_1299,In_1362);
xnor U366 (N_366,N_287,In_751);
or U367 (N_367,In_88,In_1482);
or U368 (N_368,N_284,In_710);
and U369 (N_369,In_134,In_440);
or U370 (N_370,In_419,In_463);
nand U371 (N_371,In_1232,In_5);
xnor U372 (N_372,In_1880,N_176);
nand U373 (N_373,In_1320,In_1902);
xnor U374 (N_374,In_1957,In_1613);
xnor U375 (N_375,In_985,In_987);
or U376 (N_376,In_681,In_1516);
nand U377 (N_377,In_1102,In_71);
nand U378 (N_378,In_51,In_1713);
or U379 (N_379,In_185,In_83);
or U380 (N_380,In_1527,In_1206);
nand U381 (N_381,N_266,In_197);
xnor U382 (N_382,In_484,In_932);
xor U383 (N_383,In_403,In_1106);
nor U384 (N_384,In_1759,In_1089);
or U385 (N_385,In_1750,In_1019);
xor U386 (N_386,In_1444,N_197);
nand U387 (N_387,N_236,In_1982);
or U388 (N_388,In_1676,In_1061);
xnor U389 (N_389,In_1107,In_1311);
nor U390 (N_390,In_1569,In_1711);
xnor U391 (N_391,In_1407,N_134);
and U392 (N_392,In_1610,In_871);
nor U393 (N_393,In_1696,In_1097);
and U394 (N_394,In_226,In_518);
xnor U395 (N_395,In_927,In_1605);
xnor U396 (N_396,N_288,In_571);
xor U397 (N_397,In_31,In_863);
or U398 (N_398,In_1187,In_853);
or U399 (N_399,In_1234,In_950);
xnor U400 (N_400,In_1691,In_175);
xor U401 (N_401,In_663,In_282);
nand U402 (N_402,In_1014,In_1281);
nor U403 (N_403,In_1639,In_187);
or U404 (N_404,In_511,In_1116);
xnor U405 (N_405,In_37,In_700);
nor U406 (N_406,In_984,N_182);
nand U407 (N_407,In_989,In_1626);
nand U408 (N_408,In_561,In_465);
and U409 (N_409,N_146,In_12);
nand U410 (N_410,In_576,In_618);
nand U411 (N_411,In_140,In_351);
nor U412 (N_412,In_65,In_339);
and U413 (N_413,In_367,In_61);
nor U414 (N_414,In_418,N_93);
and U415 (N_415,In_1082,In_1190);
or U416 (N_416,In_1451,In_1772);
or U417 (N_417,In_1006,In_830);
nor U418 (N_418,In_846,N_250);
nand U419 (N_419,In_712,In_711);
or U420 (N_420,In_1695,In_1113);
nand U421 (N_421,N_306,In_1716);
xor U422 (N_422,In_1422,In_585);
or U423 (N_423,In_593,In_172);
nor U424 (N_424,In_885,In_1667);
nor U425 (N_425,In_1498,N_315);
and U426 (N_426,In_1410,In_606);
and U427 (N_427,N_239,In_1443);
and U428 (N_428,In_466,In_1959);
nand U429 (N_429,In_610,In_1374);
or U430 (N_430,In_1788,In_844);
nand U431 (N_431,In_1603,N_56);
nor U432 (N_432,In_75,In_1977);
or U433 (N_433,In_1035,N_272);
and U434 (N_434,In_688,N_70);
nor U435 (N_435,In_734,N_277);
xnor U436 (N_436,In_714,In_1245);
nand U437 (N_437,N_201,In_584);
nor U438 (N_438,In_1792,In_411);
nor U439 (N_439,In_344,In_329);
or U440 (N_440,N_114,In_319);
nand U441 (N_441,In_391,In_1179);
and U442 (N_442,In_16,In_1176);
nand U443 (N_443,In_373,In_1191);
xor U444 (N_444,N_225,In_1908);
or U445 (N_445,In_1517,In_422);
and U446 (N_446,In_1156,In_1381);
xor U447 (N_447,In_632,In_923);
or U448 (N_448,In_1240,In_1270);
xnor U449 (N_449,In_1730,N_37);
nand U450 (N_450,In_814,In_205);
nor U451 (N_451,In_829,In_1508);
xor U452 (N_452,In_1559,N_184);
or U453 (N_453,In_85,In_1905);
xnor U454 (N_454,In_1829,In_235);
or U455 (N_455,In_1745,In_1924);
and U456 (N_456,In_982,In_1007);
and U457 (N_457,In_1819,In_706);
or U458 (N_458,In_635,In_1546);
xnor U459 (N_459,In_486,In_349);
nor U460 (N_460,In_620,N_129);
nor U461 (N_461,N_145,In_355);
xor U462 (N_462,In_1861,In_777);
and U463 (N_463,In_697,In_902);
and U464 (N_464,In_23,In_532);
nor U465 (N_465,N_49,In_1348);
or U466 (N_466,In_455,In_1878);
and U467 (N_467,In_432,N_85);
or U468 (N_468,In_835,In_477);
nand U469 (N_469,N_300,In_1085);
xnor U470 (N_470,In_1565,N_282);
and U471 (N_471,In_742,In_948);
nor U472 (N_472,In_1105,N_274);
xor U473 (N_473,In_1778,In_978);
nor U474 (N_474,In_1433,In_251);
nand U475 (N_475,In_1347,In_590);
nand U476 (N_476,In_1806,In_520);
or U477 (N_477,In_1632,In_1117);
nand U478 (N_478,In_1552,In_1678);
or U479 (N_479,In_95,N_251);
and U480 (N_480,N_175,In_146);
and U481 (N_481,In_1328,In_1143);
xnor U482 (N_482,N_229,In_1026);
nand U483 (N_483,N_84,In_1133);
or U484 (N_484,In_1894,N_10);
nand U485 (N_485,N_360,In_768);
nand U486 (N_486,In_1144,In_1675);
and U487 (N_487,N_177,In_1198);
or U488 (N_488,In_896,N_245);
nand U489 (N_489,In_974,N_291);
xnor U490 (N_490,In_1009,In_1434);
and U491 (N_491,In_1627,In_1385);
nand U492 (N_492,In_488,In_13);
nor U493 (N_493,In_1200,In_1185);
or U494 (N_494,In_1964,In_1661);
nor U495 (N_495,In_1566,In_87);
and U496 (N_496,N_211,In_1315);
nand U497 (N_497,In_778,In_318);
nor U498 (N_498,In_1210,In_1648);
nand U499 (N_499,In_1057,N_130);
nor U500 (N_500,N_101,N_165);
or U501 (N_501,In_1521,In_1244);
nor U502 (N_502,In_372,In_1519);
and U503 (N_503,In_245,In_933);
and U504 (N_504,In_1986,In_364);
nand U505 (N_505,N_383,N_443);
nor U506 (N_506,N_445,In_828);
and U507 (N_507,N_327,In_581);
nand U508 (N_508,N_262,In_753);
nand U509 (N_509,In_541,In_242);
nand U510 (N_510,In_204,In_1050);
or U511 (N_511,In_151,In_1756);
nor U512 (N_512,In_1774,In_203);
xnor U513 (N_513,N_345,In_949);
and U514 (N_514,In_1305,N_185);
nand U515 (N_515,N_392,In_1845);
or U516 (N_516,N_439,In_1099);
xnor U517 (N_517,In_353,N_246);
nor U518 (N_518,In_648,In_303);
xor U519 (N_519,N_178,In_1607);
and U520 (N_520,In_595,In_565);
nand U521 (N_521,In_1970,In_1134);
nand U522 (N_522,In_825,N_54);
xor U523 (N_523,N_369,In_945);
xnor U524 (N_524,In_168,N_209);
nand U525 (N_525,In_608,In_1321);
nor U526 (N_526,In_1188,N_390);
or U527 (N_527,N_207,N_405);
or U528 (N_528,In_1368,N_326);
nor U529 (N_529,In_628,N_347);
and U530 (N_530,N_278,In_1442);
xor U531 (N_531,In_244,N_472);
nand U532 (N_532,N_415,In_966);
and U533 (N_533,In_1161,In_1370);
nand U534 (N_534,In_1120,In_1933);
nor U535 (N_535,In_1956,N_309);
nand U536 (N_536,In_1704,In_732);
nor U537 (N_537,In_1807,In_1553);
xnor U538 (N_538,In_441,In_1039);
or U539 (N_539,In_1490,In_647);
xnor U540 (N_540,In_301,In_467);
nand U541 (N_541,In_237,N_191);
or U542 (N_542,In_448,N_9);
or U543 (N_543,N_330,In_1590);
xor U544 (N_544,In_1457,In_1196);
or U545 (N_545,N_73,In_1509);
nand U546 (N_546,In_1383,In_1121);
and U547 (N_547,In_666,In_1473);
or U548 (N_548,In_1707,In_1870);
or U549 (N_549,N_192,In_1969);
xnor U550 (N_550,N_431,In_142);
nand U551 (N_551,In_366,In_1981);
nand U552 (N_552,In_1862,N_14);
nand U553 (N_553,In_1545,N_364);
nor U554 (N_554,In_100,In_1137);
or U555 (N_555,In_1650,In_464);
and U556 (N_556,In_554,In_137);
or U557 (N_557,In_627,In_437);
nand U558 (N_558,N_408,In_1388);
nor U559 (N_559,In_1207,In_903);
and U560 (N_560,In_1955,In_672);
nand U561 (N_561,In_1242,In_1925);
nand U562 (N_562,In_1502,N_428);
xnor U563 (N_563,In_642,In_1637);
nor U564 (N_564,In_1356,In_415);
and U565 (N_565,N_45,N_6);
nor U566 (N_566,In_1067,In_240);
nand U567 (N_567,In_589,N_63);
nor U568 (N_568,N_74,In_1746);
nor U569 (N_569,In_1463,In_1735);
nand U570 (N_570,N_321,In_1733);
and U571 (N_571,N_232,In_873);
and U572 (N_572,In_1261,N_409);
and U573 (N_573,In_623,In_880);
nand U574 (N_574,N_235,N_386);
nor U575 (N_575,In_946,In_809);
nor U576 (N_576,In_111,In_116);
nand U577 (N_577,N_438,In_1301);
or U578 (N_578,In_682,N_152);
and U579 (N_579,In_258,In_659);
and U580 (N_580,In_1585,N_179);
or U581 (N_581,N_324,In_69);
nand U582 (N_582,In_1051,N_459);
xnor U583 (N_583,In_1853,N_442);
xnor U584 (N_584,In_57,N_356);
xnor U585 (N_585,N_110,N_237);
nor U586 (N_586,N_318,In_1763);
nand U587 (N_587,In_1087,In_1523);
nor U588 (N_588,N_153,In_1233);
xor U589 (N_589,N_22,In_1762);
nor U590 (N_590,In_1405,In_726);
or U591 (N_591,N_91,In_670);
nand U592 (N_592,In_1727,In_1225);
nor U593 (N_593,N_258,In_549);
or U594 (N_594,N_55,N_410);
nand U595 (N_595,In_969,N_449);
nor U596 (N_596,N_370,In_646);
xor U597 (N_597,In_819,In_817);
and U598 (N_598,In_961,In_1411);
nor U599 (N_599,In_1712,In_1436);
nand U600 (N_600,In_1437,In_1115);
xnor U601 (N_601,N_329,In_1263);
and U602 (N_602,In_1075,In_1999);
xnor U603 (N_603,In_662,N_354);
nand U604 (N_604,In_35,In_730);
xor U605 (N_605,N_170,In_963);
nand U606 (N_606,N_425,In_1450);
or U607 (N_607,In_207,In_1462);
and U608 (N_608,In_1002,In_1549);
xnor U609 (N_609,In_21,In_1582);
nand U610 (N_610,In_1972,In_1148);
xor U611 (N_611,In_1158,N_308);
xor U612 (N_612,N_379,N_34);
nand U613 (N_613,N_1,In_1852);
nand U614 (N_614,In_1415,N_275);
and U615 (N_615,N_59,N_419);
or U616 (N_616,In_1114,N_357);
and U617 (N_617,In_395,In_1783);
and U618 (N_618,In_1946,In_1859);
and U619 (N_619,In_442,In_1495);
nand U620 (N_620,In_1332,In_1029);
nor U621 (N_621,N_264,N_240);
or U622 (N_622,In_598,In_692);
xor U623 (N_623,N_263,In_574);
nand U624 (N_624,In_334,In_1086);
nand U625 (N_625,In_1611,In_913);
and U626 (N_626,N_388,In_728);
or U627 (N_627,In_1576,N_384);
or U628 (N_628,In_834,In_1291);
nand U629 (N_629,In_545,N_121);
xor U630 (N_630,In_785,In_1330);
xnor U631 (N_631,N_372,In_556);
and U632 (N_632,N_249,In_1885);
or U633 (N_633,In_1335,In_1997);
nor U634 (N_634,In_332,In_970);
and U635 (N_635,N_98,In_380);
or U636 (N_636,In_1420,In_1917);
or U637 (N_637,In_864,In_333);
or U638 (N_638,In_1855,In_1555);
or U639 (N_639,In_1379,N_462);
or U640 (N_640,In_337,In_1258);
or U641 (N_641,N_181,In_772);
nand U642 (N_642,N_501,In_1396);
or U643 (N_643,In_1427,In_971);
nand U644 (N_644,In_225,In_725);
nor U645 (N_645,N_137,In_262);
or U646 (N_646,N_292,In_274);
and U647 (N_647,N_188,In_983);
nand U648 (N_648,In_1980,In_1944);
or U649 (N_649,N_285,N_342);
or U650 (N_650,In_658,N_103);
xnor U651 (N_651,In_1149,N_639);
and U652 (N_652,N_526,In_1284);
nor U653 (N_653,In_888,N_618);
nand U654 (N_654,In_831,N_424);
nand U655 (N_655,N_381,N_463);
xnor U656 (N_656,In_1920,N_555);
nor U657 (N_657,In_1954,N_310);
and U658 (N_658,N_603,N_214);
nor U659 (N_659,In_1402,In_1491);
nor U660 (N_660,In_1341,N_362);
and U661 (N_661,N_633,In_346);
nand U662 (N_662,In_575,N_602);
nor U663 (N_663,In_1505,In_1850);
nand U664 (N_664,In_631,In_926);
and U665 (N_665,In_1949,In_722);
nand U666 (N_666,In_793,In_1352);
or U667 (N_667,N_118,N_508);
or U668 (N_668,In_1973,In_1391);
xnor U669 (N_669,N_626,In_1539);
or U670 (N_670,In_1342,N_476);
nor U671 (N_671,In_272,In_1048);
or U672 (N_672,N_113,In_826);
nand U673 (N_673,N_551,In_860);
xor U674 (N_674,N_148,In_1801);
nand U675 (N_675,N_189,N_485);
xnor U676 (N_676,In_1851,In_248);
and U677 (N_677,In_1467,In_1001);
nor U678 (N_678,In_1791,In_1813);
or U679 (N_679,In_794,N_216);
xnor U680 (N_680,In_236,In_1211);
and U681 (N_681,N_563,N_365);
xnor U682 (N_682,In_537,In_220);
xor U683 (N_683,In_1432,In_471);
and U684 (N_684,In_1212,In_1858);
or U685 (N_685,In_1345,In_66);
or U686 (N_686,N_414,N_195);
or U687 (N_687,In_1003,In_123);
and U688 (N_688,N_550,N_406);
nand U689 (N_689,In_758,In_914);
and U690 (N_690,In_58,N_349);
or U691 (N_691,In_476,In_1474);
nand U692 (N_692,N_541,In_270);
nor U693 (N_693,In_675,In_1077);
and U694 (N_694,N_494,In_754);
xnor U695 (N_695,In_1439,N_7);
and U696 (N_696,N_46,In_645);
xor U697 (N_697,In_456,N_483);
nand U698 (N_698,In_1882,N_186);
and U699 (N_699,In_1609,In_120);
and U700 (N_700,In_1622,In_1583);
xor U701 (N_701,In_298,In_1589);
and U702 (N_702,In_1419,N_173);
xor U703 (N_703,In_739,N_228);
and U704 (N_704,N_554,N_221);
and U705 (N_705,N_99,N_446);
or U706 (N_706,In_957,N_556);
nand U707 (N_707,N_88,In_1616);
xnor U708 (N_708,In_1510,In_1264);
and U709 (N_709,In_398,N_125);
nand U710 (N_710,In_1201,In_1409);
and U711 (N_711,In_1817,In_1044);
or U712 (N_712,N_334,In_1931);
xor U713 (N_713,In_135,In_1540);
or U714 (N_714,In_821,In_219);
nand U715 (N_715,In_256,In_104);
nand U716 (N_716,In_1963,In_1282);
and U717 (N_717,In_703,In_278);
or U718 (N_718,In_478,In_1897);
nor U719 (N_719,In_879,In_1484);
xnor U720 (N_720,N_257,In_975);
nor U721 (N_721,In_1890,In_1558);
nand U722 (N_722,In_908,N_171);
or U723 (N_723,In_705,N_465);
nor U724 (N_724,In_1794,N_536);
nand U725 (N_725,In_383,In_588);
nand U726 (N_726,In_322,In_493);
or U727 (N_727,N_202,In_859);
xnor U728 (N_728,In_1732,In_850);
and U729 (N_729,In_898,N_30);
nor U730 (N_730,N_562,N_572);
nor U731 (N_731,N_621,In_1773);
or U732 (N_732,N_163,N_546);
nand U733 (N_733,In_1866,N_468);
or U734 (N_734,N_154,In_1272);
nand U735 (N_735,In_115,In_1888);
or U736 (N_736,In_1702,In_1464);
xnor U737 (N_737,N_493,In_1426);
nor U738 (N_738,In_500,N_391);
xor U739 (N_739,In_1818,In_105);
xnor U740 (N_740,In_1367,N_374);
or U741 (N_741,In_797,N_27);
nor U742 (N_742,N_590,In_653);
or U743 (N_743,In_1629,In_1739);
nor U744 (N_744,In_1091,In_577);
nand U745 (N_745,In_1943,In_461);
nand U746 (N_746,N_517,In_1122);
xor U747 (N_747,In_227,N_15);
nand U748 (N_748,In_7,In_1790);
or U749 (N_749,In_1929,In_1758);
or U750 (N_750,N_519,In_354);
or U751 (N_751,In_1293,N_487);
xnor U752 (N_752,In_1780,In_1624);
or U753 (N_753,In_414,In_1728);
and U754 (N_754,In_232,In_1038);
nand U755 (N_755,In_833,N_123);
and U756 (N_756,N_448,In_1548);
and U757 (N_757,In_1204,In_745);
or U758 (N_758,In_1349,In_1159);
or U759 (N_759,In_702,N_21);
and U760 (N_760,In_637,N_537);
or U761 (N_761,N_17,N_283);
and U762 (N_762,In_1318,N_566);
and U763 (N_763,In_1587,N_255);
nor U764 (N_764,In_229,N_135);
or U765 (N_765,N_40,In_1714);
or U766 (N_766,In_453,In_181);
and U767 (N_767,In_1715,In_560);
nand U768 (N_768,N_452,N_608);
or U769 (N_769,N_515,In_139);
xnor U770 (N_770,In_643,In_1706);
or U771 (N_771,In_1334,In_1775);
xor U772 (N_772,N_16,In_1684);
and U773 (N_773,In_567,N_322);
and U774 (N_774,In_917,In_1592);
or U775 (N_775,N_339,In_1856);
or U776 (N_776,In_1653,In_1633);
or U777 (N_777,In_1904,In_960);
nand U778 (N_778,In_167,In_786);
or U779 (N_779,N_488,In_552);
nor U780 (N_780,N_553,In_434);
nand U781 (N_781,In_1418,In_299);
or U782 (N_782,In_1054,In_1323);
or U783 (N_783,In_405,In_693);
or U784 (N_784,N_402,N_385);
and U785 (N_785,N_270,In_1493);
or U786 (N_786,In_1313,In_201);
and U787 (N_787,N_377,In_1618);
nor U788 (N_788,N_294,In_807);
xnor U789 (N_789,In_155,N_509);
and U790 (N_790,N_124,In_838);
or U791 (N_791,In_639,N_611);
nor U792 (N_792,In_972,N_133);
xnor U793 (N_793,N_254,N_591);
nor U794 (N_794,In_412,In_1979);
nand U795 (N_795,N_531,In_630);
nand U796 (N_796,In_1167,In_993);
nand U797 (N_797,In_1231,In_289);
nor U798 (N_798,In_304,N_100);
nor U799 (N_799,In_76,N_586);
or U800 (N_800,In_877,N_625);
or U801 (N_801,N_606,In_291);
or U802 (N_802,In_1098,In_690);
and U803 (N_803,In_41,N_187);
xnor U804 (N_804,N_157,In_1837);
or U805 (N_805,N_336,N_243);
xor U806 (N_806,N_527,In_40);
or U807 (N_807,In_1459,In_1199);
xnor U808 (N_808,In_323,In_462);
or U809 (N_809,In_655,N_490);
nand U810 (N_810,In_1088,N_686);
nand U811 (N_811,N_687,N_290);
nand U812 (N_812,N_248,In_36);
nand U813 (N_813,In_1195,In_1155);
xnor U814 (N_814,In_62,In_481);
nor U815 (N_815,N_784,N_412);
xnor U816 (N_816,In_389,In_1224);
nor U817 (N_817,N_455,N_786);
nor U818 (N_818,N_363,N_492);
nand U819 (N_819,N_713,In_920);
or U820 (N_820,In_563,N_299);
xor U821 (N_821,In_1251,In_209);
and U822 (N_822,In_1671,In_52);
or U823 (N_823,N_394,N_650);
or U824 (N_824,N_719,In_1488);
nor U825 (N_825,N_204,N_783);
nand U826 (N_826,N_547,N_529);
xor U827 (N_827,In_239,In_959);
or U828 (N_828,In_1013,N_65);
nor U829 (N_829,N_645,N_267);
nand U830 (N_830,In_955,N_644);
xnor U831 (N_831,N_92,In_1824);
or U832 (N_832,In_114,In_607);
nand U833 (N_833,In_1243,In_650);
and U834 (N_834,N_785,N_599);
nor U835 (N_835,N_760,N_624);
and U836 (N_836,In_362,In_1995);
xor U837 (N_837,In_228,N_36);
and U838 (N_838,N_538,N_115);
nand U839 (N_839,In_911,In_1597);
or U840 (N_840,N_593,In_170);
xnor U841 (N_841,N_677,In_327);
nand U842 (N_842,In_1222,In_761);
nor U843 (N_843,In_1296,In_1496);
xor U844 (N_844,In_1721,In_1682);
or U845 (N_845,In_1172,N_471);
nand U846 (N_846,In_1512,N_510);
nand U847 (N_847,In_1297,N_222);
or U848 (N_848,In_1911,N_588);
or U849 (N_849,N_241,N_710);
xnor U850 (N_850,In_285,In_715);
nor U851 (N_851,In_409,In_685);
nor U852 (N_852,N_435,In_233);
or U853 (N_853,In_328,In_1635);
or U854 (N_854,In_1827,In_1227);
and U855 (N_855,N_499,In_174);
nand U856 (N_856,In_740,N_104);
and U857 (N_857,N_641,In_1221);
and U858 (N_858,In_163,In_1657);
and U859 (N_859,In_1316,N_393);
xor U860 (N_860,N_174,In_719);
nand U861 (N_861,N_558,N_97);
nand U862 (N_862,In_1404,In_1446);
nand U863 (N_863,In_46,N_549);
nand U864 (N_864,N_500,In_1047);
xor U865 (N_865,In_1278,In_808);
and U866 (N_866,In_159,N_109);
xor U867 (N_867,In_90,N_5);
or U868 (N_868,N_316,N_736);
nor U869 (N_869,N_643,In_1398);
xnor U870 (N_870,In_96,N_495);
and U871 (N_871,In_668,In_324);
nor U872 (N_872,In_141,N_271);
xnor U873 (N_873,N_344,In_1615);
and U874 (N_874,In_770,In_539);
nand U875 (N_875,In_1095,In_1453);
and U876 (N_876,N_717,In_883);
xnor U877 (N_877,In_1743,N_589);
or U878 (N_878,In_1857,N_706);
or U879 (N_879,N_647,N_720);
xor U880 (N_880,In_901,In_109);
nand U881 (N_881,N_668,In_50);
xnor U882 (N_882,In_629,In_1140);
or U883 (N_883,N_496,In_1823);
nand U884 (N_884,N_627,In_1990);
nand U885 (N_885,N_569,N_323);
nand U886 (N_886,In_429,In_1985);
nor U887 (N_887,In_176,In_1359);
or U888 (N_888,N_585,In_891);
or U889 (N_889,In_357,N_768);
nand U890 (N_890,N_26,In_216);
xor U891 (N_891,N_696,In_1812);
or U892 (N_892,In_470,In_1036);
nor U893 (N_893,In_1747,In_930);
nand U894 (N_894,In_1071,N_744);
nor U895 (N_895,N_256,N_505);
xor U896 (N_896,N_387,In_1967);
nor U897 (N_897,N_320,In_445);
nand U898 (N_898,N_293,In_45);
or U899 (N_899,In_680,N_375);
or U900 (N_900,In_613,In_1065);
or U901 (N_901,In_1760,N_543);
nor U902 (N_902,In_126,In_779);
or U903 (N_903,N_213,In_1664);
nor U904 (N_904,N_771,N_711);
xnor U905 (N_905,In_1514,In_1889);
or U906 (N_906,N_155,In_49);
xor U907 (N_907,In_1425,N_530);
xnor U908 (N_908,N_514,N_682);
xor U909 (N_909,In_1435,N_791);
xnor U910 (N_910,N_507,In_1277);
or U911 (N_911,N_367,N_681);
or U912 (N_912,N_351,In_1351);
or U913 (N_913,In_1363,In_1742);
or U914 (N_914,N_670,In_1525);
xor U915 (N_915,N_521,In_1073);
or U916 (N_916,In_1860,N_503);
or U917 (N_917,In_749,N_142);
nand U918 (N_918,N_131,N_359);
and U919 (N_919,N_688,In_1322);
nor U920 (N_920,In_295,In_336);
or U921 (N_921,In_1588,N_787);
and U922 (N_922,N_763,In_874);
and U923 (N_923,In_1477,N_141);
nand U924 (N_924,In_1810,In_836);
xor U925 (N_925,In_1621,N_429);
or U926 (N_926,N_217,N_502);
nand U927 (N_927,N_548,In_1018);
xor U928 (N_928,In_1934,In_378);
or U929 (N_929,N_622,N_470);
xor U930 (N_930,In_1907,N_654);
and U931 (N_931,In_1871,N_355);
xnor U932 (N_932,In_890,In_815);
nor U933 (N_933,N_567,In_1875);
nor U934 (N_934,In_156,In_1068);
or U935 (N_935,In_192,N_413);
xnor U936 (N_936,In_1781,N_473);
nor U937 (N_937,N_136,N_231);
or U938 (N_938,N_631,N_87);
or U939 (N_939,In_678,N_312);
nand U940 (N_940,In_1486,N_702);
xor U941 (N_941,N_122,In_1534);
or U942 (N_942,In_1256,In_280);
and U943 (N_943,N_71,In_858);
nor U944 (N_944,N_143,In_1423);
xor U945 (N_945,In_1469,N_401);
and U946 (N_946,N_373,In_1042);
or U947 (N_947,N_313,In_1660);
nor U948 (N_948,N_685,N_683);
nor U949 (N_949,In_352,N_695);
nand U950 (N_950,In_736,N_160);
nand U951 (N_951,In_218,In_832);
or U952 (N_952,In_1782,N_436);
nor U953 (N_953,In_64,N_658);
and U954 (N_954,N_166,In_1466);
nor U955 (N_955,In_1080,In_1386);
xnor U956 (N_956,In_343,N_504);
xor U957 (N_957,In_1403,In_1303);
or U958 (N_958,N_466,In_897);
nand U959 (N_959,In_15,N_724);
nand U960 (N_960,N_437,In_756);
and U961 (N_961,In_762,N_646);
xnor U962 (N_962,N_814,N_581);
nor U963 (N_963,N_398,N_789);
nor U964 (N_964,In_1656,In_1076);
nor U965 (N_965,In_1839,N_523);
nor U966 (N_966,N_120,In_143);
nor U967 (N_967,N_610,In_1834);
nor U968 (N_968,In_1365,N_151);
nand U969 (N_969,N_954,N_38);
or U970 (N_970,In_1729,N_94);
and U971 (N_971,In_939,In_307);
and U972 (N_972,N_926,In_1751);
or U973 (N_973,N_848,N_220);
nor U974 (N_974,In_1893,In_1575);
and U975 (N_975,In_311,N_167);
nand U976 (N_976,In_524,N_664);
or U977 (N_977,In_154,In_986);
xnor U978 (N_978,N_640,N_782);
nand U979 (N_979,In_1554,In_527);
xor U980 (N_980,N_798,In_424);
xor U981 (N_981,In_59,N_892);
or U982 (N_982,N_845,N_605);
or U983 (N_983,N_756,N_755);
nor U984 (N_984,In_269,N_440);
and U985 (N_985,N_172,N_651);
nand U986 (N_986,In_516,In_1654);
and U987 (N_987,N_630,In_127);
or U988 (N_988,In_769,In_166);
nor U989 (N_989,N_335,N_108);
nand U990 (N_990,In_382,In_566);
or U991 (N_991,N_307,N_801);
xnor U992 (N_992,N_479,N_396);
nand U993 (N_993,In_934,N_657);
xnor U994 (N_994,N_434,N_303);
nand U995 (N_995,In_68,In_1928);
nand U996 (N_996,In_1606,N_361);
nand U997 (N_997,N_758,In_33);
nand U998 (N_998,In_1413,In_1249);
xor U999 (N_999,In_1560,N_656);
xnor U1000 (N_1000,N_12,In_1066);
nand U1001 (N_1001,In_1193,In_1738);
nor U1002 (N_1002,In_1454,In_1252);
nor U1003 (N_1003,In_1511,In_882);
nand U1004 (N_1004,In_535,In_515);
or U1005 (N_1005,N_609,In_1142);
and U1006 (N_1006,N_498,In_1598);
nor U1007 (N_1007,In_1679,N_797);
or U1008 (N_1008,N_648,In_1371);
and U1009 (N_1009,In_614,In_47);
and U1010 (N_1010,In_1455,In_1376);
xor U1011 (N_1011,In_1777,In_1279);
nand U1012 (N_1012,N_447,N_126);
or U1013 (N_1013,N_331,In_1992);
xor U1014 (N_1014,In_1989,In_1295);
nand U1015 (N_1015,N_882,In_1329);
or U1016 (N_1016,N_722,N_659);
or U1017 (N_1017,N_261,In_173);
nor U1018 (N_1018,N_745,N_319);
nor U1019 (N_1019,In_195,In_1030);
nand U1020 (N_1020,N_917,In_67);
nand U1021 (N_1021,N_869,N_592);
nor U1022 (N_1022,In_212,In_543);
nand U1023 (N_1023,N_302,N_353);
nor U1024 (N_1024,In_1698,In_160);
and U1025 (N_1025,N_901,N_259);
nand U1026 (N_1026,N_52,N_247);
and U1027 (N_1027,In_596,N_934);
nand U1028 (N_1028,N_959,N_403);
nor U1029 (N_1029,In_1154,N_574);
nand U1030 (N_1030,In_153,N_417);
nand U1031 (N_1031,N_366,N_524);
nor U1032 (N_1032,In_765,N_219);
nand U1033 (N_1033,In_1687,In_335);
or U1034 (N_1034,N_484,N_927);
nand U1035 (N_1035,In_447,In_129);
and U1036 (N_1036,N_169,N_407);
or U1037 (N_1037,N_450,N_311);
xor U1038 (N_1038,N_675,In_773);
xor U1039 (N_1039,N_715,N_25);
nor U1040 (N_1040,N_738,In_474);
and U1041 (N_1041,N_804,In_997);
and U1042 (N_1042,In_1058,In_1799);
nand U1043 (N_1043,N_737,In_193);
and U1044 (N_1044,In_1011,N_423);
nor U1045 (N_1045,In_392,In_1529);
nor U1046 (N_1046,N_705,In_102);
xor U1047 (N_1047,In_394,In_1052);
nand U1048 (N_1048,In_1910,In_1501);
nor U1049 (N_1049,N_460,In_1836);
nor U1050 (N_1050,N_795,In_780);
nand U1051 (N_1051,In_1414,In_791);
nand U1052 (N_1052,In_1843,N_422);
or U1053 (N_1053,N_718,In_1162);
xor U1054 (N_1054,N_79,N_595);
nand U1055 (N_1055,In_316,N_477);
xnor U1056 (N_1056,N_853,In_1004);
nor U1057 (N_1057,In_472,In_247);
nand U1058 (N_1058,In_1045,N_692);
nor U1059 (N_1059,In_215,In_674);
and U1060 (N_1060,N_777,In_3);
and U1061 (N_1061,In_1194,N_741);
xnor U1062 (N_1062,In_529,In_1596);
nor U1063 (N_1063,In_103,In_951);
nor U1064 (N_1064,In_497,In_716);
and U1065 (N_1065,In_843,In_1489);
and U1066 (N_1066,In_654,N_728);
nor U1067 (N_1067,In_542,In_1736);
and U1068 (N_1068,N_676,In_958);
nor U1069 (N_1069,N_159,In_300);
xnor U1070 (N_1070,N_680,N_11);
nand U1071 (N_1071,N_921,N_380);
or U1072 (N_1072,In_525,In_98);
and U1073 (N_1073,In_1906,N_652);
and U1074 (N_1074,N_400,N_616);
and U1075 (N_1075,N_577,In_1497);
nand U1076 (N_1076,In_1017,In_186);
and U1077 (N_1077,In_1947,N_632);
nor U1078 (N_1078,N_874,In_390);
nor U1079 (N_1079,N_458,In_1838);
nand U1080 (N_1080,In_1372,N_480);
nor U1081 (N_1081,N_456,N_729);
and U1082 (N_1082,N_164,N_649);
and U1083 (N_1083,In_1708,In_594);
nor U1084 (N_1084,N_570,N_301);
and U1085 (N_1085,N_489,N_857);
nor U1086 (N_1086,N_317,N_426);
xor U1087 (N_1087,In_469,N_860);
nand U1088 (N_1088,N_847,N_619);
and U1089 (N_1089,In_1874,N_790);
or U1090 (N_1090,N_224,In_214);
or U1091 (N_1091,In_1685,N_337);
or U1092 (N_1092,N_843,N_205);
nor U1093 (N_1093,In_79,In_182);
nand U1094 (N_1094,In_981,In_32);
nor U1095 (N_1095,N_582,N_371);
or U1096 (N_1096,N_887,N_451);
nand U1097 (N_1097,N_427,In_1602);
nand U1098 (N_1098,N_839,N_947);
nand U1099 (N_1099,In_1471,In_1757);
and U1100 (N_1100,In_42,In_1987);
and U1101 (N_1101,N_432,N_837);
or U1102 (N_1102,N_942,In_1886);
or U1103 (N_1103,In_1016,In_330);
or U1104 (N_1104,N_338,N_520);
or U1105 (N_1105,In_1557,N_761);
nor U1106 (N_1106,In_1101,N_821);
nand U1107 (N_1107,N_297,In_1139);
xnor U1108 (N_1108,N_861,N_557);
xor U1109 (N_1109,In_1652,N_749);
nand U1110 (N_1110,In_1417,In_178);
nor U1111 (N_1111,In_1731,In_302);
xnor U1112 (N_1112,In_375,N_899);
or U1113 (N_1113,In_1465,In_1357);
and U1114 (N_1114,In_202,N_828);
nor U1115 (N_1115,N_855,In_99);
nand U1116 (N_1116,N_842,N_560);
or U1117 (N_1117,N_568,N_348);
nand U1118 (N_1118,In_60,N_834);
nand U1119 (N_1119,N_807,In_1815);
nand U1120 (N_1120,In_840,N_865);
and U1121 (N_1121,In_1912,N_704);
nor U1122 (N_1122,N_826,In_28);
or U1123 (N_1123,N_889,In_1840);
and U1124 (N_1124,In_747,N_199);
nand U1125 (N_1125,N_754,N_888);
and U1126 (N_1126,In_1387,N_920);
and U1127 (N_1127,In_439,N_296);
and U1128 (N_1128,N_1071,In_443);
and U1129 (N_1129,In_255,In_238);
or U1130 (N_1130,N_1049,In_1689);
and U1131 (N_1131,In_224,N_932);
nand U1132 (N_1132,In_1551,In_633);
or U1133 (N_1133,In_1530,In_599);
and U1134 (N_1134,N_1074,N_571);
xor U1135 (N_1135,N_678,In_1968);
or U1136 (N_1136,N_852,In_1238);
nand U1137 (N_1137,In_721,N_62);
nand U1138 (N_1138,In_22,In_1481);
or U1139 (N_1139,N_1033,In_152);
nor U1140 (N_1140,N_827,N_168);
xor U1141 (N_1141,In_669,In_915);
nand U1142 (N_1142,N_1022,In_1124);
nor U1143 (N_1143,In_1709,N_573);
nor U1144 (N_1144,N_565,N_700);
xor U1145 (N_1145,N_957,In_1828);
nand U1146 (N_1146,In_1841,N_776);
and U1147 (N_1147,N_516,In_1217);
nand U1148 (N_1148,N_1048,In_1128);
and U1149 (N_1149,In_1438,N_111);
nand U1150 (N_1150,In_1571,In_118);
and U1151 (N_1151,In_1903,N_914);
nor U1152 (N_1152,In_673,In_616);
and U1153 (N_1153,In_641,N_817);
nor U1154 (N_1154,N_575,In_1412);
and U1155 (N_1155,In_401,In_1723);
xor U1156 (N_1156,N_227,In_942);
xor U1157 (N_1157,N_269,N_667);
or U1158 (N_1158,N_982,N_697);
nor U1159 (N_1159,N_642,N_350);
or U1160 (N_1160,N_1064,N_880);
nand U1161 (N_1161,N_89,N_535);
and U1162 (N_1162,In_1670,In_1993);
or U1163 (N_1163,N_1113,In_1666);
or U1164 (N_1164,N_1039,N_420);
nor U1165 (N_1165,N_699,N_389);
and U1166 (N_1166,N_1059,N_304);
and U1167 (N_1167,N_482,In_84);
nor U1168 (N_1168,N_730,In_649);
nand U1169 (N_1169,N_835,In_1369);
xnor U1170 (N_1170,In_851,N_1011);
nor U1171 (N_1171,N_884,In_1094);
and U1172 (N_1172,In_1914,N_1092);
nor U1173 (N_1173,N_902,N_802);
nand U1174 (N_1174,In_1513,N_870);
nor U1175 (N_1175,In_784,In_551);
and U1176 (N_1176,N_1017,In_1975);
and U1177 (N_1177,N_878,N_868);
xor U1178 (N_1178,N_328,N_872);
and U1179 (N_1179,N_1101,N_128);
nand U1180 (N_1180,N_1023,N_1055);
nand U1181 (N_1181,N_533,In_1503);
nand U1182 (N_1182,N_905,N_368);
and U1183 (N_1183,In_287,N_769);
and U1184 (N_1184,In_1699,N_475);
or U1185 (N_1185,N_977,In_1802);
and U1186 (N_1186,In_1164,N_1093);
nand U1187 (N_1187,In_130,N_981);
and U1188 (N_1188,N_544,In_112);
or U1189 (N_1189,N_81,N_915);
or U1190 (N_1190,N_962,In_1659);
or U1191 (N_1191,In_1520,In_1259);
and U1192 (N_1192,In_1237,In_1069);
xor U1193 (N_1193,In_489,In_1631);
and U1194 (N_1194,N_579,N_352);
and U1195 (N_1195,N_739,N_1070);
or U1196 (N_1196,N_1056,N_960);
and U1197 (N_1197,N_596,N_638);
or U1198 (N_1198,N_1079,N_486);
or U1199 (N_1199,In_1248,In_893);
nand U1200 (N_1200,In_1138,N_382);
or U1201 (N_1201,N_1116,N_881);
xnor U1202 (N_1202,N_689,In_1260);
and U1203 (N_1203,In_1793,N_1081);
xnor U1204 (N_1204,N_1086,N_346);
or U1205 (N_1205,N_956,In_1830);
or U1206 (N_1206,N_911,In_622);
or U1207 (N_1207,N_951,In_1814);
or U1208 (N_1208,N_1082,N_669);
or U1209 (N_1209,N_223,N_800);
or U1210 (N_1210,In_1181,In_1111);
or U1211 (N_1211,N_1041,N_1063);
and U1212 (N_1212,N_1094,N_1030);
nor U1213 (N_1213,In_1236,N_1003);
nor U1214 (N_1214,N_862,In_340);
or U1215 (N_1215,In_1229,N_743);
nand U1216 (N_1216,In_1923,N_945);
or U1217 (N_1217,N_773,N_815);
or U1218 (N_1218,N_753,N_467);
xor U1219 (N_1219,N_762,N_1095);
nor U1220 (N_1220,In_707,In_795);
nor U1221 (N_1221,N_193,N_971);
nor U1222 (N_1222,N_694,In_281);
nor U1223 (N_1223,N_684,N_497);
xor U1224 (N_1224,N_858,N_1024);
nand U1225 (N_1225,In_221,N_859);
nand U1226 (N_1226,N_1100,N_1062);
xor U1227 (N_1227,N_1083,In_717);
and U1228 (N_1228,N_1040,In_1499);
nand U1229 (N_1229,In_161,N_474);
xor U1230 (N_1230,In_1717,In_1584);
nor U1231 (N_1231,N_820,N_765);
xnor U1232 (N_1232,N_96,N_832);
xnor U1233 (N_1233,N_742,In_1197);
xor U1234 (N_1234,In_1104,In_870);
nand U1235 (N_1235,N_325,N_732);
nor U1236 (N_1236,N_979,In_1280);
xor U1237 (N_1237,N_162,In_626);
nor U1238 (N_1238,N_253,N_721);
or U1239 (N_1239,N_788,N_86);
xnor U1240 (N_1240,N_823,N_879);
or U1241 (N_1241,N_844,N_18);
nor U1242 (N_1242,N_830,N_701);
nand U1243 (N_1243,N_810,N_919);
and U1244 (N_1244,N_660,N_150);
xor U1245 (N_1245,N_1072,N_513);
nor U1246 (N_1246,N_863,In_1638);
or U1247 (N_1247,In_347,N_1034);
and U1248 (N_1248,In_211,In_485);
and U1249 (N_1249,In_1580,In_1891);
and U1250 (N_1250,N_907,In_912);
nand U1251 (N_1251,In_314,N_716);
or U1252 (N_1252,In_259,In_277);
or U1253 (N_1253,N_539,In_1216);
and U1254 (N_1254,N_298,N_1012);
and U1255 (N_1255,N_1118,N_933);
nand U1256 (N_1256,In_165,N_923);
nor U1257 (N_1257,N_663,N_876);
or U1258 (N_1258,In_1881,N_909);
or U1259 (N_1259,In_1630,In_1218);
nand U1260 (N_1260,N_925,N_799);
or U1261 (N_1261,N_600,N_208);
nand U1262 (N_1262,N_464,N_867);
xor U1263 (N_1263,N_1117,N_397);
nor U1264 (N_1264,N_42,In_698);
and U1265 (N_1265,N_1104,In_1983);
and U1266 (N_1266,In_943,In_1440);
or U1267 (N_1267,N_803,N_1112);
xor U1268 (N_1268,N_39,N_286);
or U1269 (N_1269,N_774,In_1262);
nor U1270 (N_1270,N_430,N_963);
xor U1271 (N_1271,N_812,N_156);
xnor U1272 (N_1272,In_1150,In_1668);
xor U1273 (N_1273,N_824,N_949);
and U1274 (N_1274,N_779,N_238);
xor U1275 (N_1275,N_747,N_144);
nor U1276 (N_1276,N_988,N_866);
or U1277 (N_1277,In_804,N_378);
or U1278 (N_1278,In_1562,N_506);
xnor U1279 (N_1279,In_133,In_1470);
xnor U1280 (N_1280,N_849,N_672);
nor U1281 (N_1281,N_871,N_598);
nand U1282 (N_1282,In_827,N_734);
or U1283 (N_1283,In_30,N_1001);
or U1284 (N_1284,N_604,N_825);
nand U1285 (N_1285,N_980,N_260);
and U1286 (N_1286,N_1019,In_572);
nand U1287 (N_1287,In_910,In_876);
xor U1288 (N_1288,In_1269,In_1395);
nand U1289 (N_1289,N_13,In_661);
and U1290 (N_1290,N_1029,In_55);
nand U1291 (N_1291,In_1223,N_890);
and U1292 (N_1292,N_1179,N_1027);
nor U1293 (N_1293,N_1258,In_1921);
nor U1294 (N_1294,N_196,N_1152);
or U1295 (N_1295,N_61,N_1234);
and U1296 (N_1296,N_1203,In_704);
nand U1297 (N_1297,N_19,In_750);
nor U1298 (N_1298,In_796,In_1542);
nand U1299 (N_1299,In_558,N_614);
and U1300 (N_1300,N_607,N_161);
and U1301 (N_1301,N_943,N_775);
nand U1302 (N_1302,N_481,N_1066);
nand U1303 (N_1303,N_1025,N_634);
and U1304 (N_1304,N_958,In_1049);
or U1305 (N_1305,N_1107,N_772);
or U1306 (N_1306,In_1811,N_1127);
xnor U1307 (N_1307,N_1123,In_709);
or U1308 (N_1308,N_1140,N_561);
nand U1309 (N_1309,In_523,N_511);
or U1310 (N_1310,N_816,N_912);
or U1311 (N_1311,N_1243,N_200);
and U1312 (N_1312,N_276,N_985);
or U1313 (N_1313,In_125,N_1216);
xnor U1314 (N_1314,In_1074,In_848);
nand U1315 (N_1315,N_967,N_829);
or U1316 (N_1316,In_1175,N_1111);
or U1317 (N_1317,N_822,In_1205);
nand U1318 (N_1318,N_1211,N_1241);
nor U1319 (N_1319,N_811,In_1526);
nor U1320 (N_1320,N_1195,N_757);
and U1321 (N_1321,In_617,N_206);
nor U1322 (N_1322,In_1393,N_534);
and U1323 (N_1323,N_444,In_1570);
nor U1324 (N_1324,N_404,N_265);
nor U1325 (N_1325,In_1384,N_613);
and U1326 (N_1326,In_213,N_1150);
nor U1327 (N_1327,N_215,N_1173);
nand U1328 (N_1328,N_1166,N_139);
xnor U1329 (N_1329,N_1139,N_1075);
or U1330 (N_1330,In_1642,N_594);
xnor U1331 (N_1331,In_359,N_1067);
and U1332 (N_1332,In_536,N_731);
and U1333 (N_1333,N_831,N_1273);
nand U1334 (N_1334,N_1035,In_388);
nor U1335 (N_1335,In_611,In_265);
nor U1336 (N_1336,N_3,In_789);
nand U1337 (N_1337,N_117,In_73);
nand U1338 (N_1338,N_1202,N_1212);
xor U1339 (N_1339,N_453,N_418);
or U1340 (N_1340,N_1162,N_751);
or U1341 (N_1341,N_999,N_1115);
nor U1342 (N_1342,N_1247,In_1998);
nand U1343 (N_1343,In_1522,N_972);
nor U1344 (N_1344,N_522,In_1214);
and U1345 (N_1345,N_1044,N_903);
nand U1346 (N_1346,In_813,N_1047);
and U1347 (N_1347,N_32,N_76);
and U1348 (N_1348,N_767,In_1271);
and U1349 (N_1349,N_1016,In_124);
nor U1350 (N_1350,In_805,In_1697);
or U1351 (N_1351,N_978,N_1114);
nor U1352 (N_1352,N_1190,N_780);
nor U1353 (N_1353,N_1271,N_1076);
xor U1354 (N_1354,N_1102,N_127);
or U1355 (N_1355,N_940,N_1200);
and U1356 (N_1356,In_358,In_1062);
and U1357 (N_1357,N_836,N_908);
or U1358 (N_1358,In_956,N_1168);
nor U1359 (N_1359,In_56,N_78);
xnor U1360 (N_1360,N_896,N_1009);
or U1361 (N_1361,N_1148,In_952);
or U1362 (N_1362,N_948,N_792);
xnor U1363 (N_1363,N_970,N_1182);
or U1364 (N_1364,N_1224,N_1028);
xnor U1365 (N_1365,N_712,In_150);
nor U1366 (N_1366,In_1186,N_1000);
and U1367 (N_1367,In_521,N_1194);
nand U1368 (N_1368,N_1218,N_1244);
xnor U1369 (N_1369,N_138,N_1225);
nand U1370 (N_1370,N_1109,In_249);
nand U1371 (N_1371,N_709,In_1253);
nand U1372 (N_1372,N_1060,N_1133);
xnor U1373 (N_1373,In_1324,In_436);
xnor U1374 (N_1374,N_1215,N_875);
or U1375 (N_1375,N_1155,In_1690);
and U1376 (N_1376,N_1005,N_1014);
or U1377 (N_1377,N_1099,In_889);
xor U1378 (N_1378,In_954,N_491);
or U1379 (N_1379,N_234,N_1161);
nor U1380 (N_1380,In_738,In_884);
xnor U1381 (N_1381,N_399,N_210);
nor U1382 (N_1382,In_1145,N_1185);
and U1383 (N_1383,N_1233,N_1253);
and U1384 (N_1384,N_1259,In_310);
nor U1385 (N_1385,N_961,N_564);
xor U1386 (N_1386,In_94,In_1239);
nor U1387 (N_1387,N_518,N_1121);
and U1388 (N_1388,N_1054,In_1083);
nand U1389 (N_1389,In_188,In_857);
nor U1390 (N_1390,N_242,In_696);
and U1391 (N_1391,N_636,N_1138);
xor U1392 (N_1392,N_976,N_726);
nand U1393 (N_1393,N_1106,In_787);
nor U1394 (N_1394,In_555,N_1164);
xor U1395 (N_1395,In_1789,N_629);
nor U1396 (N_1396,N_796,In_6);
or U1397 (N_1397,N_268,N_1010);
nand U1398 (N_1398,N_1045,N_1231);
nor U1399 (N_1399,N_673,N_29);
nand U1400 (N_1400,N_733,N_991);
xor U1401 (N_1401,N_1251,In_918);
and U1402 (N_1402,N_1143,N_343);
nor U1403 (N_1403,In_266,N_1057);
or U1404 (N_1404,N_1052,N_906);
xnor U1405 (N_1405,N_1085,N_1220);
or U1406 (N_1406,In_746,N_1183);
nor U1407 (N_1407,N_924,In_1276);
nand U1408 (N_1408,In_665,In_924);
or U1409 (N_1409,N_708,In_592);
nor U1410 (N_1410,N_1219,N_540);
and U1411 (N_1411,N_900,N_528);
nand U1412 (N_1412,In_1960,N_289);
xnor U1413 (N_1413,N_194,N_1252);
nor U1414 (N_1414,In_1681,N_1134);
nand U1415 (N_1415,N_1242,N_1153);
and U1416 (N_1416,In_1595,N_457);
nor U1417 (N_1417,N_1223,In_1031);
nor U1418 (N_1418,N_584,In_1563);
nand U1419 (N_1419,N_1222,N_51);
and U1420 (N_1420,In_1808,N_1269);
nor U1421 (N_1421,N_838,N_395);
nor U1422 (N_1422,In_1382,In_1887);
nor U1423 (N_1423,N_1263,N_1230);
xnor U1424 (N_1424,In_1936,In_528);
and U1425 (N_1425,N_1108,In_1865);
nor U1426 (N_1426,N_965,N_714);
nand U1427 (N_1427,N_1004,N_989);
xnor U1428 (N_1428,In_1599,In_1247);
and U1429 (N_1429,N_1128,N_1037);
nor U1430 (N_1430,N_1105,N_809);
or U1431 (N_1431,N_740,In_1421);
xnor U1432 (N_1432,In_664,N_1165);
nor U1433 (N_1433,N_1237,N_1204);
xor U1434 (N_1434,N_930,In_1832);
xor U1435 (N_1435,N_376,N_1221);
or U1436 (N_1436,N_1261,N_105);
and U1437 (N_1437,N_218,N_938);
or U1438 (N_1438,N_735,N_992);
and U1439 (N_1439,N_1192,N_1068);
or U1440 (N_1440,In_1152,In_371);
xnor U1441 (N_1441,N_1283,N_1331);
nand U1442 (N_1442,N_1330,N_1136);
nor U1443 (N_1443,N_1386,N_1188);
and U1444 (N_1444,In_973,N_1350);
and U1445 (N_1445,N_1098,N_1207);
nor U1446 (N_1446,N_993,In_905);
nand U1447 (N_1447,N_1051,N_1199);
and U1448 (N_1448,N_615,N_226);
xnor U1449 (N_1449,In_292,In_1129);
or U1450 (N_1450,In_964,N_1322);
and U1451 (N_1451,N_1077,N_1318);
xnor U1452 (N_1452,In_1662,N_1174);
nor U1453 (N_1453,N_1103,N_1154);
nor U1454 (N_1454,N_805,N_746);
xnor U1455 (N_1455,N_1335,N_748);
nor U1456 (N_1456,N_1434,N_552);
or U1457 (N_1457,N_1413,N_1310);
and U1458 (N_1458,N_935,N_1205);
nand U1459 (N_1459,In_1766,N_1329);
or U1460 (N_1460,N_916,N_937);
xor U1461 (N_1461,N_1389,N_1349);
xnor U1462 (N_1462,In_331,N_1270);
nand U1463 (N_1463,N_894,N_1297);
nand U1464 (N_1464,N_662,N_1429);
or U1465 (N_1465,N_1398,N_806);
and U1466 (N_1466,N_601,N_1015);
xnor U1467 (N_1467,N_1018,N_1416);
and U1468 (N_1468,In_1319,N_1409);
nor U1469 (N_1469,N_1364,In_1309);
or U1470 (N_1470,N_1248,N_1124);
and U1471 (N_1471,N_984,N_1120);
or U1472 (N_1472,N_1306,N_1132);
nand U1473 (N_1473,N_1374,In_540);
nand U1474 (N_1474,N_1193,N_690);
nor U1475 (N_1475,N_1013,N_1341);
nor U1476 (N_1476,In_1909,N_132);
nand U1477 (N_1477,In_1524,N_1189);
and U1478 (N_1478,N_1296,N_1299);
or U1479 (N_1479,N_1284,In_1941);
nor U1480 (N_1480,In_482,In_1141);
and U1481 (N_1481,N_1361,N_1303);
xor U1482 (N_1482,N_1319,N_341);
nor U1483 (N_1483,N_1317,N_1352);
nor U1484 (N_1484,In_1310,N_1245);
nor U1485 (N_1485,In_1768,N_1332);
xnor U1486 (N_1486,N_1320,In_1822);
nand U1487 (N_1487,In_180,In_548);
nor U1488 (N_1488,N_612,N_990);
and U1489 (N_1489,N_1314,N_1380);
nor U1490 (N_1490,N_587,N_1163);
nor U1491 (N_1491,N_1144,N_808);
nand U1492 (N_1492,N_1180,N_693);
nor U1493 (N_1493,In_1110,N_1122);
or U1494 (N_1494,In_241,N_1294);
and U1495 (N_1495,N_1399,N_1309);
and U1496 (N_1496,N_1379,N_1147);
nand U1497 (N_1497,N_1336,N_512);
or U1498 (N_1498,N_1042,N_1260);
nand U1499 (N_1499,In_121,N_67);
xor U1500 (N_1500,N_666,N_1226);
or U1501 (N_1501,N_1228,N_1184);
nand U1502 (N_1502,N_1240,N_1290);
or U1503 (N_1503,N_1146,In_757);
xor U1504 (N_1504,N_1333,N_1187);
or U1505 (N_1505,In_10,N_1227);
xor U1506 (N_1506,In_999,N_454);
nor U1507 (N_1507,N_1325,N_1394);
xor U1508 (N_1508,N_1279,N_1137);
or U1509 (N_1509,N_818,N_1403);
xnor U1510 (N_1510,N_1430,N_1435);
xnor U1511 (N_1511,In_183,N_1359);
or U1512 (N_1512,N_1401,N_1286);
nor U1513 (N_1513,N_212,N_1407);
or U1514 (N_1514,N_819,N_1427);
nor U1515 (N_1515,In_1953,N_1287);
xor U1516 (N_1516,N_441,In_82);
nand U1517 (N_1517,N_433,N_766);
nor U1518 (N_1518,N_8,N_617);
or U1519 (N_1519,N_1171,N_1311);
nor U1520 (N_1520,N_944,N_559);
nor U1521 (N_1521,N_1340,N_1363);
xnor U1522 (N_1522,N_1424,N_1312);
xnor U1523 (N_1523,N_987,N_1423);
nand U1524 (N_1524,In_320,N_891);
nand U1525 (N_1525,In_1937,N_1388);
nand U1526 (N_1526,N_1141,N_1372);
xnor U1527 (N_1527,N_1422,N_1091);
nor U1528 (N_1528,N_230,In_775);
nor U1529 (N_1529,N_1383,N_1327);
or U1530 (N_1530,N_1323,N_1238);
xnor U1531 (N_1531,N_1266,N_968);
xnor U1532 (N_1532,N_1419,N_1061);
or U1533 (N_1533,N_1175,N_1097);
nor U1534 (N_1534,N_1345,N_854);
or U1535 (N_1535,N_931,N_597);
and U1536 (N_1536,N_1315,N_545);
or U1537 (N_1537,In_1578,In_223);
and U1538 (N_1538,N_1366,N_90);
nand U1539 (N_1539,N_904,N_416);
nand U1540 (N_1540,N_1217,N_983);
xor U1541 (N_1541,N_1302,In_321);
nor U1542 (N_1542,In_210,N_995);
nand U1543 (N_1543,N_1291,N_1395);
nor U1544 (N_1544,N_1169,N_1334);
and U1545 (N_1545,N_1281,In_619);
or U1546 (N_1546,N_1381,N_580);
or U1547 (N_1547,In_1325,N_1343);
nor U1548 (N_1548,N_1382,N_939);
or U1549 (N_1549,N_929,N_1362);
xor U1550 (N_1550,N_723,N_1355);
nor U1551 (N_1551,N_1073,N_358);
or U1552 (N_1552,N_781,N_244);
and U1553 (N_1553,N_1026,N_1300);
or U1554 (N_1554,N_1096,N_1324);
nor U1555 (N_1555,In_1593,N_1378);
or U1556 (N_1556,N_1326,N_1257);
and U1557 (N_1557,N_1089,N_1370);
and U1558 (N_1558,N_478,N_1080);
nor U1559 (N_1559,In_1343,N_1006);
nand U1560 (N_1560,N_674,N_1348);
or U1561 (N_1561,N_1339,N_1256);
xnor U1562 (N_1562,N_1264,N_469);
nor U1563 (N_1563,In_771,N_1369);
nand U1564 (N_1564,N_851,N_1328);
xor U1565 (N_1565,N_1131,In_473);
or U1566 (N_1566,N_31,N_1020);
and U1567 (N_1567,In_1826,N_759);
nand U1568 (N_1568,N_1181,N_48);
xnor U1569 (N_1569,N_1142,In_1163);
and U1570 (N_1570,N_679,N_1313);
xor U1571 (N_1571,N_918,In_89);
and U1572 (N_1572,N_969,N_1254);
or U1573 (N_1573,N_994,N_1426);
or U1574 (N_1574,N_1126,N_1250);
or U1575 (N_1575,N_665,N_1400);
or U1576 (N_1576,N_1214,N_1125);
xnor U1577 (N_1577,N_1065,N_305);
nor U1578 (N_1578,In_720,In_74);
nor U1579 (N_1579,In_1306,N_1285);
or U1580 (N_1580,In_393,N_1373);
nor U1581 (N_1581,N_1288,N_576);
xor U1582 (N_1582,N_794,N_850);
nand U1583 (N_1583,N_461,In_1940);
nor U1584 (N_1584,In_691,N_1420);
and U1585 (N_1585,N_628,In_1020);
xnor U1586 (N_1586,In_1568,N_1084);
nand U1587 (N_1587,N_996,In_1688);
xnor U1588 (N_1588,In_1448,N_846);
xor U1589 (N_1589,N_68,N_1396);
or U1590 (N_1590,In_92,N_1268);
nor U1591 (N_1591,In_869,In_377);
nor U1592 (N_1592,N_1196,N_1408);
and U1593 (N_1593,N_1351,N_1439);
and U1594 (N_1594,N_1437,N_1008);
nand U1595 (N_1595,N_1255,N_1275);
nand U1596 (N_1596,In_783,N_1405);
nand U1597 (N_1597,N_57,N_1119);
and U1598 (N_1598,N_1415,N_1149);
nand U1599 (N_1599,N_190,N_1078);
nor U1600 (N_1600,N_966,N_116);
nor U1601 (N_1601,In_1485,N_1547);
nor U1602 (N_1602,N_1412,N_1496);
nor U1603 (N_1603,N_4,N_1458);
and U1604 (N_1604,N_1551,N_1523);
and U1605 (N_1605,N_1574,N_1446);
nand U1606 (N_1606,N_1178,N_411);
or U1607 (N_1607,N_1476,N_1546);
nor U1608 (N_1608,N_1356,N_1462);
nor U1609 (N_1609,N_1198,N_1562);
or U1610 (N_1610,N_1582,N_1544);
and U1611 (N_1611,N_1456,N_1573);
and U1612 (N_1612,N_1497,N_1489);
xnor U1613 (N_1613,N_1032,N_1043);
xor U1614 (N_1614,N_833,N_1347);
nor U1615 (N_1615,N_1490,N_1298);
or U1616 (N_1616,N_691,In_1958);
nand U1617 (N_1617,N_1229,N_1021);
xnor U1618 (N_1618,N_1110,N_1575);
and U1619 (N_1619,N_1512,N_770);
nor U1620 (N_1620,N_764,N_1090);
nor U1621 (N_1621,N_1552,In_1915);
or U1622 (N_1622,N_1464,N_1466);
and U1623 (N_1623,In_764,N_1528);
xnor U1624 (N_1624,In_546,N_1526);
nand U1625 (N_1625,N_1433,N_698);
xor U1626 (N_1626,N_583,N_1443);
nand U1627 (N_1627,N_1524,N_1537);
and U1628 (N_1628,N_1507,N_1553);
or U1629 (N_1629,In_1171,N_1410);
nand U1630 (N_1630,N_1565,N_1514);
or U1631 (N_1631,N_910,In_1333);
and U1632 (N_1632,N_1521,N_998);
xor U1633 (N_1633,In_979,In_149);
nor U1634 (N_1634,N_623,In_904);
and U1635 (N_1635,N_1088,In_1586);
nor U1636 (N_1636,N_1556,N_1440);
xnor U1637 (N_1637,N_936,In_1673);
nand U1638 (N_1638,N_885,N_1472);
and U1639 (N_1639,N_1555,N_1087);
xnor U1640 (N_1640,N_1534,N_1598);
nand U1641 (N_1641,N_1232,In_416);
nand U1642 (N_1642,N_1421,N_1338);
xnor U1643 (N_1643,N_1404,N_655);
or U1644 (N_1644,N_1246,N_1402);
nand U1645 (N_1645,In_1177,N_1589);
xor U1646 (N_1646,N_1566,In_1250);
nand U1647 (N_1647,N_1482,N_1493);
or U1648 (N_1648,N_1572,N_913);
nor U1649 (N_1649,N_1473,N_1516);
or U1650 (N_1650,N_1444,In_171);
nor U1651 (N_1651,N_1542,In_980);
xnor U1652 (N_1652,N_1567,N_1478);
and U1653 (N_1653,In_194,N_198);
or U1654 (N_1654,N_1485,N_727);
and U1655 (N_1655,In_421,N_1321);
and U1656 (N_1656,N_1540,N_1594);
nand U1657 (N_1657,N_1518,N_1499);
xor U1658 (N_1658,N_1491,N_1365);
or U1659 (N_1659,N_1586,N_973);
xnor U1660 (N_1660,N_1197,N_1170);
nand U1661 (N_1661,N_1129,N_1344);
or U1662 (N_1662,N_707,N_1517);
or U1663 (N_1663,N_1417,N_1494);
or U1664 (N_1664,N_183,In_1406);
and U1665 (N_1665,N_1058,N_1158);
and U1666 (N_1666,N_1236,In_1103);
nand U1667 (N_1667,N_1584,N_1577);
or U1668 (N_1668,N_1474,N_1451);
nand U1669 (N_1669,N_1465,N_1428);
or U1670 (N_1670,In_677,N_1590);
or U1671 (N_1671,N_1477,N_1530);
and U1672 (N_1672,In_1939,N_1277);
and U1673 (N_1673,N_1470,N_1487);
and U1674 (N_1674,N_1449,N_1593);
nor U1675 (N_1675,N_1511,N_1301);
nor U1676 (N_1676,N_1342,N_1130);
nand U1677 (N_1677,N_1550,N_1282);
and U1678 (N_1678,N_1368,N_1280);
and U1679 (N_1679,N_620,N_1535);
nor U1680 (N_1680,N_1460,N_1592);
nor U1681 (N_1681,N_1580,N_1506);
or U1682 (N_1682,N_314,N_1397);
and U1683 (N_1683,N_1543,N_1570);
xor U1684 (N_1684,N_1069,N_1249);
nor U1685 (N_1685,N_1046,N_1157);
nand U1686 (N_1686,In_1625,N_1591);
xor U1687 (N_1687,N_873,N_1167);
xor U1688 (N_1688,N_1559,N_898);
nor U1689 (N_1689,N_1448,N_578);
or U1690 (N_1690,In_1895,N_922);
and U1691 (N_1691,N_1436,In_348);
nor U1692 (N_1692,N_1414,N_1377);
nand U1693 (N_1693,In_1350,N_793);
nand U1694 (N_1694,N_1425,N_1469);
nor U1695 (N_1695,N_895,N_1201);
or U1696 (N_1696,In_1651,N_1527);
or U1697 (N_1697,N_1545,N_1276);
xnor U1698 (N_1698,N_1272,N_1510);
or U1699 (N_1699,N_1525,N_1548);
and U1700 (N_1700,N_1160,N_1159);
nor U1701 (N_1701,N_1564,N_671);
nor U1702 (N_1702,N_1191,N_332);
nand U1703 (N_1703,N_1036,N_1305);
nor U1704 (N_1704,N_1385,N_941);
or U1705 (N_1705,N_147,N_1515);
nand U1706 (N_1706,N_986,N_525);
xor U1707 (N_1707,N_1235,N_41);
or U1708 (N_1708,N_1053,N_1384);
nor U1709 (N_1709,In_1028,N_1007);
and U1710 (N_1710,N_778,N_1557);
nand U1711 (N_1711,N_813,N_928);
or U1712 (N_1712,N_974,N_1308);
nor U1713 (N_1713,N_1583,N_856);
nor U1714 (N_1714,N_1459,N_1354);
nand U1715 (N_1715,N_1453,N_1316);
nand U1716 (N_1716,In_1647,In_1649);
xor U1717 (N_1717,N_1538,N_1353);
xnor U1718 (N_1718,N_1569,In_1010);
xnor U1719 (N_1719,N_1587,N_1387);
nor U1720 (N_1720,N_1213,N_1346);
nor U1721 (N_1721,N_1596,N_883);
nand U1722 (N_1722,N_1457,N_1509);
nand U1723 (N_1723,N_1431,N_1452);
or U1724 (N_1724,N_1480,N_1442);
or U1725 (N_1725,N_1571,N_1393);
or U1726 (N_1726,N_1471,In_1873);
or U1727 (N_1727,N_107,N_1533);
or U1728 (N_1728,N_1145,N_1522);
or U1729 (N_1729,N_1337,N_1151);
or U1730 (N_1730,N_1209,N_1445);
nand U1731 (N_1731,N_1463,N_1467);
xor U1732 (N_1732,N_1597,N_1031);
and U1733 (N_1733,N_1292,N_1176);
and U1734 (N_1734,N_1560,N_1406);
nand U1735 (N_1735,In_1119,N_653);
xnor U1736 (N_1736,N_1038,N_1441);
nor U1737 (N_1737,N_1581,In_1032);
nor U1738 (N_1738,N_1488,N_1262);
or U1739 (N_1739,N_1520,N_635);
and U1740 (N_1740,N_725,N_1495);
nor U1741 (N_1741,In_312,N_1563);
xnor U1742 (N_1742,N_955,N_1513);
or U1743 (N_1743,N_1295,N_1293);
xor U1744 (N_1744,N_1418,N_893);
xnor U1745 (N_1745,N_1501,N_1475);
and U1746 (N_1746,N_1206,N_1519);
and U1747 (N_1747,N_997,N_1376);
and U1748 (N_1748,N_1578,N_1390);
or U1749 (N_1749,N_1438,N_897);
and U1750 (N_1750,N_750,N_1585);
and U1751 (N_1751,N_637,N_841);
or U1752 (N_1752,N_1172,N_1357);
nand U1753 (N_1753,N_703,In_1182);
xnor U1754 (N_1754,In_1209,N_1588);
or U1755 (N_1755,N_1504,N_340);
nand U1756 (N_1756,N_1289,N_1135);
nor U1757 (N_1757,N_1447,N_333);
or U1758 (N_1758,In_1535,N_1532);
or U1759 (N_1759,N_1508,N_1595);
nand U1760 (N_1760,N_1705,N_1745);
xnor U1761 (N_1761,N_1651,N_1604);
and U1762 (N_1762,In_1180,N_1643);
nor U1763 (N_1763,N_1708,N_1481);
nor U1764 (N_1764,N_1626,N_1721);
xor U1765 (N_1765,N_1568,N_1669);
nand U1766 (N_1766,N_1360,N_1050);
nand U1767 (N_1767,N_1502,N_1695);
xor U1768 (N_1768,N_1455,N_1265);
and U1769 (N_1769,N_1628,N_1741);
xor U1770 (N_1770,N_1358,N_1479);
xnor U1771 (N_1771,N_1600,N_1744);
xnor U1772 (N_1772,N_1713,In_11);
and U1773 (N_1773,N_964,N_1753);
and U1774 (N_1774,N_1645,N_1720);
xor U1775 (N_1775,N_1186,N_1612);
xor U1776 (N_1776,N_1274,N_1671);
xnor U1777 (N_1777,N_1724,N_1696);
xnor U1778 (N_1778,N_1716,In_1556);
and U1779 (N_1779,N_1682,N_1549);
nand U1780 (N_1780,N_1684,N_1662);
or U1781 (N_1781,N_1531,N_1714);
or U1782 (N_1782,N_1661,N_1608);
or U1783 (N_1783,N_1667,N_1576);
and U1784 (N_1784,N_1536,N_1685);
and U1785 (N_1785,N_1613,N_1649);
nor U1786 (N_1786,N_1638,N_1492);
xnor U1787 (N_1787,N_1625,N_1707);
xnor U1788 (N_1788,N_1450,N_1411);
xor U1789 (N_1789,N_1672,N_1629);
or U1790 (N_1790,N_1541,N_1689);
and U1791 (N_1791,In_1169,N_1632);
nor U1792 (N_1792,N_1751,N_1432);
nand U1793 (N_1793,N_1610,N_1391);
xor U1794 (N_1794,N_1644,N_1648);
nand U1795 (N_1795,N_1717,N_1620);
nand U1796 (N_1796,In_1796,N_1611);
or U1797 (N_1797,N_1752,N_1683);
nor U1798 (N_1798,N_1002,N_1601);
or U1799 (N_1799,N_1723,N_1609);
xor U1800 (N_1800,N_1691,N_1666);
and U1801 (N_1801,N_1500,N_421);
or U1802 (N_1802,N_1636,N_1746);
or U1803 (N_1803,In_350,N_1710);
or U1804 (N_1804,N_1554,N_1647);
nor U1805 (N_1805,N_752,N_1758);
or U1806 (N_1806,In_491,N_1665);
nor U1807 (N_1807,N_1267,N_1239);
nor U1808 (N_1808,N_1733,N_1698);
nor U1809 (N_1809,N_1693,N_1639);
or U1810 (N_1810,N_1726,N_1728);
nor U1811 (N_1811,N_1701,N_1634);
xor U1812 (N_1812,N_1679,N_1757);
and U1813 (N_1813,N_1755,N_1635);
nor U1814 (N_1814,N_1732,N_1619);
nor U1815 (N_1815,N_1740,N_1624);
xor U1816 (N_1816,N_1653,N_1622);
xor U1817 (N_1817,N_1738,N_1668);
nand U1818 (N_1818,N_1642,N_1686);
or U1819 (N_1819,N_1735,N_952);
or U1820 (N_1820,N_1709,N_1742);
nor U1821 (N_1821,N_1605,N_1539);
xnor U1822 (N_1822,N_840,N_1641);
nand U1823 (N_1823,N_1697,N_1688);
and U1824 (N_1824,N_1392,N_1748);
nor U1825 (N_1825,N_1371,N_1660);
and U1826 (N_1826,N_1676,N_1177);
or U1827 (N_1827,N_1617,N_1529);
nor U1828 (N_1828,N_1646,N_1503);
nand U1829 (N_1829,In_1771,N_886);
nor U1830 (N_1830,N_1498,N_1704);
nor U1831 (N_1831,N_1375,N_1703);
nand U1832 (N_1832,N_1678,N_1654);
xor U1833 (N_1833,N_1278,N_1307);
and U1834 (N_1834,N_950,N_1754);
or U1835 (N_1835,N_1579,N_1663);
nor U1836 (N_1836,N_1484,N_1674);
or U1837 (N_1837,N_1607,N_953);
nor U1838 (N_1838,N_975,N_1759);
nor U1839 (N_1839,N_946,N_864);
or U1840 (N_1840,N_1631,N_1743);
nand U1841 (N_1841,In_759,N_1750);
and U1842 (N_1842,N_1658,N_1561);
nand U1843 (N_1843,N_1731,N_1690);
nand U1844 (N_1844,N_532,N_1749);
xor U1845 (N_1845,N_1734,N_1680);
nor U1846 (N_1846,In_1600,N_1675);
xnor U1847 (N_1847,N_661,N_1711);
or U1848 (N_1848,N_1729,N_1461);
nand U1849 (N_1849,N_1656,N_1739);
nand U1850 (N_1850,N_1615,N_1616);
xnor U1851 (N_1851,N_1486,N_1681);
nand U1852 (N_1852,N_1670,N_542);
xor U1853 (N_1853,N_1702,N_1627);
nand U1854 (N_1854,In_1168,N_1483);
or U1855 (N_1855,N_1715,N_1208);
nor U1856 (N_1856,N_1673,N_1712);
and U1857 (N_1857,N_1621,N_1655);
or U1858 (N_1858,N_1210,N_1367);
nand U1859 (N_1859,N_1602,N_1304);
or U1860 (N_1860,N_1623,N_1454);
nor U1861 (N_1861,N_1505,N_1468);
or U1862 (N_1862,N_1614,N_1558);
xor U1863 (N_1863,N_1599,N_1725);
xnor U1864 (N_1864,N_1637,N_1722);
nor U1865 (N_1865,N_1718,N_1719);
xor U1866 (N_1866,N_877,N_1727);
nand U1867 (N_1867,N_1692,N_1677);
and U1868 (N_1868,N_1650,N_1606);
nand U1869 (N_1869,N_1706,N_1603);
nor U1870 (N_1870,N_1699,N_1657);
nor U1871 (N_1871,N_1756,N_1700);
and U1872 (N_1872,N_1630,N_1652);
xnor U1873 (N_1873,In_264,N_1687);
or U1874 (N_1874,In_1390,N_1747);
or U1875 (N_1875,N_1640,N_1736);
and U1876 (N_1876,N_1156,N_1664);
nor U1877 (N_1877,N_1694,N_1618);
xnor U1878 (N_1878,N_1659,N_1730);
nand U1879 (N_1879,N_1737,N_1633);
xor U1880 (N_1880,N_1576,N_1734);
xnor U1881 (N_1881,N_1617,N_1742);
nor U1882 (N_1882,N_1717,N_1755);
and U1883 (N_1883,N_1208,N_1610);
nand U1884 (N_1884,N_1719,N_1690);
nand U1885 (N_1885,N_1671,N_1634);
nor U1886 (N_1886,N_964,N_1484);
nand U1887 (N_1887,N_1727,N_1675);
nor U1888 (N_1888,N_752,N_1722);
or U1889 (N_1889,N_1632,N_1613);
nand U1890 (N_1890,N_542,N_1682);
and U1891 (N_1891,N_1733,N_1683);
nor U1892 (N_1892,N_1642,N_1741);
xor U1893 (N_1893,N_1599,N_1628);
or U1894 (N_1894,N_1690,N_1639);
nand U1895 (N_1895,N_1743,N_1706);
xor U1896 (N_1896,N_1360,N_1649);
xnor U1897 (N_1897,N_1239,N_1690);
or U1898 (N_1898,N_1682,N_1640);
nand U1899 (N_1899,N_1554,N_1655);
xor U1900 (N_1900,N_1720,N_1627);
xnor U1901 (N_1901,In_1556,N_1498);
and U1902 (N_1902,N_1625,N_1679);
nand U1903 (N_1903,N_1304,N_1657);
and U1904 (N_1904,N_1678,N_661);
nand U1905 (N_1905,N_1367,N_1623);
or U1906 (N_1906,N_1274,N_1698);
nor U1907 (N_1907,In_11,N_752);
xor U1908 (N_1908,N_1177,N_1708);
or U1909 (N_1909,N_1725,N_1692);
nand U1910 (N_1910,N_1690,N_1610);
nand U1911 (N_1911,N_1632,N_1719);
xor U1912 (N_1912,N_1745,N_1614);
or U1913 (N_1913,N_1617,N_1568);
and U1914 (N_1914,N_1743,N_1752);
and U1915 (N_1915,N_1623,N_1050);
or U1916 (N_1916,N_1375,N_1502);
nand U1917 (N_1917,N_1755,N_1732);
and U1918 (N_1918,N_1670,N_1610);
nor U1919 (N_1919,N_1729,N_1483);
xnor U1920 (N_1920,N_1857,N_1872);
nor U1921 (N_1921,N_1856,N_1869);
nand U1922 (N_1922,N_1794,N_1841);
and U1923 (N_1923,N_1848,N_1771);
or U1924 (N_1924,N_1793,N_1788);
and U1925 (N_1925,N_1785,N_1839);
and U1926 (N_1926,N_1823,N_1879);
or U1927 (N_1927,N_1835,N_1908);
and U1928 (N_1928,N_1799,N_1911);
or U1929 (N_1929,N_1797,N_1824);
nor U1930 (N_1930,N_1833,N_1874);
nand U1931 (N_1931,N_1814,N_1873);
nand U1932 (N_1932,N_1822,N_1766);
nor U1933 (N_1933,N_1884,N_1801);
nand U1934 (N_1934,N_1803,N_1825);
nor U1935 (N_1935,N_1912,N_1864);
or U1936 (N_1936,N_1890,N_1807);
and U1937 (N_1937,N_1805,N_1867);
nand U1938 (N_1938,N_1896,N_1855);
xor U1939 (N_1939,N_1767,N_1893);
nor U1940 (N_1940,N_1777,N_1909);
or U1941 (N_1941,N_1903,N_1838);
nor U1942 (N_1942,N_1892,N_1829);
nor U1943 (N_1943,N_1883,N_1882);
and U1944 (N_1944,N_1791,N_1795);
nand U1945 (N_1945,N_1876,N_1844);
or U1946 (N_1946,N_1810,N_1789);
xnor U1947 (N_1947,N_1804,N_1760);
nor U1948 (N_1948,N_1891,N_1796);
or U1949 (N_1949,N_1845,N_1820);
or U1950 (N_1950,N_1846,N_1917);
or U1951 (N_1951,N_1778,N_1769);
xnor U1952 (N_1952,N_1780,N_1905);
and U1953 (N_1953,N_1837,N_1898);
nor U1954 (N_1954,N_1853,N_1815);
xnor U1955 (N_1955,N_1836,N_1871);
nor U1956 (N_1956,N_1910,N_1821);
and U1957 (N_1957,N_1842,N_1907);
or U1958 (N_1958,N_1781,N_1826);
nand U1959 (N_1959,N_1786,N_1787);
and U1960 (N_1960,N_1861,N_1798);
and U1961 (N_1961,N_1875,N_1865);
xor U1962 (N_1962,N_1862,N_1850);
nor U1963 (N_1963,N_1851,N_1868);
nand U1964 (N_1964,N_1776,N_1915);
or U1965 (N_1965,N_1765,N_1854);
and U1966 (N_1966,N_1816,N_1881);
xor U1967 (N_1967,N_1809,N_1817);
or U1968 (N_1968,N_1919,N_1770);
nand U1969 (N_1969,N_1859,N_1904);
or U1970 (N_1970,N_1763,N_1774);
xnor U1971 (N_1971,N_1790,N_1779);
nor U1972 (N_1972,N_1843,N_1852);
nor U1973 (N_1973,N_1913,N_1813);
xor U1974 (N_1974,N_1831,N_1792);
xnor U1975 (N_1975,N_1768,N_1899);
nand U1976 (N_1976,N_1858,N_1783);
or U1977 (N_1977,N_1832,N_1818);
xor U1978 (N_1978,N_1811,N_1830);
xnor U1979 (N_1979,N_1885,N_1761);
nor U1980 (N_1980,N_1847,N_1772);
nor U1981 (N_1981,N_1888,N_1762);
nor U1982 (N_1982,N_1784,N_1802);
or U1983 (N_1983,N_1887,N_1916);
or U1984 (N_1984,N_1895,N_1886);
xnor U1985 (N_1985,N_1902,N_1800);
and U1986 (N_1986,N_1812,N_1863);
nor U1987 (N_1987,N_1827,N_1906);
or U1988 (N_1988,N_1877,N_1764);
nand U1989 (N_1989,N_1840,N_1773);
and U1990 (N_1990,N_1870,N_1828);
nor U1991 (N_1991,N_1914,N_1878);
nor U1992 (N_1992,N_1806,N_1866);
xor U1993 (N_1993,N_1849,N_1775);
xnor U1994 (N_1994,N_1897,N_1782);
or U1995 (N_1995,N_1860,N_1808);
or U1996 (N_1996,N_1889,N_1834);
and U1997 (N_1997,N_1900,N_1819);
and U1998 (N_1998,N_1894,N_1880);
or U1999 (N_1999,N_1901,N_1918);
nor U2000 (N_2000,N_1897,N_1912);
nand U2001 (N_2001,N_1807,N_1765);
xor U2002 (N_2002,N_1909,N_1908);
and U2003 (N_2003,N_1876,N_1879);
and U2004 (N_2004,N_1824,N_1903);
nand U2005 (N_2005,N_1835,N_1905);
xnor U2006 (N_2006,N_1888,N_1792);
or U2007 (N_2007,N_1770,N_1819);
nand U2008 (N_2008,N_1899,N_1817);
nor U2009 (N_2009,N_1912,N_1851);
nor U2010 (N_2010,N_1870,N_1833);
or U2011 (N_2011,N_1844,N_1888);
and U2012 (N_2012,N_1844,N_1828);
and U2013 (N_2013,N_1799,N_1772);
xnor U2014 (N_2014,N_1777,N_1839);
nor U2015 (N_2015,N_1763,N_1778);
and U2016 (N_2016,N_1878,N_1889);
xor U2017 (N_2017,N_1789,N_1791);
and U2018 (N_2018,N_1821,N_1890);
or U2019 (N_2019,N_1830,N_1860);
xor U2020 (N_2020,N_1789,N_1852);
and U2021 (N_2021,N_1774,N_1878);
xnor U2022 (N_2022,N_1762,N_1807);
nor U2023 (N_2023,N_1917,N_1828);
nand U2024 (N_2024,N_1765,N_1879);
or U2025 (N_2025,N_1840,N_1897);
or U2026 (N_2026,N_1815,N_1837);
nor U2027 (N_2027,N_1901,N_1796);
or U2028 (N_2028,N_1904,N_1856);
and U2029 (N_2029,N_1789,N_1826);
and U2030 (N_2030,N_1896,N_1788);
and U2031 (N_2031,N_1890,N_1811);
xor U2032 (N_2032,N_1890,N_1848);
nor U2033 (N_2033,N_1867,N_1883);
nand U2034 (N_2034,N_1847,N_1891);
or U2035 (N_2035,N_1781,N_1906);
xnor U2036 (N_2036,N_1915,N_1770);
and U2037 (N_2037,N_1794,N_1914);
and U2038 (N_2038,N_1830,N_1901);
nand U2039 (N_2039,N_1807,N_1826);
or U2040 (N_2040,N_1794,N_1793);
nor U2041 (N_2041,N_1825,N_1850);
nor U2042 (N_2042,N_1797,N_1871);
xnor U2043 (N_2043,N_1855,N_1830);
nor U2044 (N_2044,N_1772,N_1895);
xnor U2045 (N_2045,N_1780,N_1890);
nand U2046 (N_2046,N_1867,N_1816);
nor U2047 (N_2047,N_1862,N_1853);
or U2048 (N_2048,N_1859,N_1824);
or U2049 (N_2049,N_1779,N_1794);
or U2050 (N_2050,N_1845,N_1760);
and U2051 (N_2051,N_1837,N_1785);
xor U2052 (N_2052,N_1908,N_1863);
xor U2053 (N_2053,N_1836,N_1855);
nand U2054 (N_2054,N_1816,N_1774);
and U2055 (N_2055,N_1857,N_1778);
xnor U2056 (N_2056,N_1902,N_1782);
nand U2057 (N_2057,N_1882,N_1843);
or U2058 (N_2058,N_1896,N_1884);
nor U2059 (N_2059,N_1800,N_1869);
or U2060 (N_2060,N_1885,N_1895);
and U2061 (N_2061,N_1819,N_1777);
and U2062 (N_2062,N_1761,N_1819);
nand U2063 (N_2063,N_1762,N_1869);
nor U2064 (N_2064,N_1790,N_1864);
and U2065 (N_2065,N_1848,N_1891);
or U2066 (N_2066,N_1808,N_1789);
xor U2067 (N_2067,N_1855,N_1818);
xnor U2068 (N_2068,N_1861,N_1850);
nand U2069 (N_2069,N_1853,N_1800);
xor U2070 (N_2070,N_1782,N_1887);
nand U2071 (N_2071,N_1901,N_1890);
nand U2072 (N_2072,N_1807,N_1905);
and U2073 (N_2073,N_1855,N_1805);
and U2074 (N_2074,N_1821,N_1791);
nor U2075 (N_2075,N_1886,N_1877);
xnor U2076 (N_2076,N_1852,N_1854);
and U2077 (N_2077,N_1872,N_1784);
xnor U2078 (N_2078,N_1853,N_1811);
xor U2079 (N_2079,N_1780,N_1807);
nor U2080 (N_2080,N_2003,N_2077);
and U2081 (N_2081,N_2028,N_1966);
or U2082 (N_2082,N_1974,N_2038);
nor U2083 (N_2083,N_2070,N_2048);
or U2084 (N_2084,N_2044,N_1960);
nand U2085 (N_2085,N_2075,N_1964);
xnor U2086 (N_2086,N_2061,N_1950);
xor U2087 (N_2087,N_2043,N_1990);
xor U2088 (N_2088,N_1994,N_1979);
or U2089 (N_2089,N_2057,N_1940);
nand U2090 (N_2090,N_1962,N_1920);
xor U2091 (N_2091,N_1977,N_1930);
or U2092 (N_2092,N_1969,N_1929);
nor U2093 (N_2093,N_2035,N_2053);
and U2094 (N_2094,N_1923,N_1978);
xnor U2095 (N_2095,N_2022,N_2023);
and U2096 (N_2096,N_1944,N_1926);
nand U2097 (N_2097,N_2021,N_2059);
nor U2098 (N_2098,N_1982,N_2006);
and U2099 (N_2099,N_2064,N_1987);
nand U2100 (N_2100,N_1967,N_2014);
nor U2101 (N_2101,N_2025,N_2040);
and U2102 (N_2102,N_1942,N_1932);
nor U2103 (N_2103,N_1951,N_1989);
and U2104 (N_2104,N_1993,N_2076);
nand U2105 (N_2105,N_1980,N_1922);
xor U2106 (N_2106,N_2072,N_1968);
and U2107 (N_2107,N_2069,N_1965);
or U2108 (N_2108,N_2068,N_2041);
or U2109 (N_2109,N_2020,N_2037);
nor U2110 (N_2110,N_2055,N_1972);
and U2111 (N_2111,N_2009,N_2018);
nor U2112 (N_2112,N_1931,N_1996);
and U2113 (N_2113,N_2079,N_2010);
nand U2114 (N_2114,N_1957,N_2067);
nor U2115 (N_2115,N_2060,N_1935);
nand U2116 (N_2116,N_1986,N_1949);
or U2117 (N_2117,N_1981,N_1983);
or U2118 (N_2118,N_1921,N_2039);
nor U2119 (N_2119,N_1976,N_2031);
xor U2120 (N_2120,N_2046,N_1952);
or U2121 (N_2121,N_2030,N_2011);
or U2122 (N_2122,N_1998,N_1999);
nor U2123 (N_2123,N_1946,N_2002);
nor U2124 (N_2124,N_1934,N_1939);
or U2125 (N_2125,N_1936,N_2019);
or U2126 (N_2126,N_1937,N_2065);
nand U2127 (N_2127,N_1997,N_1988);
nand U2128 (N_2128,N_1933,N_2078);
xnor U2129 (N_2129,N_2005,N_1928);
or U2130 (N_2130,N_1948,N_1973);
xnor U2131 (N_2131,N_1953,N_2063);
xnor U2132 (N_2132,N_2047,N_1961);
or U2133 (N_2133,N_2062,N_2024);
nand U2134 (N_2134,N_2052,N_2029);
nand U2135 (N_2135,N_1958,N_2032);
nor U2136 (N_2136,N_2000,N_2026);
or U2137 (N_2137,N_2027,N_1970);
nand U2138 (N_2138,N_2001,N_2071);
and U2139 (N_2139,N_1963,N_2051);
nand U2140 (N_2140,N_2012,N_1945);
and U2141 (N_2141,N_1925,N_2066);
nand U2142 (N_2142,N_2050,N_2074);
xor U2143 (N_2143,N_2008,N_1943);
nor U2144 (N_2144,N_1924,N_1956);
nand U2145 (N_2145,N_1985,N_2016);
xor U2146 (N_2146,N_1991,N_1975);
nand U2147 (N_2147,N_1941,N_2007);
nor U2148 (N_2148,N_1959,N_1927);
xnor U2149 (N_2149,N_2036,N_2017);
or U2150 (N_2150,N_2056,N_2073);
nand U2151 (N_2151,N_2042,N_1955);
nor U2152 (N_2152,N_1954,N_1984);
xnor U2153 (N_2153,N_2004,N_2058);
nor U2154 (N_2154,N_1947,N_2013);
or U2155 (N_2155,N_2049,N_2054);
nand U2156 (N_2156,N_2033,N_2034);
and U2157 (N_2157,N_1938,N_1971);
nor U2158 (N_2158,N_1992,N_1995);
nor U2159 (N_2159,N_2045,N_2015);
or U2160 (N_2160,N_1959,N_2014);
and U2161 (N_2161,N_2026,N_1927);
and U2162 (N_2162,N_2019,N_2013);
nand U2163 (N_2163,N_1953,N_2043);
or U2164 (N_2164,N_2038,N_2047);
or U2165 (N_2165,N_1963,N_2030);
nand U2166 (N_2166,N_1963,N_1984);
and U2167 (N_2167,N_1967,N_2007);
or U2168 (N_2168,N_1997,N_1986);
xnor U2169 (N_2169,N_1992,N_2019);
xnor U2170 (N_2170,N_1954,N_2027);
xor U2171 (N_2171,N_1943,N_1997);
or U2172 (N_2172,N_2018,N_1922);
and U2173 (N_2173,N_1959,N_1989);
or U2174 (N_2174,N_2052,N_1935);
and U2175 (N_2175,N_1935,N_2023);
or U2176 (N_2176,N_1959,N_2066);
nand U2177 (N_2177,N_1979,N_2021);
nor U2178 (N_2178,N_2061,N_2000);
nand U2179 (N_2179,N_2040,N_2064);
and U2180 (N_2180,N_1983,N_1993);
nand U2181 (N_2181,N_1958,N_2010);
and U2182 (N_2182,N_2004,N_1995);
xor U2183 (N_2183,N_1973,N_1933);
nand U2184 (N_2184,N_2017,N_1986);
nor U2185 (N_2185,N_2079,N_2052);
or U2186 (N_2186,N_1996,N_1952);
xnor U2187 (N_2187,N_1933,N_2052);
nand U2188 (N_2188,N_1940,N_1937);
or U2189 (N_2189,N_1948,N_2071);
and U2190 (N_2190,N_2039,N_2027);
nand U2191 (N_2191,N_2020,N_2058);
xor U2192 (N_2192,N_1943,N_1986);
nor U2193 (N_2193,N_1965,N_2027);
xnor U2194 (N_2194,N_1927,N_2003);
and U2195 (N_2195,N_1963,N_2034);
or U2196 (N_2196,N_1978,N_1957);
or U2197 (N_2197,N_1924,N_1969);
nor U2198 (N_2198,N_1990,N_2029);
nand U2199 (N_2199,N_2053,N_2025);
nor U2200 (N_2200,N_2064,N_1996);
nor U2201 (N_2201,N_1966,N_2002);
xor U2202 (N_2202,N_1994,N_1923);
or U2203 (N_2203,N_2062,N_1941);
or U2204 (N_2204,N_1945,N_1937);
and U2205 (N_2205,N_2021,N_2046);
and U2206 (N_2206,N_2048,N_2005);
nor U2207 (N_2207,N_2053,N_2065);
or U2208 (N_2208,N_2005,N_1939);
xnor U2209 (N_2209,N_2055,N_1920);
nand U2210 (N_2210,N_1923,N_2011);
nand U2211 (N_2211,N_2030,N_2028);
nand U2212 (N_2212,N_1939,N_2044);
or U2213 (N_2213,N_1928,N_1925);
nor U2214 (N_2214,N_1977,N_1988);
nor U2215 (N_2215,N_1950,N_1930);
xor U2216 (N_2216,N_2032,N_1974);
and U2217 (N_2217,N_1987,N_2063);
nor U2218 (N_2218,N_2033,N_1944);
nand U2219 (N_2219,N_2000,N_2037);
nand U2220 (N_2220,N_2067,N_1990);
or U2221 (N_2221,N_2006,N_2034);
nand U2222 (N_2222,N_1950,N_1943);
or U2223 (N_2223,N_1987,N_2018);
and U2224 (N_2224,N_2050,N_2029);
and U2225 (N_2225,N_1955,N_2010);
and U2226 (N_2226,N_2055,N_2006);
nor U2227 (N_2227,N_1982,N_1945);
and U2228 (N_2228,N_1945,N_2021);
and U2229 (N_2229,N_2015,N_1946);
nor U2230 (N_2230,N_1980,N_1920);
and U2231 (N_2231,N_1943,N_2065);
xnor U2232 (N_2232,N_2008,N_1958);
nand U2233 (N_2233,N_2007,N_2043);
nand U2234 (N_2234,N_2042,N_2033);
nor U2235 (N_2235,N_1941,N_2004);
nor U2236 (N_2236,N_1985,N_1954);
or U2237 (N_2237,N_2076,N_2032);
nand U2238 (N_2238,N_2023,N_2008);
nand U2239 (N_2239,N_1935,N_2018);
xnor U2240 (N_2240,N_2146,N_2196);
nand U2241 (N_2241,N_2179,N_2171);
or U2242 (N_2242,N_2163,N_2177);
or U2243 (N_2243,N_2159,N_2148);
nor U2244 (N_2244,N_2087,N_2116);
or U2245 (N_2245,N_2180,N_2213);
xor U2246 (N_2246,N_2115,N_2147);
nor U2247 (N_2247,N_2142,N_2155);
nand U2248 (N_2248,N_2096,N_2141);
xnor U2249 (N_2249,N_2164,N_2118);
and U2250 (N_2250,N_2190,N_2088);
xnor U2251 (N_2251,N_2110,N_2083);
or U2252 (N_2252,N_2099,N_2134);
or U2253 (N_2253,N_2193,N_2175);
or U2254 (N_2254,N_2227,N_2168);
or U2255 (N_2255,N_2231,N_2086);
nand U2256 (N_2256,N_2184,N_2174);
nor U2257 (N_2257,N_2122,N_2121);
and U2258 (N_2258,N_2172,N_2217);
nand U2259 (N_2259,N_2204,N_2080);
nand U2260 (N_2260,N_2199,N_2239);
xor U2261 (N_2261,N_2150,N_2205);
nand U2262 (N_2262,N_2100,N_2212);
nand U2263 (N_2263,N_2166,N_2145);
or U2264 (N_2264,N_2136,N_2181);
and U2265 (N_2265,N_2149,N_2229);
xnor U2266 (N_2266,N_2089,N_2173);
and U2267 (N_2267,N_2207,N_2151);
nor U2268 (N_2268,N_2206,N_2197);
or U2269 (N_2269,N_2108,N_2143);
and U2270 (N_2270,N_2123,N_2084);
or U2271 (N_2271,N_2201,N_2152);
nand U2272 (N_2272,N_2176,N_2219);
and U2273 (N_2273,N_2234,N_2183);
nand U2274 (N_2274,N_2178,N_2191);
nand U2275 (N_2275,N_2104,N_2119);
nand U2276 (N_2276,N_2117,N_2228);
nor U2277 (N_2277,N_2235,N_2156);
nand U2278 (N_2278,N_2097,N_2107);
xnor U2279 (N_2279,N_2182,N_2124);
xor U2280 (N_2280,N_2202,N_2113);
nand U2281 (N_2281,N_2216,N_2198);
nand U2282 (N_2282,N_2232,N_2167);
or U2283 (N_2283,N_2126,N_2082);
nand U2284 (N_2284,N_2165,N_2161);
nor U2285 (N_2285,N_2162,N_2132);
or U2286 (N_2286,N_2220,N_2209);
xnor U2287 (N_2287,N_2157,N_2192);
xor U2288 (N_2288,N_2169,N_2114);
or U2289 (N_2289,N_2106,N_2139);
or U2290 (N_2290,N_2131,N_2233);
nand U2291 (N_2291,N_2238,N_2185);
or U2292 (N_2292,N_2111,N_2128);
nand U2293 (N_2293,N_2153,N_2154);
nand U2294 (N_2294,N_2127,N_2222);
xnor U2295 (N_2295,N_2138,N_2214);
and U2296 (N_2296,N_2092,N_2189);
nor U2297 (N_2297,N_2109,N_2130);
xnor U2298 (N_2298,N_2102,N_2223);
nand U2299 (N_2299,N_2125,N_2160);
and U2300 (N_2300,N_2195,N_2094);
nand U2301 (N_2301,N_2133,N_2203);
and U2302 (N_2302,N_2103,N_2098);
xnor U2303 (N_2303,N_2158,N_2144);
or U2304 (N_2304,N_2188,N_2186);
xnor U2305 (N_2305,N_2237,N_2226);
and U2306 (N_2306,N_2101,N_2105);
nor U2307 (N_2307,N_2208,N_2230);
and U2308 (N_2308,N_2120,N_2236);
xor U2309 (N_2309,N_2129,N_2221);
nand U2310 (N_2310,N_2218,N_2091);
nor U2311 (N_2311,N_2093,N_2224);
or U2312 (N_2312,N_2211,N_2137);
or U2313 (N_2313,N_2085,N_2090);
nand U2314 (N_2314,N_2215,N_2210);
and U2315 (N_2315,N_2170,N_2187);
or U2316 (N_2316,N_2112,N_2081);
and U2317 (N_2317,N_2194,N_2095);
nand U2318 (N_2318,N_2140,N_2225);
nor U2319 (N_2319,N_2135,N_2200);
or U2320 (N_2320,N_2160,N_2183);
nor U2321 (N_2321,N_2239,N_2096);
xnor U2322 (N_2322,N_2097,N_2110);
or U2323 (N_2323,N_2130,N_2160);
xor U2324 (N_2324,N_2211,N_2163);
or U2325 (N_2325,N_2119,N_2108);
xor U2326 (N_2326,N_2209,N_2096);
or U2327 (N_2327,N_2100,N_2196);
and U2328 (N_2328,N_2087,N_2239);
xnor U2329 (N_2329,N_2157,N_2094);
nand U2330 (N_2330,N_2094,N_2171);
or U2331 (N_2331,N_2157,N_2155);
nand U2332 (N_2332,N_2152,N_2114);
xnor U2333 (N_2333,N_2169,N_2186);
nand U2334 (N_2334,N_2104,N_2224);
nand U2335 (N_2335,N_2172,N_2150);
nor U2336 (N_2336,N_2165,N_2230);
nand U2337 (N_2337,N_2125,N_2080);
nor U2338 (N_2338,N_2192,N_2191);
nand U2339 (N_2339,N_2185,N_2087);
or U2340 (N_2340,N_2185,N_2123);
and U2341 (N_2341,N_2137,N_2221);
or U2342 (N_2342,N_2177,N_2162);
nand U2343 (N_2343,N_2094,N_2193);
nand U2344 (N_2344,N_2174,N_2098);
and U2345 (N_2345,N_2081,N_2150);
xnor U2346 (N_2346,N_2168,N_2101);
xnor U2347 (N_2347,N_2125,N_2176);
and U2348 (N_2348,N_2223,N_2155);
nor U2349 (N_2349,N_2184,N_2145);
xnor U2350 (N_2350,N_2190,N_2145);
nand U2351 (N_2351,N_2116,N_2182);
xor U2352 (N_2352,N_2148,N_2190);
and U2353 (N_2353,N_2104,N_2211);
nand U2354 (N_2354,N_2139,N_2209);
xor U2355 (N_2355,N_2187,N_2203);
or U2356 (N_2356,N_2109,N_2101);
nor U2357 (N_2357,N_2157,N_2144);
nand U2358 (N_2358,N_2101,N_2108);
or U2359 (N_2359,N_2119,N_2224);
and U2360 (N_2360,N_2154,N_2211);
nor U2361 (N_2361,N_2159,N_2211);
xor U2362 (N_2362,N_2104,N_2198);
or U2363 (N_2363,N_2232,N_2145);
or U2364 (N_2364,N_2088,N_2218);
nor U2365 (N_2365,N_2084,N_2175);
nor U2366 (N_2366,N_2087,N_2114);
and U2367 (N_2367,N_2102,N_2174);
xor U2368 (N_2368,N_2092,N_2214);
and U2369 (N_2369,N_2116,N_2132);
xor U2370 (N_2370,N_2181,N_2205);
nand U2371 (N_2371,N_2184,N_2100);
nand U2372 (N_2372,N_2103,N_2147);
nand U2373 (N_2373,N_2177,N_2118);
xnor U2374 (N_2374,N_2183,N_2162);
or U2375 (N_2375,N_2174,N_2186);
nor U2376 (N_2376,N_2226,N_2229);
or U2377 (N_2377,N_2148,N_2225);
nor U2378 (N_2378,N_2144,N_2234);
nor U2379 (N_2379,N_2133,N_2164);
xnor U2380 (N_2380,N_2156,N_2158);
or U2381 (N_2381,N_2209,N_2165);
and U2382 (N_2382,N_2147,N_2092);
and U2383 (N_2383,N_2199,N_2176);
xor U2384 (N_2384,N_2185,N_2152);
xnor U2385 (N_2385,N_2093,N_2085);
xor U2386 (N_2386,N_2123,N_2109);
nand U2387 (N_2387,N_2136,N_2237);
and U2388 (N_2388,N_2161,N_2190);
xnor U2389 (N_2389,N_2102,N_2156);
nand U2390 (N_2390,N_2236,N_2082);
nor U2391 (N_2391,N_2204,N_2118);
or U2392 (N_2392,N_2092,N_2141);
nor U2393 (N_2393,N_2218,N_2228);
nand U2394 (N_2394,N_2237,N_2176);
xor U2395 (N_2395,N_2096,N_2162);
or U2396 (N_2396,N_2158,N_2114);
xor U2397 (N_2397,N_2238,N_2234);
nor U2398 (N_2398,N_2163,N_2179);
and U2399 (N_2399,N_2170,N_2147);
nand U2400 (N_2400,N_2317,N_2357);
nor U2401 (N_2401,N_2271,N_2286);
nand U2402 (N_2402,N_2291,N_2372);
xnor U2403 (N_2403,N_2264,N_2385);
or U2404 (N_2404,N_2359,N_2305);
nor U2405 (N_2405,N_2248,N_2350);
nor U2406 (N_2406,N_2282,N_2329);
and U2407 (N_2407,N_2325,N_2366);
and U2408 (N_2408,N_2367,N_2396);
nor U2409 (N_2409,N_2254,N_2364);
or U2410 (N_2410,N_2277,N_2321);
and U2411 (N_2411,N_2395,N_2334);
xor U2412 (N_2412,N_2267,N_2293);
or U2413 (N_2413,N_2273,N_2344);
and U2414 (N_2414,N_2285,N_2240);
and U2415 (N_2415,N_2301,N_2353);
xor U2416 (N_2416,N_2393,N_2298);
xnor U2417 (N_2417,N_2390,N_2352);
nand U2418 (N_2418,N_2318,N_2360);
or U2419 (N_2419,N_2268,N_2260);
nor U2420 (N_2420,N_2332,N_2311);
or U2421 (N_2421,N_2243,N_2276);
xor U2422 (N_2422,N_2275,N_2375);
nor U2423 (N_2423,N_2245,N_2322);
nand U2424 (N_2424,N_2369,N_2287);
xnor U2425 (N_2425,N_2269,N_2341);
and U2426 (N_2426,N_2255,N_2336);
and U2427 (N_2427,N_2278,N_2250);
nand U2428 (N_2428,N_2378,N_2331);
nand U2429 (N_2429,N_2398,N_2347);
xnor U2430 (N_2430,N_2288,N_2251);
nand U2431 (N_2431,N_2241,N_2339);
xor U2432 (N_2432,N_2380,N_2302);
nand U2433 (N_2433,N_2361,N_2328);
xor U2434 (N_2434,N_2354,N_2296);
and U2435 (N_2435,N_2356,N_2368);
or U2436 (N_2436,N_2306,N_2299);
xor U2437 (N_2437,N_2326,N_2307);
xor U2438 (N_2438,N_2274,N_2379);
nand U2439 (N_2439,N_2397,N_2242);
xnor U2440 (N_2440,N_2300,N_2358);
nor U2441 (N_2441,N_2391,N_2244);
xor U2442 (N_2442,N_2387,N_2297);
and U2443 (N_2443,N_2309,N_2363);
nand U2444 (N_2444,N_2280,N_2371);
nand U2445 (N_2445,N_2365,N_2374);
nor U2446 (N_2446,N_2383,N_2289);
xnor U2447 (N_2447,N_2247,N_2290);
or U2448 (N_2448,N_2304,N_2257);
nor U2449 (N_2449,N_2388,N_2266);
and U2450 (N_2450,N_2263,N_2381);
or U2451 (N_2451,N_2335,N_2308);
nor U2452 (N_2452,N_2310,N_2265);
nand U2453 (N_2453,N_2323,N_2386);
nor U2454 (N_2454,N_2370,N_2258);
or U2455 (N_2455,N_2252,N_2303);
or U2456 (N_2456,N_2340,N_2373);
and U2457 (N_2457,N_2342,N_2249);
nand U2458 (N_2458,N_2382,N_2389);
nand U2459 (N_2459,N_2262,N_2355);
or U2460 (N_2460,N_2376,N_2279);
nand U2461 (N_2461,N_2315,N_2324);
nand U2462 (N_2462,N_2349,N_2316);
xnor U2463 (N_2463,N_2377,N_2333);
or U2464 (N_2464,N_2246,N_2283);
nand U2465 (N_2465,N_2394,N_2346);
xnor U2466 (N_2466,N_2384,N_2337);
xnor U2467 (N_2467,N_2259,N_2292);
or U2468 (N_2468,N_2320,N_2256);
xor U2469 (N_2469,N_2284,N_2314);
and U2470 (N_2470,N_2313,N_2281);
nor U2471 (N_2471,N_2348,N_2272);
or U2472 (N_2472,N_2319,N_2327);
and U2473 (N_2473,N_2253,N_2312);
xor U2474 (N_2474,N_2392,N_2338);
xnor U2475 (N_2475,N_2362,N_2399);
xor U2476 (N_2476,N_2343,N_2270);
and U2477 (N_2477,N_2345,N_2295);
and U2478 (N_2478,N_2351,N_2294);
nor U2479 (N_2479,N_2330,N_2261);
nand U2480 (N_2480,N_2337,N_2249);
or U2481 (N_2481,N_2319,N_2249);
xnor U2482 (N_2482,N_2247,N_2253);
xor U2483 (N_2483,N_2338,N_2350);
or U2484 (N_2484,N_2331,N_2258);
nor U2485 (N_2485,N_2308,N_2246);
and U2486 (N_2486,N_2314,N_2247);
and U2487 (N_2487,N_2301,N_2241);
or U2488 (N_2488,N_2265,N_2361);
or U2489 (N_2489,N_2381,N_2300);
or U2490 (N_2490,N_2367,N_2310);
or U2491 (N_2491,N_2354,N_2395);
nand U2492 (N_2492,N_2366,N_2268);
xor U2493 (N_2493,N_2355,N_2395);
nand U2494 (N_2494,N_2250,N_2383);
and U2495 (N_2495,N_2357,N_2390);
nor U2496 (N_2496,N_2385,N_2338);
xor U2497 (N_2497,N_2280,N_2350);
nand U2498 (N_2498,N_2243,N_2347);
nor U2499 (N_2499,N_2281,N_2352);
nor U2500 (N_2500,N_2276,N_2267);
and U2501 (N_2501,N_2246,N_2269);
nor U2502 (N_2502,N_2302,N_2269);
nand U2503 (N_2503,N_2334,N_2286);
nand U2504 (N_2504,N_2392,N_2336);
xor U2505 (N_2505,N_2293,N_2336);
xnor U2506 (N_2506,N_2357,N_2265);
nand U2507 (N_2507,N_2325,N_2358);
and U2508 (N_2508,N_2277,N_2343);
and U2509 (N_2509,N_2366,N_2282);
nor U2510 (N_2510,N_2321,N_2310);
and U2511 (N_2511,N_2260,N_2312);
nor U2512 (N_2512,N_2355,N_2329);
nor U2513 (N_2513,N_2369,N_2382);
nor U2514 (N_2514,N_2270,N_2395);
and U2515 (N_2515,N_2333,N_2345);
xnor U2516 (N_2516,N_2254,N_2385);
xnor U2517 (N_2517,N_2321,N_2385);
and U2518 (N_2518,N_2375,N_2334);
and U2519 (N_2519,N_2279,N_2274);
xnor U2520 (N_2520,N_2315,N_2262);
or U2521 (N_2521,N_2362,N_2318);
nor U2522 (N_2522,N_2379,N_2317);
or U2523 (N_2523,N_2303,N_2251);
nand U2524 (N_2524,N_2268,N_2299);
xor U2525 (N_2525,N_2283,N_2287);
nand U2526 (N_2526,N_2288,N_2325);
and U2527 (N_2527,N_2252,N_2357);
xnor U2528 (N_2528,N_2242,N_2337);
or U2529 (N_2529,N_2288,N_2384);
or U2530 (N_2530,N_2256,N_2285);
nand U2531 (N_2531,N_2396,N_2332);
nor U2532 (N_2532,N_2323,N_2304);
nand U2533 (N_2533,N_2379,N_2299);
and U2534 (N_2534,N_2338,N_2293);
and U2535 (N_2535,N_2338,N_2279);
xor U2536 (N_2536,N_2314,N_2277);
and U2537 (N_2537,N_2385,N_2279);
or U2538 (N_2538,N_2279,N_2297);
and U2539 (N_2539,N_2250,N_2245);
nand U2540 (N_2540,N_2250,N_2377);
nand U2541 (N_2541,N_2392,N_2387);
or U2542 (N_2542,N_2395,N_2287);
and U2543 (N_2543,N_2250,N_2292);
nand U2544 (N_2544,N_2399,N_2299);
or U2545 (N_2545,N_2336,N_2298);
and U2546 (N_2546,N_2359,N_2345);
nand U2547 (N_2547,N_2240,N_2283);
nor U2548 (N_2548,N_2248,N_2310);
nand U2549 (N_2549,N_2322,N_2292);
and U2550 (N_2550,N_2270,N_2260);
and U2551 (N_2551,N_2343,N_2323);
xor U2552 (N_2552,N_2260,N_2367);
nand U2553 (N_2553,N_2334,N_2387);
or U2554 (N_2554,N_2399,N_2283);
xor U2555 (N_2555,N_2361,N_2338);
and U2556 (N_2556,N_2290,N_2310);
xnor U2557 (N_2557,N_2296,N_2395);
or U2558 (N_2558,N_2348,N_2395);
and U2559 (N_2559,N_2296,N_2314);
nor U2560 (N_2560,N_2540,N_2459);
nand U2561 (N_2561,N_2521,N_2458);
and U2562 (N_2562,N_2439,N_2505);
or U2563 (N_2563,N_2514,N_2545);
and U2564 (N_2564,N_2492,N_2450);
xor U2565 (N_2565,N_2552,N_2474);
nor U2566 (N_2566,N_2435,N_2461);
and U2567 (N_2567,N_2468,N_2426);
nor U2568 (N_2568,N_2408,N_2478);
or U2569 (N_2569,N_2511,N_2462);
and U2570 (N_2570,N_2463,N_2529);
nor U2571 (N_2571,N_2436,N_2416);
or U2572 (N_2572,N_2472,N_2424);
or U2573 (N_2573,N_2465,N_2479);
nand U2574 (N_2574,N_2440,N_2525);
and U2575 (N_2575,N_2473,N_2453);
or U2576 (N_2576,N_2464,N_2486);
xnor U2577 (N_2577,N_2510,N_2509);
nor U2578 (N_2578,N_2410,N_2490);
and U2579 (N_2579,N_2541,N_2536);
xnor U2580 (N_2580,N_2412,N_2523);
and U2581 (N_2581,N_2409,N_2415);
and U2582 (N_2582,N_2497,N_2498);
nor U2583 (N_2583,N_2522,N_2423);
and U2584 (N_2584,N_2420,N_2488);
nor U2585 (N_2585,N_2475,N_2407);
nand U2586 (N_2586,N_2531,N_2542);
and U2587 (N_2587,N_2553,N_2516);
nand U2588 (N_2588,N_2451,N_2437);
and U2589 (N_2589,N_2487,N_2452);
or U2590 (N_2590,N_2538,N_2454);
and U2591 (N_2591,N_2419,N_2499);
or U2592 (N_2592,N_2433,N_2449);
or U2593 (N_2593,N_2403,N_2432);
nand U2594 (N_2594,N_2405,N_2512);
or U2595 (N_2595,N_2485,N_2548);
and U2596 (N_2596,N_2556,N_2513);
and U2597 (N_2597,N_2500,N_2429);
nand U2598 (N_2598,N_2491,N_2400);
nor U2599 (N_2599,N_2425,N_2554);
or U2600 (N_2600,N_2406,N_2528);
and U2601 (N_2601,N_2413,N_2504);
or U2602 (N_2602,N_2550,N_2508);
nor U2603 (N_2603,N_2418,N_2480);
or U2604 (N_2604,N_2460,N_2414);
nand U2605 (N_2605,N_2441,N_2506);
nor U2606 (N_2606,N_2448,N_2447);
and U2607 (N_2607,N_2481,N_2484);
xnor U2608 (N_2608,N_2430,N_2466);
and U2609 (N_2609,N_2535,N_2421);
and U2610 (N_2610,N_2549,N_2537);
and U2611 (N_2611,N_2476,N_2530);
nor U2612 (N_2612,N_2434,N_2526);
or U2613 (N_2613,N_2493,N_2477);
and U2614 (N_2614,N_2558,N_2470);
and U2615 (N_2615,N_2457,N_2524);
xnor U2616 (N_2616,N_2483,N_2551);
nand U2617 (N_2617,N_2442,N_2444);
and U2618 (N_2618,N_2456,N_2559);
nand U2619 (N_2619,N_2489,N_2527);
nor U2620 (N_2620,N_2402,N_2532);
and U2621 (N_2621,N_2557,N_2496);
nor U2622 (N_2622,N_2431,N_2427);
or U2623 (N_2623,N_2411,N_2539);
and U2624 (N_2624,N_2534,N_2494);
nor U2625 (N_2625,N_2517,N_2546);
xor U2626 (N_2626,N_2555,N_2544);
xnor U2627 (N_2627,N_2469,N_2533);
xnor U2628 (N_2628,N_2547,N_2482);
or U2629 (N_2629,N_2422,N_2543);
and U2630 (N_2630,N_2455,N_2501);
nand U2631 (N_2631,N_2515,N_2445);
nor U2632 (N_2632,N_2467,N_2507);
or U2633 (N_2633,N_2520,N_2471);
nor U2634 (N_2634,N_2438,N_2519);
nor U2635 (N_2635,N_2428,N_2446);
xor U2636 (N_2636,N_2503,N_2404);
nand U2637 (N_2637,N_2518,N_2401);
or U2638 (N_2638,N_2495,N_2502);
nand U2639 (N_2639,N_2443,N_2417);
and U2640 (N_2640,N_2507,N_2408);
and U2641 (N_2641,N_2423,N_2488);
xor U2642 (N_2642,N_2436,N_2454);
nand U2643 (N_2643,N_2435,N_2521);
nor U2644 (N_2644,N_2559,N_2527);
nor U2645 (N_2645,N_2469,N_2467);
or U2646 (N_2646,N_2474,N_2453);
nand U2647 (N_2647,N_2549,N_2492);
nand U2648 (N_2648,N_2548,N_2460);
xor U2649 (N_2649,N_2483,N_2530);
xnor U2650 (N_2650,N_2480,N_2497);
or U2651 (N_2651,N_2424,N_2544);
nand U2652 (N_2652,N_2418,N_2495);
nand U2653 (N_2653,N_2505,N_2523);
and U2654 (N_2654,N_2485,N_2410);
xor U2655 (N_2655,N_2481,N_2515);
or U2656 (N_2656,N_2401,N_2505);
xor U2657 (N_2657,N_2464,N_2432);
or U2658 (N_2658,N_2427,N_2406);
or U2659 (N_2659,N_2430,N_2503);
nor U2660 (N_2660,N_2488,N_2482);
or U2661 (N_2661,N_2515,N_2486);
nand U2662 (N_2662,N_2423,N_2497);
nand U2663 (N_2663,N_2525,N_2526);
nor U2664 (N_2664,N_2559,N_2499);
or U2665 (N_2665,N_2423,N_2489);
xnor U2666 (N_2666,N_2504,N_2407);
xnor U2667 (N_2667,N_2449,N_2476);
xor U2668 (N_2668,N_2500,N_2454);
nor U2669 (N_2669,N_2474,N_2497);
xor U2670 (N_2670,N_2417,N_2456);
or U2671 (N_2671,N_2554,N_2505);
and U2672 (N_2672,N_2526,N_2557);
nand U2673 (N_2673,N_2534,N_2440);
nor U2674 (N_2674,N_2437,N_2543);
nand U2675 (N_2675,N_2517,N_2530);
nor U2676 (N_2676,N_2459,N_2520);
xor U2677 (N_2677,N_2408,N_2500);
and U2678 (N_2678,N_2548,N_2419);
xnor U2679 (N_2679,N_2500,N_2442);
nand U2680 (N_2680,N_2484,N_2445);
nand U2681 (N_2681,N_2532,N_2459);
or U2682 (N_2682,N_2437,N_2493);
nand U2683 (N_2683,N_2442,N_2493);
xor U2684 (N_2684,N_2556,N_2529);
or U2685 (N_2685,N_2529,N_2424);
or U2686 (N_2686,N_2443,N_2449);
and U2687 (N_2687,N_2550,N_2441);
xor U2688 (N_2688,N_2497,N_2435);
or U2689 (N_2689,N_2465,N_2413);
and U2690 (N_2690,N_2515,N_2557);
or U2691 (N_2691,N_2475,N_2430);
xor U2692 (N_2692,N_2546,N_2513);
nand U2693 (N_2693,N_2462,N_2417);
nand U2694 (N_2694,N_2451,N_2423);
or U2695 (N_2695,N_2467,N_2500);
nor U2696 (N_2696,N_2518,N_2460);
xnor U2697 (N_2697,N_2548,N_2480);
xnor U2698 (N_2698,N_2542,N_2457);
or U2699 (N_2699,N_2503,N_2526);
or U2700 (N_2700,N_2417,N_2420);
nand U2701 (N_2701,N_2556,N_2491);
xor U2702 (N_2702,N_2403,N_2469);
nand U2703 (N_2703,N_2515,N_2459);
xor U2704 (N_2704,N_2533,N_2502);
or U2705 (N_2705,N_2413,N_2531);
and U2706 (N_2706,N_2401,N_2549);
xor U2707 (N_2707,N_2468,N_2518);
and U2708 (N_2708,N_2426,N_2479);
nand U2709 (N_2709,N_2479,N_2461);
or U2710 (N_2710,N_2431,N_2429);
xor U2711 (N_2711,N_2514,N_2457);
xnor U2712 (N_2712,N_2442,N_2488);
nand U2713 (N_2713,N_2541,N_2400);
nand U2714 (N_2714,N_2504,N_2414);
or U2715 (N_2715,N_2510,N_2540);
xnor U2716 (N_2716,N_2498,N_2503);
or U2717 (N_2717,N_2473,N_2442);
and U2718 (N_2718,N_2559,N_2486);
nand U2719 (N_2719,N_2430,N_2486);
xor U2720 (N_2720,N_2648,N_2685);
and U2721 (N_2721,N_2677,N_2643);
nand U2722 (N_2722,N_2609,N_2702);
or U2723 (N_2723,N_2708,N_2655);
nand U2724 (N_2724,N_2680,N_2638);
xnor U2725 (N_2725,N_2651,N_2584);
or U2726 (N_2726,N_2713,N_2717);
or U2727 (N_2727,N_2691,N_2593);
and U2728 (N_2728,N_2616,N_2647);
or U2729 (N_2729,N_2591,N_2642);
xnor U2730 (N_2730,N_2620,N_2590);
nand U2731 (N_2731,N_2703,N_2574);
or U2732 (N_2732,N_2649,N_2573);
or U2733 (N_2733,N_2603,N_2633);
xor U2734 (N_2734,N_2694,N_2576);
or U2735 (N_2735,N_2704,N_2653);
nor U2736 (N_2736,N_2560,N_2661);
nand U2737 (N_2737,N_2636,N_2596);
nor U2738 (N_2738,N_2567,N_2663);
nand U2739 (N_2739,N_2598,N_2606);
nor U2740 (N_2740,N_2707,N_2645);
nand U2741 (N_2741,N_2571,N_2610);
nor U2742 (N_2742,N_2656,N_2632);
xnor U2743 (N_2743,N_2607,N_2627);
nor U2744 (N_2744,N_2563,N_2624);
xnor U2745 (N_2745,N_2582,N_2618);
nand U2746 (N_2746,N_2568,N_2673);
nor U2747 (N_2747,N_2601,N_2681);
nor U2748 (N_2748,N_2565,N_2562);
nand U2749 (N_2749,N_2639,N_2604);
or U2750 (N_2750,N_2577,N_2668);
nand U2751 (N_2751,N_2715,N_2682);
or U2752 (N_2752,N_2689,N_2697);
nand U2753 (N_2753,N_2602,N_2611);
and U2754 (N_2754,N_2660,N_2587);
and U2755 (N_2755,N_2619,N_2629);
or U2756 (N_2756,N_2637,N_2688);
and U2757 (N_2757,N_2613,N_2646);
or U2758 (N_2758,N_2622,N_2695);
nor U2759 (N_2759,N_2561,N_2672);
nor U2760 (N_2760,N_2667,N_2706);
nand U2761 (N_2761,N_2634,N_2712);
and U2762 (N_2762,N_2714,N_2696);
or U2763 (N_2763,N_2719,N_2625);
xnor U2764 (N_2764,N_2569,N_2583);
and U2765 (N_2765,N_2705,N_2614);
xnor U2766 (N_2766,N_2631,N_2710);
and U2767 (N_2767,N_2617,N_2630);
nand U2768 (N_2768,N_2670,N_2658);
or U2769 (N_2769,N_2687,N_2671);
nand U2770 (N_2770,N_2701,N_2659);
nor U2771 (N_2771,N_2575,N_2580);
and U2772 (N_2772,N_2652,N_2581);
and U2773 (N_2773,N_2566,N_2654);
nor U2774 (N_2774,N_2678,N_2586);
nand U2775 (N_2775,N_2675,N_2676);
nor U2776 (N_2776,N_2628,N_2626);
nor U2777 (N_2777,N_2683,N_2644);
and U2778 (N_2778,N_2608,N_2595);
or U2779 (N_2779,N_2592,N_2564);
nor U2780 (N_2780,N_2579,N_2621);
nand U2781 (N_2781,N_2679,N_2605);
and U2782 (N_2782,N_2662,N_2588);
xor U2783 (N_2783,N_2599,N_2594);
nand U2784 (N_2784,N_2692,N_2572);
nand U2785 (N_2785,N_2711,N_2640);
nor U2786 (N_2786,N_2674,N_2666);
nand U2787 (N_2787,N_2641,N_2615);
and U2788 (N_2788,N_2686,N_2612);
xor U2789 (N_2789,N_2578,N_2570);
nor U2790 (N_2790,N_2669,N_2600);
nand U2791 (N_2791,N_2698,N_2716);
or U2792 (N_2792,N_2693,N_2684);
xor U2793 (N_2793,N_2657,N_2664);
xnor U2794 (N_2794,N_2699,N_2700);
xor U2795 (N_2795,N_2589,N_2709);
nor U2796 (N_2796,N_2718,N_2623);
or U2797 (N_2797,N_2665,N_2690);
nor U2798 (N_2798,N_2635,N_2650);
and U2799 (N_2799,N_2585,N_2597);
or U2800 (N_2800,N_2609,N_2601);
nand U2801 (N_2801,N_2571,N_2649);
nor U2802 (N_2802,N_2674,N_2658);
and U2803 (N_2803,N_2686,N_2716);
xor U2804 (N_2804,N_2636,N_2626);
nand U2805 (N_2805,N_2688,N_2583);
or U2806 (N_2806,N_2604,N_2602);
nor U2807 (N_2807,N_2623,N_2563);
and U2808 (N_2808,N_2569,N_2587);
or U2809 (N_2809,N_2699,N_2577);
xnor U2810 (N_2810,N_2628,N_2710);
nor U2811 (N_2811,N_2626,N_2676);
or U2812 (N_2812,N_2603,N_2703);
nand U2813 (N_2813,N_2604,N_2666);
nor U2814 (N_2814,N_2664,N_2638);
or U2815 (N_2815,N_2631,N_2562);
nor U2816 (N_2816,N_2643,N_2641);
xor U2817 (N_2817,N_2707,N_2580);
xor U2818 (N_2818,N_2581,N_2578);
or U2819 (N_2819,N_2628,N_2618);
and U2820 (N_2820,N_2687,N_2717);
nor U2821 (N_2821,N_2565,N_2632);
and U2822 (N_2822,N_2665,N_2712);
nand U2823 (N_2823,N_2701,N_2678);
xnor U2824 (N_2824,N_2622,N_2713);
nand U2825 (N_2825,N_2596,N_2705);
and U2826 (N_2826,N_2587,N_2562);
or U2827 (N_2827,N_2710,N_2695);
nor U2828 (N_2828,N_2651,N_2681);
nand U2829 (N_2829,N_2615,N_2681);
nor U2830 (N_2830,N_2597,N_2690);
xor U2831 (N_2831,N_2635,N_2596);
nor U2832 (N_2832,N_2566,N_2592);
or U2833 (N_2833,N_2654,N_2698);
or U2834 (N_2834,N_2626,N_2698);
nor U2835 (N_2835,N_2560,N_2691);
nand U2836 (N_2836,N_2560,N_2714);
xnor U2837 (N_2837,N_2667,N_2710);
nand U2838 (N_2838,N_2575,N_2685);
or U2839 (N_2839,N_2562,N_2632);
xor U2840 (N_2840,N_2571,N_2679);
nand U2841 (N_2841,N_2687,N_2648);
xnor U2842 (N_2842,N_2621,N_2708);
xor U2843 (N_2843,N_2576,N_2661);
and U2844 (N_2844,N_2562,N_2592);
and U2845 (N_2845,N_2711,N_2584);
xnor U2846 (N_2846,N_2606,N_2690);
nor U2847 (N_2847,N_2642,N_2580);
xnor U2848 (N_2848,N_2587,N_2683);
or U2849 (N_2849,N_2633,N_2592);
xnor U2850 (N_2850,N_2695,N_2635);
and U2851 (N_2851,N_2669,N_2639);
nand U2852 (N_2852,N_2640,N_2694);
xor U2853 (N_2853,N_2561,N_2692);
and U2854 (N_2854,N_2711,N_2650);
nor U2855 (N_2855,N_2678,N_2580);
and U2856 (N_2856,N_2715,N_2663);
nor U2857 (N_2857,N_2642,N_2632);
or U2858 (N_2858,N_2693,N_2618);
and U2859 (N_2859,N_2651,N_2591);
nand U2860 (N_2860,N_2570,N_2663);
xor U2861 (N_2861,N_2701,N_2692);
xor U2862 (N_2862,N_2604,N_2625);
or U2863 (N_2863,N_2608,N_2664);
nor U2864 (N_2864,N_2586,N_2591);
and U2865 (N_2865,N_2695,N_2640);
nand U2866 (N_2866,N_2681,N_2595);
or U2867 (N_2867,N_2667,N_2634);
nor U2868 (N_2868,N_2667,N_2677);
and U2869 (N_2869,N_2657,N_2696);
nand U2870 (N_2870,N_2587,N_2674);
nor U2871 (N_2871,N_2645,N_2704);
nor U2872 (N_2872,N_2590,N_2637);
nand U2873 (N_2873,N_2600,N_2572);
nor U2874 (N_2874,N_2660,N_2626);
xnor U2875 (N_2875,N_2600,N_2649);
xor U2876 (N_2876,N_2656,N_2696);
or U2877 (N_2877,N_2598,N_2563);
xnor U2878 (N_2878,N_2587,N_2576);
xor U2879 (N_2879,N_2653,N_2595);
nor U2880 (N_2880,N_2866,N_2806);
or U2881 (N_2881,N_2829,N_2877);
or U2882 (N_2882,N_2779,N_2751);
and U2883 (N_2883,N_2721,N_2725);
nand U2884 (N_2884,N_2747,N_2805);
and U2885 (N_2885,N_2850,N_2809);
nor U2886 (N_2886,N_2851,N_2836);
nand U2887 (N_2887,N_2788,N_2838);
and U2888 (N_2888,N_2773,N_2798);
and U2889 (N_2889,N_2874,N_2879);
xor U2890 (N_2890,N_2864,N_2857);
nor U2891 (N_2891,N_2731,N_2828);
nor U2892 (N_2892,N_2765,N_2755);
and U2893 (N_2893,N_2786,N_2768);
nand U2894 (N_2894,N_2812,N_2826);
and U2895 (N_2895,N_2872,N_2837);
nand U2896 (N_2896,N_2834,N_2816);
nand U2897 (N_2897,N_2817,N_2776);
nor U2898 (N_2898,N_2796,N_2784);
xor U2899 (N_2899,N_2761,N_2754);
and U2900 (N_2900,N_2859,N_2744);
and U2901 (N_2901,N_2832,N_2760);
or U2902 (N_2902,N_2759,N_2750);
nor U2903 (N_2903,N_2801,N_2726);
nand U2904 (N_2904,N_2808,N_2763);
and U2905 (N_2905,N_2827,N_2794);
xor U2906 (N_2906,N_2831,N_2791);
and U2907 (N_2907,N_2736,N_2793);
nor U2908 (N_2908,N_2840,N_2800);
xnor U2909 (N_2909,N_2771,N_2739);
or U2910 (N_2910,N_2847,N_2862);
nor U2911 (N_2911,N_2875,N_2873);
or U2912 (N_2912,N_2858,N_2799);
nor U2913 (N_2913,N_2743,N_2766);
nor U2914 (N_2914,N_2839,N_2803);
and U2915 (N_2915,N_2752,N_2749);
xor U2916 (N_2916,N_2753,N_2748);
nor U2917 (N_2917,N_2738,N_2822);
or U2918 (N_2918,N_2856,N_2767);
or U2919 (N_2919,N_2815,N_2804);
and U2920 (N_2920,N_2819,N_2846);
nand U2921 (N_2921,N_2865,N_2848);
xnor U2922 (N_2922,N_2841,N_2835);
nand U2923 (N_2923,N_2729,N_2811);
nand U2924 (N_2924,N_2724,N_2842);
nor U2925 (N_2925,N_2833,N_2869);
and U2926 (N_2926,N_2780,N_2789);
and U2927 (N_2927,N_2782,N_2756);
nand U2928 (N_2928,N_2762,N_2860);
nor U2929 (N_2929,N_2734,N_2777);
nor U2930 (N_2930,N_2870,N_2787);
xor U2931 (N_2931,N_2720,N_2740);
or U2932 (N_2932,N_2797,N_2820);
nor U2933 (N_2933,N_2830,N_2795);
or U2934 (N_2934,N_2863,N_2730);
and U2935 (N_2935,N_2741,N_2813);
nor U2936 (N_2936,N_2871,N_2845);
and U2937 (N_2937,N_2732,N_2742);
nand U2938 (N_2938,N_2745,N_2843);
nor U2939 (N_2939,N_2737,N_2849);
xnor U2940 (N_2940,N_2781,N_2728);
or U2941 (N_2941,N_2823,N_2844);
xor U2942 (N_2942,N_2867,N_2868);
or U2943 (N_2943,N_2746,N_2727);
nand U2944 (N_2944,N_2825,N_2757);
xnor U2945 (N_2945,N_2818,N_2802);
xnor U2946 (N_2946,N_2876,N_2769);
and U2947 (N_2947,N_2824,N_2878);
nor U2948 (N_2948,N_2722,N_2855);
xnor U2949 (N_2949,N_2770,N_2723);
xor U2950 (N_2950,N_2778,N_2854);
or U2951 (N_2951,N_2772,N_2814);
and U2952 (N_2952,N_2792,N_2783);
nor U2953 (N_2953,N_2861,N_2821);
nor U2954 (N_2954,N_2733,N_2774);
nand U2955 (N_2955,N_2735,N_2807);
nor U2956 (N_2956,N_2785,N_2810);
nor U2957 (N_2957,N_2852,N_2764);
or U2958 (N_2958,N_2790,N_2853);
or U2959 (N_2959,N_2775,N_2758);
and U2960 (N_2960,N_2861,N_2749);
and U2961 (N_2961,N_2856,N_2771);
nand U2962 (N_2962,N_2747,N_2830);
xnor U2963 (N_2963,N_2746,N_2738);
nand U2964 (N_2964,N_2816,N_2764);
xnor U2965 (N_2965,N_2746,N_2728);
and U2966 (N_2966,N_2776,N_2745);
nor U2967 (N_2967,N_2819,N_2863);
xor U2968 (N_2968,N_2787,N_2730);
xnor U2969 (N_2969,N_2807,N_2811);
or U2970 (N_2970,N_2812,N_2853);
nand U2971 (N_2971,N_2867,N_2775);
nand U2972 (N_2972,N_2841,N_2816);
and U2973 (N_2973,N_2797,N_2726);
nor U2974 (N_2974,N_2775,N_2776);
xor U2975 (N_2975,N_2733,N_2817);
nor U2976 (N_2976,N_2791,N_2731);
nor U2977 (N_2977,N_2736,N_2731);
xor U2978 (N_2978,N_2823,N_2741);
nor U2979 (N_2979,N_2768,N_2813);
nand U2980 (N_2980,N_2809,N_2786);
nand U2981 (N_2981,N_2857,N_2729);
nor U2982 (N_2982,N_2785,N_2786);
xor U2983 (N_2983,N_2781,N_2849);
and U2984 (N_2984,N_2744,N_2819);
nor U2985 (N_2985,N_2776,N_2748);
xor U2986 (N_2986,N_2761,N_2744);
xnor U2987 (N_2987,N_2748,N_2762);
and U2988 (N_2988,N_2847,N_2756);
or U2989 (N_2989,N_2727,N_2754);
nor U2990 (N_2990,N_2857,N_2825);
or U2991 (N_2991,N_2747,N_2875);
or U2992 (N_2992,N_2879,N_2801);
nor U2993 (N_2993,N_2815,N_2844);
or U2994 (N_2994,N_2766,N_2733);
and U2995 (N_2995,N_2879,N_2754);
nand U2996 (N_2996,N_2796,N_2732);
or U2997 (N_2997,N_2827,N_2725);
xor U2998 (N_2998,N_2753,N_2810);
nand U2999 (N_2999,N_2753,N_2791);
nand U3000 (N_3000,N_2746,N_2737);
nand U3001 (N_3001,N_2816,N_2868);
nor U3002 (N_3002,N_2872,N_2816);
nand U3003 (N_3003,N_2836,N_2867);
nor U3004 (N_3004,N_2877,N_2776);
xor U3005 (N_3005,N_2749,N_2720);
xnor U3006 (N_3006,N_2752,N_2829);
nor U3007 (N_3007,N_2767,N_2722);
or U3008 (N_3008,N_2793,N_2757);
nor U3009 (N_3009,N_2814,N_2729);
or U3010 (N_3010,N_2769,N_2777);
xnor U3011 (N_3011,N_2727,N_2813);
xnor U3012 (N_3012,N_2728,N_2733);
and U3013 (N_3013,N_2720,N_2854);
xor U3014 (N_3014,N_2738,N_2848);
nand U3015 (N_3015,N_2725,N_2747);
xor U3016 (N_3016,N_2843,N_2762);
nand U3017 (N_3017,N_2842,N_2727);
xor U3018 (N_3018,N_2830,N_2802);
nand U3019 (N_3019,N_2863,N_2766);
xor U3020 (N_3020,N_2813,N_2873);
nor U3021 (N_3021,N_2835,N_2849);
nand U3022 (N_3022,N_2730,N_2741);
or U3023 (N_3023,N_2804,N_2805);
nand U3024 (N_3024,N_2811,N_2830);
and U3025 (N_3025,N_2723,N_2821);
nand U3026 (N_3026,N_2740,N_2781);
nor U3027 (N_3027,N_2853,N_2784);
and U3028 (N_3028,N_2721,N_2854);
nor U3029 (N_3029,N_2740,N_2761);
or U3030 (N_3030,N_2814,N_2790);
xor U3031 (N_3031,N_2738,N_2803);
and U3032 (N_3032,N_2781,N_2823);
nor U3033 (N_3033,N_2774,N_2798);
xnor U3034 (N_3034,N_2776,N_2846);
nor U3035 (N_3035,N_2794,N_2758);
and U3036 (N_3036,N_2876,N_2785);
nand U3037 (N_3037,N_2854,N_2789);
and U3038 (N_3038,N_2772,N_2803);
and U3039 (N_3039,N_2862,N_2799);
and U3040 (N_3040,N_2881,N_3039);
nand U3041 (N_3041,N_2938,N_2901);
and U3042 (N_3042,N_2957,N_2944);
or U3043 (N_3043,N_2891,N_3004);
or U3044 (N_3044,N_2961,N_2931);
nor U3045 (N_3045,N_2937,N_2933);
or U3046 (N_3046,N_2897,N_2893);
xnor U3047 (N_3047,N_2887,N_2998);
xnor U3048 (N_3048,N_3018,N_3008);
and U3049 (N_3049,N_3027,N_2971);
xor U3050 (N_3050,N_2895,N_3001);
or U3051 (N_3051,N_2941,N_3037);
xor U3052 (N_3052,N_2978,N_3033);
and U3053 (N_3053,N_2880,N_2885);
and U3054 (N_3054,N_2994,N_2995);
nor U3055 (N_3055,N_2980,N_3036);
xor U3056 (N_3056,N_2888,N_2913);
nand U3057 (N_3057,N_2904,N_2958);
nand U3058 (N_3058,N_2935,N_2919);
and U3059 (N_3059,N_2925,N_2907);
and U3060 (N_3060,N_3017,N_2927);
and U3061 (N_3061,N_2906,N_3011);
nor U3062 (N_3062,N_2920,N_2984);
or U3063 (N_3063,N_2890,N_2950);
and U3064 (N_3064,N_2974,N_2922);
nor U3065 (N_3065,N_3010,N_2928);
and U3066 (N_3066,N_2970,N_2900);
and U3067 (N_3067,N_2945,N_2955);
nand U3068 (N_3068,N_2926,N_2882);
or U3069 (N_3069,N_2997,N_2948);
and U3070 (N_3070,N_2883,N_2921);
or U3071 (N_3071,N_3028,N_2967);
or U3072 (N_3072,N_2989,N_3024);
and U3073 (N_3073,N_2979,N_3022);
or U3074 (N_3074,N_2910,N_3019);
nand U3075 (N_3075,N_2999,N_2902);
nor U3076 (N_3076,N_2936,N_3015);
nand U3077 (N_3077,N_2939,N_3003);
or U3078 (N_3078,N_2953,N_2908);
nor U3079 (N_3079,N_2923,N_2929);
nor U3080 (N_3080,N_3020,N_2934);
nand U3081 (N_3081,N_2960,N_2988);
and U3082 (N_3082,N_2981,N_2965);
and U3083 (N_3083,N_2951,N_2905);
nor U3084 (N_3084,N_2987,N_2894);
or U3085 (N_3085,N_2954,N_2962);
nor U3086 (N_3086,N_2976,N_3007);
nand U3087 (N_3087,N_2991,N_2985);
nand U3088 (N_3088,N_2972,N_2959);
xnor U3089 (N_3089,N_3016,N_2911);
and U3090 (N_3090,N_3029,N_2886);
or U3091 (N_3091,N_2940,N_2986);
or U3092 (N_3092,N_2912,N_3038);
and U3093 (N_3093,N_2946,N_2992);
nand U3094 (N_3094,N_2964,N_3035);
nor U3095 (N_3095,N_2993,N_3023);
and U3096 (N_3096,N_2896,N_2956);
nor U3097 (N_3097,N_3006,N_2963);
xnor U3098 (N_3098,N_3030,N_2947);
xor U3099 (N_3099,N_2884,N_2917);
or U3100 (N_3100,N_2973,N_2918);
or U3101 (N_3101,N_2899,N_2916);
xor U3102 (N_3102,N_3014,N_2892);
nor U3103 (N_3103,N_3032,N_3013);
xnor U3104 (N_3104,N_3034,N_2969);
and U3105 (N_3105,N_2889,N_2924);
nor U3106 (N_3106,N_3005,N_3009);
or U3107 (N_3107,N_2968,N_2977);
xnor U3108 (N_3108,N_2903,N_2942);
nand U3109 (N_3109,N_2975,N_2915);
xnor U3110 (N_3110,N_2932,N_3021);
or U3111 (N_3111,N_3002,N_2996);
and U3112 (N_3112,N_2909,N_2966);
or U3113 (N_3113,N_2914,N_2930);
nand U3114 (N_3114,N_3000,N_2943);
and U3115 (N_3115,N_2990,N_3026);
and U3116 (N_3116,N_2952,N_3031);
xnor U3117 (N_3117,N_2949,N_3012);
nand U3118 (N_3118,N_2982,N_2898);
nor U3119 (N_3119,N_3025,N_2983);
nor U3120 (N_3120,N_2949,N_2995);
nor U3121 (N_3121,N_2954,N_3002);
or U3122 (N_3122,N_2889,N_2971);
nor U3123 (N_3123,N_2918,N_2913);
nor U3124 (N_3124,N_2944,N_2952);
xnor U3125 (N_3125,N_2977,N_2995);
nand U3126 (N_3126,N_3001,N_2982);
nor U3127 (N_3127,N_2997,N_2984);
and U3128 (N_3128,N_2961,N_2970);
nor U3129 (N_3129,N_2941,N_2994);
and U3130 (N_3130,N_2919,N_2907);
nor U3131 (N_3131,N_2956,N_3020);
nand U3132 (N_3132,N_2999,N_2998);
nand U3133 (N_3133,N_2965,N_2999);
nand U3134 (N_3134,N_2894,N_2892);
nor U3135 (N_3135,N_2927,N_2937);
and U3136 (N_3136,N_2910,N_3006);
nand U3137 (N_3137,N_2991,N_3036);
xnor U3138 (N_3138,N_2912,N_2938);
xor U3139 (N_3139,N_3004,N_3020);
nor U3140 (N_3140,N_2941,N_3016);
or U3141 (N_3141,N_2965,N_2958);
nand U3142 (N_3142,N_2919,N_2957);
or U3143 (N_3143,N_2969,N_2930);
nand U3144 (N_3144,N_3007,N_2948);
nor U3145 (N_3145,N_2888,N_3035);
nand U3146 (N_3146,N_2957,N_2986);
xnor U3147 (N_3147,N_2914,N_3038);
nor U3148 (N_3148,N_2937,N_2956);
nand U3149 (N_3149,N_2944,N_2900);
nand U3150 (N_3150,N_2915,N_3009);
xor U3151 (N_3151,N_2989,N_3022);
nor U3152 (N_3152,N_2914,N_2932);
nand U3153 (N_3153,N_2957,N_2958);
xnor U3154 (N_3154,N_2949,N_2963);
nand U3155 (N_3155,N_2891,N_2962);
xor U3156 (N_3156,N_2888,N_3006);
xor U3157 (N_3157,N_2900,N_3020);
and U3158 (N_3158,N_2933,N_3002);
nand U3159 (N_3159,N_2947,N_2933);
and U3160 (N_3160,N_3038,N_2940);
and U3161 (N_3161,N_2968,N_2915);
xnor U3162 (N_3162,N_2979,N_2978);
nor U3163 (N_3163,N_3011,N_2881);
and U3164 (N_3164,N_2936,N_2939);
nor U3165 (N_3165,N_2947,N_2982);
xnor U3166 (N_3166,N_2957,N_3000);
nor U3167 (N_3167,N_2893,N_2919);
xor U3168 (N_3168,N_2919,N_3022);
nand U3169 (N_3169,N_2952,N_2905);
nand U3170 (N_3170,N_2957,N_3031);
nor U3171 (N_3171,N_2965,N_3030);
and U3172 (N_3172,N_2974,N_2979);
or U3173 (N_3173,N_2890,N_2978);
nand U3174 (N_3174,N_3032,N_3001);
nor U3175 (N_3175,N_2982,N_2886);
nand U3176 (N_3176,N_2987,N_2886);
nand U3177 (N_3177,N_2951,N_2947);
nand U3178 (N_3178,N_2891,N_2951);
xor U3179 (N_3179,N_2923,N_2992);
and U3180 (N_3180,N_2966,N_2939);
nor U3181 (N_3181,N_3002,N_3010);
nand U3182 (N_3182,N_2924,N_2937);
nand U3183 (N_3183,N_2884,N_2897);
or U3184 (N_3184,N_2927,N_2932);
nor U3185 (N_3185,N_3039,N_3032);
and U3186 (N_3186,N_2976,N_2958);
or U3187 (N_3187,N_2909,N_2918);
nand U3188 (N_3188,N_2974,N_2948);
nand U3189 (N_3189,N_2959,N_2990);
xnor U3190 (N_3190,N_2890,N_3015);
nor U3191 (N_3191,N_2997,N_2937);
nor U3192 (N_3192,N_2958,N_2886);
nor U3193 (N_3193,N_2963,N_2992);
and U3194 (N_3194,N_2907,N_3002);
or U3195 (N_3195,N_2967,N_2902);
or U3196 (N_3196,N_2901,N_3021);
nor U3197 (N_3197,N_2921,N_2946);
xor U3198 (N_3198,N_2947,N_2967);
nand U3199 (N_3199,N_2958,N_2962);
or U3200 (N_3200,N_3120,N_3106);
xnor U3201 (N_3201,N_3047,N_3199);
nand U3202 (N_3202,N_3044,N_3089);
or U3203 (N_3203,N_3146,N_3187);
or U3204 (N_3204,N_3159,N_3045);
nor U3205 (N_3205,N_3157,N_3069);
nor U3206 (N_3206,N_3129,N_3160);
and U3207 (N_3207,N_3158,N_3154);
xnor U3208 (N_3208,N_3074,N_3176);
or U3209 (N_3209,N_3198,N_3058);
nor U3210 (N_3210,N_3168,N_3172);
or U3211 (N_3211,N_3184,N_3061);
or U3212 (N_3212,N_3185,N_3054);
nor U3213 (N_3213,N_3156,N_3131);
xnor U3214 (N_3214,N_3093,N_3189);
nand U3215 (N_3215,N_3107,N_3060);
xnor U3216 (N_3216,N_3071,N_3092);
xnor U3217 (N_3217,N_3183,N_3086);
and U3218 (N_3218,N_3163,N_3155);
nand U3219 (N_3219,N_3164,N_3113);
nand U3220 (N_3220,N_3090,N_3197);
xor U3221 (N_3221,N_3121,N_3181);
nor U3222 (N_3222,N_3126,N_3143);
or U3223 (N_3223,N_3094,N_3178);
nand U3224 (N_3224,N_3171,N_3080);
nand U3225 (N_3225,N_3049,N_3103);
nor U3226 (N_3226,N_3072,N_3174);
or U3227 (N_3227,N_3125,N_3065);
nand U3228 (N_3228,N_3165,N_3105);
nor U3229 (N_3229,N_3188,N_3051);
nor U3230 (N_3230,N_3170,N_3057);
and U3231 (N_3231,N_3084,N_3191);
xor U3232 (N_3232,N_3050,N_3134);
or U3233 (N_3233,N_3133,N_3195);
and U3234 (N_3234,N_3112,N_3040);
nand U3235 (N_3235,N_3076,N_3180);
or U3236 (N_3236,N_3175,N_3148);
or U3237 (N_3237,N_3097,N_3147);
or U3238 (N_3238,N_3041,N_3110);
nor U3239 (N_3239,N_3109,N_3087);
xor U3240 (N_3240,N_3101,N_3102);
xnor U3241 (N_3241,N_3114,N_3118);
nor U3242 (N_3242,N_3070,N_3169);
xor U3243 (N_3243,N_3052,N_3075);
or U3244 (N_3244,N_3166,N_3139);
nand U3245 (N_3245,N_3123,N_3062);
or U3246 (N_3246,N_3081,N_3190);
nor U3247 (N_3247,N_3141,N_3108);
nand U3248 (N_3248,N_3098,N_3152);
xor U3249 (N_3249,N_3048,N_3063);
and U3250 (N_3250,N_3079,N_3186);
or U3251 (N_3251,N_3056,N_3130);
or U3252 (N_3252,N_3173,N_3117);
or U3253 (N_3253,N_3142,N_3085);
nand U3254 (N_3254,N_3151,N_3116);
and U3255 (N_3255,N_3104,N_3091);
nand U3256 (N_3256,N_3132,N_3179);
xnor U3257 (N_3257,N_3055,N_3115);
or U3258 (N_3258,N_3073,N_3127);
nor U3259 (N_3259,N_3067,N_3144);
or U3260 (N_3260,N_3088,N_3119);
nand U3261 (N_3261,N_3082,N_3053);
or U3262 (N_3262,N_3124,N_3150);
and U3263 (N_3263,N_3162,N_3066);
nand U3264 (N_3264,N_3096,N_3194);
and U3265 (N_3265,N_3100,N_3128);
xnor U3266 (N_3266,N_3149,N_3192);
and U3267 (N_3267,N_3182,N_3161);
and U3268 (N_3268,N_3167,N_3064);
or U3269 (N_3269,N_3153,N_3043);
nand U3270 (N_3270,N_3046,N_3059);
or U3271 (N_3271,N_3138,N_3042);
nor U3272 (N_3272,N_3196,N_3095);
xnor U3273 (N_3273,N_3122,N_3193);
and U3274 (N_3274,N_3137,N_3136);
or U3275 (N_3275,N_3078,N_3145);
and U3276 (N_3276,N_3099,N_3068);
xnor U3277 (N_3277,N_3083,N_3111);
nor U3278 (N_3278,N_3077,N_3177);
nor U3279 (N_3279,N_3140,N_3135);
nor U3280 (N_3280,N_3130,N_3128);
and U3281 (N_3281,N_3156,N_3178);
nor U3282 (N_3282,N_3115,N_3093);
nor U3283 (N_3283,N_3058,N_3114);
nor U3284 (N_3284,N_3164,N_3059);
nor U3285 (N_3285,N_3085,N_3190);
and U3286 (N_3286,N_3162,N_3052);
xor U3287 (N_3287,N_3081,N_3107);
xor U3288 (N_3288,N_3118,N_3176);
nand U3289 (N_3289,N_3173,N_3140);
nand U3290 (N_3290,N_3096,N_3137);
nand U3291 (N_3291,N_3126,N_3139);
nor U3292 (N_3292,N_3078,N_3129);
nand U3293 (N_3293,N_3158,N_3092);
or U3294 (N_3294,N_3043,N_3109);
nand U3295 (N_3295,N_3075,N_3186);
xnor U3296 (N_3296,N_3180,N_3043);
nand U3297 (N_3297,N_3128,N_3179);
nor U3298 (N_3298,N_3155,N_3143);
or U3299 (N_3299,N_3155,N_3110);
nand U3300 (N_3300,N_3192,N_3122);
nand U3301 (N_3301,N_3127,N_3183);
and U3302 (N_3302,N_3097,N_3154);
nor U3303 (N_3303,N_3182,N_3067);
xor U3304 (N_3304,N_3095,N_3185);
and U3305 (N_3305,N_3082,N_3134);
xor U3306 (N_3306,N_3168,N_3103);
and U3307 (N_3307,N_3122,N_3043);
and U3308 (N_3308,N_3168,N_3147);
nand U3309 (N_3309,N_3108,N_3069);
xnor U3310 (N_3310,N_3065,N_3134);
nor U3311 (N_3311,N_3124,N_3071);
nand U3312 (N_3312,N_3065,N_3128);
xnor U3313 (N_3313,N_3094,N_3090);
nand U3314 (N_3314,N_3071,N_3184);
and U3315 (N_3315,N_3109,N_3199);
nor U3316 (N_3316,N_3173,N_3191);
or U3317 (N_3317,N_3169,N_3148);
and U3318 (N_3318,N_3090,N_3162);
xor U3319 (N_3319,N_3059,N_3044);
nand U3320 (N_3320,N_3125,N_3159);
nand U3321 (N_3321,N_3065,N_3122);
nand U3322 (N_3322,N_3180,N_3191);
or U3323 (N_3323,N_3151,N_3149);
xor U3324 (N_3324,N_3103,N_3182);
and U3325 (N_3325,N_3073,N_3128);
nand U3326 (N_3326,N_3170,N_3078);
nor U3327 (N_3327,N_3160,N_3042);
xor U3328 (N_3328,N_3120,N_3040);
or U3329 (N_3329,N_3190,N_3176);
nor U3330 (N_3330,N_3094,N_3067);
nand U3331 (N_3331,N_3065,N_3108);
nand U3332 (N_3332,N_3070,N_3146);
and U3333 (N_3333,N_3057,N_3051);
xnor U3334 (N_3334,N_3073,N_3040);
xor U3335 (N_3335,N_3070,N_3178);
or U3336 (N_3336,N_3049,N_3136);
nor U3337 (N_3337,N_3164,N_3090);
or U3338 (N_3338,N_3134,N_3170);
nor U3339 (N_3339,N_3165,N_3087);
nand U3340 (N_3340,N_3051,N_3065);
or U3341 (N_3341,N_3198,N_3062);
nand U3342 (N_3342,N_3186,N_3089);
or U3343 (N_3343,N_3047,N_3117);
nand U3344 (N_3344,N_3097,N_3046);
and U3345 (N_3345,N_3152,N_3078);
and U3346 (N_3346,N_3119,N_3074);
and U3347 (N_3347,N_3158,N_3185);
or U3348 (N_3348,N_3143,N_3099);
nand U3349 (N_3349,N_3089,N_3042);
or U3350 (N_3350,N_3177,N_3064);
and U3351 (N_3351,N_3089,N_3088);
or U3352 (N_3352,N_3120,N_3154);
nor U3353 (N_3353,N_3188,N_3194);
nor U3354 (N_3354,N_3048,N_3098);
or U3355 (N_3355,N_3085,N_3040);
nand U3356 (N_3356,N_3054,N_3128);
nor U3357 (N_3357,N_3123,N_3114);
and U3358 (N_3358,N_3175,N_3117);
nor U3359 (N_3359,N_3160,N_3131);
xor U3360 (N_3360,N_3225,N_3269);
and U3361 (N_3361,N_3342,N_3311);
nor U3362 (N_3362,N_3237,N_3253);
or U3363 (N_3363,N_3350,N_3344);
nor U3364 (N_3364,N_3345,N_3259);
xor U3365 (N_3365,N_3294,N_3288);
xnor U3366 (N_3366,N_3291,N_3270);
or U3367 (N_3367,N_3213,N_3250);
xor U3368 (N_3368,N_3347,N_3310);
and U3369 (N_3369,N_3289,N_3333);
and U3370 (N_3370,N_3275,N_3290);
nand U3371 (N_3371,N_3292,N_3234);
or U3372 (N_3372,N_3260,N_3331);
or U3373 (N_3373,N_3206,N_3302);
and U3374 (N_3374,N_3305,N_3231);
xor U3375 (N_3375,N_3351,N_3352);
nand U3376 (N_3376,N_3319,N_3271);
nor U3377 (N_3377,N_3293,N_3203);
nor U3378 (N_3378,N_3211,N_3249);
xnor U3379 (N_3379,N_3278,N_3210);
xor U3380 (N_3380,N_3287,N_3279);
xor U3381 (N_3381,N_3258,N_3348);
xor U3382 (N_3382,N_3264,N_3245);
or U3383 (N_3383,N_3318,N_3228);
nand U3384 (N_3384,N_3248,N_3208);
nor U3385 (N_3385,N_3357,N_3215);
or U3386 (N_3386,N_3358,N_3227);
xnor U3387 (N_3387,N_3327,N_3354);
nor U3388 (N_3388,N_3246,N_3286);
and U3389 (N_3389,N_3243,N_3336);
nor U3390 (N_3390,N_3209,N_3359);
nand U3391 (N_3391,N_3267,N_3244);
nand U3392 (N_3392,N_3316,N_3337);
nor U3393 (N_3393,N_3326,N_3321);
xnor U3394 (N_3394,N_3315,N_3202);
and U3395 (N_3395,N_3282,N_3340);
nor U3396 (N_3396,N_3328,N_3299);
or U3397 (N_3397,N_3221,N_3251);
and U3398 (N_3398,N_3273,N_3303);
or U3399 (N_3399,N_3307,N_3236);
and U3400 (N_3400,N_3223,N_3281);
and U3401 (N_3401,N_3266,N_3200);
nor U3402 (N_3402,N_3317,N_3207);
and U3403 (N_3403,N_3323,N_3205);
and U3404 (N_3404,N_3296,N_3226);
and U3405 (N_3405,N_3263,N_3309);
nor U3406 (N_3406,N_3339,N_3283);
xnor U3407 (N_3407,N_3308,N_3300);
and U3408 (N_3408,N_3272,N_3220);
and U3409 (N_3409,N_3346,N_3274);
and U3410 (N_3410,N_3261,N_3295);
nand U3411 (N_3411,N_3301,N_3276);
or U3412 (N_3412,N_3284,N_3232);
xor U3413 (N_3413,N_3239,N_3353);
nor U3414 (N_3414,N_3338,N_3322);
nor U3415 (N_3415,N_3298,N_3241);
and U3416 (N_3416,N_3280,N_3238);
nand U3417 (N_3417,N_3306,N_3335);
and U3418 (N_3418,N_3240,N_3324);
nand U3419 (N_3419,N_3320,N_3235);
xnor U3420 (N_3420,N_3212,N_3204);
xnor U3421 (N_3421,N_3297,N_3254);
nand U3422 (N_3422,N_3229,N_3277);
nor U3423 (N_3423,N_3252,N_3230);
xnor U3424 (N_3424,N_3334,N_3257);
and U3425 (N_3425,N_3341,N_3219);
nor U3426 (N_3426,N_3262,N_3356);
and U3427 (N_3427,N_3329,N_3214);
and U3428 (N_3428,N_3314,N_3313);
xor U3429 (N_3429,N_3332,N_3256);
nor U3430 (N_3430,N_3217,N_3285);
xor U3431 (N_3431,N_3349,N_3247);
nand U3432 (N_3432,N_3312,N_3355);
xor U3433 (N_3433,N_3201,N_3265);
xnor U3434 (N_3434,N_3218,N_3268);
and U3435 (N_3435,N_3325,N_3242);
or U3436 (N_3436,N_3233,N_3222);
xor U3437 (N_3437,N_3330,N_3224);
nor U3438 (N_3438,N_3343,N_3216);
and U3439 (N_3439,N_3304,N_3255);
and U3440 (N_3440,N_3316,N_3227);
nand U3441 (N_3441,N_3267,N_3291);
nand U3442 (N_3442,N_3311,N_3279);
nor U3443 (N_3443,N_3348,N_3260);
nor U3444 (N_3444,N_3247,N_3342);
xor U3445 (N_3445,N_3318,N_3316);
nand U3446 (N_3446,N_3344,N_3262);
and U3447 (N_3447,N_3243,N_3218);
or U3448 (N_3448,N_3230,N_3216);
or U3449 (N_3449,N_3357,N_3339);
and U3450 (N_3450,N_3239,N_3229);
or U3451 (N_3451,N_3212,N_3227);
xor U3452 (N_3452,N_3276,N_3286);
nor U3453 (N_3453,N_3204,N_3218);
nor U3454 (N_3454,N_3290,N_3351);
or U3455 (N_3455,N_3238,N_3303);
or U3456 (N_3456,N_3247,N_3225);
and U3457 (N_3457,N_3319,N_3247);
nor U3458 (N_3458,N_3346,N_3344);
nor U3459 (N_3459,N_3346,N_3259);
nand U3460 (N_3460,N_3238,N_3339);
and U3461 (N_3461,N_3330,N_3213);
nand U3462 (N_3462,N_3288,N_3330);
nor U3463 (N_3463,N_3331,N_3283);
and U3464 (N_3464,N_3240,N_3264);
xor U3465 (N_3465,N_3219,N_3302);
nor U3466 (N_3466,N_3255,N_3202);
and U3467 (N_3467,N_3234,N_3329);
xnor U3468 (N_3468,N_3280,N_3228);
xnor U3469 (N_3469,N_3296,N_3274);
nor U3470 (N_3470,N_3354,N_3251);
nand U3471 (N_3471,N_3315,N_3343);
nand U3472 (N_3472,N_3322,N_3218);
and U3473 (N_3473,N_3306,N_3351);
and U3474 (N_3474,N_3231,N_3346);
and U3475 (N_3475,N_3321,N_3277);
xnor U3476 (N_3476,N_3291,N_3245);
xor U3477 (N_3477,N_3358,N_3218);
or U3478 (N_3478,N_3265,N_3271);
nand U3479 (N_3479,N_3205,N_3219);
nor U3480 (N_3480,N_3254,N_3300);
and U3481 (N_3481,N_3333,N_3227);
or U3482 (N_3482,N_3223,N_3350);
and U3483 (N_3483,N_3357,N_3223);
nand U3484 (N_3484,N_3307,N_3345);
and U3485 (N_3485,N_3300,N_3227);
nand U3486 (N_3486,N_3249,N_3215);
and U3487 (N_3487,N_3292,N_3233);
nor U3488 (N_3488,N_3279,N_3225);
nor U3489 (N_3489,N_3265,N_3277);
or U3490 (N_3490,N_3300,N_3307);
nand U3491 (N_3491,N_3209,N_3247);
nor U3492 (N_3492,N_3226,N_3208);
or U3493 (N_3493,N_3205,N_3295);
nor U3494 (N_3494,N_3264,N_3339);
nor U3495 (N_3495,N_3213,N_3280);
nor U3496 (N_3496,N_3233,N_3274);
or U3497 (N_3497,N_3277,N_3235);
and U3498 (N_3498,N_3310,N_3219);
nor U3499 (N_3499,N_3331,N_3316);
nor U3500 (N_3500,N_3320,N_3295);
xnor U3501 (N_3501,N_3319,N_3229);
nand U3502 (N_3502,N_3321,N_3355);
and U3503 (N_3503,N_3349,N_3298);
or U3504 (N_3504,N_3263,N_3265);
xor U3505 (N_3505,N_3275,N_3205);
nor U3506 (N_3506,N_3201,N_3318);
nand U3507 (N_3507,N_3202,N_3227);
nand U3508 (N_3508,N_3355,N_3309);
and U3509 (N_3509,N_3207,N_3333);
and U3510 (N_3510,N_3247,N_3283);
and U3511 (N_3511,N_3328,N_3247);
xnor U3512 (N_3512,N_3271,N_3314);
xor U3513 (N_3513,N_3200,N_3210);
and U3514 (N_3514,N_3294,N_3329);
or U3515 (N_3515,N_3244,N_3210);
xnor U3516 (N_3516,N_3326,N_3300);
nand U3517 (N_3517,N_3358,N_3274);
and U3518 (N_3518,N_3210,N_3214);
or U3519 (N_3519,N_3241,N_3248);
nand U3520 (N_3520,N_3463,N_3455);
xnor U3521 (N_3521,N_3385,N_3389);
and U3522 (N_3522,N_3410,N_3494);
or U3523 (N_3523,N_3497,N_3404);
xnor U3524 (N_3524,N_3440,N_3454);
xor U3525 (N_3525,N_3437,N_3450);
and U3526 (N_3526,N_3444,N_3369);
xnor U3527 (N_3527,N_3431,N_3516);
xor U3528 (N_3528,N_3393,N_3400);
nand U3529 (N_3529,N_3408,N_3403);
xnor U3530 (N_3530,N_3387,N_3451);
nand U3531 (N_3531,N_3447,N_3501);
xnor U3532 (N_3532,N_3378,N_3519);
and U3533 (N_3533,N_3390,N_3492);
and U3534 (N_3534,N_3443,N_3413);
nand U3535 (N_3535,N_3513,N_3414);
and U3536 (N_3536,N_3517,N_3491);
nor U3537 (N_3537,N_3479,N_3461);
and U3538 (N_3538,N_3504,N_3490);
and U3539 (N_3539,N_3379,N_3417);
or U3540 (N_3540,N_3367,N_3416);
and U3541 (N_3541,N_3406,N_3421);
or U3542 (N_3542,N_3496,N_3449);
nor U3543 (N_3543,N_3388,N_3398);
or U3544 (N_3544,N_3372,N_3481);
xnor U3545 (N_3545,N_3361,N_3475);
xor U3546 (N_3546,N_3473,N_3508);
and U3547 (N_3547,N_3493,N_3433);
nor U3548 (N_3548,N_3515,N_3459);
nor U3549 (N_3549,N_3370,N_3384);
nor U3550 (N_3550,N_3395,N_3422);
xor U3551 (N_3551,N_3482,N_3364);
and U3552 (N_3552,N_3411,N_3471);
and U3553 (N_3553,N_3442,N_3412);
xnor U3554 (N_3554,N_3418,N_3474);
and U3555 (N_3555,N_3456,N_3396);
nor U3556 (N_3556,N_3377,N_3480);
nor U3557 (N_3557,N_3363,N_3506);
nor U3558 (N_3558,N_3509,N_3446);
xor U3559 (N_3559,N_3477,N_3430);
xnor U3560 (N_3560,N_3436,N_3429);
xnor U3561 (N_3561,N_3469,N_3498);
and U3562 (N_3562,N_3453,N_3362);
and U3563 (N_3563,N_3391,N_3434);
xnor U3564 (N_3564,N_3420,N_3438);
xor U3565 (N_3565,N_3374,N_3427);
nor U3566 (N_3566,N_3483,N_3448);
nor U3567 (N_3567,N_3476,N_3441);
xnor U3568 (N_3568,N_3478,N_3486);
xor U3569 (N_3569,N_3465,N_3472);
nor U3570 (N_3570,N_3485,N_3383);
and U3571 (N_3571,N_3488,N_3360);
nand U3572 (N_3572,N_3392,N_3376);
or U3573 (N_3573,N_3425,N_3401);
or U3574 (N_3574,N_3510,N_3381);
nor U3575 (N_3575,N_3458,N_3382);
nand U3576 (N_3576,N_3435,N_3415);
and U3577 (N_3577,N_3495,N_3445);
nand U3578 (N_3578,N_3466,N_3409);
nor U3579 (N_3579,N_3507,N_3375);
nand U3580 (N_3580,N_3428,N_3405);
nand U3581 (N_3581,N_3424,N_3365);
nand U3582 (N_3582,N_3464,N_3503);
nand U3583 (N_3583,N_3484,N_3419);
nand U3584 (N_3584,N_3462,N_3373);
or U3585 (N_3585,N_3386,N_3432);
nand U3586 (N_3586,N_3487,N_3511);
nand U3587 (N_3587,N_3505,N_3460);
nand U3588 (N_3588,N_3394,N_3518);
xor U3589 (N_3589,N_3514,N_3402);
or U3590 (N_3590,N_3426,N_3407);
nand U3591 (N_3591,N_3452,N_3489);
nor U3592 (N_3592,N_3457,N_3468);
xor U3593 (N_3593,N_3397,N_3500);
or U3594 (N_3594,N_3439,N_3380);
nand U3595 (N_3595,N_3366,N_3423);
or U3596 (N_3596,N_3399,N_3499);
or U3597 (N_3597,N_3467,N_3368);
nand U3598 (N_3598,N_3502,N_3512);
nor U3599 (N_3599,N_3470,N_3371);
or U3600 (N_3600,N_3502,N_3465);
xor U3601 (N_3601,N_3424,N_3517);
nor U3602 (N_3602,N_3418,N_3368);
xnor U3603 (N_3603,N_3441,N_3422);
nor U3604 (N_3604,N_3365,N_3467);
xor U3605 (N_3605,N_3458,N_3403);
nand U3606 (N_3606,N_3447,N_3391);
nor U3607 (N_3607,N_3372,N_3434);
nand U3608 (N_3608,N_3467,N_3367);
nor U3609 (N_3609,N_3467,N_3495);
and U3610 (N_3610,N_3432,N_3431);
nor U3611 (N_3611,N_3457,N_3519);
or U3612 (N_3612,N_3465,N_3468);
or U3613 (N_3613,N_3421,N_3508);
nor U3614 (N_3614,N_3450,N_3388);
nor U3615 (N_3615,N_3418,N_3519);
and U3616 (N_3616,N_3456,N_3491);
and U3617 (N_3617,N_3493,N_3424);
nor U3618 (N_3618,N_3496,N_3419);
nor U3619 (N_3619,N_3458,N_3481);
or U3620 (N_3620,N_3487,N_3471);
nand U3621 (N_3621,N_3491,N_3407);
or U3622 (N_3622,N_3488,N_3452);
nand U3623 (N_3623,N_3457,N_3418);
and U3624 (N_3624,N_3443,N_3470);
nor U3625 (N_3625,N_3506,N_3384);
xnor U3626 (N_3626,N_3365,N_3476);
and U3627 (N_3627,N_3450,N_3511);
or U3628 (N_3628,N_3413,N_3445);
or U3629 (N_3629,N_3508,N_3416);
and U3630 (N_3630,N_3455,N_3391);
or U3631 (N_3631,N_3449,N_3378);
nor U3632 (N_3632,N_3429,N_3497);
nor U3633 (N_3633,N_3423,N_3389);
nor U3634 (N_3634,N_3374,N_3493);
xnor U3635 (N_3635,N_3415,N_3380);
or U3636 (N_3636,N_3436,N_3400);
nand U3637 (N_3637,N_3366,N_3410);
nor U3638 (N_3638,N_3472,N_3457);
and U3639 (N_3639,N_3462,N_3402);
nand U3640 (N_3640,N_3419,N_3466);
or U3641 (N_3641,N_3431,N_3401);
xnor U3642 (N_3642,N_3501,N_3475);
and U3643 (N_3643,N_3394,N_3422);
and U3644 (N_3644,N_3367,N_3430);
xor U3645 (N_3645,N_3439,N_3514);
nand U3646 (N_3646,N_3461,N_3398);
nor U3647 (N_3647,N_3515,N_3383);
nand U3648 (N_3648,N_3442,N_3362);
nand U3649 (N_3649,N_3409,N_3398);
and U3650 (N_3650,N_3462,N_3363);
and U3651 (N_3651,N_3462,N_3485);
nor U3652 (N_3652,N_3456,N_3431);
and U3653 (N_3653,N_3450,N_3491);
xor U3654 (N_3654,N_3446,N_3370);
and U3655 (N_3655,N_3494,N_3445);
and U3656 (N_3656,N_3407,N_3460);
nand U3657 (N_3657,N_3512,N_3504);
nor U3658 (N_3658,N_3371,N_3505);
nand U3659 (N_3659,N_3514,N_3476);
and U3660 (N_3660,N_3427,N_3425);
and U3661 (N_3661,N_3386,N_3456);
nand U3662 (N_3662,N_3475,N_3490);
xor U3663 (N_3663,N_3472,N_3372);
xnor U3664 (N_3664,N_3421,N_3481);
xor U3665 (N_3665,N_3392,N_3460);
and U3666 (N_3666,N_3439,N_3512);
and U3667 (N_3667,N_3439,N_3462);
xnor U3668 (N_3668,N_3383,N_3440);
xor U3669 (N_3669,N_3399,N_3502);
nand U3670 (N_3670,N_3479,N_3500);
and U3671 (N_3671,N_3365,N_3433);
or U3672 (N_3672,N_3453,N_3374);
nand U3673 (N_3673,N_3460,N_3378);
xor U3674 (N_3674,N_3487,N_3378);
nor U3675 (N_3675,N_3384,N_3477);
or U3676 (N_3676,N_3509,N_3424);
and U3677 (N_3677,N_3468,N_3404);
nand U3678 (N_3678,N_3394,N_3501);
nand U3679 (N_3679,N_3459,N_3462);
and U3680 (N_3680,N_3639,N_3597);
or U3681 (N_3681,N_3592,N_3544);
nand U3682 (N_3682,N_3554,N_3665);
and U3683 (N_3683,N_3525,N_3574);
and U3684 (N_3684,N_3651,N_3591);
nor U3685 (N_3685,N_3631,N_3578);
xnor U3686 (N_3686,N_3534,N_3657);
and U3687 (N_3687,N_3600,N_3625);
nor U3688 (N_3688,N_3543,N_3527);
or U3689 (N_3689,N_3618,N_3595);
or U3690 (N_3690,N_3610,N_3523);
or U3691 (N_3691,N_3620,N_3627);
nor U3692 (N_3692,N_3557,N_3561);
nand U3693 (N_3693,N_3535,N_3575);
and U3694 (N_3694,N_3529,N_3643);
or U3695 (N_3695,N_3577,N_3632);
xnor U3696 (N_3696,N_3599,N_3616);
nand U3697 (N_3697,N_3565,N_3677);
or U3698 (N_3698,N_3556,N_3559);
and U3699 (N_3699,N_3640,N_3552);
nand U3700 (N_3700,N_3650,N_3536);
xor U3701 (N_3701,N_3545,N_3568);
nor U3702 (N_3702,N_3675,N_3562);
nor U3703 (N_3703,N_3629,N_3564);
nand U3704 (N_3704,N_3621,N_3602);
and U3705 (N_3705,N_3623,N_3652);
nand U3706 (N_3706,N_3641,N_3569);
xor U3707 (N_3707,N_3678,N_3603);
or U3708 (N_3708,N_3645,N_3630);
and U3709 (N_3709,N_3670,N_3526);
or U3710 (N_3710,N_3663,N_3679);
nor U3711 (N_3711,N_3537,N_3533);
nand U3712 (N_3712,N_3522,N_3653);
xnor U3713 (N_3713,N_3667,N_3606);
nor U3714 (N_3714,N_3584,N_3560);
and U3715 (N_3715,N_3648,N_3676);
or U3716 (N_3716,N_3570,N_3656);
nor U3717 (N_3717,N_3538,N_3634);
or U3718 (N_3718,N_3541,N_3540);
nor U3719 (N_3719,N_3531,N_3674);
nand U3720 (N_3720,N_3590,N_3671);
and U3721 (N_3721,N_3587,N_3598);
nor U3722 (N_3722,N_3547,N_3580);
nand U3723 (N_3723,N_3572,N_3649);
or U3724 (N_3724,N_3548,N_3614);
and U3725 (N_3725,N_3609,N_3601);
nand U3726 (N_3726,N_3642,N_3532);
xor U3727 (N_3727,N_3528,N_3635);
xnor U3728 (N_3728,N_3655,N_3567);
or U3729 (N_3729,N_3636,N_3551);
xnor U3730 (N_3730,N_3583,N_3542);
and U3731 (N_3731,N_3573,N_3662);
nor U3732 (N_3732,N_3576,N_3608);
or U3733 (N_3733,N_3617,N_3571);
or U3734 (N_3734,N_3638,N_3624);
or U3735 (N_3735,N_3612,N_3646);
xnor U3736 (N_3736,N_3654,N_3604);
nand U3737 (N_3737,N_3669,N_3647);
or U3738 (N_3738,N_3586,N_3539);
or U3739 (N_3739,N_3673,N_3579);
and U3740 (N_3740,N_3550,N_3521);
nor U3741 (N_3741,N_3622,N_3605);
nand U3742 (N_3742,N_3637,N_3660);
and U3743 (N_3743,N_3661,N_3615);
xnor U3744 (N_3744,N_3582,N_3644);
xor U3745 (N_3745,N_3581,N_3659);
nor U3746 (N_3746,N_3596,N_3546);
and U3747 (N_3747,N_3668,N_3628);
nor U3748 (N_3748,N_3664,N_3672);
and U3749 (N_3749,N_3553,N_3530);
and U3750 (N_3750,N_3588,N_3520);
nor U3751 (N_3751,N_3594,N_3633);
nor U3752 (N_3752,N_3611,N_3585);
xor U3753 (N_3753,N_3549,N_3613);
and U3754 (N_3754,N_3563,N_3626);
nand U3755 (N_3755,N_3666,N_3558);
xnor U3756 (N_3756,N_3658,N_3593);
xnor U3757 (N_3757,N_3524,N_3607);
and U3758 (N_3758,N_3555,N_3619);
nor U3759 (N_3759,N_3589,N_3566);
nor U3760 (N_3760,N_3627,N_3602);
nand U3761 (N_3761,N_3581,N_3543);
nor U3762 (N_3762,N_3566,N_3595);
nand U3763 (N_3763,N_3674,N_3588);
xnor U3764 (N_3764,N_3581,N_3523);
and U3765 (N_3765,N_3532,N_3522);
nand U3766 (N_3766,N_3563,N_3568);
nor U3767 (N_3767,N_3635,N_3618);
nand U3768 (N_3768,N_3607,N_3661);
xnor U3769 (N_3769,N_3655,N_3669);
and U3770 (N_3770,N_3590,N_3651);
nand U3771 (N_3771,N_3643,N_3645);
nor U3772 (N_3772,N_3539,N_3605);
nor U3773 (N_3773,N_3556,N_3670);
nand U3774 (N_3774,N_3572,N_3582);
xnor U3775 (N_3775,N_3571,N_3631);
or U3776 (N_3776,N_3612,N_3585);
nand U3777 (N_3777,N_3661,N_3528);
and U3778 (N_3778,N_3580,N_3564);
nor U3779 (N_3779,N_3643,N_3521);
and U3780 (N_3780,N_3619,N_3662);
nor U3781 (N_3781,N_3643,N_3524);
or U3782 (N_3782,N_3532,N_3540);
or U3783 (N_3783,N_3670,N_3648);
or U3784 (N_3784,N_3526,N_3659);
or U3785 (N_3785,N_3625,N_3618);
xnor U3786 (N_3786,N_3573,N_3599);
xor U3787 (N_3787,N_3635,N_3662);
xnor U3788 (N_3788,N_3604,N_3668);
nor U3789 (N_3789,N_3529,N_3661);
nor U3790 (N_3790,N_3581,N_3563);
xnor U3791 (N_3791,N_3613,N_3595);
xnor U3792 (N_3792,N_3521,N_3669);
and U3793 (N_3793,N_3677,N_3609);
xor U3794 (N_3794,N_3552,N_3624);
xnor U3795 (N_3795,N_3566,N_3559);
nor U3796 (N_3796,N_3661,N_3574);
or U3797 (N_3797,N_3562,N_3558);
nor U3798 (N_3798,N_3610,N_3639);
nor U3799 (N_3799,N_3607,N_3619);
xor U3800 (N_3800,N_3575,N_3673);
nor U3801 (N_3801,N_3629,N_3610);
or U3802 (N_3802,N_3635,N_3566);
xor U3803 (N_3803,N_3557,N_3548);
nor U3804 (N_3804,N_3595,N_3676);
nand U3805 (N_3805,N_3564,N_3605);
xor U3806 (N_3806,N_3645,N_3625);
xor U3807 (N_3807,N_3582,N_3645);
nor U3808 (N_3808,N_3609,N_3527);
nor U3809 (N_3809,N_3520,N_3648);
and U3810 (N_3810,N_3665,N_3625);
nand U3811 (N_3811,N_3556,N_3606);
or U3812 (N_3812,N_3651,N_3659);
or U3813 (N_3813,N_3617,N_3663);
and U3814 (N_3814,N_3612,N_3555);
or U3815 (N_3815,N_3632,N_3672);
nand U3816 (N_3816,N_3651,N_3655);
or U3817 (N_3817,N_3600,N_3610);
nand U3818 (N_3818,N_3561,N_3573);
and U3819 (N_3819,N_3637,N_3604);
nor U3820 (N_3820,N_3648,N_3533);
nand U3821 (N_3821,N_3560,N_3665);
nor U3822 (N_3822,N_3617,N_3629);
nand U3823 (N_3823,N_3540,N_3564);
and U3824 (N_3824,N_3522,N_3541);
and U3825 (N_3825,N_3541,N_3662);
nor U3826 (N_3826,N_3558,N_3677);
nand U3827 (N_3827,N_3562,N_3587);
xor U3828 (N_3828,N_3592,N_3588);
or U3829 (N_3829,N_3631,N_3547);
and U3830 (N_3830,N_3560,N_3604);
and U3831 (N_3831,N_3534,N_3599);
or U3832 (N_3832,N_3547,N_3539);
nor U3833 (N_3833,N_3569,N_3578);
xnor U3834 (N_3834,N_3572,N_3670);
xnor U3835 (N_3835,N_3585,N_3649);
nand U3836 (N_3836,N_3654,N_3644);
nor U3837 (N_3837,N_3537,N_3539);
or U3838 (N_3838,N_3595,N_3530);
nand U3839 (N_3839,N_3591,N_3657);
and U3840 (N_3840,N_3831,N_3743);
or U3841 (N_3841,N_3832,N_3742);
nor U3842 (N_3842,N_3727,N_3732);
nor U3843 (N_3843,N_3797,N_3747);
nand U3844 (N_3844,N_3781,N_3691);
nand U3845 (N_3845,N_3765,N_3768);
nor U3846 (N_3846,N_3839,N_3821);
nor U3847 (N_3847,N_3750,N_3681);
and U3848 (N_3848,N_3739,N_3769);
and U3849 (N_3849,N_3751,N_3779);
nand U3850 (N_3850,N_3760,N_3692);
nor U3851 (N_3851,N_3787,N_3726);
xnor U3852 (N_3852,N_3753,N_3687);
or U3853 (N_3853,N_3680,N_3702);
nor U3854 (N_3854,N_3826,N_3708);
nand U3855 (N_3855,N_3686,N_3764);
nor U3856 (N_3856,N_3761,N_3685);
or U3857 (N_3857,N_3815,N_3799);
or U3858 (N_3858,N_3706,N_3705);
or U3859 (N_3859,N_3715,N_3804);
and U3860 (N_3860,N_3837,N_3794);
nor U3861 (N_3861,N_3713,N_3721);
or U3862 (N_3862,N_3682,N_3836);
or U3863 (N_3863,N_3694,N_3735);
nor U3864 (N_3864,N_3693,N_3683);
xor U3865 (N_3865,N_3766,N_3699);
nor U3866 (N_3866,N_3783,N_3785);
xor U3867 (N_3867,N_3824,N_3806);
nor U3868 (N_3868,N_3688,N_3711);
and U3869 (N_3869,N_3734,N_3812);
or U3870 (N_3870,N_3701,N_3774);
or U3871 (N_3871,N_3801,N_3723);
nand U3872 (N_3872,N_3767,N_3823);
xnor U3873 (N_3873,N_3703,N_3704);
nor U3874 (N_3874,N_3717,N_3745);
nor U3875 (N_3875,N_3762,N_3825);
nor U3876 (N_3876,N_3814,N_3773);
or U3877 (N_3877,N_3754,N_3782);
nor U3878 (N_3878,N_3789,N_3811);
nor U3879 (N_3879,N_3808,N_3802);
and U3880 (N_3880,N_3698,N_3712);
and U3881 (N_3881,N_3736,N_3755);
and U3882 (N_3882,N_3738,N_3813);
and U3883 (N_3883,N_3722,N_3796);
and U3884 (N_3884,N_3700,N_3756);
nand U3885 (N_3885,N_3780,N_3778);
nor U3886 (N_3886,N_3795,N_3791);
or U3887 (N_3887,N_3748,N_3809);
xnor U3888 (N_3888,N_3807,N_3752);
nand U3889 (N_3889,N_3740,N_3805);
xnor U3890 (N_3890,N_3790,N_3757);
nor U3891 (N_3891,N_3835,N_3720);
and U3892 (N_3892,N_3776,N_3749);
nand U3893 (N_3893,N_3725,N_3793);
nand U3894 (N_3894,N_3770,N_3684);
nor U3895 (N_3895,N_3758,N_3827);
or U3896 (N_3896,N_3800,N_3690);
nor U3897 (N_3897,N_3830,N_3689);
or U3898 (N_3898,N_3772,N_3817);
nand U3899 (N_3899,N_3771,N_3834);
xor U3900 (N_3900,N_3829,N_3709);
xnor U3901 (N_3901,N_3737,N_3810);
xnor U3902 (N_3902,N_3833,N_3710);
xor U3903 (N_3903,N_3719,N_3707);
and U3904 (N_3904,N_3784,N_3816);
or U3905 (N_3905,N_3818,N_3822);
and U3906 (N_3906,N_3786,N_3838);
nor U3907 (N_3907,N_3828,N_3803);
or U3908 (N_3908,N_3733,N_3714);
nor U3909 (N_3909,N_3741,N_3695);
or U3910 (N_3910,N_3759,N_3730);
nand U3911 (N_3911,N_3716,N_3777);
nand U3912 (N_3912,N_3729,N_3798);
xnor U3913 (N_3913,N_3718,N_3697);
nor U3914 (N_3914,N_3744,N_3819);
and U3915 (N_3915,N_3728,N_3775);
nor U3916 (N_3916,N_3820,N_3731);
or U3917 (N_3917,N_3696,N_3792);
xnor U3918 (N_3918,N_3746,N_3763);
nand U3919 (N_3919,N_3788,N_3724);
nand U3920 (N_3920,N_3826,N_3696);
or U3921 (N_3921,N_3701,N_3722);
or U3922 (N_3922,N_3790,N_3806);
xnor U3923 (N_3923,N_3696,N_3694);
xor U3924 (N_3924,N_3765,N_3716);
nor U3925 (N_3925,N_3715,N_3738);
or U3926 (N_3926,N_3811,N_3815);
or U3927 (N_3927,N_3740,N_3804);
and U3928 (N_3928,N_3805,N_3819);
and U3929 (N_3929,N_3716,N_3745);
nand U3930 (N_3930,N_3784,N_3771);
nor U3931 (N_3931,N_3793,N_3825);
nor U3932 (N_3932,N_3808,N_3790);
and U3933 (N_3933,N_3686,N_3726);
nor U3934 (N_3934,N_3700,N_3730);
nor U3935 (N_3935,N_3703,N_3767);
or U3936 (N_3936,N_3796,N_3687);
nand U3937 (N_3937,N_3775,N_3773);
or U3938 (N_3938,N_3810,N_3804);
xnor U3939 (N_3939,N_3719,N_3747);
and U3940 (N_3940,N_3728,N_3839);
and U3941 (N_3941,N_3804,N_3684);
nand U3942 (N_3942,N_3681,N_3831);
and U3943 (N_3943,N_3835,N_3772);
or U3944 (N_3944,N_3820,N_3780);
or U3945 (N_3945,N_3800,N_3757);
and U3946 (N_3946,N_3726,N_3799);
xnor U3947 (N_3947,N_3815,N_3722);
nand U3948 (N_3948,N_3707,N_3791);
or U3949 (N_3949,N_3715,N_3686);
and U3950 (N_3950,N_3709,N_3828);
nor U3951 (N_3951,N_3788,N_3761);
xnor U3952 (N_3952,N_3727,N_3720);
or U3953 (N_3953,N_3693,N_3682);
and U3954 (N_3954,N_3726,N_3776);
xnor U3955 (N_3955,N_3836,N_3722);
nand U3956 (N_3956,N_3742,N_3736);
nor U3957 (N_3957,N_3780,N_3792);
nand U3958 (N_3958,N_3754,N_3808);
or U3959 (N_3959,N_3824,N_3832);
and U3960 (N_3960,N_3686,N_3736);
or U3961 (N_3961,N_3691,N_3702);
nor U3962 (N_3962,N_3810,N_3694);
and U3963 (N_3963,N_3763,N_3757);
nor U3964 (N_3964,N_3700,N_3827);
xor U3965 (N_3965,N_3695,N_3716);
xor U3966 (N_3966,N_3774,N_3809);
nor U3967 (N_3967,N_3755,N_3799);
nand U3968 (N_3968,N_3731,N_3787);
nor U3969 (N_3969,N_3787,N_3729);
xnor U3970 (N_3970,N_3715,N_3786);
nand U3971 (N_3971,N_3693,N_3755);
nand U3972 (N_3972,N_3768,N_3733);
nand U3973 (N_3973,N_3756,N_3816);
xnor U3974 (N_3974,N_3710,N_3796);
nand U3975 (N_3975,N_3694,N_3682);
nand U3976 (N_3976,N_3760,N_3836);
and U3977 (N_3977,N_3825,N_3699);
nand U3978 (N_3978,N_3733,N_3782);
or U3979 (N_3979,N_3703,N_3729);
and U3980 (N_3980,N_3732,N_3820);
or U3981 (N_3981,N_3700,N_3818);
nor U3982 (N_3982,N_3743,N_3725);
and U3983 (N_3983,N_3698,N_3808);
and U3984 (N_3984,N_3683,N_3699);
and U3985 (N_3985,N_3803,N_3754);
or U3986 (N_3986,N_3803,N_3839);
and U3987 (N_3987,N_3685,N_3774);
xnor U3988 (N_3988,N_3731,N_3713);
and U3989 (N_3989,N_3779,N_3794);
and U3990 (N_3990,N_3807,N_3782);
or U3991 (N_3991,N_3829,N_3807);
and U3992 (N_3992,N_3741,N_3805);
or U3993 (N_3993,N_3684,N_3798);
nor U3994 (N_3994,N_3720,N_3729);
and U3995 (N_3995,N_3721,N_3837);
or U3996 (N_3996,N_3776,N_3760);
xnor U3997 (N_3997,N_3709,N_3766);
xor U3998 (N_3998,N_3697,N_3710);
or U3999 (N_3999,N_3705,N_3825);
nand U4000 (N_4000,N_3929,N_3934);
nor U4001 (N_4001,N_3919,N_3848);
xor U4002 (N_4002,N_3884,N_3946);
xor U4003 (N_4003,N_3882,N_3841);
nand U4004 (N_4004,N_3890,N_3977);
and U4005 (N_4005,N_3980,N_3904);
nor U4006 (N_4006,N_3849,N_3953);
nor U4007 (N_4007,N_3924,N_3976);
nand U4008 (N_4008,N_3950,N_3911);
nor U4009 (N_4009,N_3973,N_3843);
nor U4010 (N_4010,N_3966,N_3889);
or U4011 (N_4011,N_3888,N_3887);
xor U4012 (N_4012,N_3864,N_3920);
nor U4013 (N_4013,N_3931,N_3858);
nand U4014 (N_4014,N_3952,N_3925);
or U4015 (N_4015,N_3846,N_3874);
nor U4016 (N_4016,N_3989,N_3986);
and U4017 (N_4017,N_3855,N_3886);
or U4018 (N_4018,N_3939,N_3942);
nand U4019 (N_4019,N_3965,N_3972);
nand U4020 (N_4020,N_3892,N_3860);
nand U4021 (N_4021,N_3851,N_3967);
nand U4022 (N_4022,N_3932,N_3871);
xnor U4023 (N_4023,N_3913,N_3987);
or U4024 (N_4024,N_3974,N_3927);
and U4025 (N_4025,N_3970,N_3903);
nor U4026 (N_4026,N_3981,N_3964);
nand U4027 (N_4027,N_3854,N_3909);
nand U4028 (N_4028,N_3865,N_3936);
or U4029 (N_4029,N_3951,N_3945);
xnor U4030 (N_4030,N_3968,N_3940);
nor U4031 (N_4031,N_3960,N_3955);
xor U4032 (N_4032,N_3877,N_3875);
xnor U4033 (N_4033,N_3881,N_3862);
or U4034 (N_4034,N_3869,N_3961);
nand U4035 (N_4035,N_3859,N_3897);
nor U4036 (N_4036,N_3891,N_3917);
or U4037 (N_4037,N_3947,N_3856);
and U4038 (N_4038,N_3866,N_3840);
nor U4039 (N_4039,N_3908,N_3957);
or U4040 (N_4040,N_3985,N_3845);
xnor U4041 (N_4041,N_3914,N_3943);
nor U4042 (N_4042,N_3933,N_3861);
or U4043 (N_4043,N_3959,N_3906);
or U4044 (N_4044,N_3954,N_3992);
xor U4045 (N_4045,N_3844,N_3873);
and U4046 (N_4046,N_3857,N_3899);
and U4047 (N_4047,N_3993,N_3937);
nor U4048 (N_4048,N_3983,N_3979);
nand U4049 (N_4049,N_3923,N_3900);
nor U4050 (N_4050,N_3915,N_3901);
xnor U4051 (N_4051,N_3998,N_3930);
xnor U4052 (N_4052,N_3893,N_3894);
and U4053 (N_4053,N_3896,N_3921);
nor U4054 (N_4054,N_3853,N_3958);
xor U4055 (N_4055,N_3918,N_3852);
nor U4056 (N_4056,N_3928,N_3898);
nor U4057 (N_4057,N_3870,N_3948);
xor U4058 (N_4058,N_3971,N_3912);
nand U4059 (N_4059,N_3885,N_3922);
or U4060 (N_4060,N_3880,N_3876);
and U4061 (N_4061,N_3878,N_3999);
nor U4062 (N_4062,N_3969,N_3926);
nor U4063 (N_4063,N_3975,N_3938);
nand U4064 (N_4064,N_3994,N_3872);
and U4065 (N_4065,N_3990,N_3902);
xor U4066 (N_4066,N_3941,N_3978);
xor U4067 (N_4067,N_3962,N_3982);
nand U4068 (N_4068,N_3883,N_3916);
or U4069 (N_4069,N_3905,N_3944);
xnor U4070 (N_4070,N_3988,N_3956);
or U4071 (N_4071,N_3867,N_3963);
nand U4072 (N_4072,N_3847,N_3850);
xnor U4073 (N_4073,N_3991,N_3868);
nand U4074 (N_4074,N_3949,N_3842);
nor U4075 (N_4075,N_3910,N_3895);
or U4076 (N_4076,N_3879,N_3935);
xor U4077 (N_4077,N_3984,N_3995);
nor U4078 (N_4078,N_3997,N_3907);
nor U4079 (N_4079,N_3996,N_3863);
xor U4080 (N_4080,N_3885,N_3846);
and U4081 (N_4081,N_3961,N_3969);
and U4082 (N_4082,N_3946,N_3914);
nor U4083 (N_4083,N_3982,N_3942);
xnor U4084 (N_4084,N_3967,N_3843);
xnor U4085 (N_4085,N_3865,N_3983);
nand U4086 (N_4086,N_3964,N_3842);
or U4087 (N_4087,N_3927,N_3907);
and U4088 (N_4088,N_3942,N_3930);
or U4089 (N_4089,N_3961,N_3856);
xor U4090 (N_4090,N_3922,N_3943);
nor U4091 (N_4091,N_3892,N_3926);
and U4092 (N_4092,N_3930,N_3877);
or U4093 (N_4093,N_3842,N_3958);
nand U4094 (N_4094,N_3990,N_3841);
nand U4095 (N_4095,N_3967,N_3854);
xnor U4096 (N_4096,N_3872,N_3890);
and U4097 (N_4097,N_3944,N_3997);
or U4098 (N_4098,N_3881,N_3982);
nor U4099 (N_4099,N_3924,N_3959);
nand U4100 (N_4100,N_3943,N_3998);
xnor U4101 (N_4101,N_3907,N_3862);
xor U4102 (N_4102,N_3929,N_3909);
or U4103 (N_4103,N_3953,N_3888);
nand U4104 (N_4104,N_3951,N_3893);
nor U4105 (N_4105,N_3850,N_3854);
nand U4106 (N_4106,N_3881,N_3938);
nand U4107 (N_4107,N_3936,N_3964);
nor U4108 (N_4108,N_3850,N_3994);
nand U4109 (N_4109,N_3981,N_3971);
or U4110 (N_4110,N_3866,N_3925);
nor U4111 (N_4111,N_3951,N_3860);
or U4112 (N_4112,N_3955,N_3926);
and U4113 (N_4113,N_3952,N_3858);
and U4114 (N_4114,N_3891,N_3910);
nor U4115 (N_4115,N_3867,N_3899);
nor U4116 (N_4116,N_3868,N_3950);
and U4117 (N_4117,N_3993,N_3970);
xnor U4118 (N_4118,N_3870,N_3983);
nand U4119 (N_4119,N_3898,N_3847);
nor U4120 (N_4120,N_3917,N_3925);
xnor U4121 (N_4121,N_3992,N_3948);
nor U4122 (N_4122,N_3918,N_3842);
or U4123 (N_4123,N_3944,N_3931);
and U4124 (N_4124,N_3905,N_3900);
and U4125 (N_4125,N_3854,N_3980);
nand U4126 (N_4126,N_3973,N_3913);
and U4127 (N_4127,N_3945,N_3925);
and U4128 (N_4128,N_3867,N_3976);
nor U4129 (N_4129,N_3998,N_3936);
nand U4130 (N_4130,N_3930,N_3872);
or U4131 (N_4131,N_3924,N_3880);
and U4132 (N_4132,N_3969,N_3877);
nand U4133 (N_4133,N_3910,N_3921);
or U4134 (N_4134,N_3983,N_3995);
and U4135 (N_4135,N_3850,N_3915);
and U4136 (N_4136,N_3916,N_3902);
and U4137 (N_4137,N_3896,N_3931);
nor U4138 (N_4138,N_3969,N_3903);
nand U4139 (N_4139,N_3876,N_3850);
nand U4140 (N_4140,N_3982,N_3966);
or U4141 (N_4141,N_3854,N_3999);
and U4142 (N_4142,N_3992,N_3981);
and U4143 (N_4143,N_3980,N_3869);
and U4144 (N_4144,N_3920,N_3996);
or U4145 (N_4145,N_3993,N_3895);
or U4146 (N_4146,N_3861,N_3889);
or U4147 (N_4147,N_3871,N_3847);
or U4148 (N_4148,N_3958,N_3971);
nand U4149 (N_4149,N_3995,N_3884);
nor U4150 (N_4150,N_3899,N_3965);
nor U4151 (N_4151,N_3932,N_3952);
nand U4152 (N_4152,N_3997,N_3953);
or U4153 (N_4153,N_3878,N_3914);
or U4154 (N_4154,N_3999,N_3913);
nand U4155 (N_4155,N_3932,N_3930);
or U4156 (N_4156,N_3842,N_3990);
or U4157 (N_4157,N_3939,N_3965);
or U4158 (N_4158,N_3989,N_3947);
nor U4159 (N_4159,N_3934,N_3841);
and U4160 (N_4160,N_4066,N_4133);
nand U4161 (N_4161,N_4095,N_4042);
nand U4162 (N_4162,N_4143,N_4037);
xor U4163 (N_4163,N_4137,N_4138);
and U4164 (N_4164,N_4076,N_4038);
and U4165 (N_4165,N_4053,N_4086);
xor U4166 (N_4166,N_4114,N_4050);
or U4167 (N_4167,N_4052,N_4039);
or U4168 (N_4168,N_4004,N_4005);
xor U4169 (N_4169,N_4113,N_4088);
nand U4170 (N_4170,N_4067,N_4146);
nand U4171 (N_4171,N_4079,N_4156);
and U4172 (N_4172,N_4012,N_4151);
nor U4173 (N_4173,N_4158,N_4058);
nor U4174 (N_4174,N_4064,N_4069);
nor U4175 (N_4175,N_4089,N_4002);
or U4176 (N_4176,N_4071,N_4136);
or U4177 (N_4177,N_4013,N_4142);
and U4178 (N_4178,N_4027,N_4025);
and U4179 (N_4179,N_4118,N_4017);
nand U4180 (N_4180,N_4157,N_4087);
xor U4181 (N_4181,N_4129,N_4123);
and U4182 (N_4182,N_4131,N_4015);
nor U4183 (N_4183,N_4135,N_4041);
nand U4184 (N_4184,N_4081,N_4006);
and U4185 (N_4185,N_4096,N_4080);
xnor U4186 (N_4186,N_4097,N_4154);
and U4187 (N_4187,N_4044,N_4105);
or U4188 (N_4188,N_4147,N_4102);
nor U4189 (N_4189,N_4083,N_4057);
or U4190 (N_4190,N_4007,N_4024);
or U4191 (N_4191,N_4101,N_4132);
or U4192 (N_4192,N_4141,N_4120);
xor U4193 (N_4193,N_4054,N_4034);
or U4194 (N_4194,N_4001,N_4010);
xnor U4195 (N_4195,N_4103,N_4032);
and U4196 (N_4196,N_4073,N_4144);
nor U4197 (N_4197,N_4082,N_4029);
nand U4198 (N_4198,N_4127,N_4048);
nand U4199 (N_4199,N_4099,N_4085);
and U4200 (N_4200,N_4056,N_4119);
xnor U4201 (N_4201,N_4023,N_4030);
nand U4202 (N_4202,N_4026,N_4104);
xnor U4203 (N_4203,N_4060,N_4051);
nor U4204 (N_4204,N_4159,N_4070);
xnor U4205 (N_4205,N_4028,N_4074);
xnor U4206 (N_4206,N_4098,N_4112);
nand U4207 (N_4207,N_4078,N_4155);
or U4208 (N_4208,N_4106,N_4090);
and U4209 (N_4209,N_4110,N_4084);
nor U4210 (N_4210,N_4020,N_4036);
xor U4211 (N_4211,N_4016,N_4059);
nand U4212 (N_4212,N_4008,N_4062);
or U4213 (N_4213,N_4046,N_4014);
or U4214 (N_4214,N_4068,N_4108);
nand U4215 (N_4215,N_4111,N_4117);
nor U4216 (N_4216,N_4145,N_4149);
or U4217 (N_4217,N_4043,N_4018);
and U4218 (N_4218,N_4031,N_4091);
nand U4219 (N_4219,N_4035,N_4109);
and U4220 (N_4220,N_4093,N_4094);
xor U4221 (N_4221,N_4116,N_4122);
and U4222 (N_4222,N_4140,N_4011);
nand U4223 (N_4223,N_4033,N_4003);
and U4224 (N_4224,N_4072,N_4022);
and U4225 (N_4225,N_4130,N_4125);
or U4226 (N_4226,N_4040,N_4063);
or U4227 (N_4227,N_4092,N_4139);
xor U4228 (N_4228,N_4126,N_4061);
and U4229 (N_4229,N_4128,N_4077);
and U4230 (N_4230,N_4107,N_4152);
xor U4231 (N_4231,N_4115,N_4153);
nor U4232 (N_4232,N_4100,N_4148);
xnor U4233 (N_4233,N_4045,N_4021);
nor U4234 (N_4234,N_4049,N_4019);
xnor U4235 (N_4235,N_4121,N_4047);
and U4236 (N_4236,N_4065,N_4150);
nor U4237 (N_4237,N_4055,N_4000);
xnor U4238 (N_4238,N_4134,N_4075);
nand U4239 (N_4239,N_4009,N_4124);
xor U4240 (N_4240,N_4052,N_4151);
nor U4241 (N_4241,N_4066,N_4004);
xnor U4242 (N_4242,N_4001,N_4157);
and U4243 (N_4243,N_4134,N_4143);
nand U4244 (N_4244,N_4129,N_4069);
or U4245 (N_4245,N_4069,N_4083);
or U4246 (N_4246,N_4056,N_4128);
and U4247 (N_4247,N_4048,N_4003);
and U4248 (N_4248,N_4021,N_4011);
nand U4249 (N_4249,N_4138,N_4116);
or U4250 (N_4250,N_4019,N_4122);
or U4251 (N_4251,N_4137,N_4053);
and U4252 (N_4252,N_4044,N_4041);
nor U4253 (N_4253,N_4092,N_4048);
and U4254 (N_4254,N_4074,N_4018);
nor U4255 (N_4255,N_4003,N_4130);
and U4256 (N_4256,N_4004,N_4080);
or U4257 (N_4257,N_4036,N_4157);
and U4258 (N_4258,N_4137,N_4003);
or U4259 (N_4259,N_4020,N_4001);
nand U4260 (N_4260,N_4082,N_4051);
and U4261 (N_4261,N_4155,N_4087);
and U4262 (N_4262,N_4034,N_4079);
xor U4263 (N_4263,N_4032,N_4098);
nor U4264 (N_4264,N_4078,N_4070);
xnor U4265 (N_4265,N_4010,N_4072);
nand U4266 (N_4266,N_4038,N_4126);
nand U4267 (N_4267,N_4037,N_4052);
nor U4268 (N_4268,N_4123,N_4060);
xnor U4269 (N_4269,N_4045,N_4026);
and U4270 (N_4270,N_4125,N_4038);
or U4271 (N_4271,N_4108,N_4136);
nor U4272 (N_4272,N_4042,N_4064);
and U4273 (N_4273,N_4083,N_4027);
and U4274 (N_4274,N_4033,N_4025);
nor U4275 (N_4275,N_4146,N_4154);
nand U4276 (N_4276,N_4026,N_4013);
and U4277 (N_4277,N_4081,N_4119);
and U4278 (N_4278,N_4024,N_4027);
nor U4279 (N_4279,N_4129,N_4101);
xnor U4280 (N_4280,N_4112,N_4068);
xnor U4281 (N_4281,N_4077,N_4134);
or U4282 (N_4282,N_4102,N_4001);
or U4283 (N_4283,N_4037,N_4121);
xnor U4284 (N_4284,N_4140,N_4084);
or U4285 (N_4285,N_4085,N_4006);
nor U4286 (N_4286,N_4095,N_4076);
and U4287 (N_4287,N_4118,N_4152);
nor U4288 (N_4288,N_4011,N_4097);
xnor U4289 (N_4289,N_4035,N_4055);
nor U4290 (N_4290,N_4055,N_4007);
or U4291 (N_4291,N_4052,N_4032);
and U4292 (N_4292,N_4014,N_4159);
nand U4293 (N_4293,N_4082,N_4073);
nand U4294 (N_4294,N_4126,N_4091);
and U4295 (N_4295,N_4075,N_4080);
and U4296 (N_4296,N_4095,N_4014);
nand U4297 (N_4297,N_4019,N_4100);
nand U4298 (N_4298,N_4027,N_4009);
and U4299 (N_4299,N_4099,N_4094);
nor U4300 (N_4300,N_4131,N_4060);
or U4301 (N_4301,N_4107,N_4112);
nor U4302 (N_4302,N_4107,N_4093);
xnor U4303 (N_4303,N_4020,N_4140);
xor U4304 (N_4304,N_4052,N_4086);
or U4305 (N_4305,N_4076,N_4044);
nand U4306 (N_4306,N_4086,N_4060);
nor U4307 (N_4307,N_4115,N_4015);
xor U4308 (N_4308,N_4104,N_4046);
or U4309 (N_4309,N_4134,N_4122);
nand U4310 (N_4310,N_4010,N_4113);
or U4311 (N_4311,N_4007,N_4158);
nor U4312 (N_4312,N_4158,N_4017);
or U4313 (N_4313,N_4064,N_4037);
or U4314 (N_4314,N_4114,N_4111);
nand U4315 (N_4315,N_4023,N_4087);
or U4316 (N_4316,N_4140,N_4142);
and U4317 (N_4317,N_4142,N_4002);
or U4318 (N_4318,N_4088,N_4133);
xor U4319 (N_4319,N_4028,N_4143);
nor U4320 (N_4320,N_4259,N_4244);
nand U4321 (N_4321,N_4313,N_4204);
and U4322 (N_4322,N_4209,N_4247);
nor U4323 (N_4323,N_4275,N_4175);
nand U4324 (N_4324,N_4190,N_4165);
or U4325 (N_4325,N_4292,N_4220);
or U4326 (N_4326,N_4283,N_4245);
nand U4327 (N_4327,N_4201,N_4253);
or U4328 (N_4328,N_4246,N_4173);
xnor U4329 (N_4329,N_4225,N_4200);
and U4330 (N_4330,N_4298,N_4186);
xnor U4331 (N_4331,N_4314,N_4172);
nor U4332 (N_4332,N_4174,N_4315);
or U4333 (N_4333,N_4176,N_4169);
and U4334 (N_4334,N_4260,N_4181);
xnor U4335 (N_4335,N_4239,N_4316);
and U4336 (N_4336,N_4297,N_4170);
and U4337 (N_4337,N_4262,N_4163);
nor U4338 (N_4338,N_4290,N_4303);
xnor U4339 (N_4339,N_4268,N_4301);
nand U4340 (N_4340,N_4226,N_4274);
nand U4341 (N_4341,N_4212,N_4305);
xor U4342 (N_4342,N_4236,N_4276);
and U4343 (N_4343,N_4265,N_4230);
nor U4344 (N_4344,N_4307,N_4271);
nand U4345 (N_4345,N_4278,N_4289);
xor U4346 (N_4346,N_4218,N_4256);
nor U4347 (N_4347,N_4264,N_4280);
xor U4348 (N_4348,N_4224,N_4219);
or U4349 (N_4349,N_4167,N_4232);
xor U4350 (N_4350,N_4185,N_4233);
or U4351 (N_4351,N_4300,N_4319);
and U4352 (N_4352,N_4309,N_4296);
or U4353 (N_4353,N_4195,N_4310);
and U4354 (N_4354,N_4242,N_4192);
and U4355 (N_4355,N_4168,N_4272);
or U4356 (N_4356,N_4235,N_4258);
xnor U4357 (N_4357,N_4308,N_4255);
and U4358 (N_4358,N_4284,N_4248);
or U4359 (N_4359,N_4304,N_4291);
xnor U4360 (N_4360,N_4281,N_4213);
and U4361 (N_4361,N_4203,N_4288);
and U4362 (N_4362,N_4270,N_4217);
nor U4363 (N_4363,N_4227,N_4197);
and U4364 (N_4364,N_4206,N_4238);
xnor U4365 (N_4365,N_4261,N_4194);
nand U4366 (N_4366,N_4214,N_4207);
xor U4367 (N_4367,N_4180,N_4184);
or U4368 (N_4368,N_4252,N_4178);
or U4369 (N_4369,N_4299,N_4179);
and U4370 (N_4370,N_4229,N_4211);
xor U4371 (N_4371,N_4263,N_4222);
xor U4372 (N_4372,N_4221,N_4166);
xor U4373 (N_4373,N_4182,N_4277);
or U4374 (N_4374,N_4295,N_4164);
nor U4375 (N_4375,N_4210,N_4234);
nand U4376 (N_4376,N_4285,N_4311);
nand U4377 (N_4377,N_4279,N_4243);
or U4378 (N_4378,N_4241,N_4215);
or U4379 (N_4379,N_4282,N_4171);
and U4380 (N_4380,N_4161,N_4269);
xor U4381 (N_4381,N_4208,N_4293);
xor U4382 (N_4382,N_4317,N_4250);
and U4383 (N_4383,N_4254,N_4205);
nor U4384 (N_4384,N_4177,N_4187);
nand U4385 (N_4385,N_4228,N_4198);
or U4386 (N_4386,N_4199,N_4266);
and U4387 (N_4387,N_4216,N_4237);
nand U4388 (N_4388,N_4294,N_4257);
nand U4389 (N_4389,N_4286,N_4287);
nand U4390 (N_4390,N_4318,N_4306);
or U4391 (N_4391,N_4240,N_4191);
xnor U4392 (N_4392,N_4202,N_4196);
xnor U4393 (N_4393,N_4193,N_4251);
and U4394 (N_4394,N_4162,N_4189);
and U4395 (N_4395,N_4312,N_4231);
and U4396 (N_4396,N_4188,N_4223);
nand U4397 (N_4397,N_4267,N_4302);
xnor U4398 (N_4398,N_4249,N_4273);
nor U4399 (N_4399,N_4160,N_4183);
nor U4400 (N_4400,N_4273,N_4219);
and U4401 (N_4401,N_4222,N_4319);
xor U4402 (N_4402,N_4200,N_4233);
nand U4403 (N_4403,N_4291,N_4224);
nand U4404 (N_4404,N_4276,N_4241);
xnor U4405 (N_4405,N_4223,N_4182);
and U4406 (N_4406,N_4306,N_4296);
nand U4407 (N_4407,N_4252,N_4183);
nand U4408 (N_4408,N_4289,N_4231);
nor U4409 (N_4409,N_4173,N_4231);
nand U4410 (N_4410,N_4239,N_4285);
and U4411 (N_4411,N_4270,N_4277);
or U4412 (N_4412,N_4259,N_4224);
nor U4413 (N_4413,N_4226,N_4304);
or U4414 (N_4414,N_4292,N_4177);
nand U4415 (N_4415,N_4165,N_4296);
nand U4416 (N_4416,N_4266,N_4194);
xnor U4417 (N_4417,N_4230,N_4315);
xnor U4418 (N_4418,N_4245,N_4280);
nand U4419 (N_4419,N_4258,N_4277);
nand U4420 (N_4420,N_4188,N_4246);
nand U4421 (N_4421,N_4317,N_4176);
xor U4422 (N_4422,N_4293,N_4160);
nor U4423 (N_4423,N_4182,N_4165);
and U4424 (N_4424,N_4177,N_4247);
nor U4425 (N_4425,N_4247,N_4197);
nor U4426 (N_4426,N_4290,N_4197);
or U4427 (N_4427,N_4226,N_4282);
nand U4428 (N_4428,N_4193,N_4182);
or U4429 (N_4429,N_4284,N_4272);
or U4430 (N_4430,N_4298,N_4308);
or U4431 (N_4431,N_4195,N_4215);
and U4432 (N_4432,N_4175,N_4198);
and U4433 (N_4433,N_4294,N_4305);
xnor U4434 (N_4434,N_4172,N_4220);
and U4435 (N_4435,N_4306,N_4165);
nand U4436 (N_4436,N_4232,N_4161);
xor U4437 (N_4437,N_4310,N_4184);
and U4438 (N_4438,N_4246,N_4175);
xnor U4439 (N_4439,N_4201,N_4232);
nand U4440 (N_4440,N_4226,N_4291);
xor U4441 (N_4441,N_4160,N_4280);
and U4442 (N_4442,N_4163,N_4218);
and U4443 (N_4443,N_4295,N_4174);
or U4444 (N_4444,N_4173,N_4179);
nand U4445 (N_4445,N_4296,N_4189);
and U4446 (N_4446,N_4270,N_4227);
nand U4447 (N_4447,N_4295,N_4246);
nand U4448 (N_4448,N_4283,N_4195);
xnor U4449 (N_4449,N_4248,N_4279);
nor U4450 (N_4450,N_4173,N_4238);
nor U4451 (N_4451,N_4277,N_4167);
nand U4452 (N_4452,N_4211,N_4184);
nor U4453 (N_4453,N_4176,N_4184);
or U4454 (N_4454,N_4298,N_4250);
and U4455 (N_4455,N_4282,N_4169);
xor U4456 (N_4456,N_4234,N_4292);
or U4457 (N_4457,N_4255,N_4276);
nor U4458 (N_4458,N_4160,N_4255);
nand U4459 (N_4459,N_4279,N_4289);
nand U4460 (N_4460,N_4294,N_4313);
and U4461 (N_4461,N_4194,N_4214);
xor U4462 (N_4462,N_4184,N_4307);
or U4463 (N_4463,N_4305,N_4197);
xnor U4464 (N_4464,N_4188,N_4318);
xor U4465 (N_4465,N_4175,N_4209);
nand U4466 (N_4466,N_4296,N_4263);
nand U4467 (N_4467,N_4196,N_4317);
nand U4468 (N_4468,N_4241,N_4282);
nand U4469 (N_4469,N_4163,N_4299);
or U4470 (N_4470,N_4223,N_4191);
xnor U4471 (N_4471,N_4247,N_4285);
nor U4472 (N_4472,N_4222,N_4314);
and U4473 (N_4473,N_4305,N_4198);
nand U4474 (N_4474,N_4270,N_4273);
nand U4475 (N_4475,N_4277,N_4293);
nand U4476 (N_4476,N_4166,N_4199);
nor U4477 (N_4477,N_4169,N_4265);
and U4478 (N_4478,N_4199,N_4227);
nor U4479 (N_4479,N_4261,N_4241);
nand U4480 (N_4480,N_4394,N_4357);
nand U4481 (N_4481,N_4358,N_4346);
nor U4482 (N_4482,N_4439,N_4473);
or U4483 (N_4483,N_4415,N_4467);
xnor U4484 (N_4484,N_4426,N_4441);
and U4485 (N_4485,N_4339,N_4360);
or U4486 (N_4486,N_4354,N_4388);
or U4487 (N_4487,N_4455,N_4366);
nand U4488 (N_4488,N_4373,N_4361);
nor U4489 (N_4489,N_4468,N_4352);
xor U4490 (N_4490,N_4380,N_4396);
nor U4491 (N_4491,N_4343,N_4347);
xor U4492 (N_4492,N_4353,N_4436);
nand U4493 (N_4493,N_4342,N_4433);
nand U4494 (N_4494,N_4404,N_4381);
xnor U4495 (N_4495,N_4376,N_4417);
nor U4496 (N_4496,N_4398,N_4446);
nor U4497 (N_4497,N_4335,N_4400);
xor U4498 (N_4498,N_4375,N_4413);
or U4499 (N_4499,N_4359,N_4397);
nand U4500 (N_4500,N_4401,N_4372);
nor U4501 (N_4501,N_4356,N_4364);
nand U4502 (N_4502,N_4457,N_4387);
nand U4503 (N_4503,N_4419,N_4408);
xnor U4504 (N_4504,N_4466,N_4389);
nor U4505 (N_4505,N_4325,N_4423);
nor U4506 (N_4506,N_4362,N_4420);
and U4507 (N_4507,N_4355,N_4399);
and U4508 (N_4508,N_4464,N_4437);
nor U4509 (N_4509,N_4435,N_4327);
nor U4510 (N_4510,N_4418,N_4363);
and U4511 (N_4511,N_4365,N_4448);
xor U4512 (N_4512,N_4474,N_4456);
nand U4513 (N_4513,N_4458,N_4465);
nor U4514 (N_4514,N_4451,N_4333);
and U4515 (N_4515,N_4410,N_4412);
and U4516 (N_4516,N_4478,N_4348);
and U4517 (N_4517,N_4344,N_4336);
or U4518 (N_4518,N_4321,N_4383);
or U4519 (N_4519,N_4447,N_4427);
xor U4520 (N_4520,N_4322,N_4349);
nor U4521 (N_4521,N_4479,N_4445);
xnor U4522 (N_4522,N_4450,N_4460);
xnor U4523 (N_4523,N_4449,N_4328);
nand U4524 (N_4524,N_4462,N_4428);
or U4525 (N_4525,N_4326,N_4429);
xor U4526 (N_4526,N_4371,N_4320);
nor U4527 (N_4527,N_4422,N_4341);
or U4528 (N_4528,N_4367,N_4402);
and U4529 (N_4529,N_4471,N_4386);
or U4530 (N_4530,N_4351,N_4324);
nor U4531 (N_4531,N_4370,N_4390);
nand U4532 (N_4532,N_4403,N_4395);
or U4533 (N_4533,N_4377,N_4475);
or U4534 (N_4534,N_4405,N_4459);
xnor U4535 (N_4535,N_4425,N_4391);
xor U4536 (N_4536,N_4470,N_4431);
xor U4537 (N_4537,N_4382,N_4432);
or U4538 (N_4538,N_4384,N_4379);
or U4539 (N_4539,N_4469,N_4434);
nand U4540 (N_4540,N_4330,N_4438);
nor U4541 (N_4541,N_4421,N_4454);
nor U4542 (N_4542,N_4442,N_4409);
nor U4543 (N_4543,N_4424,N_4461);
and U4544 (N_4544,N_4430,N_4411);
or U4545 (N_4545,N_4338,N_4452);
and U4546 (N_4546,N_4443,N_4477);
xor U4547 (N_4547,N_4332,N_4374);
and U4548 (N_4548,N_4323,N_4472);
and U4549 (N_4549,N_4378,N_4453);
and U4550 (N_4550,N_4414,N_4393);
and U4551 (N_4551,N_4476,N_4416);
nand U4552 (N_4552,N_4440,N_4340);
xor U4553 (N_4553,N_4350,N_4345);
xor U4554 (N_4554,N_4369,N_4407);
xor U4555 (N_4555,N_4392,N_4406);
and U4556 (N_4556,N_4329,N_4334);
nor U4557 (N_4557,N_4385,N_4331);
or U4558 (N_4558,N_4368,N_4463);
and U4559 (N_4559,N_4337,N_4444);
or U4560 (N_4560,N_4348,N_4374);
and U4561 (N_4561,N_4423,N_4331);
and U4562 (N_4562,N_4330,N_4456);
or U4563 (N_4563,N_4383,N_4359);
and U4564 (N_4564,N_4400,N_4418);
or U4565 (N_4565,N_4355,N_4455);
and U4566 (N_4566,N_4336,N_4447);
nand U4567 (N_4567,N_4465,N_4423);
or U4568 (N_4568,N_4381,N_4375);
nor U4569 (N_4569,N_4330,N_4339);
nor U4570 (N_4570,N_4462,N_4382);
nand U4571 (N_4571,N_4459,N_4358);
or U4572 (N_4572,N_4435,N_4400);
xnor U4573 (N_4573,N_4474,N_4361);
or U4574 (N_4574,N_4393,N_4394);
and U4575 (N_4575,N_4467,N_4339);
nor U4576 (N_4576,N_4389,N_4374);
nand U4577 (N_4577,N_4338,N_4369);
and U4578 (N_4578,N_4354,N_4369);
or U4579 (N_4579,N_4472,N_4435);
or U4580 (N_4580,N_4368,N_4454);
xor U4581 (N_4581,N_4383,N_4459);
nand U4582 (N_4582,N_4375,N_4334);
nand U4583 (N_4583,N_4367,N_4413);
or U4584 (N_4584,N_4390,N_4468);
and U4585 (N_4585,N_4354,N_4373);
xor U4586 (N_4586,N_4426,N_4401);
xor U4587 (N_4587,N_4329,N_4376);
or U4588 (N_4588,N_4392,N_4425);
and U4589 (N_4589,N_4431,N_4354);
or U4590 (N_4590,N_4441,N_4410);
xor U4591 (N_4591,N_4408,N_4338);
nor U4592 (N_4592,N_4347,N_4391);
nor U4593 (N_4593,N_4412,N_4390);
nand U4594 (N_4594,N_4321,N_4386);
and U4595 (N_4595,N_4401,N_4343);
and U4596 (N_4596,N_4466,N_4436);
nor U4597 (N_4597,N_4363,N_4413);
xnor U4598 (N_4598,N_4357,N_4368);
and U4599 (N_4599,N_4433,N_4414);
xor U4600 (N_4600,N_4330,N_4378);
xor U4601 (N_4601,N_4433,N_4325);
and U4602 (N_4602,N_4366,N_4459);
xnor U4603 (N_4603,N_4463,N_4455);
nor U4604 (N_4604,N_4450,N_4386);
nor U4605 (N_4605,N_4382,N_4447);
nand U4606 (N_4606,N_4322,N_4448);
xnor U4607 (N_4607,N_4408,N_4366);
and U4608 (N_4608,N_4351,N_4417);
nor U4609 (N_4609,N_4448,N_4474);
xnor U4610 (N_4610,N_4368,N_4388);
xnor U4611 (N_4611,N_4357,N_4433);
or U4612 (N_4612,N_4407,N_4327);
nand U4613 (N_4613,N_4447,N_4385);
xnor U4614 (N_4614,N_4381,N_4471);
nand U4615 (N_4615,N_4412,N_4326);
nand U4616 (N_4616,N_4400,N_4448);
and U4617 (N_4617,N_4327,N_4432);
nand U4618 (N_4618,N_4380,N_4368);
and U4619 (N_4619,N_4449,N_4341);
xnor U4620 (N_4620,N_4327,N_4328);
nand U4621 (N_4621,N_4359,N_4391);
nor U4622 (N_4622,N_4326,N_4320);
xnor U4623 (N_4623,N_4354,N_4447);
nand U4624 (N_4624,N_4369,N_4371);
xnor U4625 (N_4625,N_4422,N_4479);
nor U4626 (N_4626,N_4404,N_4385);
nor U4627 (N_4627,N_4435,N_4360);
nor U4628 (N_4628,N_4452,N_4451);
nand U4629 (N_4629,N_4323,N_4334);
and U4630 (N_4630,N_4419,N_4407);
and U4631 (N_4631,N_4351,N_4356);
nor U4632 (N_4632,N_4361,N_4442);
and U4633 (N_4633,N_4430,N_4439);
nand U4634 (N_4634,N_4419,N_4428);
and U4635 (N_4635,N_4425,N_4410);
nand U4636 (N_4636,N_4345,N_4373);
or U4637 (N_4637,N_4342,N_4364);
nor U4638 (N_4638,N_4436,N_4365);
nor U4639 (N_4639,N_4421,N_4320);
and U4640 (N_4640,N_4607,N_4618);
and U4641 (N_4641,N_4638,N_4566);
xor U4642 (N_4642,N_4511,N_4589);
and U4643 (N_4643,N_4595,N_4611);
nand U4644 (N_4644,N_4541,N_4540);
or U4645 (N_4645,N_4533,N_4612);
and U4646 (N_4646,N_4556,N_4604);
and U4647 (N_4647,N_4490,N_4531);
nor U4648 (N_4648,N_4507,N_4623);
and U4649 (N_4649,N_4510,N_4588);
nor U4650 (N_4650,N_4543,N_4495);
nand U4651 (N_4651,N_4622,N_4572);
nand U4652 (N_4652,N_4485,N_4577);
or U4653 (N_4653,N_4512,N_4516);
nor U4654 (N_4654,N_4505,N_4621);
and U4655 (N_4655,N_4606,N_4601);
nand U4656 (N_4656,N_4628,N_4527);
and U4657 (N_4657,N_4591,N_4608);
and U4658 (N_4658,N_4635,N_4487);
and U4659 (N_4659,N_4552,N_4500);
nor U4660 (N_4660,N_4548,N_4626);
nor U4661 (N_4661,N_4596,N_4528);
nor U4662 (N_4662,N_4633,N_4494);
nand U4663 (N_4663,N_4598,N_4561);
or U4664 (N_4664,N_4491,N_4605);
or U4665 (N_4665,N_4587,N_4590);
or U4666 (N_4666,N_4619,N_4594);
xnor U4667 (N_4667,N_4536,N_4522);
xor U4668 (N_4668,N_4597,N_4538);
or U4669 (N_4669,N_4625,N_4488);
or U4670 (N_4670,N_4486,N_4515);
and U4671 (N_4671,N_4547,N_4639);
and U4672 (N_4672,N_4545,N_4503);
nand U4673 (N_4673,N_4569,N_4574);
xnor U4674 (N_4674,N_4519,N_4497);
nor U4675 (N_4675,N_4537,N_4482);
nand U4676 (N_4676,N_4629,N_4489);
xor U4677 (N_4677,N_4636,N_4514);
and U4678 (N_4678,N_4544,N_4513);
or U4679 (N_4679,N_4565,N_4508);
nand U4680 (N_4680,N_4571,N_4483);
or U4681 (N_4681,N_4480,N_4509);
or U4682 (N_4682,N_4524,N_4521);
nor U4683 (N_4683,N_4570,N_4616);
or U4684 (N_4684,N_4539,N_4484);
and U4685 (N_4685,N_4564,N_4554);
or U4686 (N_4686,N_4578,N_4492);
xor U4687 (N_4687,N_4602,N_4610);
xor U4688 (N_4688,N_4501,N_4632);
and U4689 (N_4689,N_4581,N_4575);
nand U4690 (N_4690,N_4599,N_4624);
nor U4691 (N_4691,N_4614,N_4620);
nor U4692 (N_4692,N_4603,N_4549);
nor U4693 (N_4693,N_4520,N_4613);
nand U4694 (N_4694,N_4615,N_4567);
or U4695 (N_4695,N_4560,N_4584);
and U4696 (N_4696,N_4526,N_4532);
nor U4697 (N_4697,N_4593,N_4546);
nand U4698 (N_4698,N_4583,N_4517);
xor U4699 (N_4699,N_4559,N_4634);
nor U4700 (N_4700,N_4529,N_4637);
and U4701 (N_4701,N_4542,N_4631);
xnor U4702 (N_4702,N_4562,N_4585);
and U4703 (N_4703,N_4558,N_4600);
xor U4704 (N_4704,N_4557,N_4563);
nand U4705 (N_4705,N_4530,N_4502);
or U4706 (N_4706,N_4496,N_4481);
nand U4707 (N_4707,N_4617,N_4553);
or U4708 (N_4708,N_4518,N_4499);
nand U4709 (N_4709,N_4525,N_4493);
and U4710 (N_4710,N_4498,N_4580);
or U4711 (N_4711,N_4579,N_4551);
nand U4712 (N_4712,N_4586,N_4582);
nor U4713 (N_4713,N_4535,N_4550);
nand U4714 (N_4714,N_4627,N_4504);
nor U4715 (N_4715,N_4506,N_4523);
xor U4716 (N_4716,N_4576,N_4568);
nor U4717 (N_4717,N_4592,N_4573);
or U4718 (N_4718,N_4534,N_4630);
xnor U4719 (N_4719,N_4609,N_4555);
or U4720 (N_4720,N_4536,N_4501);
or U4721 (N_4721,N_4633,N_4637);
and U4722 (N_4722,N_4502,N_4557);
xor U4723 (N_4723,N_4507,N_4627);
and U4724 (N_4724,N_4570,N_4537);
nor U4725 (N_4725,N_4537,N_4581);
nor U4726 (N_4726,N_4587,N_4542);
nand U4727 (N_4727,N_4569,N_4616);
or U4728 (N_4728,N_4553,N_4638);
nand U4729 (N_4729,N_4550,N_4506);
and U4730 (N_4730,N_4543,N_4542);
xor U4731 (N_4731,N_4506,N_4554);
nor U4732 (N_4732,N_4552,N_4514);
nor U4733 (N_4733,N_4578,N_4623);
nor U4734 (N_4734,N_4576,N_4599);
nand U4735 (N_4735,N_4539,N_4496);
and U4736 (N_4736,N_4575,N_4627);
or U4737 (N_4737,N_4531,N_4487);
or U4738 (N_4738,N_4503,N_4538);
xnor U4739 (N_4739,N_4503,N_4508);
xor U4740 (N_4740,N_4490,N_4625);
xor U4741 (N_4741,N_4622,N_4515);
xor U4742 (N_4742,N_4497,N_4569);
nor U4743 (N_4743,N_4516,N_4570);
and U4744 (N_4744,N_4537,N_4604);
or U4745 (N_4745,N_4495,N_4602);
nor U4746 (N_4746,N_4628,N_4548);
xor U4747 (N_4747,N_4545,N_4550);
or U4748 (N_4748,N_4599,N_4614);
nand U4749 (N_4749,N_4587,N_4545);
or U4750 (N_4750,N_4629,N_4486);
xnor U4751 (N_4751,N_4580,N_4588);
nand U4752 (N_4752,N_4567,N_4549);
nor U4753 (N_4753,N_4501,N_4527);
nor U4754 (N_4754,N_4529,N_4521);
and U4755 (N_4755,N_4543,N_4582);
and U4756 (N_4756,N_4633,N_4486);
nor U4757 (N_4757,N_4600,N_4634);
and U4758 (N_4758,N_4609,N_4612);
nand U4759 (N_4759,N_4572,N_4528);
and U4760 (N_4760,N_4504,N_4551);
nor U4761 (N_4761,N_4619,N_4604);
or U4762 (N_4762,N_4612,N_4483);
nor U4763 (N_4763,N_4490,N_4511);
or U4764 (N_4764,N_4554,N_4492);
or U4765 (N_4765,N_4485,N_4546);
xnor U4766 (N_4766,N_4538,N_4587);
nor U4767 (N_4767,N_4618,N_4623);
xor U4768 (N_4768,N_4615,N_4605);
or U4769 (N_4769,N_4559,N_4535);
or U4770 (N_4770,N_4504,N_4585);
nor U4771 (N_4771,N_4620,N_4597);
nor U4772 (N_4772,N_4525,N_4599);
nor U4773 (N_4773,N_4606,N_4513);
or U4774 (N_4774,N_4612,N_4506);
and U4775 (N_4775,N_4605,N_4547);
and U4776 (N_4776,N_4521,N_4542);
and U4777 (N_4777,N_4522,N_4575);
nor U4778 (N_4778,N_4530,N_4600);
xor U4779 (N_4779,N_4541,N_4487);
nor U4780 (N_4780,N_4591,N_4604);
nor U4781 (N_4781,N_4590,N_4568);
or U4782 (N_4782,N_4608,N_4619);
nand U4783 (N_4783,N_4544,N_4487);
nand U4784 (N_4784,N_4524,N_4622);
and U4785 (N_4785,N_4600,N_4506);
nor U4786 (N_4786,N_4639,N_4582);
xor U4787 (N_4787,N_4584,N_4581);
nor U4788 (N_4788,N_4511,N_4582);
xnor U4789 (N_4789,N_4546,N_4604);
nand U4790 (N_4790,N_4512,N_4639);
nor U4791 (N_4791,N_4529,N_4527);
and U4792 (N_4792,N_4625,N_4624);
xnor U4793 (N_4793,N_4614,N_4587);
nand U4794 (N_4794,N_4540,N_4501);
or U4795 (N_4795,N_4605,N_4569);
xor U4796 (N_4796,N_4601,N_4639);
nor U4797 (N_4797,N_4526,N_4553);
nor U4798 (N_4798,N_4629,N_4628);
nor U4799 (N_4799,N_4592,N_4525);
xnor U4800 (N_4800,N_4665,N_4753);
xor U4801 (N_4801,N_4744,N_4731);
nor U4802 (N_4802,N_4766,N_4687);
xnor U4803 (N_4803,N_4751,N_4728);
nor U4804 (N_4804,N_4694,N_4795);
or U4805 (N_4805,N_4649,N_4693);
or U4806 (N_4806,N_4733,N_4793);
or U4807 (N_4807,N_4797,N_4770);
nor U4808 (N_4808,N_4792,N_4708);
nand U4809 (N_4809,N_4703,N_4763);
nand U4810 (N_4810,N_4768,N_4757);
xor U4811 (N_4811,N_4787,N_4683);
xnor U4812 (N_4812,N_4655,N_4765);
or U4813 (N_4813,N_4775,N_4739);
nand U4814 (N_4814,N_4781,N_4764);
nand U4815 (N_4815,N_4715,N_4661);
nor U4816 (N_4816,N_4656,N_4719);
nor U4817 (N_4817,N_4674,N_4729);
or U4818 (N_4818,N_4760,N_4667);
nand U4819 (N_4819,N_4672,N_4713);
nor U4820 (N_4820,N_4796,N_4706);
nand U4821 (N_4821,N_4700,N_4690);
and U4822 (N_4822,N_4666,N_4784);
xnor U4823 (N_4823,N_4788,N_4684);
or U4824 (N_4824,N_4720,N_4722);
nor U4825 (N_4825,N_4685,N_4642);
xnor U4826 (N_4826,N_4704,N_4747);
xor U4827 (N_4827,N_4725,N_4756);
nand U4828 (N_4828,N_4698,N_4758);
nand U4829 (N_4829,N_4738,N_4783);
nand U4830 (N_4830,N_4707,N_4794);
xor U4831 (N_4831,N_4699,N_4679);
xnor U4832 (N_4832,N_4741,N_4651);
or U4833 (N_4833,N_4681,N_4780);
nand U4834 (N_4834,N_4671,N_4740);
and U4835 (N_4835,N_4790,N_4652);
and U4836 (N_4836,N_4688,N_4723);
nor U4837 (N_4837,N_4748,N_4734);
and U4838 (N_4838,N_4745,N_4798);
xor U4839 (N_4839,N_4771,N_4697);
and U4840 (N_4840,N_4742,N_4647);
xor U4841 (N_4841,N_4767,N_4657);
nor U4842 (N_4842,N_4754,N_4658);
or U4843 (N_4843,N_4779,N_4746);
nor U4844 (N_4844,N_4778,N_4730);
nand U4845 (N_4845,N_4718,N_4721);
nor U4846 (N_4846,N_4673,N_4759);
or U4847 (N_4847,N_4732,N_4772);
nor U4848 (N_4848,N_4646,N_4752);
nand U4849 (N_4849,N_4662,N_4743);
and U4850 (N_4850,N_4689,N_4659);
nor U4851 (N_4851,N_4643,N_4664);
nor U4852 (N_4852,N_4701,N_4785);
nand U4853 (N_4853,N_4726,N_4789);
or U4854 (N_4854,N_4692,N_4709);
or U4855 (N_4855,N_4676,N_4711);
xor U4856 (N_4856,N_4737,N_4680);
or U4857 (N_4857,N_4670,N_4645);
or U4858 (N_4858,N_4735,N_4717);
nand U4859 (N_4859,N_4755,N_4677);
or U4860 (N_4860,N_4750,N_4782);
nand U4861 (N_4861,N_4663,N_4686);
or U4862 (N_4862,N_4786,N_4716);
or U4863 (N_4863,N_4654,N_4791);
nand U4864 (N_4864,N_4710,N_4640);
nor U4865 (N_4865,N_4762,N_4736);
nor U4866 (N_4866,N_4705,N_4695);
nor U4867 (N_4867,N_4682,N_4678);
nor U4868 (N_4868,N_4648,N_4653);
or U4869 (N_4869,N_4727,N_4777);
or U4870 (N_4870,N_4749,N_4696);
nand U4871 (N_4871,N_4660,N_4668);
xor U4872 (N_4872,N_4761,N_4650);
nand U4873 (N_4873,N_4776,N_4669);
or U4874 (N_4874,N_4774,N_4691);
nand U4875 (N_4875,N_4675,N_4714);
nor U4876 (N_4876,N_4712,N_4641);
or U4877 (N_4877,N_4769,N_4644);
nand U4878 (N_4878,N_4799,N_4773);
nor U4879 (N_4879,N_4702,N_4724);
nand U4880 (N_4880,N_4765,N_4683);
or U4881 (N_4881,N_4765,N_4671);
nor U4882 (N_4882,N_4663,N_4671);
or U4883 (N_4883,N_4795,N_4719);
and U4884 (N_4884,N_4690,N_4679);
or U4885 (N_4885,N_4669,N_4641);
and U4886 (N_4886,N_4759,N_4691);
and U4887 (N_4887,N_4785,N_4721);
xnor U4888 (N_4888,N_4694,N_4688);
nor U4889 (N_4889,N_4734,N_4763);
nand U4890 (N_4890,N_4710,N_4740);
nand U4891 (N_4891,N_4781,N_4762);
xnor U4892 (N_4892,N_4685,N_4679);
nand U4893 (N_4893,N_4707,N_4667);
xor U4894 (N_4894,N_4645,N_4640);
nor U4895 (N_4895,N_4771,N_4646);
nand U4896 (N_4896,N_4700,N_4762);
or U4897 (N_4897,N_4756,N_4726);
or U4898 (N_4898,N_4758,N_4671);
nor U4899 (N_4899,N_4648,N_4796);
nand U4900 (N_4900,N_4797,N_4686);
xnor U4901 (N_4901,N_4646,N_4672);
xnor U4902 (N_4902,N_4693,N_4756);
nor U4903 (N_4903,N_4752,N_4660);
nor U4904 (N_4904,N_4645,N_4714);
nand U4905 (N_4905,N_4771,N_4756);
xor U4906 (N_4906,N_4715,N_4705);
or U4907 (N_4907,N_4658,N_4719);
nand U4908 (N_4908,N_4646,N_4695);
nand U4909 (N_4909,N_4683,N_4650);
or U4910 (N_4910,N_4679,N_4695);
or U4911 (N_4911,N_4666,N_4798);
and U4912 (N_4912,N_4729,N_4723);
xor U4913 (N_4913,N_4725,N_4734);
or U4914 (N_4914,N_4750,N_4790);
and U4915 (N_4915,N_4660,N_4735);
nand U4916 (N_4916,N_4764,N_4695);
and U4917 (N_4917,N_4739,N_4717);
or U4918 (N_4918,N_4666,N_4645);
and U4919 (N_4919,N_4648,N_4681);
and U4920 (N_4920,N_4651,N_4771);
xnor U4921 (N_4921,N_4786,N_4681);
or U4922 (N_4922,N_4798,N_4789);
nand U4923 (N_4923,N_4771,N_4648);
nor U4924 (N_4924,N_4644,N_4701);
xnor U4925 (N_4925,N_4738,N_4759);
and U4926 (N_4926,N_4693,N_4725);
nand U4927 (N_4927,N_4740,N_4756);
or U4928 (N_4928,N_4750,N_4769);
or U4929 (N_4929,N_4687,N_4769);
xor U4930 (N_4930,N_4680,N_4725);
or U4931 (N_4931,N_4717,N_4729);
xor U4932 (N_4932,N_4795,N_4775);
xor U4933 (N_4933,N_4788,N_4691);
xor U4934 (N_4934,N_4669,N_4791);
xor U4935 (N_4935,N_4702,N_4679);
xnor U4936 (N_4936,N_4671,N_4774);
nor U4937 (N_4937,N_4692,N_4706);
xnor U4938 (N_4938,N_4680,N_4645);
and U4939 (N_4939,N_4656,N_4791);
xnor U4940 (N_4940,N_4677,N_4757);
and U4941 (N_4941,N_4728,N_4644);
nand U4942 (N_4942,N_4696,N_4797);
and U4943 (N_4943,N_4651,N_4714);
and U4944 (N_4944,N_4677,N_4727);
and U4945 (N_4945,N_4765,N_4739);
and U4946 (N_4946,N_4759,N_4780);
and U4947 (N_4947,N_4759,N_4765);
nor U4948 (N_4948,N_4692,N_4792);
and U4949 (N_4949,N_4784,N_4669);
xor U4950 (N_4950,N_4642,N_4644);
xnor U4951 (N_4951,N_4648,N_4693);
and U4952 (N_4952,N_4671,N_4787);
and U4953 (N_4953,N_4710,N_4782);
or U4954 (N_4954,N_4789,N_4764);
and U4955 (N_4955,N_4788,N_4736);
xor U4956 (N_4956,N_4766,N_4701);
nor U4957 (N_4957,N_4799,N_4739);
or U4958 (N_4958,N_4778,N_4690);
nand U4959 (N_4959,N_4784,N_4725);
nor U4960 (N_4960,N_4882,N_4950);
nand U4961 (N_4961,N_4910,N_4850);
nand U4962 (N_4962,N_4904,N_4833);
or U4963 (N_4963,N_4837,N_4844);
and U4964 (N_4964,N_4846,N_4845);
nand U4965 (N_4965,N_4928,N_4841);
nor U4966 (N_4966,N_4941,N_4920);
and U4967 (N_4967,N_4956,N_4861);
and U4968 (N_4968,N_4802,N_4842);
nor U4969 (N_4969,N_4951,N_4892);
xor U4970 (N_4970,N_4817,N_4902);
or U4971 (N_4971,N_4893,N_4889);
nand U4972 (N_4972,N_4839,N_4923);
nor U4973 (N_4973,N_4914,N_4911);
or U4974 (N_4974,N_4942,N_4822);
and U4975 (N_4975,N_4947,N_4866);
nand U4976 (N_4976,N_4849,N_4917);
nor U4977 (N_4977,N_4948,N_4880);
nor U4978 (N_4978,N_4940,N_4819);
nor U4979 (N_4979,N_4898,N_4934);
nand U4980 (N_4980,N_4901,N_4958);
nor U4981 (N_4981,N_4815,N_4831);
nor U4982 (N_4982,N_4903,N_4812);
xnor U4983 (N_4983,N_4926,N_4938);
or U4984 (N_4984,N_4908,N_4811);
and U4985 (N_4985,N_4804,N_4927);
xnor U4986 (N_4986,N_4825,N_4879);
xor U4987 (N_4987,N_4943,N_4883);
and U4988 (N_4988,N_4945,N_4877);
xor U4989 (N_4989,N_4888,N_4873);
nand U4990 (N_4990,N_4946,N_4868);
nor U4991 (N_4991,N_4924,N_4847);
xnor U4992 (N_4992,N_4890,N_4854);
or U4993 (N_4993,N_4929,N_4939);
nor U4994 (N_4994,N_4807,N_4878);
or U4995 (N_4995,N_4870,N_4955);
nor U4996 (N_4996,N_4801,N_4918);
nand U4997 (N_4997,N_4823,N_4810);
nand U4998 (N_4998,N_4897,N_4949);
or U4999 (N_4999,N_4875,N_4858);
or U5000 (N_5000,N_4835,N_4957);
nand U5001 (N_5001,N_4916,N_4824);
nor U5002 (N_5002,N_4816,N_4891);
nor U5003 (N_5003,N_4836,N_4921);
nand U5004 (N_5004,N_4912,N_4872);
nand U5005 (N_5005,N_4874,N_4922);
xor U5006 (N_5006,N_4809,N_4820);
nor U5007 (N_5007,N_4863,N_4906);
nand U5008 (N_5008,N_4907,N_4855);
xnor U5009 (N_5009,N_4853,N_4859);
xnor U5010 (N_5010,N_4867,N_4856);
nand U5011 (N_5011,N_4851,N_4885);
nor U5012 (N_5012,N_4919,N_4813);
or U5013 (N_5013,N_4864,N_4959);
and U5014 (N_5014,N_4803,N_4857);
or U5015 (N_5015,N_4935,N_4805);
xnor U5016 (N_5016,N_4936,N_4937);
nor U5017 (N_5017,N_4827,N_4832);
nand U5018 (N_5018,N_4840,N_4930);
xnor U5019 (N_5019,N_4800,N_4899);
nor U5020 (N_5020,N_4884,N_4894);
nand U5021 (N_5021,N_4860,N_4952);
nand U5022 (N_5022,N_4896,N_4826);
xnor U5023 (N_5023,N_4834,N_4944);
nand U5024 (N_5024,N_4829,N_4954);
and U5025 (N_5025,N_4905,N_4818);
or U5026 (N_5026,N_4953,N_4900);
and U5027 (N_5027,N_4821,N_4876);
nand U5028 (N_5028,N_4886,N_4869);
nand U5029 (N_5029,N_4881,N_4925);
or U5030 (N_5030,N_4806,N_4933);
or U5031 (N_5031,N_4913,N_4848);
and U5032 (N_5032,N_4865,N_4895);
and U5033 (N_5033,N_4814,N_4887);
or U5034 (N_5034,N_4909,N_4808);
or U5035 (N_5035,N_4843,N_4871);
and U5036 (N_5036,N_4932,N_4852);
nand U5037 (N_5037,N_4915,N_4830);
or U5038 (N_5038,N_4838,N_4862);
nor U5039 (N_5039,N_4828,N_4931);
xnor U5040 (N_5040,N_4938,N_4875);
nor U5041 (N_5041,N_4821,N_4877);
xor U5042 (N_5042,N_4818,N_4920);
nand U5043 (N_5043,N_4908,N_4848);
or U5044 (N_5044,N_4943,N_4813);
and U5045 (N_5045,N_4903,N_4934);
nor U5046 (N_5046,N_4827,N_4943);
or U5047 (N_5047,N_4854,N_4917);
nand U5048 (N_5048,N_4886,N_4800);
or U5049 (N_5049,N_4870,N_4949);
xor U5050 (N_5050,N_4847,N_4829);
or U5051 (N_5051,N_4882,N_4934);
and U5052 (N_5052,N_4873,N_4869);
xor U5053 (N_5053,N_4929,N_4876);
and U5054 (N_5054,N_4847,N_4805);
or U5055 (N_5055,N_4843,N_4928);
and U5056 (N_5056,N_4819,N_4875);
and U5057 (N_5057,N_4889,N_4933);
or U5058 (N_5058,N_4808,N_4915);
or U5059 (N_5059,N_4870,N_4848);
nor U5060 (N_5060,N_4844,N_4830);
nor U5061 (N_5061,N_4921,N_4902);
and U5062 (N_5062,N_4867,N_4926);
and U5063 (N_5063,N_4922,N_4863);
or U5064 (N_5064,N_4921,N_4933);
xnor U5065 (N_5065,N_4917,N_4851);
nor U5066 (N_5066,N_4849,N_4874);
xnor U5067 (N_5067,N_4888,N_4957);
xor U5068 (N_5068,N_4954,N_4900);
or U5069 (N_5069,N_4879,N_4817);
nand U5070 (N_5070,N_4898,N_4852);
nor U5071 (N_5071,N_4855,N_4936);
and U5072 (N_5072,N_4890,N_4878);
nand U5073 (N_5073,N_4803,N_4844);
nor U5074 (N_5074,N_4891,N_4896);
nor U5075 (N_5075,N_4830,N_4839);
and U5076 (N_5076,N_4887,N_4907);
and U5077 (N_5077,N_4953,N_4929);
nand U5078 (N_5078,N_4929,N_4928);
and U5079 (N_5079,N_4872,N_4919);
nand U5080 (N_5080,N_4947,N_4877);
xor U5081 (N_5081,N_4874,N_4843);
and U5082 (N_5082,N_4885,N_4854);
or U5083 (N_5083,N_4857,N_4927);
nand U5084 (N_5084,N_4886,N_4890);
or U5085 (N_5085,N_4801,N_4853);
xnor U5086 (N_5086,N_4931,N_4909);
and U5087 (N_5087,N_4870,N_4868);
nor U5088 (N_5088,N_4879,N_4883);
nor U5089 (N_5089,N_4824,N_4897);
nand U5090 (N_5090,N_4854,N_4901);
nand U5091 (N_5091,N_4855,N_4898);
nand U5092 (N_5092,N_4801,N_4941);
nor U5093 (N_5093,N_4883,N_4826);
xnor U5094 (N_5094,N_4902,N_4863);
and U5095 (N_5095,N_4817,N_4860);
or U5096 (N_5096,N_4952,N_4927);
nor U5097 (N_5097,N_4882,N_4854);
xor U5098 (N_5098,N_4935,N_4823);
or U5099 (N_5099,N_4934,N_4909);
or U5100 (N_5100,N_4877,N_4940);
or U5101 (N_5101,N_4892,N_4880);
nand U5102 (N_5102,N_4879,N_4899);
and U5103 (N_5103,N_4884,N_4927);
or U5104 (N_5104,N_4847,N_4940);
and U5105 (N_5105,N_4853,N_4880);
and U5106 (N_5106,N_4955,N_4889);
xor U5107 (N_5107,N_4893,N_4814);
nor U5108 (N_5108,N_4820,N_4912);
or U5109 (N_5109,N_4896,N_4843);
nand U5110 (N_5110,N_4831,N_4942);
or U5111 (N_5111,N_4820,N_4902);
nand U5112 (N_5112,N_4870,N_4890);
xnor U5113 (N_5113,N_4813,N_4914);
and U5114 (N_5114,N_4801,N_4908);
nand U5115 (N_5115,N_4858,N_4833);
nand U5116 (N_5116,N_4950,N_4884);
nand U5117 (N_5117,N_4899,N_4824);
or U5118 (N_5118,N_4931,N_4816);
or U5119 (N_5119,N_4863,N_4865);
nor U5120 (N_5120,N_5099,N_5075);
and U5121 (N_5121,N_5092,N_4976);
nand U5122 (N_5122,N_4980,N_5047);
nand U5123 (N_5123,N_5029,N_5090);
nand U5124 (N_5124,N_4974,N_4990);
or U5125 (N_5125,N_5072,N_5021);
nand U5126 (N_5126,N_5111,N_5070);
and U5127 (N_5127,N_5015,N_5002);
nor U5128 (N_5128,N_5008,N_4965);
nand U5129 (N_5129,N_5071,N_5112);
nor U5130 (N_5130,N_4999,N_4993);
or U5131 (N_5131,N_5105,N_5058);
nor U5132 (N_5132,N_5096,N_5083);
nor U5133 (N_5133,N_5025,N_4972);
or U5134 (N_5134,N_5016,N_4967);
nand U5135 (N_5135,N_5011,N_5010);
nor U5136 (N_5136,N_5118,N_5078);
or U5137 (N_5137,N_4987,N_5062);
xor U5138 (N_5138,N_5098,N_4984);
nor U5139 (N_5139,N_5088,N_5086);
nand U5140 (N_5140,N_5028,N_5110);
nor U5141 (N_5141,N_5039,N_5109);
nor U5142 (N_5142,N_5017,N_5026);
nor U5143 (N_5143,N_4979,N_5082);
xnor U5144 (N_5144,N_4964,N_5030);
or U5145 (N_5145,N_5041,N_4982);
or U5146 (N_5146,N_5007,N_4962);
nor U5147 (N_5147,N_5065,N_5051);
xnor U5148 (N_5148,N_4971,N_5012);
or U5149 (N_5149,N_5085,N_5059);
and U5150 (N_5150,N_4969,N_5003);
or U5151 (N_5151,N_5093,N_5023);
or U5152 (N_5152,N_4975,N_5104);
or U5153 (N_5153,N_5080,N_5004);
and U5154 (N_5154,N_5081,N_5038);
xor U5155 (N_5155,N_5089,N_4995);
nand U5156 (N_5156,N_5046,N_5014);
or U5157 (N_5157,N_5066,N_5061);
and U5158 (N_5158,N_5114,N_5107);
nand U5159 (N_5159,N_5005,N_4997);
and U5160 (N_5160,N_4985,N_4977);
nand U5161 (N_5161,N_5044,N_5077);
nand U5162 (N_5162,N_5031,N_5064);
nand U5163 (N_5163,N_5097,N_5019);
xnor U5164 (N_5164,N_5102,N_5040);
nand U5165 (N_5165,N_5033,N_5000);
nor U5166 (N_5166,N_5022,N_5079);
nor U5167 (N_5167,N_5063,N_4998);
nand U5168 (N_5168,N_5043,N_5009);
xor U5169 (N_5169,N_5018,N_5045);
xor U5170 (N_5170,N_5091,N_5074);
or U5171 (N_5171,N_5032,N_4992);
nand U5172 (N_5172,N_4994,N_5060);
and U5173 (N_5173,N_5069,N_5034);
xor U5174 (N_5174,N_5108,N_4983);
or U5175 (N_5175,N_5073,N_4986);
and U5176 (N_5176,N_5036,N_5052);
xor U5177 (N_5177,N_5101,N_5020);
or U5178 (N_5178,N_5042,N_5053);
and U5179 (N_5179,N_5115,N_5084);
nand U5180 (N_5180,N_5067,N_5056);
xnor U5181 (N_5181,N_4989,N_5048);
nand U5182 (N_5182,N_5117,N_5037);
xor U5183 (N_5183,N_5035,N_5094);
or U5184 (N_5184,N_5054,N_4996);
nor U5185 (N_5185,N_4991,N_5116);
nand U5186 (N_5186,N_5113,N_4970);
or U5187 (N_5187,N_5001,N_4981);
nand U5188 (N_5188,N_4978,N_5055);
and U5189 (N_5189,N_4973,N_5095);
and U5190 (N_5190,N_5087,N_5006);
xnor U5191 (N_5191,N_5068,N_4960);
nor U5192 (N_5192,N_5013,N_5106);
and U5193 (N_5193,N_4988,N_5103);
and U5194 (N_5194,N_5100,N_5076);
or U5195 (N_5195,N_4961,N_5024);
nand U5196 (N_5196,N_5027,N_4966);
nor U5197 (N_5197,N_5119,N_5049);
nor U5198 (N_5198,N_4968,N_5050);
nor U5199 (N_5199,N_4963,N_5057);
or U5200 (N_5200,N_4980,N_4987);
nand U5201 (N_5201,N_4978,N_5106);
or U5202 (N_5202,N_5030,N_5051);
nand U5203 (N_5203,N_5034,N_5110);
and U5204 (N_5204,N_5020,N_5003);
or U5205 (N_5205,N_5104,N_5012);
xor U5206 (N_5206,N_4988,N_4974);
xor U5207 (N_5207,N_4978,N_5082);
nand U5208 (N_5208,N_5106,N_5099);
and U5209 (N_5209,N_5016,N_4985);
xor U5210 (N_5210,N_5045,N_4967);
xor U5211 (N_5211,N_4989,N_5119);
nor U5212 (N_5212,N_4972,N_5103);
nand U5213 (N_5213,N_5088,N_5051);
nor U5214 (N_5214,N_5036,N_5002);
or U5215 (N_5215,N_5003,N_5057);
and U5216 (N_5216,N_5069,N_5090);
xor U5217 (N_5217,N_5090,N_4991);
nor U5218 (N_5218,N_5020,N_5038);
or U5219 (N_5219,N_5077,N_4990);
nand U5220 (N_5220,N_5107,N_4971);
xnor U5221 (N_5221,N_5043,N_5073);
nand U5222 (N_5222,N_5037,N_5003);
and U5223 (N_5223,N_4976,N_4999);
nor U5224 (N_5224,N_4997,N_5073);
xnor U5225 (N_5225,N_4990,N_5067);
or U5226 (N_5226,N_4996,N_4985);
nand U5227 (N_5227,N_5119,N_4974);
xor U5228 (N_5228,N_4984,N_5109);
nor U5229 (N_5229,N_5070,N_4972);
xnor U5230 (N_5230,N_4976,N_5034);
nor U5231 (N_5231,N_4982,N_5026);
or U5232 (N_5232,N_5010,N_5078);
and U5233 (N_5233,N_5085,N_4983);
nor U5234 (N_5234,N_5008,N_4997);
nand U5235 (N_5235,N_5100,N_5054);
nand U5236 (N_5236,N_5104,N_5041);
or U5237 (N_5237,N_5115,N_4976);
and U5238 (N_5238,N_5036,N_5093);
nor U5239 (N_5239,N_5051,N_5012);
nand U5240 (N_5240,N_5059,N_5101);
and U5241 (N_5241,N_5027,N_5105);
nor U5242 (N_5242,N_5113,N_5010);
nand U5243 (N_5243,N_5077,N_5035);
and U5244 (N_5244,N_5057,N_5079);
and U5245 (N_5245,N_5084,N_4972);
nand U5246 (N_5246,N_5020,N_5114);
or U5247 (N_5247,N_4972,N_4989);
nor U5248 (N_5248,N_4985,N_5034);
or U5249 (N_5249,N_5033,N_5106);
nor U5250 (N_5250,N_5073,N_5089);
xor U5251 (N_5251,N_5010,N_5116);
nor U5252 (N_5252,N_5072,N_5056);
nor U5253 (N_5253,N_4969,N_4988);
xor U5254 (N_5254,N_5071,N_5009);
xnor U5255 (N_5255,N_4986,N_5086);
or U5256 (N_5256,N_5022,N_4994);
nor U5257 (N_5257,N_4985,N_5114);
nor U5258 (N_5258,N_5006,N_5062);
nand U5259 (N_5259,N_4965,N_5056);
xnor U5260 (N_5260,N_4992,N_5050);
and U5261 (N_5261,N_5118,N_5043);
nor U5262 (N_5262,N_5011,N_5078);
and U5263 (N_5263,N_4993,N_5108);
xnor U5264 (N_5264,N_5087,N_5106);
and U5265 (N_5265,N_5059,N_4983);
and U5266 (N_5266,N_5024,N_5051);
and U5267 (N_5267,N_5069,N_4992);
nand U5268 (N_5268,N_5030,N_5006);
nor U5269 (N_5269,N_5056,N_5068);
nor U5270 (N_5270,N_5060,N_4972);
and U5271 (N_5271,N_4994,N_5071);
and U5272 (N_5272,N_5065,N_5058);
and U5273 (N_5273,N_5025,N_5021);
xnor U5274 (N_5274,N_5082,N_5074);
nor U5275 (N_5275,N_4984,N_4979);
or U5276 (N_5276,N_5104,N_4989);
or U5277 (N_5277,N_5059,N_5094);
or U5278 (N_5278,N_5038,N_5116);
xnor U5279 (N_5279,N_5087,N_5058);
xnor U5280 (N_5280,N_5224,N_5251);
xor U5281 (N_5281,N_5180,N_5137);
xor U5282 (N_5282,N_5147,N_5272);
nor U5283 (N_5283,N_5149,N_5209);
xor U5284 (N_5284,N_5187,N_5260);
and U5285 (N_5285,N_5218,N_5244);
nor U5286 (N_5286,N_5219,N_5141);
or U5287 (N_5287,N_5253,N_5173);
nand U5288 (N_5288,N_5239,N_5151);
nor U5289 (N_5289,N_5133,N_5157);
nor U5290 (N_5290,N_5197,N_5127);
xor U5291 (N_5291,N_5206,N_5158);
nor U5292 (N_5292,N_5203,N_5262);
nor U5293 (N_5293,N_5257,N_5276);
xnor U5294 (N_5294,N_5123,N_5190);
nand U5295 (N_5295,N_5215,N_5225);
or U5296 (N_5296,N_5125,N_5271);
nand U5297 (N_5297,N_5177,N_5200);
nand U5298 (N_5298,N_5242,N_5196);
or U5299 (N_5299,N_5132,N_5234);
or U5300 (N_5300,N_5217,N_5179);
or U5301 (N_5301,N_5148,N_5230);
and U5302 (N_5302,N_5183,N_5162);
nand U5303 (N_5303,N_5226,N_5266);
xnor U5304 (N_5304,N_5256,N_5172);
nor U5305 (N_5305,N_5274,N_5204);
or U5306 (N_5306,N_5258,N_5176);
nand U5307 (N_5307,N_5229,N_5249);
and U5308 (N_5308,N_5191,N_5238);
and U5309 (N_5309,N_5202,N_5134);
nor U5310 (N_5310,N_5232,N_5216);
and U5311 (N_5311,N_5228,N_5174);
and U5312 (N_5312,N_5163,N_5184);
nand U5313 (N_5313,N_5277,N_5245);
nand U5314 (N_5314,N_5171,N_5146);
xnor U5315 (N_5315,N_5152,N_5124);
nor U5316 (N_5316,N_5139,N_5188);
or U5317 (N_5317,N_5178,N_5213);
or U5318 (N_5318,N_5243,N_5159);
nor U5319 (N_5319,N_5129,N_5128);
nor U5320 (N_5320,N_5221,N_5201);
nor U5321 (N_5321,N_5273,N_5150);
nor U5322 (N_5322,N_5235,N_5165);
nand U5323 (N_5323,N_5186,N_5212);
and U5324 (N_5324,N_5198,N_5126);
xnor U5325 (N_5325,N_5208,N_5153);
nor U5326 (N_5326,N_5120,N_5143);
or U5327 (N_5327,N_5138,N_5205);
or U5328 (N_5328,N_5182,N_5136);
and U5329 (N_5329,N_5194,N_5161);
nor U5330 (N_5330,N_5189,N_5241);
and U5331 (N_5331,N_5265,N_5195);
or U5332 (N_5332,N_5193,N_5270);
and U5333 (N_5333,N_5233,N_5268);
nor U5334 (N_5334,N_5122,N_5154);
nor U5335 (N_5335,N_5248,N_5167);
xnor U5336 (N_5336,N_5142,N_5220);
xnor U5337 (N_5337,N_5131,N_5210);
and U5338 (N_5338,N_5269,N_5259);
nor U5339 (N_5339,N_5166,N_5261);
xnor U5340 (N_5340,N_5279,N_5156);
or U5341 (N_5341,N_5278,N_5247);
and U5342 (N_5342,N_5130,N_5214);
nand U5343 (N_5343,N_5255,N_5135);
nand U5344 (N_5344,N_5254,N_5192);
xnor U5345 (N_5345,N_5275,N_5231);
nor U5346 (N_5346,N_5246,N_5170);
nor U5347 (N_5347,N_5164,N_5169);
xor U5348 (N_5348,N_5237,N_5250);
xnor U5349 (N_5349,N_5175,N_5211);
nand U5350 (N_5350,N_5227,N_5140);
nand U5351 (N_5351,N_5207,N_5199);
xor U5352 (N_5352,N_5181,N_5264);
and U5353 (N_5353,N_5252,N_5240);
and U5354 (N_5354,N_5223,N_5155);
xnor U5355 (N_5355,N_5222,N_5267);
nor U5356 (N_5356,N_5263,N_5145);
or U5357 (N_5357,N_5160,N_5121);
nor U5358 (N_5358,N_5185,N_5144);
or U5359 (N_5359,N_5168,N_5236);
nand U5360 (N_5360,N_5156,N_5258);
or U5361 (N_5361,N_5179,N_5146);
or U5362 (N_5362,N_5159,N_5274);
xor U5363 (N_5363,N_5156,N_5248);
xnor U5364 (N_5364,N_5147,N_5188);
or U5365 (N_5365,N_5222,N_5135);
and U5366 (N_5366,N_5180,N_5242);
and U5367 (N_5367,N_5197,N_5200);
nor U5368 (N_5368,N_5211,N_5261);
and U5369 (N_5369,N_5205,N_5243);
or U5370 (N_5370,N_5227,N_5250);
or U5371 (N_5371,N_5181,N_5124);
nor U5372 (N_5372,N_5233,N_5192);
or U5373 (N_5373,N_5274,N_5229);
xor U5374 (N_5374,N_5245,N_5192);
or U5375 (N_5375,N_5267,N_5258);
and U5376 (N_5376,N_5144,N_5172);
nand U5377 (N_5377,N_5243,N_5120);
or U5378 (N_5378,N_5265,N_5155);
nor U5379 (N_5379,N_5227,N_5209);
nor U5380 (N_5380,N_5133,N_5189);
nand U5381 (N_5381,N_5165,N_5229);
nor U5382 (N_5382,N_5142,N_5126);
and U5383 (N_5383,N_5274,N_5136);
or U5384 (N_5384,N_5126,N_5139);
or U5385 (N_5385,N_5225,N_5258);
nor U5386 (N_5386,N_5219,N_5218);
and U5387 (N_5387,N_5235,N_5255);
and U5388 (N_5388,N_5208,N_5154);
nor U5389 (N_5389,N_5198,N_5277);
xnor U5390 (N_5390,N_5125,N_5217);
nor U5391 (N_5391,N_5205,N_5120);
and U5392 (N_5392,N_5270,N_5121);
nand U5393 (N_5393,N_5143,N_5162);
nor U5394 (N_5394,N_5207,N_5192);
and U5395 (N_5395,N_5275,N_5230);
and U5396 (N_5396,N_5271,N_5196);
and U5397 (N_5397,N_5137,N_5159);
or U5398 (N_5398,N_5152,N_5153);
nand U5399 (N_5399,N_5188,N_5278);
xnor U5400 (N_5400,N_5157,N_5164);
and U5401 (N_5401,N_5157,N_5257);
and U5402 (N_5402,N_5207,N_5166);
and U5403 (N_5403,N_5199,N_5236);
nand U5404 (N_5404,N_5152,N_5195);
or U5405 (N_5405,N_5152,N_5123);
or U5406 (N_5406,N_5252,N_5268);
nor U5407 (N_5407,N_5133,N_5201);
and U5408 (N_5408,N_5245,N_5200);
or U5409 (N_5409,N_5250,N_5213);
nor U5410 (N_5410,N_5272,N_5170);
or U5411 (N_5411,N_5266,N_5210);
nand U5412 (N_5412,N_5136,N_5120);
and U5413 (N_5413,N_5130,N_5224);
and U5414 (N_5414,N_5262,N_5188);
nand U5415 (N_5415,N_5184,N_5211);
nor U5416 (N_5416,N_5252,N_5136);
nor U5417 (N_5417,N_5248,N_5256);
xnor U5418 (N_5418,N_5251,N_5150);
or U5419 (N_5419,N_5194,N_5146);
nor U5420 (N_5420,N_5179,N_5207);
nor U5421 (N_5421,N_5162,N_5255);
xor U5422 (N_5422,N_5226,N_5140);
and U5423 (N_5423,N_5157,N_5134);
xor U5424 (N_5424,N_5220,N_5231);
or U5425 (N_5425,N_5198,N_5160);
xnor U5426 (N_5426,N_5160,N_5149);
nand U5427 (N_5427,N_5268,N_5182);
and U5428 (N_5428,N_5179,N_5251);
xnor U5429 (N_5429,N_5166,N_5181);
nand U5430 (N_5430,N_5220,N_5265);
xnor U5431 (N_5431,N_5250,N_5267);
or U5432 (N_5432,N_5160,N_5216);
nand U5433 (N_5433,N_5120,N_5132);
xor U5434 (N_5434,N_5215,N_5222);
nor U5435 (N_5435,N_5223,N_5211);
nor U5436 (N_5436,N_5194,N_5261);
and U5437 (N_5437,N_5145,N_5239);
nor U5438 (N_5438,N_5199,N_5205);
xnor U5439 (N_5439,N_5153,N_5122);
or U5440 (N_5440,N_5296,N_5388);
nand U5441 (N_5441,N_5379,N_5387);
or U5442 (N_5442,N_5302,N_5325);
nand U5443 (N_5443,N_5316,N_5386);
and U5444 (N_5444,N_5412,N_5338);
nand U5445 (N_5445,N_5405,N_5283);
or U5446 (N_5446,N_5361,N_5428);
or U5447 (N_5447,N_5352,N_5301);
nor U5448 (N_5448,N_5318,N_5403);
xnor U5449 (N_5449,N_5335,N_5400);
nor U5450 (N_5450,N_5417,N_5294);
nand U5451 (N_5451,N_5320,N_5374);
and U5452 (N_5452,N_5398,N_5292);
nor U5453 (N_5453,N_5434,N_5311);
nor U5454 (N_5454,N_5280,N_5423);
xor U5455 (N_5455,N_5366,N_5392);
or U5456 (N_5456,N_5436,N_5418);
and U5457 (N_5457,N_5310,N_5340);
nor U5458 (N_5458,N_5401,N_5342);
and U5459 (N_5459,N_5383,N_5399);
nor U5460 (N_5460,N_5429,N_5426);
xnor U5461 (N_5461,N_5375,N_5373);
and U5462 (N_5462,N_5389,N_5390);
xor U5463 (N_5463,N_5350,N_5416);
xor U5464 (N_5464,N_5349,N_5363);
or U5465 (N_5465,N_5327,N_5360);
nand U5466 (N_5466,N_5393,N_5365);
nor U5467 (N_5467,N_5435,N_5300);
nor U5468 (N_5468,N_5346,N_5289);
nor U5469 (N_5469,N_5420,N_5306);
nand U5470 (N_5470,N_5427,N_5319);
nand U5471 (N_5471,N_5395,N_5305);
or U5472 (N_5472,N_5371,N_5282);
xnor U5473 (N_5473,N_5432,N_5425);
and U5474 (N_5474,N_5359,N_5362);
or U5475 (N_5475,N_5333,N_5424);
nand U5476 (N_5476,N_5380,N_5376);
and U5477 (N_5477,N_5351,N_5329);
or U5478 (N_5478,N_5323,N_5295);
nand U5479 (N_5479,N_5406,N_5337);
and U5480 (N_5480,N_5367,N_5437);
xnor U5481 (N_5481,N_5378,N_5288);
xnor U5482 (N_5482,N_5339,N_5347);
and U5483 (N_5483,N_5382,N_5321);
and U5484 (N_5484,N_5317,N_5328);
and U5485 (N_5485,N_5345,N_5397);
or U5486 (N_5486,N_5369,N_5299);
nand U5487 (N_5487,N_5414,N_5408);
xor U5488 (N_5488,N_5324,N_5355);
nor U5489 (N_5489,N_5394,N_5402);
and U5490 (N_5490,N_5286,N_5344);
or U5491 (N_5491,N_5396,N_5356);
xnor U5492 (N_5492,N_5303,N_5413);
and U5493 (N_5493,N_5385,N_5326);
nand U5494 (N_5494,N_5309,N_5322);
or U5495 (N_5495,N_5431,N_5430);
or U5496 (N_5496,N_5281,N_5411);
nor U5497 (N_5497,N_5348,N_5358);
nand U5498 (N_5498,N_5368,N_5410);
nand U5499 (N_5499,N_5381,N_5377);
nand U5500 (N_5500,N_5415,N_5330);
nor U5501 (N_5501,N_5370,N_5343);
xor U5502 (N_5502,N_5419,N_5404);
and U5503 (N_5503,N_5433,N_5364);
or U5504 (N_5504,N_5372,N_5409);
nor U5505 (N_5505,N_5439,N_5315);
nor U5506 (N_5506,N_5297,N_5422);
nand U5507 (N_5507,N_5384,N_5332);
nand U5508 (N_5508,N_5298,N_5391);
nor U5509 (N_5509,N_5336,N_5314);
and U5510 (N_5510,N_5284,N_5438);
and U5511 (N_5511,N_5341,N_5421);
nor U5512 (N_5512,N_5407,N_5291);
or U5513 (N_5513,N_5312,N_5331);
and U5514 (N_5514,N_5308,N_5293);
xor U5515 (N_5515,N_5285,N_5313);
or U5516 (N_5516,N_5304,N_5353);
nor U5517 (N_5517,N_5334,N_5287);
and U5518 (N_5518,N_5354,N_5290);
nand U5519 (N_5519,N_5357,N_5307);
nand U5520 (N_5520,N_5409,N_5354);
xor U5521 (N_5521,N_5305,N_5371);
and U5522 (N_5522,N_5433,N_5354);
nor U5523 (N_5523,N_5427,N_5439);
xor U5524 (N_5524,N_5413,N_5283);
xor U5525 (N_5525,N_5320,N_5370);
or U5526 (N_5526,N_5395,N_5383);
and U5527 (N_5527,N_5336,N_5369);
xor U5528 (N_5528,N_5417,N_5354);
nor U5529 (N_5529,N_5365,N_5404);
xor U5530 (N_5530,N_5398,N_5421);
or U5531 (N_5531,N_5331,N_5388);
and U5532 (N_5532,N_5296,N_5364);
nand U5533 (N_5533,N_5431,N_5357);
or U5534 (N_5534,N_5375,N_5353);
xor U5535 (N_5535,N_5296,N_5322);
or U5536 (N_5536,N_5328,N_5340);
and U5537 (N_5537,N_5311,N_5403);
and U5538 (N_5538,N_5409,N_5398);
and U5539 (N_5539,N_5368,N_5322);
nand U5540 (N_5540,N_5394,N_5364);
nor U5541 (N_5541,N_5380,N_5338);
nor U5542 (N_5542,N_5280,N_5369);
or U5543 (N_5543,N_5285,N_5383);
or U5544 (N_5544,N_5357,N_5339);
nor U5545 (N_5545,N_5393,N_5285);
nand U5546 (N_5546,N_5339,N_5363);
nor U5547 (N_5547,N_5284,N_5385);
and U5548 (N_5548,N_5343,N_5335);
xor U5549 (N_5549,N_5377,N_5401);
nand U5550 (N_5550,N_5341,N_5297);
nor U5551 (N_5551,N_5433,N_5399);
nor U5552 (N_5552,N_5362,N_5378);
nand U5553 (N_5553,N_5375,N_5420);
xnor U5554 (N_5554,N_5435,N_5432);
nor U5555 (N_5555,N_5284,N_5389);
and U5556 (N_5556,N_5290,N_5334);
nand U5557 (N_5557,N_5402,N_5314);
nand U5558 (N_5558,N_5372,N_5382);
or U5559 (N_5559,N_5422,N_5294);
xnor U5560 (N_5560,N_5316,N_5373);
and U5561 (N_5561,N_5321,N_5358);
nor U5562 (N_5562,N_5340,N_5409);
and U5563 (N_5563,N_5307,N_5383);
nor U5564 (N_5564,N_5345,N_5322);
and U5565 (N_5565,N_5318,N_5405);
nor U5566 (N_5566,N_5401,N_5385);
nor U5567 (N_5567,N_5285,N_5339);
nor U5568 (N_5568,N_5336,N_5412);
or U5569 (N_5569,N_5411,N_5312);
and U5570 (N_5570,N_5302,N_5329);
and U5571 (N_5571,N_5324,N_5419);
nor U5572 (N_5572,N_5321,N_5346);
xor U5573 (N_5573,N_5285,N_5368);
and U5574 (N_5574,N_5327,N_5405);
xor U5575 (N_5575,N_5360,N_5325);
nand U5576 (N_5576,N_5368,N_5435);
xor U5577 (N_5577,N_5296,N_5298);
xnor U5578 (N_5578,N_5286,N_5399);
nor U5579 (N_5579,N_5347,N_5401);
and U5580 (N_5580,N_5397,N_5331);
or U5581 (N_5581,N_5354,N_5327);
nor U5582 (N_5582,N_5350,N_5391);
or U5583 (N_5583,N_5306,N_5409);
xnor U5584 (N_5584,N_5361,N_5394);
or U5585 (N_5585,N_5433,N_5419);
or U5586 (N_5586,N_5388,N_5280);
nor U5587 (N_5587,N_5329,N_5378);
nor U5588 (N_5588,N_5422,N_5389);
xor U5589 (N_5589,N_5375,N_5360);
or U5590 (N_5590,N_5385,N_5403);
or U5591 (N_5591,N_5297,N_5420);
or U5592 (N_5592,N_5335,N_5288);
xor U5593 (N_5593,N_5298,N_5324);
or U5594 (N_5594,N_5301,N_5287);
nand U5595 (N_5595,N_5329,N_5401);
nand U5596 (N_5596,N_5299,N_5335);
and U5597 (N_5597,N_5348,N_5311);
xor U5598 (N_5598,N_5381,N_5400);
or U5599 (N_5599,N_5428,N_5338);
xor U5600 (N_5600,N_5453,N_5510);
nor U5601 (N_5601,N_5515,N_5448);
nand U5602 (N_5602,N_5497,N_5581);
nand U5603 (N_5603,N_5508,N_5494);
and U5604 (N_5604,N_5487,N_5504);
nand U5605 (N_5605,N_5468,N_5568);
or U5606 (N_5606,N_5520,N_5511);
and U5607 (N_5607,N_5560,N_5483);
and U5608 (N_5608,N_5489,N_5443);
xnor U5609 (N_5609,N_5519,N_5579);
nor U5610 (N_5610,N_5580,N_5481);
or U5611 (N_5611,N_5595,N_5527);
and U5612 (N_5612,N_5478,N_5540);
nand U5613 (N_5613,N_5591,N_5463);
nand U5614 (N_5614,N_5523,N_5528);
nor U5615 (N_5615,N_5496,N_5451);
nand U5616 (N_5616,N_5537,N_5596);
xnor U5617 (N_5617,N_5590,N_5492);
or U5618 (N_5618,N_5462,N_5564);
nor U5619 (N_5619,N_5495,N_5460);
nor U5620 (N_5620,N_5479,N_5456);
and U5621 (N_5621,N_5507,N_5441);
xnor U5622 (N_5622,N_5522,N_5502);
or U5623 (N_5623,N_5573,N_5567);
nand U5624 (N_5624,N_5445,N_5534);
nor U5625 (N_5625,N_5473,N_5525);
nor U5626 (N_5626,N_5529,N_5446);
nand U5627 (N_5627,N_5465,N_5535);
or U5628 (N_5628,N_5578,N_5449);
nand U5629 (N_5629,N_5440,N_5597);
and U5630 (N_5630,N_5532,N_5552);
or U5631 (N_5631,N_5442,N_5485);
xnor U5632 (N_5632,N_5554,N_5471);
and U5633 (N_5633,N_5500,N_5536);
nor U5634 (N_5634,N_5547,N_5541);
xnor U5635 (N_5635,N_5498,N_5542);
xnor U5636 (N_5636,N_5548,N_5521);
and U5637 (N_5637,N_5533,N_5582);
or U5638 (N_5638,N_5553,N_5539);
nand U5639 (N_5639,N_5454,N_5513);
and U5640 (N_5640,N_5549,N_5505);
and U5641 (N_5641,N_5572,N_5531);
or U5642 (N_5642,N_5583,N_5484);
nor U5643 (N_5643,N_5458,N_5474);
nor U5644 (N_5644,N_5464,N_5526);
or U5645 (N_5645,N_5588,N_5503);
nand U5646 (N_5646,N_5516,N_5576);
xnor U5647 (N_5647,N_5559,N_5491);
nand U5648 (N_5648,N_5566,N_5530);
xnor U5649 (N_5649,N_5593,N_5486);
and U5650 (N_5650,N_5558,N_5466);
nor U5651 (N_5651,N_5599,N_5545);
and U5652 (N_5652,N_5514,N_5480);
xnor U5653 (N_5653,N_5509,N_5517);
or U5654 (N_5654,N_5524,N_5561);
xor U5655 (N_5655,N_5598,N_5584);
xor U5656 (N_5656,N_5550,N_5472);
or U5657 (N_5657,N_5459,N_5577);
xor U5658 (N_5658,N_5574,N_5470);
nand U5659 (N_5659,N_5546,N_5457);
or U5660 (N_5660,N_5551,N_5575);
nor U5661 (N_5661,N_5569,N_5452);
xor U5662 (N_5662,N_5476,N_5488);
nand U5663 (N_5663,N_5587,N_5450);
xnor U5664 (N_5664,N_5493,N_5477);
nor U5665 (N_5665,N_5455,N_5544);
nand U5666 (N_5666,N_5555,N_5556);
and U5667 (N_5667,N_5444,N_5563);
and U5668 (N_5668,N_5543,N_5447);
nor U5669 (N_5669,N_5501,N_5562);
nand U5670 (N_5670,N_5469,N_5565);
xor U5671 (N_5671,N_5585,N_5557);
or U5672 (N_5672,N_5570,N_5499);
or U5673 (N_5673,N_5461,N_5589);
and U5674 (N_5674,N_5482,N_5475);
nand U5675 (N_5675,N_5538,N_5594);
nand U5676 (N_5676,N_5571,N_5586);
xor U5677 (N_5677,N_5592,N_5518);
or U5678 (N_5678,N_5506,N_5467);
nand U5679 (N_5679,N_5512,N_5490);
or U5680 (N_5680,N_5504,N_5460);
or U5681 (N_5681,N_5564,N_5501);
xnor U5682 (N_5682,N_5467,N_5544);
nor U5683 (N_5683,N_5529,N_5484);
nand U5684 (N_5684,N_5568,N_5492);
nor U5685 (N_5685,N_5564,N_5590);
nor U5686 (N_5686,N_5547,N_5579);
and U5687 (N_5687,N_5562,N_5536);
nor U5688 (N_5688,N_5568,N_5594);
and U5689 (N_5689,N_5527,N_5557);
or U5690 (N_5690,N_5495,N_5487);
or U5691 (N_5691,N_5536,N_5463);
or U5692 (N_5692,N_5563,N_5470);
nand U5693 (N_5693,N_5572,N_5485);
nor U5694 (N_5694,N_5572,N_5578);
xnor U5695 (N_5695,N_5518,N_5447);
nor U5696 (N_5696,N_5512,N_5531);
nand U5697 (N_5697,N_5545,N_5465);
nand U5698 (N_5698,N_5551,N_5548);
nand U5699 (N_5699,N_5587,N_5529);
nor U5700 (N_5700,N_5485,N_5464);
xor U5701 (N_5701,N_5441,N_5473);
nor U5702 (N_5702,N_5529,N_5471);
and U5703 (N_5703,N_5560,N_5494);
or U5704 (N_5704,N_5455,N_5578);
nor U5705 (N_5705,N_5524,N_5546);
nor U5706 (N_5706,N_5444,N_5587);
xor U5707 (N_5707,N_5462,N_5576);
xnor U5708 (N_5708,N_5599,N_5444);
nand U5709 (N_5709,N_5465,N_5500);
nor U5710 (N_5710,N_5492,N_5518);
and U5711 (N_5711,N_5537,N_5590);
nor U5712 (N_5712,N_5562,N_5471);
and U5713 (N_5713,N_5452,N_5507);
nand U5714 (N_5714,N_5576,N_5494);
nand U5715 (N_5715,N_5554,N_5589);
nand U5716 (N_5716,N_5503,N_5540);
xnor U5717 (N_5717,N_5531,N_5536);
nand U5718 (N_5718,N_5468,N_5516);
and U5719 (N_5719,N_5513,N_5571);
nor U5720 (N_5720,N_5598,N_5503);
and U5721 (N_5721,N_5526,N_5528);
nor U5722 (N_5722,N_5509,N_5481);
or U5723 (N_5723,N_5558,N_5493);
nand U5724 (N_5724,N_5548,N_5586);
and U5725 (N_5725,N_5573,N_5511);
xor U5726 (N_5726,N_5448,N_5533);
nand U5727 (N_5727,N_5562,N_5484);
nor U5728 (N_5728,N_5507,N_5472);
nand U5729 (N_5729,N_5586,N_5500);
nor U5730 (N_5730,N_5591,N_5479);
xnor U5731 (N_5731,N_5507,N_5467);
and U5732 (N_5732,N_5540,N_5553);
nor U5733 (N_5733,N_5450,N_5507);
nor U5734 (N_5734,N_5541,N_5487);
nand U5735 (N_5735,N_5476,N_5574);
xnor U5736 (N_5736,N_5562,N_5561);
or U5737 (N_5737,N_5594,N_5471);
nor U5738 (N_5738,N_5517,N_5546);
xor U5739 (N_5739,N_5451,N_5581);
nand U5740 (N_5740,N_5578,N_5514);
and U5741 (N_5741,N_5537,N_5566);
nor U5742 (N_5742,N_5539,N_5469);
xor U5743 (N_5743,N_5578,N_5553);
or U5744 (N_5744,N_5597,N_5558);
and U5745 (N_5745,N_5598,N_5478);
nor U5746 (N_5746,N_5513,N_5458);
nand U5747 (N_5747,N_5597,N_5534);
and U5748 (N_5748,N_5560,N_5593);
and U5749 (N_5749,N_5523,N_5535);
xor U5750 (N_5750,N_5474,N_5490);
nor U5751 (N_5751,N_5465,N_5523);
and U5752 (N_5752,N_5578,N_5590);
nand U5753 (N_5753,N_5506,N_5515);
and U5754 (N_5754,N_5576,N_5565);
nand U5755 (N_5755,N_5536,N_5464);
xnor U5756 (N_5756,N_5462,N_5445);
or U5757 (N_5757,N_5518,N_5499);
nor U5758 (N_5758,N_5593,N_5499);
nor U5759 (N_5759,N_5525,N_5450);
xor U5760 (N_5760,N_5739,N_5609);
nand U5761 (N_5761,N_5725,N_5605);
xor U5762 (N_5762,N_5654,N_5625);
xnor U5763 (N_5763,N_5669,N_5620);
nor U5764 (N_5764,N_5626,N_5702);
or U5765 (N_5765,N_5735,N_5617);
or U5766 (N_5766,N_5743,N_5731);
nand U5767 (N_5767,N_5699,N_5667);
nand U5768 (N_5768,N_5672,N_5656);
and U5769 (N_5769,N_5757,N_5643);
or U5770 (N_5770,N_5621,N_5631);
nand U5771 (N_5771,N_5646,N_5706);
nor U5772 (N_5772,N_5710,N_5634);
nor U5773 (N_5773,N_5641,N_5652);
nor U5774 (N_5774,N_5683,N_5622);
or U5775 (N_5775,N_5696,N_5693);
xnor U5776 (N_5776,N_5687,N_5684);
nor U5777 (N_5777,N_5653,N_5613);
nor U5778 (N_5778,N_5749,N_5727);
and U5779 (N_5779,N_5633,N_5750);
or U5780 (N_5780,N_5677,N_5737);
nor U5781 (N_5781,N_5741,N_5637);
or U5782 (N_5782,N_5648,N_5651);
and U5783 (N_5783,N_5628,N_5742);
xor U5784 (N_5784,N_5675,N_5665);
and U5785 (N_5785,N_5714,N_5688);
or U5786 (N_5786,N_5666,N_5748);
nor U5787 (N_5787,N_5718,N_5670);
nand U5788 (N_5788,N_5671,N_5676);
nand U5789 (N_5789,N_5717,N_5645);
nor U5790 (N_5790,N_5673,N_5664);
nor U5791 (N_5791,N_5638,N_5623);
nor U5792 (N_5792,N_5612,N_5619);
or U5793 (N_5793,N_5630,N_5657);
and U5794 (N_5794,N_5627,N_5650);
or U5795 (N_5795,N_5695,N_5719);
or U5796 (N_5796,N_5690,N_5618);
and U5797 (N_5797,N_5658,N_5660);
or U5798 (N_5798,N_5711,N_5635);
or U5799 (N_5799,N_5709,N_5639);
nand U5800 (N_5800,N_5746,N_5624);
nor U5801 (N_5801,N_5682,N_5734);
or U5802 (N_5802,N_5722,N_5640);
and U5803 (N_5803,N_5659,N_5751);
or U5804 (N_5804,N_5655,N_5756);
xor U5805 (N_5805,N_5611,N_5733);
and U5806 (N_5806,N_5694,N_5712);
and U5807 (N_5807,N_5698,N_5680);
or U5808 (N_5808,N_5663,N_5661);
and U5809 (N_5809,N_5668,N_5728);
and U5810 (N_5810,N_5715,N_5610);
nor U5811 (N_5811,N_5723,N_5755);
and U5812 (N_5812,N_5704,N_5721);
nor U5813 (N_5813,N_5729,N_5685);
or U5814 (N_5814,N_5615,N_5679);
nor U5815 (N_5815,N_5744,N_5607);
and U5816 (N_5816,N_5732,N_5700);
nor U5817 (N_5817,N_5697,N_5616);
and U5818 (N_5818,N_5629,N_5708);
xnor U5819 (N_5819,N_5642,N_5745);
nor U5820 (N_5820,N_5738,N_5703);
or U5821 (N_5821,N_5692,N_5686);
or U5822 (N_5822,N_5736,N_5636);
nand U5823 (N_5823,N_5604,N_5600);
nand U5824 (N_5824,N_5603,N_5747);
nand U5825 (N_5825,N_5662,N_5753);
or U5826 (N_5826,N_5602,N_5730);
and U5827 (N_5827,N_5754,N_5707);
xor U5828 (N_5828,N_5759,N_5681);
nor U5829 (N_5829,N_5720,N_5608);
xnor U5830 (N_5830,N_5606,N_5632);
and U5831 (N_5831,N_5678,N_5713);
nor U5832 (N_5832,N_5758,N_5644);
xnor U5833 (N_5833,N_5614,N_5740);
xnor U5834 (N_5834,N_5716,N_5724);
nand U5835 (N_5835,N_5705,N_5701);
and U5836 (N_5836,N_5649,N_5647);
xor U5837 (N_5837,N_5601,N_5689);
or U5838 (N_5838,N_5752,N_5726);
xnor U5839 (N_5839,N_5691,N_5674);
or U5840 (N_5840,N_5740,N_5636);
and U5841 (N_5841,N_5756,N_5659);
nand U5842 (N_5842,N_5700,N_5665);
and U5843 (N_5843,N_5738,N_5650);
xor U5844 (N_5844,N_5670,N_5719);
nand U5845 (N_5845,N_5613,N_5711);
nand U5846 (N_5846,N_5608,N_5664);
xor U5847 (N_5847,N_5713,N_5716);
nand U5848 (N_5848,N_5716,N_5688);
nand U5849 (N_5849,N_5657,N_5713);
nand U5850 (N_5850,N_5673,N_5601);
nand U5851 (N_5851,N_5615,N_5614);
xor U5852 (N_5852,N_5748,N_5736);
nand U5853 (N_5853,N_5713,N_5618);
nand U5854 (N_5854,N_5685,N_5720);
and U5855 (N_5855,N_5672,N_5624);
or U5856 (N_5856,N_5613,N_5647);
nor U5857 (N_5857,N_5628,N_5640);
nor U5858 (N_5858,N_5630,N_5660);
and U5859 (N_5859,N_5656,N_5622);
or U5860 (N_5860,N_5617,N_5665);
and U5861 (N_5861,N_5747,N_5726);
or U5862 (N_5862,N_5637,N_5738);
xor U5863 (N_5863,N_5682,N_5665);
and U5864 (N_5864,N_5659,N_5736);
nand U5865 (N_5865,N_5671,N_5690);
nor U5866 (N_5866,N_5639,N_5740);
nand U5867 (N_5867,N_5611,N_5665);
nand U5868 (N_5868,N_5676,N_5649);
and U5869 (N_5869,N_5722,N_5637);
nand U5870 (N_5870,N_5695,N_5721);
nand U5871 (N_5871,N_5723,N_5753);
nand U5872 (N_5872,N_5638,N_5625);
or U5873 (N_5873,N_5704,N_5665);
xnor U5874 (N_5874,N_5614,N_5742);
nand U5875 (N_5875,N_5752,N_5713);
nor U5876 (N_5876,N_5694,N_5720);
nor U5877 (N_5877,N_5693,N_5675);
xnor U5878 (N_5878,N_5636,N_5733);
nor U5879 (N_5879,N_5707,N_5732);
nor U5880 (N_5880,N_5626,N_5749);
nor U5881 (N_5881,N_5602,N_5648);
or U5882 (N_5882,N_5741,N_5617);
or U5883 (N_5883,N_5601,N_5710);
xnor U5884 (N_5884,N_5718,N_5758);
or U5885 (N_5885,N_5731,N_5618);
nor U5886 (N_5886,N_5718,N_5687);
or U5887 (N_5887,N_5726,N_5657);
nor U5888 (N_5888,N_5650,N_5724);
xor U5889 (N_5889,N_5667,N_5728);
and U5890 (N_5890,N_5681,N_5724);
nor U5891 (N_5891,N_5605,N_5723);
xnor U5892 (N_5892,N_5707,N_5619);
nand U5893 (N_5893,N_5681,N_5684);
nor U5894 (N_5894,N_5720,N_5745);
nand U5895 (N_5895,N_5742,N_5601);
nor U5896 (N_5896,N_5706,N_5703);
nor U5897 (N_5897,N_5682,N_5654);
and U5898 (N_5898,N_5748,N_5702);
nor U5899 (N_5899,N_5613,N_5625);
nor U5900 (N_5900,N_5629,N_5626);
xnor U5901 (N_5901,N_5676,N_5735);
xnor U5902 (N_5902,N_5695,N_5677);
and U5903 (N_5903,N_5608,N_5621);
xnor U5904 (N_5904,N_5618,N_5614);
xor U5905 (N_5905,N_5605,N_5742);
xnor U5906 (N_5906,N_5636,N_5726);
and U5907 (N_5907,N_5651,N_5695);
xnor U5908 (N_5908,N_5613,N_5627);
nand U5909 (N_5909,N_5710,N_5698);
or U5910 (N_5910,N_5646,N_5681);
nand U5911 (N_5911,N_5684,N_5616);
xor U5912 (N_5912,N_5724,N_5730);
xor U5913 (N_5913,N_5678,N_5668);
xor U5914 (N_5914,N_5736,N_5710);
xnor U5915 (N_5915,N_5723,N_5738);
or U5916 (N_5916,N_5612,N_5653);
and U5917 (N_5917,N_5660,N_5605);
and U5918 (N_5918,N_5720,N_5689);
or U5919 (N_5919,N_5727,N_5651);
xor U5920 (N_5920,N_5858,N_5829);
and U5921 (N_5921,N_5814,N_5796);
and U5922 (N_5922,N_5806,N_5852);
xor U5923 (N_5923,N_5914,N_5841);
xnor U5924 (N_5924,N_5873,N_5916);
or U5925 (N_5925,N_5804,N_5878);
nand U5926 (N_5926,N_5785,N_5812);
or U5927 (N_5927,N_5893,N_5815);
nor U5928 (N_5928,N_5890,N_5898);
or U5929 (N_5929,N_5882,N_5854);
xor U5930 (N_5930,N_5847,N_5883);
xor U5931 (N_5931,N_5781,N_5911);
xor U5932 (N_5932,N_5813,N_5855);
xor U5933 (N_5933,N_5903,N_5770);
xor U5934 (N_5934,N_5799,N_5767);
nand U5935 (N_5935,N_5792,N_5768);
or U5936 (N_5936,N_5798,N_5809);
nand U5937 (N_5937,N_5877,N_5889);
or U5938 (N_5938,N_5825,N_5848);
nor U5939 (N_5939,N_5902,N_5900);
nor U5940 (N_5940,N_5778,N_5771);
xor U5941 (N_5941,N_5840,N_5836);
nor U5942 (N_5942,N_5800,N_5761);
and U5943 (N_5943,N_5888,N_5894);
nor U5944 (N_5944,N_5786,N_5795);
nor U5945 (N_5945,N_5919,N_5850);
nand U5946 (N_5946,N_5896,N_5760);
or U5947 (N_5947,N_5834,N_5784);
and U5948 (N_5948,N_5915,N_5872);
and U5949 (N_5949,N_5762,N_5886);
nand U5950 (N_5950,N_5822,N_5862);
nor U5951 (N_5951,N_5803,N_5909);
and U5952 (N_5952,N_5791,N_5772);
xnor U5953 (N_5953,N_5861,N_5763);
or U5954 (N_5954,N_5827,N_5777);
nor U5955 (N_5955,N_5764,N_5787);
nor U5956 (N_5956,N_5846,N_5776);
nand U5957 (N_5957,N_5790,N_5913);
xnor U5958 (N_5958,N_5807,N_5856);
xor U5959 (N_5959,N_5899,N_5870);
nor U5960 (N_5960,N_5793,N_5810);
and U5961 (N_5961,N_5816,N_5875);
xor U5962 (N_5962,N_5766,N_5904);
xnor U5963 (N_5963,N_5811,N_5851);
nor U5964 (N_5964,N_5892,N_5908);
or U5965 (N_5965,N_5887,N_5783);
or U5966 (N_5966,N_5818,N_5833);
and U5967 (N_5967,N_5769,N_5906);
or U5968 (N_5968,N_5794,N_5830);
nor U5969 (N_5969,N_5788,N_5837);
xnor U5970 (N_5970,N_5839,N_5845);
and U5971 (N_5971,N_5857,N_5901);
nand U5972 (N_5972,N_5864,N_5917);
xor U5973 (N_5973,N_5779,N_5895);
nand U5974 (N_5974,N_5835,N_5775);
nand U5975 (N_5975,N_5808,N_5871);
xor U5976 (N_5976,N_5918,N_5819);
nand U5977 (N_5977,N_5824,N_5831);
or U5978 (N_5978,N_5823,N_5912);
nand U5979 (N_5979,N_5843,N_5821);
and U5980 (N_5980,N_5884,N_5879);
and U5981 (N_5981,N_5860,N_5838);
nor U5982 (N_5982,N_5826,N_5885);
and U5983 (N_5983,N_5817,N_5820);
xor U5984 (N_5984,N_5853,N_5802);
nand U5985 (N_5985,N_5876,N_5844);
nor U5986 (N_5986,N_5774,N_5867);
nand U5987 (N_5987,N_5866,N_5881);
xor U5988 (N_5988,N_5880,N_5891);
or U5989 (N_5989,N_5865,N_5868);
and U5990 (N_5990,N_5780,N_5828);
and U5991 (N_5991,N_5765,N_5874);
nand U5992 (N_5992,N_5773,N_5859);
nand U5993 (N_5993,N_5789,N_5910);
xor U5994 (N_5994,N_5897,N_5849);
and U5995 (N_5995,N_5863,N_5869);
xnor U5996 (N_5996,N_5801,N_5842);
or U5997 (N_5997,N_5907,N_5782);
or U5998 (N_5998,N_5805,N_5905);
and U5999 (N_5999,N_5797,N_5832);
xnor U6000 (N_6000,N_5765,N_5914);
and U6001 (N_6001,N_5779,N_5813);
xnor U6002 (N_6002,N_5857,N_5813);
nor U6003 (N_6003,N_5850,N_5873);
nor U6004 (N_6004,N_5864,N_5879);
or U6005 (N_6005,N_5900,N_5885);
xor U6006 (N_6006,N_5845,N_5780);
nand U6007 (N_6007,N_5789,N_5851);
xnor U6008 (N_6008,N_5823,N_5846);
nand U6009 (N_6009,N_5842,N_5788);
nor U6010 (N_6010,N_5910,N_5905);
xor U6011 (N_6011,N_5906,N_5885);
nor U6012 (N_6012,N_5836,N_5809);
or U6013 (N_6013,N_5822,N_5864);
and U6014 (N_6014,N_5843,N_5888);
and U6015 (N_6015,N_5838,N_5764);
or U6016 (N_6016,N_5795,N_5852);
nand U6017 (N_6017,N_5836,N_5812);
xnor U6018 (N_6018,N_5917,N_5771);
nand U6019 (N_6019,N_5855,N_5831);
xnor U6020 (N_6020,N_5897,N_5829);
and U6021 (N_6021,N_5917,N_5796);
nor U6022 (N_6022,N_5832,N_5811);
nand U6023 (N_6023,N_5851,N_5902);
or U6024 (N_6024,N_5917,N_5880);
xnor U6025 (N_6025,N_5874,N_5766);
xor U6026 (N_6026,N_5853,N_5847);
nor U6027 (N_6027,N_5817,N_5865);
nor U6028 (N_6028,N_5862,N_5840);
nand U6029 (N_6029,N_5919,N_5865);
and U6030 (N_6030,N_5843,N_5912);
xnor U6031 (N_6031,N_5844,N_5917);
or U6032 (N_6032,N_5859,N_5805);
or U6033 (N_6033,N_5832,N_5886);
or U6034 (N_6034,N_5798,N_5901);
nand U6035 (N_6035,N_5903,N_5839);
and U6036 (N_6036,N_5894,N_5813);
nor U6037 (N_6037,N_5826,N_5833);
xor U6038 (N_6038,N_5779,N_5796);
and U6039 (N_6039,N_5841,N_5769);
or U6040 (N_6040,N_5917,N_5905);
nor U6041 (N_6041,N_5902,N_5812);
nor U6042 (N_6042,N_5795,N_5813);
nor U6043 (N_6043,N_5784,N_5840);
nor U6044 (N_6044,N_5816,N_5836);
or U6045 (N_6045,N_5781,N_5859);
and U6046 (N_6046,N_5852,N_5803);
nor U6047 (N_6047,N_5801,N_5784);
or U6048 (N_6048,N_5879,N_5843);
and U6049 (N_6049,N_5778,N_5797);
xnor U6050 (N_6050,N_5766,N_5854);
or U6051 (N_6051,N_5888,N_5835);
or U6052 (N_6052,N_5791,N_5811);
or U6053 (N_6053,N_5876,N_5909);
or U6054 (N_6054,N_5836,N_5876);
nand U6055 (N_6055,N_5840,N_5813);
and U6056 (N_6056,N_5781,N_5898);
xnor U6057 (N_6057,N_5778,N_5768);
nor U6058 (N_6058,N_5831,N_5766);
nor U6059 (N_6059,N_5894,N_5766);
and U6060 (N_6060,N_5861,N_5913);
nand U6061 (N_6061,N_5763,N_5810);
and U6062 (N_6062,N_5802,N_5851);
or U6063 (N_6063,N_5904,N_5868);
nand U6064 (N_6064,N_5851,N_5899);
and U6065 (N_6065,N_5810,N_5789);
xnor U6066 (N_6066,N_5807,N_5803);
nor U6067 (N_6067,N_5904,N_5815);
and U6068 (N_6068,N_5846,N_5879);
nand U6069 (N_6069,N_5838,N_5843);
nand U6070 (N_6070,N_5863,N_5896);
or U6071 (N_6071,N_5863,N_5806);
nor U6072 (N_6072,N_5890,N_5799);
and U6073 (N_6073,N_5903,N_5842);
and U6074 (N_6074,N_5845,N_5825);
nand U6075 (N_6075,N_5797,N_5891);
nand U6076 (N_6076,N_5862,N_5878);
and U6077 (N_6077,N_5801,N_5906);
xor U6078 (N_6078,N_5850,N_5801);
nand U6079 (N_6079,N_5876,N_5807);
or U6080 (N_6080,N_6076,N_5970);
nor U6081 (N_6081,N_5948,N_6041);
xnor U6082 (N_6082,N_6050,N_5978);
and U6083 (N_6083,N_6056,N_5994);
xnor U6084 (N_6084,N_5965,N_6045);
and U6085 (N_6085,N_5934,N_6040);
nor U6086 (N_6086,N_5993,N_6072);
and U6087 (N_6087,N_5984,N_5946);
xnor U6088 (N_6088,N_5942,N_6062);
and U6089 (N_6089,N_5938,N_6068);
and U6090 (N_6090,N_5976,N_5931);
or U6091 (N_6091,N_5921,N_5985);
xor U6092 (N_6092,N_5964,N_5952);
nand U6093 (N_6093,N_5924,N_5979);
and U6094 (N_6094,N_6039,N_6031);
and U6095 (N_6095,N_5928,N_5959);
or U6096 (N_6096,N_6003,N_5932);
or U6097 (N_6097,N_5926,N_6019);
or U6098 (N_6098,N_6022,N_6069);
nand U6099 (N_6099,N_6002,N_6007);
nor U6100 (N_6100,N_6024,N_5977);
xor U6101 (N_6101,N_6027,N_5935);
nor U6102 (N_6102,N_5949,N_5958);
nand U6103 (N_6103,N_6052,N_6044);
and U6104 (N_6104,N_6063,N_6008);
nand U6105 (N_6105,N_5943,N_5940);
or U6106 (N_6106,N_5922,N_5953);
xor U6107 (N_6107,N_5963,N_6079);
xor U6108 (N_6108,N_5999,N_6070);
nand U6109 (N_6109,N_5933,N_6033);
and U6110 (N_6110,N_6035,N_5951);
nand U6111 (N_6111,N_6053,N_6061);
nand U6112 (N_6112,N_6048,N_5941);
nor U6113 (N_6113,N_6054,N_5937);
and U6114 (N_6114,N_6025,N_6004);
xor U6115 (N_6115,N_5968,N_5986);
or U6116 (N_6116,N_5966,N_6037);
nand U6117 (N_6117,N_5956,N_5936);
nor U6118 (N_6118,N_6043,N_5925);
nand U6119 (N_6119,N_6057,N_5991);
xnor U6120 (N_6120,N_5955,N_5971);
nand U6121 (N_6121,N_6074,N_6030);
xnor U6122 (N_6122,N_6012,N_5927);
or U6123 (N_6123,N_6001,N_5957);
nor U6124 (N_6124,N_6028,N_5975);
or U6125 (N_6125,N_5982,N_6059);
or U6126 (N_6126,N_6009,N_6073);
nand U6127 (N_6127,N_5973,N_6049);
and U6128 (N_6128,N_5990,N_6005);
nand U6129 (N_6129,N_6036,N_6065);
or U6130 (N_6130,N_6077,N_6000);
xnor U6131 (N_6131,N_6021,N_6032);
nand U6132 (N_6132,N_5998,N_6064);
or U6133 (N_6133,N_5939,N_6023);
or U6134 (N_6134,N_5983,N_6067);
or U6135 (N_6135,N_6011,N_6017);
nand U6136 (N_6136,N_5997,N_6034);
nand U6137 (N_6137,N_6029,N_5967);
or U6138 (N_6138,N_5969,N_5947);
xor U6139 (N_6139,N_6047,N_5988);
xor U6140 (N_6140,N_6015,N_5980);
nor U6141 (N_6141,N_5972,N_6038);
xor U6142 (N_6142,N_6013,N_5961);
nand U6143 (N_6143,N_5944,N_5954);
xnor U6144 (N_6144,N_6051,N_5962);
nor U6145 (N_6145,N_5992,N_6026);
or U6146 (N_6146,N_5923,N_6006);
or U6147 (N_6147,N_5920,N_6071);
and U6148 (N_6148,N_6058,N_5996);
or U6149 (N_6149,N_5960,N_6055);
nand U6150 (N_6150,N_5950,N_5930);
xor U6151 (N_6151,N_5995,N_5981);
and U6152 (N_6152,N_5974,N_6016);
nor U6153 (N_6153,N_6010,N_6060);
and U6154 (N_6154,N_6014,N_6020);
nand U6155 (N_6155,N_5987,N_5929);
and U6156 (N_6156,N_6018,N_5945);
xor U6157 (N_6157,N_5989,N_6046);
or U6158 (N_6158,N_6066,N_6075);
nor U6159 (N_6159,N_6042,N_6078);
nor U6160 (N_6160,N_5938,N_6065);
or U6161 (N_6161,N_6023,N_6005);
xnor U6162 (N_6162,N_6026,N_6050);
nor U6163 (N_6163,N_6037,N_6077);
and U6164 (N_6164,N_5955,N_6070);
or U6165 (N_6165,N_5985,N_5988);
nor U6166 (N_6166,N_6063,N_6001);
xnor U6167 (N_6167,N_6025,N_6021);
and U6168 (N_6168,N_5996,N_6044);
or U6169 (N_6169,N_5985,N_6055);
and U6170 (N_6170,N_5941,N_5922);
or U6171 (N_6171,N_5992,N_6037);
and U6172 (N_6172,N_6008,N_5976);
or U6173 (N_6173,N_5920,N_6046);
xor U6174 (N_6174,N_6066,N_6068);
and U6175 (N_6175,N_5925,N_6008);
and U6176 (N_6176,N_6052,N_6046);
or U6177 (N_6177,N_5956,N_5951);
xor U6178 (N_6178,N_6019,N_6013);
nand U6179 (N_6179,N_5932,N_5968);
or U6180 (N_6180,N_6050,N_5959);
and U6181 (N_6181,N_5988,N_5930);
and U6182 (N_6182,N_6061,N_5963);
xnor U6183 (N_6183,N_6016,N_6007);
xnor U6184 (N_6184,N_6066,N_6071);
or U6185 (N_6185,N_6021,N_5990);
xnor U6186 (N_6186,N_6055,N_6041);
or U6187 (N_6187,N_6046,N_6073);
and U6188 (N_6188,N_5972,N_5970);
xnor U6189 (N_6189,N_5938,N_6008);
and U6190 (N_6190,N_5924,N_6038);
or U6191 (N_6191,N_5929,N_6023);
xnor U6192 (N_6192,N_5973,N_5950);
nand U6193 (N_6193,N_6056,N_6001);
nor U6194 (N_6194,N_6015,N_6074);
nand U6195 (N_6195,N_5964,N_5943);
nor U6196 (N_6196,N_5922,N_5925);
nor U6197 (N_6197,N_5939,N_6006);
xnor U6198 (N_6198,N_5947,N_6057);
nand U6199 (N_6199,N_6028,N_5984);
and U6200 (N_6200,N_5980,N_6057);
xor U6201 (N_6201,N_5979,N_5933);
and U6202 (N_6202,N_6051,N_6073);
nor U6203 (N_6203,N_6038,N_5938);
and U6204 (N_6204,N_5972,N_6027);
nor U6205 (N_6205,N_6077,N_6032);
or U6206 (N_6206,N_6000,N_5976);
and U6207 (N_6207,N_6013,N_6079);
or U6208 (N_6208,N_5975,N_6002);
and U6209 (N_6209,N_5948,N_5975);
and U6210 (N_6210,N_5937,N_6005);
nor U6211 (N_6211,N_6056,N_5932);
xor U6212 (N_6212,N_5941,N_6012);
and U6213 (N_6213,N_6046,N_6010);
nor U6214 (N_6214,N_6010,N_6037);
nand U6215 (N_6215,N_5990,N_6010);
xnor U6216 (N_6216,N_6003,N_6020);
nand U6217 (N_6217,N_5940,N_5946);
nor U6218 (N_6218,N_6018,N_5924);
nand U6219 (N_6219,N_5954,N_6015);
xor U6220 (N_6220,N_5941,N_5959);
and U6221 (N_6221,N_6013,N_6022);
xnor U6222 (N_6222,N_5946,N_5987);
and U6223 (N_6223,N_5955,N_5968);
nor U6224 (N_6224,N_5963,N_6036);
nand U6225 (N_6225,N_5966,N_6005);
or U6226 (N_6226,N_6056,N_5974);
xnor U6227 (N_6227,N_6045,N_5997);
nor U6228 (N_6228,N_5964,N_6030);
or U6229 (N_6229,N_6052,N_5947);
or U6230 (N_6230,N_6000,N_5968);
nor U6231 (N_6231,N_6044,N_5981);
and U6232 (N_6232,N_5995,N_5987);
nand U6233 (N_6233,N_5922,N_5956);
and U6234 (N_6234,N_6010,N_6062);
or U6235 (N_6235,N_6055,N_5947);
or U6236 (N_6236,N_6007,N_5960);
or U6237 (N_6237,N_5950,N_5997);
or U6238 (N_6238,N_5951,N_5992);
nor U6239 (N_6239,N_5923,N_5953);
and U6240 (N_6240,N_6113,N_6201);
xnor U6241 (N_6241,N_6138,N_6107);
or U6242 (N_6242,N_6163,N_6185);
and U6243 (N_6243,N_6217,N_6187);
or U6244 (N_6244,N_6146,N_6101);
or U6245 (N_6245,N_6196,N_6143);
or U6246 (N_6246,N_6086,N_6115);
xor U6247 (N_6247,N_6127,N_6211);
xor U6248 (N_6248,N_6102,N_6093);
nand U6249 (N_6249,N_6083,N_6198);
or U6250 (N_6250,N_6117,N_6150);
xor U6251 (N_6251,N_6091,N_6237);
xor U6252 (N_6252,N_6154,N_6189);
and U6253 (N_6253,N_6088,N_6195);
or U6254 (N_6254,N_6109,N_6222);
nand U6255 (N_6255,N_6145,N_6200);
xor U6256 (N_6256,N_6188,N_6202);
nand U6257 (N_6257,N_6173,N_6136);
nor U6258 (N_6258,N_6218,N_6129);
and U6259 (N_6259,N_6206,N_6183);
and U6260 (N_6260,N_6179,N_6209);
nor U6261 (N_6261,N_6157,N_6124);
nor U6262 (N_6262,N_6172,N_6090);
xor U6263 (N_6263,N_6223,N_6147);
nor U6264 (N_6264,N_6190,N_6126);
nand U6265 (N_6265,N_6153,N_6235);
and U6266 (N_6266,N_6155,N_6122);
xor U6267 (N_6267,N_6132,N_6212);
or U6268 (N_6268,N_6181,N_6215);
or U6269 (N_6269,N_6229,N_6207);
nand U6270 (N_6270,N_6168,N_6148);
xor U6271 (N_6271,N_6213,N_6110);
and U6272 (N_6272,N_6084,N_6118);
or U6273 (N_6273,N_6192,N_6231);
nand U6274 (N_6274,N_6099,N_6175);
or U6275 (N_6275,N_6162,N_6100);
nor U6276 (N_6276,N_6139,N_6226);
and U6277 (N_6277,N_6186,N_6120);
nand U6278 (N_6278,N_6210,N_6141);
or U6279 (N_6279,N_6177,N_6149);
nor U6280 (N_6280,N_6197,N_6097);
xor U6281 (N_6281,N_6236,N_6089);
nor U6282 (N_6282,N_6178,N_6135);
nor U6283 (N_6283,N_6142,N_6131);
nor U6284 (N_6284,N_6080,N_6214);
and U6285 (N_6285,N_6199,N_6152);
and U6286 (N_6286,N_6105,N_6161);
nor U6287 (N_6287,N_6221,N_6121);
and U6288 (N_6288,N_6230,N_6116);
and U6289 (N_6289,N_6176,N_6219);
xor U6290 (N_6290,N_6140,N_6158);
nand U6291 (N_6291,N_6194,N_6232);
and U6292 (N_6292,N_6166,N_6239);
xnor U6293 (N_6293,N_6167,N_6106);
nand U6294 (N_6294,N_6238,N_6111);
and U6295 (N_6295,N_6169,N_6160);
xor U6296 (N_6296,N_6159,N_6191);
xnor U6297 (N_6297,N_6227,N_6108);
xnor U6298 (N_6298,N_6096,N_6092);
or U6299 (N_6299,N_6225,N_6208);
nor U6300 (N_6300,N_6228,N_6234);
nor U6301 (N_6301,N_6220,N_6174);
or U6302 (N_6302,N_6233,N_6125);
nor U6303 (N_6303,N_6204,N_6184);
nor U6304 (N_6304,N_6180,N_6137);
xor U6305 (N_6305,N_6164,N_6203);
nand U6306 (N_6306,N_6151,N_6095);
and U6307 (N_6307,N_6123,N_6165);
xnor U6308 (N_6308,N_6104,N_6171);
xnor U6309 (N_6309,N_6224,N_6144);
nand U6310 (N_6310,N_6098,N_6133);
or U6311 (N_6311,N_6103,N_6114);
and U6312 (N_6312,N_6119,N_6081);
nand U6313 (N_6313,N_6085,N_6134);
and U6314 (N_6314,N_6087,N_6216);
nor U6315 (N_6315,N_6128,N_6170);
and U6316 (N_6316,N_6205,N_6094);
xnor U6317 (N_6317,N_6112,N_6156);
or U6318 (N_6318,N_6193,N_6082);
xor U6319 (N_6319,N_6182,N_6130);
or U6320 (N_6320,N_6082,N_6136);
xor U6321 (N_6321,N_6140,N_6108);
nand U6322 (N_6322,N_6123,N_6087);
or U6323 (N_6323,N_6111,N_6117);
xor U6324 (N_6324,N_6206,N_6215);
nor U6325 (N_6325,N_6156,N_6145);
xor U6326 (N_6326,N_6146,N_6164);
xor U6327 (N_6327,N_6114,N_6112);
or U6328 (N_6328,N_6080,N_6082);
nand U6329 (N_6329,N_6144,N_6119);
nor U6330 (N_6330,N_6184,N_6225);
or U6331 (N_6331,N_6167,N_6218);
and U6332 (N_6332,N_6208,N_6107);
nand U6333 (N_6333,N_6222,N_6166);
nand U6334 (N_6334,N_6120,N_6194);
nand U6335 (N_6335,N_6221,N_6107);
and U6336 (N_6336,N_6164,N_6209);
xor U6337 (N_6337,N_6211,N_6228);
and U6338 (N_6338,N_6213,N_6186);
xnor U6339 (N_6339,N_6168,N_6215);
xnor U6340 (N_6340,N_6209,N_6231);
and U6341 (N_6341,N_6155,N_6198);
xor U6342 (N_6342,N_6089,N_6138);
or U6343 (N_6343,N_6100,N_6222);
nand U6344 (N_6344,N_6134,N_6225);
or U6345 (N_6345,N_6171,N_6120);
xor U6346 (N_6346,N_6186,N_6087);
xor U6347 (N_6347,N_6149,N_6160);
nor U6348 (N_6348,N_6130,N_6219);
or U6349 (N_6349,N_6082,N_6225);
and U6350 (N_6350,N_6213,N_6091);
nand U6351 (N_6351,N_6237,N_6176);
nor U6352 (N_6352,N_6126,N_6161);
nor U6353 (N_6353,N_6100,N_6191);
xnor U6354 (N_6354,N_6179,N_6103);
nor U6355 (N_6355,N_6158,N_6236);
nor U6356 (N_6356,N_6207,N_6224);
or U6357 (N_6357,N_6131,N_6080);
xnor U6358 (N_6358,N_6197,N_6163);
and U6359 (N_6359,N_6126,N_6169);
nor U6360 (N_6360,N_6208,N_6163);
or U6361 (N_6361,N_6141,N_6145);
nor U6362 (N_6362,N_6219,N_6141);
nand U6363 (N_6363,N_6122,N_6180);
nand U6364 (N_6364,N_6090,N_6196);
or U6365 (N_6365,N_6209,N_6109);
nand U6366 (N_6366,N_6120,N_6109);
nor U6367 (N_6367,N_6125,N_6166);
and U6368 (N_6368,N_6138,N_6234);
nand U6369 (N_6369,N_6158,N_6111);
and U6370 (N_6370,N_6233,N_6219);
nand U6371 (N_6371,N_6203,N_6124);
and U6372 (N_6372,N_6238,N_6187);
nand U6373 (N_6373,N_6086,N_6212);
nand U6374 (N_6374,N_6193,N_6156);
nor U6375 (N_6375,N_6109,N_6198);
xor U6376 (N_6376,N_6130,N_6166);
or U6377 (N_6377,N_6105,N_6210);
and U6378 (N_6378,N_6201,N_6128);
and U6379 (N_6379,N_6143,N_6183);
or U6380 (N_6380,N_6114,N_6169);
nand U6381 (N_6381,N_6148,N_6187);
nand U6382 (N_6382,N_6215,N_6194);
xor U6383 (N_6383,N_6114,N_6226);
nand U6384 (N_6384,N_6089,N_6140);
xor U6385 (N_6385,N_6160,N_6138);
nor U6386 (N_6386,N_6187,N_6085);
nand U6387 (N_6387,N_6231,N_6174);
or U6388 (N_6388,N_6193,N_6121);
xor U6389 (N_6389,N_6210,N_6122);
nor U6390 (N_6390,N_6234,N_6139);
nor U6391 (N_6391,N_6096,N_6200);
xnor U6392 (N_6392,N_6111,N_6174);
or U6393 (N_6393,N_6231,N_6107);
xor U6394 (N_6394,N_6162,N_6157);
or U6395 (N_6395,N_6182,N_6189);
xnor U6396 (N_6396,N_6099,N_6193);
nand U6397 (N_6397,N_6123,N_6210);
xor U6398 (N_6398,N_6152,N_6233);
or U6399 (N_6399,N_6136,N_6154);
nand U6400 (N_6400,N_6325,N_6319);
and U6401 (N_6401,N_6350,N_6278);
or U6402 (N_6402,N_6361,N_6302);
nor U6403 (N_6403,N_6253,N_6348);
and U6404 (N_6404,N_6321,N_6250);
xor U6405 (N_6405,N_6313,N_6264);
xnor U6406 (N_6406,N_6341,N_6267);
xnor U6407 (N_6407,N_6329,N_6291);
nor U6408 (N_6408,N_6293,N_6245);
xnor U6409 (N_6409,N_6330,N_6399);
and U6410 (N_6410,N_6275,N_6266);
and U6411 (N_6411,N_6339,N_6360);
and U6412 (N_6412,N_6284,N_6377);
nor U6413 (N_6413,N_6337,N_6340);
nor U6414 (N_6414,N_6323,N_6298);
and U6415 (N_6415,N_6391,N_6347);
nor U6416 (N_6416,N_6270,N_6306);
and U6417 (N_6417,N_6381,N_6255);
nor U6418 (N_6418,N_6285,N_6286);
nand U6419 (N_6419,N_6297,N_6371);
nand U6420 (N_6420,N_6390,N_6367);
nand U6421 (N_6421,N_6261,N_6307);
nor U6422 (N_6422,N_6383,N_6276);
and U6423 (N_6423,N_6300,N_6355);
nand U6424 (N_6424,N_6343,N_6310);
xnor U6425 (N_6425,N_6395,N_6331);
or U6426 (N_6426,N_6356,N_6254);
nor U6427 (N_6427,N_6387,N_6320);
or U6428 (N_6428,N_6370,N_6246);
xor U6429 (N_6429,N_6368,N_6338);
xnor U6430 (N_6430,N_6296,N_6256);
or U6431 (N_6431,N_6259,N_6268);
nor U6432 (N_6432,N_6389,N_6375);
xnor U6433 (N_6433,N_6362,N_6366);
xor U6434 (N_6434,N_6369,N_6384);
xnor U6435 (N_6435,N_6248,N_6277);
or U6436 (N_6436,N_6282,N_6363);
and U6437 (N_6437,N_6358,N_6392);
xnor U6438 (N_6438,N_6327,N_6333);
nand U6439 (N_6439,N_6315,N_6295);
nor U6440 (N_6440,N_6376,N_6289);
or U6441 (N_6441,N_6394,N_6280);
xor U6442 (N_6442,N_6257,N_6326);
xnor U6443 (N_6443,N_6322,N_6382);
or U6444 (N_6444,N_6269,N_6260);
nand U6445 (N_6445,N_6249,N_6346);
and U6446 (N_6446,N_6272,N_6290);
or U6447 (N_6447,N_6251,N_6308);
xor U6448 (N_6448,N_6317,N_6351);
or U6449 (N_6449,N_6396,N_6301);
nand U6450 (N_6450,N_6292,N_6397);
xor U6451 (N_6451,N_6352,N_6309);
nand U6452 (N_6452,N_6273,N_6364);
xor U6453 (N_6453,N_6265,N_6385);
nor U6454 (N_6454,N_6305,N_6242);
nand U6455 (N_6455,N_6318,N_6328);
nor U6456 (N_6456,N_6342,N_6247);
nor U6457 (N_6457,N_6316,N_6334);
xor U6458 (N_6458,N_6274,N_6372);
and U6459 (N_6459,N_6304,N_6240);
nor U6460 (N_6460,N_6349,N_6303);
xnor U6461 (N_6461,N_6379,N_6271);
or U6462 (N_6462,N_6288,N_6359);
and U6463 (N_6463,N_6258,N_6312);
xor U6464 (N_6464,N_6354,N_6241);
nand U6465 (N_6465,N_6314,N_6294);
nor U6466 (N_6466,N_6299,N_6311);
and U6467 (N_6467,N_6283,N_6353);
nor U6468 (N_6468,N_6287,N_6388);
or U6469 (N_6469,N_6332,N_6243);
or U6470 (N_6470,N_6398,N_6393);
xnor U6471 (N_6471,N_6262,N_6344);
xnor U6472 (N_6472,N_6357,N_6263);
or U6473 (N_6473,N_6279,N_6386);
or U6474 (N_6474,N_6252,N_6335);
nor U6475 (N_6475,N_6373,N_6378);
nor U6476 (N_6476,N_6374,N_6281);
xor U6477 (N_6477,N_6380,N_6365);
or U6478 (N_6478,N_6336,N_6324);
or U6479 (N_6479,N_6345,N_6244);
or U6480 (N_6480,N_6387,N_6376);
and U6481 (N_6481,N_6385,N_6342);
xor U6482 (N_6482,N_6356,N_6288);
xor U6483 (N_6483,N_6318,N_6316);
xnor U6484 (N_6484,N_6288,N_6321);
xnor U6485 (N_6485,N_6244,N_6293);
nand U6486 (N_6486,N_6399,N_6380);
xnor U6487 (N_6487,N_6247,N_6257);
and U6488 (N_6488,N_6319,N_6393);
nor U6489 (N_6489,N_6268,N_6245);
nor U6490 (N_6490,N_6300,N_6383);
nand U6491 (N_6491,N_6258,N_6337);
or U6492 (N_6492,N_6383,N_6289);
nor U6493 (N_6493,N_6295,N_6304);
nand U6494 (N_6494,N_6293,N_6308);
and U6495 (N_6495,N_6389,N_6352);
nand U6496 (N_6496,N_6371,N_6308);
nor U6497 (N_6497,N_6321,N_6261);
or U6498 (N_6498,N_6251,N_6286);
nor U6499 (N_6499,N_6285,N_6303);
and U6500 (N_6500,N_6390,N_6351);
xnor U6501 (N_6501,N_6246,N_6308);
nor U6502 (N_6502,N_6325,N_6386);
or U6503 (N_6503,N_6300,N_6389);
or U6504 (N_6504,N_6276,N_6251);
and U6505 (N_6505,N_6350,N_6291);
and U6506 (N_6506,N_6300,N_6345);
xnor U6507 (N_6507,N_6279,N_6311);
nand U6508 (N_6508,N_6295,N_6314);
xnor U6509 (N_6509,N_6267,N_6359);
or U6510 (N_6510,N_6286,N_6276);
and U6511 (N_6511,N_6285,N_6332);
xor U6512 (N_6512,N_6334,N_6357);
or U6513 (N_6513,N_6370,N_6329);
nand U6514 (N_6514,N_6324,N_6264);
nor U6515 (N_6515,N_6249,N_6303);
nor U6516 (N_6516,N_6349,N_6383);
nor U6517 (N_6517,N_6245,N_6394);
xor U6518 (N_6518,N_6318,N_6390);
and U6519 (N_6519,N_6346,N_6335);
or U6520 (N_6520,N_6299,N_6293);
nor U6521 (N_6521,N_6251,N_6304);
xor U6522 (N_6522,N_6353,N_6297);
and U6523 (N_6523,N_6345,N_6333);
nand U6524 (N_6524,N_6387,N_6368);
nor U6525 (N_6525,N_6397,N_6374);
xnor U6526 (N_6526,N_6299,N_6351);
xor U6527 (N_6527,N_6265,N_6280);
and U6528 (N_6528,N_6283,N_6332);
nor U6529 (N_6529,N_6303,N_6244);
xor U6530 (N_6530,N_6383,N_6282);
nor U6531 (N_6531,N_6278,N_6341);
nor U6532 (N_6532,N_6334,N_6363);
nor U6533 (N_6533,N_6298,N_6352);
and U6534 (N_6534,N_6321,N_6339);
xor U6535 (N_6535,N_6299,N_6268);
or U6536 (N_6536,N_6275,N_6354);
xnor U6537 (N_6537,N_6283,N_6342);
nand U6538 (N_6538,N_6269,N_6362);
nor U6539 (N_6539,N_6276,N_6299);
or U6540 (N_6540,N_6398,N_6255);
xor U6541 (N_6541,N_6369,N_6269);
nor U6542 (N_6542,N_6275,N_6251);
xnor U6543 (N_6543,N_6297,N_6335);
nand U6544 (N_6544,N_6284,N_6265);
or U6545 (N_6545,N_6285,N_6329);
xnor U6546 (N_6546,N_6354,N_6287);
xnor U6547 (N_6547,N_6255,N_6358);
nand U6548 (N_6548,N_6350,N_6296);
nand U6549 (N_6549,N_6390,N_6262);
nor U6550 (N_6550,N_6396,N_6299);
nor U6551 (N_6551,N_6347,N_6367);
xor U6552 (N_6552,N_6382,N_6303);
nor U6553 (N_6553,N_6376,N_6276);
or U6554 (N_6554,N_6285,N_6242);
or U6555 (N_6555,N_6380,N_6393);
xor U6556 (N_6556,N_6314,N_6389);
nor U6557 (N_6557,N_6358,N_6259);
and U6558 (N_6558,N_6264,N_6244);
nand U6559 (N_6559,N_6242,N_6322);
nand U6560 (N_6560,N_6476,N_6546);
nor U6561 (N_6561,N_6435,N_6436);
nor U6562 (N_6562,N_6517,N_6420);
nor U6563 (N_6563,N_6479,N_6441);
or U6564 (N_6564,N_6478,N_6445);
nor U6565 (N_6565,N_6432,N_6493);
and U6566 (N_6566,N_6498,N_6450);
nor U6567 (N_6567,N_6511,N_6469);
nand U6568 (N_6568,N_6447,N_6508);
and U6569 (N_6569,N_6426,N_6497);
nand U6570 (N_6570,N_6408,N_6439);
or U6571 (N_6571,N_6440,N_6530);
or U6572 (N_6572,N_6434,N_6475);
or U6573 (N_6573,N_6552,N_6416);
xor U6574 (N_6574,N_6405,N_6422);
or U6575 (N_6575,N_6502,N_6461);
nand U6576 (N_6576,N_6510,N_6543);
or U6577 (N_6577,N_6526,N_6443);
nand U6578 (N_6578,N_6438,N_6427);
nor U6579 (N_6579,N_6402,N_6407);
or U6580 (N_6580,N_6471,N_6509);
or U6581 (N_6581,N_6548,N_6406);
and U6582 (N_6582,N_6522,N_6444);
nand U6583 (N_6583,N_6520,N_6462);
nor U6584 (N_6584,N_6554,N_6477);
and U6585 (N_6585,N_6431,N_6538);
or U6586 (N_6586,N_6413,N_6531);
and U6587 (N_6587,N_6480,N_6521);
nand U6588 (N_6588,N_6536,N_6425);
nor U6589 (N_6589,N_6421,N_6401);
nor U6590 (N_6590,N_6513,N_6418);
and U6591 (N_6591,N_6448,N_6412);
nand U6592 (N_6592,N_6458,N_6472);
or U6593 (N_6593,N_6430,N_6446);
nor U6594 (N_6594,N_6500,N_6454);
nor U6595 (N_6595,N_6488,N_6400);
xor U6596 (N_6596,N_6417,N_6542);
and U6597 (N_6597,N_6501,N_6491);
xnor U6598 (N_6598,N_6483,N_6468);
nor U6599 (N_6599,N_6528,N_6499);
xor U6600 (N_6600,N_6541,N_6525);
nor U6601 (N_6601,N_6534,N_6544);
or U6602 (N_6602,N_6424,N_6423);
or U6603 (N_6603,N_6545,N_6505);
xnor U6604 (N_6604,N_6455,N_6464);
and U6605 (N_6605,N_6555,N_6467);
xor U6606 (N_6606,N_6539,N_6492);
and U6607 (N_6607,N_6519,N_6459);
nand U6608 (N_6608,N_6465,N_6512);
and U6609 (N_6609,N_6527,N_6460);
or U6610 (N_6610,N_6414,N_6504);
nor U6611 (N_6611,N_6533,N_6456);
nor U6612 (N_6612,N_6419,N_6540);
nor U6613 (N_6613,N_6518,N_6486);
and U6614 (N_6614,N_6466,N_6474);
and U6615 (N_6615,N_6433,N_6556);
or U6616 (N_6616,N_6549,N_6410);
or U6617 (N_6617,N_6496,N_6484);
and U6618 (N_6618,N_6551,N_6449);
or U6619 (N_6619,N_6489,N_6482);
nand U6620 (N_6620,N_6494,N_6457);
nand U6621 (N_6621,N_6437,N_6428);
or U6622 (N_6622,N_6524,N_6550);
nand U6623 (N_6623,N_6559,N_6470);
xor U6624 (N_6624,N_6490,N_6403);
or U6625 (N_6625,N_6503,N_6507);
or U6626 (N_6626,N_6529,N_6463);
or U6627 (N_6627,N_6453,N_6523);
and U6628 (N_6628,N_6481,N_6558);
nor U6629 (N_6629,N_6404,N_6514);
nand U6630 (N_6630,N_6409,N_6487);
xnor U6631 (N_6631,N_6506,N_6411);
nor U6632 (N_6632,N_6473,N_6515);
and U6633 (N_6633,N_6485,N_6415);
nand U6634 (N_6634,N_6495,N_6537);
xor U6635 (N_6635,N_6452,N_6516);
nand U6636 (N_6636,N_6429,N_6553);
and U6637 (N_6637,N_6547,N_6557);
nor U6638 (N_6638,N_6535,N_6532);
nor U6639 (N_6639,N_6442,N_6451);
or U6640 (N_6640,N_6523,N_6541);
nor U6641 (N_6641,N_6502,N_6428);
or U6642 (N_6642,N_6455,N_6533);
or U6643 (N_6643,N_6401,N_6433);
and U6644 (N_6644,N_6544,N_6418);
nand U6645 (N_6645,N_6404,N_6513);
nand U6646 (N_6646,N_6404,N_6525);
xnor U6647 (N_6647,N_6549,N_6461);
xor U6648 (N_6648,N_6516,N_6427);
nor U6649 (N_6649,N_6442,N_6504);
and U6650 (N_6650,N_6413,N_6400);
nand U6651 (N_6651,N_6533,N_6450);
xor U6652 (N_6652,N_6547,N_6490);
xor U6653 (N_6653,N_6553,N_6539);
nor U6654 (N_6654,N_6529,N_6490);
and U6655 (N_6655,N_6403,N_6510);
or U6656 (N_6656,N_6417,N_6411);
xnor U6657 (N_6657,N_6552,N_6435);
and U6658 (N_6658,N_6522,N_6451);
and U6659 (N_6659,N_6525,N_6400);
nor U6660 (N_6660,N_6513,N_6500);
nor U6661 (N_6661,N_6504,N_6412);
xnor U6662 (N_6662,N_6518,N_6462);
or U6663 (N_6663,N_6545,N_6537);
and U6664 (N_6664,N_6462,N_6491);
nor U6665 (N_6665,N_6502,N_6514);
nor U6666 (N_6666,N_6495,N_6477);
nand U6667 (N_6667,N_6540,N_6550);
or U6668 (N_6668,N_6530,N_6479);
or U6669 (N_6669,N_6429,N_6515);
xnor U6670 (N_6670,N_6524,N_6423);
nor U6671 (N_6671,N_6431,N_6441);
nand U6672 (N_6672,N_6442,N_6465);
nand U6673 (N_6673,N_6497,N_6550);
and U6674 (N_6674,N_6554,N_6525);
nor U6675 (N_6675,N_6432,N_6499);
nor U6676 (N_6676,N_6520,N_6460);
xnor U6677 (N_6677,N_6496,N_6456);
nor U6678 (N_6678,N_6548,N_6442);
and U6679 (N_6679,N_6466,N_6453);
or U6680 (N_6680,N_6459,N_6551);
nand U6681 (N_6681,N_6521,N_6461);
xor U6682 (N_6682,N_6441,N_6541);
and U6683 (N_6683,N_6410,N_6420);
nor U6684 (N_6684,N_6402,N_6454);
nand U6685 (N_6685,N_6545,N_6425);
xnor U6686 (N_6686,N_6516,N_6458);
nand U6687 (N_6687,N_6549,N_6523);
or U6688 (N_6688,N_6500,N_6504);
nor U6689 (N_6689,N_6506,N_6412);
nor U6690 (N_6690,N_6517,N_6408);
nand U6691 (N_6691,N_6418,N_6440);
and U6692 (N_6692,N_6489,N_6417);
or U6693 (N_6693,N_6520,N_6505);
xnor U6694 (N_6694,N_6496,N_6477);
or U6695 (N_6695,N_6553,N_6400);
nor U6696 (N_6696,N_6524,N_6402);
nand U6697 (N_6697,N_6410,N_6423);
nor U6698 (N_6698,N_6403,N_6541);
nor U6699 (N_6699,N_6499,N_6521);
nor U6700 (N_6700,N_6444,N_6532);
xnor U6701 (N_6701,N_6553,N_6436);
or U6702 (N_6702,N_6516,N_6536);
and U6703 (N_6703,N_6428,N_6429);
and U6704 (N_6704,N_6519,N_6486);
nor U6705 (N_6705,N_6496,N_6409);
and U6706 (N_6706,N_6471,N_6547);
nand U6707 (N_6707,N_6481,N_6535);
xor U6708 (N_6708,N_6459,N_6523);
and U6709 (N_6709,N_6536,N_6523);
or U6710 (N_6710,N_6509,N_6531);
and U6711 (N_6711,N_6502,N_6414);
nand U6712 (N_6712,N_6441,N_6409);
nor U6713 (N_6713,N_6461,N_6453);
xnor U6714 (N_6714,N_6522,N_6427);
xnor U6715 (N_6715,N_6456,N_6457);
xnor U6716 (N_6716,N_6489,N_6512);
or U6717 (N_6717,N_6420,N_6484);
xor U6718 (N_6718,N_6524,N_6466);
xnor U6719 (N_6719,N_6489,N_6538);
and U6720 (N_6720,N_6575,N_6648);
or U6721 (N_6721,N_6593,N_6675);
xnor U6722 (N_6722,N_6695,N_6677);
and U6723 (N_6723,N_6701,N_6646);
and U6724 (N_6724,N_6706,N_6687);
nand U6725 (N_6725,N_6622,N_6641);
xor U6726 (N_6726,N_6716,N_6608);
xor U6727 (N_6727,N_6634,N_6659);
xnor U6728 (N_6728,N_6671,N_6614);
and U6729 (N_6729,N_6697,N_6637);
nor U6730 (N_6730,N_6649,N_6655);
xor U6731 (N_6731,N_6615,N_6632);
and U6732 (N_6732,N_6696,N_6678);
or U6733 (N_6733,N_6656,N_6621);
nand U6734 (N_6734,N_6606,N_6709);
or U6735 (N_6735,N_6564,N_6693);
xor U6736 (N_6736,N_6662,N_6581);
nor U6737 (N_6737,N_6660,N_6570);
and U6738 (N_6738,N_6638,N_6616);
nor U6739 (N_6739,N_6610,N_6674);
nor U6740 (N_6740,N_6651,N_6639);
xnor U6741 (N_6741,N_6580,N_6684);
or U6742 (N_6742,N_6718,N_6635);
nor U6743 (N_6743,N_6563,N_6604);
nor U6744 (N_6744,N_6661,N_6682);
nand U6745 (N_6745,N_6699,N_6653);
xor U6746 (N_6746,N_6607,N_6681);
nor U6747 (N_6747,N_6618,N_6667);
or U6748 (N_6748,N_6663,N_6573);
and U6749 (N_6749,N_6600,N_6700);
and U6750 (N_6750,N_6691,N_6599);
nand U6751 (N_6751,N_6692,N_6715);
or U6752 (N_6752,N_6710,N_6589);
xor U6753 (N_6753,N_6586,N_6628);
xor U6754 (N_6754,N_6666,N_6576);
xor U6755 (N_6755,N_6711,N_6670);
nand U6756 (N_6756,N_6668,N_6623);
nor U6757 (N_6757,N_6567,N_6679);
xor U6758 (N_6758,N_6609,N_6590);
and U6759 (N_6759,N_6703,N_6571);
and U6760 (N_6760,N_6626,N_6582);
xnor U6761 (N_6761,N_6717,N_6713);
or U6762 (N_6762,N_6657,N_6603);
nor U6763 (N_6763,N_6591,N_6688);
nand U6764 (N_6764,N_6652,N_6644);
or U6765 (N_6765,N_6636,N_6605);
and U6766 (N_6766,N_6630,N_6704);
nor U6767 (N_6767,N_6572,N_6598);
nand U6768 (N_6768,N_6627,N_6676);
and U6769 (N_6769,N_6579,N_6642);
or U6770 (N_6770,N_6633,N_6650);
and U6771 (N_6771,N_6617,N_6707);
nor U6772 (N_6772,N_6566,N_6624);
nor U6773 (N_6773,N_6584,N_6645);
xnor U6774 (N_6774,N_6665,N_6654);
nor U6775 (N_6775,N_6583,N_6698);
nor U6776 (N_6776,N_6585,N_6664);
xnor U6777 (N_6777,N_6647,N_6562);
nand U6778 (N_6778,N_6561,N_6694);
and U6779 (N_6779,N_6613,N_6560);
nand U6780 (N_6780,N_6574,N_6611);
nand U6781 (N_6781,N_6568,N_6620);
nand U6782 (N_6782,N_6669,N_6702);
nor U6783 (N_6783,N_6629,N_6683);
and U6784 (N_6784,N_6592,N_6673);
nor U6785 (N_6785,N_6708,N_6643);
nand U6786 (N_6786,N_6625,N_6640);
nand U6787 (N_6787,N_6631,N_6587);
xnor U6788 (N_6788,N_6612,N_6578);
nor U6789 (N_6789,N_6658,N_6595);
or U6790 (N_6790,N_6719,N_6712);
nand U6791 (N_6791,N_6619,N_6601);
or U6792 (N_6792,N_6686,N_6602);
and U6793 (N_6793,N_6597,N_6588);
nand U6794 (N_6794,N_6672,N_6685);
nand U6795 (N_6795,N_6569,N_6577);
nand U6796 (N_6796,N_6714,N_6689);
or U6797 (N_6797,N_6680,N_6594);
or U6798 (N_6798,N_6565,N_6690);
xor U6799 (N_6799,N_6596,N_6705);
and U6800 (N_6800,N_6617,N_6597);
nand U6801 (N_6801,N_6701,N_6580);
nand U6802 (N_6802,N_6602,N_6641);
and U6803 (N_6803,N_6593,N_6648);
and U6804 (N_6804,N_6606,N_6632);
xor U6805 (N_6805,N_6645,N_6646);
and U6806 (N_6806,N_6643,N_6584);
or U6807 (N_6807,N_6625,N_6715);
or U6808 (N_6808,N_6572,N_6625);
xnor U6809 (N_6809,N_6624,N_6632);
xor U6810 (N_6810,N_6698,N_6612);
nor U6811 (N_6811,N_6651,N_6654);
or U6812 (N_6812,N_6709,N_6607);
nand U6813 (N_6813,N_6628,N_6574);
and U6814 (N_6814,N_6704,N_6628);
xor U6815 (N_6815,N_6642,N_6633);
and U6816 (N_6816,N_6638,N_6691);
or U6817 (N_6817,N_6587,N_6695);
nand U6818 (N_6818,N_6561,N_6577);
nor U6819 (N_6819,N_6607,N_6574);
nor U6820 (N_6820,N_6715,N_6681);
and U6821 (N_6821,N_6703,N_6676);
xor U6822 (N_6822,N_6651,N_6667);
xor U6823 (N_6823,N_6713,N_6695);
nor U6824 (N_6824,N_6677,N_6674);
nand U6825 (N_6825,N_6695,N_6631);
xnor U6826 (N_6826,N_6702,N_6714);
and U6827 (N_6827,N_6688,N_6685);
or U6828 (N_6828,N_6659,N_6695);
nor U6829 (N_6829,N_6645,N_6575);
or U6830 (N_6830,N_6635,N_6591);
xnor U6831 (N_6831,N_6632,N_6576);
and U6832 (N_6832,N_6587,N_6690);
nand U6833 (N_6833,N_6659,N_6617);
or U6834 (N_6834,N_6577,N_6679);
nand U6835 (N_6835,N_6656,N_6617);
or U6836 (N_6836,N_6655,N_6587);
or U6837 (N_6837,N_6710,N_6717);
nor U6838 (N_6838,N_6663,N_6703);
and U6839 (N_6839,N_6585,N_6615);
nor U6840 (N_6840,N_6595,N_6669);
nor U6841 (N_6841,N_6716,N_6642);
or U6842 (N_6842,N_6644,N_6565);
and U6843 (N_6843,N_6638,N_6636);
nor U6844 (N_6844,N_6695,N_6706);
or U6845 (N_6845,N_6629,N_6587);
nor U6846 (N_6846,N_6701,N_6641);
xor U6847 (N_6847,N_6627,N_6695);
nand U6848 (N_6848,N_6719,N_6711);
or U6849 (N_6849,N_6679,N_6568);
or U6850 (N_6850,N_6565,N_6632);
and U6851 (N_6851,N_6668,N_6652);
or U6852 (N_6852,N_6570,N_6643);
nand U6853 (N_6853,N_6657,N_6560);
xnor U6854 (N_6854,N_6567,N_6675);
nand U6855 (N_6855,N_6672,N_6682);
or U6856 (N_6856,N_6576,N_6661);
nor U6857 (N_6857,N_6563,N_6588);
xnor U6858 (N_6858,N_6693,N_6702);
xor U6859 (N_6859,N_6607,N_6658);
and U6860 (N_6860,N_6665,N_6588);
or U6861 (N_6861,N_6716,N_6700);
nand U6862 (N_6862,N_6622,N_6662);
xnor U6863 (N_6863,N_6664,N_6595);
and U6864 (N_6864,N_6596,N_6709);
and U6865 (N_6865,N_6665,N_6585);
or U6866 (N_6866,N_6562,N_6682);
xor U6867 (N_6867,N_6596,N_6617);
nor U6868 (N_6868,N_6713,N_6618);
nand U6869 (N_6869,N_6600,N_6583);
xor U6870 (N_6870,N_6658,N_6561);
or U6871 (N_6871,N_6655,N_6697);
nand U6872 (N_6872,N_6640,N_6648);
or U6873 (N_6873,N_6688,N_6619);
nor U6874 (N_6874,N_6712,N_6564);
or U6875 (N_6875,N_6667,N_6680);
xnor U6876 (N_6876,N_6642,N_6617);
nor U6877 (N_6877,N_6683,N_6666);
or U6878 (N_6878,N_6560,N_6716);
or U6879 (N_6879,N_6712,N_6633);
nand U6880 (N_6880,N_6786,N_6772);
and U6881 (N_6881,N_6744,N_6859);
xor U6882 (N_6882,N_6759,N_6766);
nor U6883 (N_6883,N_6858,N_6720);
nand U6884 (N_6884,N_6737,N_6855);
nor U6885 (N_6885,N_6745,N_6808);
nand U6886 (N_6886,N_6799,N_6877);
nor U6887 (N_6887,N_6754,N_6760);
and U6888 (N_6888,N_6804,N_6724);
xor U6889 (N_6889,N_6853,N_6820);
or U6890 (N_6890,N_6733,N_6755);
or U6891 (N_6891,N_6729,N_6735);
nor U6892 (N_6892,N_6844,N_6774);
xor U6893 (N_6893,N_6838,N_6812);
xnor U6894 (N_6894,N_6725,N_6753);
and U6895 (N_6895,N_6782,N_6834);
xnor U6896 (N_6896,N_6768,N_6835);
or U6897 (N_6897,N_6852,N_6878);
nor U6898 (N_6898,N_6762,N_6815);
nand U6899 (N_6899,N_6831,N_6795);
xnor U6900 (N_6900,N_6829,N_6765);
or U6901 (N_6901,N_6867,N_6806);
or U6902 (N_6902,N_6865,N_6741);
or U6903 (N_6903,N_6814,N_6781);
and U6904 (N_6904,N_6739,N_6784);
xor U6905 (N_6905,N_6860,N_6872);
nand U6906 (N_6906,N_6749,N_6803);
nand U6907 (N_6907,N_6863,N_6792);
xor U6908 (N_6908,N_6790,N_6746);
nor U6909 (N_6909,N_6726,N_6805);
nor U6910 (N_6910,N_6779,N_6847);
xor U6911 (N_6911,N_6777,N_6848);
and U6912 (N_6912,N_6798,N_6824);
xor U6913 (N_6913,N_6827,N_6832);
or U6914 (N_6914,N_6787,N_6742);
nand U6915 (N_6915,N_6730,N_6828);
xor U6916 (N_6916,N_6861,N_6841);
xnor U6917 (N_6917,N_6833,N_6796);
xor U6918 (N_6918,N_6722,N_6721);
nor U6919 (N_6919,N_6748,N_6738);
xor U6920 (N_6920,N_6870,N_6761);
xnor U6921 (N_6921,N_6727,N_6869);
xor U6922 (N_6922,N_6871,N_6846);
and U6923 (N_6923,N_6797,N_6840);
nor U6924 (N_6924,N_6757,N_6843);
nand U6925 (N_6925,N_6773,N_6758);
or U6926 (N_6926,N_6818,N_6771);
nand U6927 (N_6927,N_6750,N_6822);
or U6928 (N_6928,N_6817,N_6837);
xnor U6929 (N_6929,N_6868,N_6788);
or U6930 (N_6930,N_6874,N_6816);
nor U6931 (N_6931,N_6876,N_6845);
or U6932 (N_6932,N_6791,N_6810);
xnor U6933 (N_6933,N_6794,N_6747);
or U6934 (N_6934,N_6836,N_6740);
and U6935 (N_6935,N_6851,N_6785);
nand U6936 (N_6936,N_6780,N_6778);
xor U6937 (N_6937,N_6775,N_6821);
xnor U6938 (N_6938,N_6728,N_6864);
or U6939 (N_6939,N_6875,N_6830);
xnor U6940 (N_6940,N_6825,N_6763);
nor U6941 (N_6941,N_6732,N_6857);
nand U6942 (N_6942,N_6734,N_6769);
nand U6943 (N_6943,N_6879,N_6862);
xor U6944 (N_6944,N_6743,N_6826);
xnor U6945 (N_6945,N_6823,N_6801);
xnor U6946 (N_6946,N_6811,N_6849);
nor U6947 (N_6947,N_6767,N_6856);
nor U6948 (N_6948,N_6723,N_6839);
xnor U6949 (N_6949,N_6854,N_6800);
nand U6950 (N_6950,N_6866,N_6731);
nand U6951 (N_6951,N_6873,N_6793);
xnor U6952 (N_6952,N_6850,N_6752);
nor U6953 (N_6953,N_6813,N_6776);
xor U6954 (N_6954,N_6783,N_6751);
and U6955 (N_6955,N_6802,N_6756);
and U6956 (N_6956,N_6789,N_6842);
xnor U6957 (N_6957,N_6819,N_6807);
and U6958 (N_6958,N_6764,N_6809);
xnor U6959 (N_6959,N_6770,N_6736);
or U6960 (N_6960,N_6722,N_6756);
nand U6961 (N_6961,N_6740,N_6805);
nand U6962 (N_6962,N_6742,N_6740);
nor U6963 (N_6963,N_6766,N_6727);
xor U6964 (N_6964,N_6724,N_6732);
or U6965 (N_6965,N_6787,N_6839);
nor U6966 (N_6966,N_6864,N_6759);
xnor U6967 (N_6967,N_6727,N_6872);
xnor U6968 (N_6968,N_6808,N_6854);
or U6969 (N_6969,N_6830,N_6821);
or U6970 (N_6970,N_6877,N_6864);
xor U6971 (N_6971,N_6793,N_6841);
and U6972 (N_6972,N_6783,N_6871);
or U6973 (N_6973,N_6751,N_6835);
or U6974 (N_6974,N_6864,N_6841);
nor U6975 (N_6975,N_6788,N_6879);
nor U6976 (N_6976,N_6858,N_6782);
or U6977 (N_6977,N_6872,N_6745);
and U6978 (N_6978,N_6772,N_6842);
nor U6979 (N_6979,N_6846,N_6842);
xor U6980 (N_6980,N_6763,N_6793);
nand U6981 (N_6981,N_6733,N_6791);
nand U6982 (N_6982,N_6814,N_6827);
nand U6983 (N_6983,N_6851,N_6793);
and U6984 (N_6984,N_6777,N_6806);
xnor U6985 (N_6985,N_6800,N_6723);
nor U6986 (N_6986,N_6775,N_6741);
nand U6987 (N_6987,N_6724,N_6801);
or U6988 (N_6988,N_6732,N_6832);
nand U6989 (N_6989,N_6879,N_6878);
xnor U6990 (N_6990,N_6820,N_6876);
or U6991 (N_6991,N_6803,N_6826);
nand U6992 (N_6992,N_6867,N_6752);
nand U6993 (N_6993,N_6817,N_6839);
or U6994 (N_6994,N_6854,N_6738);
xor U6995 (N_6995,N_6832,N_6745);
xnor U6996 (N_6996,N_6802,N_6813);
nand U6997 (N_6997,N_6731,N_6824);
and U6998 (N_6998,N_6734,N_6853);
nand U6999 (N_6999,N_6867,N_6799);
nand U7000 (N_7000,N_6835,N_6867);
xor U7001 (N_7001,N_6727,N_6832);
xnor U7002 (N_7002,N_6801,N_6857);
nand U7003 (N_7003,N_6800,N_6855);
xnor U7004 (N_7004,N_6817,N_6768);
nand U7005 (N_7005,N_6813,N_6781);
xor U7006 (N_7006,N_6822,N_6785);
nor U7007 (N_7007,N_6858,N_6851);
nor U7008 (N_7008,N_6845,N_6801);
and U7009 (N_7009,N_6759,N_6746);
nand U7010 (N_7010,N_6751,N_6840);
nor U7011 (N_7011,N_6757,N_6839);
xnor U7012 (N_7012,N_6728,N_6815);
or U7013 (N_7013,N_6740,N_6842);
and U7014 (N_7014,N_6728,N_6788);
nor U7015 (N_7015,N_6762,N_6827);
xor U7016 (N_7016,N_6791,N_6780);
xnor U7017 (N_7017,N_6871,N_6863);
and U7018 (N_7018,N_6735,N_6797);
and U7019 (N_7019,N_6756,N_6867);
xor U7020 (N_7020,N_6857,N_6848);
xnor U7021 (N_7021,N_6873,N_6868);
nor U7022 (N_7022,N_6781,N_6735);
and U7023 (N_7023,N_6860,N_6762);
nor U7024 (N_7024,N_6783,N_6818);
or U7025 (N_7025,N_6776,N_6732);
xor U7026 (N_7026,N_6862,N_6759);
nand U7027 (N_7027,N_6756,N_6845);
xor U7028 (N_7028,N_6721,N_6731);
xnor U7029 (N_7029,N_6771,N_6859);
and U7030 (N_7030,N_6864,N_6762);
or U7031 (N_7031,N_6725,N_6867);
xnor U7032 (N_7032,N_6831,N_6871);
or U7033 (N_7033,N_6850,N_6878);
xor U7034 (N_7034,N_6732,N_6767);
nor U7035 (N_7035,N_6756,N_6720);
and U7036 (N_7036,N_6871,N_6813);
nand U7037 (N_7037,N_6792,N_6783);
nor U7038 (N_7038,N_6774,N_6776);
nand U7039 (N_7039,N_6815,N_6817);
or U7040 (N_7040,N_6880,N_7036);
or U7041 (N_7041,N_6942,N_6975);
or U7042 (N_7042,N_6992,N_6967);
nand U7043 (N_7043,N_7037,N_6987);
and U7044 (N_7044,N_7016,N_7020);
nor U7045 (N_7045,N_6928,N_6890);
and U7046 (N_7046,N_7003,N_7025);
xor U7047 (N_7047,N_6905,N_7012);
xor U7048 (N_7048,N_7023,N_7008);
and U7049 (N_7049,N_6956,N_7035);
and U7050 (N_7050,N_6965,N_7029);
nor U7051 (N_7051,N_6953,N_6952);
nor U7052 (N_7052,N_7005,N_6969);
nor U7053 (N_7053,N_6909,N_7006);
xnor U7054 (N_7054,N_6897,N_7024);
nand U7055 (N_7055,N_6936,N_6949);
xnor U7056 (N_7056,N_6892,N_7002);
xnor U7057 (N_7057,N_6925,N_6889);
xor U7058 (N_7058,N_7030,N_6973);
nor U7059 (N_7059,N_7000,N_6908);
nor U7060 (N_7060,N_7022,N_6903);
nor U7061 (N_7061,N_6955,N_6923);
or U7062 (N_7062,N_6950,N_6886);
nand U7063 (N_7063,N_6896,N_6900);
nor U7064 (N_7064,N_7028,N_6982);
and U7065 (N_7065,N_6996,N_6984);
or U7066 (N_7066,N_6995,N_7019);
nand U7067 (N_7067,N_7031,N_6977);
xnor U7068 (N_7068,N_6957,N_6913);
xnor U7069 (N_7069,N_6948,N_7034);
nor U7070 (N_7070,N_6986,N_7014);
nor U7071 (N_7071,N_6993,N_7004);
and U7072 (N_7072,N_7021,N_6976);
or U7073 (N_7073,N_6902,N_6914);
nor U7074 (N_7074,N_6971,N_6947);
nor U7075 (N_7075,N_7017,N_6893);
and U7076 (N_7076,N_6933,N_7009);
nor U7077 (N_7077,N_6916,N_6990);
xor U7078 (N_7078,N_6959,N_6911);
or U7079 (N_7079,N_7038,N_6962);
nand U7080 (N_7080,N_6921,N_6985);
or U7081 (N_7081,N_6887,N_6970);
or U7082 (N_7082,N_6968,N_6974);
or U7083 (N_7083,N_6932,N_6972);
or U7084 (N_7084,N_6898,N_6978);
nor U7085 (N_7085,N_6934,N_6960);
nor U7086 (N_7086,N_6951,N_6904);
nand U7087 (N_7087,N_6901,N_6991);
xor U7088 (N_7088,N_6888,N_6918);
nor U7089 (N_7089,N_6899,N_6927);
nand U7090 (N_7090,N_7015,N_6894);
xor U7091 (N_7091,N_6958,N_6883);
xor U7092 (N_7092,N_6907,N_6961);
or U7093 (N_7093,N_7010,N_7039);
and U7094 (N_7094,N_6912,N_6944);
xor U7095 (N_7095,N_6989,N_6924);
xor U7096 (N_7096,N_6998,N_7032);
or U7097 (N_7097,N_6938,N_6915);
nor U7098 (N_7098,N_6885,N_6963);
or U7099 (N_7099,N_6997,N_6964);
nor U7100 (N_7100,N_6999,N_6920);
and U7101 (N_7101,N_6943,N_6930);
or U7102 (N_7102,N_6966,N_6954);
and U7103 (N_7103,N_6917,N_6906);
nand U7104 (N_7104,N_6929,N_6895);
nor U7105 (N_7105,N_6937,N_7033);
xnor U7106 (N_7106,N_7001,N_6983);
xnor U7107 (N_7107,N_6994,N_6882);
nand U7108 (N_7108,N_6926,N_6941);
nand U7109 (N_7109,N_7026,N_7007);
and U7110 (N_7110,N_6910,N_6919);
or U7111 (N_7111,N_6945,N_6981);
nand U7112 (N_7112,N_7018,N_6946);
nand U7113 (N_7113,N_6988,N_6979);
xnor U7114 (N_7114,N_7011,N_6884);
xor U7115 (N_7115,N_7013,N_6980);
nand U7116 (N_7116,N_6935,N_6922);
or U7117 (N_7117,N_6891,N_6940);
xnor U7118 (N_7118,N_6881,N_6931);
and U7119 (N_7119,N_7027,N_6939);
xnor U7120 (N_7120,N_6915,N_6909);
nand U7121 (N_7121,N_6980,N_6953);
xor U7122 (N_7122,N_6905,N_6897);
nand U7123 (N_7123,N_6929,N_6896);
or U7124 (N_7124,N_7019,N_6925);
nand U7125 (N_7125,N_6956,N_6906);
xnor U7126 (N_7126,N_6991,N_6952);
nor U7127 (N_7127,N_6993,N_7009);
nand U7128 (N_7128,N_6900,N_7015);
or U7129 (N_7129,N_6944,N_7009);
or U7130 (N_7130,N_6925,N_6946);
xor U7131 (N_7131,N_7018,N_6890);
nand U7132 (N_7132,N_6909,N_6920);
xor U7133 (N_7133,N_6969,N_6982);
xor U7134 (N_7134,N_6895,N_6881);
or U7135 (N_7135,N_6916,N_6887);
xor U7136 (N_7136,N_7029,N_6964);
xnor U7137 (N_7137,N_6887,N_6898);
nor U7138 (N_7138,N_6943,N_6999);
or U7139 (N_7139,N_6936,N_6932);
xnor U7140 (N_7140,N_6976,N_6961);
or U7141 (N_7141,N_7002,N_7011);
xnor U7142 (N_7142,N_6929,N_6954);
xnor U7143 (N_7143,N_7017,N_6981);
nand U7144 (N_7144,N_7014,N_6896);
xor U7145 (N_7145,N_6965,N_6995);
nor U7146 (N_7146,N_7038,N_6926);
nand U7147 (N_7147,N_6946,N_6972);
xor U7148 (N_7148,N_7014,N_6898);
xor U7149 (N_7149,N_6912,N_6993);
or U7150 (N_7150,N_6976,N_6918);
or U7151 (N_7151,N_6917,N_6965);
and U7152 (N_7152,N_7020,N_7022);
xor U7153 (N_7153,N_6913,N_6960);
or U7154 (N_7154,N_6932,N_7036);
or U7155 (N_7155,N_6935,N_7033);
or U7156 (N_7156,N_6922,N_6998);
nand U7157 (N_7157,N_6973,N_6991);
nand U7158 (N_7158,N_7014,N_6959);
nor U7159 (N_7159,N_7027,N_6926);
xor U7160 (N_7160,N_6918,N_6993);
and U7161 (N_7161,N_6952,N_6972);
and U7162 (N_7162,N_6892,N_6912);
and U7163 (N_7163,N_6904,N_7017);
and U7164 (N_7164,N_6921,N_6957);
nand U7165 (N_7165,N_7001,N_6939);
and U7166 (N_7166,N_6910,N_6898);
or U7167 (N_7167,N_6995,N_7021);
xnor U7168 (N_7168,N_7000,N_6942);
nor U7169 (N_7169,N_6981,N_7028);
nand U7170 (N_7170,N_6957,N_6917);
nor U7171 (N_7171,N_6895,N_7008);
and U7172 (N_7172,N_7005,N_6962);
nor U7173 (N_7173,N_7031,N_6909);
nand U7174 (N_7174,N_6922,N_6999);
xnor U7175 (N_7175,N_6927,N_6975);
or U7176 (N_7176,N_6933,N_7001);
nand U7177 (N_7177,N_6916,N_6926);
nor U7178 (N_7178,N_6907,N_6929);
nand U7179 (N_7179,N_6929,N_6988);
xor U7180 (N_7180,N_6906,N_6908);
and U7181 (N_7181,N_7037,N_6957);
nand U7182 (N_7182,N_6976,N_6912);
nand U7183 (N_7183,N_6983,N_7011);
nand U7184 (N_7184,N_6943,N_6948);
or U7185 (N_7185,N_6929,N_6985);
or U7186 (N_7186,N_6907,N_6916);
and U7187 (N_7187,N_6905,N_6919);
nor U7188 (N_7188,N_6987,N_7029);
nand U7189 (N_7189,N_6931,N_6900);
and U7190 (N_7190,N_6924,N_6985);
and U7191 (N_7191,N_7021,N_6901);
nand U7192 (N_7192,N_6973,N_6938);
nand U7193 (N_7193,N_7006,N_6882);
or U7194 (N_7194,N_6951,N_7034);
nor U7195 (N_7195,N_6955,N_6919);
and U7196 (N_7196,N_7035,N_6998);
nor U7197 (N_7197,N_7024,N_6990);
xnor U7198 (N_7198,N_6936,N_7009);
and U7199 (N_7199,N_6919,N_6911);
or U7200 (N_7200,N_7047,N_7117);
xor U7201 (N_7201,N_7150,N_7146);
or U7202 (N_7202,N_7085,N_7115);
and U7203 (N_7203,N_7070,N_7098);
and U7204 (N_7204,N_7162,N_7155);
xor U7205 (N_7205,N_7169,N_7105);
nor U7206 (N_7206,N_7195,N_7175);
and U7207 (N_7207,N_7109,N_7176);
and U7208 (N_7208,N_7174,N_7072);
nand U7209 (N_7209,N_7164,N_7188);
nor U7210 (N_7210,N_7140,N_7060);
nor U7211 (N_7211,N_7048,N_7066);
and U7212 (N_7212,N_7199,N_7193);
and U7213 (N_7213,N_7071,N_7139);
nor U7214 (N_7214,N_7108,N_7178);
and U7215 (N_7215,N_7165,N_7043);
nand U7216 (N_7216,N_7064,N_7143);
or U7217 (N_7217,N_7159,N_7076);
xnor U7218 (N_7218,N_7172,N_7045);
xor U7219 (N_7219,N_7086,N_7126);
or U7220 (N_7220,N_7197,N_7182);
nand U7221 (N_7221,N_7121,N_7107);
nor U7222 (N_7222,N_7183,N_7112);
nand U7223 (N_7223,N_7061,N_7106);
and U7224 (N_7224,N_7145,N_7099);
or U7225 (N_7225,N_7161,N_7113);
and U7226 (N_7226,N_7100,N_7144);
or U7227 (N_7227,N_7073,N_7111);
xor U7228 (N_7228,N_7180,N_7130);
xor U7229 (N_7229,N_7148,N_7138);
nand U7230 (N_7230,N_7095,N_7079);
and U7231 (N_7231,N_7080,N_7185);
nand U7232 (N_7232,N_7055,N_7198);
and U7233 (N_7233,N_7120,N_7181);
or U7234 (N_7234,N_7189,N_7094);
nor U7235 (N_7235,N_7135,N_7096);
or U7236 (N_7236,N_7054,N_7127);
or U7237 (N_7237,N_7184,N_7058);
xor U7238 (N_7238,N_7152,N_7104);
nor U7239 (N_7239,N_7186,N_7166);
nand U7240 (N_7240,N_7087,N_7053);
or U7241 (N_7241,N_7077,N_7062);
nand U7242 (N_7242,N_7083,N_7119);
nand U7243 (N_7243,N_7170,N_7133);
xnor U7244 (N_7244,N_7116,N_7049);
xnor U7245 (N_7245,N_7041,N_7173);
nor U7246 (N_7246,N_7131,N_7081);
nand U7247 (N_7247,N_7040,N_7067);
xor U7248 (N_7248,N_7046,N_7124);
nor U7249 (N_7249,N_7114,N_7153);
nand U7250 (N_7250,N_7160,N_7142);
and U7251 (N_7251,N_7134,N_7102);
xnor U7252 (N_7252,N_7158,N_7059);
and U7253 (N_7253,N_7074,N_7042);
or U7254 (N_7254,N_7190,N_7044);
and U7255 (N_7255,N_7163,N_7110);
xor U7256 (N_7256,N_7089,N_7123);
xnor U7257 (N_7257,N_7129,N_7101);
and U7258 (N_7258,N_7141,N_7052);
nor U7259 (N_7259,N_7191,N_7051);
or U7260 (N_7260,N_7118,N_7082);
and U7261 (N_7261,N_7154,N_7075);
xor U7262 (N_7262,N_7156,N_7068);
nor U7263 (N_7263,N_7147,N_7151);
nor U7264 (N_7264,N_7149,N_7157);
and U7265 (N_7265,N_7091,N_7065);
or U7266 (N_7266,N_7103,N_7137);
nor U7267 (N_7267,N_7093,N_7050);
nand U7268 (N_7268,N_7078,N_7125);
nor U7269 (N_7269,N_7084,N_7179);
nand U7270 (N_7270,N_7057,N_7171);
and U7271 (N_7271,N_7128,N_7168);
or U7272 (N_7272,N_7090,N_7187);
and U7273 (N_7273,N_7136,N_7063);
and U7274 (N_7274,N_7092,N_7097);
nor U7275 (N_7275,N_7196,N_7088);
nand U7276 (N_7276,N_7069,N_7177);
and U7277 (N_7277,N_7056,N_7122);
xnor U7278 (N_7278,N_7132,N_7167);
xnor U7279 (N_7279,N_7192,N_7194);
nor U7280 (N_7280,N_7150,N_7087);
xnor U7281 (N_7281,N_7123,N_7162);
or U7282 (N_7282,N_7131,N_7137);
xor U7283 (N_7283,N_7060,N_7182);
nor U7284 (N_7284,N_7180,N_7162);
and U7285 (N_7285,N_7050,N_7181);
nor U7286 (N_7286,N_7060,N_7105);
and U7287 (N_7287,N_7131,N_7152);
and U7288 (N_7288,N_7087,N_7184);
nor U7289 (N_7289,N_7092,N_7153);
nor U7290 (N_7290,N_7087,N_7156);
xnor U7291 (N_7291,N_7057,N_7086);
xor U7292 (N_7292,N_7173,N_7125);
or U7293 (N_7293,N_7185,N_7045);
xor U7294 (N_7294,N_7189,N_7092);
xor U7295 (N_7295,N_7171,N_7179);
and U7296 (N_7296,N_7153,N_7094);
nand U7297 (N_7297,N_7041,N_7116);
nand U7298 (N_7298,N_7128,N_7059);
or U7299 (N_7299,N_7190,N_7153);
and U7300 (N_7300,N_7042,N_7064);
or U7301 (N_7301,N_7050,N_7165);
and U7302 (N_7302,N_7177,N_7160);
nand U7303 (N_7303,N_7102,N_7071);
nand U7304 (N_7304,N_7161,N_7079);
xnor U7305 (N_7305,N_7112,N_7140);
nor U7306 (N_7306,N_7065,N_7080);
nor U7307 (N_7307,N_7120,N_7171);
nand U7308 (N_7308,N_7135,N_7108);
xnor U7309 (N_7309,N_7060,N_7108);
and U7310 (N_7310,N_7108,N_7165);
and U7311 (N_7311,N_7094,N_7097);
xor U7312 (N_7312,N_7068,N_7127);
xor U7313 (N_7313,N_7125,N_7145);
nand U7314 (N_7314,N_7181,N_7069);
xnor U7315 (N_7315,N_7126,N_7161);
nand U7316 (N_7316,N_7117,N_7085);
and U7317 (N_7317,N_7098,N_7075);
nand U7318 (N_7318,N_7128,N_7045);
or U7319 (N_7319,N_7042,N_7154);
nand U7320 (N_7320,N_7073,N_7048);
or U7321 (N_7321,N_7170,N_7107);
and U7322 (N_7322,N_7088,N_7127);
xor U7323 (N_7323,N_7059,N_7108);
nand U7324 (N_7324,N_7188,N_7152);
xor U7325 (N_7325,N_7152,N_7059);
nand U7326 (N_7326,N_7078,N_7042);
and U7327 (N_7327,N_7145,N_7053);
xor U7328 (N_7328,N_7190,N_7194);
xor U7329 (N_7329,N_7130,N_7195);
xnor U7330 (N_7330,N_7137,N_7071);
nand U7331 (N_7331,N_7185,N_7138);
and U7332 (N_7332,N_7088,N_7122);
nor U7333 (N_7333,N_7130,N_7163);
and U7334 (N_7334,N_7089,N_7069);
and U7335 (N_7335,N_7133,N_7044);
and U7336 (N_7336,N_7173,N_7166);
or U7337 (N_7337,N_7055,N_7042);
nor U7338 (N_7338,N_7138,N_7109);
xor U7339 (N_7339,N_7103,N_7181);
nand U7340 (N_7340,N_7083,N_7118);
or U7341 (N_7341,N_7059,N_7166);
xor U7342 (N_7342,N_7150,N_7184);
or U7343 (N_7343,N_7163,N_7180);
or U7344 (N_7344,N_7074,N_7048);
or U7345 (N_7345,N_7177,N_7173);
nor U7346 (N_7346,N_7186,N_7054);
nand U7347 (N_7347,N_7186,N_7104);
nor U7348 (N_7348,N_7134,N_7130);
nor U7349 (N_7349,N_7098,N_7170);
nor U7350 (N_7350,N_7061,N_7131);
xnor U7351 (N_7351,N_7160,N_7114);
nor U7352 (N_7352,N_7162,N_7196);
nor U7353 (N_7353,N_7129,N_7119);
and U7354 (N_7354,N_7058,N_7148);
xor U7355 (N_7355,N_7089,N_7199);
nor U7356 (N_7356,N_7135,N_7055);
and U7357 (N_7357,N_7150,N_7130);
or U7358 (N_7358,N_7068,N_7179);
and U7359 (N_7359,N_7106,N_7081);
nor U7360 (N_7360,N_7332,N_7301);
or U7361 (N_7361,N_7270,N_7343);
and U7362 (N_7362,N_7353,N_7218);
nor U7363 (N_7363,N_7355,N_7222);
nand U7364 (N_7364,N_7302,N_7297);
nor U7365 (N_7365,N_7305,N_7235);
and U7366 (N_7366,N_7225,N_7217);
xor U7367 (N_7367,N_7313,N_7293);
xor U7368 (N_7368,N_7358,N_7249);
and U7369 (N_7369,N_7203,N_7333);
and U7370 (N_7370,N_7321,N_7295);
nand U7371 (N_7371,N_7221,N_7340);
and U7372 (N_7372,N_7334,N_7344);
and U7373 (N_7373,N_7245,N_7226);
xor U7374 (N_7374,N_7207,N_7335);
nand U7375 (N_7375,N_7350,N_7261);
or U7376 (N_7376,N_7288,N_7247);
nor U7377 (N_7377,N_7357,N_7312);
and U7378 (N_7378,N_7338,N_7346);
nand U7379 (N_7379,N_7291,N_7205);
or U7380 (N_7380,N_7352,N_7204);
or U7381 (N_7381,N_7265,N_7224);
xor U7382 (N_7382,N_7267,N_7330);
nand U7383 (N_7383,N_7317,N_7231);
nand U7384 (N_7384,N_7213,N_7239);
nand U7385 (N_7385,N_7264,N_7228);
or U7386 (N_7386,N_7215,N_7345);
or U7387 (N_7387,N_7274,N_7242);
nor U7388 (N_7388,N_7342,N_7243);
nand U7389 (N_7389,N_7262,N_7292);
and U7390 (N_7390,N_7303,N_7287);
xnor U7391 (N_7391,N_7266,N_7285);
nand U7392 (N_7392,N_7256,N_7223);
xnor U7393 (N_7393,N_7209,N_7227);
and U7394 (N_7394,N_7331,N_7329);
nor U7395 (N_7395,N_7210,N_7282);
nor U7396 (N_7396,N_7253,N_7351);
nand U7397 (N_7397,N_7319,N_7233);
and U7398 (N_7398,N_7212,N_7324);
xnor U7399 (N_7399,N_7259,N_7252);
xnor U7400 (N_7400,N_7281,N_7220);
xor U7401 (N_7401,N_7237,N_7298);
or U7402 (N_7402,N_7279,N_7339);
or U7403 (N_7403,N_7219,N_7254);
xor U7404 (N_7404,N_7310,N_7251);
xor U7405 (N_7405,N_7286,N_7208);
nor U7406 (N_7406,N_7269,N_7202);
or U7407 (N_7407,N_7234,N_7258);
or U7408 (N_7408,N_7216,N_7246);
or U7409 (N_7409,N_7277,N_7325);
nand U7410 (N_7410,N_7236,N_7314);
nor U7411 (N_7411,N_7296,N_7309);
xor U7412 (N_7412,N_7276,N_7229);
or U7413 (N_7413,N_7348,N_7308);
xor U7414 (N_7414,N_7318,N_7257);
nand U7415 (N_7415,N_7290,N_7241);
or U7416 (N_7416,N_7271,N_7349);
xnor U7417 (N_7417,N_7206,N_7322);
and U7418 (N_7418,N_7230,N_7304);
nor U7419 (N_7419,N_7201,N_7328);
nor U7420 (N_7420,N_7300,N_7248);
and U7421 (N_7421,N_7275,N_7278);
nand U7422 (N_7422,N_7240,N_7356);
nand U7423 (N_7423,N_7268,N_7200);
nor U7424 (N_7424,N_7359,N_7323);
nand U7425 (N_7425,N_7284,N_7347);
or U7426 (N_7426,N_7294,N_7214);
xor U7427 (N_7427,N_7283,N_7273);
nand U7428 (N_7428,N_7280,N_7341);
xor U7429 (N_7429,N_7336,N_7307);
and U7430 (N_7430,N_7354,N_7316);
or U7431 (N_7431,N_7211,N_7232);
and U7432 (N_7432,N_7327,N_7326);
and U7433 (N_7433,N_7289,N_7311);
nand U7434 (N_7434,N_7263,N_7315);
nor U7435 (N_7435,N_7306,N_7272);
and U7436 (N_7436,N_7238,N_7299);
xor U7437 (N_7437,N_7320,N_7260);
nand U7438 (N_7438,N_7255,N_7244);
or U7439 (N_7439,N_7250,N_7337);
and U7440 (N_7440,N_7239,N_7200);
nand U7441 (N_7441,N_7301,N_7231);
xnor U7442 (N_7442,N_7330,N_7336);
or U7443 (N_7443,N_7244,N_7281);
xor U7444 (N_7444,N_7300,N_7354);
and U7445 (N_7445,N_7278,N_7292);
or U7446 (N_7446,N_7254,N_7232);
nor U7447 (N_7447,N_7243,N_7256);
and U7448 (N_7448,N_7346,N_7305);
or U7449 (N_7449,N_7333,N_7286);
nand U7450 (N_7450,N_7244,N_7276);
nand U7451 (N_7451,N_7249,N_7276);
xor U7452 (N_7452,N_7277,N_7333);
or U7453 (N_7453,N_7326,N_7325);
xnor U7454 (N_7454,N_7259,N_7323);
xor U7455 (N_7455,N_7335,N_7264);
and U7456 (N_7456,N_7319,N_7260);
nand U7457 (N_7457,N_7267,N_7351);
or U7458 (N_7458,N_7228,N_7218);
nor U7459 (N_7459,N_7337,N_7295);
nor U7460 (N_7460,N_7210,N_7243);
xnor U7461 (N_7461,N_7210,N_7236);
and U7462 (N_7462,N_7283,N_7206);
xor U7463 (N_7463,N_7333,N_7295);
and U7464 (N_7464,N_7327,N_7208);
xnor U7465 (N_7465,N_7276,N_7214);
xor U7466 (N_7466,N_7325,N_7297);
and U7467 (N_7467,N_7224,N_7264);
nand U7468 (N_7468,N_7282,N_7237);
nand U7469 (N_7469,N_7302,N_7345);
or U7470 (N_7470,N_7295,N_7223);
nor U7471 (N_7471,N_7243,N_7261);
and U7472 (N_7472,N_7277,N_7278);
nor U7473 (N_7473,N_7271,N_7251);
and U7474 (N_7474,N_7353,N_7340);
xnor U7475 (N_7475,N_7214,N_7355);
or U7476 (N_7476,N_7210,N_7214);
nor U7477 (N_7477,N_7231,N_7359);
xnor U7478 (N_7478,N_7233,N_7262);
nor U7479 (N_7479,N_7232,N_7222);
nand U7480 (N_7480,N_7229,N_7254);
xor U7481 (N_7481,N_7253,N_7290);
or U7482 (N_7482,N_7352,N_7288);
nand U7483 (N_7483,N_7303,N_7229);
and U7484 (N_7484,N_7242,N_7284);
and U7485 (N_7485,N_7315,N_7250);
xor U7486 (N_7486,N_7250,N_7307);
or U7487 (N_7487,N_7320,N_7327);
nor U7488 (N_7488,N_7356,N_7232);
nand U7489 (N_7489,N_7274,N_7271);
and U7490 (N_7490,N_7202,N_7309);
xnor U7491 (N_7491,N_7238,N_7235);
and U7492 (N_7492,N_7257,N_7272);
and U7493 (N_7493,N_7335,N_7334);
nor U7494 (N_7494,N_7293,N_7259);
and U7495 (N_7495,N_7206,N_7310);
nand U7496 (N_7496,N_7282,N_7234);
nor U7497 (N_7497,N_7219,N_7348);
xnor U7498 (N_7498,N_7288,N_7356);
or U7499 (N_7499,N_7351,N_7259);
xor U7500 (N_7500,N_7207,N_7206);
nand U7501 (N_7501,N_7350,N_7317);
xor U7502 (N_7502,N_7202,N_7205);
and U7503 (N_7503,N_7225,N_7342);
and U7504 (N_7504,N_7317,N_7338);
xnor U7505 (N_7505,N_7358,N_7288);
nor U7506 (N_7506,N_7272,N_7241);
and U7507 (N_7507,N_7329,N_7279);
nor U7508 (N_7508,N_7333,N_7216);
or U7509 (N_7509,N_7272,N_7210);
nor U7510 (N_7510,N_7309,N_7321);
nand U7511 (N_7511,N_7268,N_7329);
xnor U7512 (N_7512,N_7202,N_7324);
or U7513 (N_7513,N_7267,N_7292);
nand U7514 (N_7514,N_7245,N_7333);
nand U7515 (N_7515,N_7353,N_7267);
nor U7516 (N_7516,N_7254,N_7313);
and U7517 (N_7517,N_7278,N_7294);
and U7518 (N_7518,N_7231,N_7259);
and U7519 (N_7519,N_7326,N_7332);
nor U7520 (N_7520,N_7397,N_7462);
nand U7521 (N_7521,N_7499,N_7437);
nand U7522 (N_7522,N_7360,N_7458);
nor U7523 (N_7523,N_7387,N_7472);
and U7524 (N_7524,N_7488,N_7408);
or U7525 (N_7525,N_7477,N_7423);
xor U7526 (N_7526,N_7413,N_7382);
nor U7527 (N_7527,N_7398,N_7506);
or U7528 (N_7528,N_7438,N_7420);
xnor U7529 (N_7529,N_7431,N_7485);
and U7530 (N_7530,N_7516,N_7426);
or U7531 (N_7531,N_7491,N_7367);
nor U7532 (N_7532,N_7518,N_7374);
or U7533 (N_7533,N_7368,N_7419);
or U7534 (N_7534,N_7452,N_7505);
and U7535 (N_7535,N_7492,N_7464);
nand U7536 (N_7536,N_7370,N_7441);
nand U7537 (N_7537,N_7376,N_7473);
and U7538 (N_7538,N_7468,N_7509);
and U7539 (N_7539,N_7510,N_7489);
nor U7540 (N_7540,N_7500,N_7502);
or U7541 (N_7541,N_7519,N_7475);
and U7542 (N_7542,N_7504,N_7384);
or U7543 (N_7543,N_7386,N_7372);
or U7544 (N_7544,N_7471,N_7383);
or U7545 (N_7545,N_7493,N_7400);
nand U7546 (N_7546,N_7385,N_7416);
nand U7547 (N_7547,N_7361,N_7483);
xnor U7548 (N_7548,N_7381,N_7402);
nand U7549 (N_7549,N_7453,N_7389);
xnor U7550 (N_7550,N_7494,N_7508);
or U7551 (N_7551,N_7414,N_7495);
xnor U7552 (N_7552,N_7394,N_7364);
xor U7553 (N_7553,N_7448,N_7478);
or U7554 (N_7554,N_7362,N_7399);
nor U7555 (N_7555,N_7430,N_7380);
and U7556 (N_7556,N_7435,N_7517);
and U7557 (N_7557,N_7422,N_7439);
nand U7558 (N_7558,N_7424,N_7403);
xnor U7559 (N_7559,N_7490,N_7487);
or U7560 (N_7560,N_7404,N_7444);
xor U7561 (N_7561,N_7465,N_7445);
nand U7562 (N_7562,N_7486,N_7451);
and U7563 (N_7563,N_7363,N_7480);
and U7564 (N_7564,N_7456,N_7371);
xnor U7565 (N_7565,N_7469,N_7421);
xnor U7566 (N_7566,N_7467,N_7474);
nor U7567 (N_7567,N_7406,N_7391);
and U7568 (N_7568,N_7513,N_7410);
nand U7569 (N_7569,N_7375,N_7440);
xnor U7570 (N_7570,N_7425,N_7482);
nor U7571 (N_7571,N_7390,N_7412);
xnor U7572 (N_7572,N_7377,N_7470);
and U7573 (N_7573,N_7395,N_7393);
xor U7574 (N_7574,N_7476,N_7411);
nand U7575 (N_7575,N_7378,N_7511);
xor U7576 (N_7576,N_7457,N_7432);
nor U7577 (N_7577,N_7479,N_7442);
xnor U7578 (N_7578,N_7466,N_7455);
xnor U7579 (N_7579,N_7436,N_7514);
and U7580 (N_7580,N_7461,N_7396);
nand U7581 (N_7581,N_7459,N_7501);
nand U7582 (N_7582,N_7407,N_7481);
and U7583 (N_7583,N_7460,N_7388);
and U7584 (N_7584,N_7507,N_7405);
nor U7585 (N_7585,N_7433,N_7515);
xnor U7586 (N_7586,N_7365,N_7418);
nand U7587 (N_7587,N_7409,N_7369);
and U7588 (N_7588,N_7496,N_7415);
and U7589 (N_7589,N_7512,N_7428);
xor U7590 (N_7590,N_7366,N_7434);
or U7591 (N_7591,N_7447,N_7497);
or U7592 (N_7592,N_7401,N_7449);
or U7593 (N_7593,N_7417,N_7450);
nand U7594 (N_7594,N_7427,N_7484);
nand U7595 (N_7595,N_7446,N_7379);
and U7596 (N_7596,N_7429,N_7498);
xnor U7597 (N_7597,N_7392,N_7463);
nand U7598 (N_7598,N_7454,N_7443);
and U7599 (N_7599,N_7503,N_7373);
or U7600 (N_7600,N_7465,N_7494);
and U7601 (N_7601,N_7460,N_7459);
xor U7602 (N_7602,N_7420,N_7374);
or U7603 (N_7603,N_7483,N_7378);
nand U7604 (N_7604,N_7386,N_7425);
xor U7605 (N_7605,N_7478,N_7495);
nor U7606 (N_7606,N_7452,N_7497);
nor U7607 (N_7607,N_7488,N_7367);
and U7608 (N_7608,N_7382,N_7486);
or U7609 (N_7609,N_7442,N_7451);
or U7610 (N_7610,N_7451,N_7498);
nand U7611 (N_7611,N_7436,N_7453);
or U7612 (N_7612,N_7364,N_7482);
xor U7613 (N_7613,N_7376,N_7501);
or U7614 (N_7614,N_7382,N_7510);
or U7615 (N_7615,N_7421,N_7500);
nor U7616 (N_7616,N_7378,N_7405);
xnor U7617 (N_7617,N_7481,N_7396);
and U7618 (N_7618,N_7410,N_7459);
xor U7619 (N_7619,N_7470,N_7366);
nor U7620 (N_7620,N_7444,N_7518);
xor U7621 (N_7621,N_7417,N_7477);
nor U7622 (N_7622,N_7469,N_7386);
nor U7623 (N_7623,N_7473,N_7420);
xor U7624 (N_7624,N_7445,N_7456);
nor U7625 (N_7625,N_7492,N_7439);
and U7626 (N_7626,N_7388,N_7509);
xor U7627 (N_7627,N_7451,N_7472);
nand U7628 (N_7628,N_7492,N_7502);
and U7629 (N_7629,N_7499,N_7383);
nand U7630 (N_7630,N_7502,N_7416);
or U7631 (N_7631,N_7398,N_7501);
or U7632 (N_7632,N_7478,N_7470);
nor U7633 (N_7633,N_7516,N_7469);
and U7634 (N_7634,N_7443,N_7372);
and U7635 (N_7635,N_7422,N_7428);
xnor U7636 (N_7636,N_7486,N_7360);
xnor U7637 (N_7637,N_7398,N_7406);
nand U7638 (N_7638,N_7447,N_7467);
or U7639 (N_7639,N_7503,N_7513);
xor U7640 (N_7640,N_7402,N_7473);
nand U7641 (N_7641,N_7414,N_7428);
xor U7642 (N_7642,N_7506,N_7391);
nor U7643 (N_7643,N_7402,N_7415);
or U7644 (N_7644,N_7504,N_7405);
or U7645 (N_7645,N_7485,N_7519);
xnor U7646 (N_7646,N_7442,N_7375);
or U7647 (N_7647,N_7496,N_7416);
and U7648 (N_7648,N_7391,N_7501);
xor U7649 (N_7649,N_7489,N_7504);
nand U7650 (N_7650,N_7437,N_7408);
nand U7651 (N_7651,N_7457,N_7369);
or U7652 (N_7652,N_7456,N_7422);
and U7653 (N_7653,N_7499,N_7400);
nor U7654 (N_7654,N_7409,N_7425);
and U7655 (N_7655,N_7371,N_7501);
or U7656 (N_7656,N_7512,N_7489);
and U7657 (N_7657,N_7466,N_7464);
nand U7658 (N_7658,N_7403,N_7515);
and U7659 (N_7659,N_7400,N_7438);
or U7660 (N_7660,N_7400,N_7451);
nor U7661 (N_7661,N_7488,N_7497);
nand U7662 (N_7662,N_7492,N_7380);
xnor U7663 (N_7663,N_7504,N_7465);
xnor U7664 (N_7664,N_7441,N_7388);
nor U7665 (N_7665,N_7403,N_7417);
and U7666 (N_7666,N_7424,N_7418);
and U7667 (N_7667,N_7455,N_7379);
nand U7668 (N_7668,N_7477,N_7450);
and U7669 (N_7669,N_7419,N_7423);
nor U7670 (N_7670,N_7420,N_7518);
xnor U7671 (N_7671,N_7369,N_7500);
xor U7672 (N_7672,N_7386,N_7367);
xnor U7673 (N_7673,N_7402,N_7502);
nand U7674 (N_7674,N_7479,N_7383);
xor U7675 (N_7675,N_7492,N_7453);
and U7676 (N_7676,N_7399,N_7419);
xor U7677 (N_7677,N_7389,N_7377);
nor U7678 (N_7678,N_7463,N_7514);
nand U7679 (N_7679,N_7426,N_7420);
nor U7680 (N_7680,N_7534,N_7642);
xor U7681 (N_7681,N_7582,N_7672);
nor U7682 (N_7682,N_7538,N_7613);
nand U7683 (N_7683,N_7541,N_7654);
nor U7684 (N_7684,N_7599,N_7609);
nand U7685 (N_7685,N_7675,N_7676);
nor U7686 (N_7686,N_7547,N_7602);
nor U7687 (N_7687,N_7583,N_7567);
or U7688 (N_7688,N_7542,N_7604);
or U7689 (N_7689,N_7625,N_7590);
or U7690 (N_7690,N_7563,N_7608);
nand U7691 (N_7691,N_7656,N_7624);
nor U7692 (N_7692,N_7611,N_7657);
xnor U7693 (N_7693,N_7537,N_7647);
or U7694 (N_7694,N_7655,N_7557);
nand U7695 (N_7695,N_7545,N_7548);
xor U7696 (N_7696,N_7650,N_7559);
and U7697 (N_7697,N_7635,N_7525);
or U7698 (N_7698,N_7522,N_7575);
and U7699 (N_7699,N_7673,N_7619);
or U7700 (N_7700,N_7598,N_7528);
xnor U7701 (N_7701,N_7668,N_7586);
nor U7702 (N_7702,N_7531,N_7651);
nor U7703 (N_7703,N_7580,N_7550);
or U7704 (N_7704,N_7544,N_7562);
nand U7705 (N_7705,N_7576,N_7627);
and U7706 (N_7706,N_7595,N_7622);
nor U7707 (N_7707,N_7593,N_7539);
or U7708 (N_7708,N_7558,N_7589);
nor U7709 (N_7709,N_7520,N_7612);
xnor U7710 (N_7710,N_7653,N_7596);
nand U7711 (N_7711,N_7638,N_7665);
or U7712 (N_7712,N_7588,N_7618);
nor U7713 (N_7713,N_7524,N_7570);
xnor U7714 (N_7714,N_7597,N_7523);
or U7715 (N_7715,N_7561,N_7662);
nor U7716 (N_7716,N_7551,N_7643);
and U7717 (N_7717,N_7664,N_7636);
xor U7718 (N_7718,N_7634,N_7587);
nand U7719 (N_7719,N_7565,N_7535);
or U7720 (N_7720,N_7584,N_7614);
nor U7721 (N_7721,N_7617,N_7637);
xor U7722 (N_7722,N_7574,N_7641);
nor U7723 (N_7723,N_7639,N_7526);
nor U7724 (N_7724,N_7601,N_7566);
or U7725 (N_7725,N_7629,N_7573);
nand U7726 (N_7726,N_7667,N_7671);
xor U7727 (N_7727,N_7533,N_7630);
or U7728 (N_7728,N_7530,N_7615);
and U7729 (N_7729,N_7646,N_7555);
nor U7730 (N_7730,N_7592,N_7652);
and U7731 (N_7731,N_7633,N_7677);
xnor U7732 (N_7732,N_7577,N_7674);
nand U7733 (N_7733,N_7554,N_7564);
xnor U7734 (N_7734,N_7594,N_7591);
nand U7735 (N_7735,N_7581,N_7628);
nand U7736 (N_7736,N_7670,N_7659);
and U7737 (N_7737,N_7529,N_7623);
nor U7738 (N_7738,N_7666,N_7663);
and U7739 (N_7739,N_7521,N_7600);
xnor U7740 (N_7740,N_7532,N_7556);
nor U7741 (N_7741,N_7669,N_7540);
or U7742 (N_7742,N_7632,N_7527);
or U7743 (N_7743,N_7585,N_7605);
xnor U7744 (N_7744,N_7536,N_7571);
nor U7745 (N_7745,N_7640,N_7660);
nand U7746 (N_7746,N_7607,N_7661);
and U7747 (N_7747,N_7616,N_7644);
nand U7748 (N_7748,N_7645,N_7678);
or U7749 (N_7749,N_7560,N_7648);
xnor U7750 (N_7750,N_7631,N_7621);
nor U7751 (N_7751,N_7572,N_7626);
and U7752 (N_7752,N_7569,N_7603);
nor U7753 (N_7753,N_7543,N_7679);
or U7754 (N_7754,N_7620,N_7579);
nand U7755 (N_7755,N_7610,N_7549);
xnor U7756 (N_7756,N_7606,N_7649);
nor U7757 (N_7757,N_7568,N_7578);
xnor U7758 (N_7758,N_7553,N_7552);
nand U7759 (N_7759,N_7658,N_7546);
nor U7760 (N_7760,N_7522,N_7606);
nand U7761 (N_7761,N_7673,N_7592);
xnor U7762 (N_7762,N_7554,N_7567);
or U7763 (N_7763,N_7555,N_7664);
nor U7764 (N_7764,N_7596,N_7542);
xnor U7765 (N_7765,N_7520,N_7646);
nor U7766 (N_7766,N_7545,N_7587);
and U7767 (N_7767,N_7539,N_7660);
or U7768 (N_7768,N_7567,N_7607);
nor U7769 (N_7769,N_7535,N_7587);
nand U7770 (N_7770,N_7670,N_7587);
nor U7771 (N_7771,N_7612,N_7580);
nand U7772 (N_7772,N_7644,N_7538);
nand U7773 (N_7773,N_7592,N_7626);
nor U7774 (N_7774,N_7663,N_7535);
xor U7775 (N_7775,N_7555,N_7586);
nor U7776 (N_7776,N_7658,N_7607);
xnor U7777 (N_7777,N_7618,N_7675);
xnor U7778 (N_7778,N_7559,N_7525);
xnor U7779 (N_7779,N_7580,N_7552);
nor U7780 (N_7780,N_7612,N_7654);
and U7781 (N_7781,N_7613,N_7571);
or U7782 (N_7782,N_7618,N_7615);
nand U7783 (N_7783,N_7592,N_7607);
xnor U7784 (N_7784,N_7580,N_7538);
xnor U7785 (N_7785,N_7553,N_7576);
and U7786 (N_7786,N_7593,N_7639);
and U7787 (N_7787,N_7568,N_7607);
nand U7788 (N_7788,N_7630,N_7635);
or U7789 (N_7789,N_7612,N_7615);
nand U7790 (N_7790,N_7579,N_7527);
nand U7791 (N_7791,N_7522,N_7566);
and U7792 (N_7792,N_7630,N_7634);
xor U7793 (N_7793,N_7554,N_7649);
nor U7794 (N_7794,N_7601,N_7609);
or U7795 (N_7795,N_7665,N_7643);
xor U7796 (N_7796,N_7636,N_7576);
nor U7797 (N_7797,N_7605,N_7610);
nand U7798 (N_7798,N_7606,N_7550);
or U7799 (N_7799,N_7607,N_7610);
or U7800 (N_7800,N_7617,N_7566);
and U7801 (N_7801,N_7662,N_7677);
and U7802 (N_7802,N_7549,N_7619);
or U7803 (N_7803,N_7579,N_7665);
nand U7804 (N_7804,N_7617,N_7528);
and U7805 (N_7805,N_7673,N_7542);
nand U7806 (N_7806,N_7544,N_7598);
nand U7807 (N_7807,N_7528,N_7534);
xor U7808 (N_7808,N_7555,N_7616);
and U7809 (N_7809,N_7598,N_7623);
nor U7810 (N_7810,N_7539,N_7622);
nor U7811 (N_7811,N_7541,N_7564);
and U7812 (N_7812,N_7524,N_7589);
nand U7813 (N_7813,N_7679,N_7576);
or U7814 (N_7814,N_7674,N_7645);
xnor U7815 (N_7815,N_7611,N_7599);
nor U7816 (N_7816,N_7606,N_7577);
nand U7817 (N_7817,N_7539,N_7608);
nor U7818 (N_7818,N_7599,N_7657);
xor U7819 (N_7819,N_7654,N_7552);
nor U7820 (N_7820,N_7647,N_7667);
and U7821 (N_7821,N_7582,N_7649);
nand U7822 (N_7822,N_7566,N_7567);
xnor U7823 (N_7823,N_7614,N_7568);
nor U7824 (N_7824,N_7528,N_7557);
nor U7825 (N_7825,N_7523,N_7532);
nor U7826 (N_7826,N_7525,N_7659);
xnor U7827 (N_7827,N_7563,N_7541);
nand U7828 (N_7828,N_7537,N_7660);
xor U7829 (N_7829,N_7555,N_7658);
xor U7830 (N_7830,N_7521,N_7565);
and U7831 (N_7831,N_7565,N_7677);
nor U7832 (N_7832,N_7645,N_7561);
or U7833 (N_7833,N_7585,N_7592);
and U7834 (N_7834,N_7627,N_7539);
or U7835 (N_7835,N_7549,N_7572);
nand U7836 (N_7836,N_7602,N_7620);
or U7837 (N_7837,N_7582,N_7529);
nand U7838 (N_7838,N_7562,N_7664);
or U7839 (N_7839,N_7586,N_7588);
nor U7840 (N_7840,N_7834,N_7783);
or U7841 (N_7841,N_7757,N_7761);
xor U7842 (N_7842,N_7787,N_7755);
xor U7843 (N_7843,N_7770,N_7774);
nor U7844 (N_7844,N_7736,N_7717);
or U7845 (N_7845,N_7709,N_7752);
and U7846 (N_7846,N_7792,N_7700);
or U7847 (N_7847,N_7695,N_7747);
nand U7848 (N_7848,N_7714,N_7782);
xnor U7849 (N_7849,N_7828,N_7748);
nor U7850 (N_7850,N_7772,N_7708);
or U7851 (N_7851,N_7825,N_7735);
nand U7852 (N_7852,N_7687,N_7703);
nand U7853 (N_7853,N_7730,N_7771);
or U7854 (N_7854,N_7765,N_7740);
xnor U7855 (N_7855,N_7822,N_7727);
or U7856 (N_7856,N_7820,N_7753);
nor U7857 (N_7857,N_7726,N_7724);
or U7858 (N_7858,N_7722,N_7713);
or U7859 (N_7859,N_7759,N_7811);
or U7860 (N_7860,N_7728,N_7816);
nor U7861 (N_7861,N_7710,N_7680);
or U7862 (N_7862,N_7694,N_7784);
or U7863 (N_7863,N_7763,N_7777);
nor U7864 (N_7864,N_7821,N_7810);
nand U7865 (N_7865,N_7809,N_7804);
nor U7866 (N_7866,N_7684,N_7795);
and U7867 (N_7867,N_7823,N_7829);
and U7868 (N_7868,N_7781,N_7775);
nor U7869 (N_7869,N_7754,N_7734);
nand U7870 (N_7870,N_7723,N_7690);
and U7871 (N_7871,N_7686,N_7705);
or U7872 (N_7872,N_7788,N_7746);
and U7873 (N_7873,N_7815,N_7762);
or U7874 (N_7874,N_7803,N_7769);
nor U7875 (N_7875,N_7702,N_7758);
nor U7876 (N_7876,N_7779,N_7812);
xor U7877 (N_7877,N_7786,N_7701);
nor U7878 (N_7878,N_7835,N_7744);
or U7879 (N_7879,N_7760,N_7745);
and U7880 (N_7880,N_7827,N_7793);
nor U7881 (N_7881,N_7737,N_7826);
nand U7882 (N_7882,N_7798,N_7729);
and U7883 (N_7883,N_7718,N_7790);
nand U7884 (N_7884,N_7682,N_7692);
nand U7885 (N_7885,N_7697,N_7824);
and U7886 (N_7886,N_7768,N_7681);
nor U7887 (N_7887,N_7807,N_7685);
nor U7888 (N_7888,N_7691,N_7813);
or U7889 (N_7889,N_7805,N_7696);
xor U7890 (N_7890,N_7808,N_7741);
or U7891 (N_7891,N_7756,N_7800);
or U7892 (N_7892,N_7789,N_7731);
and U7893 (N_7893,N_7819,N_7716);
nand U7894 (N_7894,N_7780,N_7721);
nand U7895 (N_7895,N_7720,N_7725);
or U7896 (N_7896,N_7683,N_7773);
and U7897 (N_7897,N_7833,N_7806);
xnor U7898 (N_7898,N_7719,N_7839);
nor U7899 (N_7899,N_7818,N_7704);
or U7900 (N_7900,N_7832,N_7776);
or U7901 (N_7901,N_7796,N_7711);
nor U7902 (N_7902,N_7698,N_7739);
xnor U7903 (N_7903,N_7688,N_7764);
nand U7904 (N_7904,N_7794,N_7751);
nor U7905 (N_7905,N_7732,N_7814);
or U7906 (N_7906,N_7699,N_7749);
nand U7907 (N_7907,N_7785,N_7743);
nand U7908 (N_7908,N_7837,N_7766);
nor U7909 (N_7909,N_7838,N_7801);
nand U7910 (N_7910,N_7767,N_7707);
or U7911 (N_7911,N_7706,N_7830);
nor U7912 (N_7912,N_7715,N_7836);
nand U7913 (N_7913,N_7750,N_7712);
nand U7914 (N_7914,N_7791,N_7778);
and U7915 (N_7915,N_7733,N_7742);
nor U7916 (N_7916,N_7738,N_7693);
xnor U7917 (N_7917,N_7802,N_7797);
nor U7918 (N_7918,N_7689,N_7799);
nor U7919 (N_7919,N_7831,N_7817);
nand U7920 (N_7920,N_7738,N_7720);
nand U7921 (N_7921,N_7687,N_7757);
or U7922 (N_7922,N_7720,N_7689);
nor U7923 (N_7923,N_7797,N_7781);
nand U7924 (N_7924,N_7715,N_7807);
nand U7925 (N_7925,N_7752,N_7760);
nand U7926 (N_7926,N_7691,N_7745);
and U7927 (N_7927,N_7812,N_7734);
xnor U7928 (N_7928,N_7695,N_7833);
or U7929 (N_7929,N_7704,N_7759);
nand U7930 (N_7930,N_7804,N_7783);
and U7931 (N_7931,N_7715,N_7749);
nor U7932 (N_7932,N_7680,N_7744);
nor U7933 (N_7933,N_7695,N_7717);
or U7934 (N_7934,N_7816,N_7741);
and U7935 (N_7935,N_7835,N_7721);
nor U7936 (N_7936,N_7819,N_7743);
xor U7937 (N_7937,N_7704,N_7765);
nor U7938 (N_7938,N_7707,N_7689);
nor U7939 (N_7939,N_7759,N_7793);
nor U7940 (N_7940,N_7685,N_7710);
or U7941 (N_7941,N_7831,N_7774);
xor U7942 (N_7942,N_7732,N_7734);
nand U7943 (N_7943,N_7765,N_7766);
xnor U7944 (N_7944,N_7691,N_7690);
nor U7945 (N_7945,N_7706,N_7773);
nor U7946 (N_7946,N_7764,N_7740);
xnor U7947 (N_7947,N_7695,N_7701);
nor U7948 (N_7948,N_7751,N_7704);
xnor U7949 (N_7949,N_7739,N_7757);
xnor U7950 (N_7950,N_7784,N_7824);
xnor U7951 (N_7951,N_7828,N_7760);
nand U7952 (N_7952,N_7726,N_7828);
xor U7953 (N_7953,N_7707,N_7747);
or U7954 (N_7954,N_7700,N_7702);
and U7955 (N_7955,N_7826,N_7772);
or U7956 (N_7956,N_7782,N_7721);
or U7957 (N_7957,N_7824,N_7707);
nor U7958 (N_7958,N_7769,N_7693);
and U7959 (N_7959,N_7774,N_7751);
nor U7960 (N_7960,N_7701,N_7809);
and U7961 (N_7961,N_7709,N_7687);
nor U7962 (N_7962,N_7690,N_7686);
nor U7963 (N_7963,N_7712,N_7710);
and U7964 (N_7964,N_7717,N_7710);
xor U7965 (N_7965,N_7684,N_7753);
or U7966 (N_7966,N_7704,N_7827);
xor U7967 (N_7967,N_7827,N_7744);
or U7968 (N_7968,N_7784,N_7819);
xor U7969 (N_7969,N_7747,N_7832);
xnor U7970 (N_7970,N_7788,N_7771);
and U7971 (N_7971,N_7713,N_7824);
and U7972 (N_7972,N_7746,N_7711);
xor U7973 (N_7973,N_7742,N_7763);
and U7974 (N_7974,N_7706,N_7814);
xnor U7975 (N_7975,N_7729,N_7741);
nand U7976 (N_7976,N_7720,N_7742);
and U7977 (N_7977,N_7792,N_7707);
and U7978 (N_7978,N_7811,N_7817);
nand U7979 (N_7979,N_7727,N_7763);
nor U7980 (N_7980,N_7727,N_7735);
and U7981 (N_7981,N_7716,N_7780);
nor U7982 (N_7982,N_7824,N_7821);
nor U7983 (N_7983,N_7834,N_7823);
and U7984 (N_7984,N_7681,N_7803);
nand U7985 (N_7985,N_7682,N_7817);
xor U7986 (N_7986,N_7739,N_7785);
or U7987 (N_7987,N_7730,N_7806);
or U7988 (N_7988,N_7838,N_7820);
xnor U7989 (N_7989,N_7804,N_7767);
nand U7990 (N_7990,N_7760,N_7764);
nand U7991 (N_7991,N_7726,N_7765);
and U7992 (N_7992,N_7743,N_7700);
xnor U7993 (N_7993,N_7685,N_7735);
nand U7994 (N_7994,N_7794,N_7791);
nor U7995 (N_7995,N_7807,N_7832);
nor U7996 (N_7996,N_7781,N_7808);
xnor U7997 (N_7997,N_7808,N_7715);
or U7998 (N_7998,N_7762,N_7775);
nor U7999 (N_7999,N_7699,N_7692);
nand U8000 (N_8000,N_7934,N_7981);
or U8001 (N_8001,N_7841,N_7988);
and U8002 (N_8002,N_7983,N_7850);
xnor U8003 (N_8003,N_7951,N_7987);
nand U8004 (N_8004,N_7902,N_7868);
nor U8005 (N_8005,N_7991,N_7974);
or U8006 (N_8006,N_7979,N_7944);
nor U8007 (N_8007,N_7863,N_7899);
xnor U8008 (N_8008,N_7845,N_7886);
or U8009 (N_8009,N_7962,N_7923);
and U8010 (N_8010,N_7905,N_7939);
nor U8011 (N_8011,N_7970,N_7954);
nor U8012 (N_8012,N_7937,N_7892);
nand U8013 (N_8013,N_7842,N_7897);
and U8014 (N_8014,N_7953,N_7906);
nor U8015 (N_8015,N_7921,N_7877);
or U8016 (N_8016,N_7949,N_7948);
nand U8017 (N_8017,N_7849,N_7919);
xnor U8018 (N_8018,N_7881,N_7958);
and U8019 (N_8019,N_7967,N_7916);
or U8020 (N_8020,N_7992,N_7936);
and U8021 (N_8021,N_7858,N_7920);
xor U8022 (N_8022,N_7993,N_7990);
xor U8023 (N_8023,N_7903,N_7908);
or U8024 (N_8024,N_7853,N_7888);
nand U8025 (N_8025,N_7966,N_7938);
nand U8026 (N_8026,N_7895,N_7940);
nor U8027 (N_8027,N_7980,N_7866);
nand U8028 (N_8028,N_7932,N_7875);
nand U8029 (N_8029,N_7865,N_7977);
nor U8030 (N_8030,N_7880,N_7896);
or U8031 (N_8031,N_7976,N_7843);
xor U8032 (N_8032,N_7887,N_7969);
nor U8033 (N_8033,N_7847,N_7885);
nand U8034 (N_8034,N_7846,N_7884);
nor U8035 (N_8035,N_7960,N_7848);
and U8036 (N_8036,N_7851,N_7869);
and U8037 (N_8037,N_7968,N_7947);
and U8038 (N_8038,N_7931,N_7874);
xor U8039 (N_8039,N_7894,N_7956);
xor U8040 (N_8040,N_7864,N_7942);
and U8041 (N_8041,N_7996,N_7840);
xor U8042 (N_8042,N_7889,N_7882);
or U8043 (N_8043,N_7891,N_7873);
or U8044 (N_8044,N_7964,N_7989);
and U8045 (N_8045,N_7860,N_7898);
and U8046 (N_8046,N_7872,N_7900);
xor U8047 (N_8047,N_7867,N_7876);
or U8048 (N_8048,N_7859,N_7998);
nand U8049 (N_8049,N_7972,N_7924);
or U8050 (N_8050,N_7963,N_7950);
nand U8051 (N_8051,N_7878,N_7943);
and U8052 (N_8052,N_7984,N_7922);
nor U8053 (N_8053,N_7999,N_7927);
xor U8054 (N_8054,N_7933,N_7925);
and U8055 (N_8055,N_7857,N_7883);
xor U8056 (N_8056,N_7852,N_7854);
xnor U8057 (N_8057,N_7971,N_7918);
xnor U8058 (N_8058,N_7870,N_7911);
xor U8059 (N_8059,N_7965,N_7862);
nand U8060 (N_8060,N_7909,N_7904);
nor U8061 (N_8061,N_7890,N_7959);
nand U8062 (N_8062,N_7945,N_7941);
or U8063 (N_8063,N_7844,N_7926);
nand U8064 (N_8064,N_7861,N_7997);
xnor U8065 (N_8065,N_7871,N_7917);
nand U8066 (N_8066,N_7982,N_7957);
or U8067 (N_8067,N_7907,N_7978);
nor U8068 (N_8068,N_7893,N_7955);
and U8069 (N_8069,N_7912,N_7973);
xnor U8070 (N_8070,N_7986,N_7901);
xor U8071 (N_8071,N_7995,N_7946);
and U8072 (N_8072,N_7914,N_7855);
and U8073 (N_8073,N_7935,N_7915);
or U8074 (N_8074,N_7913,N_7985);
nor U8075 (N_8075,N_7856,N_7929);
nand U8076 (N_8076,N_7952,N_7910);
and U8077 (N_8077,N_7961,N_7975);
xnor U8078 (N_8078,N_7928,N_7930);
xor U8079 (N_8079,N_7879,N_7994);
or U8080 (N_8080,N_7924,N_7881);
nand U8081 (N_8081,N_7948,N_7864);
or U8082 (N_8082,N_7912,N_7872);
xor U8083 (N_8083,N_7969,N_7954);
and U8084 (N_8084,N_7884,N_7865);
nor U8085 (N_8085,N_7931,N_7960);
and U8086 (N_8086,N_7841,N_7850);
or U8087 (N_8087,N_7916,N_7989);
nor U8088 (N_8088,N_7914,N_7875);
xor U8089 (N_8089,N_7995,N_7871);
xnor U8090 (N_8090,N_7900,N_7844);
and U8091 (N_8091,N_7927,N_7920);
nor U8092 (N_8092,N_7957,N_7859);
nand U8093 (N_8093,N_7885,N_7891);
nor U8094 (N_8094,N_7899,N_7918);
nand U8095 (N_8095,N_7845,N_7987);
and U8096 (N_8096,N_7980,N_7957);
xnor U8097 (N_8097,N_7966,N_7891);
xnor U8098 (N_8098,N_7954,N_7876);
nand U8099 (N_8099,N_7973,N_7905);
or U8100 (N_8100,N_7966,N_7985);
xnor U8101 (N_8101,N_7894,N_7899);
and U8102 (N_8102,N_7991,N_7891);
xnor U8103 (N_8103,N_7992,N_7942);
nand U8104 (N_8104,N_7916,N_7998);
nand U8105 (N_8105,N_7927,N_7985);
nor U8106 (N_8106,N_7888,N_7917);
nor U8107 (N_8107,N_7967,N_7948);
or U8108 (N_8108,N_7977,N_7949);
nor U8109 (N_8109,N_7858,N_7851);
xnor U8110 (N_8110,N_7845,N_7950);
nor U8111 (N_8111,N_7869,N_7938);
xnor U8112 (N_8112,N_7928,N_7882);
xnor U8113 (N_8113,N_7855,N_7929);
xor U8114 (N_8114,N_7907,N_7859);
nand U8115 (N_8115,N_7934,N_7962);
nand U8116 (N_8116,N_7899,N_7980);
or U8117 (N_8117,N_7859,N_7840);
xnor U8118 (N_8118,N_7896,N_7871);
and U8119 (N_8119,N_7873,N_7862);
nor U8120 (N_8120,N_7907,N_7869);
nor U8121 (N_8121,N_7909,N_7940);
xor U8122 (N_8122,N_7956,N_7927);
nand U8123 (N_8123,N_7958,N_7918);
xnor U8124 (N_8124,N_7895,N_7941);
xor U8125 (N_8125,N_7862,N_7856);
nor U8126 (N_8126,N_7889,N_7848);
xnor U8127 (N_8127,N_7901,N_7984);
xnor U8128 (N_8128,N_7975,N_7984);
nand U8129 (N_8129,N_7988,N_7979);
nor U8130 (N_8130,N_7855,N_7938);
or U8131 (N_8131,N_7871,N_7983);
nor U8132 (N_8132,N_7974,N_7851);
and U8133 (N_8133,N_7991,N_7951);
or U8134 (N_8134,N_7909,N_7910);
or U8135 (N_8135,N_7957,N_7911);
nor U8136 (N_8136,N_7939,N_7880);
and U8137 (N_8137,N_7875,N_7841);
or U8138 (N_8138,N_7943,N_7914);
nand U8139 (N_8139,N_7895,N_7844);
and U8140 (N_8140,N_7935,N_7869);
nand U8141 (N_8141,N_7859,N_7982);
or U8142 (N_8142,N_7983,N_7928);
nor U8143 (N_8143,N_7869,N_7972);
and U8144 (N_8144,N_7902,N_7951);
or U8145 (N_8145,N_7852,N_7976);
xor U8146 (N_8146,N_7938,N_7879);
or U8147 (N_8147,N_7971,N_7879);
xor U8148 (N_8148,N_7862,N_7933);
nor U8149 (N_8149,N_7874,N_7893);
nor U8150 (N_8150,N_7975,N_7884);
nor U8151 (N_8151,N_7974,N_7928);
nor U8152 (N_8152,N_7913,N_7980);
nand U8153 (N_8153,N_7849,N_7879);
or U8154 (N_8154,N_7844,N_7986);
and U8155 (N_8155,N_7861,N_7955);
or U8156 (N_8156,N_7845,N_7854);
and U8157 (N_8157,N_7944,N_7966);
nor U8158 (N_8158,N_7940,N_7971);
xor U8159 (N_8159,N_7993,N_7954);
and U8160 (N_8160,N_8091,N_8151);
and U8161 (N_8161,N_8002,N_8017);
xnor U8162 (N_8162,N_8059,N_8090);
xnor U8163 (N_8163,N_8148,N_8044);
or U8164 (N_8164,N_8115,N_8133);
and U8165 (N_8165,N_8086,N_8088);
nor U8166 (N_8166,N_8014,N_8146);
nor U8167 (N_8167,N_8049,N_8134);
nand U8168 (N_8168,N_8104,N_8031);
xnor U8169 (N_8169,N_8008,N_8034);
nand U8170 (N_8170,N_8022,N_8021);
and U8171 (N_8171,N_8157,N_8046);
nand U8172 (N_8172,N_8035,N_8135);
nand U8173 (N_8173,N_8120,N_8058);
nor U8174 (N_8174,N_8089,N_8041);
xnor U8175 (N_8175,N_8142,N_8095);
or U8176 (N_8176,N_8074,N_8042);
or U8177 (N_8177,N_8145,N_8079);
xnor U8178 (N_8178,N_8136,N_8103);
nor U8179 (N_8179,N_8124,N_8073);
nor U8180 (N_8180,N_8101,N_8153);
nand U8181 (N_8181,N_8139,N_8118);
nand U8182 (N_8182,N_8123,N_8083);
or U8183 (N_8183,N_8030,N_8040);
xnor U8184 (N_8184,N_8075,N_8102);
or U8185 (N_8185,N_8077,N_8066);
or U8186 (N_8186,N_8043,N_8117);
xnor U8187 (N_8187,N_8070,N_8098);
xor U8188 (N_8188,N_8093,N_8019);
or U8189 (N_8189,N_8149,N_8111);
nand U8190 (N_8190,N_8065,N_8011);
nand U8191 (N_8191,N_8045,N_8025);
and U8192 (N_8192,N_8023,N_8147);
and U8193 (N_8193,N_8051,N_8055);
and U8194 (N_8194,N_8010,N_8052);
xnor U8195 (N_8195,N_8009,N_8027);
nand U8196 (N_8196,N_8116,N_8112);
nor U8197 (N_8197,N_8105,N_8140);
xnor U8198 (N_8198,N_8080,N_8039);
or U8199 (N_8199,N_8113,N_8012);
xnor U8200 (N_8200,N_8015,N_8159);
or U8201 (N_8201,N_8057,N_8024);
xor U8202 (N_8202,N_8053,N_8128);
or U8203 (N_8203,N_8050,N_8082);
and U8204 (N_8204,N_8106,N_8003);
or U8205 (N_8205,N_8069,N_8028);
nand U8206 (N_8206,N_8063,N_8132);
or U8207 (N_8207,N_8006,N_8062);
or U8208 (N_8208,N_8097,N_8158);
and U8209 (N_8209,N_8000,N_8130);
nor U8210 (N_8210,N_8122,N_8054);
or U8211 (N_8211,N_8143,N_8068);
nor U8212 (N_8212,N_8016,N_8005);
and U8213 (N_8213,N_8129,N_8107);
nand U8214 (N_8214,N_8141,N_8131);
and U8215 (N_8215,N_8036,N_8154);
xnor U8216 (N_8216,N_8020,N_8018);
and U8217 (N_8217,N_8108,N_8109);
xor U8218 (N_8218,N_8047,N_8144);
and U8219 (N_8219,N_8152,N_8156);
and U8220 (N_8220,N_8138,N_8007);
nand U8221 (N_8221,N_8067,N_8061);
xor U8222 (N_8222,N_8004,N_8032);
nand U8223 (N_8223,N_8064,N_8110);
nand U8224 (N_8224,N_8126,N_8084);
xnor U8225 (N_8225,N_8085,N_8076);
and U8226 (N_8226,N_8001,N_8078);
nor U8227 (N_8227,N_8155,N_8121);
xnor U8228 (N_8228,N_8026,N_8100);
xor U8229 (N_8229,N_8013,N_8094);
or U8230 (N_8230,N_8033,N_8137);
nor U8231 (N_8231,N_8071,N_8127);
or U8232 (N_8232,N_8087,N_8081);
or U8233 (N_8233,N_8038,N_8125);
or U8234 (N_8234,N_8056,N_8060);
nor U8235 (N_8235,N_8092,N_8048);
xnor U8236 (N_8236,N_8114,N_8119);
and U8237 (N_8237,N_8072,N_8099);
nand U8238 (N_8238,N_8029,N_8037);
or U8239 (N_8239,N_8150,N_8096);
and U8240 (N_8240,N_8100,N_8090);
and U8241 (N_8241,N_8108,N_8159);
xnor U8242 (N_8242,N_8030,N_8092);
nor U8243 (N_8243,N_8037,N_8106);
nand U8244 (N_8244,N_8053,N_8055);
or U8245 (N_8245,N_8077,N_8146);
or U8246 (N_8246,N_8097,N_8036);
or U8247 (N_8247,N_8084,N_8121);
and U8248 (N_8248,N_8120,N_8004);
and U8249 (N_8249,N_8116,N_8104);
nor U8250 (N_8250,N_8145,N_8070);
nand U8251 (N_8251,N_8059,N_8031);
nand U8252 (N_8252,N_8129,N_8143);
or U8253 (N_8253,N_8030,N_8071);
and U8254 (N_8254,N_8060,N_8015);
xnor U8255 (N_8255,N_8044,N_8037);
nand U8256 (N_8256,N_8005,N_8000);
nor U8257 (N_8257,N_8019,N_8084);
and U8258 (N_8258,N_8031,N_8112);
and U8259 (N_8259,N_8020,N_8101);
nand U8260 (N_8260,N_8047,N_8135);
or U8261 (N_8261,N_8069,N_8015);
and U8262 (N_8262,N_8025,N_8090);
or U8263 (N_8263,N_8151,N_8093);
nand U8264 (N_8264,N_8152,N_8083);
nand U8265 (N_8265,N_8063,N_8009);
or U8266 (N_8266,N_8048,N_8021);
nand U8267 (N_8267,N_8005,N_8135);
nor U8268 (N_8268,N_8003,N_8024);
xnor U8269 (N_8269,N_8074,N_8072);
nand U8270 (N_8270,N_8050,N_8132);
nor U8271 (N_8271,N_8031,N_8060);
xor U8272 (N_8272,N_8061,N_8158);
nor U8273 (N_8273,N_8117,N_8084);
and U8274 (N_8274,N_8070,N_8102);
or U8275 (N_8275,N_8031,N_8078);
or U8276 (N_8276,N_8135,N_8158);
nor U8277 (N_8277,N_8105,N_8123);
or U8278 (N_8278,N_8106,N_8108);
xnor U8279 (N_8279,N_8024,N_8109);
or U8280 (N_8280,N_8030,N_8016);
nand U8281 (N_8281,N_8054,N_8095);
and U8282 (N_8282,N_8105,N_8088);
nand U8283 (N_8283,N_8120,N_8082);
nand U8284 (N_8284,N_8071,N_8113);
or U8285 (N_8285,N_8129,N_8005);
nor U8286 (N_8286,N_8026,N_8088);
nor U8287 (N_8287,N_8082,N_8159);
and U8288 (N_8288,N_8017,N_8053);
nor U8289 (N_8289,N_8131,N_8064);
nand U8290 (N_8290,N_8134,N_8009);
nor U8291 (N_8291,N_8046,N_8114);
xnor U8292 (N_8292,N_8049,N_8023);
nor U8293 (N_8293,N_8023,N_8146);
and U8294 (N_8294,N_8084,N_8012);
xor U8295 (N_8295,N_8149,N_8082);
or U8296 (N_8296,N_8033,N_8153);
nand U8297 (N_8297,N_8001,N_8114);
nand U8298 (N_8298,N_8037,N_8077);
and U8299 (N_8299,N_8076,N_8136);
and U8300 (N_8300,N_8157,N_8120);
xnor U8301 (N_8301,N_8144,N_8027);
nand U8302 (N_8302,N_8022,N_8113);
and U8303 (N_8303,N_8072,N_8109);
or U8304 (N_8304,N_8033,N_8094);
nor U8305 (N_8305,N_8123,N_8121);
nand U8306 (N_8306,N_8124,N_8153);
and U8307 (N_8307,N_8154,N_8043);
or U8308 (N_8308,N_8035,N_8003);
nand U8309 (N_8309,N_8012,N_8131);
xnor U8310 (N_8310,N_8074,N_8019);
nand U8311 (N_8311,N_8076,N_8084);
nand U8312 (N_8312,N_8121,N_8012);
and U8313 (N_8313,N_8124,N_8063);
nor U8314 (N_8314,N_8150,N_8139);
or U8315 (N_8315,N_8064,N_8126);
nor U8316 (N_8316,N_8048,N_8084);
or U8317 (N_8317,N_8004,N_8146);
nor U8318 (N_8318,N_8149,N_8136);
nor U8319 (N_8319,N_8137,N_8122);
nand U8320 (N_8320,N_8191,N_8245);
nand U8321 (N_8321,N_8319,N_8196);
nor U8322 (N_8322,N_8175,N_8195);
nor U8323 (N_8323,N_8273,N_8225);
or U8324 (N_8324,N_8298,N_8295);
or U8325 (N_8325,N_8262,N_8186);
or U8326 (N_8326,N_8258,N_8270);
or U8327 (N_8327,N_8251,N_8274);
or U8328 (N_8328,N_8250,N_8279);
nor U8329 (N_8329,N_8170,N_8254);
nand U8330 (N_8330,N_8162,N_8236);
or U8331 (N_8331,N_8198,N_8306);
and U8332 (N_8332,N_8311,N_8315);
xnor U8333 (N_8333,N_8210,N_8242);
nand U8334 (N_8334,N_8266,N_8228);
nand U8335 (N_8335,N_8163,N_8260);
nor U8336 (N_8336,N_8271,N_8265);
nand U8337 (N_8337,N_8207,N_8220);
xor U8338 (N_8338,N_8178,N_8215);
or U8339 (N_8339,N_8172,N_8256);
xor U8340 (N_8340,N_8278,N_8310);
xor U8341 (N_8341,N_8253,N_8219);
nor U8342 (N_8342,N_8307,N_8272);
nor U8343 (N_8343,N_8188,N_8283);
or U8344 (N_8344,N_8249,N_8232);
nand U8345 (N_8345,N_8229,N_8248);
nor U8346 (N_8346,N_8259,N_8177);
nand U8347 (N_8347,N_8240,N_8282);
xor U8348 (N_8348,N_8281,N_8230);
nor U8349 (N_8349,N_8200,N_8314);
xor U8350 (N_8350,N_8164,N_8287);
xnor U8351 (N_8351,N_8189,N_8179);
nand U8352 (N_8352,N_8199,N_8174);
and U8353 (N_8353,N_8204,N_8197);
xor U8354 (N_8354,N_8261,N_8194);
nand U8355 (N_8355,N_8302,N_8277);
xor U8356 (N_8356,N_8161,N_8231);
and U8357 (N_8357,N_8305,N_8297);
nor U8358 (N_8358,N_8268,N_8214);
or U8359 (N_8359,N_8203,N_8299);
nor U8360 (N_8360,N_8185,N_8289);
xnor U8361 (N_8361,N_8309,N_8316);
xnor U8362 (N_8362,N_8171,N_8290);
nand U8363 (N_8363,N_8317,N_8224);
nor U8364 (N_8364,N_8184,N_8233);
and U8365 (N_8365,N_8255,N_8308);
and U8366 (N_8366,N_8166,N_8180);
and U8367 (N_8367,N_8201,N_8173);
and U8368 (N_8368,N_8280,N_8226);
nand U8369 (N_8369,N_8167,N_8190);
nand U8370 (N_8370,N_8304,N_8244);
xor U8371 (N_8371,N_8264,N_8303);
nor U8372 (N_8372,N_8318,N_8252);
or U8373 (N_8373,N_8294,N_8176);
nand U8374 (N_8374,N_8227,N_8206);
or U8375 (N_8375,N_8243,N_8312);
nand U8376 (N_8376,N_8285,N_8181);
or U8377 (N_8377,N_8218,N_8241);
nand U8378 (N_8378,N_8238,N_8239);
nand U8379 (N_8379,N_8301,N_8237);
and U8380 (N_8380,N_8183,N_8288);
nor U8381 (N_8381,N_8292,N_8205);
xnor U8382 (N_8382,N_8182,N_8257);
and U8383 (N_8383,N_8269,N_8234);
or U8384 (N_8384,N_8276,N_8275);
or U8385 (N_8385,N_8216,N_8217);
nand U8386 (N_8386,N_8209,N_8160);
nor U8387 (N_8387,N_8263,N_8202);
or U8388 (N_8388,N_8313,N_8213);
and U8389 (N_8389,N_8193,N_8267);
and U8390 (N_8390,N_8247,N_8296);
nor U8391 (N_8391,N_8187,N_8223);
xor U8392 (N_8392,N_8165,N_8291);
and U8393 (N_8393,N_8221,N_8212);
nor U8394 (N_8394,N_8246,N_8222);
and U8395 (N_8395,N_8235,N_8300);
nor U8396 (N_8396,N_8211,N_8169);
nor U8397 (N_8397,N_8284,N_8168);
or U8398 (N_8398,N_8208,N_8192);
xnor U8399 (N_8399,N_8293,N_8286);
xnor U8400 (N_8400,N_8163,N_8222);
or U8401 (N_8401,N_8166,N_8238);
xnor U8402 (N_8402,N_8312,N_8317);
or U8403 (N_8403,N_8248,N_8192);
nor U8404 (N_8404,N_8293,N_8304);
nand U8405 (N_8405,N_8207,N_8208);
and U8406 (N_8406,N_8246,N_8319);
nor U8407 (N_8407,N_8227,N_8274);
nor U8408 (N_8408,N_8315,N_8192);
and U8409 (N_8409,N_8195,N_8166);
nor U8410 (N_8410,N_8301,N_8259);
and U8411 (N_8411,N_8319,N_8219);
nor U8412 (N_8412,N_8270,N_8264);
nor U8413 (N_8413,N_8319,N_8311);
xnor U8414 (N_8414,N_8171,N_8208);
nor U8415 (N_8415,N_8295,N_8288);
nand U8416 (N_8416,N_8293,N_8213);
xnor U8417 (N_8417,N_8273,N_8253);
or U8418 (N_8418,N_8196,N_8247);
nand U8419 (N_8419,N_8162,N_8271);
or U8420 (N_8420,N_8186,N_8160);
nor U8421 (N_8421,N_8273,N_8218);
and U8422 (N_8422,N_8266,N_8283);
or U8423 (N_8423,N_8303,N_8233);
nand U8424 (N_8424,N_8264,N_8283);
nor U8425 (N_8425,N_8299,N_8230);
nor U8426 (N_8426,N_8296,N_8269);
and U8427 (N_8427,N_8243,N_8279);
xor U8428 (N_8428,N_8245,N_8228);
xnor U8429 (N_8429,N_8242,N_8237);
nand U8430 (N_8430,N_8223,N_8196);
nor U8431 (N_8431,N_8197,N_8191);
and U8432 (N_8432,N_8293,N_8275);
and U8433 (N_8433,N_8176,N_8226);
nand U8434 (N_8434,N_8207,N_8196);
nor U8435 (N_8435,N_8309,N_8206);
and U8436 (N_8436,N_8257,N_8319);
xnor U8437 (N_8437,N_8176,N_8284);
xor U8438 (N_8438,N_8206,N_8268);
or U8439 (N_8439,N_8234,N_8279);
and U8440 (N_8440,N_8201,N_8291);
or U8441 (N_8441,N_8304,N_8261);
xnor U8442 (N_8442,N_8288,N_8191);
xnor U8443 (N_8443,N_8259,N_8169);
or U8444 (N_8444,N_8239,N_8269);
or U8445 (N_8445,N_8239,N_8202);
xor U8446 (N_8446,N_8285,N_8315);
xnor U8447 (N_8447,N_8224,N_8288);
and U8448 (N_8448,N_8222,N_8183);
xor U8449 (N_8449,N_8313,N_8265);
xnor U8450 (N_8450,N_8221,N_8209);
and U8451 (N_8451,N_8207,N_8246);
and U8452 (N_8452,N_8242,N_8172);
and U8453 (N_8453,N_8244,N_8197);
and U8454 (N_8454,N_8241,N_8268);
or U8455 (N_8455,N_8306,N_8278);
nand U8456 (N_8456,N_8241,N_8260);
nor U8457 (N_8457,N_8176,N_8248);
nand U8458 (N_8458,N_8234,N_8222);
xnor U8459 (N_8459,N_8172,N_8235);
and U8460 (N_8460,N_8278,N_8181);
and U8461 (N_8461,N_8215,N_8225);
and U8462 (N_8462,N_8297,N_8201);
or U8463 (N_8463,N_8206,N_8241);
nor U8464 (N_8464,N_8170,N_8173);
nor U8465 (N_8465,N_8262,N_8260);
xnor U8466 (N_8466,N_8232,N_8299);
and U8467 (N_8467,N_8285,N_8316);
or U8468 (N_8468,N_8300,N_8178);
nand U8469 (N_8469,N_8280,N_8307);
and U8470 (N_8470,N_8245,N_8301);
or U8471 (N_8471,N_8214,N_8160);
nor U8472 (N_8472,N_8303,N_8249);
and U8473 (N_8473,N_8200,N_8245);
nor U8474 (N_8474,N_8213,N_8285);
xnor U8475 (N_8475,N_8223,N_8195);
or U8476 (N_8476,N_8168,N_8262);
and U8477 (N_8477,N_8289,N_8222);
nand U8478 (N_8478,N_8220,N_8284);
nand U8479 (N_8479,N_8188,N_8262);
or U8480 (N_8480,N_8474,N_8390);
nand U8481 (N_8481,N_8436,N_8462);
nor U8482 (N_8482,N_8472,N_8378);
or U8483 (N_8483,N_8381,N_8428);
nand U8484 (N_8484,N_8404,N_8401);
or U8485 (N_8485,N_8322,N_8418);
and U8486 (N_8486,N_8456,N_8422);
nor U8487 (N_8487,N_8446,N_8426);
nor U8488 (N_8488,N_8415,N_8324);
xor U8489 (N_8489,N_8377,N_8445);
and U8490 (N_8490,N_8343,N_8367);
nor U8491 (N_8491,N_8361,N_8414);
and U8492 (N_8492,N_8452,N_8321);
and U8493 (N_8493,N_8346,N_8339);
nand U8494 (N_8494,N_8337,N_8368);
nor U8495 (N_8495,N_8443,N_8475);
or U8496 (N_8496,N_8429,N_8478);
or U8497 (N_8497,N_8357,N_8435);
xnor U8498 (N_8498,N_8387,N_8326);
or U8499 (N_8499,N_8396,N_8420);
xnor U8500 (N_8500,N_8331,N_8402);
nor U8501 (N_8501,N_8416,N_8391);
and U8502 (N_8502,N_8458,N_8385);
nor U8503 (N_8503,N_8364,N_8388);
or U8504 (N_8504,N_8374,N_8406);
xor U8505 (N_8505,N_8354,N_8350);
and U8506 (N_8506,N_8338,N_8463);
and U8507 (N_8507,N_8470,N_8469);
or U8508 (N_8508,N_8425,N_8461);
nand U8509 (N_8509,N_8379,N_8464);
xnor U8510 (N_8510,N_8359,N_8448);
nand U8511 (N_8511,N_8467,N_8408);
nand U8512 (N_8512,N_8392,N_8423);
xor U8513 (N_8513,N_8410,N_8449);
or U8514 (N_8514,N_8457,N_8444);
xor U8515 (N_8515,N_8413,N_8356);
xnor U8516 (N_8516,N_8330,N_8333);
nand U8517 (N_8517,N_8382,N_8434);
nand U8518 (N_8518,N_8348,N_8431);
nand U8519 (N_8519,N_8440,N_8328);
xnor U8520 (N_8520,N_8439,N_8340);
and U8521 (N_8521,N_8427,N_8366);
or U8522 (N_8522,N_8351,N_8369);
nand U8523 (N_8523,N_8344,N_8471);
nor U8524 (N_8524,N_8375,N_8355);
nor U8525 (N_8525,N_8332,N_8373);
or U8526 (N_8526,N_8384,N_8336);
or U8527 (N_8527,N_8419,N_8397);
or U8528 (N_8528,N_8454,N_8399);
xnor U8529 (N_8529,N_8451,N_8409);
xor U8530 (N_8530,N_8342,N_8335);
or U8531 (N_8531,N_8400,N_8447);
nand U8532 (N_8532,N_8412,N_8341);
nor U8533 (N_8533,N_8479,N_8398);
nand U8534 (N_8534,N_8386,N_8365);
xnor U8535 (N_8535,N_8353,N_8352);
and U8536 (N_8536,N_8349,N_8421);
nand U8537 (N_8537,N_8380,N_8320);
nor U8538 (N_8538,N_8459,N_8395);
or U8539 (N_8539,N_8473,N_8468);
xor U8540 (N_8540,N_8477,N_8327);
or U8541 (N_8541,N_8433,N_8325);
or U8542 (N_8542,N_8389,N_8363);
and U8543 (N_8543,N_8323,N_8358);
nor U8544 (N_8544,N_8460,N_8405);
nor U8545 (N_8545,N_8371,N_8432);
or U8546 (N_8546,N_8394,N_8362);
nand U8547 (N_8547,N_8372,N_8441);
nor U8548 (N_8548,N_8424,N_8437);
nor U8549 (N_8549,N_8360,N_8403);
xnor U8550 (N_8550,N_8466,N_8370);
nor U8551 (N_8551,N_8442,N_8376);
nand U8552 (N_8552,N_8455,N_8465);
nor U8553 (N_8553,N_8417,N_8430);
and U8554 (N_8554,N_8347,N_8453);
or U8555 (N_8555,N_8450,N_8345);
nand U8556 (N_8556,N_8476,N_8393);
xor U8557 (N_8557,N_8438,N_8334);
nor U8558 (N_8558,N_8329,N_8383);
xnor U8559 (N_8559,N_8407,N_8411);
xor U8560 (N_8560,N_8423,N_8446);
and U8561 (N_8561,N_8341,N_8437);
xor U8562 (N_8562,N_8424,N_8350);
xor U8563 (N_8563,N_8477,N_8408);
or U8564 (N_8564,N_8474,N_8445);
xor U8565 (N_8565,N_8442,N_8455);
or U8566 (N_8566,N_8404,N_8341);
nor U8567 (N_8567,N_8448,N_8376);
xor U8568 (N_8568,N_8408,N_8434);
nor U8569 (N_8569,N_8416,N_8448);
or U8570 (N_8570,N_8336,N_8343);
or U8571 (N_8571,N_8377,N_8419);
and U8572 (N_8572,N_8464,N_8425);
or U8573 (N_8573,N_8424,N_8341);
xnor U8574 (N_8574,N_8360,N_8392);
and U8575 (N_8575,N_8456,N_8392);
or U8576 (N_8576,N_8340,N_8459);
and U8577 (N_8577,N_8432,N_8451);
xor U8578 (N_8578,N_8434,N_8457);
or U8579 (N_8579,N_8421,N_8391);
nor U8580 (N_8580,N_8367,N_8377);
xor U8581 (N_8581,N_8476,N_8391);
or U8582 (N_8582,N_8395,N_8412);
nor U8583 (N_8583,N_8372,N_8394);
or U8584 (N_8584,N_8383,N_8399);
and U8585 (N_8585,N_8358,N_8429);
or U8586 (N_8586,N_8410,N_8382);
and U8587 (N_8587,N_8323,N_8346);
nand U8588 (N_8588,N_8479,N_8329);
nand U8589 (N_8589,N_8330,N_8353);
or U8590 (N_8590,N_8421,N_8371);
and U8591 (N_8591,N_8425,N_8466);
xnor U8592 (N_8592,N_8460,N_8388);
and U8593 (N_8593,N_8473,N_8400);
nor U8594 (N_8594,N_8351,N_8458);
xnor U8595 (N_8595,N_8385,N_8436);
nand U8596 (N_8596,N_8357,N_8436);
or U8597 (N_8597,N_8384,N_8405);
nor U8598 (N_8598,N_8338,N_8390);
nor U8599 (N_8599,N_8465,N_8429);
nand U8600 (N_8600,N_8362,N_8345);
or U8601 (N_8601,N_8443,N_8442);
xor U8602 (N_8602,N_8448,N_8378);
nand U8603 (N_8603,N_8442,N_8396);
and U8604 (N_8604,N_8350,N_8431);
or U8605 (N_8605,N_8438,N_8423);
nand U8606 (N_8606,N_8340,N_8350);
or U8607 (N_8607,N_8396,N_8364);
nand U8608 (N_8608,N_8357,N_8321);
or U8609 (N_8609,N_8422,N_8325);
and U8610 (N_8610,N_8360,N_8387);
nand U8611 (N_8611,N_8425,N_8321);
nor U8612 (N_8612,N_8433,N_8321);
nor U8613 (N_8613,N_8452,N_8400);
and U8614 (N_8614,N_8394,N_8468);
xnor U8615 (N_8615,N_8455,N_8458);
and U8616 (N_8616,N_8327,N_8377);
nand U8617 (N_8617,N_8340,N_8358);
or U8618 (N_8618,N_8398,N_8362);
or U8619 (N_8619,N_8434,N_8385);
xnor U8620 (N_8620,N_8399,N_8451);
nand U8621 (N_8621,N_8446,N_8420);
or U8622 (N_8622,N_8349,N_8368);
and U8623 (N_8623,N_8397,N_8321);
nor U8624 (N_8624,N_8342,N_8422);
and U8625 (N_8625,N_8400,N_8389);
and U8626 (N_8626,N_8367,N_8411);
nand U8627 (N_8627,N_8387,N_8473);
and U8628 (N_8628,N_8450,N_8364);
xor U8629 (N_8629,N_8362,N_8353);
xor U8630 (N_8630,N_8390,N_8340);
nor U8631 (N_8631,N_8361,N_8432);
or U8632 (N_8632,N_8416,N_8376);
and U8633 (N_8633,N_8383,N_8458);
xnor U8634 (N_8634,N_8367,N_8478);
xor U8635 (N_8635,N_8389,N_8436);
nor U8636 (N_8636,N_8320,N_8405);
or U8637 (N_8637,N_8378,N_8466);
xnor U8638 (N_8638,N_8414,N_8374);
nand U8639 (N_8639,N_8418,N_8468);
xor U8640 (N_8640,N_8524,N_8558);
and U8641 (N_8641,N_8488,N_8588);
or U8642 (N_8642,N_8570,N_8516);
nand U8643 (N_8643,N_8624,N_8487);
nand U8644 (N_8644,N_8493,N_8636);
nor U8645 (N_8645,N_8566,N_8629);
nor U8646 (N_8646,N_8618,N_8527);
or U8647 (N_8647,N_8557,N_8484);
xor U8648 (N_8648,N_8633,N_8546);
or U8649 (N_8649,N_8512,N_8500);
nor U8650 (N_8650,N_8571,N_8533);
and U8651 (N_8651,N_8578,N_8601);
nor U8652 (N_8652,N_8537,N_8483);
nor U8653 (N_8653,N_8604,N_8541);
nor U8654 (N_8654,N_8494,N_8631);
and U8655 (N_8655,N_8506,N_8559);
nor U8656 (N_8656,N_8606,N_8562);
nand U8657 (N_8657,N_8542,N_8563);
nand U8658 (N_8658,N_8591,N_8523);
nand U8659 (N_8659,N_8637,N_8485);
and U8660 (N_8660,N_8480,N_8583);
nor U8661 (N_8661,N_8622,N_8498);
xnor U8662 (N_8662,N_8535,N_8615);
and U8663 (N_8663,N_8551,N_8573);
and U8664 (N_8664,N_8518,N_8491);
and U8665 (N_8665,N_8540,N_8539);
or U8666 (N_8666,N_8611,N_8590);
xnor U8667 (N_8667,N_8554,N_8536);
or U8668 (N_8668,N_8505,N_8628);
nor U8669 (N_8669,N_8592,N_8585);
xnor U8670 (N_8670,N_8482,N_8587);
and U8671 (N_8671,N_8614,N_8577);
xor U8672 (N_8672,N_8575,N_8579);
nor U8673 (N_8673,N_8596,N_8555);
and U8674 (N_8674,N_8502,N_8620);
xnor U8675 (N_8675,N_8564,N_8553);
and U8676 (N_8676,N_8521,N_8589);
xnor U8677 (N_8677,N_8621,N_8602);
nor U8678 (N_8678,N_8632,N_8567);
xnor U8679 (N_8679,N_8584,N_8515);
nand U8680 (N_8680,N_8513,N_8581);
nor U8681 (N_8681,N_8509,N_8550);
xnor U8682 (N_8682,N_8595,N_8528);
nand U8683 (N_8683,N_8538,N_8625);
and U8684 (N_8684,N_8569,N_8490);
nor U8685 (N_8685,N_8598,N_8489);
or U8686 (N_8686,N_8608,N_8607);
nand U8687 (N_8687,N_8568,N_8499);
and U8688 (N_8688,N_8612,N_8481);
and U8689 (N_8689,N_8630,N_8545);
and U8690 (N_8690,N_8508,N_8507);
nor U8691 (N_8691,N_8531,N_8639);
nand U8692 (N_8692,N_8603,N_8560);
and U8693 (N_8693,N_8617,N_8501);
nor U8694 (N_8694,N_8552,N_8548);
nor U8695 (N_8695,N_8549,N_8544);
or U8696 (N_8696,N_8580,N_8511);
and U8697 (N_8697,N_8486,N_8600);
and U8698 (N_8698,N_8634,N_8605);
nor U8699 (N_8699,N_8547,N_8635);
or U8700 (N_8700,N_8593,N_8503);
or U8701 (N_8701,N_8619,N_8530);
nand U8702 (N_8702,N_8532,N_8597);
nor U8703 (N_8703,N_8543,N_8576);
and U8704 (N_8704,N_8594,N_8556);
or U8705 (N_8705,N_8613,N_8517);
nand U8706 (N_8706,N_8510,N_8526);
nand U8707 (N_8707,N_8522,N_8525);
and U8708 (N_8708,N_8582,N_8609);
nand U8709 (N_8709,N_8504,N_8529);
nor U8710 (N_8710,N_8565,N_8561);
or U8711 (N_8711,N_8626,N_8627);
nor U8712 (N_8712,N_8520,N_8495);
nand U8713 (N_8713,N_8514,N_8519);
or U8714 (N_8714,N_8534,N_8638);
or U8715 (N_8715,N_8574,N_8496);
nand U8716 (N_8716,N_8497,N_8572);
or U8717 (N_8717,N_8586,N_8610);
xor U8718 (N_8718,N_8616,N_8599);
or U8719 (N_8719,N_8623,N_8492);
xnor U8720 (N_8720,N_8589,N_8593);
or U8721 (N_8721,N_8566,N_8484);
and U8722 (N_8722,N_8495,N_8517);
or U8723 (N_8723,N_8612,N_8579);
or U8724 (N_8724,N_8563,N_8624);
xnor U8725 (N_8725,N_8521,N_8634);
xnor U8726 (N_8726,N_8630,N_8543);
nor U8727 (N_8727,N_8506,N_8510);
nor U8728 (N_8728,N_8493,N_8629);
xor U8729 (N_8729,N_8553,N_8588);
nor U8730 (N_8730,N_8557,N_8639);
and U8731 (N_8731,N_8603,N_8629);
nor U8732 (N_8732,N_8504,N_8514);
nand U8733 (N_8733,N_8555,N_8578);
xnor U8734 (N_8734,N_8513,N_8611);
and U8735 (N_8735,N_8572,N_8629);
nor U8736 (N_8736,N_8605,N_8626);
and U8737 (N_8737,N_8585,N_8555);
nand U8738 (N_8738,N_8481,N_8579);
or U8739 (N_8739,N_8627,N_8611);
and U8740 (N_8740,N_8549,N_8588);
and U8741 (N_8741,N_8488,N_8594);
or U8742 (N_8742,N_8490,N_8507);
and U8743 (N_8743,N_8593,N_8596);
and U8744 (N_8744,N_8578,N_8548);
or U8745 (N_8745,N_8630,N_8599);
nor U8746 (N_8746,N_8519,N_8621);
nor U8747 (N_8747,N_8504,N_8563);
nor U8748 (N_8748,N_8504,N_8618);
nor U8749 (N_8749,N_8576,N_8503);
nand U8750 (N_8750,N_8551,N_8495);
xnor U8751 (N_8751,N_8622,N_8570);
nor U8752 (N_8752,N_8515,N_8490);
nand U8753 (N_8753,N_8549,N_8605);
nand U8754 (N_8754,N_8512,N_8612);
nor U8755 (N_8755,N_8620,N_8551);
nand U8756 (N_8756,N_8514,N_8589);
and U8757 (N_8757,N_8506,N_8633);
xnor U8758 (N_8758,N_8630,N_8618);
and U8759 (N_8759,N_8544,N_8587);
nor U8760 (N_8760,N_8549,N_8572);
or U8761 (N_8761,N_8576,N_8511);
nor U8762 (N_8762,N_8526,N_8586);
and U8763 (N_8763,N_8622,N_8547);
and U8764 (N_8764,N_8607,N_8585);
nand U8765 (N_8765,N_8596,N_8627);
nand U8766 (N_8766,N_8616,N_8535);
xor U8767 (N_8767,N_8532,N_8544);
nor U8768 (N_8768,N_8621,N_8565);
and U8769 (N_8769,N_8618,N_8492);
xor U8770 (N_8770,N_8581,N_8572);
or U8771 (N_8771,N_8518,N_8554);
or U8772 (N_8772,N_8499,N_8612);
nor U8773 (N_8773,N_8625,N_8505);
or U8774 (N_8774,N_8579,N_8484);
nor U8775 (N_8775,N_8616,N_8630);
xor U8776 (N_8776,N_8631,N_8622);
and U8777 (N_8777,N_8524,N_8596);
nor U8778 (N_8778,N_8565,N_8492);
nor U8779 (N_8779,N_8577,N_8631);
nor U8780 (N_8780,N_8494,N_8612);
nor U8781 (N_8781,N_8512,N_8561);
or U8782 (N_8782,N_8546,N_8621);
and U8783 (N_8783,N_8629,N_8595);
and U8784 (N_8784,N_8584,N_8587);
nor U8785 (N_8785,N_8534,N_8634);
xnor U8786 (N_8786,N_8519,N_8585);
xnor U8787 (N_8787,N_8497,N_8507);
or U8788 (N_8788,N_8602,N_8506);
nand U8789 (N_8789,N_8634,N_8483);
or U8790 (N_8790,N_8517,N_8588);
xnor U8791 (N_8791,N_8617,N_8534);
or U8792 (N_8792,N_8489,N_8619);
or U8793 (N_8793,N_8553,N_8635);
nor U8794 (N_8794,N_8576,N_8625);
and U8795 (N_8795,N_8561,N_8521);
or U8796 (N_8796,N_8635,N_8537);
nand U8797 (N_8797,N_8547,N_8490);
and U8798 (N_8798,N_8492,N_8559);
or U8799 (N_8799,N_8533,N_8576);
or U8800 (N_8800,N_8655,N_8685);
nor U8801 (N_8801,N_8703,N_8731);
xor U8802 (N_8802,N_8799,N_8708);
xnor U8803 (N_8803,N_8645,N_8663);
xnor U8804 (N_8804,N_8691,N_8762);
xnor U8805 (N_8805,N_8719,N_8758);
nor U8806 (N_8806,N_8756,N_8748);
nor U8807 (N_8807,N_8672,N_8650);
and U8808 (N_8808,N_8767,N_8796);
or U8809 (N_8809,N_8751,N_8694);
or U8810 (N_8810,N_8732,N_8724);
or U8811 (N_8811,N_8782,N_8714);
and U8812 (N_8812,N_8723,N_8797);
and U8813 (N_8813,N_8693,N_8681);
nand U8814 (N_8814,N_8749,N_8772);
nand U8815 (N_8815,N_8669,N_8664);
and U8816 (N_8816,N_8705,N_8690);
nand U8817 (N_8817,N_8730,N_8649);
or U8818 (N_8818,N_8768,N_8752);
or U8819 (N_8819,N_8774,N_8753);
nor U8820 (N_8820,N_8786,N_8793);
nand U8821 (N_8821,N_8735,N_8750);
or U8822 (N_8822,N_8795,N_8670);
and U8823 (N_8823,N_8711,N_8736);
or U8824 (N_8824,N_8646,N_8780);
nand U8825 (N_8825,N_8757,N_8783);
nor U8826 (N_8826,N_8653,N_8744);
nand U8827 (N_8827,N_8746,N_8642);
xor U8828 (N_8828,N_8759,N_8682);
and U8829 (N_8829,N_8671,N_8665);
or U8830 (N_8830,N_8721,N_8687);
xnor U8831 (N_8831,N_8712,N_8716);
and U8832 (N_8832,N_8688,N_8773);
nand U8833 (N_8833,N_8728,N_8722);
and U8834 (N_8834,N_8674,N_8769);
or U8835 (N_8835,N_8792,N_8763);
nand U8836 (N_8836,N_8738,N_8689);
nand U8837 (N_8837,N_8741,N_8779);
nor U8838 (N_8838,N_8745,N_8656);
and U8839 (N_8839,N_8776,N_8733);
nor U8840 (N_8840,N_8755,N_8666);
nor U8841 (N_8841,N_8676,N_8675);
nand U8842 (N_8842,N_8720,N_8704);
nand U8843 (N_8843,N_8667,N_8640);
nor U8844 (N_8844,N_8726,N_8789);
or U8845 (N_8845,N_8643,N_8775);
and U8846 (N_8846,N_8709,N_8662);
xnor U8847 (N_8847,N_8784,N_8654);
nor U8848 (N_8848,N_8700,N_8659);
or U8849 (N_8849,N_8715,N_8678);
or U8850 (N_8850,N_8686,N_8696);
and U8851 (N_8851,N_8760,N_8684);
nor U8852 (N_8852,N_8740,N_8707);
xor U8853 (N_8853,N_8764,N_8657);
nand U8854 (N_8854,N_8713,N_8699);
or U8855 (N_8855,N_8697,N_8641);
or U8856 (N_8856,N_8698,N_8710);
nand U8857 (N_8857,N_8771,N_8729);
xnor U8858 (N_8858,N_8677,N_8765);
nor U8859 (N_8859,N_8652,N_8647);
nand U8860 (N_8860,N_8701,N_8660);
and U8861 (N_8861,N_8785,N_8651);
or U8862 (N_8862,N_8798,N_8788);
and U8863 (N_8863,N_8787,N_8737);
nand U8864 (N_8864,N_8702,N_8692);
nand U8865 (N_8865,N_8742,N_8661);
nor U8866 (N_8866,N_8778,N_8747);
and U8867 (N_8867,N_8754,N_8790);
xnor U8868 (N_8868,N_8761,N_8770);
nand U8869 (N_8869,N_8734,N_8668);
or U8870 (N_8870,N_8743,N_8791);
nor U8871 (N_8871,N_8739,N_8644);
or U8872 (N_8872,N_8683,N_8725);
nor U8873 (N_8873,N_8673,N_8727);
or U8874 (N_8874,N_8781,N_8766);
and U8875 (N_8875,N_8794,N_8679);
nor U8876 (N_8876,N_8706,N_8695);
or U8877 (N_8877,N_8777,N_8658);
nand U8878 (N_8878,N_8680,N_8648);
or U8879 (N_8879,N_8718,N_8717);
xor U8880 (N_8880,N_8686,N_8672);
xnor U8881 (N_8881,N_8775,N_8662);
or U8882 (N_8882,N_8656,N_8701);
xnor U8883 (N_8883,N_8700,N_8731);
nand U8884 (N_8884,N_8758,N_8716);
xor U8885 (N_8885,N_8655,N_8787);
nor U8886 (N_8886,N_8796,N_8708);
nand U8887 (N_8887,N_8663,N_8771);
nand U8888 (N_8888,N_8737,N_8777);
xor U8889 (N_8889,N_8640,N_8735);
xor U8890 (N_8890,N_8679,N_8719);
or U8891 (N_8891,N_8792,N_8749);
nand U8892 (N_8892,N_8675,N_8709);
or U8893 (N_8893,N_8764,N_8694);
nor U8894 (N_8894,N_8720,N_8640);
xnor U8895 (N_8895,N_8702,N_8774);
nor U8896 (N_8896,N_8663,N_8653);
nor U8897 (N_8897,N_8687,N_8707);
and U8898 (N_8898,N_8663,N_8752);
or U8899 (N_8899,N_8728,N_8659);
xor U8900 (N_8900,N_8647,N_8727);
and U8901 (N_8901,N_8661,N_8751);
nand U8902 (N_8902,N_8697,N_8688);
nand U8903 (N_8903,N_8701,N_8677);
and U8904 (N_8904,N_8787,N_8679);
nor U8905 (N_8905,N_8699,N_8642);
or U8906 (N_8906,N_8680,N_8713);
or U8907 (N_8907,N_8665,N_8676);
nor U8908 (N_8908,N_8733,N_8694);
nor U8909 (N_8909,N_8666,N_8644);
or U8910 (N_8910,N_8746,N_8790);
nand U8911 (N_8911,N_8773,N_8726);
nand U8912 (N_8912,N_8770,N_8672);
and U8913 (N_8913,N_8699,N_8766);
nand U8914 (N_8914,N_8777,N_8669);
and U8915 (N_8915,N_8779,N_8718);
xor U8916 (N_8916,N_8760,N_8773);
nand U8917 (N_8917,N_8641,N_8707);
xnor U8918 (N_8918,N_8730,N_8698);
xor U8919 (N_8919,N_8748,N_8712);
nand U8920 (N_8920,N_8700,N_8709);
xor U8921 (N_8921,N_8672,N_8692);
or U8922 (N_8922,N_8761,N_8661);
and U8923 (N_8923,N_8714,N_8772);
xnor U8924 (N_8924,N_8715,N_8755);
nor U8925 (N_8925,N_8782,N_8699);
xor U8926 (N_8926,N_8779,N_8730);
or U8927 (N_8927,N_8664,N_8793);
nor U8928 (N_8928,N_8695,N_8795);
xor U8929 (N_8929,N_8711,N_8752);
nand U8930 (N_8930,N_8778,N_8791);
or U8931 (N_8931,N_8715,N_8651);
xor U8932 (N_8932,N_8745,N_8661);
nand U8933 (N_8933,N_8659,N_8737);
xor U8934 (N_8934,N_8684,N_8770);
nor U8935 (N_8935,N_8703,N_8728);
or U8936 (N_8936,N_8756,N_8710);
xnor U8937 (N_8937,N_8707,N_8661);
nand U8938 (N_8938,N_8756,N_8793);
xnor U8939 (N_8939,N_8731,N_8799);
nor U8940 (N_8940,N_8747,N_8757);
or U8941 (N_8941,N_8722,N_8693);
and U8942 (N_8942,N_8766,N_8701);
or U8943 (N_8943,N_8771,N_8662);
xnor U8944 (N_8944,N_8688,N_8721);
nor U8945 (N_8945,N_8784,N_8723);
or U8946 (N_8946,N_8786,N_8741);
and U8947 (N_8947,N_8744,N_8707);
or U8948 (N_8948,N_8744,N_8683);
xnor U8949 (N_8949,N_8677,N_8743);
nand U8950 (N_8950,N_8760,N_8706);
nor U8951 (N_8951,N_8745,N_8647);
nor U8952 (N_8952,N_8729,N_8783);
nor U8953 (N_8953,N_8784,N_8737);
or U8954 (N_8954,N_8691,N_8783);
nand U8955 (N_8955,N_8653,N_8718);
nand U8956 (N_8956,N_8768,N_8730);
nand U8957 (N_8957,N_8648,N_8786);
nor U8958 (N_8958,N_8724,N_8752);
nor U8959 (N_8959,N_8795,N_8664);
or U8960 (N_8960,N_8865,N_8958);
and U8961 (N_8961,N_8919,N_8935);
nand U8962 (N_8962,N_8916,N_8895);
or U8963 (N_8963,N_8898,N_8870);
nand U8964 (N_8964,N_8823,N_8806);
nor U8965 (N_8965,N_8856,N_8913);
or U8966 (N_8966,N_8908,N_8836);
nand U8967 (N_8967,N_8910,N_8938);
and U8968 (N_8968,N_8905,N_8860);
nor U8969 (N_8969,N_8940,N_8876);
xor U8970 (N_8970,N_8909,N_8899);
or U8971 (N_8971,N_8877,N_8821);
and U8972 (N_8972,N_8805,N_8944);
xor U8973 (N_8973,N_8888,N_8816);
xnor U8974 (N_8974,N_8803,N_8897);
nand U8975 (N_8975,N_8858,N_8901);
and U8976 (N_8976,N_8873,N_8955);
nor U8977 (N_8977,N_8952,N_8892);
or U8978 (N_8978,N_8937,N_8850);
or U8979 (N_8979,N_8894,N_8887);
or U8980 (N_8980,N_8884,N_8934);
or U8981 (N_8981,N_8866,N_8801);
or U8982 (N_8982,N_8815,N_8819);
or U8983 (N_8983,N_8959,N_8918);
or U8984 (N_8984,N_8904,N_8829);
nand U8985 (N_8985,N_8817,N_8811);
or U8986 (N_8986,N_8890,N_8878);
nor U8987 (N_8987,N_8893,N_8924);
nand U8988 (N_8988,N_8889,N_8822);
nand U8989 (N_8989,N_8868,N_8885);
nand U8990 (N_8990,N_8922,N_8840);
xnor U8991 (N_8991,N_8917,N_8953);
nand U8992 (N_8992,N_8925,N_8902);
nor U8993 (N_8993,N_8930,N_8863);
xnor U8994 (N_8994,N_8869,N_8948);
and U8995 (N_8995,N_8820,N_8891);
nand U8996 (N_8996,N_8914,N_8841);
xor U8997 (N_8997,N_8825,N_8861);
nor U8998 (N_8998,N_8882,N_8951);
and U8999 (N_8999,N_8871,N_8831);
xor U9000 (N_9000,N_8931,N_8929);
or U9001 (N_9001,N_8859,N_8883);
nor U9002 (N_9002,N_8879,N_8818);
nor U9003 (N_9003,N_8833,N_8954);
nand U9004 (N_9004,N_8941,N_8839);
nor U9005 (N_9005,N_8838,N_8851);
nand U9006 (N_9006,N_8843,N_8800);
and U9007 (N_9007,N_8881,N_8835);
nand U9008 (N_9008,N_8945,N_8923);
nor U9009 (N_9009,N_8903,N_8906);
and U9010 (N_9010,N_8864,N_8855);
nor U9011 (N_9011,N_8834,N_8804);
and U9012 (N_9012,N_8826,N_8915);
nand U9013 (N_9013,N_8857,N_8814);
and U9014 (N_9014,N_8847,N_8949);
or U9015 (N_9015,N_8900,N_8853);
or U9016 (N_9016,N_8867,N_8874);
nand U9017 (N_9017,N_8832,N_8880);
and U9018 (N_9018,N_8828,N_8946);
nor U9019 (N_9019,N_8926,N_8928);
and U9020 (N_9020,N_8842,N_8950);
nor U9021 (N_9021,N_8921,N_8808);
xor U9022 (N_9022,N_8852,N_8957);
nor U9023 (N_9023,N_8802,N_8848);
nand U9024 (N_9024,N_8896,N_8911);
xnor U9025 (N_9025,N_8845,N_8854);
nor U9026 (N_9026,N_8846,N_8813);
nand U9027 (N_9027,N_8943,N_8956);
nor U9028 (N_9028,N_8875,N_8809);
or U9029 (N_9029,N_8810,N_8807);
and U9030 (N_9030,N_8947,N_8862);
nor U9031 (N_9031,N_8942,N_8912);
or U9032 (N_9032,N_8812,N_8844);
xor U9033 (N_9033,N_8907,N_8920);
xnor U9034 (N_9034,N_8872,N_8837);
nor U9035 (N_9035,N_8932,N_8886);
nand U9036 (N_9036,N_8936,N_8827);
and U9037 (N_9037,N_8939,N_8830);
and U9038 (N_9038,N_8824,N_8849);
nand U9039 (N_9039,N_8927,N_8933);
or U9040 (N_9040,N_8923,N_8844);
xor U9041 (N_9041,N_8847,N_8895);
nor U9042 (N_9042,N_8856,N_8802);
xnor U9043 (N_9043,N_8906,N_8881);
and U9044 (N_9044,N_8885,N_8901);
xnor U9045 (N_9045,N_8825,N_8872);
and U9046 (N_9046,N_8860,N_8846);
and U9047 (N_9047,N_8946,N_8892);
nand U9048 (N_9048,N_8819,N_8870);
nand U9049 (N_9049,N_8955,N_8910);
or U9050 (N_9050,N_8880,N_8882);
and U9051 (N_9051,N_8823,N_8856);
nor U9052 (N_9052,N_8898,N_8822);
nor U9053 (N_9053,N_8831,N_8959);
nor U9054 (N_9054,N_8842,N_8870);
and U9055 (N_9055,N_8853,N_8922);
and U9056 (N_9056,N_8927,N_8956);
nand U9057 (N_9057,N_8846,N_8895);
or U9058 (N_9058,N_8824,N_8943);
and U9059 (N_9059,N_8849,N_8819);
xor U9060 (N_9060,N_8929,N_8895);
and U9061 (N_9061,N_8851,N_8952);
nand U9062 (N_9062,N_8906,N_8878);
and U9063 (N_9063,N_8927,N_8935);
or U9064 (N_9064,N_8939,N_8882);
nor U9065 (N_9065,N_8800,N_8930);
and U9066 (N_9066,N_8953,N_8830);
xnor U9067 (N_9067,N_8890,N_8959);
or U9068 (N_9068,N_8814,N_8820);
and U9069 (N_9069,N_8859,N_8868);
and U9070 (N_9070,N_8916,N_8801);
nor U9071 (N_9071,N_8835,N_8820);
and U9072 (N_9072,N_8956,N_8891);
xnor U9073 (N_9073,N_8870,N_8835);
or U9074 (N_9074,N_8906,N_8844);
nand U9075 (N_9075,N_8873,N_8878);
xnor U9076 (N_9076,N_8942,N_8827);
or U9077 (N_9077,N_8838,N_8921);
or U9078 (N_9078,N_8847,N_8800);
and U9079 (N_9079,N_8908,N_8804);
nand U9080 (N_9080,N_8883,N_8841);
and U9081 (N_9081,N_8822,N_8953);
nand U9082 (N_9082,N_8832,N_8869);
or U9083 (N_9083,N_8923,N_8818);
or U9084 (N_9084,N_8910,N_8909);
xor U9085 (N_9085,N_8896,N_8916);
nor U9086 (N_9086,N_8957,N_8823);
and U9087 (N_9087,N_8957,N_8855);
xor U9088 (N_9088,N_8867,N_8916);
nor U9089 (N_9089,N_8858,N_8862);
nand U9090 (N_9090,N_8915,N_8907);
or U9091 (N_9091,N_8916,N_8950);
and U9092 (N_9092,N_8920,N_8871);
xor U9093 (N_9093,N_8866,N_8918);
or U9094 (N_9094,N_8954,N_8810);
and U9095 (N_9095,N_8800,N_8879);
or U9096 (N_9096,N_8958,N_8922);
nand U9097 (N_9097,N_8896,N_8810);
xnor U9098 (N_9098,N_8847,N_8836);
nand U9099 (N_9099,N_8916,N_8805);
xor U9100 (N_9100,N_8936,N_8803);
or U9101 (N_9101,N_8915,N_8958);
xor U9102 (N_9102,N_8850,N_8846);
nand U9103 (N_9103,N_8932,N_8949);
xor U9104 (N_9104,N_8929,N_8860);
nand U9105 (N_9105,N_8835,N_8862);
xor U9106 (N_9106,N_8907,N_8812);
xnor U9107 (N_9107,N_8875,N_8825);
nor U9108 (N_9108,N_8807,N_8820);
nor U9109 (N_9109,N_8819,N_8951);
xor U9110 (N_9110,N_8931,N_8907);
nand U9111 (N_9111,N_8805,N_8894);
nand U9112 (N_9112,N_8873,N_8823);
nor U9113 (N_9113,N_8944,N_8902);
or U9114 (N_9114,N_8876,N_8816);
and U9115 (N_9115,N_8895,N_8828);
xor U9116 (N_9116,N_8832,N_8860);
and U9117 (N_9117,N_8959,N_8943);
nand U9118 (N_9118,N_8904,N_8861);
and U9119 (N_9119,N_8873,N_8917);
or U9120 (N_9120,N_8968,N_8976);
xnor U9121 (N_9121,N_9096,N_9002);
and U9122 (N_9122,N_9062,N_9110);
nand U9123 (N_9123,N_9033,N_8973);
nor U9124 (N_9124,N_9014,N_9049);
and U9125 (N_9125,N_8986,N_9080);
and U9126 (N_9126,N_9012,N_9113);
or U9127 (N_9127,N_9019,N_9007);
xnor U9128 (N_9128,N_8998,N_9044);
or U9129 (N_9129,N_9026,N_8960);
or U9130 (N_9130,N_8985,N_8978);
nand U9131 (N_9131,N_9087,N_9053);
xor U9132 (N_9132,N_9079,N_8980);
nand U9133 (N_9133,N_9003,N_8991);
nor U9134 (N_9134,N_9050,N_9058);
nor U9135 (N_9135,N_9061,N_9047);
or U9136 (N_9136,N_9051,N_9073);
nor U9137 (N_9137,N_8972,N_9095);
and U9138 (N_9138,N_9076,N_9032);
nor U9139 (N_9139,N_8962,N_9109);
and U9140 (N_9140,N_9038,N_9023);
or U9141 (N_9141,N_9066,N_9085);
xor U9142 (N_9142,N_9037,N_9052);
xor U9143 (N_9143,N_9000,N_8995);
and U9144 (N_9144,N_9048,N_9088);
nor U9145 (N_9145,N_8961,N_9015);
and U9146 (N_9146,N_9108,N_9041);
nor U9147 (N_9147,N_9024,N_9070);
xor U9148 (N_9148,N_9063,N_9101);
and U9149 (N_9149,N_9068,N_9029);
and U9150 (N_9150,N_9078,N_8993);
and U9151 (N_9151,N_8975,N_9081);
and U9152 (N_9152,N_9083,N_8990);
or U9153 (N_9153,N_9105,N_8984);
or U9154 (N_9154,N_9084,N_8964);
or U9155 (N_9155,N_9069,N_9055);
xnor U9156 (N_9156,N_9042,N_9056);
or U9157 (N_9157,N_9018,N_9008);
and U9158 (N_9158,N_9090,N_9030);
and U9159 (N_9159,N_8979,N_9111);
and U9160 (N_9160,N_9013,N_9021);
xor U9161 (N_9161,N_9020,N_9004);
and U9162 (N_9162,N_9065,N_9001);
xnor U9163 (N_9163,N_9025,N_9075);
xor U9164 (N_9164,N_9107,N_9009);
nor U9165 (N_9165,N_8965,N_9022);
or U9166 (N_9166,N_9010,N_9031);
xor U9167 (N_9167,N_9064,N_8971);
or U9168 (N_9168,N_9006,N_9027);
xor U9169 (N_9169,N_9005,N_9039);
or U9170 (N_9170,N_8981,N_8966);
or U9171 (N_9171,N_8983,N_9086);
and U9172 (N_9172,N_9082,N_9092);
xor U9173 (N_9173,N_8967,N_9103);
and U9174 (N_9174,N_9071,N_9060);
nor U9175 (N_9175,N_9040,N_9112);
nand U9176 (N_9176,N_8996,N_9045);
xnor U9177 (N_9177,N_9119,N_8970);
xnor U9178 (N_9178,N_9102,N_9097);
nor U9179 (N_9179,N_8994,N_9116);
and U9180 (N_9180,N_9059,N_9118);
or U9181 (N_9181,N_9094,N_9077);
and U9182 (N_9182,N_9054,N_9057);
and U9183 (N_9183,N_9117,N_8969);
and U9184 (N_9184,N_8974,N_9046);
and U9185 (N_9185,N_9074,N_9034);
nor U9186 (N_9186,N_9028,N_9035);
or U9187 (N_9187,N_9011,N_9072);
nor U9188 (N_9188,N_9100,N_8997);
nand U9189 (N_9189,N_9016,N_9099);
nor U9190 (N_9190,N_9098,N_9043);
and U9191 (N_9191,N_8999,N_9067);
or U9192 (N_9192,N_8977,N_9106);
and U9193 (N_9193,N_9017,N_8987);
and U9194 (N_9194,N_9114,N_8982);
nand U9195 (N_9195,N_9115,N_8992);
or U9196 (N_9196,N_9036,N_9093);
nand U9197 (N_9197,N_8989,N_8988);
nor U9198 (N_9198,N_9089,N_8963);
xnor U9199 (N_9199,N_9104,N_9091);
nand U9200 (N_9200,N_9088,N_9056);
nor U9201 (N_9201,N_8961,N_9009);
nor U9202 (N_9202,N_9096,N_9064);
and U9203 (N_9203,N_9111,N_8990);
xor U9204 (N_9204,N_9016,N_9046);
or U9205 (N_9205,N_8997,N_8983);
and U9206 (N_9206,N_9119,N_8999);
or U9207 (N_9207,N_9074,N_9058);
or U9208 (N_9208,N_9044,N_9020);
and U9209 (N_9209,N_9025,N_9097);
nor U9210 (N_9210,N_9057,N_8984);
nand U9211 (N_9211,N_8965,N_9090);
nor U9212 (N_9212,N_9052,N_9059);
or U9213 (N_9213,N_9076,N_9054);
and U9214 (N_9214,N_8981,N_9009);
and U9215 (N_9215,N_9117,N_9048);
nor U9216 (N_9216,N_8971,N_8993);
xnor U9217 (N_9217,N_8990,N_8981);
xnor U9218 (N_9218,N_9002,N_9111);
or U9219 (N_9219,N_9105,N_9022);
nand U9220 (N_9220,N_8994,N_8981);
or U9221 (N_9221,N_9059,N_8977);
xnor U9222 (N_9222,N_9028,N_9077);
or U9223 (N_9223,N_9094,N_9060);
and U9224 (N_9224,N_9053,N_9031);
or U9225 (N_9225,N_9026,N_9105);
xnor U9226 (N_9226,N_9079,N_9048);
xor U9227 (N_9227,N_9098,N_9076);
or U9228 (N_9228,N_9088,N_9098);
nor U9229 (N_9229,N_8964,N_9054);
or U9230 (N_9230,N_9045,N_8986);
and U9231 (N_9231,N_9052,N_9062);
nand U9232 (N_9232,N_9075,N_9066);
and U9233 (N_9233,N_9021,N_9037);
and U9234 (N_9234,N_9080,N_9093);
xnor U9235 (N_9235,N_9109,N_9094);
nand U9236 (N_9236,N_8999,N_8962);
nor U9237 (N_9237,N_8960,N_9057);
xor U9238 (N_9238,N_9093,N_8978);
or U9239 (N_9239,N_9009,N_9058);
nand U9240 (N_9240,N_9091,N_9030);
or U9241 (N_9241,N_9011,N_9055);
nand U9242 (N_9242,N_9027,N_8993);
or U9243 (N_9243,N_9061,N_8967);
nand U9244 (N_9244,N_9012,N_8989);
nor U9245 (N_9245,N_8996,N_9087);
xor U9246 (N_9246,N_9087,N_9069);
and U9247 (N_9247,N_9001,N_9112);
xnor U9248 (N_9248,N_9026,N_9055);
nand U9249 (N_9249,N_9028,N_9031);
nor U9250 (N_9250,N_9113,N_9021);
nand U9251 (N_9251,N_9011,N_8968);
and U9252 (N_9252,N_9030,N_8980);
nand U9253 (N_9253,N_9081,N_8964);
and U9254 (N_9254,N_9070,N_8972);
and U9255 (N_9255,N_9000,N_9064);
nor U9256 (N_9256,N_9022,N_9017);
or U9257 (N_9257,N_9029,N_9031);
or U9258 (N_9258,N_9064,N_9072);
nor U9259 (N_9259,N_9036,N_9027);
xnor U9260 (N_9260,N_8991,N_9068);
nand U9261 (N_9261,N_9085,N_9007);
or U9262 (N_9262,N_9021,N_8988);
and U9263 (N_9263,N_9053,N_9011);
nand U9264 (N_9264,N_9078,N_8986);
xor U9265 (N_9265,N_9087,N_8990);
and U9266 (N_9266,N_9026,N_9078);
nor U9267 (N_9267,N_9095,N_9002);
nand U9268 (N_9268,N_9090,N_9117);
nor U9269 (N_9269,N_8995,N_9050);
nor U9270 (N_9270,N_9078,N_9090);
xor U9271 (N_9271,N_9070,N_9028);
xnor U9272 (N_9272,N_9020,N_9073);
xnor U9273 (N_9273,N_9113,N_9028);
and U9274 (N_9274,N_9093,N_9050);
or U9275 (N_9275,N_9067,N_9033);
xor U9276 (N_9276,N_9050,N_8991);
nor U9277 (N_9277,N_9084,N_9039);
nand U9278 (N_9278,N_9087,N_9044);
nand U9279 (N_9279,N_9007,N_9101);
nand U9280 (N_9280,N_9127,N_9214);
nand U9281 (N_9281,N_9265,N_9142);
nand U9282 (N_9282,N_9249,N_9257);
nor U9283 (N_9283,N_9217,N_9206);
or U9284 (N_9284,N_9186,N_9145);
nand U9285 (N_9285,N_9176,N_9163);
and U9286 (N_9286,N_9233,N_9129);
and U9287 (N_9287,N_9250,N_9261);
or U9288 (N_9288,N_9192,N_9134);
or U9289 (N_9289,N_9224,N_9133);
nand U9290 (N_9290,N_9137,N_9157);
nor U9291 (N_9291,N_9221,N_9264);
and U9292 (N_9292,N_9126,N_9174);
or U9293 (N_9293,N_9246,N_9204);
nor U9294 (N_9294,N_9228,N_9179);
nor U9295 (N_9295,N_9160,N_9189);
and U9296 (N_9296,N_9207,N_9259);
xnor U9297 (N_9297,N_9242,N_9254);
nor U9298 (N_9298,N_9121,N_9251);
and U9299 (N_9299,N_9212,N_9165);
nand U9300 (N_9300,N_9123,N_9234);
or U9301 (N_9301,N_9152,N_9122);
nor U9302 (N_9302,N_9182,N_9267);
or U9303 (N_9303,N_9181,N_9146);
xnor U9304 (N_9304,N_9230,N_9268);
nand U9305 (N_9305,N_9138,N_9240);
and U9306 (N_9306,N_9244,N_9200);
nand U9307 (N_9307,N_9271,N_9135);
xor U9308 (N_9308,N_9252,N_9247);
and U9309 (N_9309,N_9219,N_9180);
nand U9310 (N_9310,N_9202,N_9213);
nand U9311 (N_9311,N_9172,N_9203);
nand U9312 (N_9312,N_9232,N_9153);
nor U9313 (N_9313,N_9236,N_9222);
and U9314 (N_9314,N_9270,N_9173);
and U9315 (N_9315,N_9253,N_9258);
xnor U9316 (N_9316,N_9159,N_9272);
and U9317 (N_9317,N_9161,N_9274);
nor U9318 (N_9318,N_9156,N_9149);
nor U9319 (N_9319,N_9162,N_9166);
and U9320 (N_9320,N_9266,N_9144);
nand U9321 (N_9321,N_9185,N_9194);
xnor U9322 (N_9322,N_9276,N_9255);
nor U9323 (N_9323,N_9170,N_9210);
xnor U9324 (N_9324,N_9130,N_9208);
nand U9325 (N_9325,N_9154,N_9169);
and U9326 (N_9326,N_9241,N_9226);
and U9327 (N_9327,N_9239,N_9275);
xor U9328 (N_9328,N_9196,N_9177);
nand U9329 (N_9329,N_9231,N_9248);
or U9330 (N_9330,N_9273,N_9225);
or U9331 (N_9331,N_9164,N_9140);
and U9332 (N_9332,N_9256,N_9215);
nand U9333 (N_9333,N_9120,N_9269);
and U9334 (N_9334,N_9262,N_9143);
or U9335 (N_9335,N_9218,N_9197);
xor U9336 (N_9336,N_9277,N_9199);
nor U9337 (N_9337,N_9216,N_9227);
nor U9338 (N_9338,N_9279,N_9175);
nand U9339 (N_9339,N_9209,N_9198);
or U9340 (N_9340,N_9168,N_9223);
nor U9341 (N_9341,N_9183,N_9167);
nand U9342 (N_9342,N_9171,N_9151);
xor U9343 (N_9343,N_9190,N_9155);
or U9344 (N_9344,N_9278,N_9245);
or U9345 (N_9345,N_9188,N_9237);
nand U9346 (N_9346,N_9220,N_9132);
xor U9347 (N_9347,N_9184,N_9263);
and U9348 (N_9348,N_9131,N_9147);
xor U9349 (N_9349,N_9139,N_9187);
xor U9350 (N_9350,N_9243,N_9124);
or U9351 (N_9351,N_9235,N_9229);
xnor U9352 (N_9352,N_9205,N_9125);
nor U9353 (N_9353,N_9260,N_9148);
nand U9354 (N_9354,N_9158,N_9150);
or U9355 (N_9355,N_9136,N_9201);
xnor U9356 (N_9356,N_9191,N_9193);
and U9357 (N_9357,N_9128,N_9178);
nand U9358 (N_9358,N_9195,N_9141);
or U9359 (N_9359,N_9238,N_9211);
nand U9360 (N_9360,N_9209,N_9217);
xor U9361 (N_9361,N_9190,N_9200);
or U9362 (N_9362,N_9167,N_9141);
nor U9363 (N_9363,N_9223,N_9131);
nand U9364 (N_9364,N_9150,N_9123);
xor U9365 (N_9365,N_9239,N_9135);
xor U9366 (N_9366,N_9264,N_9216);
xnor U9367 (N_9367,N_9267,N_9254);
nand U9368 (N_9368,N_9263,N_9244);
and U9369 (N_9369,N_9140,N_9194);
nand U9370 (N_9370,N_9259,N_9241);
xnor U9371 (N_9371,N_9277,N_9271);
and U9372 (N_9372,N_9241,N_9129);
nor U9373 (N_9373,N_9165,N_9136);
nor U9374 (N_9374,N_9146,N_9209);
nor U9375 (N_9375,N_9209,N_9274);
xnor U9376 (N_9376,N_9223,N_9220);
nand U9377 (N_9377,N_9184,N_9235);
nand U9378 (N_9378,N_9218,N_9154);
nand U9379 (N_9379,N_9234,N_9265);
nor U9380 (N_9380,N_9224,N_9275);
nor U9381 (N_9381,N_9154,N_9258);
and U9382 (N_9382,N_9275,N_9122);
nand U9383 (N_9383,N_9170,N_9233);
xnor U9384 (N_9384,N_9229,N_9176);
and U9385 (N_9385,N_9250,N_9227);
and U9386 (N_9386,N_9279,N_9240);
nand U9387 (N_9387,N_9275,N_9166);
nand U9388 (N_9388,N_9144,N_9218);
nand U9389 (N_9389,N_9260,N_9195);
or U9390 (N_9390,N_9230,N_9277);
nor U9391 (N_9391,N_9277,N_9210);
xnor U9392 (N_9392,N_9217,N_9139);
or U9393 (N_9393,N_9137,N_9183);
or U9394 (N_9394,N_9202,N_9215);
nand U9395 (N_9395,N_9129,N_9251);
xor U9396 (N_9396,N_9248,N_9129);
and U9397 (N_9397,N_9228,N_9241);
nor U9398 (N_9398,N_9161,N_9158);
xnor U9399 (N_9399,N_9168,N_9145);
xnor U9400 (N_9400,N_9126,N_9224);
and U9401 (N_9401,N_9129,N_9126);
or U9402 (N_9402,N_9202,N_9237);
xnor U9403 (N_9403,N_9207,N_9221);
xor U9404 (N_9404,N_9184,N_9157);
nor U9405 (N_9405,N_9237,N_9145);
and U9406 (N_9406,N_9147,N_9278);
and U9407 (N_9407,N_9166,N_9182);
xor U9408 (N_9408,N_9186,N_9170);
nor U9409 (N_9409,N_9148,N_9139);
nand U9410 (N_9410,N_9279,N_9163);
and U9411 (N_9411,N_9246,N_9203);
nor U9412 (N_9412,N_9165,N_9259);
xor U9413 (N_9413,N_9251,N_9255);
xnor U9414 (N_9414,N_9125,N_9132);
or U9415 (N_9415,N_9159,N_9261);
nand U9416 (N_9416,N_9174,N_9226);
or U9417 (N_9417,N_9270,N_9177);
or U9418 (N_9418,N_9139,N_9252);
nand U9419 (N_9419,N_9214,N_9209);
or U9420 (N_9420,N_9257,N_9130);
and U9421 (N_9421,N_9136,N_9198);
and U9422 (N_9422,N_9193,N_9259);
or U9423 (N_9423,N_9155,N_9127);
nand U9424 (N_9424,N_9142,N_9174);
and U9425 (N_9425,N_9170,N_9218);
nor U9426 (N_9426,N_9139,N_9172);
nand U9427 (N_9427,N_9157,N_9231);
xnor U9428 (N_9428,N_9122,N_9172);
and U9429 (N_9429,N_9139,N_9268);
nand U9430 (N_9430,N_9235,N_9171);
and U9431 (N_9431,N_9209,N_9145);
xor U9432 (N_9432,N_9183,N_9136);
nand U9433 (N_9433,N_9247,N_9185);
nand U9434 (N_9434,N_9215,N_9174);
xor U9435 (N_9435,N_9273,N_9226);
or U9436 (N_9436,N_9234,N_9218);
xnor U9437 (N_9437,N_9270,N_9184);
and U9438 (N_9438,N_9128,N_9197);
nor U9439 (N_9439,N_9268,N_9136);
or U9440 (N_9440,N_9430,N_9353);
xor U9441 (N_9441,N_9387,N_9282);
or U9442 (N_9442,N_9309,N_9372);
xnor U9443 (N_9443,N_9301,N_9349);
xnor U9444 (N_9444,N_9423,N_9390);
nor U9445 (N_9445,N_9287,N_9429);
and U9446 (N_9446,N_9437,N_9391);
and U9447 (N_9447,N_9347,N_9362);
and U9448 (N_9448,N_9280,N_9324);
nor U9449 (N_9449,N_9389,N_9428);
xnor U9450 (N_9450,N_9299,N_9402);
nor U9451 (N_9451,N_9361,N_9438);
nor U9452 (N_9452,N_9295,N_9424);
nor U9453 (N_9453,N_9293,N_9407);
and U9454 (N_9454,N_9298,N_9406);
nand U9455 (N_9455,N_9416,N_9393);
xnor U9456 (N_9456,N_9392,N_9399);
nor U9457 (N_9457,N_9421,N_9436);
and U9458 (N_9458,N_9415,N_9404);
or U9459 (N_9459,N_9316,N_9281);
xor U9460 (N_9460,N_9386,N_9371);
nand U9461 (N_9461,N_9286,N_9369);
or U9462 (N_9462,N_9370,N_9354);
and U9463 (N_9463,N_9408,N_9377);
nand U9464 (N_9464,N_9373,N_9289);
and U9465 (N_9465,N_9419,N_9325);
xor U9466 (N_9466,N_9306,N_9337);
nand U9467 (N_9467,N_9374,N_9314);
nand U9468 (N_9468,N_9384,N_9396);
nand U9469 (N_9469,N_9300,N_9338);
xnor U9470 (N_9470,N_9379,N_9405);
or U9471 (N_9471,N_9398,N_9303);
and U9472 (N_9472,N_9360,N_9395);
nand U9473 (N_9473,N_9291,N_9422);
nor U9474 (N_9474,N_9336,N_9313);
nor U9475 (N_9475,N_9315,N_9427);
or U9476 (N_9476,N_9317,N_9412);
and U9477 (N_9477,N_9311,N_9323);
and U9478 (N_9478,N_9350,N_9388);
and U9479 (N_9479,N_9426,N_9285);
nand U9480 (N_9480,N_9439,N_9366);
nand U9481 (N_9481,N_9345,N_9294);
and U9482 (N_9482,N_9290,N_9292);
and U9483 (N_9483,N_9340,N_9328);
nand U9484 (N_9484,N_9381,N_9380);
nand U9485 (N_9485,N_9341,N_9378);
and U9486 (N_9486,N_9401,N_9376);
and U9487 (N_9487,N_9433,N_9319);
nand U9488 (N_9488,N_9308,N_9358);
or U9489 (N_9489,N_9339,N_9357);
nor U9490 (N_9490,N_9320,N_9326);
or U9491 (N_9491,N_9356,N_9321);
xor U9492 (N_9492,N_9283,N_9296);
nor U9493 (N_9493,N_9312,N_9332);
xnor U9494 (N_9494,N_9383,N_9409);
nor U9495 (N_9495,N_9431,N_9327);
xor U9496 (N_9496,N_9432,N_9331);
nor U9497 (N_9497,N_9322,N_9288);
xnor U9498 (N_9498,N_9403,N_9434);
xor U9499 (N_9499,N_9397,N_9368);
and U9500 (N_9500,N_9304,N_9363);
nor U9501 (N_9501,N_9330,N_9413);
xnor U9502 (N_9502,N_9318,N_9346);
xor U9503 (N_9503,N_9410,N_9355);
nand U9504 (N_9504,N_9375,N_9342);
and U9505 (N_9505,N_9364,N_9348);
nor U9506 (N_9506,N_9302,N_9333);
or U9507 (N_9507,N_9400,N_9411);
and U9508 (N_9508,N_9310,N_9385);
nand U9509 (N_9509,N_9365,N_9307);
nor U9510 (N_9510,N_9329,N_9367);
and U9511 (N_9511,N_9382,N_9344);
and U9512 (N_9512,N_9417,N_9420);
nand U9513 (N_9513,N_9334,N_9284);
nor U9514 (N_9514,N_9418,N_9425);
or U9515 (N_9515,N_9305,N_9414);
nor U9516 (N_9516,N_9343,N_9394);
nand U9517 (N_9517,N_9335,N_9351);
nand U9518 (N_9518,N_9435,N_9297);
nand U9519 (N_9519,N_9359,N_9352);
nand U9520 (N_9520,N_9292,N_9351);
nor U9521 (N_9521,N_9423,N_9429);
nor U9522 (N_9522,N_9327,N_9305);
xnor U9523 (N_9523,N_9384,N_9427);
nor U9524 (N_9524,N_9315,N_9429);
or U9525 (N_9525,N_9414,N_9284);
nor U9526 (N_9526,N_9297,N_9307);
nor U9527 (N_9527,N_9351,N_9401);
xnor U9528 (N_9528,N_9425,N_9422);
nor U9529 (N_9529,N_9365,N_9331);
nand U9530 (N_9530,N_9367,N_9282);
or U9531 (N_9531,N_9360,N_9340);
nor U9532 (N_9532,N_9392,N_9292);
and U9533 (N_9533,N_9350,N_9345);
xor U9534 (N_9534,N_9322,N_9326);
nor U9535 (N_9535,N_9377,N_9420);
xor U9536 (N_9536,N_9435,N_9319);
nand U9537 (N_9537,N_9434,N_9369);
xnor U9538 (N_9538,N_9420,N_9354);
nor U9539 (N_9539,N_9433,N_9357);
xnor U9540 (N_9540,N_9439,N_9329);
nor U9541 (N_9541,N_9323,N_9291);
and U9542 (N_9542,N_9351,N_9372);
nor U9543 (N_9543,N_9345,N_9411);
nand U9544 (N_9544,N_9427,N_9300);
or U9545 (N_9545,N_9350,N_9370);
nand U9546 (N_9546,N_9374,N_9293);
and U9547 (N_9547,N_9360,N_9324);
and U9548 (N_9548,N_9313,N_9416);
xnor U9549 (N_9549,N_9324,N_9330);
nand U9550 (N_9550,N_9370,N_9306);
nand U9551 (N_9551,N_9304,N_9302);
or U9552 (N_9552,N_9335,N_9401);
xor U9553 (N_9553,N_9386,N_9429);
and U9554 (N_9554,N_9297,N_9387);
xnor U9555 (N_9555,N_9349,N_9297);
nand U9556 (N_9556,N_9398,N_9292);
nand U9557 (N_9557,N_9397,N_9375);
and U9558 (N_9558,N_9325,N_9324);
and U9559 (N_9559,N_9344,N_9374);
or U9560 (N_9560,N_9404,N_9394);
or U9561 (N_9561,N_9430,N_9434);
or U9562 (N_9562,N_9341,N_9385);
xnor U9563 (N_9563,N_9330,N_9335);
nor U9564 (N_9564,N_9365,N_9410);
nor U9565 (N_9565,N_9294,N_9364);
and U9566 (N_9566,N_9363,N_9439);
nor U9567 (N_9567,N_9353,N_9355);
nand U9568 (N_9568,N_9405,N_9371);
xor U9569 (N_9569,N_9281,N_9372);
nand U9570 (N_9570,N_9425,N_9284);
and U9571 (N_9571,N_9401,N_9365);
nand U9572 (N_9572,N_9378,N_9413);
nand U9573 (N_9573,N_9301,N_9295);
xor U9574 (N_9574,N_9316,N_9307);
and U9575 (N_9575,N_9293,N_9358);
nor U9576 (N_9576,N_9411,N_9282);
xnor U9577 (N_9577,N_9413,N_9307);
nand U9578 (N_9578,N_9422,N_9293);
xnor U9579 (N_9579,N_9397,N_9417);
nor U9580 (N_9580,N_9417,N_9387);
nand U9581 (N_9581,N_9394,N_9400);
xnor U9582 (N_9582,N_9351,N_9323);
nor U9583 (N_9583,N_9347,N_9283);
or U9584 (N_9584,N_9334,N_9354);
nand U9585 (N_9585,N_9376,N_9351);
and U9586 (N_9586,N_9338,N_9343);
or U9587 (N_9587,N_9398,N_9411);
nand U9588 (N_9588,N_9305,N_9328);
or U9589 (N_9589,N_9370,N_9325);
nand U9590 (N_9590,N_9285,N_9401);
and U9591 (N_9591,N_9360,N_9315);
nand U9592 (N_9592,N_9331,N_9286);
xnor U9593 (N_9593,N_9379,N_9319);
nand U9594 (N_9594,N_9282,N_9376);
nor U9595 (N_9595,N_9284,N_9306);
and U9596 (N_9596,N_9411,N_9341);
nor U9597 (N_9597,N_9406,N_9315);
and U9598 (N_9598,N_9304,N_9404);
or U9599 (N_9599,N_9363,N_9425);
xor U9600 (N_9600,N_9474,N_9517);
and U9601 (N_9601,N_9563,N_9461);
or U9602 (N_9602,N_9587,N_9488);
xnor U9603 (N_9603,N_9594,N_9486);
or U9604 (N_9604,N_9519,N_9545);
nor U9605 (N_9605,N_9525,N_9485);
or U9606 (N_9606,N_9515,N_9458);
or U9607 (N_9607,N_9521,N_9503);
nor U9608 (N_9608,N_9459,N_9523);
or U9609 (N_9609,N_9505,N_9552);
and U9610 (N_9610,N_9547,N_9504);
or U9611 (N_9611,N_9445,N_9443);
or U9612 (N_9612,N_9534,N_9506);
nand U9613 (N_9613,N_9453,N_9558);
nor U9614 (N_9614,N_9524,N_9583);
nand U9615 (N_9615,N_9507,N_9568);
or U9616 (N_9616,N_9489,N_9480);
nor U9617 (N_9617,N_9527,N_9448);
or U9618 (N_9618,N_9564,N_9472);
xor U9619 (N_9619,N_9441,N_9473);
or U9620 (N_9620,N_9593,N_9455);
nor U9621 (N_9621,N_9582,N_9497);
or U9622 (N_9622,N_9578,N_9496);
or U9623 (N_9623,N_9493,N_9541);
xnor U9624 (N_9624,N_9508,N_9562);
xor U9625 (N_9625,N_9444,N_9491);
xor U9626 (N_9626,N_9509,N_9586);
and U9627 (N_9627,N_9535,N_9451);
xor U9628 (N_9628,N_9464,N_9442);
nand U9629 (N_9629,N_9581,N_9516);
xnor U9630 (N_9630,N_9574,N_9567);
nand U9631 (N_9631,N_9554,N_9598);
and U9632 (N_9632,N_9501,N_9560);
nand U9633 (N_9633,N_9469,N_9579);
or U9634 (N_9634,N_9476,N_9589);
nand U9635 (N_9635,N_9475,N_9452);
nand U9636 (N_9636,N_9573,N_9457);
or U9637 (N_9637,N_9576,N_9546);
nand U9638 (N_9638,N_9571,N_9447);
nor U9639 (N_9639,N_9553,N_9518);
and U9640 (N_9640,N_9440,N_9595);
nand U9641 (N_9641,N_9572,N_9483);
nor U9642 (N_9642,N_9561,N_9536);
nand U9643 (N_9643,N_9533,N_9592);
xnor U9644 (N_9644,N_9477,N_9514);
or U9645 (N_9645,N_9544,N_9492);
xor U9646 (N_9646,N_9449,N_9511);
and U9647 (N_9647,N_9467,N_9502);
nand U9648 (N_9648,N_9454,N_9538);
xnor U9649 (N_9649,N_9470,N_9487);
or U9650 (N_9650,N_9550,N_9466);
nand U9651 (N_9651,N_9494,N_9481);
or U9652 (N_9652,N_9512,N_9450);
nor U9653 (N_9653,N_9498,N_9597);
or U9654 (N_9654,N_9528,N_9542);
or U9655 (N_9655,N_9468,N_9462);
nand U9656 (N_9656,N_9482,N_9537);
or U9657 (N_9657,N_9590,N_9577);
and U9658 (N_9658,N_9529,N_9549);
nand U9659 (N_9659,N_9490,N_9570);
nor U9660 (N_9660,N_9484,N_9556);
and U9661 (N_9661,N_9599,N_9565);
or U9662 (N_9662,N_9551,N_9584);
nor U9663 (N_9663,N_9569,N_9463);
nor U9664 (N_9664,N_9566,N_9539);
nand U9665 (N_9665,N_9540,N_9532);
and U9666 (N_9666,N_9591,N_9500);
nand U9667 (N_9667,N_9555,N_9479);
xor U9668 (N_9668,N_9522,N_9531);
xor U9669 (N_9669,N_9460,N_9580);
and U9670 (N_9670,N_9513,N_9575);
nand U9671 (N_9671,N_9526,N_9530);
nand U9672 (N_9672,N_9520,N_9557);
nand U9673 (N_9673,N_9471,N_9588);
or U9674 (N_9674,N_9499,N_9596);
and U9675 (N_9675,N_9465,N_9456);
xor U9676 (N_9676,N_9548,N_9510);
and U9677 (N_9677,N_9543,N_9478);
and U9678 (N_9678,N_9585,N_9495);
xor U9679 (N_9679,N_9446,N_9559);
and U9680 (N_9680,N_9586,N_9445);
and U9681 (N_9681,N_9465,N_9447);
nor U9682 (N_9682,N_9545,N_9588);
and U9683 (N_9683,N_9468,N_9553);
nand U9684 (N_9684,N_9563,N_9590);
nand U9685 (N_9685,N_9505,N_9521);
and U9686 (N_9686,N_9460,N_9561);
nand U9687 (N_9687,N_9480,N_9455);
nand U9688 (N_9688,N_9519,N_9510);
nand U9689 (N_9689,N_9473,N_9507);
nor U9690 (N_9690,N_9577,N_9582);
nor U9691 (N_9691,N_9556,N_9521);
xor U9692 (N_9692,N_9518,N_9575);
xor U9693 (N_9693,N_9463,N_9512);
nor U9694 (N_9694,N_9565,N_9537);
or U9695 (N_9695,N_9586,N_9522);
and U9696 (N_9696,N_9585,N_9497);
and U9697 (N_9697,N_9492,N_9532);
nor U9698 (N_9698,N_9457,N_9540);
nand U9699 (N_9699,N_9507,N_9573);
xnor U9700 (N_9700,N_9589,N_9537);
and U9701 (N_9701,N_9565,N_9470);
xor U9702 (N_9702,N_9550,N_9441);
nor U9703 (N_9703,N_9452,N_9493);
nand U9704 (N_9704,N_9569,N_9521);
nand U9705 (N_9705,N_9568,N_9578);
nand U9706 (N_9706,N_9565,N_9484);
nor U9707 (N_9707,N_9492,N_9450);
or U9708 (N_9708,N_9479,N_9475);
nor U9709 (N_9709,N_9444,N_9587);
nand U9710 (N_9710,N_9570,N_9498);
xor U9711 (N_9711,N_9588,N_9585);
or U9712 (N_9712,N_9471,N_9510);
or U9713 (N_9713,N_9556,N_9594);
or U9714 (N_9714,N_9576,N_9516);
or U9715 (N_9715,N_9588,N_9568);
nor U9716 (N_9716,N_9446,N_9491);
nand U9717 (N_9717,N_9484,N_9479);
or U9718 (N_9718,N_9595,N_9497);
nor U9719 (N_9719,N_9477,N_9451);
and U9720 (N_9720,N_9442,N_9496);
and U9721 (N_9721,N_9542,N_9447);
and U9722 (N_9722,N_9597,N_9476);
xor U9723 (N_9723,N_9552,N_9470);
and U9724 (N_9724,N_9479,N_9511);
or U9725 (N_9725,N_9501,N_9599);
or U9726 (N_9726,N_9593,N_9506);
xnor U9727 (N_9727,N_9444,N_9597);
nand U9728 (N_9728,N_9452,N_9504);
xnor U9729 (N_9729,N_9578,N_9536);
nand U9730 (N_9730,N_9535,N_9452);
and U9731 (N_9731,N_9479,N_9581);
and U9732 (N_9732,N_9495,N_9447);
nor U9733 (N_9733,N_9534,N_9579);
or U9734 (N_9734,N_9544,N_9518);
or U9735 (N_9735,N_9510,N_9494);
nor U9736 (N_9736,N_9584,N_9550);
or U9737 (N_9737,N_9539,N_9568);
and U9738 (N_9738,N_9458,N_9517);
and U9739 (N_9739,N_9563,N_9572);
xor U9740 (N_9740,N_9474,N_9522);
and U9741 (N_9741,N_9576,N_9455);
nand U9742 (N_9742,N_9556,N_9462);
nand U9743 (N_9743,N_9471,N_9445);
or U9744 (N_9744,N_9556,N_9548);
nor U9745 (N_9745,N_9488,N_9474);
and U9746 (N_9746,N_9465,N_9471);
and U9747 (N_9747,N_9498,N_9511);
xor U9748 (N_9748,N_9593,N_9558);
and U9749 (N_9749,N_9534,N_9501);
xnor U9750 (N_9750,N_9450,N_9452);
xnor U9751 (N_9751,N_9444,N_9594);
nor U9752 (N_9752,N_9469,N_9538);
and U9753 (N_9753,N_9582,N_9517);
and U9754 (N_9754,N_9494,N_9469);
nand U9755 (N_9755,N_9590,N_9519);
nor U9756 (N_9756,N_9544,N_9534);
nor U9757 (N_9757,N_9442,N_9484);
xor U9758 (N_9758,N_9596,N_9487);
and U9759 (N_9759,N_9525,N_9550);
xor U9760 (N_9760,N_9662,N_9704);
nand U9761 (N_9761,N_9618,N_9623);
nor U9762 (N_9762,N_9738,N_9735);
nor U9763 (N_9763,N_9644,N_9753);
xor U9764 (N_9764,N_9732,N_9654);
xor U9765 (N_9765,N_9620,N_9628);
or U9766 (N_9766,N_9667,N_9663);
nor U9767 (N_9767,N_9734,N_9683);
xnor U9768 (N_9768,N_9702,N_9710);
nand U9769 (N_9769,N_9679,N_9682);
nor U9770 (N_9770,N_9649,N_9657);
and U9771 (N_9771,N_9638,N_9627);
nand U9772 (N_9772,N_9680,N_9757);
or U9773 (N_9773,N_9720,N_9642);
and U9774 (N_9774,N_9717,N_9645);
or U9775 (N_9775,N_9725,N_9748);
and U9776 (N_9776,N_9668,N_9664);
nor U9777 (N_9777,N_9676,N_9700);
nand U9778 (N_9778,N_9606,N_9711);
xor U9779 (N_9779,N_9721,N_9724);
nand U9780 (N_9780,N_9705,N_9731);
xnor U9781 (N_9781,N_9636,N_9646);
and U9782 (N_9782,N_9707,N_9625);
nand U9783 (N_9783,N_9730,N_9743);
xnor U9784 (N_9784,N_9714,N_9626);
nor U9785 (N_9785,N_9703,N_9684);
or U9786 (N_9786,N_9696,N_9741);
nand U9787 (N_9787,N_9602,N_9733);
xnor U9788 (N_9788,N_9652,N_9675);
or U9789 (N_9789,N_9617,N_9712);
and U9790 (N_9790,N_9665,N_9744);
nand U9791 (N_9791,N_9648,N_9759);
xnor U9792 (N_9792,N_9672,N_9630);
nand U9793 (N_9793,N_9637,N_9656);
and U9794 (N_9794,N_9699,N_9752);
xor U9795 (N_9795,N_9698,N_9653);
and U9796 (N_9796,N_9661,N_9677);
nor U9797 (N_9797,N_9692,N_9709);
and U9798 (N_9798,N_9633,N_9600);
and U9799 (N_9799,N_9697,N_9659);
and U9800 (N_9800,N_9673,N_9723);
nor U9801 (N_9801,N_9681,N_9650);
nand U9802 (N_9802,N_9695,N_9634);
nor U9803 (N_9803,N_9736,N_9693);
nor U9804 (N_9804,N_9750,N_9621);
or U9805 (N_9805,N_9613,N_9751);
or U9806 (N_9806,N_9610,N_9641);
or U9807 (N_9807,N_9745,N_9601);
xnor U9808 (N_9808,N_9718,N_9639);
nand U9809 (N_9809,N_9689,N_9749);
nor U9810 (N_9810,N_9685,N_9615);
or U9811 (N_9811,N_9687,N_9716);
nor U9812 (N_9812,N_9666,N_9729);
and U9813 (N_9813,N_9726,N_9624);
nor U9814 (N_9814,N_9611,N_9701);
and U9815 (N_9815,N_9631,N_9694);
or U9816 (N_9816,N_9747,N_9713);
or U9817 (N_9817,N_9671,N_9691);
xor U9818 (N_9818,N_9678,N_9755);
nand U9819 (N_9819,N_9658,N_9608);
nand U9820 (N_9820,N_9670,N_9632);
and U9821 (N_9821,N_9616,N_9607);
xnor U9822 (N_9822,N_9655,N_9609);
and U9823 (N_9823,N_9674,N_9669);
nor U9824 (N_9824,N_9651,N_9758);
xnor U9825 (N_9825,N_9622,N_9746);
or U9826 (N_9826,N_9612,N_9715);
nor U9827 (N_9827,N_9686,N_9640);
and U9828 (N_9828,N_9647,N_9635);
nand U9829 (N_9829,N_9756,N_9660);
xor U9830 (N_9830,N_9706,N_9614);
nand U9831 (N_9831,N_9740,N_9605);
nor U9832 (N_9832,N_9722,N_9727);
xor U9833 (N_9833,N_9742,N_9737);
xnor U9834 (N_9834,N_9629,N_9619);
and U9835 (N_9835,N_9643,N_9739);
xor U9836 (N_9836,N_9688,N_9728);
nand U9837 (N_9837,N_9719,N_9690);
nand U9838 (N_9838,N_9603,N_9604);
nand U9839 (N_9839,N_9708,N_9754);
xnor U9840 (N_9840,N_9614,N_9691);
nor U9841 (N_9841,N_9743,N_9713);
and U9842 (N_9842,N_9609,N_9729);
xor U9843 (N_9843,N_9714,N_9752);
xor U9844 (N_9844,N_9673,N_9749);
xnor U9845 (N_9845,N_9634,N_9705);
nor U9846 (N_9846,N_9617,N_9734);
nand U9847 (N_9847,N_9600,N_9730);
nor U9848 (N_9848,N_9698,N_9690);
nand U9849 (N_9849,N_9730,N_9708);
and U9850 (N_9850,N_9738,N_9710);
nand U9851 (N_9851,N_9611,N_9758);
or U9852 (N_9852,N_9700,N_9608);
xor U9853 (N_9853,N_9656,N_9642);
nand U9854 (N_9854,N_9731,N_9671);
xnor U9855 (N_9855,N_9664,N_9646);
nor U9856 (N_9856,N_9633,N_9650);
xnor U9857 (N_9857,N_9639,N_9621);
and U9858 (N_9858,N_9626,N_9726);
nor U9859 (N_9859,N_9690,N_9642);
or U9860 (N_9860,N_9709,N_9630);
and U9861 (N_9861,N_9647,N_9629);
xnor U9862 (N_9862,N_9711,N_9626);
nor U9863 (N_9863,N_9673,N_9624);
nand U9864 (N_9864,N_9715,N_9663);
and U9865 (N_9865,N_9629,N_9634);
and U9866 (N_9866,N_9746,N_9704);
nor U9867 (N_9867,N_9653,N_9625);
nor U9868 (N_9868,N_9609,N_9690);
or U9869 (N_9869,N_9632,N_9706);
and U9870 (N_9870,N_9658,N_9670);
or U9871 (N_9871,N_9758,N_9626);
and U9872 (N_9872,N_9691,N_9718);
nor U9873 (N_9873,N_9729,N_9665);
or U9874 (N_9874,N_9699,N_9656);
nor U9875 (N_9875,N_9742,N_9622);
xnor U9876 (N_9876,N_9623,N_9746);
xnor U9877 (N_9877,N_9649,N_9624);
or U9878 (N_9878,N_9744,N_9630);
nor U9879 (N_9879,N_9668,N_9631);
nor U9880 (N_9880,N_9669,N_9626);
xnor U9881 (N_9881,N_9659,N_9604);
nand U9882 (N_9882,N_9673,N_9747);
or U9883 (N_9883,N_9741,N_9699);
nor U9884 (N_9884,N_9661,N_9715);
xor U9885 (N_9885,N_9638,N_9667);
nor U9886 (N_9886,N_9619,N_9674);
nand U9887 (N_9887,N_9663,N_9610);
or U9888 (N_9888,N_9752,N_9665);
and U9889 (N_9889,N_9694,N_9647);
or U9890 (N_9890,N_9647,N_9737);
or U9891 (N_9891,N_9660,N_9634);
nor U9892 (N_9892,N_9708,N_9689);
nand U9893 (N_9893,N_9694,N_9657);
nor U9894 (N_9894,N_9692,N_9686);
xor U9895 (N_9895,N_9609,N_9732);
or U9896 (N_9896,N_9637,N_9718);
or U9897 (N_9897,N_9727,N_9686);
nor U9898 (N_9898,N_9753,N_9721);
nor U9899 (N_9899,N_9639,N_9697);
nand U9900 (N_9900,N_9648,N_9604);
and U9901 (N_9901,N_9736,N_9643);
or U9902 (N_9902,N_9630,N_9700);
nor U9903 (N_9903,N_9651,N_9616);
nor U9904 (N_9904,N_9651,N_9629);
or U9905 (N_9905,N_9725,N_9728);
nand U9906 (N_9906,N_9721,N_9602);
and U9907 (N_9907,N_9733,N_9672);
and U9908 (N_9908,N_9681,N_9606);
nand U9909 (N_9909,N_9714,N_9690);
nor U9910 (N_9910,N_9684,N_9706);
nand U9911 (N_9911,N_9645,N_9602);
xnor U9912 (N_9912,N_9655,N_9630);
xor U9913 (N_9913,N_9616,N_9718);
or U9914 (N_9914,N_9659,N_9732);
and U9915 (N_9915,N_9630,N_9623);
nor U9916 (N_9916,N_9754,N_9707);
and U9917 (N_9917,N_9716,N_9697);
or U9918 (N_9918,N_9702,N_9634);
and U9919 (N_9919,N_9748,N_9747);
nor U9920 (N_9920,N_9818,N_9804);
and U9921 (N_9921,N_9849,N_9806);
or U9922 (N_9922,N_9797,N_9910);
and U9923 (N_9923,N_9793,N_9764);
nand U9924 (N_9924,N_9809,N_9892);
and U9925 (N_9925,N_9863,N_9816);
nand U9926 (N_9926,N_9912,N_9811);
xor U9927 (N_9927,N_9817,N_9763);
or U9928 (N_9928,N_9865,N_9831);
or U9929 (N_9929,N_9789,N_9827);
xnor U9930 (N_9930,N_9821,N_9768);
nor U9931 (N_9931,N_9779,N_9862);
nand U9932 (N_9932,N_9832,N_9870);
and U9933 (N_9933,N_9904,N_9770);
nor U9934 (N_9934,N_9864,N_9810);
and U9935 (N_9935,N_9909,N_9767);
nor U9936 (N_9936,N_9900,N_9896);
xnor U9937 (N_9937,N_9891,N_9778);
nor U9938 (N_9938,N_9919,N_9785);
nor U9939 (N_9939,N_9895,N_9906);
nor U9940 (N_9940,N_9840,N_9824);
and U9941 (N_9941,N_9799,N_9901);
xnor U9942 (N_9942,N_9781,N_9825);
and U9943 (N_9943,N_9802,N_9869);
xnor U9944 (N_9944,N_9918,N_9813);
nor U9945 (N_9945,N_9888,N_9775);
nor U9946 (N_9946,N_9805,N_9783);
nand U9947 (N_9947,N_9842,N_9815);
nor U9948 (N_9948,N_9847,N_9776);
nor U9949 (N_9949,N_9907,N_9800);
or U9950 (N_9950,N_9860,N_9866);
nor U9951 (N_9951,N_9780,N_9791);
or U9952 (N_9952,N_9852,N_9856);
nor U9953 (N_9953,N_9871,N_9889);
nor U9954 (N_9954,N_9769,N_9880);
nand U9955 (N_9955,N_9808,N_9845);
nand U9956 (N_9956,N_9803,N_9854);
and U9957 (N_9957,N_9873,N_9857);
or U9958 (N_9958,N_9858,N_9872);
and U9959 (N_9959,N_9877,N_9807);
nand U9960 (N_9960,N_9830,N_9826);
and U9961 (N_9961,N_9834,N_9848);
or U9962 (N_9962,N_9794,N_9894);
xnor U9963 (N_9963,N_9801,N_9792);
nor U9964 (N_9964,N_9773,N_9843);
or U9965 (N_9965,N_9878,N_9874);
and U9966 (N_9966,N_9814,N_9837);
xnor U9967 (N_9967,N_9885,N_9823);
or U9968 (N_9968,N_9887,N_9908);
nor U9969 (N_9969,N_9876,N_9771);
nor U9970 (N_9970,N_9846,N_9890);
or U9971 (N_9971,N_9886,N_9820);
xnor U9972 (N_9972,N_9881,N_9774);
xor U9973 (N_9973,N_9844,N_9828);
nand U9974 (N_9974,N_9784,N_9859);
nor U9975 (N_9975,N_9787,N_9777);
or U9976 (N_9976,N_9913,N_9812);
xnor U9977 (N_9977,N_9796,N_9790);
or U9978 (N_9978,N_9822,N_9760);
or U9979 (N_9979,N_9902,N_9850);
xnor U9980 (N_9980,N_9761,N_9861);
and U9981 (N_9981,N_9851,N_9897);
nand U9982 (N_9982,N_9841,N_9899);
or U9983 (N_9983,N_9762,N_9786);
nand U9984 (N_9984,N_9795,N_9883);
nor U9985 (N_9985,N_9855,N_9868);
or U9986 (N_9986,N_9884,N_9839);
nand U9987 (N_9987,N_9766,N_9875);
and U9988 (N_9988,N_9835,N_9882);
xor U9989 (N_9989,N_9867,N_9819);
and U9990 (N_9990,N_9917,N_9914);
nand U9991 (N_9991,N_9879,N_9916);
xor U9992 (N_9992,N_9903,N_9853);
and U9993 (N_9993,N_9836,N_9905);
xnor U9994 (N_9994,N_9772,N_9782);
nor U9995 (N_9995,N_9911,N_9798);
nor U9996 (N_9996,N_9915,N_9765);
or U9997 (N_9997,N_9829,N_9898);
or U9998 (N_9998,N_9833,N_9788);
and U9999 (N_9999,N_9893,N_9838);
nor U10000 (N_10000,N_9898,N_9770);
or U10001 (N_10001,N_9824,N_9878);
and U10002 (N_10002,N_9846,N_9802);
nor U10003 (N_10003,N_9811,N_9775);
xnor U10004 (N_10004,N_9903,N_9808);
and U10005 (N_10005,N_9877,N_9888);
or U10006 (N_10006,N_9898,N_9918);
nand U10007 (N_10007,N_9793,N_9880);
and U10008 (N_10008,N_9839,N_9886);
nand U10009 (N_10009,N_9786,N_9772);
or U10010 (N_10010,N_9845,N_9765);
and U10011 (N_10011,N_9849,N_9859);
and U10012 (N_10012,N_9793,N_9763);
or U10013 (N_10013,N_9834,N_9915);
and U10014 (N_10014,N_9832,N_9848);
or U10015 (N_10015,N_9894,N_9861);
xor U10016 (N_10016,N_9810,N_9852);
or U10017 (N_10017,N_9886,N_9805);
or U10018 (N_10018,N_9785,N_9874);
and U10019 (N_10019,N_9892,N_9783);
nor U10020 (N_10020,N_9870,N_9771);
nor U10021 (N_10021,N_9796,N_9774);
xor U10022 (N_10022,N_9780,N_9787);
xor U10023 (N_10023,N_9804,N_9849);
and U10024 (N_10024,N_9914,N_9875);
xnor U10025 (N_10025,N_9779,N_9834);
nor U10026 (N_10026,N_9831,N_9779);
nor U10027 (N_10027,N_9860,N_9859);
nor U10028 (N_10028,N_9874,N_9867);
or U10029 (N_10029,N_9910,N_9839);
nand U10030 (N_10030,N_9760,N_9772);
nand U10031 (N_10031,N_9856,N_9868);
nor U10032 (N_10032,N_9880,N_9798);
and U10033 (N_10033,N_9795,N_9906);
nor U10034 (N_10034,N_9785,N_9912);
nand U10035 (N_10035,N_9910,N_9761);
nand U10036 (N_10036,N_9865,N_9855);
and U10037 (N_10037,N_9891,N_9789);
nor U10038 (N_10038,N_9874,N_9811);
or U10039 (N_10039,N_9764,N_9874);
xor U10040 (N_10040,N_9813,N_9907);
nand U10041 (N_10041,N_9814,N_9838);
or U10042 (N_10042,N_9767,N_9789);
or U10043 (N_10043,N_9908,N_9812);
and U10044 (N_10044,N_9818,N_9793);
nor U10045 (N_10045,N_9907,N_9764);
nand U10046 (N_10046,N_9877,N_9863);
xnor U10047 (N_10047,N_9828,N_9911);
nor U10048 (N_10048,N_9906,N_9769);
xnor U10049 (N_10049,N_9761,N_9766);
nand U10050 (N_10050,N_9772,N_9915);
and U10051 (N_10051,N_9919,N_9880);
xor U10052 (N_10052,N_9816,N_9769);
xnor U10053 (N_10053,N_9903,N_9836);
nor U10054 (N_10054,N_9858,N_9878);
xor U10055 (N_10055,N_9904,N_9772);
and U10056 (N_10056,N_9862,N_9881);
nand U10057 (N_10057,N_9836,N_9909);
and U10058 (N_10058,N_9802,N_9902);
nor U10059 (N_10059,N_9918,N_9913);
xor U10060 (N_10060,N_9780,N_9907);
nor U10061 (N_10061,N_9890,N_9793);
or U10062 (N_10062,N_9886,N_9904);
or U10063 (N_10063,N_9887,N_9844);
nor U10064 (N_10064,N_9885,N_9812);
nand U10065 (N_10065,N_9851,N_9860);
xnor U10066 (N_10066,N_9912,N_9905);
and U10067 (N_10067,N_9872,N_9826);
nor U10068 (N_10068,N_9763,N_9916);
nand U10069 (N_10069,N_9834,N_9802);
nand U10070 (N_10070,N_9804,N_9882);
xnor U10071 (N_10071,N_9773,N_9855);
and U10072 (N_10072,N_9825,N_9799);
nor U10073 (N_10073,N_9882,N_9763);
xor U10074 (N_10074,N_9894,N_9783);
nand U10075 (N_10075,N_9826,N_9828);
nor U10076 (N_10076,N_9918,N_9800);
or U10077 (N_10077,N_9783,N_9878);
nor U10078 (N_10078,N_9826,N_9884);
or U10079 (N_10079,N_9788,N_9894);
or U10080 (N_10080,N_10019,N_10035);
nor U10081 (N_10081,N_9996,N_10048);
nor U10082 (N_10082,N_9936,N_9924);
or U10083 (N_10083,N_10040,N_10001);
xor U10084 (N_10084,N_10014,N_10054);
nor U10085 (N_10085,N_10007,N_9920);
or U10086 (N_10086,N_9953,N_9923);
nor U10087 (N_10087,N_10036,N_10004);
nor U10088 (N_10088,N_9932,N_9997);
or U10089 (N_10089,N_9955,N_9956);
xnor U10090 (N_10090,N_9976,N_10031);
and U10091 (N_10091,N_9922,N_9945);
nor U10092 (N_10092,N_9967,N_10015);
xnor U10093 (N_10093,N_10030,N_10065);
nor U10094 (N_10094,N_10060,N_10066);
or U10095 (N_10095,N_10037,N_10057);
or U10096 (N_10096,N_9950,N_10072);
nor U10097 (N_10097,N_9987,N_9954);
or U10098 (N_10098,N_10075,N_9988);
and U10099 (N_10099,N_9999,N_9938);
nand U10100 (N_10100,N_10028,N_10011);
nand U10101 (N_10101,N_10008,N_9975);
nand U10102 (N_10102,N_10047,N_10049);
nor U10103 (N_10103,N_10023,N_9931);
nor U10104 (N_10104,N_9926,N_10029);
or U10105 (N_10105,N_9971,N_10022);
xor U10106 (N_10106,N_10016,N_10002);
or U10107 (N_10107,N_9947,N_10073);
nor U10108 (N_10108,N_9948,N_10064);
and U10109 (N_10109,N_10071,N_10010);
or U10110 (N_10110,N_9928,N_9992);
xor U10111 (N_10111,N_9959,N_10017);
or U10112 (N_10112,N_9964,N_9972);
xnor U10113 (N_10113,N_9962,N_10013);
nor U10114 (N_10114,N_10009,N_10056);
nor U10115 (N_10115,N_10039,N_9968);
or U10116 (N_10116,N_9985,N_10050);
and U10117 (N_10117,N_10067,N_10038);
xnor U10118 (N_10118,N_9951,N_10069);
or U10119 (N_10119,N_10003,N_10079);
xnor U10120 (N_10120,N_10078,N_9933);
xor U10121 (N_10121,N_9963,N_9991);
nor U10122 (N_10122,N_9978,N_10034);
nand U10123 (N_10123,N_10005,N_10044);
or U10124 (N_10124,N_9977,N_9989);
or U10125 (N_10125,N_9966,N_10063);
xnor U10126 (N_10126,N_10024,N_9981);
nand U10127 (N_10127,N_10000,N_10018);
nor U10128 (N_10128,N_10027,N_9980);
xnor U10129 (N_10129,N_9943,N_10042);
nand U10130 (N_10130,N_9944,N_9958);
xnor U10131 (N_10131,N_9952,N_10074);
and U10132 (N_10132,N_9946,N_10041);
and U10133 (N_10133,N_9973,N_10021);
and U10134 (N_10134,N_9942,N_10025);
nor U10135 (N_10135,N_9930,N_10068);
nor U10136 (N_10136,N_10077,N_10076);
xnor U10137 (N_10137,N_9990,N_9927);
xor U10138 (N_10138,N_10062,N_9939);
or U10139 (N_10139,N_9929,N_9979);
nand U10140 (N_10140,N_9941,N_10051);
nand U10141 (N_10141,N_9970,N_9957);
xnor U10142 (N_10142,N_10043,N_9974);
and U10143 (N_10143,N_10046,N_10055);
nor U10144 (N_10144,N_9937,N_9965);
and U10145 (N_10145,N_10061,N_9934);
or U10146 (N_10146,N_9969,N_10033);
nor U10147 (N_10147,N_10059,N_9983);
and U10148 (N_10148,N_9940,N_9935);
xnor U10149 (N_10149,N_10012,N_9982);
and U10150 (N_10150,N_10053,N_9993);
or U10151 (N_10151,N_9986,N_9961);
xor U10152 (N_10152,N_10052,N_9921);
xor U10153 (N_10153,N_9995,N_9984);
or U10154 (N_10154,N_10045,N_10058);
and U10155 (N_10155,N_9960,N_9949);
nor U10156 (N_10156,N_10020,N_9998);
xor U10157 (N_10157,N_10026,N_9925);
nand U10158 (N_10158,N_9994,N_10006);
xnor U10159 (N_10159,N_10032,N_10070);
nor U10160 (N_10160,N_10074,N_10046);
xnor U10161 (N_10161,N_9980,N_9958);
nand U10162 (N_10162,N_9951,N_9929);
nand U10163 (N_10163,N_9941,N_10008);
and U10164 (N_10164,N_9930,N_9979);
or U10165 (N_10165,N_10044,N_10030);
or U10166 (N_10166,N_9939,N_9956);
and U10167 (N_10167,N_9999,N_9959);
nand U10168 (N_10168,N_9939,N_10030);
and U10169 (N_10169,N_10013,N_10071);
nand U10170 (N_10170,N_9994,N_9978);
and U10171 (N_10171,N_10013,N_10026);
nor U10172 (N_10172,N_10069,N_10076);
xnor U10173 (N_10173,N_9988,N_10029);
or U10174 (N_10174,N_10065,N_10028);
xor U10175 (N_10175,N_10007,N_9951);
nor U10176 (N_10176,N_9964,N_9968);
xor U10177 (N_10177,N_9930,N_10001);
xnor U10178 (N_10178,N_9941,N_10053);
nor U10179 (N_10179,N_10053,N_10052);
nand U10180 (N_10180,N_10019,N_10072);
xnor U10181 (N_10181,N_9948,N_9935);
and U10182 (N_10182,N_10063,N_9933);
and U10183 (N_10183,N_9961,N_10019);
xor U10184 (N_10184,N_10028,N_9947);
xnor U10185 (N_10185,N_9926,N_10056);
or U10186 (N_10186,N_9967,N_9970);
and U10187 (N_10187,N_9941,N_10058);
nor U10188 (N_10188,N_10039,N_9937);
and U10189 (N_10189,N_9923,N_9967);
nand U10190 (N_10190,N_10014,N_9969);
nand U10191 (N_10191,N_10069,N_10068);
nand U10192 (N_10192,N_9976,N_9984);
and U10193 (N_10193,N_9967,N_10038);
nand U10194 (N_10194,N_9952,N_9999);
nor U10195 (N_10195,N_10052,N_9985);
nand U10196 (N_10196,N_10048,N_9979);
nand U10197 (N_10197,N_9996,N_9920);
and U10198 (N_10198,N_10041,N_9994);
nand U10199 (N_10199,N_9986,N_9970);
or U10200 (N_10200,N_9983,N_9928);
and U10201 (N_10201,N_9995,N_10059);
or U10202 (N_10202,N_10022,N_10074);
xnor U10203 (N_10203,N_10045,N_10005);
and U10204 (N_10204,N_10012,N_9987);
nand U10205 (N_10205,N_10015,N_9953);
and U10206 (N_10206,N_10062,N_10016);
or U10207 (N_10207,N_10008,N_9939);
xor U10208 (N_10208,N_9989,N_10035);
nor U10209 (N_10209,N_10071,N_10077);
nor U10210 (N_10210,N_9941,N_9960);
xnor U10211 (N_10211,N_9988,N_10004);
or U10212 (N_10212,N_9984,N_9949);
or U10213 (N_10213,N_9956,N_9927);
xnor U10214 (N_10214,N_9973,N_9944);
xor U10215 (N_10215,N_10027,N_10021);
nand U10216 (N_10216,N_9967,N_9992);
xor U10217 (N_10217,N_10057,N_10048);
or U10218 (N_10218,N_10056,N_10000);
nor U10219 (N_10219,N_9978,N_9922);
or U10220 (N_10220,N_10021,N_10009);
xnor U10221 (N_10221,N_10079,N_10043);
xnor U10222 (N_10222,N_10020,N_9962);
and U10223 (N_10223,N_10007,N_9961);
xnor U10224 (N_10224,N_9995,N_9964);
and U10225 (N_10225,N_9935,N_10005);
xor U10226 (N_10226,N_10041,N_10069);
or U10227 (N_10227,N_9934,N_10017);
xor U10228 (N_10228,N_9926,N_9982);
nand U10229 (N_10229,N_9986,N_10054);
nor U10230 (N_10230,N_10019,N_9937);
or U10231 (N_10231,N_10050,N_9974);
nor U10232 (N_10232,N_9956,N_10038);
nor U10233 (N_10233,N_10045,N_9995);
xor U10234 (N_10234,N_9973,N_10025);
xor U10235 (N_10235,N_9948,N_10033);
nand U10236 (N_10236,N_10040,N_10050);
or U10237 (N_10237,N_10066,N_9951);
nor U10238 (N_10238,N_9931,N_10059);
or U10239 (N_10239,N_9976,N_9959);
nand U10240 (N_10240,N_10177,N_10090);
nor U10241 (N_10241,N_10227,N_10136);
nand U10242 (N_10242,N_10230,N_10186);
xor U10243 (N_10243,N_10133,N_10150);
or U10244 (N_10244,N_10106,N_10143);
and U10245 (N_10245,N_10094,N_10174);
xor U10246 (N_10246,N_10134,N_10115);
xor U10247 (N_10247,N_10221,N_10180);
nor U10248 (N_10248,N_10110,N_10122);
nand U10249 (N_10249,N_10140,N_10225);
xor U10250 (N_10250,N_10200,N_10109);
or U10251 (N_10251,N_10183,N_10100);
or U10252 (N_10252,N_10193,N_10154);
and U10253 (N_10253,N_10214,N_10147);
nand U10254 (N_10254,N_10121,N_10219);
nand U10255 (N_10255,N_10162,N_10172);
and U10256 (N_10256,N_10080,N_10210);
xor U10257 (N_10257,N_10197,N_10223);
xnor U10258 (N_10258,N_10199,N_10169);
nor U10259 (N_10259,N_10222,N_10152);
xor U10260 (N_10260,N_10141,N_10085);
or U10261 (N_10261,N_10168,N_10101);
and U10262 (N_10262,N_10204,N_10086);
and U10263 (N_10263,N_10120,N_10153);
nor U10264 (N_10264,N_10108,N_10132);
nor U10265 (N_10265,N_10159,N_10087);
nor U10266 (N_10266,N_10170,N_10192);
nand U10267 (N_10267,N_10190,N_10194);
nor U10268 (N_10268,N_10083,N_10182);
or U10269 (N_10269,N_10158,N_10217);
nor U10270 (N_10270,N_10178,N_10187);
nor U10271 (N_10271,N_10232,N_10220);
nand U10272 (N_10272,N_10111,N_10179);
xor U10273 (N_10273,N_10216,N_10104);
or U10274 (N_10274,N_10116,N_10119);
and U10275 (N_10275,N_10139,N_10195);
and U10276 (N_10276,N_10185,N_10099);
or U10277 (N_10277,N_10123,N_10117);
or U10278 (N_10278,N_10184,N_10157);
and U10279 (N_10279,N_10093,N_10163);
and U10280 (N_10280,N_10175,N_10207);
nor U10281 (N_10281,N_10088,N_10084);
and U10282 (N_10282,N_10126,N_10129);
xnor U10283 (N_10283,N_10107,N_10124);
nand U10284 (N_10284,N_10130,N_10092);
xor U10285 (N_10285,N_10226,N_10224);
nand U10286 (N_10286,N_10156,N_10173);
and U10287 (N_10287,N_10128,N_10238);
and U10288 (N_10288,N_10202,N_10098);
xor U10289 (N_10289,N_10161,N_10114);
nand U10290 (N_10290,N_10196,N_10105);
and U10291 (N_10291,N_10148,N_10205);
and U10292 (N_10292,N_10137,N_10164);
or U10293 (N_10293,N_10138,N_10082);
nand U10294 (N_10294,N_10228,N_10096);
nor U10295 (N_10295,N_10176,N_10089);
xnor U10296 (N_10296,N_10081,N_10229);
nor U10297 (N_10297,N_10125,N_10237);
xnor U10298 (N_10298,N_10239,N_10135);
or U10299 (N_10299,N_10131,N_10112);
and U10300 (N_10300,N_10095,N_10145);
nand U10301 (N_10301,N_10206,N_10103);
xnor U10302 (N_10302,N_10091,N_10102);
xnor U10303 (N_10303,N_10213,N_10208);
xor U10304 (N_10304,N_10171,N_10203);
and U10305 (N_10305,N_10151,N_10160);
and U10306 (N_10306,N_10149,N_10189);
or U10307 (N_10307,N_10211,N_10215);
xor U10308 (N_10308,N_10167,N_10155);
xnor U10309 (N_10309,N_10235,N_10146);
nor U10310 (N_10310,N_10181,N_10209);
nand U10311 (N_10311,N_10127,N_10231);
xor U10312 (N_10312,N_10144,N_10191);
xnor U10313 (N_10313,N_10234,N_10118);
and U10314 (N_10314,N_10113,N_10165);
xor U10315 (N_10315,N_10166,N_10142);
nor U10316 (N_10316,N_10233,N_10236);
xnor U10317 (N_10317,N_10218,N_10097);
and U10318 (N_10318,N_10188,N_10201);
or U10319 (N_10319,N_10198,N_10212);
xnor U10320 (N_10320,N_10081,N_10235);
or U10321 (N_10321,N_10174,N_10208);
or U10322 (N_10322,N_10089,N_10108);
and U10323 (N_10323,N_10128,N_10227);
or U10324 (N_10324,N_10116,N_10091);
or U10325 (N_10325,N_10132,N_10101);
and U10326 (N_10326,N_10088,N_10206);
xor U10327 (N_10327,N_10140,N_10227);
nor U10328 (N_10328,N_10173,N_10100);
and U10329 (N_10329,N_10157,N_10218);
nand U10330 (N_10330,N_10208,N_10169);
nor U10331 (N_10331,N_10186,N_10193);
xnor U10332 (N_10332,N_10236,N_10134);
nand U10333 (N_10333,N_10174,N_10211);
and U10334 (N_10334,N_10122,N_10139);
xnor U10335 (N_10335,N_10151,N_10090);
xor U10336 (N_10336,N_10159,N_10152);
and U10337 (N_10337,N_10151,N_10165);
nand U10338 (N_10338,N_10144,N_10146);
nor U10339 (N_10339,N_10107,N_10096);
nor U10340 (N_10340,N_10210,N_10189);
nand U10341 (N_10341,N_10207,N_10198);
nand U10342 (N_10342,N_10235,N_10113);
xnor U10343 (N_10343,N_10215,N_10172);
nand U10344 (N_10344,N_10090,N_10211);
and U10345 (N_10345,N_10204,N_10147);
xor U10346 (N_10346,N_10080,N_10238);
nand U10347 (N_10347,N_10095,N_10116);
nand U10348 (N_10348,N_10092,N_10204);
nor U10349 (N_10349,N_10172,N_10148);
xnor U10350 (N_10350,N_10151,N_10182);
or U10351 (N_10351,N_10217,N_10202);
or U10352 (N_10352,N_10223,N_10135);
and U10353 (N_10353,N_10129,N_10236);
nand U10354 (N_10354,N_10134,N_10227);
and U10355 (N_10355,N_10116,N_10168);
nor U10356 (N_10356,N_10208,N_10117);
xor U10357 (N_10357,N_10199,N_10177);
and U10358 (N_10358,N_10230,N_10139);
nand U10359 (N_10359,N_10149,N_10081);
nor U10360 (N_10360,N_10101,N_10205);
xnor U10361 (N_10361,N_10159,N_10162);
xnor U10362 (N_10362,N_10147,N_10111);
and U10363 (N_10363,N_10163,N_10152);
nand U10364 (N_10364,N_10128,N_10228);
and U10365 (N_10365,N_10194,N_10220);
nor U10366 (N_10366,N_10229,N_10226);
nand U10367 (N_10367,N_10186,N_10084);
nand U10368 (N_10368,N_10141,N_10111);
xnor U10369 (N_10369,N_10190,N_10168);
nor U10370 (N_10370,N_10214,N_10092);
and U10371 (N_10371,N_10174,N_10122);
nand U10372 (N_10372,N_10165,N_10223);
or U10373 (N_10373,N_10215,N_10132);
and U10374 (N_10374,N_10098,N_10114);
nand U10375 (N_10375,N_10082,N_10094);
nor U10376 (N_10376,N_10121,N_10160);
and U10377 (N_10377,N_10142,N_10090);
nor U10378 (N_10378,N_10228,N_10194);
nand U10379 (N_10379,N_10223,N_10120);
and U10380 (N_10380,N_10114,N_10137);
nand U10381 (N_10381,N_10102,N_10122);
xor U10382 (N_10382,N_10116,N_10205);
xor U10383 (N_10383,N_10114,N_10224);
or U10384 (N_10384,N_10212,N_10166);
or U10385 (N_10385,N_10209,N_10235);
nand U10386 (N_10386,N_10208,N_10235);
or U10387 (N_10387,N_10163,N_10208);
nand U10388 (N_10388,N_10132,N_10186);
nand U10389 (N_10389,N_10224,N_10142);
and U10390 (N_10390,N_10084,N_10219);
nor U10391 (N_10391,N_10190,N_10152);
and U10392 (N_10392,N_10198,N_10178);
nand U10393 (N_10393,N_10150,N_10125);
or U10394 (N_10394,N_10103,N_10239);
nand U10395 (N_10395,N_10235,N_10204);
nand U10396 (N_10396,N_10136,N_10085);
and U10397 (N_10397,N_10092,N_10210);
nor U10398 (N_10398,N_10239,N_10124);
xor U10399 (N_10399,N_10229,N_10082);
or U10400 (N_10400,N_10365,N_10288);
xnor U10401 (N_10401,N_10350,N_10281);
nand U10402 (N_10402,N_10260,N_10352);
and U10403 (N_10403,N_10266,N_10251);
nor U10404 (N_10404,N_10318,N_10290);
and U10405 (N_10405,N_10277,N_10264);
xor U10406 (N_10406,N_10245,N_10397);
and U10407 (N_10407,N_10341,N_10354);
nand U10408 (N_10408,N_10263,N_10301);
or U10409 (N_10409,N_10374,N_10310);
nor U10410 (N_10410,N_10314,N_10346);
or U10411 (N_10411,N_10246,N_10317);
or U10412 (N_10412,N_10391,N_10345);
and U10413 (N_10413,N_10329,N_10387);
and U10414 (N_10414,N_10243,N_10366);
and U10415 (N_10415,N_10254,N_10364);
and U10416 (N_10416,N_10315,N_10340);
or U10417 (N_10417,N_10355,N_10271);
and U10418 (N_10418,N_10291,N_10383);
xnor U10419 (N_10419,N_10344,N_10368);
and U10420 (N_10420,N_10381,N_10392);
nand U10421 (N_10421,N_10363,N_10370);
xor U10422 (N_10422,N_10250,N_10375);
nand U10423 (N_10423,N_10295,N_10362);
nor U10424 (N_10424,N_10268,N_10393);
or U10425 (N_10425,N_10316,N_10303);
nor U10426 (N_10426,N_10358,N_10371);
and U10427 (N_10427,N_10379,N_10388);
nor U10428 (N_10428,N_10322,N_10247);
and U10429 (N_10429,N_10382,N_10339);
nand U10430 (N_10430,N_10267,N_10289);
or U10431 (N_10431,N_10256,N_10279);
nand U10432 (N_10432,N_10257,N_10385);
and U10433 (N_10433,N_10321,N_10262);
xnor U10434 (N_10434,N_10324,N_10276);
nand U10435 (N_10435,N_10356,N_10330);
xor U10436 (N_10436,N_10286,N_10376);
xor U10437 (N_10437,N_10325,N_10309);
or U10438 (N_10438,N_10394,N_10326);
and U10439 (N_10439,N_10328,N_10361);
nand U10440 (N_10440,N_10274,N_10304);
nand U10441 (N_10441,N_10311,N_10248);
xor U10442 (N_10442,N_10283,N_10265);
xor U10443 (N_10443,N_10269,N_10259);
nor U10444 (N_10444,N_10360,N_10395);
nand U10445 (N_10445,N_10313,N_10242);
and U10446 (N_10446,N_10386,N_10398);
and U10447 (N_10447,N_10396,N_10323);
nor U10448 (N_10448,N_10333,N_10327);
xnor U10449 (N_10449,N_10390,N_10338);
or U10450 (N_10450,N_10253,N_10320);
xor U10451 (N_10451,N_10336,N_10319);
xor U10452 (N_10452,N_10351,N_10299);
xor U10453 (N_10453,N_10273,N_10252);
or U10454 (N_10454,N_10305,N_10284);
nor U10455 (N_10455,N_10308,N_10240);
nor U10456 (N_10456,N_10297,N_10302);
xor U10457 (N_10457,N_10300,N_10380);
nand U10458 (N_10458,N_10367,N_10292);
nand U10459 (N_10459,N_10278,N_10270);
and U10460 (N_10460,N_10384,N_10399);
nor U10461 (N_10461,N_10335,N_10275);
xnor U10462 (N_10462,N_10369,N_10306);
or U10463 (N_10463,N_10287,N_10241);
nor U10464 (N_10464,N_10334,N_10296);
or U10465 (N_10465,N_10353,N_10347);
nor U10466 (N_10466,N_10342,N_10348);
and U10467 (N_10467,N_10337,N_10244);
xnor U10468 (N_10468,N_10294,N_10359);
and U10469 (N_10469,N_10389,N_10357);
nand U10470 (N_10470,N_10378,N_10377);
nand U10471 (N_10471,N_10331,N_10249);
and U10472 (N_10472,N_10373,N_10293);
xnor U10473 (N_10473,N_10349,N_10298);
or U10474 (N_10474,N_10282,N_10312);
xnor U10475 (N_10475,N_10307,N_10255);
and U10476 (N_10476,N_10343,N_10372);
or U10477 (N_10477,N_10280,N_10258);
nand U10478 (N_10478,N_10272,N_10261);
nor U10479 (N_10479,N_10285,N_10332);
nor U10480 (N_10480,N_10271,N_10309);
nor U10481 (N_10481,N_10276,N_10302);
nor U10482 (N_10482,N_10308,N_10356);
and U10483 (N_10483,N_10347,N_10313);
and U10484 (N_10484,N_10362,N_10303);
nand U10485 (N_10485,N_10270,N_10262);
nor U10486 (N_10486,N_10385,N_10351);
and U10487 (N_10487,N_10387,N_10282);
nand U10488 (N_10488,N_10288,N_10386);
xor U10489 (N_10489,N_10393,N_10315);
or U10490 (N_10490,N_10359,N_10346);
nor U10491 (N_10491,N_10378,N_10313);
nor U10492 (N_10492,N_10250,N_10311);
xor U10493 (N_10493,N_10296,N_10274);
or U10494 (N_10494,N_10277,N_10371);
xor U10495 (N_10495,N_10267,N_10240);
xnor U10496 (N_10496,N_10347,N_10397);
nand U10497 (N_10497,N_10287,N_10358);
nor U10498 (N_10498,N_10332,N_10329);
nor U10499 (N_10499,N_10318,N_10320);
or U10500 (N_10500,N_10338,N_10359);
xnor U10501 (N_10501,N_10323,N_10319);
or U10502 (N_10502,N_10356,N_10248);
nand U10503 (N_10503,N_10346,N_10356);
and U10504 (N_10504,N_10319,N_10379);
or U10505 (N_10505,N_10355,N_10384);
nand U10506 (N_10506,N_10312,N_10391);
and U10507 (N_10507,N_10397,N_10261);
nor U10508 (N_10508,N_10313,N_10250);
and U10509 (N_10509,N_10374,N_10326);
or U10510 (N_10510,N_10280,N_10363);
nor U10511 (N_10511,N_10311,N_10368);
or U10512 (N_10512,N_10335,N_10384);
xnor U10513 (N_10513,N_10399,N_10377);
and U10514 (N_10514,N_10333,N_10312);
or U10515 (N_10515,N_10396,N_10321);
or U10516 (N_10516,N_10300,N_10326);
or U10517 (N_10517,N_10288,N_10378);
or U10518 (N_10518,N_10363,N_10316);
nor U10519 (N_10519,N_10284,N_10277);
xnor U10520 (N_10520,N_10317,N_10384);
and U10521 (N_10521,N_10362,N_10316);
nand U10522 (N_10522,N_10253,N_10294);
or U10523 (N_10523,N_10320,N_10357);
xnor U10524 (N_10524,N_10318,N_10277);
and U10525 (N_10525,N_10242,N_10397);
nand U10526 (N_10526,N_10333,N_10334);
and U10527 (N_10527,N_10339,N_10282);
and U10528 (N_10528,N_10396,N_10287);
and U10529 (N_10529,N_10304,N_10314);
and U10530 (N_10530,N_10299,N_10290);
xnor U10531 (N_10531,N_10299,N_10385);
or U10532 (N_10532,N_10374,N_10360);
nor U10533 (N_10533,N_10354,N_10353);
xor U10534 (N_10534,N_10289,N_10323);
xor U10535 (N_10535,N_10329,N_10257);
and U10536 (N_10536,N_10271,N_10314);
nor U10537 (N_10537,N_10296,N_10394);
or U10538 (N_10538,N_10243,N_10274);
nor U10539 (N_10539,N_10253,N_10336);
nand U10540 (N_10540,N_10341,N_10299);
or U10541 (N_10541,N_10364,N_10329);
nand U10542 (N_10542,N_10335,N_10320);
nor U10543 (N_10543,N_10247,N_10377);
and U10544 (N_10544,N_10266,N_10353);
nor U10545 (N_10545,N_10306,N_10349);
nor U10546 (N_10546,N_10301,N_10387);
and U10547 (N_10547,N_10309,N_10288);
nand U10548 (N_10548,N_10268,N_10343);
nor U10549 (N_10549,N_10332,N_10342);
nand U10550 (N_10550,N_10348,N_10254);
nor U10551 (N_10551,N_10265,N_10388);
or U10552 (N_10552,N_10336,N_10293);
nor U10553 (N_10553,N_10245,N_10352);
nand U10554 (N_10554,N_10261,N_10375);
nand U10555 (N_10555,N_10240,N_10328);
or U10556 (N_10556,N_10370,N_10318);
and U10557 (N_10557,N_10302,N_10251);
nand U10558 (N_10558,N_10352,N_10325);
nand U10559 (N_10559,N_10363,N_10346);
and U10560 (N_10560,N_10423,N_10416);
and U10561 (N_10561,N_10476,N_10458);
or U10562 (N_10562,N_10486,N_10403);
or U10563 (N_10563,N_10537,N_10530);
nor U10564 (N_10564,N_10503,N_10527);
nor U10565 (N_10565,N_10519,N_10495);
or U10566 (N_10566,N_10426,N_10415);
and U10567 (N_10567,N_10522,N_10524);
or U10568 (N_10568,N_10494,N_10454);
nor U10569 (N_10569,N_10430,N_10433);
xor U10570 (N_10570,N_10501,N_10437);
nor U10571 (N_10571,N_10513,N_10472);
or U10572 (N_10572,N_10462,N_10531);
and U10573 (N_10573,N_10525,N_10457);
or U10574 (N_10574,N_10424,N_10410);
or U10575 (N_10575,N_10490,N_10523);
and U10576 (N_10576,N_10418,N_10404);
and U10577 (N_10577,N_10460,N_10409);
or U10578 (N_10578,N_10496,N_10540);
or U10579 (N_10579,N_10507,N_10548);
nor U10580 (N_10580,N_10413,N_10480);
xnor U10581 (N_10581,N_10556,N_10508);
and U10582 (N_10582,N_10559,N_10474);
or U10583 (N_10583,N_10401,N_10434);
nand U10584 (N_10584,N_10557,N_10478);
nor U10585 (N_10585,N_10493,N_10541);
or U10586 (N_10586,N_10431,N_10505);
nor U10587 (N_10587,N_10445,N_10506);
nand U10588 (N_10588,N_10482,N_10533);
nand U10589 (N_10589,N_10544,N_10439);
nand U10590 (N_10590,N_10481,N_10411);
and U10591 (N_10591,N_10528,N_10488);
and U10592 (N_10592,N_10517,N_10449);
nand U10593 (N_10593,N_10440,N_10498);
xor U10594 (N_10594,N_10516,N_10463);
xnor U10595 (N_10595,N_10470,N_10412);
xor U10596 (N_10596,N_10536,N_10405);
nand U10597 (N_10597,N_10421,N_10538);
xnor U10598 (N_10598,N_10558,N_10499);
or U10599 (N_10599,N_10497,N_10444);
nand U10600 (N_10600,N_10436,N_10402);
nor U10601 (N_10601,N_10465,N_10448);
or U10602 (N_10602,N_10500,N_10492);
nor U10603 (N_10603,N_10429,N_10441);
xnor U10604 (N_10604,N_10443,N_10514);
and U10605 (N_10605,N_10502,N_10475);
or U10606 (N_10606,N_10504,N_10483);
or U10607 (N_10607,N_10529,N_10408);
and U10608 (N_10608,N_10451,N_10442);
xnor U10609 (N_10609,N_10555,N_10487);
and U10610 (N_10610,N_10471,N_10521);
or U10611 (N_10611,N_10468,N_10464);
or U10612 (N_10612,N_10406,N_10477);
or U10613 (N_10613,N_10489,N_10512);
nor U10614 (N_10614,N_10547,N_10414);
xnor U10615 (N_10615,N_10435,N_10420);
nand U10616 (N_10616,N_10450,N_10438);
and U10617 (N_10617,N_10550,N_10509);
or U10618 (N_10618,N_10552,N_10485);
and U10619 (N_10619,N_10427,N_10526);
nor U10620 (N_10620,N_10539,N_10425);
and U10621 (N_10621,N_10520,N_10551);
xor U10622 (N_10622,N_10428,N_10546);
and U10623 (N_10623,N_10510,N_10473);
nand U10624 (N_10624,N_10400,N_10461);
or U10625 (N_10625,N_10432,N_10452);
and U10626 (N_10626,N_10419,N_10549);
and U10627 (N_10627,N_10535,N_10456);
nor U10628 (N_10628,N_10515,N_10447);
or U10629 (N_10629,N_10484,N_10417);
and U10630 (N_10630,N_10518,N_10511);
xor U10631 (N_10631,N_10446,N_10545);
nand U10632 (N_10632,N_10491,N_10554);
nand U10633 (N_10633,N_10459,N_10469);
or U10634 (N_10634,N_10455,N_10542);
and U10635 (N_10635,N_10553,N_10453);
nand U10636 (N_10636,N_10532,N_10479);
nor U10637 (N_10637,N_10422,N_10543);
nand U10638 (N_10638,N_10467,N_10466);
or U10639 (N_10639,N_10534,N_10407);
xnor U10640 (N_10640,N_10516,N_10552);
or U10641 (N_10641,N_10409,N_10497);
or U10642 (N_10642,N_10530,N_10541);
or U10643 (N_10643,N_10487,N_10511);
or U10644 (N_10644,N_10401,N_10531);
nor U10645 (N_10645,N_10522,N_10471);
or U10646 (N_10646,N_10558,N_10544);
xnor U10647 (N_10647,N_10411,N_10517);
or U10648 (N_10648,N_10442,N_10482);
xnor U10649 (N_10649,N_10484,N_10537);
xor U10650 (N_10650,N_10525,N_10448);
nand U10651 (N_10651,N_10533,N_10522);
nor U10652 (N_10652,N_10544,N_10505);
nor U10653 (N_10653,N_10489,N_10455);
and U10654 (N_10654,N_10549,N_10408);
xnor U10655 (N_10655,N_10516,N_10545);
nand U10656 (N_10656,N_10413,N_10502);
nand U10657 (N_10657,N_10445,N_10426);
xor U10658 (N_10658,N_10410,N_10459);
or U10659 (N_10659,N_10405,N_10437);
and U10660 (N_10660,N_10448,N_10498);
nor U10661 (N_10661,N_10402,N_10478);
or U10662 (N_10662,N_10546,N_10462);
nand U10663 (N_10663,N_10445,N_10450);
xnor U10664 (N_10664,N_10534,N_10463);
nor U10665 (N_10665,N_10444,N_10419);
xnor U10666 (N_10666,N_10559,N_10558);
nand U10667 (N_10667,N_10475,N_10461);
nor U10668 (N_10668,N_10468,N_10512);
or U10669 (N_10669,N_10452,N_10508);
or U10670 (N_10670,N_10461,N_10469);
and U10671 (N_10671,N_10457,N_10494);
nor U10672 (N_10672,N_10514,N_10484);
and U10673 (N_10673,N_10553,N_10427);
nor U10674 (N_10674,N_10469,N_10422);
and U10675 (N_10675,N_10415,N_10475);
xnor U10676 (N_10676,N_10539,N_10405);
xnor U10677 (N_10677,N_10401,N_10484);
xnor U10678 (N_10678,N_10476,N_10462);
and U10679 (N_10679,N_10432,N_10507);
nor U10680 (N_10680,N_10479,N_10441);
xor U10681 (N_10681,N_10528,N_10514);
nor U10682 (N_10682,N_10544,N_10538);
or U10683 (N_10683,N_10476,N_10556);
nor U10684 (N_10684,N_10439,N_10504);
or U10685 (N_10685,N_10481,N_10429);
nor U10686 (N_10686,N_10407,N_10519);
nand U10687 (N_10687,N_10524,N_10437);
nand U10688 (N_10688,N_10482,N_10432);
nand U10689 (N_10689,N_10428,N_10458);
nand U10690 (N_10690,N_10497,N_10549);
nor U10691 (N_10691,N_10401,N_10407);
nor U10692 (N_10692,N_10452,N_10555);
or U10693 (N_10693,N_10446,N_10408);
nand U10694 (N_10694,N_10484,N_10420);
and U10695 (N_10695,N_10452,N_10414);
and U10696 (N_10696,N_10472,N_10499);
nor U10697 (N_10697,N_10411,N_10547);
or U10698 (N_10698,N_10541,N_10479);
and U10699 (N_10699,N_10489,N_10480);
and U10700 (N_10700,N_10430,N_10445);
xor U10701 (N_10701,N_10536,N_10433);
nand U10702 (N_10702,N_10493,N_10487);
or U10703 (N_10703,N_10534,N_10442);
nor U10704 (N_10704,N_10442,N_10477);
and U10705 (N_10705,N_10495,N_10486);
and U10706 (N_10706,N_10524,N_10480);
or U10707 (N_10707,N_10518,N_10445);
and U10708 (N_10708,N_10464,N_10465);
nand U10709 (N_10709,N_10549,N_10410);
and U10710 (N_10710,N_10491,N_10409);
or U10711 (N_10711,N_10433,N_10445);
nand U10712 (N_10712,N_10488,N_10535);
xnor U10713 (N_10713,N_10457,N_10526);
xor U10714 (N_10714,N_10480,N_10452);
and U10715 (N_10715,N_10506,N_10466);
or U10716 (N_10716,N_10473,N_10502);
nand U10717 (N_10717,N_10404,N_10421);
nor U10718 (N_10718,N_10419,N_10447);
xnor U10719 (N_10719,N_10512,N_10446);
or U10720 (N_10720,N_10569,N_10581);
and U10721 (N_10721,N_10627,N_10639);
nand U10722 (N_10722,N_10573,N_10629);
or U10723 (N_10723,N_10649,N_10718);
xnor U10724 (N_10724,N_10621,N_10689);
nand U10725 (N_10725,N_10697,N_10575);
xor U10726 (N_10726,N_10567,N_10713);
nand U10727 (N_10727,N_10626,N_10669);
nor U10728 (N_10728,N_10591,N_10623);
nor U10729 (N_10729,N_10578,N_10609);
nor U10730 (N_10730,N_10692,N_10565);
nand U10731 (N_10731,N_10696,N_10657);
or U10732 (N_10732,N_10600,N_10691);
xnor U10733 (N_10733,N_10704,N_10579);
nand U10734 (N_10734,N_10676,N_10642);
or U10735 (N_10735,N_10717,N_10641);
or U10736 (N_10736,N_10615,N_10614);
nand U10737 (N_10737,N_10708,N_10570);
nor U10738 (N_10738,N_10606,N_10706);
xor U10739 (N_10739,N_10571,N_10564);
nor U10740 (N_10740,N_10563,N_10598);
xnor U10741 (N_10741,N_10656,N_10572);
or U10742 (N_10742,N_10643,N_10577);
or U10743 (N_10743,N_10667,N_10599);
xor U10744 (N_10744,N_10635,N_10701);
or U10745 (N_10745,N_10703,N_10677);
xor U10746 (N_10746,N_10678,N_10576);
xnor U10747 (N_10747,N_10680,N_10624);
nand U10748 (N_10748,N_10647,N_10601);
xor U10749 (N_10749,N_10584,N_10674);
and U10750 (N_10750,N_10662,N_10588);
nor U10751 (N_10751,N_10640,N_10589);
and U10752 (N_10752,N_10638,N_10670);
or U10753 (N_10753,N_10597,N_10688);
nand U10754 (N_10754,N_10580,N_10664);
or U10755 (N_10755,N_10709,N_10710);
nand U10756 (N_10756,N_10566,N_10604);
nor U10757 (N_10757,N_10716,N_10613);
xnor U10758 (N_10758,N_10585,N_10594);
xnor U10759 (N_10759,N_10634,N_10561);
xnor U10760 (N_10760,N_10684,N_10690);
and U10761 (N_10761,N_10616,N_10665);
or U10762 (N_10762,N_10574,N_10582);
or U10763 (N_10763,N_10686,N_10602);
xor U10764 (N_10764,N_10661,N_10611);
and U10765 (N_10765,N_10707,N_10630);
or U10766 (N_10766,N_10659,N_10622);
or U10767 (N_10767,N_10653,N_10645);
or U10768 (N_10768,N_10632,N_10694);
or U10769 (N_10769,N_10612,N_10673);
nand U10770 (N_10770,N_10628,N_10655);
xor U10771 (N_10771,N_10633,N_10668);
xor U10772 (N_10772,N_10671,N_10714);
nor U10773 (N_10773,N_10595,N_10675);
nand U10774 (N_10774,N_10650,N_10715);
and U10775 (N_10775,N_10637,N_10654);
or U10776 (N_10776,N_10651,N_10618);
and U10777 (N_10777,N_10719,N_10663);
nand U10778 (N_10778,N_10695,N_10687);
nor U10779 (N_10779,N_10605,N_10607);
nand U10780 (N_10780,N_10693,N_10592);
nor U10781 (N_10781,N_10712,N_10700);
nor U10782 (N_10782,N_10658,N_10648);
xnor U10783 (N_10783,N_10593,N_10562);
or U10784 (N_10784,N_10702,N_10685);
or U10785 (N_10785,N_10636,N_10666);
and U10786 (N_10786,N_10610,N_10619);
and U10787 (N_10787,N_10682,N_10560);
and U10788 (N_10788,N_10590,N_10568);
and U10789 (N_10789,N_10672,N_10620);
nor U10790 (N_10790,N_10644,N_10705);
xor U10791 (N_10791,N_10679,N_10698);
or U10792 (N_10792,N_10583,N_10603);
or U10793 (N_10793,N_10652,N_10586);
or U10794 (N_10794,N_10596,N_10646);
or U10795 (N_10795,N_10617,N_10683);
nand U10796 (N_10796,N_10699,N_10608);
xor U10797 (N_10797,N_10660,N_10587);
xor U10798 (N_10798,N_10625,N_10631);
xor U10799 (N_10799,N_10681,N_10711);
xnor U10800 (N_10800,N_10713,N_10637);
nor U10801 (N_10801,N_10589,N_10711);
and U10802 (N_10802,N_10611,N_10659);
nor U10803 (N_10803,N_10711,N_10612);
or U10804 (N_10804,N_10631,N_10669);
xnor U10805 (N_10805,N_10707,N_10585);
nor U10806 (N_10806,N_10666,N_10610);
nor U10807 (N_10807,N_10597,N_10677);
and U10808 (N_10808,N_10566,N_10584);
nor U10809 (N_10809,N_10645,N_10690);
nand U10810 (N_10810,N_10651,N_10626);
nand U10811 (N_10811,N_10684,N_10603);
or U10812 (N_10812,N_10613,N_10582);
nand U10813 (N_10813,N_10593,N_10621);
nor U10814 (N_10814,N_10704,N_10610);
nor U10815 (N_10815,N_10566,N_10692);
nor U10816 (N_10816,N_10681,N_10651);
and U10817 (N_10817,N_10683,N_10707);
or U10818 (N_10818,N_10602,N_10637);
or U10819 (N_10819,N_10645,N_10713);
xnor U10820 (N_10820,N_10607,N_10691);
or U10821 (N_10821,N_10684,N_10608);
nand U10822 (N_10822,N_10599,N_10592);
nor U10823 (N_10823,N_10655,N_10573);
xnor U10824 (N_10824,N_10684,N_10680);
or U10825 (N_10825,N_10718,N_10703);
xnor U10826 (N_10826,N_10562,N_10692);
nand U10827 (N_10827,N_10617,N_10597);
nand U10828 (N_10828,N_10678,N_10631);
or U10829 (N_10829,N_10629,N_10593);
xnor U10830 (N_10830,N_10649,N_10575);
and U10831 (N_10831,N_10574,N_10719);
and U10832 (N_10832,N_10592,N_10618);
nand U10833 (N_10833,N_10561,N_10606);
xnor U10834 (N_10834,N_10634,N_10596);
xor U10835 (N_10835,N_10702,N_10696);
nor U10836 (N_10836,N_10581,N_10578);
nor U10837 (N_10837,N_10702,N_10670);
nor U10838 (N_10838,N_10613,N_10605);
or U10839 (N_10839,N_10684,N_10631);
nand U10840 (N_10840,N_10680,N_10604);
nand U10841 (N_10841,N_10678,N_10652);
xor U10842 (N_10842,N_10700,N_10678);
nand U10843 (N_10843,N_10694,N_10666);
and U10844 (N_10844,N_10704,N_10671);
nand U10845 (N_10845,N_10627,N_10576);
nor U10846 (N_10846,N_10706,N_10593);
xor U10847 (N_10847,N_10588,N_10647);
nor U10848 (N_10848,N_10611,N_10600);
and U10849 (N_10849,N_10644,N_10659);
or U10850 (N_10850,N_10622,N_10664);
xnor U10851 (N_10851,N_10604,N_10584);
nor U10852 (N_10852,N_10604,N_10682);
xnor U10853 (N_10853,N_10714,N_10620);
and U10854 (N_10854,N_10651,N_10656);
and U10855 (N_10855,N_10708,N_10632);
nor U10856 (N_10856,N_10591,N_10595);
and U10857 (N_10857,N_10670,N_10678);
or U10858 (N_10858,N_10714,N_10643);
and U10859 (N_10859,N_10601,N_10635);
xnor U10860 (N_10860,N_10709,N_10676);
nor U10861 (N_10861,N_10664,N_10647);
and U10862 (N_10862,N_10609,N_10613);
or U10863 (N_10863,N_10702,N_10597);
nor U10864 (N_10864,N_10640,N_10648);
or U10865 (N_10865,N_10582,N_10715);
nand U10866 (N_10866,N_10671,N_10632);
or U10867 (N_10867,N_10603,N_10697);
or U10868 (N_10868,N_10688,N_10602);
and U10869 (N_10869,N_10715,N_10561);
xor U10870 (N_10870,N_10561,N_10580);
xor U10871 (N_10871,N_10601,N_10582);
or U10872 (N_10872,N_10669,N_10586);
and U10873 (N_10873,N_10598,N_10583);
nand U10874 (N_10874,N_10694,N_10674);
nand U10875 (N_10875,N_10655,N_10713);
or U10876 (N_10876,N_10577,N_10670);
nand U10877 (N_10877,N_10682,N_10673);
xnor U10878 (N_10878,N_10609,N_10662);
nor U10879 (N_10879,N_10639,N_10564);
and U10880 (N_10880,N_10846,N_10868);
and U10881 (N_10881,N_10809,N_10748);
nand U10882 (N_10882,N_10832,N_10826);
nor U10883 (N_10883,N_10857,N_10842);
or U10884 (N_10884,N_10856,N_10736);
or U10885 (N_10885,N_10851,N_10739);
nor U10886 (N_10886,N_10738,N_10755);
or U10887 (N_10887,N_10729,N_10835);
xnor U10888 (N_10888,N_10721,N_10830);
xor U10889 (N_10889,N_10848,N_10818);
xnor U10890 (N_10890,N_10795,N_10840);
or U10891 (N_10891,N_10811,N_10794);
nor U10892 (N_10892,N_10810,N_10754);
nand U10893 (N_10893,N_10749,N_10775);
nor U10894 (N_10894,N_10841,N_10825);
or U10895 (N_10895,N_10878,N_10798);
and U10896 (N_10896,N_10780,N_10759);
nor U10897 (N_10897,N_10859,N_10860);
or U10898 (N_10898,N_10735,N_10787);
or U10899 (N_10899,N_10763,N_10764);
nand U10900 (N_10900,N_10854,N_10769);
and U10901 (N_10901,N_10731,N_10804);
or U10902 (N_10902,N_10720,N_10761);
and U10903 (N_10903,N_10766,N_10740);
nand U10904 (N_10904,N_10872,N_10765);
xnor U10905 (N_10905,N_10803,N_10849);
or U10906 (N_10906,N_10870,N_10762);
xor U10907 (N_10907,N_10844,N_10876);
nor U10908 (N_10908,N_10820,N_10789);
or U10909 (N_10909,N_10728,N_10732);
xor U10910 (N_10910,N_10799,N_10836);
nand U10911 (N_10911,N_10858,N_10744);
nand U10912 (N_10912,N_10772,N_10837);
nand U10913 (N_10913,N_10779,N_10785);
xnor U10914 (N_10914,N_10808,N_10867);
and U10915 (N_10915,N_10737,N_10816);
and U10916 (N_10916,N_10833,N_10853);
xnor U10917 (N_10917,N_10805,N_10861);
xnor U10918 (N_10918,N_10864,N_10750);
nand U10919 (N_10919,N_10722,N_10733);
and U10920 (N_10920,N_10824,N_10768);
nand U10921 (N_10921,N_10797,N_10869);
nand U10922 (N_10922,N_10777,N_10725);
nand U10923 (N_10923,N_10852,N_10806);
xnor U10924 (N_10924,N_10745,N_10855);
or U10925 (N_10925,N_10843,N_10800);
nor U10926 (N_10926,N_10845,N_10741);
and U10927 (N_10927,N_10817,N_10863);
nand U10928 (N_10928,N_10742,N_10819);
xnor U10929 (N_10929,N_10839,N_10726);
xor U10930 (N_10930,N_10847,N_10814);
or U10931 (N_10931,N_10791,N_10758);
xor U10932 (N_10932,N_10774,N_10724);
and U10933 (N_10933,N_10828,N_10784);
xor U10934 (N_10934,N_10815,N_10778);
or U10935 (N_10935,N_10792,N_10751);
xnor U10936 (N_10936,N_10874,N_10862);
and U10937 (N_10937,N_10822,N_10875);
and U10938 (N_10938,N_10866,N_10813);
nor U10939 (N_10939,N_10788,N_10873);
nor U10940 (N_10940,N_10801,N_10879);
xor U10941 (N_10941,N_10757,N_10821);
nor U10942 (N_10942,N_10723,N_10783);
and U10943 (N_10943,N_10770,N_10756);
or U10944 (N_10944,N_10850,N_10752);
and U10945 (N_10945,N_10812,N_10773);
xnor U10946 (N_10946,N_10760,N_10734);
xnor U10947 (N_10947,N_10827,N_10786);
nor U10948 (N_10948,N_10782,N_10871);
nand U10949 (N_10949,N_10747,N_10793);
nand U10950 (N_10950,N_10781,N_10727);
nand U10951 (N_10951,N_10796,N_10865);
xnor U10952 (N_10952,N_10834,N_10877);
xnor U10953 (N_10953,N_10807,N_10829);
nand U10954 (N_10954,N_10831,N_10771);
or U10955 (N_10955,N_10753,N_10767);
xor U10956 (N_10956,N_10776,N_10730);
and U10957 (N_10957,N_10838,N_10823);
xnor U10958 (N_10958,N_10790,N_10746);
or U10959 (N_10959,N_10743,N_10802);
and U10960 (N_10960,N_10810,N_10847);
nor U10961 (N_10961,N_10763,N_10829);
and U10962 (N_10962,N_10737,N_10724);
or U10963 (N_10963,N_10787,N_10807);
xnor U10964 (N_10964,N_10724,N_10772);
or U10965 (N_10965,N_10731,N_10790);
nand U10966 (N_10966,N_10754,N_10747);
nand U10967 (N_10967,N_10865,N_10743);
and U10968 (N_10968,N_10875,N_10818);
or U10969 (N_10969,N_10820,N_10819);
nand U10970 (N_10970,N_10720,N_10722);
xnor U10971 (N_10971,N_10798,N_10800);
nand U10972 (N_10972,N_10864,N_10816);
nand U10973 (N_10973,N_10768,N_10736);
and U10974 (N_10974,N_10862,N_10766);
or U10975 (N_10975,N_10749,N_10792);
nand U10976 (N_10976,N_10855,N_10848);
and U10977 (N_10977,N_10813,N_10791);
nor U10978 (N_10978,N_10816,N_10789);
nor U10979 (N_10979,N_10850,N_10732);
xor U10980 (N_10980,N_10820,N_10832);
or U10981 (N_10981,N_10858,N_10756);
xnor U10982 (N_10982,N_10729,N_10808);
nor U10983 (N_10983,N_10844,N_10854);
nand U10984 (N_10984,N_10846,N_10812);
xor U10985 (N_10985,N_10782,N_10836);
nand U10986 (N_10986,N_10782,N_10746);
nor U10987 (N_10987,N_10723,N_10721);
or U10988 (N_10988,N_10874,N_10777);
nor U10989 (N_10989,N_10814,N_10744);
nand U10990 (N_10990,N_10730,N_10746);
nand U10991 (N_10991,N_10738,N_10763);
or U10992 (N_10992,N_10833,N_10775);
nand U10993 (N_10993,N_10745,N_10793);
xor U10994 (N_10994,N_10855,N_10793);
and U10995 (N_10995,N_10832,N_10737);
nand U10996 (N_10996,N_10874,N_10805);
xor U10997 (N_10997,N_10721,N_10789);
xor U10998 (N_10998,N_10822,N_10770);
xor U10999 (N_10999,N_10753,N_10874);
nand U11000 (N_11000,N_10782,N_10761);
xnor U11001 (N_11001,N_10849,N_10848);
nor U11002 (N_11002,N_10815,N_10785);
and U11003 (N_11003,N_10729,N_10873);
xnor U11004 (N_11004,N_10780,N_10754);
nand U11005 (N_11005,N_10732,N_10753);
xor U11006 (N_11006,N_10753,N_10836);
or U11007 (N_11007,N_10795,N_10747);
and U11008 (N_11008,N_10732,N_10756);
xor U11009 (N_11009,N_10831,N_10806);
or U11010 (N_11010,N_10837,N_10730);
and U11011 (N_11011,N_10800,N_10833);
nand U11012 (N_11012,N_10732,N_10763);
nor U11013 (N_11013,N_10850,N_10820);
nor U11014 (N_11014,N_10741,N_10739);
xor U11015 (N_11015,N_10720,N_10870);
and U11016 (N_11016,N_10824,N_10811);
nand U11017 (N_11017,N_10787,N_10804);
nand U11018 (N_11018,N_10851,N_10785);
or U11019 (N_11019,N_10777,N_10815);
xor U11020 (N_11020,N_10831,N_10736);
and U11021 (N_11021,N_10808,N_10778);
nand U11022 (N_11022,N_10836,N_10742);
xnor U11023 (N_11023,N_10871,N_10749);
nand U11024 (N_11024,N_10754,N_10876);
xnor U11025 (N_11025,N_10864,N_10792);
nor U11026 (N_11026,N_10755,N_10732);
or U11027 (N_11027,N_10779,N_10818);
nand U11028 (N_11028,N_10730,N_10844);
or U11029 (N_11029,N_10804,N_10777);
and U11030 (N_11030,N_10760,N_10822);
nor U11031 (N_11031,N_10765,N_10738);
xor U11032 (N_11032,N_10819,N_10743);
or U11033 (N_11033,N_10825,N_10745);
or U11034 (N_11034,N_10788,N_10849);
nand U11035 (N_11035,N_10828,N_10847);
nor U11036 (N_11036,N_10867,N_10796);
nor U11037 (N_11037,N_10782,N_10803);
or U11038 (N_11038,N_10774,N_10729);
xor U11039 (N_11039,N_10750,N_10748);
and U11040 (N_11040,N_11013,N_10883);
and U11041 (N_11041,N_10977,N_10953);
nand U11042 (N_11042,N_11001,N_10971);
nand U11043 (N_11043,N_10887,N_10969);
and U11044 (N_11044,N_10891,N_10893);
and U11045 (N_11045,N_11035,N_10921);
or U11046 (N_11046,N_10986,N_11022);
xor U11047 (N_11047,N_10982,N_10890);
or U11048 (N_11048,N_11016,N_10915);
xor U11049 (N_11049,N_10892,N_10929);
and U11050 (N_11050,N_10918,N_10980);
nor U11051 (N_11051,N_10895,N_11026);
nor U11052 (N_11052,N_10912,N_10973);
or U11053 (N_11053,N_10936,N_10974);
and U11054 (N_11054,N_10884,N_11007);
xor U11055 (N_11055,N_10984,N_10940);
or U11056 (N_11056,N_10939,N_10968);
nand U11057 (N_11057,N_11002,N_11038);
and U11058 (N_11058,N_10933,N_10899);
nor U11059 (N_11059,N_11000,N_10950);
nor U11060 (N_11060,N_11018,N_10901);
nor U11061 (N_11061,N_10956,N_11030);
or U11062 (N_11062,N_10978,N_10945);
and U11063 (N_11063,N_10927,N_10994);
and U11064 (N_11064,N_10996,N_10967);
nand U11065 (N_11065,N_10910,N_10952);
or U11066 (N_11066,N_10880,N_10905);
or U11067 (N_11067,N_10926,N_11027);
nor U11068 (N_11068,N_10897,N_10907);
nor U11069 (N_11069,N_10985,N_10987);
nand U11070 (N_11070,N_10917,N_10894);
xnor U11071 (N_11071,N_10970,N_10920);
nor U11072 (N_11072,N_10923,N_10944);
and U11073 (N_11073,N_10922,N_10916);
and U11074 (N_11074,N_10934,N_10911);
nor U11075 (N_11075,N_11032,N_10966);
and U11076 (N_11076,N_11025,N_10941);
nand U11077 (N_11077,N_10998,N_10991);
nand U11078 (N_11078,N_10903,N_10924);
and U11079 (N_11079,N_10914,N_10947);
nor U11080 (N_11080,N_11021,N_11015);
nor U11081 (N_11081,N_11024,N_10930);
or U11082 (N_11082,N_10881,N_10896);
nor U11083 (N_11083,N_11004,N_10949);
nor U11084 (N_11084,N_10989,N_10932);
xor U11085 (N_11085,N_10904,N_10938);
nand U11086 (N_11086,N_10992,N_10963);
and U11087 (N_11087,N_11031,N_10898);
nand U11088 (N_11088,N_10931,N_10960);
and U11089 (N_11089,N_11005,N_10888);
and U11090 (N_11090,N_10993,N_10906);
or U11091 (N_11091,N_10885,N_11034);
xnor U11092 (N_11092,N_10964,N_10975);
and U11093 (N_11093,N_11029,N_10942);
xor U11094 (N_11094,N_10902,N_10955);
and U11095 (N_11095,N_10928,N_10948);
nor U11096 (N_11096,N_10954,N_11017);
and U11097 (N_11097,N_10961,N_10900);
xnor U11098 (N_11098,N_11014,N_10962);
or U11099 (N_11099,N_11003,N_10965);
xnor U11100 (N_11100,N_10958,N_11019);
and U11101 (N_11101,N_10919,N_10935);
nor U11102 (N_11102,N_11036,N_10886);
and U11103 (N_11103,N_10981,N_10988);
nor U11104 (N_11104,N_11006,N_10997);
xnor U11105 (N_11105,N_11028,N_10946);
and U11106 (N_11106,N_11020,N_11010);
or U11107 (N_11107,N_11012,N_11023);
or U11108 (N_11108,N_10951,N_10990);
and U11109 (N_11109,N_11039,N_11037);
xnor U11110 (N_11110,N_10943,N_10983);
nor U11111 (N_11111,N_10913,N_10908);
and U11112 (N_11112,N_11008,N_10972);
or U11113 (N_11113,N_10959,N_10995);
and U11114 (N_11114,N_10937,N_11033);
nor U11115 (N_11115,N_11009,N_10909);
xnor U11116 (N_11116,N_10979,N_10925);
and U11117 (N_11117,N_10882,N_10957);
nand U11118 (N_11118,N_10999,N_11011);
nand U11119 (N_11119,N_10976,N_10889);
nor U11120 (N_11120,N_11023,N_11016);
nand U11121 (N_11121,N_10898,N_10959);
and U11122 (N_11122,N_10958,N_10922);
or U11123 (N_11123,N_10961,N_10908);
nor U11124 (N_11124,N_10898,N_10970);
nor U11125 (N_11125,N_10903,N_10949);
and U11126 (N_11126,N_11023,N_11039);
xnor U11127 (N_11127,N_11008,N_10913);
and U11128 (N_11128,N_10880,N_10985);
and U11129 (N_11129,N_10966,N_11011);
nor U11130 (N_11130,N_10889,N_10910);
nor U11131 (N_11131,N_11027,N_10896);
nor U11132 (N_11132,N_10989,N_11007);
nand U11133 (N_11133,N_10961,N_10944);
or U11134 (N_11134,N_11027,N_10887);
nand U11135 (N_11135,N_10946,N_10912);
or U11136 (N_11136,N_10964,N_10905);
nand U11137 (N_11137,N_10945,N_10910);
and U11138 (N_11138,N_10943,N_10882);
and U11139 (N_11139,N_11035,N_11002);
nand U11140 (N_11140,N_10994,N_10973);
or U11141 (N_11141,N_10999,N_11018);
nor U11142 (N_11142,N_10937,N_10921);
and U11143 (N_11143,N_11008,N_11006);
nand U11144 (N_11144,N_11014,N_11022);
nor U11145 (N_11145,N_11017,N_10904);
nor U11146 (N_11146,N_10885,N_10987);
nand U11147 (N_11147,N_10935,N_10973);
xor U11148 (N_11148,N_10956,N_10890);
xnor U11149 (N_11149,N_10911,N_11024);
nor U11150 (N_11150,N_10925,N_10909);
nand U11151 (N_11151,N_10888,N_11015);
and U11152 (N_11152,N_11017,N_11039);
and U11153 (N_11153,N_11019,N_10900);
nor U11154 (N_11154,N_10930,N_10931);
or U11155 (N_11155,N_10914,N_10897);
or U11156 (N_11156,N_11021,N_11009);
nor U11157 (N_11157,N_10909,N_11039);
nor U11158 (N_11158,N_10942,N_10903);
nand U11159 (N_11159,N_10946,N_10971);
and U11160 (N_11160,N_10967,N_10943);
and U11161 (N_11161,N_10944,N_10927);
nor U11162 (N_11162,N_10977,N_10952);
xnor U11163 (N_11163,N_11031,N_11012);
nand U11164 (N_11164,N_10929,N_10982);
nand U11165 (N_11165,N_10983,N_11012);
or U11166 (N_11166,N_11030,N_11003);
or U11167 (N_11167,N_10914,N_11034);
xnor U11168 (N_11168,N_11006,N_10982);
nand U11169 (N_11169,N_11009,N_10895);
nand U11170 (N_11170,N_10881,N_10977);
nor U11171 (N_11171,N_10978,N_10963);
or U11172 (N_11172,N_10975,N_11033);
or U11173 (N_11173,N_11011,N_10925);
xnor U11174 (N_11174,N_10890,N_10976);
and U11175 (N_11175,N_10984,N_10947);
nor U11176 (N_11176,N_10963,N_10935);
nand U11177 (N_11177,N_10968,N_11029);
xor U11178 (N_11178,N_10949,N_10953);
nand U11179 (N_11179,N_10920,N_11030);
xor U11180 (N_11180,N_10935,N_10888);
and U11181 (N_11181,N_11036,N_10943);
nand U11182 (N_11182,N_11024,N_10988);
nand U11183 (N_11183,N_10890,N_11001);
nand U11184 (N_11184,N_10987,N_10936);
or U11185 (N_11185,N_11010,N_11014);
nor U11186 (N_11186,N_10931,N_10967);
nor U11187 (N_11187,N_10928,N_11029);
or U11188 (N_11188,N_10951,N_11020);
and U11189 (N_11189,N_10897,N_10921);
and U11190 (N_11190,N_11002,N_10983);
nand U11191 (N_11191,N_10958,N_10972);
nand U11192 (N_11192,N_10902,N_10980);
nor U11193 (N_11193,N_10957,N_10963);
or U11194 (N_11194,N_10933,N_11008);
nor U11195 (N_11195,N_10881,N_10942);
nor U11196 (N_11196,N_10898,N_10892);
or U11197 (N_11197,N_10895,N_10923);
and U11198 (N_11198,N_10940,N_10990);
nor U11199 (N_11199,N_11016,N_10941);
nand U11200 (N_11200,N_11081,N_11127);
and U11201 (N_11201,N_11142,N_11106);
or U11202 (N_11202,N_11077,N_11110);
nor U11203 (N_11203,N_11088,N_11190);
and U11204 (N_11204,N_11070,N_11073);
nand U11205 (N_11205,N_11129,N_11114);
nor U11206 (N_11206,N_11109,N_11082);
nand U11207 (N_11207,N_11158,N_11199);
nor U11208 (N_11208,N_11093,N_11125);
nand U11209 (N_11209,N_11052,N_11163);
xnor U11210 (N_11210,N_11122,N_11167);
and U11211 (N_11211,N_11054,N_11173);
and U11212 (N_11212,N_11099,N_11188);
and U11213 (N_11213,N_11183,N_11041);
nor U11214 (N_11214,N_11195,N_11162);
nand U11215 (N_11215,N_11112,N_11172);
or U11216 (N_11216,N_11150,N_11168);
nand U11217 (N_11217,N_11056,N_11059);
nand U11218 (N_11218,N_11108,N_11133);
xor U11219 (N_11219,N_11102,N_11107);
and U11220 (N_11220,N_11148,N_11089);
nand U11221 (N_11221,N_11050,N_11184);
nand U11222 (N_11222,N_11058,N_11064);
or U11223 (N_11223,N_11130,N_11040);
or U11224 (N_11224,N_11189,N_11042);
and U11225 (N_11225,N_11111,N_11147);
or U11226 (N_11226,N_11078,N_11103);
and U11227 (N_11227,N_11047,N_11105);
and U11228 (N_11228,N_11159,N_11098);
xnor U11229 (N_11229,N_11079,N_11123);
xnor U11230 (N_11230,N_11194,N_11179);
and U11231 (N_11231,N_11174,N_11063);
and U11232 (N_11232,N_11180,N_11053);
nor U11233 (N_11233,N_11115,N_11138);
nand U11234 (N_11234,N_11141,N_11156);
and U11235 (N_11235,N_11043,N_11196);
or U11236 (N_11236,N_11157,N_11090);
nand U11237 (N_11237,N_11071,N_11149);
or U11238 (N_11238,N_11057,N_11140);
and U11239 (N_11239,N_11074,N_11134);
xnor U11240 (N_11240,N_11067,N_11072);
xnor U11241 (N_11241,N_11083,N_11061);
xor U11242 (N_11242,N_11197,N_11060);
and U11243 (N_11243,N_11169,N_11068);
nor U11244 (N_11244,N_11121,N_11066);
nor U11245 (N_11245,N_11143,N_11131);
nand U11246 (N_11246,N_11161,N_11119);
or U11247 (N_11247,N_11062,N_11155);
or U11248 (N_11248,N_11154,N_11175);
nand U11249 (N_11249,N_11124,N_11132);
nand U11250 (N_11250,N_11193,N_11049);
nor U11251 (N_11251,N_11046,N_11087);
or U11252 (N_11252,N_11091,N_11095);
and U11253 (N_11253,N_11187,N_11139);
and U11254 (N_11254,N_11186,N_11181);
and U11255 (N_11255,N_11045,N_11152);
nor U11256 (N_11256,N_11136,N_11113);
nor U11257 (N_11257,N_11065,N_11044);
nand U11258 (N_11258,N_11104,N_11094);
nor U11259 (N_11259,N_11145,N_11126);
or U11260 (N_11260,N_11137,N_11084);
and U11261 (N_11261,N_11198,N_11176);
xor U11262 (N_11262,N_11166,N_11100);
nand U11263 (N_11263,N_11076,N_11055);
nand U11264 (N_11264,N_11144,N_11075);
nor U11265 (N_11265,N_11117,N_11101);
nand U11266 (N_11266,N_11178,N_11085);
and U11267 (N_11267,N_11151,N_11069);
or U11268 (N_11268,N_11160,N_11165);
or U11269 (N_11269,N_11086,N_11146);
and U11270 (N_11270,N_11080,N_11185);
or U11271 (N_11271,N_11096,N_11116);
nand U11272 (N_11272,N_11192,N_11051);
and U11273 (N_11273,N_11170,N_11128);
or U11274 (N_11274,N_11097,N_11118);
xnor U11275 (N_11275,N_11191,N_11120);
nand U11276 (N_11276,N_11092,N_11171);
and U11277 (N_11277,N_11177,N_11182);
nor U11278 (N_11278,N_11048,N_11164);
nand U11279 (N_11279,N_11153,N_11135);
xor U11280 (N_11280,N_11187,N_11066);
nor U11281 (N_11281,N_11140,N_11170);
nor U11282 (N_11282,N_11066,N_11158);
nand U11283 (N_11283,N_11112,N_11134);
or U11284 (N_11284,N_11046,N_11125);
nand U11285 (N_11285,N_11081,N_11093);
nand U11286 (N_11286,N_11147,N_11066);
and U11287 (N_11287,N_11147,N_11043);
nor U11288 (N_11288,N_11080,N_11061);
nor U11289 (N_11289,N_11133,N_11190);
or U11290 (N_11290,N_11089,N_11123);
nor U11291 (N_11291,N_11041,N_11099);
xnor U11292 (N_11292,N_11102,N_11091);
and U11293 (N_11293,N_11065,N_11110);
nor U11294 (N_11294,N_11136,N_11151);
xor U11295 (N_11295,N_11155,N_11189);
and U11296 (N_11296,N_11057,N_11172);
and U11297 (N_11297,N_11152,N_11172);
or U11298 (N_11298,N_11120,N_11143);
or U11299 (N_11299,N_11187,N_11189);
and U11300 (N_11300,N_11068,N_11190);
nor U11301 (N_11301,N_11141,N_11153);
or U11302 (N_11302,N_11137,N_11111);
or U11303 (N_11303,N_11196,N_11129);
nor U11304 (N_11304,N_11158,N_11172);
nor U11305 (N_11305,N_11173,N_11109);
or U11306 (N_11306,N_11197,N_11068);
and U11307 (N_11307,N_11107,N_11153);
or U11308 (N_11308,N_11093,N_11134);
nand U11309 (N_11309,N_11192,N_11148);
or U11310 (N_11310,N_11136,N_11164);
or U11311 (N_11311,N_11146,N_11059);
nand U11312 (N_11312,N_11131,N_11102);
xor U11313 (N_11313,N_11040,N_11051);
and U11314 (N_11314,N_11105,N_11076);
nor U11315 (N_11315,N_11185,N_11079);
nand U11316 (N_11316,N_11071,N_11192);
xor U11317 (N_11317,N_11177,N_11179);
xnor U11318 (N_11318,N_11052,N_11065);
nand U11319 (N_11319,N_11191,N_11165);
nand U11320 (N_11320,N_11144,N_11112);
or U11321 (N_11321,N_11043,N_11117);
nor U11322 (N_11322,N_11164,N_11171);
and U11323 (N_11323,N_11179,N_11170);
or U11324 (N_11324,N_11100,N_11156);
xnor U11325 (N_11325,N_11116,N_11127);
and U11326 (N_11326,N_11167,N_11078);
or U11327 (N_11327,N_11088,N_11059);
or U11328 (N_11328,N_11145,N_11161);
xor U11329 (N_11329,N_11044,N_11179);
or U11330 (N_11330,N_11186,N_11084);
or U11331 (N_11331,N_11172,N_11134);
and U11332 (N_11332,N_11087,N_11054);
nor U11333 (N_11333,N_11157,N_11061);
or U11334 (N_11334,N_11123,N_11076);
nand U11335 (N_11335,N_11143,N_11164);
and U11336 (N_11336,N_11152,N_11089);
or U11337 (N_11337,N_11070,N_11163);
and U11338 (N_11338,N_11158,N_11109);
and U11339 (N_11339,N_11149,N_11107);
xnor U11340 (N_11340,N_11168,N_11141);
or U11341 (N_11341,N_11135,N_11081);
nor U11342 (N_11342,N_11117,N_11089);
or U11343 (N_11343,N_11088,N_11127);
nor U11344 (N_11344,N_11054,N_11137);
or U11345 (N_11345,N_11118,N_11148);
xnor U11346 (N_11346,N_11057,N_11124);
xor U11347 (N_11347,N_11117,N_11198);
nor U11348 (N_11348,N_11153,N_11145);
xor U11349 (N_11349,N_11195,N_11164);
or U11350 (N_11350,N_11073,N_11049);
or U11351 (N_11351,N_11050,N_11071);
xnor U11352 (N_11352,N_11196,N_11199);
or U11353 (N_11353,N_11158,N_11133);
nor U11354 (N_11354,N_11134,N_11136);
or U11355 (N_11355,N_11171,N_11110);
nand U11356 (N_11356,N_11175,N_11158);
nor U11357 (N_11357,N_11105,N_11142);
or U11358 (N_11358,N_11158,N_11140);
nor U11359 (N_11359,N_11143,N_11062);
nor U11360 (N_11360,N_11322,N_11330);
or U11361 (N_11361,N_11255,N_11319);
and U11362 (N_11362,N_11347,N_11251);
nand U11363 (N_11363,N_11301,N_11265);
or U11364 (N_11364,N_11341,N_11356);
and U11365 (N_11365,N_11208,N_11200);
and U11366 (N_11366,N_11267,N_11309);
nand U11367 (N_11367,N_11323,N_11256);
or U11368 (N_11368,N_11226,N_11333);
or U11369 (N_11369,N_11314,N_11324);
and U11370 (N_11370,N_11291,N_11282);
and U11371 (N_11371,N_11338,N_11293);
or U11372 (N_11372,N_11216,N_11295);
nand U11373 (N_11373,N_11296,N_11339);
or U11374 (N_11374,N_11286,N_11212);
or U11375 (N_11375,N_11266,N_11275);
or U11376 (N_11376,N_11239,N_11305);
nor U11377 (N_11377,N_11261,N_11272);
and U11378 (N_11378,N_11229,N_11355);
xnor U11379 (N_11379,N_11289,N_11277);
or U11380 (N_11380,N_11318,N_11202);
nand U11381 (N_11381,N_11235,N_11351);
and U11382 (N_11382,N_11335,N_11237);
nand U11383 (N_11383,N_11273,N_11352);
xor U11384 (N_11384,N_11358,N_11240);
nand U11385 (N_11385,N_11274,N_11346);
or U11386 (N_11386,N_11221,N_11328);
and U11387 (N_11387,N_11278,N_11292);
nor U11388 (N_11388,N_11234,N_11252);
or U11389 (N_11389,N_11340,N_11349);
nor U11390 (N_11390,N_11313,N_11262);
nand U11391 (N_11391,N_11231,N_11317);
and U11392 (N_11392,N_11308,N_11270);
and U11393 (N_11393,N_11225,N_11236);
nand U11394 (N_11394,N_11294,N_11345);
xnor U11395 (N_11395,N_11332,N_11222);
and U11396 (N_11396,N_11213,N_11331);
xnor U11397 (N_11397,N_11211,N_11268);
and U11398 (N_11398,N_11257,N_11253);
xnor U11399 (N_11399,N_11219,N_11300);
nor U11400 (N_11400,N_11205,N_11312);
and U11401 (N_11401,N_11280,N_11223);
or U11402 (N_11402,N_11203,N_11204);
xor U11403 (N_11403,N_11241,N_11350);
nor U11404 (N_11404,N_11247,N_11343);
xor U11405 (N_11405,N_11238,N_11230);
xnor U11406 (N_11406,N_11243,N_11327);
or U11407 (N_11407,N_11337,N_11326);
or U11408 (N_11408,N_11285,N_11250);
xnor U11409 (N_11409,N_11310,N_11304);
nand U11410 (N_11410,N_11210,N_11201);
and U11411 (N_11411,N_11217,N_11271);
xor U11412 (N_11412,N_11228,N_11299);
nand U11413 (N_11413,N_11232,N_11359);
or U11414 (N_11414,N_11242,N_11209);
or U11415 (N_11415,N_11303,N_11329);
nor U11416 (N_11416,N_11248,N_11321);
and U11417 (N_11417,N_11281,N_11244);
nor U11418 (N_11418,N_11334,N_11306);
or U11419 (N_11419,N_11218,N_11342);
nand U11420 (N_11420,N_11336,N_11206);
nand U11421 (N_11421,N_11298,N_11259);
nor U11422 (N_11422,N_11279,N_11307);
nand U11423 (N_11423,N_11276,N_11260);
nand U11424 (N_11424,N_11320,N_11316);
nand U11425 (N_11425,N_11353,N_11290);
nor U11426 (N_11426,N_11215,N_11325);
and U11427 (N_11427,N_11254,N_11207);
xor U11428 (N_11428,N_11246,N_11283);
and U11429 (N_11429,N_11214,N_11227);
nor U11430 (N_11430,N_11315,N_11224);
and U11431 (N_11431,N_11311,N_11287);
or U11432 (N_11432,N_11354,N_11249);
xnor U11433 (N_11433,N_11344,N_11264);
and U11434 (N_11434,N_11245,N_11288);
or U11435 (N_11435,N_11297,N_11348);
or U11436 (N_11436,N_11357,N_11284);
xnor U11437 (N_11437,N_11269,N_11233);
nand U11438 (N_11438,N_11258,N_11220);
or U11439 (N_11439,N_11263,N_11302);
nor U11440 (N_11440,N_11316,N_11245);
xnor U11441 (N_11441,N_11268,N_11256);
nor U11442 (N_11442,N_11281,N_11229);
nand U11443 (N_11443,N_11290,N_11208);
nor U11444 (N_11444,N_11254,N_11314);
and U11445 (N_11445,N_11323,N_11335);
and U11446 (N_11446,N_11229,N_11277);
and U11447 (N_11447,N_11292,N_11301);
or U11448 (N_11448,N_11252,N_11357);
nor U11449 (N_11449,N_11359,N_11228);
nand U11450 (N_11450,N_11240,N_11325);
xnor U11451 (N_11451,N_11268,N_11291);
nand U11452 (N_11452,N_11231,N_11238);
nor U11453 (N_11453,N_11348,N_11250);
xnor U11454 (N_11454,N_11313,N_11294);
xor U11455 (N_11455,N_11240,N_11230);
or U11456 (N_11456,N_11221,N_11255);
xnor U11457 (N_11457,N_11292,N_11318);
nor U11458 (N_11458,N_11263,N_11274);
nand U11459 (N_11459,N_11359,N_11239);
and U11460 (N_11460,N_11314,N_11277);
xor U11461 (N_11461,N_11331,N_11359);
or U11462 (N_11462,N_11326,N_11211);
nand U11463 (N_11463,N_11358,N_11278);
xor U11464 (N_11464,N_11327,N_11244);
and U11465 (N_11465,N_11283,N_11277);
nand U11466 (N_11466,N_11280,N_11220);
nor U11467 (N_11467,N_11304,N_11346);
and U11468 (N_11468,N_11264,N_11314);
nand U11469 (N_11469,N_11331,N_11338);
and U11470 (N_11470,N_11234,N_11300);
nand U11471 (N_11471,N_11350,N_11223);
nand U11472 (N_11472,N_11271,N_11326);
nand U11473 (N_11473,N_11285,N_11242);
xor U11474 (N_11474,N_11241,N_11338);
nand U11475 (N_11475,N_11288,N_11347);
nor U11476 (N_11476,N_11343,N_11272);
and U11477 (N_11477,N_11247,N_11317);
and U11478 (N_11478,N_11268,N_11218);
nand U11479 (N_11479,N_11242,N_11248);
nor U11480 (N_11480,N_11258,N_11206);
xor U11481 (N_11481,N_11282,N_11236);
nor U11482 (N_11482,N_11298,N_11284);
nand U11483 (N_11483,N_11330,N_11262);
or U11484 (N_11484,N_11321,N_11207);
xor U11485 (N_11485,N_11295,N_11226);
xor U11486 (N_11486,N_11303,N_11320);
xnor U11487 (N_11487,N_11285,N_11298);
and U11488 (N_11488,N_11268,N_11212);
and U11489 (N_11489,N_11251,N_11207);
or U11490 (N_11490,N_11331,N_11253);
nand U11491 (N_11491,N_11322,N_11265);
nor U11492 (N_11492,N_11290,N_11342);
xor U11493 (N_11493,N_11305,N_11222);
nand U11494 (N_11494,N_11307,N_11348);
or U11495 (N_11495,N_11235,N_11201);
xnor U11496 (N_11496,N_11222,N_11219);
xor U11497 (N_11497,N_11250,N_11252);
xor U11498 (N_11498,N_11330,N_11212);
nand U11499 (N_11499,N_11216,N_11215);
and U11500 (N_11500,N_11250,N_11222);
and U11501 (N_11501,N_11344,N_11255);
nor U11502 (N_11502,N_11214,N_11308);
nand U11503 (N_11503,N_11229,N_11309);
or U11504 (N_11504,N_11252,N_11203);
and U11505 (N_11505,N_11350,N_11226);
nand U11506 (N_11506,N_11245,N_11218);
or U11507 (N_11507,N_11248,N_11299);
and U11508 (N_11508,N_11237,N_11229);
and U11509 (N_11509,N_11353,N_11240);
and U11510 (N_11510,N_11226,N_11233);
and U11511 (N_11511,N_11336,N_11331);
or U11512 (N_11512,N_11299,N_11309);
and U11513 (N_11513,N_11220,N_11356);
nand U11514 (N_11514,N_11295,N_11219);
nor U11515 (N_11515,N_11287,N_11307);
and U11516 (N_11516,N_11279,N_11345);
nor U11517 (N_11517,N_11232,N_11269);
xnor U11518 (N_11518,N_11250,N_11202);
or U11519 (N_11519,N_11326,N_11224);
or U11520 (N_11520,N_11466,N_11385);
and U11521 (N_11521,N_11457,N_11361);
or U11522 (N_11522,N_11428,N_11423);
nor U11523 (N_11523,N_11390,N_11404);
and U11524 (N_11524,N_11452,N_11449);
xor U11525 (N_11525,N_11426,N_11475);
nor U11526 (N_11526,N_11512,N_11447);
nand U11527 (N_11527,N_11402,N_11509);
or U11528 (N_11528,N_11501,N_11460);
xor U11529 (N_11529,N_11411,N_11432);
xnor U11530 (N_11530,N_11379,N_11491);
xnor U11531 (N_11531,N_11362,N_11433);
nand U11532 (N_11532,N_11476,N_11424);
and U11533 (N_11533,N_11389,N_11472);
nor U11534 (N_11534,N_11364,N_11471);
or U11535 (N_11535,N_11497,N_11499);
xor U11536 (N_11536,N_11446,N_11500);
nand U11537 (N_11537,N_11510,N_11455);
nor U11538 (N_11538,N_11377,N_11421);
xnor U11539 (N_11539,N_11419,N_11439);
xnor U11540 (N_11540,N_11518,N_11485);
nor U11541 (N_11541,N_11360,N_11513);
or U11542 (N_11542,N_11397,N_11496);
and U11543 (N_11543,N_11467,N_11488);
or U11544 (N_11544,N_11386,N_11492);
nor U11545 (N_11545,N_11440,N_11408);
nand U11546 (N_11546,N_11392,N_11395);
nor U11547 (N_11547,N_11483,N_11372);
nand U11548 (N_11548,N_11469,N_11366);
and U11549 (N_11549,N_11454,N_11403);
xor U11550 (N_11550,N_11394,N_11489);
xor U11551 (N_11551,N_11401,N_11515);
nand U11552 (N_11552,N_11451,N_11506);
nand U11553 (N_11553,N_11400,N_11505);
nand U11554 (N_11554,N_11374,N_11380);
xnor U11555 (N_11555,N_11458,N_11507);
nand U11556 (N_11556,N_11444,N_11413);
xor U11557 (N_11557,N_11462,N_11429);
nand U11558 (N_11558,N_11498,N_11477);
xnor U11559 (N_11559,N_11479,N_11422);
xor U11560 (N_11560,N_11504,N_11371);
nor U11561 (N_11561,N_11503,N_11405);
xor U11562 (N_11562,N_11415,N_11409);
and U11563 (N_11563,N_11376,N_11470);
nand U11564 (N_11564,N_11516,N_11434);
nand U11565 (N_11565,N_11416,N_11383);
xor U11566 (N_11566,N_11459,N_11375);
nand U11567 (N_11567,N_11370,N_11378);
nor U11568 (N_11568,N_11393,N_11438);
and U11569 (N_11569,N_11490,N_11494);
or U11570 (N_11570,N_11425,N_11481);
and U11571 (N_11571,N_11420,N_11406);
or U11572 (N_11572,N_11382,N_11436);
and U11573 (N_11573,N_11407,N_11441);
and U11574 (N_11574,N_11430,N_11369);
and U11575 (N_11575,N_11399,N_11391);
xnor U11576 (N_11576,N_11511,N_11474);
nor U11577 (N_11577,N_11461,N_11410);
and U11578 (N_11578,N_11484,N_11453);
or U11579 (N_11579,N_11519,N_11456);
and U11580 (N_11580,N_11368,N_11495);
and U11581 (N_11581,N_11514,N_11435);
nor U11582 (N_11582,N_11396,N_11448);
and U11583 (N_11583,N_11508,N_11445);
nand U11584 (N_11584,N_11437,N_11473);
or U11585 (N_11585,N_11398,N_11443);
xor U11586 (N_11586,N_11487,N_11486);
or U11587 (N_11587,N_11412,N_11431);
or U11588 (N_11588,N_11482,N_11381);
and U11589 (N_11589,N_11365,N_11465);
or U11590 (N_11590,N_11478,N_11367);
and U11591 (N_11591,N_11418,N_11517);
and U11592 (N_11592,N_11480,N_11502);
nand U11593 (N_11593,N_11388,N_11384);
xor U11594 (N_11594,N_11363,N_11427);
or U11595 (N_11595,N_11468,N_11450);
or U11596 (N_11596,N_11414,N_11373);
nor U11597 (N_11597,N_11493,N_11442);
xnor U11598 (N_11598,N_11464,N_11387);
and U11599 (N_11599,N_11417,N_11463);
or U11600 (N_11600,N_11392,N_11406);
and U11601 (N_11601,N_11378,N_11422);
or U11602 (N_11602,N_11419,N_11494);
and U11603 (N_11603,N_11411,N_11471);
nand U11604 (N_11604,N_11412,N_11460);
nand U11605 (N_11605,N_11510,N_11486);
xor U11606 (N_11606,N_11427,N_11451);
nand U11607 (N_11607,N_11456,N_11497);
nor U11608 (N_11608,N_11436,N_11378);
xnor U11609 (N_11609,N_11385,N_11433);
nor U11610 (N_11610,N_11502,N_11433);
nor U11611 (N_11611,N_11417,N_11462);
nor U11612 (N_11612,N_11451,N_11364);
or U11613 (N_11613,N_11450,N_11497);
or U11614 (N_11614,N_11457,N_11427);
and U11615 (N_11615,N_11431,N_11376);
nor U11616 (N_11616,N_11458,N_11383);
nor U11617 (N_11617,N_11509,N_11475);
and U11618 (N_11618,N_11420,N_11414);
nand U11619 (N_11619,N_11516,N_11466);
nand U11620 (N_11620,N_11482,N_11455);
nand U11621 (N_11621,N_11472,N_11489);
xor U11622 (N_11622,N_11468,N_11368);
or U11623 (N_11623,N_11395,N_11397);
nand U11624 (N_11624,N_11396,N_11472);
xor U11625 (N_11625,N_11462,N_11453);
nor U11626 (N_11626,N_11416,N_11453);
and U11627 (N_11627,N_11462,N_11439);
xor U11628 (N_11628,N_11428,N_11430);
and U11629 (N_11629,N_11482,N_11433);
or U11630 (N_11630,N_11472,N_11492);
and U11631 (N_11631,N_11394,N_11514);
nor U11632 (N_11632,N_11418,N_11443);
and U11633 (N_11633,N_11454,N_11430);
nand U11634 (N_11634,N_11471,N_11395);
and U11635 (N_11635,N_11385,N_11373);
nand U11636 (N_11636,N_11502,N_11441);
and U11637 (N_11637,N_11506,N_11393);
nor U11638 (N_11638,N_11410,N_11498);
xor U11639 (N_11639,N_11457,N_11366);
nand U11640 (N_11640,N_11459,N_11507);
and U11641 (N_11641,N_11505,N_11402);
nor U11642 (N_11642,N_11495,N_11446);
nand U11643 (N_11643,N_11514,N_11487);
or U11644 (N_11644,N_11476,N_11378);
xor U11645 (N_11645,N_11377,N_11365);
xnor U11646 (N_11646,N_11455,N_11377);
nor U11647 (N_11647,N_11367,N_11369);
xor U11648 (N_11648,N_11423,N_11385);
and U11649 (N_11649,N_11498,N_11392);
nand U11650 (N_11650,N_11469,N_11454);
and U11651 (N_11651,N_11490,N_11519);
nand U11652 (N_11652,N_11362,N_11423);
and U11653 (N_11653,N_11372,N_11418);
and U11654 (N_11654,N_11414,N_11369);
xor U11655 (N_11655,N_11518,N_11382);
or U11656 (N_11656,N_11442,N_11453);
xnor U11657 (N_11657,N_11399,N_11459);
nand U11658 (N_11658,N_11451,N_11495);
xnor U11659 (N_11659,N_11463,N_11406);
and U11660 (N_11660,N_11367,N_11381);
nand U11661 (N_11661,N_11371,N_11492);
and U11662 (N_11662,N_11513,N_11458);
and U11663 (N_11663,N_11443,N_11367);
nand U11664 (N_11664,N_11438,N_11419);
xnor U11665 (N_11665,N_11455,N_11393);
nand U11666 (N_11666,N_11429,N_11400);
and U11667 (N_11667,N_11377,N_11507);
and U11668 (N_11668,N_11409,N_11410);
or U11669 (N_11669,N_11370,N_11401);
nor U11670 (N_11670,N_11364,N_11386);
and U11671 (N_11671,N_11472,N_11423);
and U11672 (N_11672,N_11503,N_11393);
nand U11673 (N_11673,N_11457,N_11505);
xnor U11674 (N_11674,N_11366,N_11490);
and U11675 (N_11675,N_11413,N_11437);
xnor U11676 (N_11676,N_11437,N_11482);
xnor U11677 (N_11677,N_11449,N_11492);
or U11678 (N_11678,N_11467,N_11370);
and U11679 (N_11679,N_11503,N_11497);
nor U11680 (N_11680,N_11604,N_11549);
and U11681 (N_11681,N_11599,N_11629);
xnor U11682 (N_11682,N_11627,N_11534);
and U11683 (N_11683,N_11630,N_11570);
or U11684 (N_11684,N_11577,N_11563);
or U11685 (N_11685,N_11618,N_11679);
and U11686 (N_11686,N_11628,N_11655);
nor U11687 (N_11687,N_11608,N_11631);
or U11688 (N_11688,N_11554,N_11601);
xor U11689 (N_11689,N_11528,N_11579);
nor U11690 (N_11690,N_11561,N_11603);
nand U11691 (N_11691,N_11605,N_11660);
nand U11692 (N_11692,N_11667,N_11658);
and U11693 (N_11693,N_11524,N_11598);
nor U11694 (N_11694,N_11595,N_11575);
nand U11695 (N_11695,N_11673,N_11639);
nor U11696 (N_11696,N_11665,N_11523);
or U11697 (N_11697,N_11632,N_11557);
and U11698 (N_11698,N_11536,N_11542);
nor U11699 (N_11699,N_11527,N_11567);
nor U11700 (N_11700,N_11572,N_11535);
nand U11701 (N_11701,N_11649,N_11586);
xnor U11702 (N_11702,N_11532,N_11522);
nor U11703 (N_11703,N_11612,N_11610);
xor U11704 (N_11704,N_11623,N_11616);
nor U11705 (N_11705,N_11648,N_11576);
nor U11706 (N_11706,N_11583,N_11677);
nor U11707 (N_11707,N_11529,N_11611);
or U11708 (N_11708,N_11600,N_11590);
and U11709 (N_11709,N_11556,N_11565);
xnor U11710 (N_11710,N_11525,N_11545);
xnor U11711 (N_11711,N_11675,N_11581);
and U11712 (N_11712,N_11584,N_11656);
xnor U11713 (N_11713,N_11569,N_11621);
nand U11714 (N_11714,N_11607,N_11650);
xor U11715 (N_11715,N_11596,N_11635);
xnor U11716 (N_11716,N_11626,N_11589);
or U11717 (N_11717,N_11633,N_11538);
xor U11718 (N_11718,N_11606,N_11676);
nor U11719 (N_11719,N_11559,N_11647);
nor U11720 (N_11720,N_11541,N_11653);
nand U11721 (N_11721,N_11664,N_11638);
or U11722 (N_11722,N_11645,N_11663);
or U11723 (N_11723,N_11602,N_11652);
nand U11724 (N_11724,N_11642,N_11620);
nand U11725 (N_11725,N_11625,N_11668);
nor U11726 (N_11726,N_11594,N_11585);
xnor U11727 (N_11727,N_11547,N_11659);
xnor U11728 (N_11728,N_11613,N_11550);
xor U11729 (N_11729,N_11588,N_11622);
nor U11730 (N_11730,N_11531,N_11637);
nand U11731 (N_11731,N_11553,N_11520);
or U11732 (N_11732,N_11562,N_11526);
and U11733 (N_11733,N_11615,N_11609);
nand U11734 (N_11734,N_11674,N_11641);
or U11735 (N_11735,N_11551,N_11580);
nor U11736 (N_11736,N_11636,N_11672);
or U11737 (N_11737,N_11558,N_11614);
or U11738 (N_11738,N_11593,N_11568);
xnor U11739 (N_11739,N_11670,N_11662);
nor U11740 (N_11740,N_11560,N_11643);
or U11741 (N_11741,N_11654,N_11571);
xnor U11742 (N_11742,N_11671,N_11548);
and U11743 (N_11743,N_11661,N_11521);
xor U11744 (N_11744,N_11537,N_11678);
xnor U11745 (N_11745,N_11666,N_11552);
nor U11746 (N_11746,N_11592,N_11566);
or U11747 (N_11747,N_11640,N_11574);
and U11748 (N_11748,N_11644,N_11544);
or U11749 (N_11749,N_11657,N_11591);
and U11750 (N_11750,N_11555,N_11530);
xnor U11751 (N_11751,N_11646,N_11617);
and U11752 (N_11752,N_11533,N_11578);
and U11753 (N_11753,N_11546,N_11543);
and U11754 (N_11754,N_11669,N_11564);
nor U11755 (N_11755,N_11624,N_11573);
nand U11756 (N_11756,N_11619,N_11587);
or U11757 (N_11757,N_11597,N_11539);
or U11758 (N_11758,N_11582,N_11540);
or U11759 (N_11759,N_11634,N_11651);
or U11760 (N_11760,N_11650,N_11572);
xor U11761 (N_11761,N_11536,N_11651);
or U11762 (N_11762,N_11534,N_11676);
nand U11763 (N_11763,N_11610,N_11636);
and U11764 (N_11764,N_11535,N_11591);
nor U11765 (N_11765,N_11555,N_11667);
xnor U11766 (N_11766,N_11642,N_11543);
xnor U11767 (N_11767,N_11610,N_11568);
nor U11768 (N_11768,N_11601,N_11634);
nor U11769 (N_11769,N_11643,N_11551);
xor U11770 (N_11770,N_11657,N_11616);
nor U11771 (N_11771,N_11574,N_11538);
xor U11772 (N_11772,N_11521,N_11605);
nand U11773 (N_11773,N_11564,N_11660);
and U11774 (N_11774,N_11577,N_11572);
nor U11775 (N_11775,N_11666,N_11672);
and U11776 (N_11776,N_11543,N_11527);
nand U11777 (N_11777,N_11581,N_11613);
or U11778 (N_11778,N_11575,N_11669);
and U11779 (N_11779,N_11654,N_11531);
and U11780 (N_11780,N_11585,N_11677);
nand U11781 (N_11781,N_11573,N_11625);
xor U11782 (N_11782,N_11630,N_11524);
and U11783 (N_11783,N_11538,N_11645);
nand U11784 (N_11784,N_11554,N_11610);
nand U11785 (N_11785,N_11669,N_11528);
nor U11786 (N_11786,N_11578,N_11539);
xor U11787 (N_11787,N_11610,N_11536);
or U11788 (N_11788,N_11523,N_11594);
nor U11789 (N_11789,N_11607,N_11547);
and U11790 (N_11790,N_11578,N_11532);
nand U11791 (N_11791,N_11599,N_11627);
and U11792 (N_11792,N_11635,N_11542);
xnor U11793 (N_11793,N_11598,N_11637);
and U11794 (N_11794,N_11593,N_11583);
nand U11795 (N_11795,N_11529,N_11565);
and U11796 (N_11796,N_11547,N_11671);
or U11797 (N_11797,N_11614,N_11541);
nand U11798 (N_11798,N_11547,N_11637);
xor U11799 (N_11799,N_11642,N_11592);
xor U11800 (N_11800,N_11551,N_11526);
and U11801 (N_11801,N_11593,N_11563);
nand U11802 (N_11802,N_11644,N_11539);
and U11803 (N_11803,N_11651,N_11570);
nand U11804 (N_11804,N_11622,N_11585);
nand U11805 (N_11805,N_11541,N_11601);
nand U11806 (N_11806,N_11571,N_11660);
nand U11807 (N_11807,N_11524,N_11550);
nand U11808 (N_11808,N_11611,N_11629);
and U11809 (N_11809,N_11553,N_11541);
nor U11810 (N_11810,N_11598,N_11628);
and U11811 (N_11811,N_11589,N_11522);
xor U11812 (N_11812,N_11555,N_11622);
nor U11813 (N_11813,N_11555,N_11670);
or U11814 (N_11814,N_11598,N_11666);
or U11815 (N_11815,N_11636,N_11577);
xor U11816 (N_11816,N_11535,N_11585);
xor U11817 (N_11817,N_11633,N_11662);
or U11818 (N_11818,N_11578,N_11626);
and U11819 (N_11819,N_11524,N_11577);
xnor U11820 (N_11820,N_11607,N_11584);
nor U11821 (N_11821,N_11532,N_11679);
nor U11822 (N_11822,N_11658,N_11572);
nand U11823 (N_11823,N_11629,N_11626);
nand U11824 (N_11824,N_11628,N_11610);
or U11825 (N_11825,N_11606,N_11605);
or U11826 (N_11826,N_11557,N_11662);
or U11827 (N_11827,N_11620,N_11652);
xnor U11828 (N_11828,N_11587,N_11586);
nor U11829 (N_11829,N_11609,N_11550);
and U11830 (N_11830,N_11661,N_11561);
or U11831 (N_11831,N_11528,N_11608);
nor U11832 (N_11832,N_11577,N_11580);
or U11833 (N_11833,N_11600,N_11555);
xor U11834 (N_11834,N_11584,N_11562);
nand U11835 (N_11835,N_11565,N_11658);
xnor U11836 (N_11836,N_11592,N_11522);
xor U11837 (N_11837,N_11677,N_11565);
nor U11838 (N_11838,N_11606,N_11607);
xnor U11839 (N_11839,N_11621,N_11676);
nand U11840 (N_11840,N_11780,N_11720);
nand U11841 (N_11841,N_11763,N_11778);
nand U11842 (N_11842,N_11775,N_11836);
nand U11843 (N_11843,N_11769,N_11779);
nand U11844 (N_11844,N_11838,N_11750);
xor U11845 (N_11845,N_11751,N_11821);
nand U11846 (N_11846,N_11802,N_11795);
nor U11847 (N_11847,N_11723,N_11712);
nand U11848 (N_11848,N_11801,N_11799);
and U11849 (N_11849,N_11793,N_11792);
or U11850 (N_11850,N_11722,N_11759);
and U11851 (N_11851,N_11697,N_11745);
xor U11852 (N_11852,N_11732,N_11761);
nor U11853 (N_11853,N_11803,N_11728);
nor U11854 (N_11854,N_11797,N_11680);
and U11855 (N_11855,N_11718,N_11812);
xor U11856 (N_11856,N_11800,N_11729);
and U11857 (N_11857,N_11706,N_11776);
nand U11858 (N_11858,N_11826,N_11777);
and U11859 (N_11859,N_11824,N_11839);
xor U11860 (N_11860,N_11796,N_11837);
xor U11861 (N_11861,N_11828,N_11707);
nor U11862 (N_11862,N_11700,N_11773);
or U11863 (N_11863,N_11699,N_11743);
or U11864 (N_11864,N_11790,N_11816);
nor U11865 (N_11865,N_11834,N_11721);
nor U11866 (N_11866,N_11810,N_11739);
and U11867 (N_11867,N_11771,N_11789);
nor U11868 (N_11868,N_11682,N_11691);
nand U11869 (N_11869,N_11783,N_11701);
nor U11870 (N_11870,N_11693,N_11829);
or U11871 (N_11871,N_11788,N_11749);
xnor U11872 (N_11872,N_11683,N_11730);
nor U11873 (N_11873,N_11756,N_11704);
and U11874 (N_11874,N_11798,N_11738);
or U11875 (N_11875,N_11708,N_11833);
xor U11876 (N_11876,N_11760,N_11762);
and U11877 (N_11877,N_11719,N_11695);
nand U11878 (N_11878,N_11767,N_11753);
and U11879 (N_11879,N_11791,N_11755);
nand U11880 (N_11880,N_11811,N_11711);
nor U11881 (N_11881,N_11702,N_11804);
xnor U11882 (N_11882,N_11757,N_11742);
nor U11883 (N_11883,N_11827,N_11808);
and U11884 (N_11884,N_11787,N_11744);
and U11885 (N_11885,N_11690,N_11716);
xor U11886 (N_11886,N_11698,N_11692);
xnor U11887 (N_11887,N_11713,N_11825);
or U11888 (N_11888,N_11731,N_11734);
nand U11889 (N_11889,N_11786,N_11817);
or U11890 (N_11890,N_11782,N_11815);
or U11891 (N_11891,N_11725,N_11703);
nor U11892 (N_11892,N_11764,N_11831);
nand U11893 (N_11893,N_11805,N_11814);
and U11894 (N_11894,N_11727,N_11784);
xnor U11895 (N_11895,N_11754,N_11726);
nor U11896 (N_11896,N_11835,N_11714);
nand U11897 (N_11897,N_11806,N_11818);
nor U11898 (N_11898,N_11781,N_11740);
nand U11899 (N_11899,N_11724,N_11768);
nor U11900 (N_11900,N_11735,N_11770);
and U11901 (N_11901,N_11822,N_11686);
or U11902 (N_11902,N_11733,N_11813);
nand U11903 (N_11903,N_11710,N_11832);
and U11904 (N_11904,N_11685,N_11709);
and U11905 (N_11905,N_11809,N_11688);
or U11906 (N_11906,N_11807,N_11746);
nor U11907 (N_11907,N_11684,N_11705);
or U11908 (N_11908,N_11737,N_11747);
or U11909 (N_11909,N_11687,N_11736);
xnor U11910 (N_11910,N_11819,N_11752);
and U11911 (N_11911,N_11820,N_11830);
xnor U11912 (N_11912,N_11766,N_11758);
xor U11913 (N_11913,N_11748,N_11794);
xnor U11914 (N_11914,N_11717,N_11823);
nor U11915 (N_11915,N_11772,N_11765);
and U11916 (N_11916,N_11715,N_11694);
xor U11917 (N_11917,N_11689,N_11681);
nor U11918 (N_11918,N_11774,N_11785);
and U11919 (N_11919,N_11741,N_11696);
and U11920 (N_11920,N_11822,N_11695);
and U11921 (N_11921,N_11779,N_11799);
nor U11922 (N_11922,N_11777,N_11839);
or U11923 (N_11923,N_11751,N_11829);
xnor U11924 (N_11924,N_11813,N_11740);
and U11925 (N_11925,N_11712,N_11705);
nor U11926 (N_11926,N_11779,N_11782);
or U11927 (N_11927,N_11729,N_11839);
nor U11928 (N_11928,N_11823,N_11736);
and U11929 (N_11929,N_11739,N_11809);
nor U11930 (N_11930,N_11688,N_11831);
or U11931 (N_11931,N_11744,N_11730);
nand U11932 (N_11932,N_11743,N_11701);
nor U11933 (N_11933,N_11819,N_11777);
xnor U11934 (N_11934,N_11782,N_11760);
and U11935 (N_11935,N_11681,N_11806);
nand U11936 (N_11936,N_11700,N_11817);
xor U11937 (N_11937,N_11745,N_11797);
nor U11938 (N_11938,N_11781,N_11832);
and U11939 (N_11939,N_11799,N_11762);
and U11940 (N_11940,N_11752,N_11770);
nor U11941 (N_11941,N_11707,N_11832);
nor U11942 (N_11942,N_11686,N_11827);
or U11943 (N_11943,N_11754,N_11748);
nand U11944 (N_11944,N_11723,N_11811);
and U11945 (N_11945,N_11812,N_11738);
xnor U11946 (N_11946,N_11696,N_11802);
nor U11947 (N_11947,N_11832,N_11714);
or U11948 (N_11948,N_11753,N_11762);
or U11949 (N_11949,N_11785,N_11756);
and U11950 (N_11950,N_11748,N_11726);
nand U11951 (N_11951,N_11808,N_11700);
nor U11952 (N_11952,N_11834,N_11727);
or U11953 (N_11953,N_11746,N_11806);
nor U11954 (N_11954,N_11759,N_11813);
or U11955 (N_11955,N_11835,N_11804);
or U11956 (N_11956,N_11728,N_11738);
and U11957 (N_11957,N_11812,N_11774);
xor U11958 (N_11958,N_11762,N_11800);
or U11959 (N_11959,N_11808,N_11750);
and U11960 (N_11960,N_11706,N_11757);
xor U11961 (N_11961,N_11747,N_11716);
xor U11962 (N_11962,N_11764,N_11731);
or U11963 (N_11963,N_11751,N_11761);
nand U11964 (N_11964,N_11767,N_11771);
and U11965 (N_11965,N_11762,N_11686);
or U11966 (N_11966,N_11803,N_11726);
xnor U11967 (N_11967,N_11789,N_11694);
or U11968 (N_11968,N_11757,N_11744);
nor U11969 (N_11969,N_11788,N_11750);
nor U11970 (N_11970,N_11807,N_11813);
nand U11971 (N_11971,N_11805,N_11687);
or U11972 (N_11972,N_11771,N_11741);
nor U11973 (N_11973,N_11690,N_11719);
nand U11974 (N_11974,N_11818,N_11748);
xnor U11975 (N_11975,N_11793,N_11744);
or U11976 (N_11976,N_11767,N_11817);
or U11977 (N_11977,N_11686,N_11825);
nand U11978 (N_11978,N_11816,N_11835);
or U11979 (N_11979,N_11737,N_11799);
nand U11980 (N_11980,N_11837,N_11784);
xnor U11981 (N_11981,N_11749,N_11823);
nand U11982 (N_11982,N_11758,N_11768);
xnor U11983 (N_11983,N_11823,N_11684);
and U11984 (N_11984,N_11788,N_11835);
and U11985 (N_11985,N_11780,N_11795);
xnor U11986 (N_11986,N_11758,N_11743);
nor U11987 (N_11987,N_11690,N_11692);
nor U11988 (N_11988,N_11755,N_11782);
xnor U11989 (N_11989,N_11831,N_11802);
nand U11990 (N_11990,N_11782,N_11682);
nor U11991 (N_11991,N_11789,N_11803);
or U11992 (N_11992,N_11755,N_11764);
nor U11993 (N_11993,N_11833,N_11812);
or U11994 (N_11994,N_11768,N_11808);
nor U11995 (N_11995,N_11686,N_11706);
nand U11996 (N_11996,N_11760,N_11700);
and U11997 (N_11997,N_11787,N_11715);
nor U11998 (N_11998,N_11717,N_11737);
and U11999 (N_11999,N_11782,N_11703);
nand U12000 (N_12000,N_11896,N_11874);
xnor U12001 (N_12001,N_11988,N_11978);
nand U12002 (N_12002,N_11956,N_11856);
nand U12003 (N_12003,N_11882,N_11916);
nor U12004 (N_12004,N_11851,N_11987);
nor U12005 (N_12005,N_11902,N_11949);
nand U12006 (N_12006,N_11940,N_11908);
and U12007 (N_12007,N_11843,N_11952);
xor U12008 (N_12008,N_11983,N_11903);
nand U12009 (N_12009,N_11871,N_11936);
and U12010 (N_12010,N_11923,N_11880);
xor U12011 (N_12011,N_11866,N_11844);
xor U12012 (N_12012,N_11979,N_11905);
xor U12013 (N_12013,N_11850,N_11971);
xnor U12014 (N_12014,N_11974,N_11964);
xnor U12015 (N_12015,N_11991,N_11841);
xor U12016 (N_12016,N_11989,N_11976);
nand U12017 (N_12017,N_11865,N_11864);
nor U12018 (N_12018,N_11924,N_11914);
nor U12019 (N_12019,N_11845,N_11953);
nand U12020 (N_12020,N_11857,N_11852);
nand U12021 (N_12021,N_11922,N_11977);
nand U12022 (N_12022,N_11901,N_11946);
nand U12023 (N_12023,N_11962,N_11873);
xor U12024 (N_12024,N_11883,N_11915);
nor U12025 (N_12025,N_11907,N_11913);
and U12026 (N_12026,N_11959,N_11981);
nor U12027 (N_12027,N_11861,N_11869);
xor U12028 (N_12028,N_11945,N_11853);
or U12029 (N_12029,N_11943,N_11994);
xor U12030 (N_12030,N_11858,N_11957);
and U12031 (N_12031,N_11878,N_11909);
or U12032 (N_12032,N_11848,N_11982);
and U12033 (N_12033,N_11842,N_11854);
or U12034 (N_12034,N_11879,N_11860);
nand U12035 (N_12035,N_11973,N_11904);
xor U12036 (N_12036,N_11855,N_11870);
nand U12037 (N_12037,N_11970,N_11931);
xnor U12038 (N_12038,N_11911,N_11872);
nor U12039 (N_12039,N_11893,N_11875);
nand U12040 (N_12040,N_11847,N_11995);
xor U12041 (N_12041,N_11906,N_11929);
nand U12042 (N_12042,N_11965,N_11985);
and U12043 (N_12043,N_11926,N_11997);
or U12044 (N_12044,N_11888,N_11963);
nor U12045 (N_12045,N_11881,N_11930);
nand U12046 (N_12046,N_11899,N_11900);
or U12047 (N_12047,N_11958,N_11910);
nor U12048 (N_12048,N_11876,N_11894);
or U12049 (N_12049,N_11898,N_11935);
nor U12050 (N_12050,N_11947,N_11927);
or U12051 (N_12051,N_11889,N_11897);
nand U12052 (N_12052,N_11950,N_11846);
and U12053 (N_12053,N_11942,N_11890);
nand U12054 (N_12054,N_11892,N_11984);
nand U12055 (N_12055,N_11919,N_11912);
nand U12056 (N_12056,N_11867,N_11941);
xnor U12057 (N_12057,N_11990,N_11938);
nand U12058 (N_12058,N_11980,N_11933);
xnor U12059 (N_12059,N_11992,N_11934);
or U12060 (N_12060,N_11921,N_11944);
nor U12061 (N_12061,N_11993,N_11895);
nand U12062 (N_12062,N_11863,N_11996);
and U12063 (N_12063,N_11939,N_11928);
xnor U12064 (N_12064,N_11961,N_11891);
xor U12065 (N_12065,N_11999,N_11877);
or U12066 (N_12066,N_11937,N_11955);
and U12067 (N_12067,N_11886,N_11849);
nor U12068 (N_12068,N_11840,N_11868);
or U12069 (N_12069,N_11986,N_11917);
or U12070 (N_12070,N_11951,N_11966);
xnor U12071 (N_12071,N_11960,N_11862);
or U12072 (N_12072,N_11975,N_11887);
nor U12073 (N_12073,N_11967,N_11954);
nor U12074 (N_12074,N_11918,N_11925);
nand U12075 (N_12075,N_11972,N_11885);
and U12076 (N_12076,N_11968,N_11969);
nand U12077 (N_12077,N_11920,N_11948);
nor U12078 (N_12078,N_11884,N_11932);
xnor U12079 (N_12079,N_11859,N_11998);
xnor U12080 (N_12080,N_11857,N_11970);
and U12081 (N_12081,N_11891,N_11926);
xor U12082 (N_12082,N_11950,N_11947);
xnor U12083 (N_12083,N_11902,N_11994);
and U12084 (N_12084,N_11934,N_11989);
nor U12085 (N_12085,N_11873,N_11997);
and U12086 (N_12086,N_11897,N_11941);
or U12087 (N_12087,N_11977,N_11868);
nand U12088 (N_12088,N_11928,N_11996);
and U12089 (N_12089,N_11920,N_11880);
nor U12090 (N_12090,N_11842,N_11933);
or U12091 (N_12091,N_11849,N_11961);
nand U12092 (N_12092,N_11950,N_11916);
nand U12093 (N_12093,N_11992,N_11925);
and U12094 (N_12094,N_11854,N_11907);
or U12095 (N_12095,N_11863,N_11841);
xnor U12096 (N_12096,N_11949,N_11857);
nor U12097 (N_12097,N_11867,N_11963);
xor U12098 (N_12098,N_11864,N_11905);
nand U12099 (N_12099,N_11929,N_11870);
or U12100 (N_12100,N_11877,N_11942);
or U12101 (N_12101,N_11851,N_11913);
nand U12102 (N_12102,N_11970,N_11868);
or U12103 (N_12103,N_11948,N_11904);
nor U12104 (N_12104,N_11937,N_11920);
and U12105 (N_12105,N_11877,N_11973);
or U12106 (N_12106,N_11881,N_11911);
nand U12107 (N_12107,N_11977,N_11971);
or U12108 (N_12108,N_11934,N_11887);
and U12109 (N_12109,N_11900,N_11858);
xnor U12110 (N_12110,N_11881,N_11986);
or U12111 (N_12111,N_11924,N_11890);
nor U12112 (N_12112,N_11925,N_11857);
and U12113 (N_12113,N_11901,N_11915);
and U12114 (N_12114,N_11979,N_11916);
and U12115 (N_12115,N_11891,N_11841);
and U12116 (N_12116,N_11866,N_11842);
xnor U12117 (N_12117,N_11906,N_11880);
and U12118 (N_12118,N_11864,N_11975);
xor U12119 (N_12119,N_11940,N_11923);
or U12120 (N_12120,N_11919,N_11935);
or U12121 (N_12121,N_11978,N_11900);
or U12122 (N_12122,N_11842,N_11948);
or U12123 (N_12123,N_11894,N_11840);
nor U12124 (N_12124,N_11911,N_11971);
and U12125 (N_12125,N_11943,N_11860);
nor U12126 (N_12126,N_11907,N_11961);
nand U12127 (N_12127,N_11977,N_11897);
nand U12128 (N_12128,N_11872,N_11855);
or U12129 (N_12129,N_11858,N_11972);
xor U12130 (N_12130,N_11924,N_11857);
nand U12131 (N_12131,N_11959,N_11896);
nor U12132 (N_12132,N_11944,N_11871);
and U12133 (N_12133,N_11907,N_11969);
nand U12134 (N_12134,N_11851,N_11963);
xnor U12135 (N_12135,N_11911,N_11932);
and U12136 (N_12136,N_11949,N_11858);
xor U12137 (N_12137,N_11942,N_11924);
nor U12138 (N_12138,N_11860,N_11865);
nand U12139 (N_12139,N_11945,N_11894);
nand U12140 (N_12140,N_11904,N_11932);
nor U12141 (N_12141,N_11862,N_11924);
and U12142 (N_12142,N_11917,N_11860);
nand U12143 (N_12143,N_11995,N_11846);
nand U12144 (N_12144,N_11992,N_11946);
nor U12145 (N_12145,N_11913,N_11994);
or U12146 (N_12146,N_11952,N_11997);
nor U12147 (N_12147,N_11977,N_11953);
nor U12148 (N_12148,N_11910,N_11900);
or U12149 (N_12149,N_11888,N_11851);
nor U12150 (N_12150,N_11978,N_11977);
nor U12151 (N_12151,N_11917,N_11960);
nor U12152 (N_12152,N_11896,N_11998);
or U12153 (N_12153,N_11926,N_11851);
or U12154 (N_12154,N_11874,N_11972);
nand U12155 (N_12155,N_11955,N_11978);
nor U12156 (N_12156,N_11930,N_11890);
nand U12157 (N_12157,N_11915,N_11878);
xnor U12158 (N_12158,N_11973,N_11873);
nor U12159 (N_12159,N_11903,N_11874);
nand U12160 (N_12160,N_12092,N_12065);
and U12161 (N_12161,N_12032,N_12104);
nor U12162 (N_12162,N_12108,N_12107);
nand U12163 (N_12163,N_12009,N_12044);
nor U12164 (N_12164,N_12057,N_12022);
nand U12165 (N_12165,N_12097,N_12091);
and U12166 (N_12166,N_12127,N_12043);
and U12167 (N_12167,N_12099,N_12025);
nor U12168 (N_12168,N_12039,N_12085);
or U12169 (N_12169,N_12008,N_12111);
nor U12170 (N_12170,N_12078,N_12142);
xnor U12171 (N_12171,N_12070,N_12136);
and U12172 (N_12172,N_12114,N_12056);
nand U12173 (N_12173,N_12115,N_12051);
xnor U12174 (N_12174,N_12081,N_12106);
nor U12175 (N_12175,N_12156,N_12030);
nor U12176 (N_12176,N_12011,N_12047);
xor U12177 (N_12177,N_12080,N_12132);
or U12178 (N_12178,N_12034,N_12068);
nand U12179 (N_12179,N_12090,N_12063);
nand U12180 (N_12180,N_12058,N_12005);
nor U12181 (N_12181,N_12024,N_12137);
nor U12182 (N_12182,N_12118,N_12098);
nand U12183 (N_12183,N_12073,N_12117);
nor U12184 (N_12184,N_12120,N_12052);
or U12185 (N_12185,N_12053,N_12149);
or U12186 (N_12186,N_12028,N_12001);
nor U12187 (N_12187,N_12101,N_12105);
or U12188 (N_12188,N_12155,N_12029);
nand U12189 (N_12189,N_12019,N_12014);
xnor U12190 (N_12190,N_12006,N_12079);
nor U12191 (N_12191,N_12093,N_12012);
xor U12192 (N_12192,N_12003,N_12017);
or U12193 (N_12193,N_12067,N_12134);
and U12194 (N_12194,N_12059,N_12074);
nor U12195 (N_12195,N_12066,N_12061);
xor U12196 (N_12196,N_12158,N_12151);
nand U12197 (N_12197,N_12145,N_12131);
or U12198 (N_12198,N_12035,N_12040);
or U12199 (N_12199,N_12086,N_12144);
nor U12200 (N_12200,N_12077,N_12013);
or U12201 (N_12201,N_12037,N_12143);
or U12202 (N_12202,N_12119,N_12159);
nand U12203 (N_12203,N_12042,N_12010);
nor U12204 (N_12204,N_12102,N_12089);
nor U12205 (N_12205,N_12153,N_12087);
nor U12206 (N_12206,N_12060,N_12064);
and U12207 (N_12207,N_12146,N_12083);
xor U12208 (N_12208,N_12157,N_12126);
and U12209 (N_12209,N_12082,N_12130);
and U12210 (N_12210,N_12129,N_12096);
or U12211 (N_12211,N_12069,N_12124);
and U12212 (N_12212,N_12041,N_12020);
and U12213 (N_12213,N_12123,N_12076);
nand U12214 (N_12214,N_12007,N_12018);
or U12215 (N_12215,N_12152,N_12055);
xor U12216 (N_12216,N_12027,N_12148);
or U12217 (N_12217,N_12103,N_12084);
or U12218 (N_12218,N_12045,N_12122);
and U12219 (N_12219,N_12113,N_12135);
nand U12220 (N_12220,N_12125,N_12049);
or U12221 (N_12221,N_12112,N_12094);
and U12222 (N_12222,N_12140,N_12033);
xor U12223 (N_12223,N_12004,N_12000);
xnor U12224 (N_12224,N_12095,N_12100);
xor U12225 (N_12225,N_12038,N_12036);
nor U12226 (N_12226,N_12075,N_12138);
nand U12227 (N_12227,N_12031,N_12147);
and U12228 (N_12228,N_12109,N_12015);
nor U12229 (N_12229,N_12062,N_12088);
xor U12230 (N_12230,N_12154,N_12121);
and U12231 (N_12231,N_12139,N_12048);
xor U12232 (N_12232,N_12071,N_12116);
nand U12233 (N_12233,N_12023,N_12016);
nor U12234 (N_12234,N_12021,N_12110);
xnor U12235 (N_12235,N_12141,N_12054);
or U12236 (N_12236,N_12046,N_12133);
nor U12237 (N_12237,N_12002,N_12050);
xor U12238 (N_12238,N_12026,N_12128);
and U12239 (N_12239,N_12072,N_12150);
or U12240 (N_12240,N_12106,N_12097);
nand U12241 (N_12241,N_12120,N_12006);
xor U12242 (N_12242,N_12109,N_12136);
nor U12243 (N_12243,N_12069,N_12004);
and U12244 (N_12244,N_12103,N_12015);
xor U12245 (N_12245,N_12024,N_12081);
and U12246 (N_12246,N_12137,N_12047);
and U12247 (N_12247,N_12149,N_12004);
nand U12248 (N_12248,N_12106,N_12104);
xor U12249 (N_12249,N_12117,N_12130);
xnor U12250 (N_12250,N_12013,N_12088);
and U12251 (N_12251,N_12107,N_12104);
and U12252 (N_12252,N_12030,N_12087);
and U12253 (N_12253,N_12119,N_12108);
or U12254 (N_12254,N_12129,N_12036);
and U12255 (N_12255,N_12104,N_12140);
and U12256 (N_12256,N_12144,N_12083);
xor U12257 (N_12257,N_12095,N_12152);
and U12258 (N_12258,N_12136,N_12087);
and U12259 (N_12259,N_12003,N_12044);
and U12260 (N_12260,N_12153,N_12002);
nand U12261 (N_12261,N_12006,N_12022);
nor U12262 (N_12262,N_12086,N_12083);
nand U12263 (N_12263,N_12052,N_12081);
nand U12264 (N_12264,N_12134,N_12027);
and U12265 (N_12265,N_12109,N_12110);
nand U12266 (N_12266,N_12029,N_12047);
or U12267 (N_12267,N_12066,N_12059);
and U12268 (N_12268,N_12042,N_12119);
xnor U12269 (N_12269,N_12036,N_12059);
nand U12270 (N_12270,N_12133,N_12060);
nand U12271 (N_12271,N_12159,N_12074);
nor U12272 (N_12272,N_12024,N_12123);
or U12273 (N_12273,N_12107,N_12036);
nand U12274 (N_12274,N_12102,N_12077);
nor U12275 (N_12275,N_12066,N_12006);
and U12276 (N_12276,N_12023,N_12114);
xnor U12277 (N_12277,N_12117,N_12129);
and U12278 (N_12278,N_12027,N_12130);
and U12279 (N_12279,N_12107,N_12052);
and U12280 (N_12280,N_12122,N_12121);
and U12281 (N_12281,N_12075,N_12083);
nor U12282 (N_12282,N_12106,N_12016);
nand U12283 (N_12283,N_12032,N_12100);
and U12284 (N_12284,N_12064,N_12019);
nand U12285 (N_12285,N_12007,N_12023);
nor U12286 (N_12286,N_12133,N_12048);
nor U12287 (N_12287,N_12104,N_12137);
xnor U12288 (N_12288,N_12043,N_12114);
xor U12289 (N_12289,N_12155,N_12118);
xnor U12290 (N_12290,N_12120,N_12125);
and U12291 (N_12291,N_12086,N_12015);
nor U12292 (N_12292,N_12106,N_12021);
nor U12293 (N_12293,N_12126,N_12141);
and U12294 (N_12294,N_12019,N_12108);
nor U12295 (N_12295,N_12150,N_12101);
nor U12296 (N_12296,N_12014,N_12023);
and U12297 (N_12297,N_12150,N_12120);
nor U12298 (N_12298,N_12070,N_12075);
nor U12299 (N_12299,N_12140,N_12109);
nor U12300 (N_12300,N_12102,N_12141);
nor U12301 (N_12301,N_12128,N_12087);
nor U12302 (N_12302,N_12153,N_12151);
and U12303 (N_12303,N_12150,N_12123);
nand U12304 (N_12304,N_12036,N_12083);
nand U12305 (N_12305,N_12128,N_12136);
or U12306 (N_12306,N_12026,N_12051);
nor U12307 (N_12307,N_12015,N_12154);
and U12308 (N_12308,N_12035,N_12055);
xnor U12309 (N_12309,N_12040,N_12041);
nor U12310 (N_12310,N_12113,N_12089);
and U12311 (N_12311,N_12013,N_12128);
xor U12312 (N_12312,N_12062,N_12102);
nand U12313 (N_12313,N_12116,N_12079);
nor U12314 (N_12314,N_12118,N_12049);
and U12315 (N_12315,N_12103,N_12075);
and U12316 (N_12316,N_12092,N_12155);
and U12317 (N_12317,N_12091,N_12019);
or U12318 (N_12318,N_12055,N_12092);
xor U12319 (N_12319,N_12043,N_12103);
xor U12320 (N_12320,N_12262,N_12210);
nand U12321 (N_12321,N_12286,N_12281);
nor U12322 (N_12322,N_12182,N_12288);
and U12323 (N_12323,N_12198,N_12278);
or U12324 (N_12324,N_12282,N_12235);
or U12325 (N_12325,N_12221,N_12174);
or U12326 (N_12326,N_12189,N_12269);
and U12327 (N_12327,N_12166,N_12305);
nand U12328 (N_12328,N_12244,N_12218);
and U12329 (N_12329,N_12181,N_12212);
xnor U12330 (N_12330,N_12161,N_12193);
or U12331 (N_12331,N_12237,N_12230);
and U12332 (N_12332,N_12162,N_12266);
or U12333 (N_12333,N_12248,N_12216);
or U12334 (N_12334,N_12294,N_12307);
nand U12335 (N_12335,N_12298,N_12309);
or U12336 (N_12336,N_12254,N_12194);
nand U12337 (N_12337,N_12208,N_12243);
nand U12338 (N_12338,N_12300,N_12213);
nand U12339 (N_12339,N_12242,N_12249);
or U12340 (N_12340,N_12241,N_12268);
nor U12341 (N_12341,N_12270,N_12238);
or U12342 (N_12342,N_12306,N_12265);
nand U12343 (N_12343,N_12257,N_12317);
or U12344 (N_12344,N_12163,N_12301);
nor U12345 (N_12345,N_12318,N_12165);
xnor U12346 (N_12346,N_12222,N_12172);
xor U12347 (N_12347,N_12173,N_12178);
nor U12348 (N_12348,N_12233,N_12180);
nor U12349 (N_12349,N_12303,N_12264);
or U12350 (N_12350,N_12292,N_12226);
and U12351 (N_12351,N_12188,N_12204);
xor U12352 (N_12352,N_12229,N_12186);
nand U12353 (N_12353,N_12315,N_12227);
nor U12354 (N_12354,N_12289,N_12250);
xnor U12355 (N_12355,N_12234,N_12160);
xor U12356 (N_12356,N_12283,N_12175);
or U12357 (N_12357,N_12184,N_12263);
or U12358 (N_12358,N_12200,N_12192);
and U12359 (N_12359,N_12253,N_12201);
or U12360 (N_12360,N_12225,N_12187);
or U12361 (N_12361,N_12319,N_12231);
nor U12362 (N_12362,N_12232,N_12314);
xor U12363 (N_12363,N_12275,N_12211);
or U12364 (N_12364,N_12195,N_12267);
nor U12365 (N_12365,N_12177,N_12293);
nor U12366 (N_12366,N_12284,N_12205);
nand U12367 (N_12367,N_12256,N_12224);
and U12368 (N_12368,N_12167,N_12302);
nand U12369 (N_12369,N_12304,N_12311);
or U12370 (N_12370,N_12272,N_12215);
nand U12371 (N_12371,N_12239,N_12228);
nand U12372 (N_12372,N_12206,N_12169);
nor U12373 (N_12373,N_12291,N_12290);
nand U12374 (N_12374,N_12310,N_12209);
and U12375 (N_12375,N_12190,N_12176);
and U12376 (N_12376,N_12297,N_12202);
or U12377 (N_12377,N_12296,N_12299);
or U12378 (N_12378,N_12258,N_12276);
xnor U12379 (N_12379,N_12274,N_12251);
and U12380 (N_12380,N_12179,N_12255);
and U12381 (N_12381,N_12316,N_12261);
xor U12382 (N_12382,N_12223,N_12219);
or U12383 (N_12383,N_12287,N_12245);
or U12384 (N_12384,N_12220,N_12197);
xnor U12385 (N_12385,N_12271,N_12312);
nand U12386 (N_12386,N_12191,N_12171);
xor U12387 (N_12387,N_12217,N_12240);
or U12388 (N_12388,N_12280,N_12183);
nand U12389 (N_12389,N_12277,N_12308);
nor U12390 (N_12390,N_12313,N_12164);
nor U12391 (N_12391,N_12273,N_12259);
and U12392 (N_12392,N_12247,N_12285);
or U12393 (N_12393,N_12203,N_12214);
nand U12394 (N_12394,N_12170,N_12246);
and U12395 (N_12395,N_12295,N_12196);
nand U12396 (N_12396,N_12279,N_12168);
nand U12397 (N_12397,N_12199,N_12252);
xor U12398 (N_12398,N_12260,N_12236);
and U12399 (N_12399,N_12207,N_12185);
xnor U12400 (N_12400,N_12226,N_12255);
nor U12401 (N_12401,N_12203,N_12269);
nor U12402 (N_12402,N_12273,N_12189);
or U12403 (N_12403,N_12196,N_12220);
or U12404 (N_12404,N_12222,N_12178);
nand U12405 (N_12405,N_12234,N_12279);
xor U12406 (N_12406,N_12318,N_12221);
or U12407 (N_12407,N_12198,N_12282);
nand U12408 (N_12408,N_12200,N_12277);
nor U12409 (N_12409,N_12190,N_12312);
xnor U12410 (N_12410,N_12243,N_12207);
xnor U12411 (N_12411,N_12163,N_12232);
or U12412 (N_12412,N_12279,N_12303);
and U12413 (N_12413,N_12165,N_12198);
and U12414 (N_12414,N_12285,N_12284);
nor U12415 (N_12415,N_12276,N_12177);
and U12416 (N_12416,N_12307,N_12309);
nor U12417 (N_12417,N_12160,N_12308);
nand U12418 (N_12418,N_12304,N_12306);
nor U12419 (N_12419,N_12201,N_12256);
and U12420 (N_12420,N_12253,N_12174);
xor U12421 (N_12421,N_12218,N_12287);
xnor U12422 (N_12422,N_12165,N_12317);
nor U12423 (N_12423,N_12248,N_12164);
nand U12424 (N_12424,N_12221,N_12212);
nand U12425 (N_12425,N_12189,N_12297);
nand U12426 (N_12426,N_12167,N_12193);
and U12427 (N_12427,N_12162,N_12276);
nor U12428 (N_12428,N_12203,N_12232);
or U12429 (N_12429,N_12260,N_12250);
xnor U12430 (N_12430,N_12218,N_12309);
and U12431 (N_12431,N_12311,N_12293);
nand U12432 (N_12432,N_12239,N_12213);
nand U12433 (N_12433,N_12311,N_12162);
or U12434 (N_12434,N_12263,N_12235);
nor U12435 (N_12435,N_12256,N_12226);
nor U12436 (N_12436,N_12289,N_12183);
and U12437 (N_12437,N_12259,N_12214);
nor U12438 (N_12438,N_12186,N_12177);
xor U12439 (N_12439,N_12263,N_12176);
or U12440 (N_12440,N_12228,N_12237);
or U12441 (N_12441,N_12192,N_12232);
nand U12442 (N_12442,N_12251,N_12283);
nor U12443 (N_12443,N_12306,N_12206);
nor U12444 (N_12444,N_12205,N_12191);
nor U12445 (N_12445,N_12245,N_12189);
xor U12446 (N_12446,N_12196,N_12188);
and U12447 (N_12447,N_12216,N_12169);
nor U12448 (N_12448,N_12255,N_12274);
xnor U12449 (N_12449,N_12177,N_12311);
and U12450 (N_12450,N_12175,N_12220);
nor U12451 (N_12451,N_12234,N_12299);
or U12452 (N_12452,N_12197,N_12185);
nand U12453 (N_12453,N_12297,N_12250);
or U12454 (N_12454,N_12166,N_12190);
xor U12455 (N_12455,N_12255,N_12233);
nand U12456 (N_12456,N_12315,N_12240);
and U12457 (N_12457,N_12166,N_12218);
nand U12458 (N_12458,N_12185,N_12315);
xor U12459 (N_12459,N_12303,N_12179);
nor U12460 (N_12460,N_12319,N_12244);
xnor U12461 (N_12461,N_12192,N_12254);
nor U12462 (N_12462,N_12220,N_12268);
xnor U12463 (N_12463,N_12203,N_12237);
xnor U12464 (N_12464,N_12175,N_12186);
nand U12465 (N_12465,N_12227,N_12231);
or U12466 (N_12466,N_12297,N_12197);
or U12467 (N_12467,N_12235,N_12266);
or U12468 (N_12468,N_12233,N_12206);
or U12469 (N_12469,N_12221,N_12293);
nand U12470 (N_12470,N_12274,N_12258);
nand U12471 (N_12471,N_12168,N_12233);
xnor U12472 (N_12472,N_12183,N_12304);
or U12473 (N_12473,N_12221,N_12312);
nor U12474 (N_12474,N_12273,N_12204);
or U12475 (N_12475,N_12191,N_12209);
xnor U12476 (N_12476,N_12219,N_12203);
nand U12477 (N_12477,N_12227,N_12309);
and U12478 (N_12478,N_12240,N_12237);
xnor U12479 (N_12479,N_12217,N_12257);
or U12480 (N_12480,N_12347,N_12475);
or U12481 (N_12481,N_12365,N_12439);
or U12482 (N_12482,N_12388,N_12399);
nor U12483 (N_12483,N_12342,N_12418);
xor U12484 (N_12484,N_12435,N_12325);
xnor U12485 (N_12485,N_12324,N_12447);
or U12486 (N_12486,N_12417,N_12355);
and U12487 (N_12487,N_12382,N_12465);
or U12488 (N_12488,N_12360,N_12460);
xor U12489 (N_12489,N_12379,N_12454);
or U12490 (N_12490,N_12459,N_12431);
nor U12491 (N_12491,N_12404,N_12366);
nand U12492 (N_12492,N_12377,N_12323);
or U12493 (N_12493,N_12478,N_12362);
and U12494 (N_12494,N_12442,N_12389);
nor U12495 (N_12495,N_12332,N_12392);
xor U12496 (N_12496,N_12443,N_12383);
or U12497 (N_12497,N_12368,N_12372);
or U12498 (N_12498,N_12353,N_12437);
or U12499 (N_12499,N_12344,N_12341);
xnor U12500 (N_12500,N_12462,N_12423);
or U12501 (N_12501,N_12376,N_12411);
nand U12502 (N_12502,N_12381,N_12410);
nand U12503 (N_12503,N_12412,N_12452);
and U12504 (N_12504,N_12384,N_12338);
nor U12505 (N_12505,N_12407,N_12340);
or U12506 (N_12506,N_12331,N_12430);
or U12507 (N_12507,N_12432,N_12337);
xnor U12508 (N_12508,N_12415,N_12390);
nor U12509 (N_12509,N_12424,N_12468);
nor U12510 (N_12510,N_12322,N_12428);
nand U12511 (N_12511,N_12393,N_12326);
or U12512 (N_12512,N_12472,N_12354);
xnor U12513 (N_12513,N_12409,N_12334);
xnor U12514 (N_12514,N_12479,N_12446);
and U12515 (N_12515,N_12473,N_12345);
nand U12516 (N_12516,N_12466,N_12364);
nand U12517 (N_12517,N_12413,N_12385);
and U12518 (N_12518,N_12421,N_12370);
nor U12519 (N_12519,N_12330,N_12441);
and U12520 (N_12520,N_12335,N_12358);
nand U12521 (N_12521,N_12422,N_12438);
xnor U12522 (N_12522,N_12350,N_12343);
and U12523 (N_12523,N_12451,N_12425);
xnor U12524 (N_12524,N_12416,N_12361);
or U12525 (N_12525,N_12455,N_12434);
and U12526 (N_12526,N_12426,N_12394);
and U12527 (N_12527,N_12433,N_12348);
or U12528 (N_12528,N_12321,N_12464);
nand U12529 (N_12529,N_12320,N_12357);
xor U12530 (N_12530,N_12386,N_12477);
nor U12531 (N_12531,N_12396,N_12374);
nand U12532 (N_12532,N_12378,N_12397);
and U12533 (N_12533,N_12402,N_12403);
xor U12534 (N_12534,N_12380,N_12359);
or U12535 (N_12535,N_12391,N_12440);
or U12536 (N_12536,N_12429,N_12327);
and U12537 (N_12537,N_12329,N_12367);
xor U12538 (N_12538,N_12474,N_12458);
nand U12539 (N_12539,N_12476,N_12436);
nand U12540 (N_12540,N_12471,N_12448);
nor U12541 (N_12541,N_12450,N_12444);
or U12542 (N_12542,N_12333,N_12339);
or U12543 (N_12543,N_12387,N_12467);
xnor U12544 (N_12544,N_12469,N_12414);
or U12545 (N_12545,N_12346,N_12336);
nor U12546 (N_12546,N_12369,N_12420);
xor U12547 (N_12547,N_12375,N_12470);
or U12548 (N_12548,N_12463,N_12405);
xor U12549 (N_12549,N_12449,N_12408);
or U12550 (N_12550,N_12461,N_12328);
or U12551 (N_12551,N_12419,N_12456);
xnor U12552 (N_12552,N_12395,N_12351);
or U12553 (N_12553,N_12349,N_12401);
nand U12554 (N_12554,N_12427,N_12373);
or U12555 (N_12555,N_12356,N_12371);
and U12556 (N_12556,N_12400,N_12363);
and U12557 (N_12557,N_12406,N_12453);
xnor U12558 (N_12558,N_12445,N_12457);
nor U12559 (N_12559,N_12352,N_12398);
or U12560 (N_12560,N_12413,N_12453);
or U12561 (N_12561,N_12384,N_12375);
xor U12562 (N_12562,N_12323,N_12479);
and U12563 (N_12563,N_12355,N_12455);
nand U12564 (N_12564,N_12472,N_12330);
or U12565 (N_12565,N_12461,N_12367);
nor U12566 (N_12566,N_12371,N_12414);
xor U12567 (N_12567,N_12467,N_12361);
or U12568 (N_12568,N_12360,N_12473);
nor U12569 (N_12569,N_12380,N_12372);
nor U12570 (N_12570,N_12437,N_12379);
or U12571 (N_12571,N_12454,N_12404);
and U12572 (N_12572,N_12361,N_12457);
nor U12573 (N_12573,N_12368,N_12402);
xor U12574 (N_12574,N_12453,N_12345);
nand U12575 (N_12575,N_12433,N_12332);
and U12576 (N_12576,N_12437,N_12325);
and U12577 (N_12577,N_12345,N_12432);
xor U12578 (N_12578,N_12447,N_12326);
and U12579 (N_12579,N_12431,N_12392);
xor U12580 (N_12580,N_12387,N_12345);
xor U12581 (N_12581,N_12448,N_12346);
and U12582 (N_12582,N_12370,N_12331);
and U12583 (N_12583,N_12413,N_12467);
nor U12584 (N_12584,N_12433,N_12390);
xor U12585 (N_12585,N_12423,N_12391);
nor U12586 (N_12586,N_12382,N_12400);
nor U12587 (N_12587,N_12443,N_12358);
xnor U12588 (N_12588,N_12456,N_12327);
nor U12589 (N_12589,N_12438,N_12374);
nand U12590 (N_12590,N_12464,N_12455);
or U12591 (N_12591,N_12471,N_12449);
and U12592 (N_12592,N_12351,N_12328);
nand U12593 (N_12593,N_12440,N_12410);
nand U12594 (N_12594,N_12456,N_12472);
xnor U12595 (N_12595,N_12424,N_12377);
xor U12596 (N_12596,N_12330,N_12366);
xor U12597 (N_12597,N_12361,N_12372);
xor U12598 (N_12598,N_12385,N_12429);
or U12599 (N_12599,N_12372,N_12433);
and U12600 (N_12600,N_12372,N_12443);
and U12601 (N_12601,N_12408,N_12369);
and U12602 (N_12602,N_12408,N_12335);
and U12603 (N_12603,N_12347,N_12324);
and U12604 (N_12604,N_12334,N_12475);
and U12605 (N_12605,N_12412,N_12328);
and U12606 (N_12606,N_12419,N_12471);
or U12607 (N_12607,N_12427,N_12414);
nor U12608 (N_12608,N_12405,N_12387);
nor U12609 (N_12609,N_12351,N_12326);
or U12610 (N_12610,N_12432,N_12423);
nand U12611 (N_12611,N_12329,N_12375);
and U12612 (N_12612,N_12348,N_12445);
nor U12613 (N_12613,N_12361,N_12432);
and U12614 (N_12614,N_12408,N_12415);
xor U12615 (N_12615,N_12461,N_12435);
nor U12616 (N_12616,N_12427,N_12452);
nand U12617 (N_12617,N_12445,N_12479);
xor U12618 (N_12618,N_12421,N_12442);
xor U12619 (N_12619,N_12326,N_12452);
xor U12620 (N_12620,N_12476,N_12429);
xor U12621 (N_12621,N_12375,N_12376);
nand U12622 (N_12622,N_12405,N_12397);
nor U12623 (N_12623,N_12334,N_12351);
nand U12624 (N_12624,N_12378,N_12373);
or U12625 (N_12625,N_12403,N_12442);
or U12626 (N_12626,N_12424,N_12445);
and U12627 (N_12627,N_12422,N_12443);
or U12628 (N_12628,N_12327,N_12425);
nand U12629 (N_12629,N_12371,N_12460);
or U12630 (N_12630,N_12371,N_12336);
and U12631 (N_12631,N_12394,N_12346);
or U12632 (N_12632,N_12462,N_12427);
or U12633 (N_12633,N_12339,N_12365);
and U12634 (N_12634,N_12363,N_12395);
and U12635 (N_12635,N_12456,N_12374);
and U12636 (N_12636,N_12474,N_12396);
or U12637 (N_12637,N_12454,N_12457);
xor U12638 (N_12638,N_12368,N_12445);
nor U12639 (N_12639,N_12323,N_12453);
and U12640 (N_12640,N_12622,N_12592);
xor U12641 (N_12641,N_12638,N_12582);
or U12642 (N_12642,N_12557,N_12480);
nand U12643 (N_12643,N_12564,N_12634);
or U12644 (N_12644,N_12586,N_12496);
xnor U12645 (N_12645,N_12539,N_12517);
nor U12646 (N_12646,N_12519,N_12533);
xor U12647 (N_12647,N_12520,N_12594);
xnor U12648 (N_12648,N_12572,N_12508);
nor U12649 (N_12649,N_12621,N_12581);
or U12650 (N_12650,N_12552,N_12525);
and U12651 (N_12651,N_12513,N_12512);
or U12652 (N_12652,N_12498,N_12534);
xor U12653 (N_12653,N_12567,N_12573);
nand U12654 (N_12654,N_12492,N_12529);
and U12655 (N_12655,N_12614,N_12509);
and U12656 (N_12656,N_12635,N_12576);
and U12657 (N_12657,N_12531,N_12486);
xor U12658 (N_12658,N_12597,N_12605);
or U12659 (N_12659,N_12488,N_12495);
nor U12660 (N_12660,N_12629,N_12503);
and U12661 (N_12661,N_12616,N_12639);
nand U12662 (N_12662,N_12506,N_12575);
nor U12663 (N_12663,N_12627,N_12545);
xnor U12664 (N_12664,N_12584,N_12504);
and U12665 (N_12665,N_12612,N_12624);
nor U12666 (N_12666,N_12499,N_12547);
nand U12667 (N_12667,N_12560,N_12631);
xor U12668 (N_12668,N_12490,N_12571);
and U12669 (N_12669,N_12628,N_12561);
and U12670 (N_12670,N_12619,N_12535);
or U12671 (N_12671,N_12523,N_12528);
nor U12672 (N_12672,N_12527,N_12483);
nor U12673 (N_12673,N_12502,N_12515);
nand U12674 (N_12674,N_12555,N_12603);
nand U12675 (N_12675,N_12518,N_12636);
xnor U12676 (N_12676,N_12497,N_12604);
nand U12677 (N_12677,N_12589,N_12630);
xnor U12678 (N_12678,N_12577,N_12568);
xor U12679 (N_12679,N_12540,N_12543);
or U12680 (N_12680,N_12611,N_12600);
nor U12681 (N_12681,N_12563,N_12632);
or U12682 (N_12682,N_12574,N_12510);
nor U12683 (N_12683,N_12532,N_12507);
nand U12684 (N_12684,N_12542,N_12615);
nand U12685 (N_12685,N_12485,N_12484);
nand U12686 (N_12686,N_12482,N_12537);
nand U12687 (N_12687,N_12613,N_12514);
nand U12688 (N_12688,N_12530,N_12585);
nand U12689 (N_12689,N_12544,N_12538);
and U12690 (N_12690,N_12566,N_12494);
nor U12691 (N_12691,N_12601,N_12580);
nor U12692 (N_12692,N_12610,N_12562);
nand U12693 (N_12693,N_12618,N_12607);
xnor U12694 (N_12694,N_12599,N_12536);
or U12695 (N_12695,N_12521,N_12620);
or U12696 (N_12696,N_12501,N_12598);
and U12697 (N_12697,N_12556,N_12541);
and U12698 (N_12698,N_12522,N_12550);
nor U12699 (N_12699,N_12565,N_12596);
xor U12700 (N_12700,N_12590,N_12587);
and U12701 (N_12701,N_12511,N_12493);
nand U12702 (N_12702,N_12553,N_12558);
nand U12703 (N_12703,N_12625,N_12608);
nor U12704 (N_12704,N_12551,N_12637);
or U12705 (N_12705,N_12505,N_12595);
nand U12706 (N_12706,N_12602,N_12516);
xor U12707 (N_12707,N_12617,N_12491);
nand U12708 (N_12708,N_12549,N_12570);
or U12709 (N_12709,N_12569,N_12583);
nor U12710 (N_12710,N_12489,N_12591);
or U12711 (N_12711,N_12626,N_12524);
and U12712 (N_12712,N_12546,N_12548);
and U12713 (N_12713,N_12578,N_12481);
nand U12714 (N_12714,N_12606,N_12633);
and U12715 (N_12715,N_12609,N_12526);
nand U12716 (N_12716,N_12554,N_12593);
or U12717 (N_12717,N_12500,N_12623);
nand U12718 (N_12718,N_12487,N_12588);
xnor U12719 (N_12719,N_12559,N_12579);
nand U12720 (N_12720,N_12621,N_12517);
nor U12721 (N_12721,N_12556,N_12609);
nor U12722 (N_12722,N_12571,N_12546);
and U12723 (N_12723,N_12612,N_12594);
nor U12724 (N_12724,N_12548,N_12622);
xnor U12725 (N_12725,N_12614,N_12505);
or U12726 (N_12726,N_12639,N_12562);
nor U12727 (N_12727,N_12485,N_12538);
or U12728 (N_12728,N_12550,N_12495);
xnor U12729 (N_12729,N_12520,N_12588);
and U12730 (N_12730,N_12632,N_12604);
and U12731 (N_12731,N_12599,N_12532);
xnor U12732 (N_12732,N_12537,N_12589);
or U12733 (N_12733,N_12562,N_12549);
and U12734 (N_12734,N_12610,N_12592);
and U12735 (N_12735,N_12501,N_12633);
or U12736 (N_12736,N_12584,N_12520);
and U12737 (N_12737,N_12590,N_12525);
nand U12738 (N_12738,N_12534,N_12493);
nand U12739 (N_12739,N_12489,N_12558);
and U12740 (N_12740,N_12497,N_12530);
and U12741 (N_12741,N_12532,N_12498);
nor U12742 (N_12742,N_12561,N_12599);
or U12743 (N_12743,N_12517,N_12606);
or U12744 (N_12744,N_12589,N_12503);
and U12745 (N_12745,N_12544,N_12534);
or U12746 (N_12746,N_12576,N_12528);
and U12747 (N_12747,N_12515,N_12629);
and U12748 (N_12748,N_12533,N_12497);
nand U12749 (N_12749,N_12576,N_12517);
nor U12750 (N_12750,N_12627,N_12579);
and U12751 (N_12751,N_12583,N_12606);
or U12752 (N_12752,N_12638,N_12603);
nor U12753 (N_12753,N_12585,N_12485);
or U12754 (N_12754,N_12621,N_12494);
nor U12755 (N_12755,N_12527,N_12628);
nor U12756 (N_12756,N_12601,N_12484);
or U12757 (N_12757,N_12498,N_12588);
or U12758 (N_12758,N_12590,N_12606);
nor U12759 (N_12759,N_12590,N_12544);
nand U12760 (N_12760,N_12500,N_12600);
nand U12761 (N_12761,N_12568,N_12604);
and U12762 (N_12762,N_12596,N_12508);
or U12763 (N_12763,N_12609,N_12615);
nor U12764 (N_12764,N_12555,N_12615);
nand U12765 (N_12765,N_12524,N_12583);
or U12766 (N_12766,N_12572,N_12624);
nor U12767 (N_12767,N_12626,N_12556);
or U12768 (N_12768,N_12606,N_12555);
nand U12769 (N_12769,N_12568,N_12633);
nand U12770 (N_12770,N_12523,N_12618);
xnor U12771 (N_12771,N_12505,N_12539);
nand U12772 (N_12772,N_12488,N_12590);
and U12773 (N_12773,N_12529,N_12497);
nand U12774 (N_12774,N_12556,N_12596);
or U12775 (N_12775,N_12601,N_12522);
nand U12776 (N_12776,N_12493,N_12607);
and U12777 (N_12777,N_12586,N_12621);
and U12778 (N_12778,N_12571,N_12628);
xnor U12779 (N_12779,N_12621,N_12495);
xor U12780 (N_12780,N_12587,N_12589);
and U12781 (N_12781,N_12609,N_12558);
or U12782 (N_12782,N_12557,N_12527);
or U12783 (N_12783,N_12533,N_12594);
nor U12784 (N_12784,N_12542,N_12600);
nand U12785 (N_12785,N_12501,N_12531);
or U12786 (N_12786,N_12564,N_12568);
nand U12787 (N_12787,N_12614,N_12557);
nand U12788 (N_12788,N_12528,N_12554);
and U12789 (N_12789,N_12534,N_12558);
nand U12790 (N_12790,N_12584,N_12635);
nor U12791 (N_12791,N_12634,N_12492);
xnor U12792 (N_12792,N_12518,N_12608);
nand U12793 (N_12793,N_12583,N_12568);
or U12794 (N_12794,N_12518,N_12496);
nand U12795 (N_12795,N_12480,N_12493);
nand U12796 (N_12796,N_12493,N_12535);
and U12797 (N_12797,N_12539,N_12585);
nand U12798 (N_12798,N_12531,N_12562);
and U12799 (N_12799,N_12605,N_12582);
and U12800 (N_12800,N_12732,N_12769);
and U12801 (N_12801,N_12695,N_12692);
nor U12802 (N_12802,N_12758,N_12781);
xor U12803 (N_12803,N_12735,N_12661);
xor U12804 (N_12804,N_12724,N_12680);
xor U12805 (N_12805,N_12737,N_12651);
or U12806 (N_12806,N_12646,N_12792);
or U12807 (N_12807,N_12678,N_12754);
xnor U12808 (N_12808,N_12702,N_12765);
nand U12809 (N_12809,N_12757,N_12772);
xnor U12810 (N_12810,N_12684,N_12753);
and U12811 (N_12811,N_12731,N_12768);
and U12812 (N_12812,N_12743,N_12783);
xor U12813 (N_12813,N_12688,N_12668);
nand U12814 (N_12814,N_12700,N_12762);
xor U12815 (N_12815,N_12701,N_12773);
or U12816 (N_12816,N_12752,N_12725);
and U12817 (N_12817,N_12777,N_12664);
nand U12818 (N_12818,N_12694,N_12687);
xor U12819 (N_12819,N_12744,N_12713);
nand U12820 (N_12820,N_12763,N_12658);
nand U12821 (N_12821,N_12789,N_12677);
nand U12822 (N_12822,N_12727,N_12775);
nand U12823 (N_12823,N_12642,N_12730);
or U12824 (N_12824,N_12793,N_12721);
nand U12825 (N_12825,N_12690,N_12653);
xor U12826 (N_12826,N_12720,N_12794);
nor U12827 (N_12827,N_12797,N_12640);
nor U12828 (N_12828,N_12656,N_12662);
nand U12829 (N_12829,N_12670,N_12708);
nand U12830 (N_12830,N_12747,N_12696);
nand U12831 (N_12831,N_12699,N_12799);
nand U12832 (N_12832,N_12649,N_12673);
and U12833 (N_12833,N_12739,N_12709);
and U12834 (N_12834,N_12648,N_12676);
xor U12835 (N_12835,N_12756,N_12693);
nor U12836 (N_12836,N_12736,N_12738);
or U12837 (N_12837,N_12654,N_12645);
or U12838 (N_12838,N_12717,N_12679);
or U12839 (N_12839,N_12712,N_12660);
nand U12840 (N_12840,N_12665,N_12726);
nand U12841 (N_12841,N_12719,N_12760);
or U12842 (N_12842,N_12766,N_12667);
nor U12843 (N_12843,N_12674,N_12671);
or U12844 (N_12844,N_12787,N_12655);
or U12845 (N_12845,N_12788,N_12776);
nand U12846 (N_12846,N_12710,N_12740);
nand U12847 (N_12847,N_12782,N_12750);
nand U12848 (N_12848,N_12759,N_12659);
nor U12849 (N_12849,N_12669,N_12644);
nor U12850 (N_12850,N_12697,N_12657);
nand U12851 (N_12851,N_12683,N_12729);
and U12852 (N_12852,N_12796,N_12795);
nand U12853 (N_12853,N_12666,N_12650);
or U12854 (N_12854,N_12698,N_12748);
and U12855 (N_12855,N_12675,N_12705);
and U12856 (N_12856,N_12785,N_12790);
xor U12857 (N_12857,N_12741,N_12761);
or U12858 (N_12858,N_12641,N_12746);
and U12859 (N_12859,N_12652,N_12718);
nor U12860 (N_12860,N_12755,N_12704);
xor U12861 (N_12861,N_12663,N_12647);
xor U12862 (N_12862,N_12733,N_12767);
nor U12863 (N_12863,N_12722,N_12742);
and U12864 (N_12864,N_12716,N_12751);
and U12865 (N_12865,N_12791,N_12672);
or U12866 (N_12866,N_12703,N_12778);
nand U12867 (N_12867,N_12691,N_12745);
xnor U12868 (N_12868,N_12734,N_12681);
or U12869 (N_12869,N_12689,N_12714);
xnor U12870 (N_12870,N_12780,N_12728);
nand U12871 (N_12871,N_12764,N_12770);
xnor U12872 (N_12872,N_12771,N_12779);
nor U12873 (N_12873,N_12749,N_12686);
xor U12874 (N_12874,N_12682,N_12711);
nand U12875 (N_12875,N_12798,N_12784);
xor U12876 (N_12876,N_12715,N_12774);
nor U12877 (N_12877,N_12707,N_12786);
nand U12878 (N_12878,N_12643,N_12706);
nor U12879 (N_12879,N_12685,N_12723);
and U12880 (N_12880,N_12693,N_12671);
nand U12881 (N_12881,N_12657,N_12738);
nand U12882 (N_12882,N_12671,N_12655);
xor U12883 (N_12883,N_12696,N_12764);
and U12884 (N_12884,N_12739,N_12716);
and U12885 (N_12885,N_12680,N_12656);
xor U12886 (N_12886,N_12684,N_12747);
nor U12887 (N_12887,N_12707,N_12717);
xnor U12888 (N_12888,N_12708,N_12684);
and U12889 (N_12889,N_12799,N_12750);
and U12890 (N_12890,N_12759,N_12702);
and U12891 (N_12891,N_12763,N_12786);
nor U12892 (N_12892,N_12737,N_12754);
xnor U12893 (N_12893,N_12790,N_12741);
nand U12894 (N_12894,N_12669,N_12677);
xor U12895 (N_12895,N_12748,N_12726);
nor U12896 (N_12896,N_12766,N_12640);
or U12897 (N_12897,N_12659,N_12643);
nor U12898 (N_12898,N_12777,N_12773);
and U12899 (N_12899,N_12667,N_12781);
nand U12900 (N_12900,N_12769,N_12685);
nand U12901 (N_12901,N_12650,N_12772);
xor U12902 (N_12902,N_12712,N_12679);
or U12903 (N_12903,N_12746,N_12749);
or U12904 (N_12904,N_12658,N_12694);
or U12905 (N_12905,N_12711,N_12766);
nor U12906 (N_12906,N_12673,N_12758);
nor U12907 (N_12907,N_12648,N_12787);
xnor U12908 (N_12908,N_12647,N_12701);
and U12909 (N_12909,N_12647,N_12749);
nor U12910 (N_12910,N_12671,N_12683);
nor U12911 (N_12911,N_12729,N_12767);
nand U12912 (N_12912,N_12799,N_12676);
and U12913 (N_12913,N_12711,N_12756);
nand U12914 (N_12914,N_12736,N_12732);
nor U12915 (N_12915,N_12778,N_12715);
nand U12916 (N_12916,N_12727,N_12792);
nor U12917 (N_12917,N_12796,N_12700);
xor U12918 (N_12918,N_12708,N_12674);
xnor U12919 (N_12919,N_12773,N_12760);
or U12920 (N_12920,N_12778,N_12645);
nand U12921 (N_12921,N_12652,N_12776);
and U12922 (N_12922,N_12686,N_12740);
nand U12923 (N_12923,N_12713,N_12737);
and U12924 (N_12924,N_12663,N_12651);
nor U12925 (N_12925,N_12784,N_12740);
nor U12926 (N_12926,N_12689,N_12645);
nand U12927 (N_12927,N_12797,N_12700);
nor U12928 (N_12928,N_12663,N_12683);
and U12929 (N_12929,N_12769,N_12764);
or U12930 (N_12930,N_12751,N_12695);
and U12931 (N_12931,N_12771,N_12753);
or U12932 (N_12932,N_12688,N_12785);
or U12933 (N_12933,N_12767,N_12764);
xor U12934 (N_12934,N_12728,N_12771);
xnor U12935 (N_12935,N_12753,N_12791);
and U12936 (N_12936,N_12657,N_12648);
nand U12937 (N_12937,N_12792,N_12715);
and U12938 (N_12938,N_12791,N_12705);
or U12939 (N_12939,N_12739,N_12791);
nor U12940 (N_12940,N_12767,N_12678);
or U12941 (N_12941,N_12686,N_12711);
or U12942 (N_12942,N_12645,N_12757);
and U12943 (N_12943,N_12691,N_12685);
and U12944 (N_12944,N_12704,N_12667);
nand U12945 (N_12945,N_12768,N_12759);
nor U12946 (N_12946,N_12646,N_12644);
xnor U12947 (N_12947,N_12794,N_12703);
and U12948 (N_12948,N_12742,N_12733);
or U12949 (N_12949,N_12747,N_12649);
xor U12950 (N_12950,N_12756,N_12785);
xor U12951 (N_12951,N_12692,N_12709);
nor U12952 (N_12952,N_12768,N_12718);
or U12953 (N_12953,N_12677,N_12680);
xor U12954 (N_12954,N_12701,N_12771);
nand U12955 (N_12955,N_12641,N_12654);
nand U12956 (N_12956,N_12718,N_12641);
xnor U12957 (N_12957,N_12711,N_12678);
nor U12958 (N_12958,N_12774,N_12797);
nor U12959 (N_12959,N_12676,N_12675);
nor U12960 (N_12960,N_12869,N_12951);
or U12961 (N_12961,N_12919,N_12959);
and U12962 (N_12962,N_12880,N_12938);
nor U12963 (N_12963,N_12818,N_12836);
xnor U12964 (N_12964,N_12826,N_12930);
nor U12965 (N_12965,N_12851,N_12939);
xnor U12966 (N_12966,N_12865,N_12823);
nand U12967 (N_12967,N_12936,N_12843);
xor U12968 (N_12968,N_12834,N_12840);
xnor U12969 (N_12969,N_12849,N_12956);
nand U12970 (N_12970,N_12872,N_12871);
or U12971 (N_12971,N_12803,N_12879);
nand U12972 (N_12972,N_12888,N_12902);
nand U12973 (N_12973,N_12864,N_12924);
and U12974 (N_12974,N_12910,N_12855);
or U12975 (N_12975,N_12937,N_12922);
and U12976 (N_12976,N_12921,N_12848);
nor U12977 (N_12977,N_12926,N_12868);
nor U12978 (N_12978,N_12893,N_12897);
nand U12979 (N_12979,N_12933,N_12911);
or U12980 (N_12980,N_12819,N_12891);
and U12981 (N_12981,N_12882,N_12809);
xnor U12982 (N_12982,N_12870,N_12808);
or U12983 (N_12983,N_12906,N_12905);
and U12984 (N_12984,N_12908,N_12913);
nor U12985 (N_12985,N_12916,N_12917);
xor U12986 (N_12986,N_12954,N_12896);
or U12987 (N_12987,N_12867,N_12831);
or U12988 (N_12988,N_12943,N_12935);
xor U12989 (N_12989,N_12806,N_12932);
or U12990 (N_12990,N_12815,N_12941);
nor U12991 (N_12991,N_12885,N_12950);
nor U12992 (N_12992,N_12949,N_12846);
xor U12993 (N_12993,N_12861,N_12862);
xnor U12994 (N_12994,N_12925,N_12946);
or U12995 (N_12995,N_12915,N_12947);
or U12996 (N_12996,N_12820,N_12801);
nor U12997 (N_12997,N_12898,N_12907);
and U12998 (N_12998,N_12838,N_12927);
xor U12999 (N_12999,N_12904,N_12845);
and U13000 (N_13000,N_12873,N_12827);
xnor U13001 (N_13001,N_12912,N_12828);
xnor U13002 (N_13002,N_12875,N_12802);
or U13003 (N_13003,N_12929,N_12816);
nor U13004 (N_13004,N_12811,N_12854);
nand U13005 (N_13005,N_12884,N_12940);
or U13006 (N_13006,N_12813,N_12881);
nor U13007 (N_13007,N_12842,N_12886);
nor U13008 (N_13008,N_12953,N_12858);
nor U13009 (N_13009,N_12957,N_12899);
and U13010 (N_13010,N_12945,N_12914);
nor U13011 (N_13011,N_12835,N_12853);
nand U13012 (N_13012,N_12856,N_12895);
and U13013 (N_13013,N_12800,N_12909);
or U13014 (N_13014,N_12807,N_12900);
nand U13015 (N_13015,N_12890,N_12874);
nand U13016 (N_13016,N_12850,N_12889);
nor U13017 (N_13017,N_12901,N_12923);
xor U13018 (N_13018,N_12859,N_12837);
nor U13019 (N_13019,N_12866,N_12844);
xor U13020 (N_13020,N_12952,N_12825);
and U13021 (N_13021,N_12894,N_12822);
xnor U13022 (N_13022,N_12830,N_12928);
nand U13023 (N_13023,N_12852,N_12817);
or U13024 (N_13024,N_12920,N_12812);
xor U13025 (N_13025,N_12944,N_12810);
and U13026 (N_13026,N_12942,N_12804);
or U13027 (N_13027,N_12955,N_12824);
and U13028 (N_13028,N_12839,N_12892);
xor U13029 (N_13029,N_12918,N_12887);
nand U13030 (N_13030,N_12805,N_12814);
and U13031 (N_13031,N_12847,N_12876);
nand U13032 (N_13032,N_12841,N_12877);
nor U13033 (N_13033,N_12829,N_12958);
nand U13034 (N_13034,N_12948,N_12931);
xor U13035 (N_13035,N_12863,N_12832);
nand U13036 (N_13036,N_12878,N_12821);
nor U13037 (N_13037,N_12934,N_12860);
or U13038 (N_13038,N_12833,N_12883);
xnor U13039 (N_13039,N_12903,N_12857);
nand U13040 (N_13040,N_12900,N_12953);
or U13041 (N_13041,N_12940,N_12839);
xor U13042 (N_13042,N_12911,N_12827);
xor U13043 (N_13043,N_12819,N_12810);
xnor U13044 (N_13044,N_12943,N_12921);
xor U13045 (N_13045,N_12836,N_12941);
nor U13046 (N_13046,N_12938,N_12890);
or U13047 (N_13047,N_12816,N_12883);
nand U13048 (N_13048,N_12867,N_12895);
and U13049 (N_13049,N_12818,N_12842);
nor U13050 (N_13050,N_12809,N_12876);
nand U13051 (N_13051,N_12859,N_12833);
nand U13052 (N_13052,N_12843,N_12935);
or U13053 (N_13053,N_12857,N_12890);
or U13054 (N_13054,N_12812,N_12872);
nor U13055 (N_13055,N_12927,N_12865);
or U13056 (N_13056,N_12873,N_12942);
nand U13057 (N_13057,N_12855,N_12866);
or U13058 (N_13058,N_12899,N_12834);
xnor U13059 (N_13059,N_12909,N_12931);
nand U13060 (N_13060,N_12913,N_12818);
xor U13061 (N_13061,N_12916,N_12864);
or U13062 (N_13062,N_12843,N_12922);
and U13063 (N_13063,N_12826,N_12823);
xnor U13064 (N_13064,N_12917,N_12818);
or U13065 (N_13065,N_12942,N_12818);
xor U13066 (N_13066,N_12855,N_12900);
nor U13067 (N_13067,N_12808,N_12849);
or U13068 (N_13068,N_12844,N_12831);
and U13069 (N_13069,N_12885,N_12931);
or U13070 (N_13070,N_12802,N_12926);
or U13071 (N_13071,N_12925,N_12896);
nand U13072 (N_13072,N_12946,N_12936);
or U13073 (N_13073,N_12800,N_12910);
nand U13074 (N_13074,N_12934,N_12932);
and U13075 (N_13075,N_12845,N_12932);
nand U13076 (N_13076,N_12935,N_12871);
nor U13077 (N_13077,N_12899,N_12941);
xor U13078 (N_13078,N_12881,N_12876);
and U13079 (N_13079,N_12880,N_12886);
nor U13080 (N_13080,N_12828,N_12928);
nand U13081 (N_13081,N_12866,N_12828);
nand U13082 (N_13082,N_12823,N_12939);
xor U13083 (N_13083,N_12883,N_12904);
or U13084 (N_13084,N_12824,N_12917);
nand U13085 (N_13085,N_12856,N_12957);
or U13086 (N_13086,N_12864,N_12818);
nand U13087 (N_13087,N_12847,N_12813);
nand U13088 (N_13088,N_12847,N_12857);
xnor U13089 (N_13089,N_12916,N_12882);
or U13090 (N_13090,N_12949,N_12854);
nand U13091 (N_13091,N_12830,N_12889);
nand U13092 (N_13092,N_12828,N_12825);
nor U13093 (N_13093,N_12808,N_12812);
nand U13094 (N_13094,N_12933,N_12923);
xor U13095 (N_13095,N_12912,N_12845);
and U13096 (N_13096,N_12911,N_12851);
or U13097 (N_13097,N_12867,N_12950);
xnor U13098 (N_13098,N_12935,N_12805);
or U13099 (N_13099,N_12880,N_12924);
nand U13100 (N_13100,N_12934,N_12881);
or U13101 (N_13101,N_12828,N_12845);
or U13102 (N_13102,N_12853,N_12812);
nor U13103 (N_13103,N_12943,N_12959);
and U13104 (N_13104,N_12804,N_12857);
nor U13105 (N_13105,N_12938,N_12846);
nor U13106 (N_13106,N_12940,N_12816);
or U13107 (N_13107,N_12828,N_12931);
nand U13108 (N_13108,N_12831,N_12908);
xor U13109 (N_13109,N_12820,N_12809);
and U13110 (N_13110,N_12835,N_12956);
nand U13111 (N_13111,N_12864,N_12808);
or U13112 (N_13112,N_12836,N_12896);
xnor U13113 (N_13113,N_12927,N_12855);
nor U13114 (N_13114,N_12804,N_12949);
nor U13115 (N_13115,N_12913,N_12925);
and U13116 (N_13116,N_12893,N_12856);
xnor U13117 (N_13117,N_12959,N_12862);
and U13118 (N_13118,N_12860,N_12806);
nor U13119 (N_13119,N_12919,N_12916);
or U13120 (N_13120,N_13045,N_13042);
nor U13121 (N_13121,N_13038,N_12976);
xor U13122 (N_13122,N_13071,N_13028);
nor U13123 (N_13123,N_13021,N_12968);
and U13124 (N_13124,N_13111,N_13067);
xor U13125 (N_13125,N_13010,N_13017);
nor U13126 (N_13126,N_12987,N_13109);
nor U13127 (N_13127,N_12990,N_13002);
and U13128 (N_13128,N_13074,N_13020);
and U13129 (N_13129,N_13029,N_12997);
or U13130 (N_13130,N_12974,N_12971);
nor U13131 (N_13131,N_13064,N_13057);
or U13132 (N_13132,N_13079,N_13014);
or U13133 (N_13133,N_13087,N_12994);
nor U13134 (N_13134,N_13030,N_13023);
and U13135 (N_13135,N_13117,N_13015);
nand U13136 (N_13136,N_13085,N_13037);
xor U13137 (N_13137,N_12978,N_12999);
xnor U13138 (N_13138,N_13033,N_13056);
nand U13139 (N_13139,N_13073,N_13040);
nor U13140 (N_13140,N_13086,N_12964);
or U13141 (N_13141,N_13006,N_13102);
nand U13142 (N_13142,N_13105,N_13092);
or U13143 (N_13143,N_12977,N_12984);
and U13144 (N_13144,N_13065,N_13022);
or U13145 (N_13145,N_13052,N_13082);
or U13146 (N_13146,N_13068,N_13093);
and U13147 (N_13147,N_13054,N_12996);
xor U13148 (N_13148,N_12966,N_13115);
or U13149 (N_13149,N_13053,N_12970);
or U13150 (N_13150,N_13066,N_13043);
and U13151 (N_13151,N_13027,N_12995);
xor U13152 (N_13152,N_12975,N_12982);
and U13153 (N_13153,N_13100,N_13091);
and U13154 (N_13154,N_13113,N_13083);
xnor U13155 (N_13155,N_12993,N_13069);
xor U13156 (N_13156,N_13110,N_13070);
xnor U13157 (N_13157,N_13118,N_13024);
and U13158 (N_13158,N_13098,N_12963);
and U13159 (N_13159,N_13039,N_13089);
or U13160 (N_13160,N_13101,N_13012);
xor U13161 (N_13161,N_13047,N_13032);
xor U13162 (N_13162,N_13019,N_12991);
xor U13163 (N_13163,N_13007,N_13011);
nand U13164 (N_13164,N_13031,N_12981);
nand U13165 (N_13165,N_12980,N_12961);
nand U13166 (N_13166,N_12973,N_13097);
nand U13167 (N_13167,N_13060,N_13075);
or U13168 (N_13168,N_12969,N_12979);
xnor U13169 (N_13169,N_13063,N_13084);
nand U13170 (N_13170,N_13050,N_13081);
and U13171 (N_13171,N_13090,N_13016);
xnor U13172 (N_13172,N_13003,N_13041);
and U13173 (N_13173,N_12985,N_13072);
nor U13174 (N_13174,N_12988,N_12960);
nand U13175 (N_13175,N_13059,N_13008);
or U13176 (N_13176,N_13077,N_12965);
and U13177 (N_13177,N_13108,N_13005);
nor U13178 (N_13178,N_13062,N_13046);
nand U13179 (N_13179,N_13026,N_12998);
and U13180 (N_13180,N_13088,N_13078);
and U13181 (N_13181,N_13107,N_13049);
nand U13182 (N_13182,N_13035,N_13048);
nor U13183 (N_13183,N_13080,N_13114);
nand U13184 (N_13184,N_13094,N_13013);
nand U13185 (N_13185,N_13004,N_13104);
or U13186 (N_13186,N_13051,N_13116);
nand U13187 (N_13187,N_12983,N_13001);
nand U13188 (N_13188,N_13009,N_13095);
xor U13189 (N_13189,N_13055,N_12989);
nor U13190 (N_13190,N_13119,N_13076);
nor U13191 (N_13191,N_13061,N_12962);
nand U13192 (N_13192,N_13034,N_12967);
nand U13193 (N_13193,N_13018,N_12972);
and U13194 (N_13194,N_12992,N_13096);
nand U13195 (N_13195,N_13025,N_13058);
xor U13196 (N_13196,N_13103,N_13106);
or U13197 (N_13197,N_13036,N_13099);
nor U13198 (N_13198,N_12986,N_13044);
nor U13199 (N_13199,N_13112,N_13000);
nand U13200 (N_13200,N_13016,N_13066);
or U13201 (N_13201,N_12990,N_13034);
and U13202 (N_13202,N_13033,N_12961);
nand U13203 (N_13203,N_13068,N_13040);
or U13204 (N_13204,N_13078,N_12994);
and U13205 (N_13205,N_13098,N_13087);
xor U13206 (N_13206,N_13073,N_12979);
and U13207 (N_13207,N_12998,N_13105);
xnor U13208 (N_13208,N_13009,N_13080);
and U13209 (N_13209,N_13014,N_13066);
xor U13210 (N_13210,N_13046,N_13096);
nor U13211 (N_13211,N_12976,N_13017);
xnor U13212 (N_13212,N_13117,N_13061);
nand U13213 (N_13213,N_13077,N_13074);
nand U13214 (N_13214,N_13001,N_13018);
nor U13215 (N_13215,N_13012,N_13042);
xnor U13216 (N_13216,N_13079,N_13066);
nor U13217 (N_13217,N_13060,N_13041);
nand U13218 (N_13218,N_13042,N_12965);
nand U13219 (N_13219,N_13116,N_13073);
and U13220 (N_13220,N_13081,N_12992);
xnor U13221 (N_13221,N_12985,N_13055);
and U13222 (N_13222,N_13106,N_13101);
nor U13223 (N_13223,N_13083,N_12970);
xor U13224 (N_13224,N_12997,N_13077);
nor U13225 (N_13225,N_12996,N_12977);
and U13226 (N_13226,N_12960,N_12968);
xnor U13227 (N_13227,N_13072,N_12993);
or U13228 (N_13228,N_13009,N_13049);
nor U13229 (N_13229,N_13069,N_12986);
and U13230 (N_13230,N_13026,N_13115);
nand U13231 (N_13231,N_13019,N_13087);
nand U13232 (N_13232,N_13088,N_13057);
nor U13233 (N_13233,N_12979,N_12968);
nor U13234 (N_13234,N_13014,N_13018);
nor U13235 (N_13235,N_13091,N_13093);
nor U13236 (N_13236,N_13099,N_13118);
xor U13237 (N_13237,N_13084,N_13114);
nor U13238 (N_13238,N_13025,N_13045);
nand U13239 (N_13239,N_13034,N_13064);
and U13240 (N_13240,N_13115,N_13119);
or U13241 (N_13241,N_13027,N_13099);
nand U13242 (N_13242,N_13039,N_13027);
nor U13243 (N_13243,N_13019,N_13039);
and U13244 (N_13244,N_12977,N_13048);
and U13245 (N_13245,N_13025,N_13047);
xor U13246 (N_13246,N_13071,N_12991);
nand U13247 (N_13247,N_13076,N_13007);
and U13248 (N_13248,N_13083,N_12996);
or U13249 (N_13249,N_12963,N_13092);
nor U13250 (N_13250,N_12965,N_12983);
and U13251 (N_13251,N_12986,N_13009);
and U13252 (N_13252,N_13003,N_13086);
xnor U13253 (N_13253,N_13032,N_13019);
nand U13254 (N_13254,N_13027,N_13043);
xnor U13255 (N_13255,N_12961,N_12977);
nor U13256 (N_13256,N_12979,N_13040);
nor U13257 (N_13257,N_13002,N_12967);
and U13258 (N_13258,N_12996,N_13063);
or U13259 (N_13259,N_13115,N_13106);
and U13260 (N_13260,N_13013,N_13113);
and U13261 (N_13261,N_13024,N_12982);
nand U13262 (N_13262,N_13007,N_13113);
xor U13263 (N_13263,N_12968,N_13010);
and U13264 (N_13264,N_13046,N_13004);
nor U13265 (N_13265,N_12973,N_12980);
nor U13266 (N_13266,N_13060,N_12965);
nand U13267 (N_13267,N_13075,N_13033);
or U13268 (N_13268,N_12984,N_13064);
and U13269 (N_13269,N_13089,N_13008);
or U13270 (N_13270,N_13108,N_13054);
or U13271 (N_13271,N_12961,N_12976);
nand U13272 (N_13272,N_13049,N_13048);
or U13273 (N_13273,N_13057,N_13046);
or U13274 (N_13274,N_13072,N_13085);
nand U13275 (N_13275,N_13050,N_13080);
nor U13276 (N_13276,N_13087,N_13055);
nand U13277 (N_13277,N_12967,N_12987);
nor U13278 (N_13278,N_13030,N_13009);
or U13279 (N_13279,N_13005,N_13015);
and U13280 (N_13280,N_13243,N_13274);
xor U13281 (N_13281,N_13279,N_13164);
and U13282 (N_13282,N_13188,N_13230);
xnor U13283 (N_13283,N_13218,N_13269);
xnor U13284 (N_13284,N_13227,N_13175);
or U13285 (N_13285,N_13237,N_13263);
or U13286 (N_13286,N_13273,N_13196);
or U13287 (N_13287,N_13204,N_13177);
nor U13288 (N_13288,N_13180,N_13264);
xnor U13289 (N_13289,N_13223,N_13252);
xor U13290 (N_13290,N_13125,N_13161);
nor U13291 (N_13291,N_13130,N_13202);
or U13292 (N_13292,N_13143,N_13261);
and U13293 (N_13293,N_13228,N_13244);
or U13294 (N_13294,N_13212,N_13179);
and U13295 (N_13295,N_13197,N_13141);
or U13296 (N_13296,N_13253,N_13201);
and U13297 (N_13297,N_13216,N_13186);
nor U13298 (N_13298,N_13126,N_13185);
or U13299 (N_13299,N_13147,N_13142);
and U13300 (N_13300,N_13128,N_13240);
and U13301 (N_13301,N_13238,N_13149);
nand U13302 (N_13302,N_13184,N_13123);
and U13303 (N_13303,N_13157,N_13174);
xnor U13304 (N_13304,N_13138,N_13209);
nor U13305 (N_13305,N_13135,N_13159);
nor U13306 (N_13306,N_13162,N_13275);
or U13307 (N_13307,N_13277,N_13156);
or U13308 (N_13308,N_13122,N_13272);
nand U13309 (N_13309,N_13158,N_13163);
and U13310 (N_13310,N_13231,N_13239);
and U13311 (N_13311,N_13134,N_13267);
xor U13312 (N_13312,N_13246,N_13245);
nand U13313 (N_13313,N_13259,N_13262);
or U13314 (N_13314,N_13127,N_13194);
and U13315 (N_13315,N_13225,N_13133);
xnor U13316 (N_13316,N_13256,N_13121);
nor U13317 (N_13317,N_13229,N_13171);
nand U13318 (N_13318,N_13233,N_13129);
or U13319 (N_13319,N_13144,N_13270);
or U13320 (N_13320,N_13205,N_13195);
and U13321 (N_13321,N_13221,N_13160);
and U13322 (N_13322,N_13211,N_13213);
nand U13323 (N_13323,N_13187,N_13170);
nand U13324 (N_13324,N_13132,N_13120);
and U13325 (N_13325,N_13247,N_13203);
or U13326 (N_13326,N_13235,N_13241);
or U13327 (N_13327,N_13136,N_13276);
or U13328 (N_13328,N_13219,N_13131);
nand U13329 (N_13329,N_13266,N_13190);
nor U13330 (N_13330,N_13260,N_13154);
nand U13331 (N_13331,N_13207,N_13139);
or U13332 (N_13332,N_13220,N_13155);
or U13333 (N_13333,N_13182,N_13208);
or U13334 (N_13334,N_13145,N_13140);
and U13335 (N_13335,N_13257,N_13224);
xnor U13336 (N_13336,N_13222,N_13258);
and U13337 (N_13337,N_13193,N_13150);
nand U13338 (N_13338,N_13192,N_13217);
nand U13339 (N_13339,N_13172,N_13178);
and U13340 (N_13340,N_13232,N_13199);
or U13341 (N_13341,N_13226,N_13198);
and U13342 (N_13342,N_13167,N_13278);
nor U13343 (N_13343,N_13242,N_13255);
or U13344 (N_13344,N_13169,N_13210);
xor U13345 (N_13345,N_13214,N_13168);
or U13346 (N_13346,N_13148,N_13173);
nand U13347 (N_13347,N_13146,N_13234);
or U13348 (N_13348,N_13271,N_13176);
nor U13349 (N_13349,N_13268,N_13189);
and U13350 (N_13350,N_13152,N_13153);
nor U13351 (N_13351,N_13215,N_13254);
and U13352 (N_13352,N_13166,N_13191);
xnor U13353 (N_13353,N_13265,N_13248);
or U13354 (N_13354,N_13183,N_13251);
nand U13355 (N_13355,N_13137,N_13250);
or U13356 (N_13356,N_13124,N_13200);
nand U13357 (N_13357,N_13165,N_13236);
or U13358 (N_13358,N_13249,N_13181);
and U13359 (N_13359,N_13206,N_13151);
nor U13360 (N_13360,N_13139,N_13153);
nor U13361 (N_13361,N_13213,N_13274);
and U13362 (N_13362,N_13248,N_13209);
xnor U13363 (N_13363,N_13164,N_13148);
and U13364 (N_13364,N_13278,N_13166);
xor U13365 (N_13365,N_13208,N_13233);
or U13366 (N_13366,N_13266,N_13129);
xor U13367 (N_13367,N_13192,N_13165);
or U13368 (N_13368,N_13205,N_13257);
xor U13369 (N_13369,N_13230,N_13194);
or U13370 (N_13370,N_13249,N_13182);
and U13371 (N_13371,N_13279,N_13195);
nor U13372 (N_13372,N_13134,N_13198);
xor U13373 (N_13373,N_13264,N_13273);
nor U13374 (N_13374,N_13250,N_13161);
and U13375 (N_13375,N_13252,N_13175);
xnor U13376 (N_13376,N_13174,N_13176);
nand U13377 (N_13377,N_13266,N_13207);
nor U13378 (N_13378,N_13136,N_13150);
xnor U13379 (N_13379,N_13243,N_13255);
xnor U13380 (N_13380,N_13263,N_13161);
nor U13381 (N_13381,N_13136,N_13263);
and U13382 (N_13382,N_13166,N_13181);
xnor U13383 (N_13383,N_13143,N_13173);
or U13384 (N_13384,N_13139,N_13225);
nor U13385 (N_13385,N_13212,N_13206);
or U13386 (N_13386,N_13142,N_13272);
or U13387 (N_13387,N_13127,N_13218);
or U13388 (N_13388,N_13145,N_13134);
nor U13389 (N_13389,N_13186,N_13207);
nor U13390 (N_13390,N_13137,N_13178);
or U13391 (N_13391,N_13202,N_13120);
and U13392 (N_13392,N_13124,N_13249);
or U13393 (N_13393,N_13156,N_13264);
nor U13394 (N_13394,N_13197,N_13223);
nand U13395 (N_13395,N_13251,N_13181);
xnor U13396 (N_13396,N_13219,N_13158);
or U13397 (N_13397,N_13126,N_13181);
and U13398 (N_13398,N_13168,N_13164);
xor U13399 (N_13399,N_13192,N_13173);
nand U13400 (N_13400,N_13212,N_13245);
or U13401 (N_13401,N_13270,N_13194);
and U13402 (N_13402,N_13139,N_13171);
and U13403 (N_13403,N_13217,N_13141);
and U13404 (N_13404,N_13246,N_13144);
and U13405 (N_13405,N_13135,N_13276);
or U13406 (N_13406,N_13145,N_13257);
or U13407 (N_13407,N_13268,N_13217);
and U13408 (N_13408,N_13142,N_13171);
xor U13409 (N_13409,N_13173,N_13279);
nor U13410 (N_13410,N_13279,N_13152);
and U13411 (N_13411,N_13237,N_13267);
or U13412 (N_13412,N_13194,N_13271);
xnor U13413 (N_13413,N_13191,N_13151);
or U13414 (N_13414,N_13272,N_13230);
nor U13415 (N_13415,N_13164,N_13261);
nand U13416 (N_13416,N_13189,N_13135);
nand U13417 (N_13417,N_13268,N_13141);
nand U13418 (N_13418,N_13275,N_13207);
and U13419 (N_13419,N_13141,N_13160);
nor U13420 (N_13420,N_13135,N_13241);
nor U13421 (N_13421,N_13171,N_13232);
xor U13422 (N_13422,N_13190,N_13171);
and U13423 (N_13423,N_13130,N_13266);
or U13424 (N_13424,N_13275,N_13246);
nor U13425 (N_13425,N_13253,N_13121);
nand U13426 (N_13426,N_13229,N_13238);
nand U13427 (N_13427,N_13170,N_13204);
and U13428 (N_13428,N_13167,N_13196);
nor U13429 (N_13429,N_13178,N_13231);
nor U13430 (N_13430,N_13133,N_13239);
or U13431 (N_13431,N_13224,N_13262);
and U13432 (N_13432,N_13266,N_13145);
and U13433 (N_13433,N_13180,N_13140);
xor U13434 (N_13434,N_13177,N_13126);
nand U13435 (N_13435,N_13187,N_13182);
xor U13436 (N_13436,N_13127,N_13262);
or U13437 (N_13437,N_13217,N_13178);
nor U13438 (N_13438,N_13201,N_13267);
and U13439 (N_13439,N_13232,N_13212);
xnor U13440 (N_13440,N_13424,N_13350);
nand U13441 (N_13441,N_13397,N_13374);
xnor U13442 (N_13442,N_13319,N_13349);
or U13443 (N_13443,N_13309,N_13431);
xnor U13444 (N_13444,N_13291,N_13436);
and U13445 (N_13445,N_13351,N_13318);
or U13446 (N_13446,N_13299,N_13387);
nand U13447 (N_13447,N_13286,N_13377);
or U13448 (N_13448,N_13434,N_13415);
xnor U13449 (N_13449,N_13308,N_13385);
nand U13450 (N_13450,N_13358,N_13307);
nand U13451 (N_13451,N_13406,N_13362);
xor U13452 (N_13452,N_13315,N_13298);
and U13453 (N_13453,N_13322,N_13371);
nand U13454 (N_13454,N_13336,N_13342);
nor U13455 (N_13455,N_13414,N_13425);
nor U13456 (N_13456,N_13394,N_13365);
and U13457 (N_13457,N_13381,N_13301);
nand U13458 (N_13458,N_13320,N_13380);
xnor U13459 (N_13459,N_13430,N_13398);
and U13460 (N_13460,N_13302,N_13413);
xnor U13461 (N_13461,N_13373,N_13366);
nand U13462 (N_13462,N_13417,N_13403);
xnor U13463 (N_13463,N_13348,N_13405);
nand U13464 (N_13464,N_13344,N_13388);
nor U13465 (N_13465,N_13422,N_13324);
xor U13466 (N_13466,N_13321,N_13343);
xnor U13467 (N_13467,N_13331,N_13392);
nor U13468 (N_13468,N_13339,N_13347);
or U13469 (N_13469,N_13345,N_13416);
xnor U13470 (N_13470,N_13390,N_13295);
xnor U13471 (N_13471,N_13384,N_13376);
xnor U13472 (N_13472,N_13341,N_13312);
nor U13473 (N_13473,N_13297,N_13420);
and U13474 (N_13474,N_13310,N_13429);
xor U13475 (N_13475,N_13379,N_13328);
xnor U13476 (N_13476,N_13411,N_13316);
xor U13477 (N_13477,N_13294,N_13332);
or U13478 (N_13478,N_13360,N_13372);
nor U13479 (N_13479,N_13367,N_13402);
nor U13480 (N_13480,N_13382,N_13433);
or U13481 (N_13481,N_13437,N_13323);
or U13482 (N_13482,N_13346,N_13306);
xor U13483 (N_13483,N_13407,N_13404);
and U13484 (N_13484,N_13325,N_13293);
nand U13485 (N_13485,N_13427,N_13399);
xor U13486 (N_13486,N_13335,N_13330);
and U13487 (N_13487,N_13300,N_13311);
nor U13488 (N_13488,N_13354,N_13340);
or U13489 (N_13489,N_13359,N_13401);
nor U13490 (N_13490,N_13428,N_13280);
and U13491 (N_13491,N_13288,N_13412);
and U13492 (N_13492,N_13419,N_13285);
and U13493 (N_13493,N_13410,N_13408);
xor U13494 (N_13494,N_13395,N_13304);
nor U13495 (N_13495,N_13370,N_13368);
and U13496 (N_13496,N_13375,N_13426);
and U13497 (N_13497,N_13303,N_13421);
nand U13498 (N_13498,N_13355,N_13389);
xnor U13499 (N_13499,N_13400,N_13313);
xor U13500 (N_13500,N_13391,N_13296);
nor U13501 (N_13501,N_13423,N_13338);
or U13502 (N_13502,N_13292,N_13438);
xnor U13503 (N_13503,N_13386,N_13334);
nor U13504 (N_13504,N_13287,N_13364);
or U13505 (N_13505,N_13326,N_13396);
nand U13506 (N_13506,N_13383,N_13290);
xnor U13507 (N_13507,N_13283,N_13363);
nand U13508 (N_13508,N_13393,N_13352);
nor U13509 (N_13509,N_13282,N_13361);
and U13510 (N_13510,N_13327,N_13439);
nand U13511 (N_13511,N_13337,N_13356);
xnor U13512 (N_13512,N_13317,N_13432);
xnor U13513 (N_13513,N_13369,N_13333);
or U13514 (N_13514,N_13435,N_13329);
nor U13515 (N_13515,N_13357,N_13281);
nand U13516 (N_13516,N_13378,N_13418);
or U13517 (N_13517,N_13284,N_13305);
or U13518 (N_13518,N_13314,N_13353);
and U13519 (N_13519,N_13289,N_13409);
nor U13520 (N_13520,N_13298,N_13393);
or U13521 (N_13521,N_13287,N_13345);
and U13522 (N_13522,N_13325,N_13351);
nand U13523 (N_13523,N_13410,N_13345);
xnor U13524 (N_13524,N_13401,N_13381);
or U13525 (N_13525,N_13387,N_13332);
xor U13526 (N_13526,N_13317,N_13335);
nand U13527 (N_13527,N_13388,N_13386);
or U13528 (N_13528,N_13393,N_13342);
or U13529 (N_13529,N_13343,N_13330);
nor U13530 (N_13530,N_13280,N_13348);
xnor U13531 (N_13531,N_13408,N_13359);
xor U13532 (N_13532,N_13405,N_13434);
nor U13533 (N_13533,N_13281,N_13358);
nor U13534 (N_13534,N_13380,N_13337);
or U13535 (N_13535,N_13379,N_13290);
nand U13536 (N_13536,N_13415,N_13338);
nand U13537 (N_13537,N_13367,N_13322);
nor U13538 (N_13538,N_13357,N_13422);
nand U13539 (N_13539,N_13334,N_13424);
or U13540 (N_13540,N_13333,N_13427);
xnor U13541 (N_13541,N_13288,N_13384);
or U13542 (N_13542,N_13321,N_13421);
or U13543 (N_13543,N_13386,N_13409);
nand U13544 (N_13544,N_13383,N_13292);
or U13545 (N_13545,N_13280,N_13335);
and U13546 (N_13546,N_13339,N_13395);
and U13547 (N_13547,N_13298,N_13314);
and U13548 (N_13548,N_13363,N_13342);
xor U13549 (N_13549,N_13347,N_13295);
nand U13550 (N_13550,N_13368,N_13295);
and U13551 (N_13551,N_13334,N_13360);
nor U13552 (N_13552,N_13358,N_13334);
xnor U13553 (N_13553,N_13410,N_13412);
nor U13554 (N_13554,N_13429,N_13288);
or U13555 (N_13555,N_13315,N_13324);
xnor U13556 (N_13556,N_13402,N_13436);
nor U13557 (N_13557,N_13292,N_13299);
nand U13558 (N_13558,N_13337,N_13344);
nor U13559 (N_13559,N_13408,N_13422);
xor U13560 (N_13560,N_13303,N_13416);
and U13561 (N_13561,N_13385,N_13309);
xnor U13562 (N_13562,N_13307,N_13431);
and U13563 (N_13563,N_13383,N_13323);
and U13564 (N_13564,N_13402,N_13419);
nor U13565 (N_13565,N_13427,N_13374);
or U13566 (N_13566,N_13348,N_13367);
or U13567 (N_13567,N_13356,N_13303);
and U13568 (N_13568,N_13405,N_13400);
or U13569 (N_13569,N_13403,N_13381);
xor U13570 (N_13570,N_13346,N_13290);
xnor U13571 (N_13571,N_13358,N_13338);
nor U13572 (N_13572,N_13325,N_13391);
nor U13573 (N_13573,N_13437,N_13384);
nand U13574 (N_13574,N_13388,N_13331);
nand U13575 (N_13575,N_13439,N_13352);
or U13576 (N_13576,N_13383,N_13386);
xnor U13577 (N_13577,N_13430,N_13418);
xor U13578 (N_13578,N_13370,N_13308);
nand U13579 (N_13579,N_13431,N_13390);
nor U13580 (N_13580,N_13316,N_13332);
xor U13581 (N_13581,N_13395,N_13373);
nand U13582 (N_13582,N_13388,N_13351);
xnor U13583 (N_13583,N_13293,N_13364);
and U13584 (N_13584,N_13422,N_13367);
nor U13585 (N_13585,N_13299,N_13397);
and U13586 (N_13586,N_13325,N_13350);
and U13587 (N_13587,N_13343,N_13357);
or U13588 (N_13588,N_13427,N_13354);
or U13589 (N_13589,N_13401,N_13382);
nor U13590 (N_13590,N_13397,N_13377);
nor U13591 (N_13591,N_13422,N_13321);
nor U13592 (N_13592,N_13357,N_13432);
nor U13593 (N_13593,N_13362,N_13341);
and U13594 (N_13594,N_13383,N_13408);
or U13595 (N_13595,N_13310,N_13295);
xor U13596 (N_13596,N_13382,N_13282);
xnor U13597 (N_13597,N_13312,N_13330);
or U13598 (N_13598,N_13369,N_13395);
and U13599 (N_13599,N_13352,N_13304);
or U13600 (N_13600,N_13585,N_13557);
nand U13601 (N_13601,N_13442,N_13470);
nand U13602 (N_13602,N_13576,N_13502);
nor U13603 (N_13603,N_13541,N_13507);
nor U13604 (N_13604,N_13465,N_13569);
nand U13605 (N_13605,N_13511,N_13530);
xor U13606 (N_13606,N_13538,N_13531);
xnor U13607 (N_13607,N_13566,N_13529);
or U13608 (N_13608,N_13524,N_13527);
xnor U13609 (N_13609,N_13452,N_13488);
and U13610 (N_13610,N_13533,N_13514);
xor U13611 (N_13611,N_13461,N_13448);
nor U13612 (N_13612,N_13560,N_13500);
nor U13613 (N_13613,N_13484,N_13464);
xnor U13614 (N_13614,N_13476,N_13532);
or U13615 (N_13615,N_13462,N_13449);
xnor U13616 (N_13616,N_13493,N_13592);
nor U13617 (N_13617,N_13572,N_13558);
and U13618 (N_13618,N_13504,N_13547);
or U13619 (N_13619,N_13595,N_13505);
nand U13620 (N_13620,N_13551,N_13479);
nor U13621 (N_13621,N_13591,N_13463);
xor U13622 (N_13622,N_13480,N_13517);
xnor U13623 (N_13623,N_13542,N_13478);
and U13624 (N_13624,N_13586,N_13496);
and U13625 (N_13625,N_13486,N_13506);
or U13626 (N_13626,N_13444,N_13467);
nor U13627 (N_13627,N_13447,N_13581);
or U13628 (N_13628,N_13473,N_13509);
or U13629 (N_13629,N_13573,N_13575);
or U13630 (N_13630,N_13440,N_13446);
xor U13631 (N_13631,N_13582,N_13598);
or U13632 (N_13632,N_13535,N_13590);
xor U13633 (N_13633,N_13534,N_13503);
and U13634 (N_13634,N_13552,N_13489);
xor U13635 (N_13635,N_13564,N_13498);
and U13636 (N_13636,N_13519,N_13565);
and U13637 (N_13637,N_13583,N_13491);
nand U13638 (N_13638,N_13578,N_13597);
xnor U13639 (N_13639,N_13510,N_13522);
and U13640 (N_13640,N_13520,N_13453);
or U13641 (N_13641,N_13483,N_13475);
xor U13642 (N_13642,N_13587,N_13471);
xnor U13643 (N_13643,N_13482,N_13589);
nand U13644 (N_13644,N_13574,N_13457);
nand U13645 (N_13645,N_13513,N_13580);
and U13646 (N_13646,N_13523,N_13540);
nor U13647 (N_13647,N_13554,N_13481);
and U13648 (N_13648,N_13495,N_13594);
nand U13649 (N_13649,N_13570,N_13521);
nor U13650 (N_13650,N_13454,N_13460);
or U13651 (N_13651,N_13472,N_13545);
nand U13652 (N_13652,N_13567,N_13588);
xnor U13653 (N_13653,N_13456,N_13512);
nor U13654 (N_13654,N_13526,N_13562);
xnor U13655 (N_13655,N_13458,N_13490);
nor U13656 (N_13656,N_13474,N_13443);
xnor U13657 (N_13657,N_13441,N_13543);
nor U13658 (N_13658,N_13599,N_13579);
or U13659 (N_13659,N_13593,N_13596);
nand U13660 (N_13660,N_13518,N_13508);
nor U13661 (N_13661,N_13556,N_13563);
or U13662 (N_13662,N_13499,N_13497);
or U13663 (N_13663,N_13528,N_13485);
nand U13664 (N_13664,N_13536,N_13455);
nand U13665 (N_13665,N_13516,N_13544);
and U13666 (N_13666,N_13515,N_13501);
nor U13667 (N_13667,N_13561,N_13568);
and U13668 (N_13668,N_13553,N_13466);
xnor U13669 (N_13669,N_13468,N_13571);
nor U13670 (N_13670,N_13577,N_13450);
or U13671 (N_13671,N_13555,N_13525);
xor U13672 (N_13672,N_13539,N_13537);
nand U13673 (N_13673,N_13549,N_13546);
xnor U13674 (N_13674,N_13548,N_13492);
and U13675 (N_13675,N_13487,N_13459);
nor U13676 (N_13676,N_13584,N_13559);
and U13677 (N_13677,N_13477,N_13445);
nor U13678 (N_13678,N_13494,N_13451);
and U13679 (N_13679,N_13550,N_13469);
or U13680 (N_13680,N_13561,N_13500);
and U13681 (N_13681,N_13540,N_13476);
nand U13682 (N_13682,N_13485,N_13483);
xnor U13683 (N_13683,N_13478,N_13495);
xor U13684 (N_13684,N_13460,N_13466);
xor U13685 (N_13685,N_13467,N_13523);
nor U13686 (N_13686,N_13465,N_13499);
or U13687 (N_13687,N_13551,N_13591);
nand U13688 (N_13688,N_13512,N_13509);
xor U13689 (N_13689,N_13582,N_13586);
or U13690 (N_13690,N_13590,N_13598);
xor U13691 (N_13691,N_13470,N_13473);
nand U13692 (N_13692,N_13543,N_13485);
or U13693 (N_13693,N_13505,N_13559);
nand U13694 (N_13694,N_13516,N_13515);
nand U13695 (N_13695,N_13588,N_13526);
nand U13696 (N_13696,N_13569,N_13477);
and U13697 (N_13697,N_13455,N_13494);
nand U13698 (N_13698,N_13522,N_13580);
nand U13699 (N_13699,N_13455,N_13443);
nand U13700 (N_13700,N_13591,N_13509);
or U13701 (N_13701,N_13575,N_13552);
xnor U13702 (N_13702,N_13597,N_13461);
nand U13703 (N_13703,N_13568,N_13549);
nor U13704 (N_13704,N_13443,N_13581);
xor U13705 (N_13705,N_13489,N_13556);
or U13706 (N_13706,N_13484,N_13491);
and U13707 (N_13707,N_13499,N_13515);
nand U13708 (N_13708,N_13574,N_13567);
nand U13709 (N_13709,N_13475,N_13534);
and U13710 (N_13710,N_13481,N_13582);
nand U13711 (N_13711,N_13457,N_13537);
and U13712 (N_13712,N_13474,N_13453);
or U13713 (N_13713,N_13581,N_13448);
xor U13714 (N_13714,N_13594,N_13571);
nand U13715 (N_13715,N_13540,N_13515);
and U13716 (N_13716,N_13472,N_13569);
xor U13717 (N_13717,N_13589,N_13484);
nand U13718 (N_13718,N_13512,N_13547);
xor U13719 (N_13719,N_13593,N_13564);
or U13720 (N_13720,N_13475,N_13486);
and U13721 (N_13721,N_13441,N_13475);
nand U13722 (N_13722,N_13555,N_13543);
or U13723 (N_13723,N_13456,N_13550);
or U13724 (N_13724,N_13572,N_13447);
and U13725 (N_13725,N_13579,N_13458);
nand U13726 (N_13726,N_13598,N_13587);
or U13727 (N_13727,N_13573,N_13559);
or U13728 (N_13728,N_13562,N_13582);
xor U13729 (N_13729,N_13490,N_13495);
xor U13730 (N_13730,N_13538,N_13565);
nand U13731 (N_13731,N_13460,N_13596);
nor U13732 (N_13732,N_13459,N_13594);
nor U13733 (N_13733,N_13520,N_13514);
or U13734 (N_13734,N_13479,N_13535);
xor U13735 (N_13735,N_13469,N_13492);
and U13736 (N_13736,N_13556,N_13558);
and U13737 (N_13737,N_13489,N_13468);
or U13738 (N_13738,N_13573,N_13543);
nand U13739 (N_13739,N_13442,N_13530);
nor U13740 (N_13740,N_13530,N_13588);
xnor U13741 (N_13741,N_13553,N_13479);
nor U13742 (N_13742,N_13529,N_13500);
and U13743 (N_13743,N_13445,N_13460);
xor U13744 (N_13744,N_13501,N_13511);
nor U13745 (N_13745,N_13572,N_13563);
and U13746 (N_13746,N_13511,N_13571);
and U13747 (N_13747,N_13466,N_13510);
xor U13748 (N_13748,N_13515,N_13451);
nand U13749 (N_13749,N_13503,N_13445);
xor U13750 (N_13750,N_13481,N_13558);
and U13751 (N_13751,N_13556,N_13539);
and U13752 (N_13752,N_13594,N_13502);
and U13753 (N_13753,N_13521,N_13563);
or U13754 (N_13754,N_13459,N_13519);
and U13755 (N_13755,N_13532,N_13550);
or U13756 (N_13756,N_13475,N_13554);
nand U13757 (N_13757,N_13550,N_13509);
and U13758 (N_13758,N_13584,N_13444);
or U13759 (N_13759,N_13532,N_13559);
nor U13760 (N_13760,N_13606,N_13725);
nand U13761 (N_13761,N_13737,N_13758);
xnor U13762 (N_13762,N_13636,N_13627);
and U13763 (N_13763,N_13700,N_13625);
nor U13764 (N_13764,N_13730,N_13742);
xor U13765 (N_13765,N_13718,N_13754);
and U13766 (N_13766,N_13662,N_13661);
nor U13767 (N_13767,N_13664,N_13727);
nand U13768 (N_13768,N_13663,N_13740);
or U13769 (N_13769,N_13643,N_13712);
or U13770 (N_13770,N_13668,N_13716);
nand U13771 (N_13771,N_13611,N_13691);
or U13772 (N_13772,N_13669,N_13638);
xnor U13773 (N_13773,N_13652,N_13706);
and U13774 (N_13774,N_13618,N_13679);
or U13775 (N_13775,N_13626,N_13644);
or U13776 (N_13776,N_13719,N_13702);
and U13777 (N_13777,N_13689,N_13648);
or U13778 (N_13778,N_13756,N_13646);
or U13779 (N_13779,N_13735,N_13747);
or U13780 (N_13780,N_13695,N_13757);
nor U13781 (N_13781,N_13722,N_13609);
nor U13782 (N_13782,N_13723,N_13632);
nand U13783 (N_13783,N_13721,N_13628);
xnor U13784 (N_13784,N_13635,N_13732);
xor U13785 (N_13785,N_13631,N_13741);
nor U13786 (N_13786,N_13647,N_13704);
nand U13787 (N_13787,N_13751,N_13743);
and U13788 (N_13788,N_13688,N_13600);
or U13789 (N_13789,N_13728,N_13634);
and U13790 (N_13790,N_13660,N_13642);
and U13791 (N_13791,N_13707,N_13653);
xnor U13792 (N_13792,N_13610,N_13755);
xor U13793 (N_13793,N_13602,N_13658);
and U13794 (N_13794,N_13619,N_13750);
xnor U13795 (N_13795,N_13680,N_13607);
nor U13796 (N_13796,N_13613,N_13729);
and U13797 (N_13797,N_13617,N_13711);
or U13798 (N_13798,N_13649,N_13614);
and U13799 (N_13799,N_13667,N_13734);
or U13800 (N_13800,N_13746,N_13605);
and U13801 (N_13801,N_13641,N_13612);
nor U13802 (N_13802,N_13713,N_13640);
nand U13803 (N_13803,N_13693,N_13659);
or U13804 (N_13804,N_13703,N_13745);
nor U13805 (N_13805,N_13615,N_13654);
and U13806 (N_13806,N_13645,N_13675);
or U13807 (N_13807,N_13604,N_13759);
or U13808 (N_13808,N_13637,N_13657);
or U13809 (N_13809,N_13753,N_13674);
nand U13810 (N_13810,N_13724,N_13692);
nand U13811 (N_13811,N_13714,N_13676);
xnor U13812 (N_13812,N_13687,N_13666);
and U13813 (N_13813,N_13685,N_13744);
and U13814 (N_13814,N_13651,N_13672);
and U13815 (N_13815,N_13621,N_13678);
xor U13816 (N_13816,N_13684,N_13733);
and U13817 (N_13817,N_13699,N_13720);
nor U13818 (N_13818,N_13748,N_13710);
and U13819 (N_13819,N_13731,N_13656);
nor U13820 (N_13820,N_13629,N_13682);
xor U13821 (N_13821,N_13698,N_13686);
nand U13822 (N_13822,N_13690,N_13603);
or U13823 (N_13823,N_13622,N_13696);
and U13824 (N_13824,N_13665,N_13601);
or U13825 (N_13825,N_13681,N_13749);
nor U13826 (N_13826,N_13738,N_13697);
xor U13827 (N_13827,N_13694,N_13705);
xnor U13828 (N_13828,N_13715,N_13655);
or U13829 (N_13829,N_13670,N_13633);
xnor U13830 (N_13830,N_13616,N_13752);
nand U13831 (N_13831,N_13623,N_13677);
and U13832 (N_13832,N_13608,N_13739);
nor U13833 (N_13833,N_13624,N_13683);
xnor U13834 (N_13834,N_13726,N_13736);
nand U13835 (N_13835,N_13673,N_13701);
nand U13836 (N_13836,N_13671,N_13620);
nor U13837 (N_13837,N_13630,N_13709);
xor U13838 (N_13838,N_13717,N_13650);
or U13839 (N_13839,N_13639,N_13708);
and U13840 (N_13840,N_13690,N_13727);
and U13841 (N_13841,N_13741,N_13695);
nand U13842 (N_13842,N_13613,N_13648);
and U13843 (N_13843,N_13629,N_13634);
and U13844 (N_13844,N_13624,N_13606);
xor U13845 (N_13845,N_13733,N_13644);
and U13846 (N_13846,N_13680,N_13641);
and U13847 (N_13847,N_13734,N_13728);
and U13848 (N_13848,N_13729,N_13737);
xor U13849 (N_13849,N_13690,N_13686);
and U13850 (N_13850,N_13658,N_13740);
nand U13851 (N_13851,N_13759,N_13757);
or U13852 (N_13852,N_13679,N_13753);
nand U13853 (N_13853,N_13719,N_13602);
and U13854 (N_13854,N_13601,N_13668);
nor U13855 (N_13855,N_13691,N_13616);
nor U13856 (N_13856,N_13752,N_13665);
and U13857 (N_13857,N_13713,N_13619);
or U13858 (N_13858,N_13609,N_13695);
or U13859 (N_13859,N_13646,N_13708);
or U13860 (N_13860,N_13703,N_13753);
nand U13861 (N_13861,N_13664,N_13623);
nor U13862 (N_13862,N_13733,N_13656);
or U13863 (N_13863,N_13650,N_13628);
nand U13864 (N_13864,N_13692,N_13718);
nor U13865 (N_13865,N_13756,N_13635);
and U13866 (N_13866,N_13718,N_13716);
and U13867 (N_13867,N_13713,N_13618);
and U13868 (N_13868,N_13639,N_13656);
xor U13869 (N_13869,N_13729,N_13703);
nand U13870 (N_13870,N_13610,N_13609);
xor U13871 (N_13871,N_13739,N_13728);
xor U13872 (N_13872,N_13669,N_13607);
or U13873 (N_13873,N_13751,N_13719);
or U13874 (N_13874,N_13623,N_13686);
nand U13875 (N_13875,N_13738,N_13717);
nand U13876 (N_13876,N_13745,N_13647);
nand U13877 (N_13877,N_13619,N_13643);
or U13878 (N_13878,N_13609,N_13746);
nor U13879 (N_13879,N_13694,N_13625);
and U13880 (N_13880,N_13645,N_13751);
nor U13881 (N_13881,N_13653,N_13740);
nand U13882 (N_13882,N_13743,N_13661);
nand U13883 (N_13883,N_13722,N_13632);
or U13884 (N_13884,N_13662,N_13601);
xnor U13885 (N_13885,N_13638,N_13741);
nor U13886 (N_13886,N_13752,N_13663);
nand U13887 (N_13887,N_13747,N_13626);
and U13888 (N_13888,N_13745,N_13668);
xor U13889 (N_13889,N_13702,N_13679);
xor U13890 (N_13890,N_13603,N_13661);
nor U13891 (N_13891,N_13685,N_13665);
or U13892 (N_13892,N_13758,N_13625);
nand U13893 (N_13893,N_13734,N_13683);
nand U13894 (N_13894,N_13708,N_13699);
nand U13895 (N_13895,N_13615,N_13727);
and U13896 (N_13896,N_13749,N_13655);
nand U13897 (N_13897,N_13723,N_13653);
nor U13898 (N_13898,N_13626,N_13663);
nand U13899 (N_13899,N_13756,N_13747);
and U13900 (N_13900,N_13716,N_13628);
and U13901 (N_13901,N_13749,N_13738);
or U13902 (N_13902,N_13619,N_13749);
and U13903 (N_13903,N_13749,N_13682);
nand U13904 (N_13904,N_13719,N_13643);
nand U13905 (N_13905,N_13758,N_13741);
nor U13906 (N_13906,N_13666,N_13653);
or U13907 (N_13907,N_13680,N_13639);
or U13908 (N_13908,N_13628,N_13649);
nand U13909 (N_13909,N_13686,N_13638);
and U13910 (N_13910,N_13658,N_13634);
xor U13911 (N_13911,N_13675,N_13720);
or U13912 (N_13912,N_13712,N_13639);
xor U13913 (N_13913,N_13677,N_13675);
and U13914 (N_13914,N_13729,N_13712);
nand U13915 (N_13915,N_13686,N_13613);
or U13916 (N_13916,N_13720,N_13673);
and U13917 (N_13917,N_13610,N_13679);
xnor U13918 (N_13918,N_13642,N_13623);
and U13919 (N_13919,N_13742,N_13676);
nor U13920 (N_13920,N_13853,N_13831);
nor U13921 (N_13921,N_13823,N_13821);
xnor U13922 (N_13922,N_13802,N_13832);
or U13923 (N_13923,N_13817,N_13768);
nor U13924 (N_13924,N_13837,N_13886);
and U13925 (N_13925,N_13855,N_13871);
xor U13926 (N_13926,N_13811,N_13892);
nor U13927 (N_13927,N_13891,N_13820);
or U13928 (N_13928,N_13884,N_13791);
or U13929 (N_13929,N_13833,N_13763);
nand U13930 (N_13930,N_13880,N_13919);
nor U13931 (N_13931,N_13876,N_13907);
or U13932 (N_13932,N_13801,N_13869);
nor U13933 (N_13933,N_13800,N_13819);
xnor U13934 (N_13934,N_13897,N_13864);
and U13935 (N_13935,N_13804,N_13781);
xnor U13936 (N_13936,N_13793,N_13896);
nor U13937 (N_13937,N_13900,N_13771);
nand U13938 (N_13938,N_13778,N_13822);
and U13939 (N_13939,N_13785,N_13769);
nand U13940 (N_13940,N_13824,N_13762);
and U13941 (N_13941,N_13879,N_13868);
nor U13942 (N_13942,N_13797,N_13773);
or U13943 (N_13943,N_13844,N_13874);
or U13944 (N_13944,N_13796,N_13851);
and U13945 (N_13945,N_13839,N_13915);
xor U13946 (N_13946,N_13875,N_13862);
and U13947 (N_13947,N_13794,N_13850);
nor U13948 (N_13948,N_13765,N_13901);
and U13949 (N_13949,N_13912,N_13843);
nor U13950 (N_13950,N_13898,N_13792);
xor U13951 (N_13951,N_13806,N_13865);
xor U13952 (N_13952,N_13788,N_13842);
nor U13953 (N_13953,N_13854,N_13770);
and U13954 (N_13954,N_13814,N_13836);
nand U13955 (N_13955,N_13775,N_13807);
xnor U13956 (N_13956,N_13858,N_13909);
and U13957 (N_13957,N_13908,N_13772);
nand U13958 (N_13958,N_13848,N_13910);
nor U13959 (N_13959,N_13905,N_13767);
or U13960 (N_13960,N_13913,N_13849);
or U13961 (N_13961,N_13803,N_13834);
nor U13962 (N_13962,N_13795,N_13838);
and U13963 (N_13963,N_13914,N_13877);
and U13964 (N_13964,N_13815,N_13918);
nand U13965 (N_13965,N_13826,N_13798);
xor U13966 (N_13966,N_13790,N_13873);
xnor U13967 (N_13967,N_13902,N_13818);
nor U13968 (N_13968,N_13887,N_13780);
or U13969 (N_13969,N_13888,N_13878);
nand U13970 (N_13970,N_13827,N_13894);
or U13971 (N_13971,N_13903,N_13856);
nand U13972 (N_13972,N_13809,N_13787);
xor U13973 (N_13973,N_13904,N_13860);
and U13974 (N_13974,N_13825,N_13881);
nand U13975 (N_13975,N_13766,N_13906);
nand U13976 (N_13976,N_13911,N_13761);
nor U13977 (N_13977,N_13799,N_13866);
or U13978 (N_13978,N_13840,N_13916);
nor U13979 (N_13979,N_13889,N_13841);
or U13980 (N_13980,N_13852,N_13782);
and U13981 (N_13981,N_13779,N_13861);
and U13982 (N_13982,N_13805,N_13890);
xor U13983 (N_13983,N_13870,N_13777);
xor U13984 (N_13984,N_13760,N_13830);
and U13985 (N_13985,N_13829,N_13828);
or U13986 (N_13986,N_13789,N_13917);
xor U13987 (N_13987,N_13893,N_13883);
nor U13988 (N_13988,N_13810,N_13845);
and U13989 (N_13989,N_13857,N_13872);
nor U13990 (N_13990,N_13867,N_13885);
nor U13991 (N_13991,N_13764,N_13808);
and U13992 (N_13992,N_13863,N_13812);
and U13993 (N_13993,N_13847,N_13774);
nand U13994 (N_13994,N_13813,N_13859);
xor U13995 (N_13995,N_13882,N_13899);
and U13996 (N_13996,N_13786,N_13895);
nor U13997 (N_13997,N_13816,N_13846);
or U13998 (N_13998,N_13835,N_13776);
and U13999 (N_13999,N_13783,N_13784);
xor U14000 (N_14000,N_13814,N_13888);
xor U14001 (N_14001,N_13878,N_13867);
nor U14002 (N_14002,N_13855,N_13904);
and U14003 (N_14003,N_13901,N_13814);
xor U14004 (N_14004,N_13803,N_13861);
xor U14005 (N_14005,N_13782,N_13763);
or U14006 (N_14006,N_13806,N_13835);
and U14007 (N_14007,N_13771,N_13866);
and U14008 (N_14008,N_13806,N_13889);
and U14009 (N_14009,N_13828,N_13770);
nand U14010 (N_14010,N_13766,N_13798);
and U14011 (N_14011,N_13799,N_13914);
xor U14012 (N_14012,N_13805,N_13896);
and U14013 (N_14013,N_13775,N_13911);
nor U14014 (N_14014,N_13897,N_13768);
and U14015 (N_14015,N_13839,N_13843);
or U14016 (N_14016,N_13824,N_13857);
and U14017 (N_14017,N_13846,N_13784);
and U14018 (N_14018,N_13844,N_13770);
nand U14019 (N_14019,N_13842,N_13896);
nor U14020 (N_14020,N_13765,N_13766);
or U14021 (N_14021,N_13806,N_13793);
nand U14022 (N_14022,N_13782,N_13904);
and U14023 (N_14023,N_13777,N_13798);
or U14024 (N_14024,N_13862,N_13850);
or U14025 (N_14025,N_13763,N_13911);
xor U14026 (N_14026,N_13854,N_13878);
nor U14027 (N_14027,N_13760,N_13901);
nor U14028 (N_14028,N_13781,N_13893);
xnor U14029 (N_14029,N_13819,N_13774);
or U14030 (N_14030,N_13852,N_13774);
nand U14031 (N_14031,N_13888,N_13834);
nor U14032 (N_14032,N_13882,N_13862);
nor U14033 (N_14033,N_13789,N_13881);
xor U14034 (N_14034,N_13830,N_13874);
or U14035 (N_14035,N_13784,N_13884);
nand U14036 (N_14036,N_13875,N_13869);
nor U14037 (N_14037,N_13805,N_13865);
or U14038 (N_14038,N_13763,N_13861);
nor U14039 (N_14039,N_13857,N_13891);
or U14040 (N_14040,N_13911,N_13836);
xor U14041 (N_14041,N_13870,N_13900);
or U14042 (N_14042,N_13893,N_13808);
xnor U14043 (N_14043,N_13784,N_13897);
and U14044 (N_14044,N_13776,N_13798);
nand U14045 (N_14045,N_13807,N_13821);
nand U14046 (N_14046,N_13917,N_13850);
and U14047 (N_14047,N_13899,N_13862);
or U14048 (N_14048,N_13804,N_13763);
and U14049 (N_14049,N_13896,N_13847);
nor U14050 (N_14050,N_13767,N_13790);
or U14051 (N_14051,N_13917,N_13787);
nor U14052 (N_14052,N_13894,N_13788);
nand U14053 (N_14053,N_13811,N_13855);
xnor U14054 (N_14054,N_13897,N_13820);
nand U14055 (N_14055,N_13876,N_13890);
nand U14056 (N_14056,N_13909,N_13861);
and U14057 (N_14057,N_13858,N_13837);
nand U14058 (N_14058,N_13828,N_13824);
nand U14059 (N_14059,N_13859,N_13837);
nor U14060 (N_14060,N_13908,N_13806);
xnor U14061 (N_14061,N_13884,N_13902);
and U14062 (N_14062,N_13898,N_13805);
and U14063 (N_14063,N_13773,N_13768);
and U14064 (N_14064,N_13892,N_13881);
and U14065 (N_14065,N_13843,N_13834);
nand U14066 (N_14066,N_13786,N_13788);
nand U14067 (N_14067,N_13792,N_13762);
nor U14068 (N_14068,N_13876,N_13805);
xnor U14069 (N_14069,N_13783,N_13808);
and U14070 (N_14070,N_13860,N_13828);
xnor U14071 (N_14071,N_13900,N_13783);
and U14072 (N_14072,N_13805,N_13829);
nor U14073 (N_14073,N_13777,N_13818);
nand U14074 (N_14074,N_13886,N_13843);
and U14075 (N_14075,N_13854,N_13809);
and U14076 (N_14076,N_13794,N_13821);
nand U14077 (N_14077,N_13853,N_13781);
nor U14078 (N_14078,N_13768,N_13786);
nor U14079 (N_14079,N_13803,N_13793);
nand U14080 (N_14080,N_13922,N_13951);
and U14081 (N_14081,N_13992,N_13943);
or U14082 (N_14082,N_13976,N_14047);
nand U14083 (N_14083,N_14052,N_13986);
nor U14084 (N_14084,N_14038,N_14009);
or U14085 (N_14085,N_13963,N_14027);
xor U14086 (N_14086,N_13921,N_14013);
xor U14087 (N_14087,N_13980,N_13956);
and U14088 (N_14088,N_13977,N_13979);
nor U14089 (N_14089,N_14031,N_13982);
nand U14090 (N_14090,N_14001,N_13999);
and U14091 (N_14091,N_13940,N_13944);
nand U14092 (N_14092,N_13925,N_14050);
and U14093 (N_14093,N_13991,N_14032);
xnor U14094 (N_14094,N_13981,N_14075);
nand U14095 (N_14095,N_13995,N_14014);
or U14096 (N_14096,N_13932,N_14060);
or U14097 (N_14097,N_13934,N_13936);
or U14098 (N_14098,N_14042,N_14003);
nand U14099 (N_14099,N_14073,N_14071);
or U14100 (N_14100,N_13947,N_14045);
or U14101 (N_14101,N_14062,N_13949);
or U14102 (N_14102,N_14034,N_14054);
xor U14103 (N_14103,N_14078,N_14069);
xnor U14104 (N_14104,N_13971,N_13984);
nor U14105 (N_14105,N_14019,N_14011);
or U14106 (N_14106,N_13997,N_14079);
or U14107 (N_14107,N_14051,N_14010);
and U14108 (N_14108,N_14028,N_13974);
nor U14109 (N_14109,N_13923,N_14041);
nand U14110 (N_14110,N_13929,N_14022);
and U14111 (N_14111,N_13993,N_14021);
or U14112 (N_14112,N_13973,N_14067);
or U14113 (N_14113,N_13989,N_13950);
nor U14114 (N_14114,N_13970,N_13962);
nand U14115 (N_14115,N_13958,N_14006);
xor U14116 (N_14116,N_14056,N_13969);
xor U14117 (N_14117,N_14012,N_13920);
or U14118 (N_14118,N_14077,N_14026);
and U14119 (N_14119,N_13988,N_14053);
nand U14120 (N_14120,N_14005,N_13955);
and U14121 (N_14121,N_14063,N_14035);
nand U14122 (N_14122,N_14057,N_13972);
and U14123 (N_14123,N_14037,N_14029);
xor U14124 (N_14124,N_14030,N_13959);
nor U14125 (N_14125,N_14068,N_14064);
xnor U14126 (N_14126,N_14004,N_13960);
and U14127 (N_14127,N_14033,N_13996);
or U14128 (N_14128,N_14066,N_13954);
or U14129 (N_14129,N_14074,N_13966);
xnor U14130 (N_14130,N_14055,N_13998);
or U14131 (N_14131,N_13933,N_13978);
or U14132 (N_14132,N_14017,N_13937);
nand U14133 (N_14133,N_13964,N_14072);
and U14134 (N_14134,N_13927,N_14048);
nand U14135 (N_14135,N_14036,N_14061);
or U14136 (N_14136,N_14020,N_14023);
nand U14137 (N_14137,N_13967,N_13968);
or U14138 (N_14138,N_13990,N_14065);
and U14139 (N_14139,N_14076,N_13948);
xnor U14140 (N_14140,N_13994,N_14024);
and U14141 (N_14141,N_13924,N_13952);
and U14142 (N_14142,N_13945,N_13985);
or U14143 (N_14143,N_13926,N_14018);
or U14144 (N_14144,N_14039,N_13987);
nand U14145 (N_14145,N_14025,N_14070);
or U14146 (N_14146,N_13931,N_13942);
nand U14147 (N_14147,N_14044,N_13935);
and U14148 (N_14148,N_14016,N_13975);
or U14149 (N_14149,N_13961,N_13957);
nand U14150 (N_14150,N_14049,N_13938);
nor U14151 (N_14151,N_13939,N_13965);
xnor U14152 (N_14152,N_13946,N_13928);
nand U14153 (N_14153,N_13930,N_14015);
nor U14154 (N_14154,N_14008,N_14043);
and U14155 (N_14155,N_13983,N_14007);
or U14156 (N_14156,N_14040,N_14058);
or U14157 (N_14157,N_14059,N_14000);
or U14158 (N_14158,N_13941,N_14046);
or U14159 (N_14159,N_14002,N_13953);
xnor U14160 (N_14160,N_14028,N_14007);
xor U14161 (N_14161,N_14004,N_14030);
or U14162 (N_14162,N_14061,N_14008);
nand U14163 (N_14163,N_14016,N_13957);
nand U14164 (N_14164,N_14069,N_14023);
or U14165 (N_14165,N_13963,N_13983);
and U14166 (N_14166,N_13991,N_13951);
nand U14167 (N_14167,N_13972,N_14048);
nor U14168 (N_14168,N_13993,N_14024);
nand U14169 (N_14169,N_14054,N_13922);
and U14170 (N_14170,N_13939,N_14048);
or U14171 (N_14171,N_13929,N_13948);
and U14172 (N_14172,N_13958,N_13981);
or U14173 (N_14173,N_13996,N_14055);
nor U14174 (N_14174,N_14033,N_13924);
or U14175 (N_14175,N_13929,N_13930);
nor U14176 (N_14176,N_14058,N_14069);
or U14177 (N_14177,N_13931,N_13967);
xor U14178 (N_14178,N_13958,N_14038);
nand U14179 (N_14179,N_14024,N_13931);
or U14180 (N_14180,N_13973,N_14063);
nor U14181 (N_14181,N_14044,N_14043);
and U14182 (N_14182,N_13973,N_13981);
and U14183 (N_14183,N_13960,N_14058);
xnor U14184 (N_14184,N_13929,N_13981);
nor U14185 (N_14185,N_13969,N_14001);
nor U14186 (N_14186,N_13998,N_14034);
and U14187 (N_14187,N_14000,N_14039);
nand U14188 (N_14188,N_13985,N_14040);
xnor U14189 (N_14189,N_13932,N_13946);
xnor U14190 (N_14190,N_13961,N_13967);
and U14191 (N_14191,N_13998,N_14011);
xnor U14192 (N_14192,N_14015,N_13925);
nand U14193 (N_14193,N_13941,N_13970);
or U14194 (N_14194,N_13925,N_14037);
nand U14195 (N_14195,N_14035,N_14060);
nor U14196 (N_14196,N_13986,N_13991);
and U14197 (N_14197,N_13933,N_14045);
or U14198 (N_14198,N_14014,N_13990);
and U14199 (N_14199,N_14033,N_13933);
and U14200 (N_14200,N_14009,N_13977);
nand U14201 (N_14201,N_14007,N_13948);
or U14202 (N_14202,N_14019,N_13959);
and U14203 (N_14203,N_14034,N_13936);
nand U14204 (N_14204,N_14034,N_14010);
and U14205 (N_14205,N_14051,N_14047);
xnor U14206 (N_14206,N_14067,N_14027);
nand U14207 (N_14207,N_14076,N_14048);
and U14208 (N_14208,N_14036,N_14040);
xnor U14209 (N_14209,N_13982,N_14004);
nand U14210 (N_14210,N_14076,N_14049);
and U14211 (N_14211,N_13934,N_13935);
and U14212 (N_14212,N_14013,N_14025);
xnor U14213 (N_14213,N_13967,N_14032);
or U14214 (N_14214,N_14002,N_13930);
xor U14215 (N_14215,N_13999,N_13944);
and U14216 (N_14216,N_13955,N_13998);
or U14217 (N_14217,N_13990,N_14062);
nand U14218 (N_14218,N_14040,N_13980);
and U14219 (N_14219,N_13939,N_13935);
xor U14220 (N_14220,N_14075,N_14033);
nor U14221 (N_14221,N_14003,N_14037);
xor U14222 (N_14222,N_13924,N_13987);
and U14223 (N_14223,N_14044,N_13984);
nor U14224 (N_14224,N_14074,N_13957);
nor U14225 (N_14225,N_13926,N_13922);
nand U14226 (N_14226,N_13989,N_14010);
nor U14227 (N_14227,N_14048,N_13991);
xor U14228 (N_14228,N_14054,N_14037);
or U14229 (N_14229,N_14036,N_14035);
nand U14230 (N_14230,N_14037,N_13977);
xor U14231 (N_14231,N_14037,N_13948);
and U14232 (N_14232,N_14044,N_14048);
xor U14233 (N_14233,N_13975,N_13981);
or U14234 (N_14234,N_14038,N_13930);
or U14235 (N_14235,N_13968,N_13936);
nand U14236 (N_14236,N_14045,N_13982);
or U14237 (N_14237,N_14008,N_13964);
xnor U14238 (N_14238,N_13986,N_14072);
and U14239 (N_14239,N_13986,N_14019);
and U14240 (N_14240,N_14168,N_14132);
nand U14241 (N_14241,N_14238,N_14110);
xor U14242 (N_14242,N_14081,N_14157);
nor U14243 (N_14243,N_14169,N_14189);
nand U14244 (N_14244,N_14119,N_14233);
nand U14245 (N_14245,N_14155,N_14196);
or U14246 (N_14246,N_14123,N_14236);
xor U14247 (N_14247,N_14203,N_14086);
nand U14248 (N_14248,N_14175,N_14235);
xnor U14249 (N_14249,N_14124,N_14223);
and U14250 (N_14250,N_14228,N_14122);
nor U14251 (N_14251,N_14229,N_14191);
or U14252 (N_14252,N_14093,N_14120);
nor U14253 (N_14253,N_14237,N_14161);
or U14254 (N_14254,N_14188,N_14104);
or U14255 (N_14255,N_14150,N_14116);
xor U14256 (N_14256,N_14239,N_14149);
nand U14257 (N_14257,N_14139,N_14129);
and U14258 (N_14258,N_14219,N_14231);
nor U14259 (N_14259,N_14209,N_14163);
nor U14260 (N_14260,N_14148,N_14230);
xnor U14261 (N_14261,N_14214,N_14173);
and U14262 (N_14262,N_14131,N_14181);
nand U14263 (N_14263,N_14172,N_14128);
nor U14264 (N_14264,N_14201,N_14216);
nand U14265 (N_14265,N_14108,N_14153);
or U14266 (N_14266,N_14085,N_14117);
xor U14267 (N_14267,N_14152,N_14127);
xnor U14268 (N_14268,N_14192,N_14179);
nor U14269 (N_14269,N_14178,N_14174);
nand U14270 (N_14270,N_14207,N_14082);
and U14271 (N_14271,N_14126,N_14100);
nor U14272 (N_14272,N_14227,N_14164);
nor U14273 (N_14273,N_14133,N_14107);
and U14274 (N_14274,N_14106,N_14176);
or U14275 (N_14275,N_14091,N_14193);
nor U14276 (N_14276,N_14099,N_14221);
nand U14277 (N_14277,N_14084,N_14142);
nand U14278 (N_14278,N_14205,N_14170);
nor U14279 (N_14279,N_14225,N_14103);
or U14280 (N_14280,N_14160,N_14184);
and U14281 (N_14281,N_14185,N_14159);
xor U14282 (N_14282,N_14166,N_14194);
nand U14283 (N_14283,N_14218,N_14198);
nor U14284 (N_14284,N_14141,N_14121);
nor U14285 (N_14285,N_14154,N_14226);
and U14286 (N_14286,N_14137,N_14105);
and U14287 (N_14287,N_14143,N_14115);
nor U14288 (N_14288,N_14092,N_14200);
nor U14289 (N_14289,N_14204,N_14083);
xor U14290 (N_14290,N_14140,N_14113);
or U14291 (N_14291,N_14135,N_14101);
or U14292 (N_14292,N_14199,N_14215);
and U14293 (N_14293,N_14202,N_14156);
nand U14294 (N_14294,N_14089,N_14190);
and U14295 (N_14295,N_14125,N_14102);
xnor U14296 (N_14296,N_14220,N_14096);
nor U14297 (N_14297,N_14144,N_14095);
xor U14298 (N_14298,N_14187,N_14210);
nor U14299 (N_14299,N_14145,N_14208);
nand U14300 (N_14300,N_14134,N_14167);
nor U14301 (N_14301,N_14183,N_14112);
and U14302 (N_14302,N_14136,N_14222);
or U14303 (N_14303,N_14151,N_14206);
nor U14304 (N_14304,N_14180,N_14090);
xnor U14305 (N_14305,N_14094,N_14213);
nor U14306 (N_14306,N_14171,N_14146);
nor U14307 (N_14307,N_14118,N_14158);
nand U14308 (N_14308,N_14197,N_14186);
or U14309 (N_14309,N_14114,N_14088);
nand U14310 (N_14310,N_14217,N_14130);
nor U14311 (N_14311,N_14109,N_14111);
nand U14312 (N_14312,N_14232,N_14224);
and U14313 (N_14313,N_14162,N_14165);
or U14314 (N_14314,N_14211,N_14234);
nand U14315 (N_14315,N_14138,N_14098);
or U14316 (N_14316,N_14097,N_14182);
or U14317 (N_14317,N_14177,N_14147);
nor U14318 (N_14318,N_14212,N_14080);
and U14319 (N_14319,N_14087,N_14195);
nor U14320 (N_14320,N_14165,N_14142);
xor U14321 (N_14321,N_14153,N_14169);
xor U14322 (N_14322,N_14136,N_14235);
nand U14323 (N_14323,N_14134,N_14176);
nor U14324 (N_14324,N_14104,N_14210);
and U14325 (N_14325,N_14149,N_14201);
nand U14326 (N_14326,N_14175,N_14134);
nand U14327 (N_14327,N_14135,N_14112);
nand U14328 (N_14328,N_14135,N_14109);
nor U14329 (N_14329,N_14135,N_14224);
or U14330 (N_14330,N_14135,N_14233);
nand U14331 (N_14331,N_14176,N_14227);
and U14332 (N_14332,N_14234,N_14176);
nand U14333 (N_14333,N_14163,N_14130);
nor U14334 (N_14334,N_14154,N_14150);
nand U14335 (N_14335,N_14204,N_14186);
xnor U14336 (N_14336,N_14116,N_14129);
and U14337 (N_14337,N_14098,N_14178);
or U14338 (N_14338,N_14236,N_14088);
and U14339 (N_14339,N_14200,N_14083);
nand U14340 (N_14340,N_14231,N_14181);
xor U14341 (N_14341,N_14230,N_14104);
xor U14342 (N_14342,N_14106,N_14149);
or U14343 (N_14343,N_14098,N_14173);
or U14344 (N_14344,N_14188,N_14201);
and U14345 (N_14345,N_14121,N_14127);
or U14346 (N_14346,N_14166,N_14104);
or U14347 (N_14347,N_14167,N_14145);
nor U14348 (N_14348,N_14136,N_14223);
or U14349 (N_14349,N_14170,N_14209);
or U14350 (N_14350,N_14113,N_14184);
nor U14351 (N_14351,N_14087,N_14229);
and U14352 (N_14352,N_14205,N_14189);
and U14353 (N_14353,N_14130,N_14171);
and U14354 (N_14354,N_14216,N_14180);
nor U14355 (N_14355,N_14125,N_14183);
and U14356 (N_14356,N_14204,N_14219);
xor U14357 (N_14357,N_14193,N_14202);
nor U14358 (N_14358,N_14204,N_14200);
nor U14359 (N_14359,N_14187,N_14212);
and U14360 (N_14360,N_14237,N_14215);
or U14361 (N_14361,N_14183,N_14092);
and U14362 (N_14362,N_14110,N_14183);
nand U14363 (N_14363,N_14087,N_14234);
and U14364 (N_14364,N_14190,N_14201);
nor U14365 (N_14365,N_14082,N_14231);
nor U14366 (N_14366,N_14104,N_14237);
nor U14367 (N_14367,N_14188,N_14169);
nor U14368 (N_14368,N_14113,N_14150);
nor U14369 (N_14369,N_14092,N_14150);
or U14370 (N_14370,N_14144,N_14200);
nor U14371 (N_14371,N_14121,N_14081);
xnor U14372 (N_14372,N_14135,N_14179);
or U14373 (N_14373,N_14178,N_14138);
nor U14374 (N_14374,N_14234,N_14138);
xor U14375 (N_14375,N_14081,N_14212);
nand U14376 (N_14376,N_14219,N_14120);
nand U14377 (N_14377,N_14081,N_14222);
nor U14378 (N_14378,N_14109,N_14103);
or U14379 (N_14379,N_14172,N_14206);
nor U14380 (N_14380,N_14134,N_14217);
xor U14381 (N_14381,N_14136,N_14165);
nor U14382 (N_14382,N_14217,N_14169);
nand U14383 (N_14383,N_14162,N_14100);
xor U14384 (N_14384,N_14164,N_14101);
or U14385 (N_14385,N_14090,N_14186);
xnor U14386 (N_14386,N_14196,N_14120);
or U14387 (N_14387,N_14207,N_14121);
nand U14388 (N_14388,N_14141,N_14157);
nand U14389 (N_14389,N_14117,N_14189);
and U14390 (N_14390,N_14182,N_14231);
xor U14391 (N_14391,N_14228,N_14213);
nor U14392 (N_14392,N_14127,N_14162);
nor U14393 (N_14393,N_14199,N_14133);
nand U14394 (N_14394,N_14101,N_14145);
xor U14395 (N_14395,N_14220,N_14198);
nor U14396 (N_14396,N_14128,N_14145);
and U14397 (N_14397,N_14149,N_14210);
nor U14398 (N_14398,N_14179,N_14090);
nand U14399 (N_14399,N_14170,N_14152);
xnor U14400 (N_14400,N_14339,N_14289);
nor U14401 (N_14401,N_14273,N_14367);
and U14402 (N_14402,N_14343,N_14398);
and U14403 (N_14403,N_14264,N_14313);
nand U14404 (N_14404,N_14291,N_14250);
nand U14405 (N_14405,N_14392,N_14260);
and U14406 (N_14406,N_14309,N_14316);
nor U14407 (N_14407,N_14263,N_14330);
nand U14408 (N_14408,N_14301,N_14360);
nand U14409 (N_14409,N_14268,N_14314);
or U14410 (N_14410,N_14279,N_14326);
or U14411 (N_14411,N_14303,N_14318);
or U14412 (N_14412,N_14375,N_14284);
nand U14413 (N_14413,N_14292,N_14337);
xnor U14414 (N_14414,N_14358,N_14241);
nor U14415 (N_14415,N_14278,N_14338);
nor U14416 (N_14416,N_14281,N_14370);
and U14417 (N_14417,N_14305,N_14383);
or U14418 (N_14418,N_14257,N_14288);
nand U14419 (N_14419,N_14267,N_14388);
or U14420 (N_14420,N_14340,N_14247);
and U14421 (N_14421,N_14275,N_14352);
xnor U14422 (N_14422,N_14310,N_14356);
nand U14423 (N_14423,N_14299,N_14293);
and U14424 (N_14424,N_14353,N_14245);
nand U14425 (N_14425,N_14302,N_14348);
nand U14426 (N_14426,N_14307,N_14320);
nor U14427 (N_14427,N_14324,N_14285);
nand U14428 (N_14428,N_14315,N_14361);
nor U14429 (N_14429,N_14393,N_14386);
or U14430 (N_14430,N_14248,N_14387);
nor U14431 (N_14431,N_14322,N_14395);
xor U14432 (N_14432,N_14300,N_14255);
and U14433 (N_14433,N_14365,N_14271);
nand U14434 (N_14434,N_14366,N_14252);
and U14435 (N_14435,N_14249,N_14297);
nor U14436 (N_14436,N_14378,N_14396);
or U14437 (N_14437,N_14369,N_14355);
xnor U14438 (N_14438,N_14251,N_14256);
nand U14439 (N_14439,N_14287,N_14282);
xor U14440 (N_14440,N_14244,N_14276);
and U14441 (N_14441,N_14351,N_14317);
or U14442 (N_14442,N_14384,N_14296);
and U14443 (N_14443,N_14359,N_14283);
nor U14444 (N_14444,N_14331,N_14311);
and U14445 (N_14445,N_14308,N_14328);
nand U14446 (N_14446,N_14254,N_14364);
nor U14447 (N_14447,N_14265,N_14258);
nand U14448 (N_14448,N_14261,N_14277);
nand U14449 (N_14449,N_14269,N_14399);
or U14450 (N_14450,N_14243,N_14346);
and U14451 (N_14451,N_14304,N_14336);
or U14452 (N_14452,N_14381,N_14272);
nand U14453 (N_14453,N_14357,N_14390);
nor U14454 (N_14454,N_14382,N_14345);
xnor U14455 (N_14455,N_14362,N_14349);
nand U14456 (N_14456,N_14319,N_14344);
or U14457 (N_14457,N_14306,N_14377);
xor U14458 (N_14458,N_14332,N_14373);
xnor U14459 (N_14459,N_14342,N_14323);
and U14460 (N_14460,N_14295,N_14298);
or U14461 (N_14461,N_14363,N_14372);
xnor U14462 (N_14462,N_14270,N_14327);
xor U14463 (N_14463,N_14341,N_14259);
nor U14464 (N_14464,N_14312,N_14389);
nor U14465 (N_14465,N_14379,N_14394);
or U14466 (N_14466,N_14385,N_14262);
or U14467 (N_14467,N_14368,N_14329);
nor U14468 (N_14468,N_14290,N_14354);
nor U14469 (N_14469,N_14274,N_14253);
nand U14470 (N_14470,N_14321,N_14280);
xnor U14471 (N_14471,N_14347,N_14380);
nand U14472 (N_14472,N_14325,N_14240);
xor U14473 (N_14473,N_14333,N_14391);
nand U14474 (N_14474,N_14286,N_14266);
or U14475 (N_14475,N_14350,N_14397);
nand U14476 (N_14476,N_14334,N_14371);
nand U14477 (N_14477,N_14246,N_14242);
and U14478 (N_14478,N_14376,N_14374);
or U14479 (N_14479,N_14294,N_14335);
nand U14480 (N_14480,N_14321,N_14355);
or U14481 (N_14481,N_14246,N_14385);
xnor U14482 (N_14482,N_14306,N_14369);
or U14483 (N_14483,N_14320,N_14372);
or U14484 (N_14484,N_14259,N_14273);
nand U14485 (N_14485,N_14375,N_14241);
and U14486 (N_14486,N_14327,N_14275);
nor U14487 (N_14487,N_14325,N_14389);
nand U14488 (N_14488,N_14342,N_14256);
and U14489 (N_14489,N_14327,N_14386);
nand U14490 (N_14490,N_14247,N_14304);
or U14491 (N_14491,N_14390,N_14255);
or U14492 (N_14492,N_14385,N_14342);
or U14493 (N_14493,N_14249,N_14316);
or U14494 (N_14494,N_14289,N_14270);
or U14495 (N_14495,N_14292,N_14323);
nand U14496 (N_14496,N_14293,N_14262);
and U14497 (N_14497,N_14398,N_14315);
or U14498 (N_14498,N_14358,N_14295);
and U14499 (N_14499,N_14387,N_14251);
or U14500 (N_14500,N_14386,N_14345);
nand U14501 (N_14501,N_14355,N_14378);
nor U14502 (N_14502,N_14324,N_14275);
and U14503 (N_14503,N_14294,N_14282);
xor U14504 (N_14504,N_14375,N_14351);
nor U14505 (N_14505,N_14253,N_14293);
or U14506 (N_14506,N_14261,N_14318);
and U14507 (N_14507,N_14348,N_14285);
nand U14508 (N_14508,N_14284,N_14289);
nor U14509 (N_14509,N_14310,N_14294);
nand U14510 (N_14510,N_14302,N_14342);
and U14511 (N_14511,N_14259,N_14377);
nor U14512 (N_14512,N_14266,N_14357);
xor U14513 (N_14513,N_14385,N_14269);
or U14514 (N_14514,N_14350,N_14362);
and U14515 (N_14515,N_14371,N_14335);
and U14516 (N_14516,N_14256,N_14250);
and U14517 (N_14517,N_14280,N_14387);
nand U14518 (N_14518,N_14271,N_14393);
nor U14519 (N_14519,N_14246,N_14308);
xnor U14520 (N_14520,N_14241,N_14291);
xnor U14521 (N_14521,N_14271,N_14336);
xnor U14522 (N_14522,N_14243,N_14353);
or U14523 (N_14523,N_14394,N_14357);
nand U14524 (N_14524,N_14393,N_14291);
xor U14525 (N_14525,N_14365,N_14265);
and U14526 (N_14526,N_14281,N_14357);
xnor U14527 (N_14527,N_14323,N_14344);
or U14528 (N_14528,N_14351,N_14354);
nor U14529 (N_14529,N_14248,N_14264);
and U14530 (N_14530,N_14363,N_14354);
nor U14531 (N_14531,N_14312,N_14381);
and U14532 (N_14532,N_14363,N_14289);
nand U14533 (N_14533,N_14371,N_14348);
and U14534 (N_14534,N_14303,N_14354);
and U14535 (N_14535,N_14260,N_14366);
nor U14536 (N_14536,N_14250,N_14280);
nand U14537 (N_14537,N_14304,N_14255);
xnor U14538 (N_14538,N_14248,N_14270);
nand U14539 (N_14539,N_14245,N_14244);
nand U14540 (N_14540,N_14377,N_14296);
and U14541 (N_14541,N_14335,N_14271);
or U14542 (N_14542,N_14251,N_14300);
or U14543 (N_14543,N_14359,N_14310);
nand U14544 (N_14544,N_14336,N_14313);
and U14545 (N_14545,N_14260,N_14343);
or U14546 (N_14546,N_14320,N_14311);
nand U14547 (N_14547,N_14329,N_14322);
nand U14548 (N_14548,N_14244,N_14314);
nand U14549 (N_14549,N_14365,N_14296);
or U14550 (N_14550,N_14271,N_14292);
and U14551 (N_14551,N_14340,N_14242);
xnor U14552 (N_14552,N_14276,N_14254);
xor U14553 (N_14553,N_14253,N_14332);
nor U14554 (N_14554,N_14304,N_14366);
and U14555 (N_14555,N_14250,N_14247);
and U14556 (N_14556,N_14399,N_14353);
nand U14557 (N_14557,N_14299,N_14391);
nor U14558 (N_14558,N_14292,N_14324);
or U14559 (N_14559,N_14262,N_14377);
nor U14560 (N_14560,N_14529,N_14459);
nor U14561 (N_14561,N_14407,N_14502);
and U14562 (N_14562,N_14498,N_14514);
nor U14563 (N_14563,N_14461,N_14518);
nor U14564 (N_14564,N_14460,N_14457);
or U14565 (N_14565,N_14527,N_14418);
xnor U14566 (N_14566,N_14417,N_14449);
and U14567 (N_14567,N_14405,N_14499);
nand U14568 (N_14568,N_14437,N_14462);
xor U14569 (N_14569,N_14517,N_14557);
or U14570 (N_14570,N_14494,N_14426);
nand U14571 (N_14571,N_14472,N_14447);
xnor U14572 (N_14572,N_14448,N_14487);
xnor U14573 (N_14573,N_14503,N_14428);
xnor U14574 (N_14574,N_14427,N_14535);
and U14575 (N_14575,N_14436,N_14492);
or U14576 (N_14576,N_14500,N_14477);
xor U14577 (N_14577,N_14455,N_14450);
xor U14578 (N_14578,N_14410,N_14516);
nor U14579 (N_14579,N_14542,N_14452);
nor U14580 (N_14580,N_14480,N_14486);
and U14581 (N_14581,N_14442,N_14401);
nor U14582 (N_14582,N_14440,N_14409);
xor U14583 (N_14583,N_14550,N_14530);
and U14584 (N_14584,N_14444,N_14478);
nor U14585 (N_14585,N_14541,N_14493);
nor U14586 (N_14586,N_14556,N_14469);
xor U14587 (N_14587,N_14470,N_14435);
or U14588 (N_14588,N_14504,N_14402);
and U14589 (N_14589,N_14429,N_14540);
and U14590 (N_14590,N_14484,N_14408);
xor U14591 (N_14591,N_14423,N_14475);
and U14592 (N_14592,N_14466,N_14422);
xor U14593 (N_14593,N_14554,N_14458);
or U14594 (N_14594,N_14505,N_14421);
or U14595 (N_14595,N_14445,N_14539);
nor U14596 (N_14596,N_14528,N_14456);
xor U14597 (N_14597,N_14548,N_14512);
nand U14598 (N_14598,N_14552,N_14439);
and U14599 (N_14599,N_14544,N_14549);
and U14600 (N_14600,N_14524,N_14431);
and U14601 (N_14601,N_14543,N_14559);
nand U14602 (N_14602,N_14522,N_14510);
and U14603 (N_14603,N_14525,N_14463);
nand U14604 (N_14604,N_14400,N_14515);
or U14605 (N_14605,N_14473,N_14558);
and U14606 (N_14606,N_14520,N_14467);
nand U14607 (N_14607,N_14419,N_14509);
xnor U14608 (N_14608,N_14438,N_14479);
or U14609 (N_14609,N_14415,N_14474);
and U14610 (N_14610,N_14416,N_14497);
nand U14611 (N_14611,N_14424,N_14521);
and U14612 (N_14612,N_14526,N_14523);
xnor U14613 (N_14613,N_14507,N_14489);
and U14614 (N_14614,N_14534,N_14545);
nand U14615 (N_14615,N_14425,N_14531);
nand U14616 (N_14616,N_14547,N_14481);
nand U14617 (N_14617,N_14404,N_14464);
xor U14618 (N_14618,N_14551,N_14485);
xnor U14619 (N_14619,N_14532,N_14533);
and U14620 (N_14620,N_14513,N_14508);
nand U14621 (N_14621,N_14412,N_14501);
xor U14622 (N_14622,N_14538,N_14451);
nor U14623 (N_14623,N_14496,N_14432);
nor U14624 (N_14624,N_14546,N_14491);
xor U14625 (N_14625,N_14420,N_14465);
and U14626 (N_14626,N_14483,N_14454);
xnor U14627 (N_14627,N_14490,N_14443);
xnor U14628 (N_14628,N_14482,N_14471);
and U14629 (N_14629,N_14511,N_14488);
nor U14630 (N_14630,N_14446,N_14476);
nor U14631 (N_14631,N_14519,N_14553);
and U14632 (N_14632,N_14506,N_14495);
or U14633 (N_14633,N_14414,N_14441);
xnor U14634 (N_14634,N_14468,N_14406);
and U14635 (N_14635,N_14430,N_14555);
nor U14636 (N_14636,N_14536,N_14413);
and U14637 (N_14637,N_14403,N_14537);
xnor U14638 (N_14638,N_14434,N_14453);
nand U14639 (N_14639,N_14411,N_14433);
nand U14640 (N_14640,N_14540,N_14490);
xnor U14641 (N_14641,N_14512,N_14524);
nor U14642 (N_14642,N_14478,N_14447);
and U14643 (N_14643,N_14501,N_14451);
xnor U14644 (N_14644,N_14508,N_14491);
nor U14645 (N_14645,N_14446,N_14530);
nand U14646 (N_14646,N_14453,N_14525);
xor U14647 (N_14647,N_14554,N_14528);
nor U14648 (N_14648,N_14522,N_14503);
xor U14649 (N_14649,N_14523,N_14559);
xor U14650 (N_14650,N_14490,N_14499);
xor U14651 (N_14651,N_14528,N_14534);
or U14652 (N_14652,N_14402,N_14545);
nand U14653 (N_14653,N_14532,N_14467);
nand U14654 (N_14654,N_14498,N_14508);
or U14655 (N_14655,N_14532,N_14404);
and U14656 (N_14656,N_14514,N_14500);
and U14657 (N_14657,N_14527,N_14432);
and U14658 (N_14658,N_14423,N_14400);
nor U14659 (N_14659,N_14442,N_14446);
nor U14660 (N_14660,N_14402,N_14469);
or U14661 (N_14661,N_14476,N_14440);
nand U14662 (N_14662,N_14436,N_14524);
xor U14663 (N_14663,N_14533,N_14488);
nor U14664 (N_14664,N_14520,N_14473);
nand U14665 (N_14665,N_14554,N_14500);
xor U14666 (N_14666,N_14558,N_14413);
nor U14667 (N_14667,N_14514,N_14488);
nor U14668 (N_14668,N_14411,N_14443);
xnor U14669 (N_14669,N_14485,N_14507);
or U14670 (N_14670,N_14498,N_14525);
xnor U14671 (N_14671,N_14453,N_14489);
xnor U14672 (N_14672,N_14501,N_14459);
nand U14673 (N_14673,N_14479,N_14415);
and U14674 (N_14674,N_14557,N_14453);
nor U14675 (N_14675,N_14551,N_14490);
nor U14676 (N_14676,N_14546,N_14427);
nor U14677 (N_14677,N_14426,N_14446);
nor U14678 (N_14678,N_14471,N_14506);
or U14679 (N_14679,N_14471,N_14450);
nor U14680 (N_14680,N_14509,N_14539);
or U14681 (N_14681,N_14502,N_14462);
nor U14682 (N_14682,N_14510,N_14521);
nor U14683 (N_14683,N_14457,N_14470);
and U14684 (N_14684,N_14431,N_14404);
and U14685 (N_14685,N_14403,N_14463);
xnor U14686 (N_14686,N_14434,N_14522);
or U14687 (N_14687,N_14522,N_14527);
xnor U14688 (N_14688,N_14448,N_14547);
xor U14689 (N_14689,N_14540,N_14477);
nand U14690 (N_14690,N_14437,N_14482);
xnor U14691 (N_14691,N_14412,N_14465);
nor U14692 (N_14692,N_14438,N_14537);
nor U14693 (N_14693,N_14498,N_14430);
xor U14694 (N_14694,N_14468,N_14538);
and U14695 (N_14695,N_14491,N_14476);
or U14696 (N_14696,N_14436,N_14488);
nor U14697 (N_14697,N_14511,N_14478);
or U14698 (N_14698,N_14520,N_14416);
nand U14699 (N_14699,N_14420,N_14442);
nor U14700 (N_14700,N_14549,N_14501);
and U14701 (N_14701,N_14511,N_14498);
and U14702 (N_14702,N_14492,N_14502);
nand U14703 (N_14703,N_14493,N_14424);
or U14704 (N_14704,N_14500,N_14540);
nor U14705 (N_14705,N_14465,N_14523);
nor U14706 (N_14706,N_14549,N_14499);
nand U14707 (N_14707,N_14480,N_14461);
xor U14708 (N_14708,N_14463,N_14544);
nand U14709 (N_14709,N_14552,N_14504);
nand U14710 (N_14710,N_14413,N_14500);
nand U14711 (N_14711,N_14449,N_14516);
xnor U14712 (N_14712,N_14525,N_14417);
and U14713 (N_14713,N_14534,N_14506);
xor U14714 (N_14714,N_14508,N_14489);
and U14715 (N_14715,N_14460,N_14417);
nand U14716 (N_14716,N_14524,N_14517);
nand U14717 (N_14717,N_14430,N_14428);
nor U14718 (N_14718,N_14451,N_14470);
nor U14719 (N_14719,N_14504,N_14529);
or U14720 (N_14720,N_14677,N_14637);
or U14721 (N_14721,N_14578,N_14670);
and U14722 (N_14722,N_14579,N_14656);
or U14723 (N_14723,N_14696,N_14594);
and U14724 (N_14724,N_14702,N_14633);
nor U14725 (N_14725,N_14713,N_14629);
and U14726 (N_14726,N_14708,N_14662);
or U14727 (N_14727,N_14631,N_14614);
nand U14728 (N_14728,N_14603,N_14680);
and U14729 (N_14729,N_14621,N_14672);
nand U14730 (N_14730,N_14688,N_14666);
nand U14731 (N_14731,N_14609,N_14620);
nor U14732 (N_14732,N_14652,N_14564);
nor U14733 (N_14733,N_14706,N_14712);
xor U14734 (N_14734,N_14560,N_14563);
xnor U14735 (N_14735,N_14583,N_14582);
nand U14736 (N_14736,N_14659,N_14570);
nor U14737 (N_14737,N_14705,N_14585);
or U14738 (N_14738,N_14684,N_14587);
xnor U14739 (N_14739,N_14648,N_14719);
xor U14740 (N_14740,N_14709,N_14695);
nor U14741 (N_14741,N_14678,N_14591);
xor U14742 (N_14742,N_14622,N_14600);
and U14743 (N_14743,N_14632,N_14580);
nor U14744 (N_14744,N_14668,N_14685);
nor U14745 (N_14745,N_14601,N_14572);
and U14746 (N_14746,N_14718,N_14595);
xnor U14747 (N_14747,N_14616,N_14665);
and U14748 (N_14748,N_14676,N_14635);
nand U14749 (N_14749,N_14649,N_14667);
or U14750 (N_14750,N_14574,N_14625);
or U14751 (N_14751,N_14673,N_14598);
or U14752 (N_14752,N_14651,N_14716);
xor U14753 (N_14753,N_14576,N_14711);
and U14754 (N_14754,N_14645,N_14671);
xor U14755 (N_14755,N_14565,N_14599);
xor U14756 (N_14756,N_14630,N_14592);
nand U14757 (N_14757,N_14715,N_14717);
nand U14758 (N_14758,N_14681,N_14596);
nand U14759 (N_14759,N_14571,N_14569);
or U14760 (N_14760,N_14704,N_14638);
and U14761 (N_14761,N_14693,N_14661);
nand U14762 (N_14762,N_14607,N_14611);
nor U14763 (N_14763,N_14605,N_14590);
xor U14764 (N_14764,N_14664,N_14608);
and U14765 (N_14765,N_14692,N_14644);
or U14766 (N_14766,N_14698,N_14627);
xor U14767 (N_14767,N_14634,N_14646);
xnor U14768 (N_14768,N_14683,N_14628);
nand U14769 (N_14769,N_14640,N_14617);
xor U14770 (N_14770,N_14624,N_14636);
and U14771 (N_14771,N_14669,N_14675);
nand U14772 (N_14772,N_14689,N_14674);
nand U14773 (N_14773,N_14690,N_14568);
or U14774 (N_14774,N_14562,N_14618);
or U14775 (N_14775,N_14697,N_14682);
nand U14776 (N_14776,N_14650,N_14679);
nor U14777 (N_14777,N_14575,N_14660);
nor U14778 (N_14778,N_14707,N_14639);
nand U14779 (N_14779,N_14703,N_14657);
xor U14780 (N_14780,N_14602,N_14663);
nand U14781 (N_14781,N_14584,N_14710);
nand U14782 (N_14782,N_14647,N_14588);
and U14783 (N_14783,N_14573,N_14714);
and U14784 (N_14784,N_14593,N_14655);
xor U14785 (N_14785,N_14643,N_14658);
nand U14786 (N_14786,N_14619,N_14701);
and U14787 (N_14787,N_14586,N_14561);
xnor U14788 (N_14788,N_14626,N_14641);
nor U14789 (N_14789,N_14694,N_14699);
or U14790 (N_14790,N_14612,N_14581);
nand U14791 (N_14791,N_14604,N_14691);
and U14792 (N_14792,N_14653,N_14577);
nor U14793 (N_14793,N_14615,N_14597);
and U14794 (N_14794,N_14589,N_14623);
nor U14795 (N_14795,N_14613,N_14567);
nor U14796 (N_14796,N_14700,N_14606);
nor U14797 (N_14797,N_14566,N_14687);
nand U14798 (N_14798,N_14686,N_14642);
xor U14799 (N_14799,N_14610,N_14654);
xor U14800 (N_14800,N_14710,N_14685);
or U14801 (N_14801,N_14586,N_14592);
and U14802 (N_14802,N_14620,N_14644);
nor U14803 (N_14803,N_14593,N_14705);
xnor U14804 (N_14804,N_14572,N_14644);
nor U14805 (N_14805,N_14699,N_14653);
or U14806 (N_14806,N_14690,N_14709);
and U14807 (N_14807,N_14575,N_14701);
nand U14808 (N_14808,N_14663,N_14697);
xnor U14809 (N_14809,N_14693,N_14692);
xnor U14810 (N_14810,N_14685,N_14599);
xor U14811 (N_14811,N_14717,N_14573);
or U14812 (N_14812,N_14639,N_14640);
and U14813 (N_14813,N_14695,N_14600);
or U14814 (N_14814,N_14629,N_14700);
or U14815 (N_14815,N_14632,N_14577);
nor U14816 (N_14816,N_14641,N_14623);
and U14817 (N_14817,N_14711,N_14696);
nor U14818 (N_14818,N_14564,N_14617);
nor U14819 (N_14819,N_14709,N_14641);
or U14820 (N_14820,N_14601,N_14669);
and U14821 (N_14821,N_14699,N_14669);
xor U14822 (N_14822,N_14561,N_14591);
or U14823 (N_14823,N_14577,N_14652);
nor U14824 (N_14824,N_14689,N_14592);
and U14825 (N_14825,N_14575,N_14667);
xnor U14826 (N_14826,N_14710,N_14663);
nor U14827 (N_14827,N_14636,N_14686);
or U14828 (N_14828,N_14711,N_14668);
and U14829 (N_14829,N_14610,N_14715);
nand U14830 (N_14830,N_14662,N_14680);
nand U14831 (N_14831,N_14585,N_14714);
and U14832 (N_14832,N_14672,N_14680);
nand U14833 (N_14833,N_14651,N_14624);
nor U14834 (N_14834,N_14669,N_14562);
xnor U14835 (N_14835,N_14685,N_14701);
or U14836 (N_14836,N_14590,N_14699);
or U14837 (N_14837,N_14564,N_14647);
and U14838 (N_14838,N_14621,N_14587);
nor U14839 (N_14839,N_14566,N_14709);
nor U14840 (N_14840,N_14607,N_14588);
xnor U14841 (N_14841,N_14601,N_14570);
xor U14842 (N_14842,N_14699,N_14618);
nor U14843 (N_14843,N_14622,N_14714);
or U14844 (N_14844,N_14641,N_14592);
xnor U14845 (N_14845,N_14582,N_14692);
xnor U14846 (N_14846,N_14577,N_14633);
nand U14847 (N_14847,N_14575,N_14685);
nand U14848 (N_14848,N_14647,N_14680);
nor U14849 (N_14849,N_14701,N_14668);
nor U14850 (N_14850,N_14603,N_14692);
or U14851 (N_14851,N_14663,N_14695);
xnor U14852 (N_14852,N_14691,N_14624);
nand U14853 (N_14853,N_14611,N_14670);
and U14854 (N_14854,N_14606,N_14692);
nor U14855 (N_14855,N_14686,N_14568);
or U14856 (N_14856,N_14629,N_14643);
nand U14857 (N_14857,N_14572,N_14608);
nand U14858 (N_14858,N_14676,N_14707);
nand U14859 (N_14859,N_14665,N_14562);
nor U14860 (N_14860,N_14673,N_14592);
xnor U14861 (N_14861,N_14641,N_14697);
nor U14862 (N_14862,N_14677,N_14664);
xor U14863 (N_14863,N_14709,N_14631);
xnor U14864 (N_14864,N_14706,N_14679);
nand U14865 (N_14865,N_14571,N_14585);
nand U14866 (N_14866,N_14599,N_14562);
xor U14867 (N_14867,N_14654,N_14566);
xnor U14868 (N_14868,N_14647,N_14571);
or U14869 (N_14869,N_14584,N_14701);
or U14870 (N_14870,N_14696,N_14624);
nand U14871 (N_14871,N_14704,N_14623);
nor U14872 (N_14872,N_14684,N_14601);
xnor U14873 (N_14873,N_14625,N_14627);
nand U14874 (N_14874,N_14565,N_14619);
or U14875 (N_14875,N_14661,N_14598);
and U14876 (N_14876,N_14634,N_14672);
xnor U14877 (N_14877,N_14676,N_14607);
nand U14878 (N_14878,N_14632,N_14635);
nor U14879 (N_14879,N_14712,N_14649);
and U14880 (N_14880,N_14763,N_14805);
or U14881 (N_14881,N_14829,N_14789);
and U14882 (N_14882,N_14826,N_14794);
nand U14883 (N_14883,N_14803,N_14855);
nand U14884 (N_14884,N_14834,N_14837);
or U14885 (N_14885,N_14864,N_14857);
xor U14886 (N_14886,N_14869,N_14754);
xnor U14887 (N_14887,N_14727,N_14755);
or U14888 (N_14888,N_14799,N_14844);
nand U14889 (N_14889,N_14796,N_14868);
or U14890 (N_14890,N_14753,N_14740);
xor U14891 (N_14891,N_14737,N_14744);
and U14892 (N_14892,N_14780,N_14759);
nor U14893 (N_14893,N_14845,N_14800);
xor U14894 (N_14894,N_14752,N_14827);
xnor U14895 (N_14895,N_14768,N_14771);
nor U14896 (N_14896,N_14860,N_14876);
and U14897 (N_14897,N_14874,N_14774);
nand U14898 (N_14898,N_14784,N_14720);
or U14899 (N_14899,N_14721,N_14854);
nand U14900 (N_14900,N_14871,N_14732);
nor U14901 (N_14901,N_14866,N_14824);
or U14902 (N_14902,N_14728,N_14762);
or U14903 (N_14903,N_14861,N_14867);
and U14904 (N_14904,N_14828,N_14757);
and U14905 (N_14905,N_14722,N_14779);
nand U14906 (N_14906,N_14830,N_14764);
and U14907 (N_14907,N_14726,N_14733);
nor U14908 (N_14908,N_14736,N_14749);
xor U14909 (N_14909,N_14817,N_14804);
xor U14910 (N_14910,N_14751,N_14831);
xnor U14911 (N_14911,N_14730,N_14782);
or U14912 (N_14912,N_14807,N_14731);
and U14913 (N_14913,N_14767,N_14842);
nor U14914 (N_14914,N_14858,N_14760);
or U14915 (N_14915,N_14843,N_14734);
xnor U14916 (N_14916,N_14738,N_14814);
nand U14917 (N_14917,N_14798,N_14849);
nor U14918 (N_14918,N_14788,N_14847);
and U14919 (N_14919,N_14851,N_14853);
nor U14920 (N_14920,N_14793,N_14818);
nand U14921 (N_14921,N_14781,N_14790);
xnor U14922 (N_14922,N_14823,N_14766);
nor U14923 (N_14923,N_14802,N_14839);
nand U14924 (N_14924,N_14777,N_14838);
xnor U14925 (N_14925,N_14840,N_14819);
and U14926 (N_14926,N_14747,N_14835);
nor U14927 (N_14927,N_14748,N_14787);
and U14928 (N_14928,N_14863,N_14832);
and U14929 (N_14929,N_14765,N_14813);
or U14930 (N_14930,N_14769,N_14870);
nand U14931 (N_14931,N_14877,N_14775);
or U14932 (N_14932,N_14850,N_14820);
and U14933 (N_14933,N_14723,N_14862);
nor U14934 (N_14934,N_14822,N_14746);
or U14935 (N_14935,N_14772,N_14741);
or U14936 (N_14936,N_14758,N_14773);
nand U14937 (N_14937,N_14852,N_14735);
nor U14938 (N_14938,N_14873,N_14865);
nor U14939 (N_14939,N_14801,N_14739);
nand U14940 (N_14940,N_14795,N_14770);
or U14941 (N_14941,N_14725,N_14778);
nand U14942 (N_14942,N_14812,N_14756);
xor U14943 (N_14943,N_14841,N_14761);
or U14944 (N_14944,N_14836,N_14785);
nand U14945 (N_14945,N_14811,N_14729);
nand U14946 (N_14946,N_14859,N_14809);
nor U14947 (N_14947,N_14872,N_14745);
and U14948 (N_14948,N_14848,N_14816);
nand U14949 (N_14949,N_14797,N_14724);
and U14950 (N_14950,N_14846,N_14792);
and U14951 (N_14951,N_14833,N_14776);
xnor U14952 (N_14952,N_14821,N_14878);
xnor U14953 (N_14953,N_14808,N_14810);
or U14954 (N_14954,N_14815,N_14791);
nand U14955 (N_14955,N_14750,N_14825);
and U14956 (N_14956,N_14786,N_14743);
nand U14957 (N_14957,N_14806,N_14783);
and U14958 (N_14958,N_14742,N_14856);
nor U14959 (N_14959,N_14879,N_14875);
or U14960 (N_14960,N_14826,N_14820);
nand U14961 (N_14961,N_14759,N_14816);
or U14962 (N_14962,N_14860,N_14817);
nand U14963 (N_14963,N_14834,N_14838);
and U14964 (N_14964,N_14864,N_14836);
nor U14965 (N_14965,N_14745,N_14803);
nand U14966 (N_14966,N_14849,N_14842);
xor U14967 (N_14967,N_14845,N_14746);
and U14968 (N_14968,N_14777,N_14875);
nand U14969 (N_14969,N_14785,N_14763);
or U14970 (N_14970,N_14776,N_14768);
nor U14971 (N_14971,N_14852,N_14745);
nor U14972 (N_14972,N_14814,N_14740);
nand U14973 (N_14973,N_14811,N_14777);
nor U14974 (N_14974,N_14783,N_14836);
xnor U14975 (N_14975,N_14870,N_14831);
xnor U14976 (N_14976,N_14838,N_14865);
or U14977 (N_14977,N_14793,N_14822);
xor U14978 (N_14978,N_14723,N_14787);
nand U14979 (N_14979,N_14748,N_14759);
or U14980 (N_14980,N_14755,N_14772);
xnor U14981 (N_14981,N_14820,N_14723);
or U14982 (N_14982,N_14790,N_14789);
or U14983 (N_14983,N_14829,N_14830);
and U14984 (N_14984,N_14765,N_14740);
or U14985 (N_14985,N_14779,N_14740);
and U14986 (N_14986,N_14781,N_14724);
nor U14987 (N_14987,N_14811,N_14838);
and U14988 (N_14988,N_14760,N_14872);
or U14989 (N_14989,N_14729,N_14766);
nor U14990 (N_14990,N_14737,N_14796);
or U14991 (N_14991,N_14814,N_14746);
nor U14992 (N_14992,N_14739,N_14779);
and U14993 (N_14993,N_14744,N_14805);
xnor U14994 (N_14994,N_14756,N_14768);
xnor U14995 (N_14995,N_14846,N_14823);
xor U14996 (N_14996,N_14846,N_14857);
and U14997 (N_14997,N_14728,N_14849);
or U14998 (N_14998,N_14824,N_14726);
xnor U14999 (N_14999,N_14806,N_14727);
xnor U15000 (N_15000,N_14780,N_14817);
or U15001 (N_15001,N_14836,N_14777);
nand U15002 (N_15002,N_14735,N_14790);
xnor U15003 (N_15003,N_14741,N_14742);
xnor U15004 (N_15004,N_14726,N_14758);
nand U15005 (N_15005,N_14758,N_14840);
xnor U15006 (N_15006,N_14844,N_14851);
or U15007 (N_15007,N_14830,N_14796);
nand U15008 (N_15008,N_14748,N_14809);
nand U15009 (N_15009,N_14742,N_14803);
nor U15010 (N_15010,N_14730,N_14741);
or U15011 (N_15011,N_14755,N_14833);
or U15012 (N_15012,N_14807,N_14814);
or U15013 (N_15013,N_14758,N_14808);
and U15014 (N_15014,N_14755,N_14824);
or U15015 (N_15015,N_14720,N_14850);
nand U15016 (N_15016,N_14874,N_14769);
nand U15017 (N_15017,N_14741,N_14745);
nor U15018 (N_15018,N_14765,N_14847);
nand U15019 (N_15019,N_14751,N_14800);
nor U15020 (N_15020,N_14767,N_14866);
nor U15021 (N_15021,N_14858,N_14728);
nand U15022 (N_15022,N_14734,N_14873);
and U15023 (N_15023,N_14847,N_14778);
nor U15024 (N_15024,N_14821,N_14783);
nor U15025 (N_15025,N_14828,N_14791);
xor U15026 (N_15026,N_14741,N_14720);
nand U15027 (N_15027,N_14779,N_14760);
nor U15028 (N_15028,N_14729,N_14860);
xor U15029 (N_15029,N_14824,N_14781);
and U15030 (N_15030,N_14752,N_14744);
nor U15031 (N_15031,N_14736,N_14846);
or U15032 (N_15032,N_14851,N_14796);
xor U15033 (N_15033,N_14850,N_14877);
nand U15034 (N_15034,N_14863,N_14802);
nand U15035 (N_15035,N_14775,N_14821);
nand U15036 (N_15036,N_14746,N_14823);
nor U15037 (N_15037,N_14862,N_14800);
or U15038 (N_15038,N_14720,N_14753);
nand U15039 (N_15039,N_14783,N_14780);
or U15040 (N_15040,N_15004,N_14984);
or U15041 (N_15041,N_14905,N_14906);
nor U15042 (N_15042,N_14925,N_14941);
nor U15043 (N_15043,N_14917,N_14896);
or U15044 (N_15044,N_15003,N_14952);
nand U15045 (N_15045,N_14933,N_15034);
xnor U15046 (N_15046,N_14926,N_14914);
or U15047 (N_15047,N_15006,N_14924);
and U15048 (N_15048,N_14948,N_14950);
or U15049 (N_15049,N_14974,N_14956);
xor U15050 (N_15050,N_15021,N_14992);
or U15051 (N_15051,N_14910,N_14985);
nor U15052 (N_15052,N_15007,N_14929);
or U15053 (N_15053,N_14889,N_14978);
nand U15054 (N_15054,N_14886,N_14884);
nand U15055 (N_15055,N_14949,N_14893);
or U15056 (N_15056,N_14918,N_14951);
and U15057 (N_15057,N_14895,N_14981);
or U15058 (N_15058,N_15001,N_14988);
and U15059 (N_15059,N_15017,N_15028);
nor U15060 (N_15060,N_14913,N_14971);
and U15061 (N_15061,N_14943,N_14937);
and U15062 (N_15062,N_14919,N_15036);
nand U15063 (N_15063,N_15005,N_14973);
nand U15064 (N_15064,N_15010,N_14885);
and U15065 (N_15065,N_14955,N_15011);
xnor U15066 (N_15066,N_14947,N_14923);
or U15067 (N_15067,N_14944,N_14907);
or U15068 (N_15068,N_15025,N_14890);
nand U15069 (N_15069,N_14922,N_14983);
or U15070 (N_15070,N_14994,N_15023);
nand U15071 (N_15071,N_14960,N_14880);
nor U15072 (N_15072,N_14927,N_14934);
xor U15073 (N_15073,N_15027,N_15009);
nand U15074 (N_15074,N_14892,N_14883);
xnor U15075 (N_15075,N_14882,N_14945);
nand U15076 (N_15076,N_14997,N_14969);
nand U15077 (N_15077,N_14964,N_15039);
nand U15078 (N_15078,N_14920,N_14921);
nand U15079 (N_15079,N_14976,N_15019);
xor U15080 (N_15080,N_14987,N_14891);
nand U15081 (N_15081,N_14972,N_14959);
and U15082 (N_15082,N_15012,N_14935);
nor U15083 (N_15083,N_14939,N_14912);
and U15084 (N_15084,N_14931,N_15002);
xor U15085 (N_15085,N_14961,N_15022);
or U15086 (N_15086,N_14909,N_14979);
nor U15087 (N_15087,N_15015,N_14901);
nand U15088 (N_15088,N_15035,N_14908);
xor U15089 (N_15089,N_14990,N_14902);
nor U15090 (N_15090,N_14928,N_14881);
and U15091 (N_15091,N_15000,N_14965);
nand U15092 (N_15092,N_14903,N_15029);
nor U15093 (N_15093,N_14887,N_14970);
nor U15094 (N_15094,N_15013,N_15024);
nor U15095 (N_15095,N_14975,N_14989);
nand U15096 (N_15096,N_14898,N_14993);
xor U15097 (N_15097,N_14932,N_14958);
nand U15098 (N_15098,N_15033,N_15026);
and U15099 (N_15099,N_14998,N_14897);
and U15100 (N_15100,N_14904,N_14940);
nand U15101 (N_15101,N_14915,N_14991);
nor U15102 (N_15102,N_14946,N_14966);
and U15103 (N_15103,N_14888,N_14938);
nor U15104 (N_15104,N_15030,N_14963);
nand U15105 (N_15105,N_14954,N_14995);
nand U15106 (N_15106,N_14957,N_14894);
nand U15107 (N_15107,N_15031,N_14996);
or U15108 (N_15108,N_14900,N_15016);
or U15109 (N_15109,N_14967,N_15008);
nand U15110 (N_15110,N_14936,N_14977);
nand U15111 (N_15111,N_14899,N_15014);
or U15112 (N_15112,N_15032,N_14916);
xnor U15113 (N_15113,N_14968,N_14962);
xnor U15114 (N_15114,N_15018,N_15020);
xor U15115 (N_15115,N_14982,N_14953);
xor U15116 (N_15116,N_15038,N_14911);
nor U15117 (N_15117,N_14999,N_14986);
and U15118 (N_15118,N_14942,N_15037);
xor U15119 (N_15119,N_14930,N_14980);
nand U15120 (N_15120,N_14901,N_14906);
nor U15121 (N_15121,N_14957,N_14991);
xor U15122 (N_15122,N_14992,N_14887);
or U15123 (N_15123,N_14996,N_15000);
nor U15124 (N_15124,N_14918,N_14884);
and U15125 (N_15125,N_14944,N_14926);
nand U15126 (N_15126,N_15026,N_15038);
or U15127 (N_15127,N_15002,N_14887);
xor U15128 (N_15128,N_14991,N_14950);
or U15129 (N_15129,N_14929,N_14979);
nand U15130 (N_15130,N_14912,N_14971);
nand U15131 (N_15131,N_15009,N_15000);
nand U15132 (N_15132,N_14950,N_15027);
and U15133 (N_15133,N_15039,N_14962);
nand U15134 (N_15134,N_14907,N_14922);
nor U15135 (N_15135,N_15000,N_14915);
xor U15136 (N_15136,N_14891,N_15005);
or U15137 (N_15137,N_14928,N_14924);
nand U15138 (N_15138,N_14952,N_15004);
xor U15139 (N_15139,N_14951,N_14890);
nor U15140 (N_15140,N_14974,N_14964);
or U15141 (N_15141,N_14931,N_14903);
nor U15142 (N_15142,N_15030,N_15035);
and U15143 (N_15143,N_14970,N_14929);
nor U15144 (N_15144,N_15005,N_15033);
xnor U15145 (N_15145,N_14883,N_14880);
nor U15146 (N_15146,N_14904,N_14942);
nand U15147 (N_15147,N_14943,N_14985);
and U15148 (N_15148,N_14882,N_15026);
xnor U15149 (N_15149,N_14903,N_14988);
and U15150 (N_15150,N_14928,N_14985);
or U15151 (N_15151,N_14977,N_14939);
xnor U15152 (N_15152,N_15028,N_14890);
nor U15153 (N_15153,N_15034,N_14993);
xnor U15154 (N_15154,N_15013,N_14995);
nor U15155 (N_15155,N_15031,N_15000);
nor U15156 (N_15156,N_14971,N_15035);
nor U15157 (N_15157,N_14908,N_14950);
or U15158 (N_15158,N_14966,N_14956);
nor U15159 (N_15159,N_14948,N_14912);
nor U15160 (N_15160,N_14956,N_15035);
nor U15161 (N_15161,N_14901,N_14909);
and U15162 (N_15162,N_14988,N_14993);
and U15163 (N_15163,N_14929,N_14881);
nor U15164 (N_15164,N_14981,N_14947);
nand U15165 (N_15165,N_14899,N_15029);
and U15166 (N_15166,N_15003,N_14972);
and U15167 (N_15167,N_14942,N_15021);
nor U15168 (N_15168,N_14899,N_15000);
and U15169 (N_15169,N_15026,N_14916);
nand U15170 (N_15170,N_14916,N_14952);
nand U15171 (N_15171,N_14955,N_14899);
or U15172 (N_15172,N_14888,N_14989);
or U15173 (N_15173,N_14905,N_14969);
and U15174 (N_15174,N_14970,N_14972);
or U15175 (N_15175,N_14961,N_15002);
nand U15176 (N_15176,N_14935,N_14895);
nand U15177 (N_15177,N_15011,N_14881);
xnor U15178 (N_15178,N_14954,N_14949);
nand U15179 (N_15179,N_15025,N_14962);
and U15180 (N_15180,N_15035,N_14924);
nor U15181 (N_15181,N_15020,N_14921);
nor U15182 (N_15182,N_14910,N_15033);
or U15183 (N_15183,N_15003,N_14979);
nor U15184 (N_15184,N_14933,N_14898);
or U15185 (N_15185,N_14931,N_15008);
and U15186 (N_15186,N_15016,N_15030);
nand U15187 (N_15187,N_15024,N_14920);
xnor U15188 (N_15188,N_14962,N_14977);
xnor U15189 (N_15189,N_14884,N_15033);
nor U15190 (N_15190,N_14960,N_14975);
and U15191 (N_15191,N_14904,N_14970);
xnor U15192 (N_15192,N_14957,N_14928);
or U15193 (N_15193,N_14946,N_14900);
or U15194 (N_15194,N_14968,N_14922);
xor U15195 (N_15195,N_14911,N_14902);
or U15196 (N_15196,N_14964,N_15023);
nor U15197 (N_15197,N_14987,N_15021);
nor U15198 (N_15198,N_14971,N_15002);
or U15199 (N_15199,N_14893,N_14956);
and U15200 (N_15200,N_15108,N_15101);
xnor U15201 (N_15201,N_15137,N_15193);
and U15202 (N_15202,N_15078,N_15094);
xor U15203 (N_15203,N_15114,N_15080);
or U15204 (N_15204,N_15163,N_15084);
or U15205 (N_15205,N_15073,N_15115);
nand U15206 (N_15206,N_15076,N_15070);
xnor U15207 (N_15207,N_15119,N_15168);
xnor U15208 (N_15208,N_15198,N_15058);
xor U15209 (N_15209,N_15071,N_15194);
and U15210 (N_15210,N_15199,N_15162);
xnor U15211 (N_15211,N_15068,N_15152);
xor U15212 (N_15212,N_15130,N_15116);
or U15213 (N_15213,N_15097,N_15063);
nand U15214 (N_15214,N_15179,N_15135);
or U15215 (N_15215,N_15173,N_15069);
or U15216 (N_15216,N_15079,N_15176);
and U15217 (N_15217,N_15118,N_15147);
and U15218 (N_15218,N_15178,N_15050);
nor U15219 (N_15219,N_15157,N_15124);
nand U15220 (N_15220,N_15110,N_15134);
xor U15221 (N_15221,N_15132,N_15169);
or U15222 (N_15222,N_15172,N_15160);
nand U15223 (N_15223,N_15123,N_15190);
xnor U15224 (N_15224,N_15133,N_15067);
or U15225 (N_15225,N_15103,N_15089);
nand U15226 (N_15226,N_15049,N_15040);
nand U15227 (N_15227,N_15141,N_15158);
nand U15228 (N_15228,N_15117,N_15091);
and U15229 (N_15229,N_15100,N_15072);
xor U15230 (N_15230,N_15183,N_15060);
nor U15231 (N_15231,N_15161,N_15047);
nand U15232 (N_15232,N_15112,N_15131);
nand U15233 (N_15233,N_15197,N_15142);
or U15234 (N_15234,N_15092,N_15095);
and U15235 (N_15235,N_15059,N_15155);
xnor U15236 (N_15236,N_15064,N_15081);
or U15237 (N_15237,N_15177,N_15104);
or U15238 (N_15238,N_15188,N_15143);
xor U15239 (N_15239,N_15164,N_15139);
or U15240 (N_15240,N_15166,N_15189);
or U15241 (N_15241,N_15061,N_15150);
or U15242 (N_15242,N_15086,N_15044);
nor U15243 (N_15243,N_15151,N_15106);
and U15244 (N_15244,N_15185,N_15056);
and U15245 (N_15245,N_15136,N_15159);
xor U15246 (N_15246,N_15170,N_15125);
nand U15247 (N_15247,N_15083,N_15066);
and U15248 (N_15248,N_15180,N_15140);
xnor U15249 (N_15249,N_15075,N_15145);
xnor U15250 (N_15250,N_15154,N_15065);
or U15251 (N_15251,N_15105,N_15156);
nand U15252 (N_15252,N_15053,N_15127);
or U15253 (N_15253,N_15088,N_15082);
nand U15254 (N_15254,N_15121,N_15111);
nor U15255 (N_15255,N_15098,N_15195);
nand U15256 (N_15256,N_15144,N_15042);
and U15257 (N_15257,N_15165,N_15077);
or U15258 (N_15258,N_15122,N_15052);
xor U15259 (N_15259,N_15149,N_15138);
and U15260 (N_15260,N_15062,N_15057);
or U15261 (N_15261,N_15174,N_15181);
xnor U15262 (N_15262,N_15041,N_15120);
nor U15263 (N_15263,N_15107,N_15129);
xor U15264 (N_15264,N_15074,N_15045);
or U15265 (N_15265,N_15146,N_15184);
nor U15266 (N_15266,N_15090,N_15055);
nand U15267 (N_15267,N_15093,N_15191);
or U15268 (N_15268,N_15099,N_15153);
nor U15269 (N_15269,N_15051,N_15182);
or U15270 (N_15270,N_15109,N_15187);
nand U15271 (N_15271,N_15167,N_15192);
and U15272 (N_15272,N_15113,N_15054);
nor U15273 (N_15273,N_15085,N_15048);
nor U15274 (N_15274,N_15186,N_15171);
and U15275 (N_15275,N_15043,N_15096);
xor U15276 (N_15276,N_15175,N_15148);
nand U15277 (N_15277,N_15087,N_15128);
or U15278 (N_15278,N_15102,N_15126);
xor U15279 (N_15279,N_15196,N_15046);
or U15280 (N_15280,N_15152,N_15050);
nand U15281 (N_15281,N_15186,N_15185);
nand U15282 (N_15282,N_15127,N_15152);
nor U15283 (N_15283,N_15091,N_15095);
nor U15284 (N_15284,N_15093,N_15188);
xnor U15285 (N_15285,N_15131,N_15071);
nand U15286 (N_15286,N_15090,N_15169);
or U15287 (N_15287,N_15078,N_15064);
nor U15288 (N_15288,N_15169,N_15156);
or U15289 (N_15289,N_15123,N_15199);
or U15290 (N_15290,N_15190,N_15163);
and U15291 (N_15291,N_15075,N_15148);
nand U15292 (N_15292,N_15132,N_15120);
xor U15293 (N_15293,N_15091,N_15191);
xor U15294 (N_15294,N_15126,N_15121);
nor U15295 (N_15295,N_15183,N_15172);
nand U15296 (N_15296,N_15046,N_15143);
xnor U15297 (N_15297,N_15183,N_15133);
or U15298 (N_15298,N_15120,N_15115);
or U15299 (N_15299,N_15180,N_15183);
and U15300 (N_15300,N_15126,N_15127);
xnor U15301 (N_15301,N_15116,N_15101);
or U15302 (N_15302,N_15124,N_15096);
nand U15303 (N_15303,N_15191,N_15140);
nor U15304 (N_15304,N_15093,N_15129);
nor U15305 (N_15305,N_15132,N_15187);
or U15306 (N_15306,N_15066,N_15154);
xor U15307 (N_15307,N_15151,N_15108);
nor U15308 (N_15308,N_15186,N_15135);
nor U15309 (N_15309,N_15185,N_15182);
or U15310 (N_15310,N_15066,N_15098);
nand U15311 (N_15311,N_15051,N_15090);
and U15312 (N_15312,N_15102,N_15106);
nand U15313 (N_15313,N_15188,N_15163);
nor U15314 (N_15314,N_15161,N_15138);
nand U15315 (N_15315,N_15113,N_15043);
or U15316 (N_15316,N_15132,N_15052);
nand U15317 (N_15317,N_15058,N_15041);
or U15318 (N_15318,N_15041,N_15077);
xor U15319 (N_15319,N_15168,N_15104);
nand U15320 (N_15320,N_15171,N_15084);
and U15321 (N_15321,N_15184,N_15078);
and U15322 (N_15322,N_15063,N_15173);
and U15323 (N_15323,N_15055,N_15085);
and U15324 (N_15324,N_15100,N_15170);
nor U15325 (N_15325,N_15164,N_15159);
nand U15326 (N_15326,N_15052,N_15156);
and U15327 (N_15327,N_15139,N_15132);
nand U15328 (N_15328,N_15109,N_15119);
nor U15329 (N_15329,N_15045,N_15178);
or U15330 (N_15330,N_15178,N_15161);
nor U15331 (N_15331,N_15156,N_15170);
nand U15332 (N_15332,N_15091,N_15041);
nand U15333 (N_15333,N_15047,N_15173);
and U15334 (N_15334,N_15175,N_15085);
nand U15335 (N_15335,N_15152,N_15049);
nor U15336 (N_15336,N_15101,N_15106);
and U15337 (N_15337,N_15040,N_15148);
nand U15338 (N_15338,N_15191,N_15131);
nand U15339 (N_15339,N_15075,N_15134);
nor U15340 (N_15340,N_15192,N_15075);
nand U15341 (N_15341,N_15056,N_15178);
xnor U15342 (N_15342,N_15148,N_15081);
and U15343 (N_15343,N_15106,N_15074);
or U15344 (N_15344,N_15044,N_15120);
or U15345 (N_15345,N_15052,N_15188);
and U15346 (N_15346,N_15066,N_15070);
and U15347 (N_15347,N_15195,N_15154);
and U15348 (N_15348,N_15180,N_15154);
and U15349 (N_15349,N_15073,N_15044);
nor U15350 (N_15350,N_15189,N_15072);
and U15351 (N_15351,N_15179,N_15119);
or U15352 (N_15352,N_15041,N_15089);
and U15353 (N_15353,N_15195,N_15062);
or U15354 (N_15354,N_15104,N_15068);
xor U15355 (N_15355,N_15194,N_15100);
xor U15356 (N_15356,N_15137,N_15094);
xor U15357 (N_15357,N_15044,N_15060);
nor U15358 (N_15358,N_15049,N_15157);
and U15359 (N_15359,N_15110,N_15166);
nor U15360 (N_15360,N_15287,N_15228);
or U15361 (N_15361,N_15315,N_15246);
and U15362 (N_15362,N_15298,N_15269);
nor U15363 (N_15363,N_15206,N_15350);
nand U15364 (N_15364,N_15279,N_15312);
nand U15365 (N_15365,N_15327,N_15204);
or U15366 (N_15366,N_15357,N_15282);
or U15367 (N_15367,N_15342,N_15321);
nor U15368 (N_15368,N_15245,N_15239);
and U15369 (N_15369,N_15233,N_15234);
xor U15370 (N_15370,N_15271,N_15274);
nand U15371 (N_15371,N_15232,N_15309);
xor U15372 (N_15372,N_15226,N_15345);
nand U15373 (N_15373,N_15248,N_15263);
nand U15374 (N_15374,N_15221,N_15349);
and U15375 (N_15375,N_15283,N_15316);
and U15376 (N_15376,N_15339,N_15218);
xnor U15377 (N_15377,N_15209,N_15241);
nand U15378 (N_15378,N_15268,N_15275);
xnor U15379 (N_15379,N_15305,N_15278);
or U15380 (N_15380,N_15277,N_15254);
or U15381 (N_15381,N_15343,N_15285);
xor U15382 (N_15382,N_15280,N_15223);
nand U15383 (N_15383,N_15205,N_15330);
nor U15384 (N_15384,N_15247,N_15208);
nor U15385 (N_15385,N_15224,N_15356);
xnor U15386 (N_15386,N_15346,N_15253);
or U15387 (N_15387,N_15212,N_15351);
or U15388 (N_15388,N_15251,N_15216);
nand U15389 (N_15389,N_15220,N_15313);
nor U15390 (N_15390,N_15261,N_15307);
xnor U15391 (N_15391,N_15272,N_15331);
or U15392 (N_15392,N_15213,N_15332);
xnor U15393 (N_15393,N_15334,N_15230);
and U15394 (N_15394,N_15352,N_15200);
nand U15395 (N_15395,N_15337,N_15244);
or U15396 (N_15396,N_15322,N_15333);
or U15397 (N_15397,N_15252,N_15243);
xor U15398 (N_15398,N_15324,N_15310);
xor U15399 (N_15399,N_15211,N_15242);
nor U15400 (N_15400,N_15266,N_15291);
or U15401 (N_15401,N_15219,N_15215);
nor U15402 (N_15402,N_15338,N_15348);
and U15403 (N_15403,N_15311,N_15264);
nor U15404 (N_15404,N_15344,N_15326);
nor U15405 (N_15405,N_15258,N_15217);
or U15406 (N_15406,N_15227,N_15329);
nor U15407 (N_15407,N_15259,N_15238);
and U15408 (N_15408,N_15340,N_15237);
xnor U15409 (N_15409,N_15301,N_15229);
xnor U15410 (N_15410,N_15202,N_15296);
nor U15411 (N_15411,N_15201,N_15265);
nand U15412 (N_15412,N_15293,N_15286);
or U15413 (N_15413,N_15308,N_15328);
xor U15414 (N_15414,N_15250,N_15323);
nand U15415 (N_15415,N_15267,N_15276);
nand U15416 (N_15416,N_15240,N_15222);
or U15417 (N_15417,N_15300,N_15347);
or U15418 (N_15418,N_15318,N_15236);
xor U15419 (N_15419,N_15292,N_15214);
nand U15420 (N_15420,N_15297,N_15358);
nor U15421 (N_15421,N_15255,N_15302);
or U15422 (N_15422,N_15325,N_15354);
and U15423 (N_15423,N_15306,N_15353);
and U15424 (N_15424,N_15335,N_15290);
or U15425 (N_15425,N_15231,N_15359);
and U15426 (N_15426,N_15262,N_15288);
nor U15427 (N_15427,N_15355,N_15207);
and U15428 (N_15428,N_15210,N_15295);
xnor U15429 (N_15429,N_15317,N_15336);
or U15430 (N_15430,N_15320,N_15294);
or U15431 (N_15431,N_15319,N_15273);
xnor U15432 (N_15432,N_15303,N_15257);
nand U15433 (N_15433,N_15284,N_15235);
or U15434 (N_15434,N_15225,N_15289);
or U15435 (N_15435,N_15270,N_15341);
xnor U15436 (N_15436,N_15281,N_15203);
and U15437 (N_15437,N_15256,N_15304);
nand U15438 (N_15438,N_15314,N_15260);
nand U15439 (N_15439,N_15299,N_15249);
and U15440 (N_15440,N_15249,N_15322);
nand U15441 (N_15441,N_15271,N_15237);
or U15442 (N_15442,N_15278,N_15204);
and U15443 (N_15443,N_15301,N_15306);
or U15444 (N_15444,N_15334,N_15325);
or U15445 (N_15445,N_15209,N_15332);
xor U15446 (N_15446,N_15276,N_15252);
nor U15447 (N_15447,N_15301,N_15311);
or U15448 (N_15448,N_15272,N_15333);
nor U15449 (N_15449,N_15264,N_15309);
nand U15450 (N_15450,N_15315,N_15312);
nand U15451 (N_15451,N_15224,N_15342);
or U15452 (N_15452,N_15254,N_15278);
nor U15453 (N_15453,N_15212,N_15263);
nor U15454 (N_15454,N_15328,N_15214);
and U15455 (N_15455,N_15296,N_15330);
and U15456 (N_15456,N_15308,N_15206);
nand U15457 (N_15457,N_15250,N_15230);
xnor U15458 (N_15458,N_15287,N_15333);
and U15459 (N_15459,N_15231,N_15241);
nor U15460 (N_15460,N_15277,N_15218);
xor U15461 (N_15461,N_15263,N_15271);
nand U15462 (N_15462,N_15233,N_15355);
and U15463 (N_15463,N_15243,N_15292);
or U15464 (N_15464,N_15210,N_15302);
or U15465 (N_15465,N_15287,N_15246);
nor U15466 (N_15466,N_15255,N_15237);
xnor U15467 (N_15467,N_15224,N_15253);
nor U15468 (N_15468,N_15349,N_15299);
nor U15469 (N_15469,N_15348,N_15304);
nand U15470 (N_15470,N_15221,N_15313);
and U15471 (N_15471,N_15326,N_15287);
xnor U15472 (N_15472,N_15299,N_15215);
or U15473 (N_15473,N_15256,N_15343);
and U15474 (N_15474,N_15253,N_15218);
and U15475 (N_15475,N_15273,N_15331);
nand U15476 (N_15476,N_15282,N_15227);
or U15477 (N_15477,N_15356,N_15234);
nor U15478 (N_15478,N_15254,N_15283);
nand U15479 (N_15479,N_15306,N_15295);
nor U15480 (N_15480,N_15288,N_15290);
or U15481 (N_15481,N_15329,N_15281);
nand U15482 (N_15482,N_15257,N_15318);
xor U15483 (N_15483,N_15252,N_15260);
xnor U15484 (N_15484,N_15284,N_15265);
xor U15485 (N_15485,N_15300,N_15267);
and U15486 (N_15486,N_15292,N_15213);
or U15487 (N_15487,N_15225,N_15304);
nand U15488 (N_15488,N_15358,N_15339);
or U15489 (N_15489,N_15245,N_15293);
xor U15490 (N_15490,N_15249,N_15310);
and U15491 (N_15491,N_15270,N_15336);
xor U15492 (N_15492,N_15345,N_15337);
nor U15493 (N_15493,N_15221,N_15348);
nor U15494 (N_15494,N_15262,N_15345);
xnor U15495 (N_15495,N_15279,N_15357);
and U15496 (N_15496,N_15290,N_15248);
nor U15497 (N_15497,N_15351,N_15345);
xor U15498 (N_15498,N_15352,N_15328);
xnor U15499 (N_15499,N_15215,N_15296);
xor U15500 (N_15500,N_15208,N_15227);
xnor U15501 (N_15501,N_15215,N_15200);
or U15502 (N_15502,N_15317,N_15258);
nand U15503 (N_15503,N_15210,N_15213);
xnor U15504 (N_15504,N_15227,N_15346);
nand U15505 (N_15505,N_15324,N_15239);
nand U15506 (N_15506,N_15264,N_15235);
nand U15507 (N_15507,N_15357,N_15274);
and U15508 (N_15508,N_15230,N_15201);
and U15509 (N_15509,N_15290,N_15302);
or U15510 (N_15510,N_15321,N_15276);
or U15511 (N_15511,N_15237,N_15280);
or U15512 (N_15512,N_15307,N_15243);
and U15513 (N_15513,N_15222,N_15234);
nand U15514 (N_15514,N_15347,N_15293);
xnor U15515 (N_15515,N_15284,N_15343);
or U15516 (N_15516,N_15224,N_15320);
nand U15517 (N_15517,N_15272,N_15239);
nand U15518 (N_15518,N_15349,N_15263);
or U15519 (N_15519,N_15327,N_15245);
and U15520 (N_15520,N_15368,N_15385);
nor U15521 (N_15521,N_15467,N_15471);
xnor U15522 (N_15522,N_15472,N_15429);
nand U15523 (N_15523,N_15482,N_15464);
or U15524 (N_15524,N_15458,N_15455);
nor U15525 (N_15525,N_15519,N_15483);
or U15526 (N_15526,N_15360,N_15364);
nor U15527 (N_15527,N_15410,N_15461);
nor U15528 (N_15528,N_15505,N_15407);
xnor U15529 (N_15529,N_15463,N_15476);
nand U15530 (N_15530,N_15431,N_15371);
or U15531 (N_15531,N_15433,N_15457);
and U15532 (N_15532,N_15511,N_15363);
xor U15533 (N_15533,N_15479,N_15456);
and U15534 (N_15534,N_15388,N_15517);
xnor U15535 (N_15535,N_15462,N_15400);
xor U15536 (N_15536,N_15512,N_15450);
nor U15537 (N_15537,N_15460,N_15379);
nor U15538 (N_15538,N_15372,N_15504);
nand U15539 (N_15539,N_15503,N_15393);
or U15540 (N_15540,N_15432,N_15397);
and U15541 (N_15541,N_15489,N_15493);
or U15542 (N_15542,N_15438,N_15436);
xor U15543 (N_15543,N_15391,N_15448);
and U15544 (N_15544,N_15477,N_15447);
nor U15545 (N_15545,N_15496,N_15497);
and U15546 (N_15546,N_15500,N_15446);
nor U15547 (N_15547,N_15405,N_15403);
nand U15548 (N_15548,N_15387,N_15492);
nor U15549 (N_15549,N_15389,N_15509);
xor U15550 (N_15550,N_15418,N_15502);
nand U15551 (N_15551,N_15424,N_15474);
and U15552 (N_15552,N_15395,N_15392);
nor U15553 (N_15553,N_15486,N_15494);
or U15554 (N_15554,N_15453,N_15430);
nor U15555 (N_15555,N_15487,N_15390);
xnor U15556 (N_15556,N_15399,N_15411);
or U15557 (N_15557,N_15484,N_15377);
or U15558 (N_15558,N_15499,N_15518);
and U15559 (N_15559,N_15480,N_15386);
nor U15560 (N_15560,N_15449,N_15401);
nand U15561 (N_15561,N_15445,N_15415);
and U15562 (N_15562,N_15382,N_15435);
or U15563 (N_15563,N_15459,N_15422);
or U15564 (N_15564,N_15485,N_15427);
and U15565 (N_15565,N_15375,N_15394);
nand U15566 (N_15566,N_15370,N_15423);
and U15567 (N_15567,N_15417,N_15369);
nand U15568 (N_15568,N_15490,N_15443);
nor U15569 (N_15569,N_15406,N_15506);
or U15570 (N_15570,N_15404,N_15426);
or U15571 (N_15571,N_15469,N_15441);
and U15572 (N_15572,N_15380,N_15473);
nand U15573 (N_15573,N_15416,N_15442);
and U15574 (N_15574,N_15381,N_15374);
xor U15575 (N_15575,N_15488,N_15398);
nor U15576 (N_15576,N_15491,N_15444);
xor U15577 (N_15577,N_15470,N_15366);
or U15578 (N_15578,N_15516,N_15454);
and U15579 (N_15579,N_15439,N_15507);
or U15580 (N_15580,N_15412,N_15373);
xor U15581 (N_15581,N_15396,N_15384);
nor U15582 (N_15582,N_15440,N_15515);
and U15583 (N_15583,N_15428,N_15437);
and U15584 (N_15584,N_15475,N_15495);
nor U15585 (N_15585,N_15452,N_15421);
xnor U15586 (N_15586,N_15513,N_15383);
xor U15587 (N_15587,N_15409,N_15465);
xnor U15588 (N_15588,N_15419,N_15466);
nor U15589 (N_15589,N_15510,N_15481);
or U15590 (N_15590,N_15420,N_15365);
nor U15591 (N_15591,N_15508,N_15367);
xnor U15592 (N_15592,N_15361,N_15402);
nand U15593 (N_15593,N_15425,N_15413);
nor U15594 (N_15594,N_15362,N_15498);
nand U15595 (N_15595,N_15434,N_15501);
or U15596 (N_15596,N_15408,N_15514);
xor U15597 (N_15597,N_15414,N_15376);
or U15598 (N_15598,N_15468,N_15478);
nor U15599 (N_15599,N_15451,N_15378);
nand U15600 (N_15600,N_15492,N_15468);
or U15601 (N_15601,N_15418,N_15481);
xnor U15602 (N_15602,N_15455,N_15507);
nor U15603 (N_15603,N_15405,N_15495);
or U15604 (N_15604,N_15452,N_15380);
nor U15605 (N_15605,N_15498,N_15437);
xor U15606 (N_15606,N_15493,N_15500);
nor U15607 (N_15607,N_15430,N_15367);
xor U15608 (N_15608,N_15400,N_15363);
xnor U15609 (N_15609,N_15501,N_15459);
or U15610 (N_15610,N_15392,N_15377);
nor U15611 (N_15611,N_15413,N_15365);
nand U15612 (N_15612,N_15434,N_15473);
xor U15613 (N_15613,N_15437,N_15499);
and U15614 (N_15614,N_15454,N_15503);
xor U15615 (N_15615,N_15372,N_15495);
nand U15616 (N_15616,N_15369,N_15436);
nand U15617 (N_15617,N_15485,N_15382);
xnor U15618 (N_15618,N_15379,N_15386);
nand U15619 (N_15619,N_15460,N_15418);
nand U15620 (N_15620,N_15397,N_15467);
nand U15621 (N_15621,N_15508,N_15446);
nor U15622 (N_15622,N_15514,N_15435);
nor U15623 (N_15623,N_15373,N_15411);
xor U15624 (N_15624,N_15490,N_15475);
nor U15625 (N_15625,N_15507,N_15395);
and U15626 (N_15626,N_15452,N_15487);
and U15627 (N_15627,N_15460,N_15387);
nand U15628 (N_15628,N_15373,N_15456);
or U15629 (N_15629,N_15365,N_15363);
and U15630 (N_15630,N_15424,N_15449);
nor U15631 (N_15631,N_15365,N_15474);
xnor U15632 (N_15632,N_15490,N_15495);
or U15633 (N_15633,N_15370,N_15392);
xnor U15634 (N_15634,N_15365,N_15490);
nand U15635 (N_15635,N_15398,N_15460);
or U15636 (N_15636,N_15491,N_15468);
or U15637 (N_15637,N_15475,N_15395);
and U15638 (N_15638,N_15492,N_15461);
xnor U15639 (N_15639,N_15383,N_15494);
and U15640 (N_15640,N_15465,N_15449);
and U15641 (N_15641,N_15425,N_15415);
xor U15642 (N_15642,N_15379,N_15510);
nor U15643 (N_15643,N_15393,N_15517);
nor U15644 (N_15644,N_15438,N_15399);
nor U15645 (N_15645,N_15449,N_15417);
nor U15646 (N_15646,N_15368,N_15390);
or U15647 (N_15647,N_15479,N_15512);
xor U15648 (N_15648,N_15477,N_15471);
nand U15649 (N_15649,N_15452,N_15428);
or U15650 (N_15650,N_15514,N_15399);
and U15651 (N_15651,N_15437,N_15432);
nand U15652 (N_15652,N_15381,N_15426);
nand U15653 (N_15653,N_15463,N_15387);
and U15654 (N_15654,N_15381,N_15369);
nand U15655 (N_15655,N_15472,N_15494);
and U15656 (N_15656,N_15394,N_15428);
or U15657 (N_15657,N_15364,N_15477);
xor U15658 (N_15658,N_15428,N_15448);
and U15659 (N_15659,N_15419,N_15437);
or U15660 (N_15660,N_15427,N_15469);
nor U15661 (N_15661,N_15480,N_15460);
nor U15662 (N_15662,N_15470,N_15392);
and U15663 (N_15663,N_15434,N_15385);
xor U15664 (N_15664,N_15454,N_15465);
nand U15665 (N_15665,N_15431,N_15408);
nor U15666 (N_15666,N_15386,N_15360);
and U15667 (N_15667,N_15486,N_15452);
or U15668 (N_15668,N_15450,N_15412);
nand U15669 (N_15669,N_15483,N_15402);
or U15670 (N_15670,N_15405,N_15457);
xor U15671 (N_15671,N_15497,N_15481);
xor U15672 (N_15672,N_15374,N_15461);
nand U15673 (N_15673,N_15484,N_15427);
nor U15674 (N_15674,N_15377,N_15410);
or U15675 (N_15675,N_15445,N_15462);
nand U15676 (N_15676,N_15378,N_15404);
nor U15677 (N_15677,N_15476,N_15414);
or U15678 (N_15678,N_15449,N_15416);
nand U15679 (N_15679,N_15388,N_15494);
or U15680 (N_15680,N_15572,N_15604);
nand U15681 (N_15681,N_15562,N_15640);
and U15682 (N_15682,N_15524,N_15593);
nand U15683 (N_15683,N_15554,N_15653);
and U15684 (N_15684,N_15590,N_15614);
nor U15685 (N_15685,N_15581,N_15664);
nor U15686 (N_15686,N_15600,N_15673);
and U15687 (N_15687,N_15676,N_15542);
nand U15688 (N_15688,N_15582,N_15547);
or U15689 (N_15689,N_15599,N_15650);
nor U15690 (N_15690,N_15571,N_15656);
nand U15691 (N_15691,N_15598,N_15669);
xor U15692 (N_15692,N_15560,N_15566);
and U15693 (N_15693,N_15548,N_15678);
xor U15694 (N_15694,N_15601,N_15521);
nand U15695 (N_15695,N_15575,N_15657);
and U15696 (N_15696,N_15567,N_15636);
nor U15697 (N_15697,N_15563,N_15674);
nand U15698 (N_15698,N_15632,N_15620);
or U15699 (N_15699,N_15606,N_15610);
or U15700 (N_15700,N_15553,N_15668);
nor U15701 (N_15701,N_15667,N_15602);
xor U15702 (N_15702,N_15580,N_15556);
nor U15703 (N_15703,N_15536,N_15534);
nand U15704 (N_15704,N_15609,N_15586);
nand U15705 (N_15705,N_15597,N_15613);
and U15706 (N_15706,N_15579,N_15647);
nor U15707 (N_15707,N_15639,N_15635);
xor U15708 (N_15708,N_15520,N_15655);
and U15709 (N_15709,N_15629,N_15659);
and U15710 (N_15710,N_15570,N_15584);
xnor U15711 (N_15711,N_15543,N_15527);
and U15712 (N_15712,N_15589,N_15555);
or U15713 (N_15713,N_15643,N_15627);
or U15714 (N_15714,N_15546,N_15612);
nor U15715 (N_15715,N_15595,N_15675);
nor U15716 (N_15716,N_15535,N_15551);
nor U15717 (N_15717,N_15622,N_15568);
nor U15718 (N_15718,N_15671,N_15644);
or U15719 (N_15719,N_15528,N_15561);
xnor U15720 (N_15720,N_15619,N_15574);
and U15721 (N_15721,N_15558,N_15523);
or U15722 (N_15722,N_15658,N_15633);
and U15723 (N_15723,N_15670,N_15615);
xnor U15724 (N_15724,N_15677,N_15578);
or U15725 (N_15725,N_15666,N_15594);
and U15726 (N_15726,N_15541,N_15611);
or U15727 (N_15727,N_15652,N_15564);
or U15728 (N_15728,N_15544,N_15565);
and U15729 (N_15729,N_15596,N_15569);
or U15730 (N_15730,N_15641,N_15645);
or U15731 (N_15731,N_15577,N_15663);
or U15732 (N_15732,N_15559,N_15625);
or U15733 (N_15733,N_15634,N_15549);
nor U15734 (N_15734,N_15646,N_15624);
nand U15735 (N_15735,N_15617,N_15616);
nor U15736 (N_15736,N_15530,N_15637);
or U15737 (N_15737,N_15607,N_15638);
nand U15738 (N_15738,N_15603,N_15679);
and U15739 (N_15739,N_15651,N_15605);
nor U15740 (N_15740,N_15533,N_15660);
nand U15741 (N_15741,N_15626,N_15592);
xor U15742 (N_15742,N_15531,N_15585);
or U15743 (N_15743,N_15608,N_15538);
or U15744 (N_15744,N_15552,N_15532);
nor U15745 (N_15745,N_15661,N_15662);
or U15746 (N_15746,N_15588,N_15583);
nor U15747 (N_15747,N_15648,N_15529);
nand U15748 (N_15748,N_15654,N_15537);
xnor U15749 (N_15749,N_15628,N_15525);
and U15750 (N_15750,N_15545,N_15621);
and U15751 (N_15751,N_15550,N_15573);
xnor U15752 (N_15752,N_15526,N_15557);
xor U15753 (N_15753,N_15672,N_15631);
nand U15754 (N_15754,N_15540,N_15618);
xnor U15755 (N_15755,N_15649,N_15665);
or U15756 (N_15756,N_15591,N_15587);
or U15757 (N_15757,N_15642,N_15623);
nand U15758 (N_15758,N_15630,N_15539);
or U15759 (N_15759,N_15522,N_15576);
nand U15760 (N_15760,N_15521,N_15583);
nor U15761 (N_15761,N_15596,N_15616);
and U15762 (N_15762,N_15582,N_15543);
nor U15763 (N_15763,N_15658,N_15651);
nand U15764 (N_15764,N_15540,N_15574);
nor U15765 (N_15765,N_15629,N_15562);
or U15766 (N_15766,N_15606,N_15599);
or U15767 (N_15767,N_15582,N_15552);
nand U15768 (N_15768,N_15623,N_15622);
nor U15769 (N_15769,N_15569,N_15523);
xor U15770 (N_15770,N_15620,N_15629);
or U15771 (N_15771,N_15647,N_15669);
nor U15772 (N_15772,N_15539,N_15578);
nor U15773 (N_15773,N_15597,N_15526);
nor U15774 (N_15774,N_15570,N_15652);
xor U15775 (N_15775,N_15600,N_15521);
or U15776 (N_15776,N_15536,N_15667);
nor U15777 (N_15777,N_15622,N_15577);
xor U15778 (N_15778,N_15521,N_15541);
nand U15779 (N_15779,N_15551,N_15656);
nand U15780 (N_15780,N_15535,N_15625);
nor U15781 (N_15781,N_15592,N_15589);
nor U15782 (N_15782,N_15582,N_15560);
xnor U15783 (N_15783,N_15634,N_15618);
nor U15784 (N_15784,N_15591,N_15647);
or U15785 (N_15785,N_15673,N_15537);
xor U15786 (N_15786,N_15538,N_15523);
or U15787 (N_15787,N_15567,N_15545);
nand U15788 (N_15788,N_15573,N_15638);
nor U15789 (N_15789,N_15611,N_15606);
or U15790 (N_15790,N_15564,N_15647);
nand U15791 (N_15791,N_15663,N_15671);
and U15792 (N_15792,N_15523,N_15585);
nand U15793 (N_15793,N_15657,N_15579);
or U15794 (N_15794,N_15649,N_15551);
nand U15795 (N_15795,N_15596,N_15552);
nand U15796 (N_15796,N_15585,N_15621);
xor U15797 (N_15797,N_15658,N_15530);
nor U15798 (N_15798,N_15636,N_15622);
nor U15799 (N_15799,N_15672,N_15639);
nor U15800 (N_15800,N_15536,N_15663);
xor U15801 (N_15801,N_15612,N_15547);
nand U15802 (N_15802,N_15549,N_15592);
nand U15803 (N_15803,N_15523,N_15608);
nor U15804 (N_15804,N_15672,N_15566);
or U15805 (N_15805,N_15658,N_15556);
or U15806 (N_15806,N_15556,N_15648);
nand U15807 (N_15807,N_15602,N_15603);
and U15808 (N_15808,N_15541,N_15673);
and U15809 (N_15809,N_15670,N_15592);
nand U15810 (N_15810,N_15599,N_15615);
or U15811 (N_15811,N_15672,N_15633);
and U15812 (N_15812,N_15606,N_15679);
xnor U15813 (N_15813,N_15668,N_15611);
or U15814 (N_15814,N_15610,N_15586);
or U15815 (N_15815,N_15520,N_15600);
and U15816 (N_15816,N_15617,N_15557);
nand U15817 (N_15817,N_15555,N_15671);
nand U15818 (N_15818,N_15677,N_15641);
xor U15819 (N_15819,N_15589,N_15649);
or U15820 (N_15820,N_15645,N_15562);
nand U15821 (N_15821,N_15629,N_15549);
and U15822 (N_15822,N_15573,N_15627);
nand U15823 (N_15823,N_15560,N_15637);
and U15824 (N_15824,N_15660,N_15575);
or U15825 (N_15825,N_15620,N_15656);
nor U15826 (N_15826,N_15602,N_15660);
nand U15827 (N_15827,N_15539,N_15587);
xnor U15828 (N_15828,N_15561,N_15525);
xnor U15829 (N_15829,N_15618,N_15599);
xnor U15830 (N_15830,N_15647,N_15523);
or U15831 (N_15831,N_15583,N_15631);
and U15832 (N_15832,N_15651,N_15617);
xnor U15833 (N_15833,N_15569,N_15620);
nand U15834 (N_15834,N_15572,N_15603);
nor U15835 (N_15835,N_15559,N_15552);
nor U15836 (N_15836,N_15600,N_15641);
nand U15837 (N_15837,N_15522,N_15558);
nor U15838 (N_15838,N_15662,N_15641);
and U15839 (N_15839,N_15662,N_15566);
xnor U15840 (N_15840,N_15749,N_15808);
or U15841 (N_15841,N_15722,N_15703);
nor U15842 (N_15842,N_15702,N_15830);
nand U15843 (N_15843,N_15762,N_15800);
nand U15844 (N_15844,N_15816,N_15799);
or U15845 (N_15845,N_15750,N_15780);
or U15846 (N_15846,N_15769,N_15701);
nand U15847 (N_15847,N_15795,N_15828);
xor U15848 (N_15848,N_15711,N_15774);
or U15849 (N_15849,N_15777,N_15687);
xnor U15850 (N_15850,N_15834,N_15747);
nand U15851 (N_15851,N_15761,N_15694);
nand U15852 (N_15852,N_15730,N_15721);
xnor U15853 (N_15853,N_15806,N_15746);
and U15854 (N_15854,N_15740,N_15832);
nand U15855 (N_15855,N_15752,N_15698);
and U15856 (N_15856,N_15801,N_15838);
and U15857 (N_15857,N_15829,N_15684);
and U15858 (N_15858,N_15712,N_15839);
or U15859 (N_15859,N_15757,N_15803);
nor U15860 (N_15860,N_15727,N_15728);
nand U15861 (N_15861,N_15734,N_15812);
nor U15862 (N_15862,N_15726,N_15741);
or U15863 (N_15863,N_15798,N_15809);
or U15864 (N_15864,N_15735,N_15778);
or U15865 (N_15865,N_15745,N_15732);
xor U15866 (N_15866,N_15715,N_15833);
xor U15867 (N_15867,N_15689,N_15725);
nand U15868 (N_15868,N_15771,N_15784);
nand U15869 (N_15869,N_15794,N_15724);
xnor U15870 (N_15870,N_15713,N_15768);
xnor U15871 (N_15871,N_15688,N_15797);
or U15872 (N_15872,N_15707,N_15737);
nand U15873 (N_15873,N_15705,N_15815);
nor U15874 (N_15874,N_15736,N_15789);
xnor U15875 (N_15875,N_15699,N_15802);
or U15876 (N_15876,N_15765,N_15779);
xnor U15877 (N_15877,N_15782,N_15739);
xnor U15878 (N_15878,N_15783,N_15720);
xor U15879 (N_15879,N_15710,N_15796);
or U15880 (N_15880,N_15755,N_15793);
nor U15881 (N_15881,N_15810,N_15743);
and U15882 (N_15882,N_15776,N_15742);
or U15883 (N_15883,N_15729,N_15763);
nor U15884 (N_15884,N_15696,N_15823);
or U15885 (N_15885,N_15824,N_15709);
or U15886 (N_15886,N_15818,N_15718);
nand U15887 (N_15887,N_15772,N_15686);
and U15888 (N_15888,N_15825,N_15773);
xor U15889 (N_15889,N_15717,N_15819);
xnor U15890 (N_15890,N_15814,N_15813);
nor U15891 (N_15891,N_15831,N_15708);
xor U15892 (N_15892,N_15682,N_15837);
and U15893 (N_15893,N_15706,N_15683);
and U15894 (N_15894,N_15822,N_15692);
xnor U15895 (N_15895,N_15754,N_15744);
nor U15896 (N_15896,N_15785,N_15690);
nor U15897 (N_15897,N_15693,N_15767);
xnor U15898 (N_15898,N_15826,N_15748);
nand U15899 (N_15899,N_15770,N_15821);
or U15900 (N_15900,N_15817,N_15805);
xor U15901 (N_15901,N_15714,N_15790);
and U15902 (N_15902,N_15716,N_15723);
or U15903 (N_15903,N_15764,N_15781);
nand U15904 (N_15904,N_15719,N_15704);
xnor U15905 (N_15905,N_15788,N_15751);
xnor U15906 (N_15906,N_15807,N_15691);
nand U15907 (N_15907,N_15820,N_15681);
and U15908 (N_15908,N_15760,N_15731);
nand U15909 (N_15909,N_15685,N_15753);
and U15910 (N_15910,N_15836,N_15738);
nor U15911 (N_15911,N_15804,N_15697);
xnor U15912 (N_15912,N_15792,N_15811);
and U15913 (N_15913,N_15695,N_15759);
nor U15914 (N_15914,N_15775,N_15733);
nand U15915 (N_15915,N_15766,N_15758);
xnor U15916 (N_15916,N_15827,N_15680);
xor U15917 (N_15917,N_15756,N_15787);
xnor U15918 (N_15918,N_15791,N_15786);
and U15919 (N_15919,N_15700,N_15835);
nand U15920 (N_15920,N_15684,N_15734);
or U15921 (N_15921,N_15816,N_15782);
or U15922 (N_15922,N_15776,N_15804);
xnor U15923 (N_15923,N_15774,N_15810);
or U15924 (N_15924,N_15727,N_15818);
nand U15925 (N_15925,N_15683,N_15760);
and U15926 (N_15926,N_15736,N_15798);
and U15927 (N_15927,N_15700,N_15690);
xor U15928 (N_15928,N_15752,N_15696);
or U15929 (N_15929,N_15772,N_15770);
or U15930 (N_15930,N_15778,N_15796);
nand U15931 (N_15931,N_15708,N_15763);
and U15932 (N_15932,N_15690,N_15789);
nor U15933 (N_15933,N_15823,N_15692);
or U15934 (N_15934,N_15834,N_15698);
nor U15935 (N_15935,N_15790,N_15809);
and U15936 (N_15936,N_15745,N_15722);
or U15937 (N_15937,N_15691,N_15802);
nor U15938 (N_15938,N_15760,N_15699);
or U15939 (N_15939,N_15808,N_15802);
and U15940 (N_15940,N_15772,N_15688);
or U15941 (N_15941,N_15805,N_15757);
or U15942 (N_15942,N_15746,N_15718);
nor U15943 (N_15943,N_15826,N_15812);
xnor U15944 (N_15944,N_15744,N_15763);
or U15945 (N_15945,N_15788,N_15754);
and U15946 (N_15946,N_15697,N_15683);
or U15947 (N_15947,N_15790,N_15833);
nor U15948 (N_15948,N_15799,N_15694);
or U15949 (N_15949,N_15790,N_15836);
nand U15950 (N_15950,N_15746,N_15808);
nor U15951 (N_15951,N_15722,N_15816);
or U15952 (N_15952,N_15738,N_15780);
nor U15953 (N_15953,N_15721,N_15739);
nor U15954 (N_15954,N_15834,N_15709);
xor U15955 (N_15955,N_15741,N_15804);
nor U15956 (N_15956,N_15815,N_15746);
nor U15957 (N_15957,N_15757,N_15786);
nor U15958 (N_15958,N_15700,N_15682);
or U15959 (N_15959,N_15683,N_15834);
nor U15960 (N_15960,N_15759,N_15694);
nand U15961 (N_15961,N_15753,N_15826);
xnor U15962 (N_15962,N_15743,N_15829);
or U15963 (N_15963,N_15711,N_15836);
xnor U15964 (N_15964,N_15695,N_15828);
and U15965 (N_15965,N_15791,N_15766);
and U15966 (N_15966,N_15814,N_15721);
and U15967 (N_15967,N_15748,N_15683);
nand U15968 (N_15968,N_15832,N_15762);
nor U15969 (N_15969,N_15683,N_15687);
xnor U15970 (N_15970,N_15820,N_15751);
nand U15971 (N_15971,N_15731,N_15699);
xnor U15972 (N_15972,N_15799,N_15743);
or U15973 (N_15973,N_15809,N_15780);
nand U15974 (N_15974,N_15827,N_15753);
and U15975 (N_15975,N_15722,N_15735);
xor U15976 (N_15976,N_15777,N_15717);
xor U15977 (N_15977,N_15834,N_15788);
nand U15978 (N_15978,N_15781,N_15748);
and U15979 (N_15979,N_15725,N_15730);
and U15980 (N_15980,N_15702,N_15738);
and U15981 (N_15981,N_15778,N_15716);
and U15982 (N_15982,N_15705,N_15691);
nor U15983 (N_15983,N_15834,N_15696);
or U15984 (N_15984,N_15727,N_15774);
or U15985 (N_15985,N_15697,N_15823);
and U15986 (N_15986,N_15748,N_15811);
nor U15987 (N_15987,N_15698,N_15729);
nor U15988 (N_15988,N_15799,N_15689);
or U15989 (N_15989,N_15746,N_15714);
and U15990 (N_15990,N_15804,N_15825);
or U15991 (N_15991,N_15828,N_15838);
and U15992 (N_15992,N_15813,N_15793);
nor U15993 (N_15993,N_15792,N_15796);
nand U15994 (N_15994,N_15814,N_15742);
or U15995 (N_15995,N_15794,N_15831);
nor U15996 (N_15996,N_15712,N_15751);
xor U15997 (N_15997,N_15743,N_15800);
or U15998 (N_15998,N_15721,N_15708);
and U15999 (N_15999,N_15723,N_15764);
nor U16000 (N_16000,N_15977,N_15852);
nor U16001 (N_16001,N_15935,N_15884);
nand U16002 (N_16002,N_15889,N_15911);
nor U16003 (N_16003,N_15849,N_15943);
or U16004 (N_16004,N_15865,N_15879);
xor U16005 (N_16005,N_15959,N_15910);
and U16006 (N_16006,N_15897,N_15895);
or U16007 (N_16007,N_15909,N_15976);
nor U16008 (N_16008,N_15987,N_15948);
nand U16009 (N_16009,N_15988,N_15929);
xnor U16010 (N_16010,N_15967,N_15860);
xor U16011 (N_16011,N_15876,N_15871);
nand U16012 (N_16012,N_15949,N_15985);
nor U16013 (N_16013,N_15961,N_15893);
nand U16014 (N_16014,N_15858,N_15844);
and U16015 (N_16015,N_15857,N_15965);
and U16016 (N_16016,N_15963,N_15957);
xnor U16017 (N_16017,N_15846,N_15850);
and U16018 (N_16018,N_15980,N_15908);
nand U16019 (N_16019,N_15989,N_15937);
nor U16020 (N_16020,N_15996,N_15950);
xor U16021 (N_16021,N_15870,N_15969);
or U16022 (N_16022,N_15966,N_15917);
or U16023 (N_16023,N_15938,N_15899);
or U16024 (N_16024,N_15962,N_15918);
or U16025 (N_16025,N_15859,N_15971);
or U16026 (N_16026,N_15984,N_15933);
nor U16027 (N_16027,N_15885,N_15873);
xnor U16028 (N_16028,N_15999,N_15974);
nand U16029 (N_16029,N_15941,N_15851);
or U16030 (N_16030,N_15880,N_15970);
or U16031 (N_16031,N_15914,N_15925);
nand U16032 (N_16032,N_15892,N_15928);
and U16033 (N_16033,N_15845,N_15923);
or U16034 (N_16034,N_15978,N_15956);
nor U16035 (N_16035,N_15993,N_15958);
xnor U16036 (N_16036,N_15866,N_15868);
or U16037 (N_16037,N_15861,N_15912);
xnor U16038 (N_16038,N_15853,N_15942);
xor U16039 (N_16039,N_15916,N_15926);
nand U16040 (N_16040,N_15875,N_15840);
and U16041 (N_16041,N_15945,N_15997);
nor U16042 (N_16042,N_15972,N_15887);
xor U16043 (N_16043,N_15924,N_15904);
nor U16044 (N_16044,N_15856,N_15964);
nand U16045 (N_16045,N_15855,N_15862);
nand U16046 (N_16046,N_15847,N_15843);
and U16047 (N_16047,N_15883,N_15952);
or U16048 (N_16048,N_15936,N_15975);
nand U16049 (N_16049,N_15901,N_15944);
nor U16050 (N_16050,N_15960,N_15932);
xor U16051 (N_16051,N_15915,N_15968);
xor U16052 (N_16052,N_15934,N_15927);
xnor U16053 (N_16053,N_15854,N_15842);
xor U16054 (N_16054,N_15869,N_15913);
and U16055 (N_16055,N_15921,N_15994);
and U16056 (N_16056,N_15905,N_15907);
or U16057 (N_16057,N_15951,N_15947);
nand U16058 (N_16058,N_15891,N_15983);
or U16059 (N_16059,N_15898,N_15848);
and U16060 (N_16060,N_15903,N_15981);
or U16061 (N_16061,N_15955,N_15864);
nor U16062 (N_16062,N_15882,N_15973);
or U16063 (N_16063,N_15881,N_15986);
or U16064 (N_16064,N_15982,N_15922);
or U16065 (N_16065,N_15878,N_15930);
and U16066 (N_16066,N_15919,N_15863);
or U16067 (N_16067,N_15939,N_15920);
xnor U16068 (N_16068,N_15890,N_15998);
or U16069 (N_16069,N_15900,N_15872);
nand U16070 (N_16070,N_15894,N_15954);
nor U16071 (N_16071,N_15953,N_15867);
xnor U16072 (N_16072,N_15979,N_15888);
nor U16073 (N_16073,N_15940,N_15886);
nand U16074 (N_16074,N_15877,N_15906);
nand U16075 (N_16075,N_15992,N_15841);
nor U16076 (N_16076,N_15990,N_15931);
and U16077 (N_16077,N_15946,N_15991);
and U16078 (N_16078,N_15874,N_15902);
xnor U16079 (N_16079,N_15995,N_15896);
xor U16080 (N_16080,N_15986,N_15947);
and U16081 (N_16081,N_15899,N_15909);
nor U16082 (N_16082,N_15910,N_15888);
nand U16083 (N_16083,N_15931,N_15851);
and U16084 (N_16084,N_15878,N_15931);
xnor U16085 (N_16085,N_15867,N_15989);
xor U16086 (N_16086,N_15918,N_15855);
and U16087 (N_16087,N_15949,N_15959);
nand U16088 (N_16088,N_15960,N_15973);
or U16089 (N_16089,N_15984,N_15915);
or U16090 (N_16090,N_15969,N_15846);
or U16091 (N_16091,N_15854,N_15965);
nor U16092 (N_16092,N_15948,N_15865);
xnor U16093 (N_16093,N_15988,N_15978);
nor U16094 (N_16094,N_15868,N_15977);
and U16095 (N_16095,N_15971,N_15994);
and U16096 (N_16096,N_15922,N_15847);
nor U16097 (N_16097,N_15849,N_15972);
nor U16098 (N_16098,N_15912,N_15862);
and U16099 (N_16099,N_15920,N_15879);
or U16100 (N_16100,N_15938,N_15890);
and U16101 (N_16101,N_15871,N_15862);
xor U16102 (N_16102,N_15892,N_15987);
nand U16103 (N_16103,N_15968,N_15903);
or U16104 (N_16104,N_15896,N_15885);
and U16105 (N_16105,N_15877,N_15946);
or U16106 (N_16106,N_15902,N_15979);
and U16107 (N_16107,N_15999,N_15905);
nand U16108 (N_16108,N_15913,N_15846);
and U16109 (N_16109,N_15963,N_15858);
xnor U16110 (N_16110,N_15925,N_15871);
nand U16111 (N_16111,N_15917,N_15844);
or U16112 (N_16112,N_15903,N_15921);
xnor U16113 (N_16113,N_15993,N_15941);
xor U16114 (N_16114,N_15918,N_15872);
xnor U16115 (N_16115,N_15840,N_15918);
and U16116 (N_16116,N_15941,N_15996);
xnor U16117 (N_16117,N_15917,N_15880);
and U16118 (N_16118,N_15908,N_15867);
nor U16119 (N_16119,N_15994,N_15846);
xor U16120 (N_16120,N_15921,N_15853);
and U16121 (N_16121,N_15964,N_15928);
nand U16122 (N_16122,N_15864,N_15988);
and U16123 (N_16123,N_15926,N_15870);
or U16124 (N_16124,N_15991,N_15969);
nor U16125 (N_16125,N_15887,N_15950);
or U16126 (N_16126,N_15962,N_15983);
nand U16127 (N_16127,N_15982,N_15840);
or U16128 (N_16128,N_15886,N_15957);
or U16129 (N_16129,N_15865,N_15861);
xnor U16130 (N_16130,N_15909,N_15962);
nand U16131 (N_16131,N_15942,N_15981);
nor U16132 (N_16132,N_15898,N_15921);
and U16133 (N_16133,N_15864,N_15859);
and U16134 (N_16134,N_15991,N_15999);
or U16135 (N_16135,N_15865,N_15894);
or U16136 (N_16136,N_15976,N_15882);
nand U16137 (N_16137,N_15939,N_15840);
nor U16138 (N_16138,N_15975,N_15974);
or U16139 (N_16139,N_15924,N_15958);
xnor U16140 (N_16140,N_15851,N_15894);
and U16141 (N_16141,N_15978,N_15951);
nand U16142 (N_16142,N_15990,N_15907);
and U16143 (N_16143,N_15871,N_15921);
or U16144 (N_16144,N_15891,N_15861);
nand U16145 (N_16145,N_15906,N_15845);
xor U16146 (N_16146,N_15937,N_15969);
or U16147 (N_16147,N_15951,N_15871);
xnor U16148 (N_16148,N_15934,N_15945);
nor U16149 (N_16149,N_15953,N_15965);
and U16150 (N_16150,N_15886,N_15903);
xnor U16151 (N_16151,N_15996,N_15843);
nor U16152 (N_16152,N_15907,N_15854);
nor U16153 (N_16153,N_15968,N_15873);
nand U16154 (N_16154,N_15911,N_15845);
nand U16155 (N_16155,N_15879,N_15896);
xnor U16156 (N_16156,N_15871,N_15997);
or U16157 (N_16157,N_15880,N_15984);
nor U16158 (N_16158,N_15862,N_15939);
or U16159 (N_16159,N_15933,N_15842);
xnor U16160 (N_16160,N_16101,N_16153);
nand U16161 (N_16161,N_16097,N_16110);
or U16162 (N_16162,N_16109,N_16134);
nor U16163 (N_16163,N_16061,N_16130);
xnor U16164 (N_16164,N_16062,N_16042);
and U16165 (N_16165,N_16142,N_16125);
or U16166 (N_16166,N_16005,N_16149);
nand U16167 (N_16167,N_16091,N_16032);
and U16168 (N_16168,N_16145,N_16148);
xnor U16169 (N_16169,N_16004,N_16045);
nand U16170 (N_16170,N_16111,N_16106);
nor U16171 (N_16171,N_16049,N_16003);
or U16172 (N_16172,N_16132,N_16117);
nor U16173 (N_16173,N_16031,N_16055);
nand U16174 (N_16174,N_16017,N_16026);
nand U16175 (N_16175,N_16126,N_16064);
xor U16176 (N_16176,N_16096,N_16120);
and U16177 (N_16177,N_16104,N_16116);
and U16178 (N_16178,N_16054,N_16113);
nor U16179 (N_16179,N_16155,N_16011);
or U16180 (N_16180,N_16006,N_16037);
and U16181 (N_16181,N_16139,N_16025);
and U16182 (N_16182,N_16123,N_16100);
or U16183 (N_16183,N_16141,N_16107);
or U16184 (N_16184,N_16090,N_16088);
nor U16185 (N_16185,N_16073,N_16119);
nand U16186 (N_16186,N_16002,N_16030);
nor U16187 (N_16187,N_16019,N_16047);
and U16188 (N_16188,N_16137,N_16093);
or U16189 (N_16189,N_16118,N_16070);
or U16190 (N_16190,N_16052,N_16035);
nor U16191 (N_16191,N_16065,N_16034);
or U16192 (N_16192,N_16074,N_16102);
nor U16193 (N_16193,N_16127,N_16103);
nor U16194 (N_16194,N_16040,N_16066);
nand U16195 (N_16195,N_16036,N_16046);
and U16196 (N_16196,N_16078,N_16094);
nand U16197 (N_16197,N_16024,N_16135);
nand U16198 (N_16198,N_16143,N_16009);
or U16199 (N_16199,N_16081,N_16041);
and U16200 (N_16200,N_16147,N_16000);
and U16201 (N_16201,N_16124,N_16067);
or U16202 (N_16202,N_16012,N_16057);
xor U16203 (N_16203,N_16121,N_16087);
or U16204 (N_16204,N_16156,N_16068);
nor U16205 (N_16205,N_16048,N_16021);
nand U16206 (N_16206,N_16131,N_16063);
nor U16207 (N_16207,N_16159,N_16086);
or U16208 (N_16208,N_16060,N_16150);
and U16209 (N_16209,N_16108,N_16115);
and U16210 (N_16210,N_16140,N_16022);
or U16211 (N_16211,N_16080,N_16077);
and U16212 (N_16212,N_16069,N_16039);
xnor U16213 (N_16213,N_16157,N_16015);
xor U16214 (N_16214,N_16027,N_16112);
and U16215 (N_16215,N_16122,N_16059);
xnor U16216 (N_16216,N_16144,N_16051);
nor U16217 (N_16217,N_16029,N_16010);
or U16218 (N_16218,N_16020,N_16136);
xor U16219 (N_16219,N_16089,N_16128);
nor U16220 (N_16220,N_16105,N_16079);
or U16221 (N_16221,N_16114,N_16072);
xor U16222 (N_16222,N_16076,N_16018);
xor U16223 (N_16223,N_16075,N_16138);
xor U16224 (N_16224,N_16152,N_16158);
nor U16225 (N_16225,N_16095,N_16099);
xor U16226 (N_16226,N_16013,N_16053);
nand U16227 (N_16227,N_16082,N_16133);
nand U16228 (N_16228,N_16083,N_16008);
nor U16229 (N_16229,N_16084,N_16016);
nand U16230 (N_16230,N_16028,N_16050);
xor U16231 (N_16231,N_16071,N_16056);
nand U16232 (N_16232,N_16085,N_16014);
or U16233 (N_16233,N_16033,N_16151);
and U16234 (N_16234,N_16001,N_16038);
nand U16235 (N_16235,N_16023,N_16092);
xnor U16236 (N_16236,N_16129,N_16146);
nor U16237 (N_16237,N_16098,N_16043);
nand U16238 (N_16238,N_16007,N_16154);
xnor U16239 (N_16239,N_16058,N_16044);
nand U16240 (N_16240,N_16149,N_16050);
and U16241 (N_16241,N_16033,N_16041);
or U16242 (N_16242,N_16119,N_16051);
xnor U16243 (N_16243,N_16131,N_16106);
xnor U16244 (N_16244,N_16118,N_16018);
nand U16245 (N_16245,N_16037,N_16145);
or U16246 (N_16246,N_16105,N_16034);
or U16247 (N_16247,N_16048,N_16147);
nand U16248 (N_16248,N_16062,N_16001);
or U16249 (N_16249,N_16152,N_16054);
nand U16250 (N_16250,N_16024,N_16083);
nor U16251 (N_16251,N_16040,N_16104);
or U16252 (N_16252,N_16132,N_16156);
or U16253 (N_16253,N_16086,N_16003);
xnor U16254 (N_16254,N_16005,N_16025);
nor U16255 (N_16255,N_16102,N_16113);
or U16256 (N_16256,N_16144,N_16082);
nand U16257 (N_16257,N_16011,N_16079);
or U16258 (N_16258,N_16011,N_16146);
nor U16259 (N_16259,N_16119,N_16085);
nor U16260 (N_16260,N_16112,N_16147);
xor U16261 (N_16261,N_16101,N_16065);
nor U16262 (N_16262,N_16114,N_16151);
or U16263 (N_16263,N_16038,N_16128);
nand U16264 (N_16264,N_16081,N_16088);
or U16265 (N_16265,N_16085,N_16136);
nand U16266 (N_16266,N_16064,N_16026);
xor U16267 (N_16267,N_16084,N_16085);
or U16268 (N_16268,N_16102,N_16010);
and U16269 (N_16269,N_16029,N_16104);
and U16270 (N_16270,N_16072,N_16073);
and U16271 (N_16271,N_16022,N_16145);
xor U16272 (N_16272,N_16073,N_16155);
xnor U16273 (N_16273,N_16134,N_16143);
or U16274 (N_16274,N_16020,N_16018);
nand U16275 (N_16275,N_16014,N_16040);
xnor U16276 (N_16276,N_16020,N_16089);
nand U16277 (N_16277,N_16118,N_16126);
and U16278 (N_16278,N_16091,N_16093);
nor U16279 (N_16279,N_16123,N_16072);
or U16280 (N_16280,N_16060,N_16008);
nand U16281 (N_16281,N_16048,N_16023);
nor U16282 (N_16282,N_16051,N_16032);
nor U16283 (N_16283,N_16152,N_16027);
and U16284 (N_16284,N_16012,N_16103);
and U16285 (N_16285,N_16055,N_16084);
nand U16286 (N_16286,N_16009,N_16022);
and U16287 (N_16287,N_16080,N_16112);
xnor U16288 (N_16288,N_16064,N_16143);
nand U16289 (N_16289,N_16013,N_16006);
or U16290 (N_16290,N_16021,N_16111);
or U16291 (N_16291,N_16122,N_16146);
xor U16292 (N_16292,N_16105,N_16149);
nor U16293 (N_16293,N_16024,N_16055);
xor U16294 (N_16294,N_16100,N_16136);
xnor U16295 (N_16295,N_16114,N_16139);
nor U16296 (N_16296,N_16038,N_16017);
xor U16297 (N_16297,N_16110,N_16046);
nor U16298 (N_16298,N_16046,N_16130);
and U16299 (N_16299,N_16019,N_16104);
xnor U16300 (N_16300,N_16145,N_16026);
xnor U16301 (N_16301,N_16110,N_16013);
nor U16302 (N_16302,N_16138,N_16119);
and U16303 (N_16303,N_16066,N_16061);
and U16304 (N_16304,N_16138,N_16115);
or U16305 (N_16305,N_16073,N_16112);
nor U16306 (N_16306,N_16062,N_16036);
nand U16307 (N_16307,N_16139,N_16015);
or U16308 (N_16308,N_16071,N_16037);
or U16309 (N_16309,N_16033,N_16015);
xor U16310 (N_16310,N_16064,N_16108);
xnor U16311 (N_16311,N_16130,N_16089);
nor U16312 (N_16312,N_16118,N_16097);
nand U16313 (N_16313,N_16004,N_16037);
or U16314 (N_16314,N_16102,N_16122);
nand U16315 (N_16315,N_16088,N_16003);
nand U16316 (N_16316,N_16043,N_16118);
nor U16317 (N_16317,N_16125,N_16037);
and U16318 (N_16318,N_16100,N_16027);
nor U16319 (N_16319,N_16110,N_16095);
or U16320 (N_16320,N_16275,N_16271);
nand U16321 (N_16321,N_16302,N_16206);
nor U16322 (N_16322,N_16304,N_16284);
xnor U16323 (N_16323,N_16203,N_16283);
and U16324 (N_16324,N_16276,N_16255);
xor U16325 (N_16325,N_16211,N_16291);
nand U16326 (N_16326,N_16272,N_16162);
xnor U16327 (N_16327,N_16213,N_16306);
and U16328 (N_16328,N_16247,N_16278);
or U16329 (N_16329,N_16225,N_16189);
or U16330 (N_16330,N_16257,N_16200);
xnor U16331 (N_16331,N_16256,N_16232);
nor U16332 (N_16332,N_16303,N_16180);
and U16333 (N_16333,N_16201,N_16165);
xor U16334 (N_16334,N_16299,N_16172);
and U16335 (N_16335,N_16163,N_16166);
nor U16336 (N_16336,N_16215,N_16227);
nor U16337 (N_16337,N_16222,N_16171);
or U16338 (N_16338,N_16298,N_16263);
nor U16339 (N_16339,N_16252,N_16300);
xor U16340 (N_16340,N_16160,N_16168);
and U16341 (N_16341,N_16191,N_16216);
or U16342 (N_16342,N_16251,N_16223);
nor U16343 (N_16343,N_16226,N_16217);
nand U16344 (N_16344,N_16265,N_16179);
and U16345 (N_16345,N_16313,N_16293);
nand U16346 (N_16346,N_16267,N_16214);
or U16347 (N_16347,N_16254,N_16207);
nand U16348 (N_16348,N_16164,N_16229);
nand U16349 (N_16349,N_16309,N_16178);
xnor U16350 (N_16350,N_16301,N_16307);
or U16351 (N_16351,N_16228,N_16209);
or U16352 (N_16352,N_16192,N_16237);
nor U16353 (N_16353,N_16183,N_16246);
and U16354 (N_16354,N_16280,N_16249);
nand U16355 (N_16355,N_16208,N_16231);
or U16356 (N_16356,N_16314,N_16295);
nor U16357 (N_16357,N_16186,N_16234);
nor U16358 (N_16358,N_16188,N_16184);
xor U16359 (N_16359,N_16277,N_16285);
and U16360 (N_16360,N_16290,N_16242);
xor U16361 (N_16361,N_16243,N_16253);
xnor U16362 (N_16362,N_16196,N_16266);
nand U16363 (N_16363,N_16269,N_16289);
nand U16364 (N_16364,N_16182,N_16170);
nand U16365 (N_16365,N_16230,N_16194);
or U16366 (N_16366,N_16238,N_16250);
xor U16367 (N_16367,N_16296,N_16187);
xor U16368 (N_16368,N_16308,N_16286);
nor U16369 (N_16369,N_16316,N_16236);
xor U16370 (N_16370,N_16297,N_16173);
or U16371 (N_16371,N_16212,N_16161);
or U16372 (N_16372,N_16220,N_16260);
nor U16373 (N_16373,N_16241,N_16202);
nand U16374 (N_16374,N_16198,N_16315);
and U16375 (N_16375,N_16292,N_16261);
and U16376 (N_16376,N_16244,N_16305);
xor U16377 (N_16377,N_16245,N_16270);
xor U16378 (N_16378,N_16259,N_16240);
xor U16379 (N_16379,N_16205,N_16281);
nor U16380 (N_16380,N_16177,N_16185);
and U16381 (N_16381,N_16175,N_16319);
and U16382 (N_16382,N_16167,N_16233);
nor U16383 (N_16383,N_16204,N_16310);
and U16384 (N_16384,N_16311,N_16218);
and U16385 (N_16385,N_16268,N_16181);
and U16386 (N_16386,N_16288,N_16239);
and U16387 (N_16387,N_16224,N_16190);
xnor U16388 (N_16388,N_16248,N_16193);
or U16389 (N_16389,N_16235,N_16199);
nor U16390 (N_16390,N_16176,N_16312);
xor U16391 (N_16391,N_16210,N_16195);
or U16392 (N_16392,N_16258,N_16264);
nand U16393 (N_16393,N_16273,N_16287);
nand U16394 (N_16394,N_16169,N_16282);
nand U16395 (N_16395,N_16318,N_16221);
or U16396 (N_16396,N_16219,N_16294);
and U16397 (N_16397,N_16274,N_16262);
nor U16398 (N_16398,N_16279,N_16174);
and U16399 (N_16399,N_16197,N_16317);
and U16400 (N_16400,N_16301,N_16206);
xor U16401 (N_16401,N_16222,N_16184);
or U16402 (N_16402,N_16234,N_16167);
nand U16403 (N_16403,N_16182,N_16263);
nand U16404 (N_16404,N_16212,N_16246);
or U16405 (N_16405,N_16239,N_16264);
xor U16406 (N_16406,N_16278,N_16234);
xor U16407 (N_16407,N_16175,N_16290);
xor U16408 (N_16408,N_16287,N_16167);
or U16409 (N_16409,N_16262,N_16220);
xnor U16410 (N_16410,N_16243,N_16319);
nor U16411 (N_16411,N_16221,N_16259);
nor U16412 (N_16412,N_16174,N_16230);
nor U16413 (N_16413,N_16210,N_16221);
and U16414 (N_16414,N_16192,N_16161);
or U16415 (N_16415,N_16312,N_16264);
nand U16416 (N_16416,N_16298,N_16174);
nor U16417 (N_16417,N_16221,N_16232);
or U16418 (N_16418,N_16271,N_16191);
xnor U16419 (N_16419,N_16292,N_16240);
nor U16420 (N_16420,N_16235,N_16273);
nor U16421 (N_16421,N_16304,N_16279);
nand U16422 (N_16422,N_16204,N_16245);
or U16423 (N_16423,N_16173,N_16255);
xor U16424 (N_16424,N_16265,N_16308);
nor U16425 (N_16425,N_16200,N_16260);
xor U16426 (N_16426,N_16218,N_16304);
nor U16427 (N_16427,N_16231,N_16271);
xnor U16428 (N_16428,N_16185,N_16166);
xor U16429 (N_16429,N_16272,N_16264);
xnor U16430 (N_16430,N_16194,N_16283);
xnor U16431 (N_16431,N_16162,N_16257);
or U16432 (N_16432,N_16233,N_16261);
nand U16433 (N_16433,N_16216,N_16308);
nor U16434 (N_16434,N_16173,N_16243);
or U16435 (N_16435,N_16265,N_16228);
nand U16436 (N_16436,N_16239,N_16259);
nor U16437 (N_16437,N_16312,N_16234);
nor U16438 (N_16438,N_16274,N_16210);
or U16439 (N_16439,N_16259,N_16255);
nor U16440 (N_16440,N_16218,N_16295);
and U16441 (N_16441,N_16172,N_16317);
and U16442 (N_16442,N_16171,N_16312);
and U16443 (N_16443,N_16198,N_16307);
nor U16444 (N_16444,N_16164,N_16278);
or U16445 (N_16445,N_16279,N_16295);
nand U16446 (N_16446,N_16292,N_16241);
nor U16447 (N_16447,N_16289,N_16245);
and U16448 (N_16448,N_16195,N_16256);
xor U16449 (N_16449,N_16197,N_16161);
and U16450 (N_16450,N_16186,N_16213);
xor U16451 (N_16451,N_16287,N_16304);
xor U16452 (N_16452,N_16196,N_16230);
nor U16453 (N_16453,N_16257,N_16219);
xor U16454 (N_16454,N_16173,N_16224);
nand U16455 (N_16455,N_16236,N_16319);
or U16456 (N_16456,N_16229,N_16213);
nor U16457 (N_16457,N_16222,N_16223);
and U16458 (N_16458,N_16244,N_16307);
nor U16459 (N_16459,N_16267,N_16211);
nor U16460 (N_16460,N_16259,N_16266);
xor U16461 (N_16461,N_16184,N_16286);
or U16462 (N_16462,N_16268,N_16309);
or U16463 (N_16463,N_16212,N_16318);
and U16464 (N_16464,N_16239,N_16297);
or U16465 (N_16465,N_16236,N_16238);
nor U16466 (N_16466,N_16239,N_16302);
and U16467 (N_16467,N_16278,N_16207);
nand U16468 (N_16468,N_16295,N_16219);
and U16469 (N_16469,N_16196,N_16253);
or U16470 (N_16470,N_16307,N_16201);
or U16471 (N_16471,N_16278,N_16290);
or U16472 (N_16472,N_16230,N_16304);
xor U16473 (N_16473,N_16225,N_16224);
and U16474 (N_16474,N_16182,N_16186);
nor U16475 (N_16475,N_16256,N_16160);
or U16476 (N_16476,N_16180,N_16205);
xnor U16477 (N_16477,N_16283,N_16191);
nor U16478 (N_16478,N_16199,N_16168);
nand U16479 (N_16479,N_16313,N_16193);
nor U16480 (N_16480,N_16414,N_16419);
xor U16481 (N_16481,N_16346,N_16468);
xor U16482 (N_16482,N_16398,N_16384);
xor U16483 (N_16483,N_16442,N_16458);
xnor U16484 (N_16484,N_16401,N_16351);
nand U16485 (N_16485,N_16392,N_16465);
nor U16486 (N_16486,N_16444,N_16412);
nor U16487 (N_16487,N_16329,N_16336);
or U16488 (N_16488,N_16344,N_16467);
nand U16489 (N_16489,N_16323,N_16477);
or U16490 (N_16490,N_16441,N_16461);
xnor U16491 (N_16491,N_16437,N_16368);
nand U16492 (N_16492,N_16418,N_16469);
nand U16493 (N_16493,N_16434,N_16420);
and U16494 (N_16494,N_16352,N_16358);
nor U16495 (N_16495,N_16416,N_16411);
nor U16496 (N_16496,N_16391,N_16429);
and U16497 (N_16497,N_16472,N_16369);
nand U16498 (N_16498,N_16359,N_16386);
and U16499 (N_16499,N_16473,N_16470);
nor U16500 (N_16500,N_16342,N_16403);
nand U16501 (N_16501,N_16340,N_16337);
xnor U16502 (N_16502,N_16479,N_16453);
xor U16503 (N_16503,N_16387,N_16376);
or U16504 (N_16504,N_16390,N_16393);
and U16505 (N_16505,N_16460,N_16354);
or U16506 (N_16506,N_16396,N_16360);
xor U16507 (N_16507,N_16327,N_16424);
or U16508 (N_16508,N_16413,N_16348);
or U16509 (N_16509,N_16421,N_16400);
nand U16510 (N_16510,N_16372,N_16328);
nand U16511 (N_16511,N_16422,N_16406);
nand U16512 (N_16512,N_16474,N_16435);
or U16513 (N_16513,N_16395,N_16456);
xnor U16514 (N_16514,N_16431,N_16380);
nand U16515 (N_16515,N_16432,N_16321);
nor U16516 (N_16516,N_16408,N_16404);
nand U16517 (N_16517,N_16343,N_16320);
and U16518 (N_16518,N_16450,N_16448);
nor U16519 (N_16519,N_16379,N_16367);
or U16520 (N_16520,N_16333,N_16402);
nor U16521 (N_16521,N_16375,N_16425);
and U16522 (N_16522,N_16370,N_16356);
or U16523 (N_16523,N_16399,N_16363);
nor U16524 (N_16524,N_16455,N_16326);
nor U16525 (N_16525,N_16454,N_16427);
nand U16526 (N_16526,N_16322,N_16471);
or U16527 (N_16527,N_16364,N_16332);
xnor U16528 (N_16528,N_16353,N_16371);
and U16529 (N_16529,N_16410,N_16409);
and U16530 (N_16530,N_16407,N_16443);
xor U16531 (N_16531,N_16451,N_16362);
nor U16532 (N_16532,N_16325,N_16378);
nor U16533 (N_16533,N_16436,N_16335);
and U16534 (N_16534,N_16373,N_16339);
nand U16535 (N_16535,N_16382,N_16440);
or U16536 (N_16536,N_16405,N_16446);
nand U16537 (N_16537,N_16345,N_16430);
and U16538 (N_16538,N_16383,N_16463);
nor U16539 (N_16539,N_16350,N_16445);
xnor U16540 (N_16540,N_16417,N_16457);
and U16541 (N_16541,N_16426,N_16449);
nand U16542 (N_16542,N_16452,N_16347);
and U16543 (N_16543,N_16365,N_16478);
xor U16544 (N_16544,N_16388,N_16464);
nand U16545 (N_16545,N_16331,N_16381);
nor U16546 (N_16546,N_16428,N_16459);
nor U16547 (N_16547,N_16466,N_16476);
xor U16548 (N_16548,N_16341,N_16397);
xor U16549 (N_16549,N_16366,N_16415);
or U16550 (N_16550,N_16433,N_16377);
or U16551 (N_16551,N_16374,N_16385);
nand U16552 (N_16552,N_16438,N_16389);
nand U16553 (N_16553,N_16394,N_16357);
nor U16554 (N_16554,N_16324,N_16361);
or U16555 (N_16555,N_16330,N_16349);
or U16556 (N_16556,N_16475,N_16447);
or U16557 (N_16557,N_16462,N_16439);
nand U16558 (N_16558,N_16334,N_16355);
nor U16559 (N_16559,N_16423,N_16338);
nand U16560 (N_16560,N_16327,N_16354);
nand U16561 (N_16561,N_16335,N_16412);
nand U16562 (N_16562,N_16471,N_16395);
nor U16563 (N_16563,N_16338,N_16327);
nor U16564 (N_16564,N_16336,N_16434);
and U16565 (N_16565,N_16426,N_16340);
xor U16566 (N_16566,N_16379,N_16370);
nand U16567 (N_16567,N_16369,N_16389);
nor U16568 (N_16568,N_16436,N_16386);
nor U16569 (N_16569,N_16353,N_16320);
nor U16570 (N_16570,N_16349,N_16407);
and U16571 (N_16571,N_16435,N_16337);
xor U16572 (N_16572,N_16417,N_16428);
or U16573 (N_16573,N_16402,N_16476);
nand U16574 (N_16574,N_16323,N_16454);
xor U16575 (N_16575,N_16432,N_16459);
nand U16576 (N_16576,N_16470,N_16379);
nand U16577 (N_16577,N_16381,N_16444);
and U16578 (N_16578,N_16323,N_16431);
nand U16579 (N_16579,N_16440,N_16360);
nand U16580 (N_16580,N_16337,N_16379);
and U16581 (N_16581,N_16468,N_16367);
or U16582 (N_16582,N_16320,N_16442);
nor U16583 (N_16583,N_16366,N_16378);
and U16584 (N_16584,N_16377,N_16341);
and U16585 (N_16585,N_16361,N_16446);
nor U16586 (N_16586,N_16464,N_16339);
or U16587 (N_16587,N_16384,N_16443);
nor U16588 (N_16588,N_16329,N_16403);
nor U16589 (N_16589,N_16419,N_16406);
nor U16590 (N_16590,N_16416,N_16355);
nor U16591 (N_16591,N_16385,N_16398);
nor U16592 (N_16592,N_16352,N_16467);
or U16593 (N_16593,N_16430,N_16364);
nor U16594 (N_16594,N_16446,N_16345);
and U16595 (N_16595,N_16394,N_16418);
xor U16596 (N_16596,N_16358,N_16325);
nor U16597 (N_16597,N_16346,N_16371);
or U16598 (N_16598,N_16395,N_16389);
nand U16599 (N_16599,N_16371,N_16375);
nor U16600 (N_16600,N_16340,N_16359);
nand U16601 (N_16601,N_16326,N_16343);
nor U16602 (N_16602,N_16370,N_16382);
or U16603 (N_16603,N_16389,N_16474);
nand U16604 (N_16604,N_16343,N_16408);
nand U16605 (N_16605,N_16382,N_16407);
xor U16606 (N_16606,N_16331,N_16354);
and U16607 (N_16607,N_16354,N_16407);
nor U16608 (N_16608,N_16455,N_16366);
and U16609 (N_16609,N_16460,N_16425);
nor U16610 (N_16610,N_16358,N_16408);
or U16611 (N_16611,N_16389,N_16383);
xnor U16612 (N_16612,N_16414,N_16330);
and U16613 (N_16613,N_16350,N_16345);
nor U16614 (N_16614,N_16447,N_16456);
or U16615 (N_16615,N_16322,N_16400);
nor U16616 (N_16616,N_16476,N_16329);
xor U16617 (N_16617,N_16369,N_16457);
and U16618 (N_16618,N_16344,N_16455);
nor U16619 (N_16619,N_16442,N_16474);
and U16620 (N_16620,N_16402,N_16331);
or U16621 (N_16621,N_16336,N_16347);
and U16622 (N_16622,N_16439,N_16417);
or U16623 (N_16623,N_16386,N_16470);
and U16624 (N_16624,N_16427,N_16469);
xor U16625 (N_16625,N_16371,N_16401);
nor U16626 (N_16626,N_16347,N_16409);
xnor U16627 (N_16627,N_16437,N_16479);
nand U16628 (N_16628,N_16337,N_16351);
xnor U16629 (N_16629,N_16404,N_16320);
xnor U16630 (N_16630,N_16449,N_16399);
nand U16631 (N_16631,N_16343,N_16459);
xnor U16632 (N_16632,N_16369,N_16320);
nand U16633 (N_16633,N_16381,N_16404);
or U16634 (N_16634,N_16359,N_16389);
nor U16635 (N_16635,N_16435,N_16454);
nand U16636 (N_16636,N_16334,N_16353);
nand U16637 (N_16637,N_16417,N_16424);
nand U16638 (N_16638,N_16375,N_16474);
nand U16639 (N_16639,N_16431,N_16342);
xor U16640 (N_16640,N_16485,N_16520);
nor U16641 (N_16641,N_16512,N_16494);
nand U16642 (N_16642,N_16600,N_16539);
and U16643 (N_16643,N_16558,N_16622);
and U16644 (N_16644,N_16594,N_16636);
nor U16645 (N_16645,N_16639,N_16580);
and U16646 (N_16646,N_16583,N_16486);
nor U16647 (N_16647,N_16569,N_16595);
xnor U16648 (N_16648,N_16586,N_16553);
and U16649 (N_16649,N_16633,N_16524);
nor U16650 (N_16650,N_16533,N_16502);
and U16651 (N_16651,N_16566,N_16489);
nor U16652 (N_16652,N_16621,N_16599);
nor U16653 (N_16653,N_16625,N_16577);
or U16654 (N_16654,N_16634,N_16560);
and U16655 (N_16655,N_16611,N_16536);
xnor U16656 (N_16656,N_16574,N_16513);
xnor U16657 (N_16657,N_16523,N_16589);
nor U16658 (N_16658,N_16525,N_16497);
xor U16659 (N_16659,N_16587,N_16554);
xnor U16660 (N_16660,N_16635,N_16534);
nor U16661 (N_16661,N_16638,N_16607);
xor U16662 (N_16662,N_16627,N_16527);
nand U16663 (N_16663,N_16612,N_16631);
or U16664 (N_16664,N_16484,N_16608);
nand U16665 (N_16665,N_16591,N_16537);
nor U16666 (N_16666,N_16480,N_16542);
xor U16667 (N_16667,N_16528,N_16543);
nor U16668 (N_16668,N_16482,N_16596);
nor U16669 (N_16669,N_16511,N_16481);
or U16670 (N_16670,N_16624,N_16550);
and U16671 (N_16671,N_16610,N_16617);
xnor U16672 (N_16672,N_16615,N_16575);
or U16673 (N_16673,N_16491,N_16496);
xnor U16674 (N_16674,N_16620,N_16637);
nor U16675 (N_16675,N_16571,N_16565);
nor U16676 (N_16676,N_16592,N_16499);
nor U16677 (N_16677,N_16570,N_16555);
nand U16678 (N_16678,N_16604,N_16582);
nor U16679 (N_16679,N_16593,N_16544);
xor U16680 (N_16680,N_16613,N_16492);
nor U16681 (N_16681,N_16585,N_16584);
and U16682 (N_16682,N_16606,N_16629);
nor U16683 (N_16683,N_16602,N_16517);
xnor U16684 (N_16684,N_16626,N_16614);
xor U16685 (N_16685,N_16632,N_16628);
xor U16686 (N_16686,N_16532,N_16573);
or U16687 (N_16687,N_16568,N_16531);
xnor U16688 (N_16688,N_16609,N_16619);
nand U16689 (N_16689,N_16488,N_16526);
nand U16690 (N_16690,N_16588,N_16540);
and U16691 (N_16691,N_16530,N_16509);
nand U16692 (N_16692,N_16547,N_16549);
or U16693 (N_16693,N_16493,N_16598);
xor U16694 (N_16694,N_16559,N_16490);
nand U16695 (N_16695,N_16501,N_16630);
or U16696 (N_16696,N_16576,N_16519);
and U16697 (N_16697,N_16529,N_16500);
nand U16698 (N_16698,N_16605,N_16510);
nand U16699 (N_16699,N_16507,N_16579);
nand U16700 (N_16700,N_16538,N_16572);
and U16701 (N_16701,N_16521,N_16522);
and U16702 (N_16702,N_16562,N_16495);
xor U16703 (N_16703,N_16546,N_16557);
nand U16704 (N_16704,N_16548,N_16487);
or U16705 (N_16705,N_16590,N_16618);
or U16706 (N_16706,N_16616,N_16561);
or U16707 (N_16707,N_16503,N_16603);
or U16708 (N_16708,N_16563,N_16498);
nor U16709 (N_16709,N_16514,N_16505);
or U16710 (N_16710,N_16567,N_16601);
or U16711 (N_16711,N_16508,N_16504);
or U16712 (N_16712,N_16545,N_16515);
nand U16713 (N_16713,N_16541,N_16551);
nor U16714 (N_16714,N_16483,N_16597);
or U16715 (N_16715,N_16623,N_16516);
and U16716 (N_16716,N_16506,N_16556);
nand U16717 (N_16717,N_16564,N_16581);
xor U16718 (N_16718,N_16535,N_16578);
and U16719 (N_16719,N_16552,N_16518);
and U16720 (N_16720,N_16619,N_16574);
nand U16721 (N_16721,N_16551,N_16484);
nand U16722 (N_16722,N_16604,N_16481);
or U16723 (N_16723,N_16506,N_16638);
nand U16724 (N_16724,N_16508,N_16623);
and U16725 (N_16725,N_16615,N_16639);
nor U16726 (N_16726,N_16550,N_16601);
xor U16727 (N_16727,N_16560,N_16495);
or U16728 (N_16728,N_16553,N_16526);
xnor U16729 (N_16729,N_16499,N_16504);
xor U16730 (N_16730,N_16611,N_16599);
and U16731 (N_16731,N_16568,N_16532);
or U16732 (N_16732,N_16524,N_16609);
xor U16733 (N_16733,N_16568,N_16623);
nand U16734 (N_16734,N_16551,N_16540);
and U16735 (N_16735,N_16574,N_16506);
or U16736 (N_16736,N_16551,N_16570);
nand U16737 (N_16737,N_16594,N_16634);
xor U16738 (N_16738,N_16542,N_16571);
and U16739 (N_16739,N_16496,N_16590);
and U16740 (N_16740,N_16569,N_16480);
and U16741 (N_16741,N_16517,N_16491);
or U16742 (N_16742,N_16560,N_16602);
or U16743 (N_16743,N_16496,N_16555);
xor U16744 (N_16744,N_16484,N_16556);
nand U16745 (N_16745,N_16582,N_16533);
and U16746 (N_16746,N_16488,N_16567);
xnor U16747 (N_16747,N_16621,N_16540);
or U16748 (N_16748,N_16502,N_16629);
and U16749 (N_16749,N_16505,N_16637);
or U16750 (N_16750,N_16576,N_16543);
xor U16751 (N_16751,N_16493,N_16519);
or U16752 (N_16752,N_16611,N_16485);
and U16753 (N_16753,N_16531,N_16544);
nor U16754 (N_16754,N_16567,N_16515);
or U16755 (N_16755,N_16605,N_16609);
and U16756 (N_16756,N_16501,N_16574);
or U16757 (N_16757,N_16581,N_16505);
nor U16758 (N_16758,N_16486,N_16576);
nand U16759 (N_16759,N_16599,N_16623);
nor U16760 (N_16760,N_16511,N_16598);
nor U16761 (N_16761,N_16561,N_16527);
nand U16762 (N_16762,N_16595,N_16584);
or U16763 (N_16763,N_16627,N_16538);
or U16764 (N_16764,N_16603,N_16566);
nor U16765 (N_16765,N_16508,N_16601);
nor U16766 (N_16766,N_16638,N_16494);
and U16767 (N_16767,N_16514,N_16491);
and U16768 (N_16768,N_16632,N_16531);
xnor U16769 (N_16769,N_16561,N_16517);
or U16770 (N_16770,N_16606,N_16635);
nand U16771 (N_16771,N_16558,N_16542);
and U16772 (N_16772,N_16579,N_16587);
or U16773 (N_16773,N_16492,N_16497);
nand U16774 (N_16774,N_16603,N_16480);
nand U16775 (N_16775,N_16594,N_16592);
xnor U16776 (N_16776,N_16635,N_16494);
nor U16777 (N_16777,N_16614,N_16631);
nand U16778 (N_16778,N_16625,N_16605);
nor U16779 (N_16779,N_16614,N_16495);
nor U16780 (N_16780,N_16564,N_16484);
nand U16781 (N_16781,N_16489,N_16574);
and U16782 (N_16782,N_16505,N_16533);
xnor U16783 (N_16783,N_16581,N_16603);
nand U16784 (N_16784,N_16556,N_16534);
and U16785 (N_16785,N_16491,N_16615);
xnor U16786 (N_16786,N_16525,N_16577);
or U16787 (N_16787,N_16585,N_16601);
xor U16788 (N_16788,N_16481,N_16600);
nor U16789 (N_16789,N_16563,N_16521);
and U16790 (N_16790,N_16486,N_16549);
xor U16791 (N_16791,N_16496,N_16580);
xor U16792 (N_16792,N_16588,N_16596);
nand U16793 (N_16793,N_16619,N_16537);
nor U16794 (N_16794,N_16560,N_16543);
or U16795 (N_16795,N_16598,N_16585);
and U16796 (N_16796,N_16581,N_16550);
or U16797 (N_16797,N_16547,N_16509);
and U16798 (N_16798,N_16545,N_16519);
nand U16799 (N_16799,N_16530,N_16569);
nor U16800 (N_16800,N_16690,N_16784);
nand U16801 (N_16801,N_16736,N_16687);
nand U16802 (N_16802,N_16716,N_16792);
nor U16803 (N_16803,N_16649,N_16785);
and U16804 (N_16804,N_16659,N_16799);
nor U16805 (N_16805,N_16730,N_16791);
nor U16806 (N_16806,N_16654,N_16775);
and U16807 (N_16807,N_16697,N_16702);
xnor U16808 (N_16808,N_16797,N_16780);
xor U16809 (N_16809,N_16725,N_16684);
xor U16810 (N_16810,N_16679,N_16790);
xnor U16811 (N_16811,N_16676,N_16650);
nor U16812 (N_16812,N_16720,N_16642);
nor U16813 (N_16813,N_16652,N_16743);
nand U16814 (N_16814,N_16680,N_16745);
nand U16815 (N_16815,N_16750,N_16671);
nor U16816 (N_16816,N_16645,N_16749);
xor U16817 (N_16817,N_16708,N_16701);
and U16818 (N_16818,N_16757,N_16640);
xor U16819 (N_16819,N_16779,N_16648);
nor U16820 (N_16820,N_16758,N_16794);
and U16821 (N_16821,N_16657,N_16741);
xnor U16822 (N_16822,N_16713,N_16728);
nor U16823 (N_16823,N_16686,N_16718);
xor U16824 (N_16824,N_16696,N_16773);
and U16825 (N_16825,N_16769,N_16783);
nor U16826 (N_16826,N_16665,N_16703);
nand U16827 (N_16827,N_16664,N_16770);
and U16828 (N_16828,N_16755,N_16709);
and U16829 (N_16829,N_16672,N_16647);
nor U16830 (N_16830,N_16742,N_16729);
nand U16831 (N_16831,N_16681,N_16691);
and U16832 (N_16832,N_16643,N_16724);
nand U16833 (N_16833,N_16712,N_16767);
or U16834 (N_16834,N_16731,N_16752);
xor U16835 (N_16835,N_16727,N_16719);
nor U16836 (N_16836,N_16644,N_16695);
and U16837 (N_16837,N_16683,N_16768);
nor U16838 (N_16838,N_16692,N_16641);
nand U16839 (N_16839,N_16698,N_16760);
nand U16840 (N_16840,N_16756,N_16667);
or U16841 (N_16841,N_16782,N_16722);
nand U16842 (N_16842,N_16796,N_16748);
and U16843 (N_16843,N_16653,N_16663);
nand U16844 (N_16844,N_16735,N_16711);
xor U16845 (N_16845,N_16738,N_16776);
nor U16846 (N_16846,N_16798,N_16688);
and U16847 (N_16847,N_16732,N_16733);
and U16848 (N_16848,N_16693,N_16694);
xnor U16849 (N_16849,N_16658,N_16740);
xnor U16850 (N_16850,N_16789,N_16781);
and U16851 (N_16851,N_16706,N_16766);
and U16852 (N_16852,N_16714,N_16751);
and U16853 (N_16853,N_16739,N_16771);
or U16854 (N_16854,N_16700,N_16705);
nor U16855 (N_16855,N_16682,N_16677);
nand U16856 (N_16856,N_16675,N_16759);
or U16857 (N_16857,N_16710,N_16737);
xnor U16858 (N_16858,N_16717,N_16673);
nand U16859 (N_16859,N_16746,N_16772);
and U16860 (N_16860,N_16761,N_16656);
nand U16861 (N_16861,N_16753,N_16668);
or U16862 (N_16862,N_16669,N_16786);
xor U16863 (N_16863,N_16674,N_16747);
nand U16864 (N_16864,N_16707,N_16726);
and U16865 (N_16865,N_16723,N_16670);
nand U16866 (N_16866,N_16765,N_16788);
or U16867 (N_16867,N_16685,N_16763);
nand U16868 (N_16868,N_16699,N_16704);
nor U16869 (N_16869,N_16678,N_16689);
xor U16870 (N_16870,N_16651,N_16661);
and U16871 (N_16871,N_16744,N_16655);
nand U16872 (N_16872,N_16778,N_16666);
nand U16873 (N_16873,N_16764,N_16795);
nand U16874 (N_16874,N_16715,N_16793);
or U16875 (N_16875,N_16777,N_16762);
xnor U16876 (N_16876,N_16754,N_16646);
or U16877 (N_16877,N_16787,N_16774);
and U16878 (N_16878,N_16734,N_16660);
and U16879 (N_16879,N_16662,N_16721);
and U16880 (N_16880,N_16694,N_16771);
nor U16881 (N_16881,N_16719,N_16655);
nor U16882 (N_16882,N_16702,N_16681);
or U16883 (N_16883,N_16647,N_16726);
xnor U16884 (N_16884,N_16684,N_16750);
xor U16885 (N_16885,N_16725,N_16783);
and U16886 (N_16886,N_16665,N_16670);
xor U16887 (N_16887,N_16795,N_16697);
or U16888 (N_16888,N_16715,N_16664);
and U16889 (N_16889,N_16666,N_16703);
and U16890 (N_16890,N_16793,N_16791);
or U16891 (N_16891,N_16650,N_16754);
nand U16892 (N_16892,N_16789,N_16696);
and U16893 (N_16893,N_16683,N_16640);
nand U16894 (N_16894,N_16676,N_16778);
xor U16895 (N_16895,N_16759,N_16672);
xnor U16896 (N_16896,N_16774,N_16674);
and U16897 (N_16897,N_16741,N_16791);
and U16898 (N_16898,N_16704,N_16701);
nor U16899 (N_16899,N_16798,N_16785);
and U16900 (N_16900,N_16673,N_16788);
or U16901 (N_16901,N_16780,N_16676);
nor U16902 (N_16902,N_16789,N_16764);
and U16903 (N_16903,N_16770,N_16672);
nor U16904 (N_16904,N_16671,N_16704);
and U16905 (N_16905,N_16776,N_16763);
or U16906 (N_16906,N_16703,N_16671);
xnor U16907 (N_16907,N_16786,N_16727);
or U16908 (N_16908,N_16655,N_16664);
and U16909 (N_16909,N_16769,N_16743);
nor U16910 (N_16910,N_16686,N_16692);
and U16911 (N_16911,N_16728,N_16708);
nand U16912 (N_16912,N_16733,N_16755);
or U16913 (N_16913,N_16712,N_16652);
nand U16914 (N_16914,N_16773,N_16689);
or U16915 (N_16915,N_16763,N_16728);
nor U16916 (N_16916,N_16694,N_16658);
and U16917 (N_16917,N_16740,N_16707);
and U16918 (N_16918,N_16653,N_16756);
or U16919 (N_16919,N_16728,N_16795);
xnor U16920 (N_16920,N_16655,N_16773);
and U16921 (N_16921,N_16701,N_16782);
nor U16922 (N_16922,N_16672,N_16643);
and U16923 (N_16923,N_16757,N_16760);
and U16924 (N_16924,N_16703,N_16754);
nor U16925 (N_16925,N_16785,N_16723);
and U16926 (N_16926,N_16775,N_16761);
xor U16927 (N_16927,N_16680,N_16678);
and U16928 (N_16928,N_16772,N_16776);
or U16929 (N_16929,N_16733,N_16727);
xor U16930 (N_16930,N_16762,N_16686);
and U16931 (N_16931,N_16719,N_16671);
or U16932 (N_16932,N_16773,N_16720);
xnor U16933 (N_16933,N_16781,N_16793);
xor U16934 (N_16934,N_16791,N_16654);
nor U16935 (N_16935,N_16787,N_16798);
and U16936 (N_16936,N_16691,N_16709);
xnor U16937 (N_16937,N_16743,N_16724);
nor U16938 (N_16938,N_16652,N_16651);
nor U16939 (N_16939,N_16784,N_16665);
xor U16940 (N_16940,N_16646,N_16660);
or U16941 (N_16941,N_16665,N_16640);
xor U16942 (N_16942,N_16650,N_16768);
nand U16943 (N_16943,N_16697,N_16771);
xor U16944 (N_16944,N_16780,N_16765);
and U16945 (N_16945,N_16686,N_16797);
nand U16946 (N_16946,N_16753,N_16696);
and U16947 (N_16947,N_16681,N_16676);
xnor U16948 (N_16948,N_16691,N_16751);
xnor U16949 (N_16949,N_16708,N_16661);
nor U16950 (N_16950,N_16686,N_16646);
xor U16951 (N_16951,N_16655,N_16721);
nor U16952 (N_16952,N_16742,N_16725);
nand U16953 (N_16953,N_16780,N_16655);
nand U16954 (N_16954,N_16773,N_16735);
nor U16955 (N_16955,N_16692,N_16684);
and U16956 (N_16956,N_16753,N_16752);
or U16957 (N_16957,N_16656,N_16671);
nor U16958 (N_16958,N_16764,N_16750);
xnor U16959 (N_16959,N_16753,N_16689);
xnor U16960 (N_16960,N_16945,N_16800);
nor U16961 (N_16961,N_16846,N_16832);
nand U16962 (N_16962,N_16817,N_16835);
and U16963 (N_16963,N_16857,N_16901);
xnor U16964 (N_16964,N_16931,N_16896);
nand U16965 (N_16965,N_16819,N_16871);
nor U16966 (N_16966,N_16954,N_16828);
and U16967 (N_16967,N_16868,N_16842);
nand U16968 (N_16968,N_16886,N_16893);
nor U16969 (N_16969,N_16877,N_16863);
and U16970 (N_16970,N_16940,N_16939);
nor U16971 (N_16971,N_16908,N_16823);
xor U16972 (N_16972,N_16865,N_16906);
and U16973 (N_16973,N_16949,N_16873);
xnor U16974 (N_16974,N_16820,N_16809);
xor U16975 (N_16975,N_16938,N_16920);
nor U16976 (N_16976,N_16933,N_16900);
and U16977 (N_16977,N_16850,N_16838);
and U16978 (N_16978,N_16891,N_16904);
nor U16979 (N_16979,N_16903,N_16811);
and U16980 (N_16980,N_16959,N_16834);
xnor U16981 (N_16981,N_16887,N_16824);
xnor U16982 (N_16982,N_16801,N_16951);
nor U16983 (N_16983,N_16888,N_16956);
or U16984 (N_16984,N_16909,N_16924);
nand U16985 (N_16985,N_16937,N_16827);
xor U16986 (N_16986,N_16874,N_16936);
nand U16987 (N_16987,N_16875,N_16853);
and U16988 (N_16988,N_16890,N_16905);
xor U16989 (N_16989,N_16913,N_16812);
nand U16990 (N_16990,N_16855,N_16942);
xnor U16991 (N_16991,N_16944,N_16870);
and U16992 (N_16992,N_16805,N_16833);
nand U16993 (N_16993,N_16957,N_16895);
nand U16994 (N_16994,N_16911,N_16930);
xnor U16995 (N_16995,N_16818,N_16837);
nor U16996 (N_16996,N_16815,N_16892);
nand U16997 (N_16997,N_16826,N_16862);
xor U16998 (N_16998,N_16860,N_16907);
nand U16999 (N_16999,N_16808,N_16854);
xor U17000 (N_17000,N_16867,N_16915);
nand U17001 (N_17001,N_16810,N_16946);
and U17002 (N_17002,N_16921,N_16925);
nand U17003 (N_17003,N_16883,N_16852);
nor U17004 (N_17004,N_16884,N_16861);
xor U17005 (N_17005,N_16918,N_16847);
and U17006 (N_17006,N_16950,N_16881);
nand U17007 (N_17007,N_16864,N_16929);
xnor U17008 (N_17008,N_16914,N_16858);
or U17009 (N_17009,N_16821,N_16848);
xnor U17010 (N_17010,N_16917,N_16947);
or U17011 (N_17011,N_16841,N_16804);
and U17012 (N_17012,N_16845,N_16912);
nand U17013 (N_17013,N_16916,N_16807);
nand U17014 (N_17014,N_16849,N_16953);
or U17015 (N_17015,N_16843,N_16803);
nor U17016 (N_17016,N_16941,N_16813);
and U17017 (N_17017,N_16898,N_16923);
nand U17018 (N_17018,N_16928,N_16816);
nor U17019 (N_17019,N_16866,N_16844);
and U17020 (N_17020,N_16948,N_16943);
nand U17021 (N_17021,N_16831,N_16856);
or U17022 (N_17022,N_16955,N_16910);
or U17023 (N_17023,N_16919,N_16840);
nand U17024 (N_17024,N_16859,N_16878);
nand U17025 (N_17025,N_16932,N_16889);
nor U17026 (N_17026,N_16927,N_16876);
and U17027 (N_17027,N_16926,N_16869);
nand U17028 (N_17028,N_16839,N_16952);
xnor U17029 (N_17029,N_16802,N_16851);
nor U17030 (N_17030,N_16958,N_16872);
nand U17031 (N_17031,N_16830,N_16829);
xnor U17032 (N_17032,N_16822,N_16902);
nand U17033 (N_17033,N_16814,N_16897);
nor U17034 (N_17034,N_16899,N_16879);
nor U17035 (N_17035,N_16894,N_16885);
or U17036 (N_17036,N_16934,N_16935);
xor U17037 (N_17037,N_16836,N_16806);
and U17038 (N_17038,N_16825,N_16880);
and U17039 (N_17039,N_16922,N_16882);
nor U17040 (N_17040,N_16956,N_16950);
nor U17041 (N_17041,N_16835,N_16869);
and U17042 (N_17042,N_16849,N_16833);
and U17043 (N_17043,N_16805,N_16952);
nor U17044 (N_17044,N_16892,N_16901);
xor U17045 (N_17045,N_16935,N_16831);
or U17046 (N_17046,N_16872,N_16876);
nor U17047 (N_17047,N_16864,N_16913);
nand U17048 (N_17048,N_16816,N_16895);
xor U17049 (N_17049,N_16837,N_16892);
nor U17050 (N_17050,N_16823,N_16911);
and U17051 (N_17051,N_16912,N_16876);
and U17052 (N_17052,N_16885,N_16875);
xor U17053 (N_17053,N_16899,N_16808);
nor U17054 (N_17054,N_16884,N_16889);
xor U17055 (N_17055,N_16921,N_16890);
and U17056 (N_17056,N_16889,N_16954);
xor U17057 (N_17057,N_16919,N_16914);
nor U17058 (N_17058,N_16890,N_16834);
nor U17059 (N_17059,N_16897,N_16876);
or U17060 (N_17060,N_16885,N_16906);
nand U17061 (N_17061,N_16872,N_16893);
nand U17062 (N_17062,N_16926,N_16850);
and U17063 (N_17063,N_16899,N_16882);
xor U17064 (N_17064,N_16804,N_16895);
or U17065 (N_17065,N_16821,N_16880);
nand U17066 (N_17066,N_16916,N_16881);
xnor U17067 (N_17067,N_16887,N_16869);
xor U17068 (N_17068,N_16809,N_16804);
nor U17069 (N_17069,N_16881,N_16931);
and U17070 (N_17070,N_16810,N_16806);
or U17071 (N_17071,N_16928,N_16809);
or U17072 (N_17072,N_16902,N_16857);
xor U17073 (N_17073,N_16892,N_16933);
or U17074 (N_17074,N_16942,N_16857);
nand U17075 (N_17075,N_16888,N_16880);
or U17076 (N_17076,N_16929,N_16946);
and U17077 (N_17077,N_16806,N_16910);
nand U17078 (N_17078,N_16955,N_16924);
or U17079 (N_17079,N_16959,N_16809);
nand U17080 (N_17080,N_16879,N_16849);
or U17081 (N_17081,N_16948,N_16840);
xor U17082 (N_17082,N_16825,N_16948);
and U17083 (N_17083,N_16847,N_16875);
nand U17084 (N_17084,N_16886,N_16807);
nand U17085 (N_17085,N_16884,N_16958);
or U17086 (N_17086,N_16920,N_16916);
xor U17087 (N_17087,N_16957,N_16936);
nand U17088 (N_17088,N_16852,N_16831);
and U17089 (N_17089,N_16861,N_16864);
nor U17090 (N_17090,N_16913,N_16901);
xor U17091 (N_17091,N_16850,N_16803);
xnor U17092 (N_17092,N_16846,N_16918);
nand U17093 (N_17093,N_16800,N_16939);
nor U17094 (N_17094,N_16954,N_16809);
xor U17095 (N_17095,N_16881,N_16944);
nand U17096 (N_17096,N_16881,N_16955);
xor U17097 (N_17097,N_16911,N_16836);
nand U17098 (N_17098,N_16820,N_16918);
xnor U17099 (N_17099,N_16949,N_16809);
or U17100 (N_17100,N_16802,N_16882);
nor U17101 (N_17101,N_16880,N_16823);
xor U17102 (N_17102,N_16818,N_16820);
nand U17103 (N_17103,N_16828,N_16885);
nor U17104 (N_17104,N_16844,N_16835);
nor U17105 (N_17105,N_16816,N_16867);
nand U17106 (N_17106,N_16899,N_16853);
nand U17107 (N_17107,N_16895,N_16822);
or U17108 (N_17108,N_16906,N_16953);
nand U17109 (N_17109,N_16818,N_16949);
nand U17110 (N_17110,N_16840,N_16917);
and U17111 (N_17111,N_16878,N_16913);
nor U17112 (N_17112,N_16870,N_16872);
nand U17113 (N_17113,N_16936,N_16843);
and U17114 (N_17114,N_16842,N_16810);
xnor U17115 (N_17115,N_16856,N_16870);
or U17116 (N_17116,N_16890,N_16818);
xor U17117 (N_17117,N_16950,N_16937);
nand U17118 (N_17118,N_16801,N_16840);
or U17119 (N_17119,N_16955,N_16916);
and U17120 (N_17120,N_16965,N_16970);
nor U17121 (N_17121,N_17022,N_16968);
xor U17122 (N_17122,N_17019,N_17044);
nor U17123 (N_17123,N_17015,N_16992);
xnor U17124 (N_17124,N_17000,N_17032);
nor U17125 (N_17125,N_16996,N_17104);
or U17126 (N_17126,N_17078,N_17114);
nor U17127 (N_17127,N_17065,N_16962);
xnor U17128 (N_17128,N_17054,N_17002);
nor U17129 (N_17129,N_16975,N_17081);
xnor U17130 (N_17130,N_17005,N_17059);
nor U17131 (N_17131,N_17010,N_17118);
nor U17132 (N_17132,N_16993,N_17004);
or U17133 (N_17133,N_17098,N_17116);
or U17134 (N_17134,N_17058,N_16963);
or U17135 (N_17135,N_16995,N_17066);
xor U17136 (N_17136,N_16982,N_17012);
xnor U17137 (N_17137,N_16969,N_17047);
and U17138 (N_17138,N_17027,N_17034);
nand U17139 (N_17139,N_17049,N_16990);
xnor U17140 (N_17140,N_17028,N_17109);
and U17141 (N_17141,N_17008,N_17083);
and U17142 (N_17142,N_17030,N_16980);
or U17143 (N_17143,N_17043,N_17040);
and U17144 (N_17144,N_17075,N_17085);
xnor U17145 (N_17145,N_16989,N_17057);
or U17146 (N_17146,N_17045,N_17096);
and U17147 (N_17147,N_16967,N_17100);
or U17148 (N_17148,N_17079,N_17067);
xor U17149 (N_17149,N_17052,N_16971);
nand U17150 (N_17150,N_17029,N_17042);
or U17151 (N_17151,N_17089,N_16991);
xnor U17152 (N_17152,N_17108,N_17020);
nand U17153 (N_17153,N_17073,N_16972);
xor U17154 (N_17154,N_17064,N_17060);
or U17155 (N_17155,N_17031,N_17024);
and U17156 (N_17156,N_17050,N_16964);
or U17157 (N_17157,N_16987,N_17069);
xor U17158 (N_17158,N_17107,N_16985);
xnor U17159 (N_17159,N_17097,N_17101);
nor U17160 (N_17160,N_16974,N_17025);
nand U17161 (N_17161,N_17091,N_17117);
xor U17162 (N_17162,N_17090,N_17077);
or U17163 (N_17163,N_17110,N_17037);
and U17164 (N_17164,N_17046,N_17063);
or U17165 (N_17165,N_16976,N_17023);
nand U17166 (N_17166,N_17056,N_16973);
nor U17167 (N_17167,N_17080,N_17062);
xor U17168 (N_17168,N_17053,N_17082);
nand U17169 (N_17169,N_17111,N_17076);
xnor U17170 (N_17170,N_17086,N_17014);
or U17171 (N_17171,N_17061,N_16994);
and U17172 (N_17172,N_17055,N_17039);
nand U17173 (N_17173,N_17068,N_17102);
nor U17174 (N_17174,N_17094,N_17099);
nand U17175 (N_17175,N_17103,N_17095);
and U17176 (N_17176,N_16961,N_17021);
nor U17177 (N_17177,N_17016,N_17092);
nor U17178 (N_17178,N_17119,N_17009);
nand U17179 (N_17179,N_17087,N_16966);
or U17180 (N_17180,N_17070,N_17007);
xor U17181 (N_17181,N_17033,N_17115);
or U17182 (N_17182,N_17088,N_16999);
xnor U17183 (N_17183,N_17003,N_16960);
nand U17184 (N_17184,N_17113,N_17084);
nand U17185 (N_17185,N_17106,N_17071);
nand U17186 (N_17186,N_17112,N_16998);
or U17187 (N_17187,N_17026,N_17036);
xor U17188 (N_17188,N_17006,N_16978);
nand U17189 (N_17189,N_17011,N_17041);
nor U17190 (N_17190,N_16977,N_17048);
nand U17191 (N_17191,N_16983,N_17038);
nand U17192 (N_17192,N_17093,N_16981);
and U17193 (N_17193,N_16997,N_17013);
or U17194 (N_17194,N_16986,N_17035);
nand U17195 (N_17195,N_17017,N_17074);
and U17196 (N_17196,N_16984,N_17018);
and U17197 (N_17197,N_16988,N_17072);
nand U17198 (N_17198,N_17051,N_17105);
nor U17199 (N_17199,N_17001,N_16979);
nand U17200 (N_17200,N_16980,N_16973);
nand U17201 (N_17201,N_16992,N_17057);
and U17202 (N_17202,N_16973,N_17042);
nand U17203 (N_17203,N_17098,N_17065);
or U17204 (N_17204,N_17035,N_17049);
xor U17205 (N_17205,N_16997,N_17100);
nor U17206 (N_17206,N_17016,N_16995);
xnor U17207 (N_17207,N_17052,N_17046);
nor U17208 (N_17208,N_17033,N_17018);
or U17209 (N_17209,N_17084,N_17104);
nand U17210 (N_17210,N_17001,N_17117);
and U17211 (N_17211,N_17053,N_17077);
xor U17212 (N_17212,N_17009,N_17068);
or U17213 (N_17213,N_17104,N_17089);
and U17214 (N_17214,N_17075,N_17009);
or U17215 (N_17215,N_17017,N_17070);
nand U17216 (N_17216,N_17015,N_17038);
xnor U17217 (N_17217,N_17038,N_17077);
xnor U17218 (N_17218,N_17100,N_17118);
or U17219 (N_17219,N_17022,N_17119);
and U17220 (N_17220,N_17031,N_16984);
and U17221 (N_17221,N_17070,N_17032);
and U17222 (N_17222,N_17094,N_17078);
or U17223 (N_17223,N_17017,N_17029);
nand U17224 (N_17224,N_17053,N_17109);
or U17225 (N_17225,N_17074,N_16968);
nand U17226 (N_17226,N_17012,N_16963);
or U17227 (N_17227,N_17055,N_17015);
xnor U17228 (N_17228,N_17064,N_17075);
xor U17229 (N_17229,N_17054,N_17004);
nor U17230 (N_17230,N_17025,N_17108);
nand U17231 (N_17231,N_17110,N_16972);
or U17232 (N_17232,N_17100,N_17015);
nand U17233 (N_17233,N_17011,N_17009);
nor U17234 (N_17234,N_17002,N_16977);
xnor U17235 (N_17235,N_17035,N_17031);
or U17236 (N_17236,N_17101,N_17039);
or U17237 (N_17237,N_17087,N_17075);
nand U17238 (N_17238,N_17018,N_16996);
nand U17239 (N_17239,N_17008,N_17014);
xnor U17240 (N_17240,N_17041,N_17061);
and U17241 (N_17241,N_17081,N_17056);
and U17242 (N_17242,N_17078,N_16961);
and U17243 (N_17243,N_17091,N_17008);
nand U17244 (N_17244,N_17025,N_17043);
xnor U17245 (N_17245,N_17030,N_17046);
nor U17246 (N_17246,N_17035,N_17119);
and U17247 (N_17247,N_16996,N_17052);
xor U17248 (N_17248,N_17056,N_17015);
nor U17249 (N_17249,N_17105,N_16990);
or U17250 (N_17250,N_17100,N_17047);
xor U17251 (N_17251,N_16970,N_17115);
nand U17252 (N_17252,N_17114,N_17062);
xnor U17253 (N_17253,N_17113,N_17076);
xnor U17254 (N_17254,N_17019,N_17063);
or U17255 (N_17255,N_16982,N_17100);
and U17256 (N_17256,N_17027,N_16963);
nor U17257 (N_17257,N_17043,N_17061);
nand U17258 (N_17258,N_17006,N_17060);
and U17259 (N_17259,N_17071,N_17096);
and U17260 (N_17260,N_17027,N_17067);
xnor U17261 (N_17261,N_17052,N_16995);
nor U17262 (N_17262,N_17040,N_17055);
nand U17263 (N_17263,N_16987,N_17111);
xnor U17264 (N_17264,N_17017,N_17053);
and U17265 (N_17265,N_17042,N_17052);
nand U17266 (N_17266,N_17029,N_17066);
nand U17267 (N_17267,N_17098,N_17087);
or U17268 (N_17268,N_17012,N_17106);
xnor U17269 (N_17269,N_16982,N_17071);
and U17270 (N_17270,N_17115,N_16964);
or U17271 (N_17271,N_16965,N_17046);
and U17272 (N_17272,N_17047,N_17099);
or U17273 (N_17273,N_17095,N_17109);
and U17274 (N_17274,N_17025,N_17021);
nor U17275 (N_17275,N_17003,N_16996);
and U17276 (N_17276,N_16978,N_16965);
and U17277 (N_17277,N_17044,N_17012);
or U17278 (N_17278,N_17109,N_16969);
xor U17279 (N_17279,N_16979,N_17098);
and U17280 (N_17280,N_17196,N_17136);
xnor U17281 (N_17281,N_17174,N_17267);
xnor U17282 (N_17282,N_17126,N_17273);
and U17283 (N_17283,N_17168,N_17182);
xor U17284 (N_17284,N_17186,N_17250);
xnor U17285 (N_17285,N_17164,N_17180);
and U17286 (N_17286,N_17233,N_17151);
xor U17287 (N_17287,N_17225,N_17253);
or U17288 (N_17288,N_17248,N_17184);
nor U17289 (N_17289,N_17192,N_17226);
or U17290 (N_17290,N_17271,N_17159);
nand U17291 (N_17291,N_17134,N_17145);
nor U17292 (N_17292,N_17244,N_17178);
or U17293 (N_17293,N_17157,N_17137);
or U17294 (N_17294,N_17139,N_17197);
nand U17295 (N_17295,N_17149,N_17142);
and U17296 (N_17296,N_17247,N_17252);
nand U17297 (N_17297,N_17125,N_17155);
xnor U17298 (N_17298,N_17239,N_17211);
xor U17299 (N_17299,N_17243,N_17123);
nor U17300 (N_17300,N_17127,N_17229);
xor U17301 (N_17301,N_17122,N_17208);
nor U17302 (N_17302,N_17275,N_17200);
and U17303 (N_17303,N_17173,N_17189);
nand U17304 (N_17304,N_17202,N_17169);
nor U17305 (N_17305,N_17195,N_17141);
xnor U17306 (N_17306,N_17236,N_17223);
xnor U17307 (N_17307,N_17261,N_17181);
xor U17308 (N_17308,N_17165,N_17170);
nor U17309 (N_17309,N_17221,N_17166);
nor U17310 (N_17310,N_17150,N_17176);
nand U17311 (N_17311,N_17190,N_17259);
xnor U17312 (N_17312,N_17160,N_17177);
and U17313 (N_17313,N_17265,N_17209);
nor U17314 (N_17314,N_17213,N_17201);
nand U17315 (N_17315,N_17228,N_17218);
and U17316 (N_17316,N_17230,N_17220);
or U17317 (N_17317,N_17272,N_17167);
nor U17318 (N_17318,N_17279,N_17234);
nand U17319 (N_17319,N_17187,N_17245);
xor U17320 (N_17320,N_17255,N_17274);
nand U17321 (N_17321,N_17144,N_17152);
nor U17322 (N_17322,N_17257,N_17162);
xor U17323 (N_17323,N_17191,N_17148);
nor U17324 (N_17324,N_17277,N_17154);
nor U17325 (N_17325,N_17256,N_17132);
nor U17326 (N_17326,N_17179,N_17217);
nor U17327 (N_17327,N_17143,N_17214);
and U17328 (N_17328,N_17237,N_17207);
and U17329 (N_17329,N_17224,N_17212);
and U17330 (N_17330,N_17249,N_17227);
or U17331 (N_17331,N_17216,N_17246);
xnor U17332 (N_17332,N_17124,N_17266);
nor U17333 (N_17333,N_17242,N_17203);
nor U17334 (N_17334,N_17240,N_17172);
or U17335 (N_17335,N_17131,N_17268);
or U17336 (N_17336,N_17146,N_17232);
nor U17337 (N_17337,N_17276,N_17262);
or U17338 (N_17338,N_17193,N_17258);
or U17339 (N_17339,N_17235,N_17171);
or U17340 (N_17340,N_17138,N_17175);
and U17341 (N_17341,N_17260,N_17161);
or U17342 (N_17342,N_17264,N_17238);
and U17343 (N_17343,N_17140,N_17278);
nand U17344 (N_17344,N_17251,N_17183);
or U17345 (N_17345,N_17219,N_17128);
nor U17346 (N_17346,N_17130,N_17204);
or U17347 (N_17347,N_17222,N_17156);
nor U17348 (N_17348,N_17206,N_17210);
and U17349 (N_17349,N_17121,N_17194);
and U17350 (N_17350,N_17231,N_17133);
and U17351 (N_17351,N_17241,N_17135);
and U17352 (N_17352,N_17188,N_17199);
xor U17353 (N_17353,N_17153,N_17270);
or U17354 (N_17354,N_17158,N_17205);
or U17355 (N_17355,N_17254,N_17185);
or U17356 (N_17356,N_17147,N_17129);
and U17357 (N_17357,N_17163,N_17269);
xor U17358 (N_17358,N_17198,N_17215);
xor U17359 (N_17359,N_17120,N_17263);
nand U17360 (N_17360,N_17229,N_17131);
or U17361 (N_17361,N_17146,N_17162);
and U17362 (N_17362,N_17194,N_17128);
xnor U17363 (N_17363,N_17219,N_17142);
or U17364 (N_17364,N_17185,N_17133);
xor U17365 (N_17365,N_17156,N_17199);
nor U17366 (N_17366,N_17227,N_17171);
or U17367 (N_17367,N_17120,N_17264);
nor U17368 (N_17368,N_17204,N_17236);
nand U17369 (N_17369,N_17244,N_17193);
nand U17370 (N_17370,N_17162,N_17136);
nand U17371 (N_17371,N_17175,N_17174);
nor U17372 (N_17372,N_17191,N_17228);
nor U17373 (N_17373,N_17154,N_17269);
nor U17374 (N_17374,N_17210,N_17150);
or U17375 (N_17375,N_17226,N_17129);
and U17376 (N_17376,N_17144,N_17269);
xnor U17377 (N_17377,N_17156,N_17168);
nor U17378 (N_17378,N_17167,N_17198);
and U17379 (N_17379,N_17135,N_17234);
xnor U17380 (N_17380,N_17153,N_17195);
and U17381 (N_17381,N_17225,N_17257);
nand U17382 (N_17382,N_17228,N_17278);
or U17383 (N_17383,N_17244,N_17222);
or U17384 (N_17384,N_17166,N_17269);
nor U17385 (N_17385,N_17225,N_17204);
xnor U17386 (N_17386,N_17198,N_17185);
xor U17387 (N_17387,N_17271,N_17195);
or U17388 (N_17388,N_17217,N_17156);
nand U17389 (N_17389,N_17211,N_17183);
or U17390 (N_17390,N_17268,N_17195);
or U17391 (N_17391,N_17177,N_17199);
nand U17392 (N_17392,N_17151,N_17279);
xnor U17393 (N_17393,N_17197,N_17252);
nand U17394 (N_17394,N_17266,N_17139);
xor U17395 (N_17395,N_17154,N_17216);
nand U17396 (N_17396,N_17204,N_17124);
nor U17397 (N_17397,N_17220,N_17136);
nand U17398 (N_17398,N_17202,N_17131);
or U17399 (N_17399,N_17247,N_17256);
and U17400 (N_17400,N_17184,N_17218);
nand U17401 (N_17401,N_17127,N_17279);
and U17402 (N_17402,N_17139,N_17188);
xnor U17403 (N_17403,N_17175,N_17269);
xor U17404 (N_17404,N_17186,N_17141);
xnor U17405 (N_17405,N_17174,N_17134);
or U17406 (N_17406,N_17189,N_17226);
nor U17407 (N_17407,N_17271,N_17243);
xnor U17408 (N_17408,N_17221,N_17120);
and U17409 (N_17409,N_17254,N_17186);
nor U17410 (N_17410,N_17137,N_17275);
nand U17411 (N_17411,N_17127,N_17132);
or U17412 (N_17412,N_17164,N_17256);
or U17413 (N_17413,N_17210,N_17141);
xnor U17414 (N_17414,N_17169,N_17148);
xor U17415 (N_17415,N_17212,N_17236);
or U17416 (N_17416,N_17133,N_17240);
or U17417 (N_17417,N_17192,N_17187);
xor U17418 (N_17418,N_17261,N_17172);
nor U17419 (N_17419,N_17220,N_17164);
and U17420 (N_17420,N_17125,N_17231);
xor U17421 (N_17421,N_17140,N_17192);
nor U17422 (N_17422,N_17143,N_17236);
nand U17423 (N_17423,N_17210,N_17146);
xnor U17424 (N_17424,N_17278,N_17273);
and U17425 (N_17425,N_17137,N_17240);
xor U17426 (N_17426,N_17167,N_17229);
xor U17427 (N_17427,N_17145,N_17178);
or U17428 (N_17428,N_17184,N_17124);
or U17429 (N_17429,N_17160,N_17191);
nand U17430 (N_17430,N_17210,N_17213);
xor U17431 (N_17431,N_17224,N_17277);
nor U17432 (N_17432,N_17170,N_17276);
or U17433 (N_17433,N_17218,N_17264);
nand U17434 (N_17434,N_17163,N_17225);
or U17435 (N_17435,N_17180,N_17268);
nor U17436 (N_17436,N_17153,N_17192);
nand U17437 (N_17437,N_17245,N_17221);
nor U17438 (N_17438,N_17239,N_17122);
nand U17439 (N_17439,N_17278,N_17237);
nand U17440 (N_17440,N_17286,N_17346);
or U17441 (N_17441,N_17316,N_17285);
nand U17442 (N_17442,N_17427,N_17412);
nand U17443 (N_17443,N_17425,N_17348);
nor U17444 (N_17444,N_17337,N_17395);
nand U17445 (N_17445,N_17290,N_17378);
nor U17446 (N_17446,N_17399,N_17380);
nor U17447 (N_17447,N_17434,N_17372);
nor U17448 (N_17448,N_17439,N_17394);
nand U17449 (N_17449,N_17367,N_17392);
xnor U17450 (N_17450,N_17357,N_17389);
or U17451 (N_17451,N_17418,N_17349);
or U17452 (N_17452,N_17342,N_17319);
nor U17453 (N_17453,N_17291,N_17364);
or U17454 (N_17454,N_17374,N_17414);
nand U17455 (N_17455,N_17386,N_17402);
xor U17456 (N_17456,N_17338,N_17363);
or U17457 (N_17457,N_17426,N_17343);
xnor U17458 (N_17458,N_17366,N_17306);
and U17459 (N_17459,N_17437,N_17300);
xnor U17460 (N_17460,N_17317,N_17391);
nand U17461 (N_17461,N_17345,N_17350);
nor U17462 (N_17462,N_17292,N_17408);
or U17463 (N_17463,N_17326,N_17359);
or U17464 (N_17464,N_17315,N_17299);
and U17465 (N_17465,N_17329,N_17323);
xnor U17466 (N_17466,N_17409,N_17407);
xor U17467 (N_17467,N_17435,N_17303);
nor U17468 (N_17468,N_17419,N_17438);
and U17469 (N_17469,N_17436,N_17301);
and U17470 (N_17470,N_17324,N_17421);
and U17471 (N_17471,N_17356,N_17281);
or U17472 (N_17472,N_17430,N_17304);
nand U17473 (N_17473,N_17293,N_17390);
or U17474 (N_17474,N_17416,N_17410);
nand U17475 (N_17475,N_17289,N_17347);
xnor U17476 (N_17476,N_17397,N_17318);
xor U17477 (N_17477,N_17354,N_17280);
or U17478 (N_17478,N_17330,N_17352);
xnor U17479 (N_17479,N_17379,N_17369);
or U17480 (N_17480,N_17313,N_17344);
nand U17481 (N_17481,N_17353,N_17432);
and U17482 (N_17482,N_17295,N_17294);
xnor U17483 (N_17483,N_17384,N_17400);
and U17484 (N_17484,N_17358,N_17305);
nor U17485 (N_17485,N_17332,N_17288);
and U17486 (N_17486,N_17321,N_17302);
xnor U17487 (N_17487,N_17371,N_17341);
or U17488 (N_17488,N_17398,N_17360);
nand U17489 (N_17489,N_17393,N_17428);
nor U17490 (N_17490,N_17355,N_17388);
and U17491 (N_17491,N_17312,N_17308);
nand U17492 (N_17492,N_17382,N_17310);
or U17493 (N_17493,N_17339,N_17429);
nor U17494 (N_17494,N_17396,N_17284);
nor U17495 (N_17495,N_17385,N_17362);
nor U17496 (N_17496,N_17327,N_17334);
or U17497 (N_17497,N_17377,N_17387);
or U17498 (N_17498,N_17336,N_17307);
nor U17499 (N_17499,N_17376,N_17322);
nor U17500 (N_17500,N_17375,N_17413);
nand U17501 (N_17501,N_17298,N_17287);
and U17502 (N_17502,N_17411,N_17404);
or U17503 (N_17503,N_17424,N_17373);
nand U17504 (N_17504,N_17331,N_17405);
and U17505 (N_17505,N_17309,N_17361);
nand U17506 (N_17506,N_17314,N_17423);
and U17507 (N_17507,N_17297,N_17335);
xor U17508 (N_17508,N_17365,N_17403);
xnor U17509 (N_17509,N_17422,N_17431);
xnor U17510 (N_17510,N_17406,N_17328);
and U17511 (N_17511,N_17320,N_17370);
xor U17512 (N_17512,N_17433,N_17296);
nand U17513 (N_17513,N_17415,N_17351);
xor U17514 (N_17514,N_17325,N_17311);
nand U17515 (N_17515,N_17368,N_17282);
xnor U17516 (N_17516,N_17383,N_17340);
nand U17517 (N_17517,N_17420,N_17381);
nand U17518 (N_17518,N_17283,N_17401);
nor U17519 (N_17519,N_17333,N_17417);
nand U17520 (N_17520,N_17379,N_17325);
or U17521 (N_17521,N_17353,N_17288);
nand U17522 (N_17522,N_17423,N_17372);
xnor U17523 (N_17523,N_17389,N_17323);
and U17524 (N_17524,N_17288,N_17403);
and U17525 (N_17525,N_17415,N_17433);
nand U17526 (N_17526,N_17329,N_17342);
xnor U17527 (N_17527,N_17380,N_17294);
or U17528 (N_17528,N_17355,N_17414);
nor U17529 (N_17529,N_17322,N_17291);
nor U17530 (N_17530,N_17360,N_17346);
nand U17531 (N_17531,N_17397,N_17394);
nor U17532 (N_17532,N_17379,N_17405);
or U17533 (N_17533,N_17285,N_17294);
nand U17534 (N_17534,N_17386,N_17287);
nor U17535 (N_17535,N_17418,N_17307);
nor U17536 (N_17536,N_17307,N_17367);
and U17537 (N_17537,N_17370,N_17322);
or U17538 (N_17538,N_17368,N_17387);
xnor U17539 (N_17539,N_17291,N_17357);
and U17540 (N_17540,N_17396,N_17397);
nor U17541 (N_17541,N_17290,N_17387);
nand U17542 (N_17542,N_17359,N_17428);
xor U17543 (N_17543,N_17346,N_17385);
or U17544 (N_17544,N_17305,N_17389);
nand U17545 (N_17545,N_17330,N_17299);
nand U17546 (N_17546,N_17359,N_17379);
or U17547 (N_17547,N_17339,N_17362);
xnor U17548 (N_17548,N_17358,N_17384);
xor U17549 (N_17549,N_17364,N_17338);
and U17550 (N_17550,N_17319,N_17306);
nand U17551 (N_17551,N_17430,N_17419);
nand U17552 (N_17552,N_17372,N_17361);
nor U17553 (N_17553,N_17394,N_17374);
and U17554 (N_17554,N_17382,N_17393);
or U17555 (N_17555,N_17309,N_17290);
nand U17556 (N_17556,N_17389,N_17290);
and U17557 (N_17557,N_17369,N_17420);
and U17558 (N_17558,N_17283,N_17348);
xor U17559 (N_17559,N_17419,N_17388);
and U17560 (N_17560,N_17420,N_17408);
nand U17561 (N_17561,N_17345,N_17432);
xnor U17562 (N_17562,N_17423,N_17343);
and U17563 (N_17563,N_17417,N_17286);
and U17564 (N_17564,N_17307,N_17399);
nand U17565 (N_17565,N_17384,N_17335);
and U17566 (N_17566,N_17365,N_17287);
nor U17567 (N_17567,N_17316,N_17309);
nor U17568 (N_17568,N_17408,N_17318);
and U17569 (N_17569,N_17434,N_17320);
or U17570 (N_17570,N_17334,N_17353);
xnor U17571 (N_17571,N_17319,N_17343);
or U17572 (N_17572,N_17334,N_17406);
xor U17573 (N_17573,N_17390,N_17285);
or U17574 (N_17574,N_17380,N_17346);
xnor U17575 (N_17575,N_17401,N_17302);
nor U17576 (N_17576,N_17367,N_17406);
and U17577 (N_17577,N_17309,N_17281);
or U17578 (N_17578,N_17432,N_17366);
or U17579 (N_17579,N_17283,N_17315);
and U17580 (N_17580,N_17402,N_17434);
and U17581 (N_17581,N_17320,N_17391);
and U17582 (N_17582,N_17354,N_17395);
or U17583 (N_17583,N_17335,N_17380);
nor U17584 (N_17584,N_17360,N_17432);
or U17585 (N_17585,N_17430,N_17316);
nor U17586 (N_17586,N_17369,N_17324);
xnor U17587 (N_17587,N_17286,N_17292);
xor U17588 (N_17588,N_17389,N_17364);
and U17589 (N_17589,N_17302,N_17284);
nor U17590 (N_17590,N_17395,N_17416);
nand U17591 (N_17591,N_17298,N_17422);
nor U17592 (N_17592,N_17367,N_17353);
xor U17593 (N_17593,N_17428,N_17311);
and U17594 (N_17594,N_17284,N_17389);
and U17595 (N_17595,N_17385,N_17329);
and U17596 (N_17596,N_17329,N_17333);
nand U17597 (N_17597,N_17304,N_17405);
nand U17598 (N_17598,N_17399,N_17409);
xnor U17599 (N_17599,N_17368,N_17413);
or U17600 (N_17600,N_17548,N_17518);
xnor U17601 (N_17601,N_17449,N_17523);
and U17602 (N_17602,N_17462,N_17470);
xor U17603 (N_17603,N_17453,N_17474);
and U17604 (N_17604,N_17461,N_17599);
or U17605 (N_17605,N_17496,N_17564);
and U17606 (N_17606,N_17469,N_17537);
xnor U17607 (N_17607,N_17509,N_17551);
xor U17608 (N_17608,N_17465,N_17570);
and U17609 (N_17609,N_17484,N_17550);
nor U17610 (N_17610,N_17479,N_17597);
nor U17611 (N_17611,N_17504,N_17573);
nor U17612 (N_17612,N_17524,N_17489);
nand U17613 (N_17613,N_17500,N_17519);
xnor U17614 (N_17614,N_17534,N_17447);
nor U17615 (N_17615,N_17522,N_17460);
and U17616 (N_17616,N_17456,N_17579);
and U17617 (N_17617,N_17546,N_17584);
or U17618 (N_17618,N_17452,N_17587);
nand U17619 (N_17619,N_17440,N_17578);
nor U17620 (N_17620,N_17580,N_17533);
or U17621 (N_17621,N_17481,N_17468);
and U17622 (N_17622,N_17464,N_17556);
nand U17623 (N_17623,N_17554,N_17486);
nand U17624 (N_17624,N_17557,N_17539);
and U17625 (N_17625,N_17574,N_17517);
and U17626 (N_17626,N_17572,N_17511);
or U17627 (N_17627,N_17506,N_17581);
or U17628 (N_17628,N_17567,N_17591);
nand U17629 (N_17629,N_17478,N_17475);
nand U17630 (N_17630,N_17476,N_17463);
or U17631 (N_17631,N_17526,N_17542);
and U17632 (N_17632,N_17592,N_17528);
xnor U17633 (N_17633,N_17515,N_17467);
nor U17634 (N_17634,N_17596,N_17483);
and U17635 (N_17635,N_17594,N_17568);
nand U17636 (N_17636,N_17491,N_17482);
nor U17637 (N_17637,N_17445,N_17493);
nand U17638 (N_17638,N_17490,N_17516);
or U17639 (N_17639,N_17569,N_17543);
nor U17640 (N_17640,N_17450,N_17590);
or U17641 (N_17641,N_17510,N_17576);
or U17642 (N_17642,N_17575,N_17558);
nor U17643 (N_17643,N_17457,N_17507);
or U17644 (N_17644,N_17583,N_17571);
xor U17645 (N_17645,N_17497,N_17565);
xor U17646 (N_17646,N_17501,N_17494);
nand U17647 (N_17647,N_17595,N_17505);
nand U17648 (N_17648,N_17598,N_17446);
nor U17649 (N_17649,N_17540,N_17536);
nor U17650 (N_17650,N_17477,N_17547);
or U17651 (N_17651,N_17552,N_17527);
nor U17652 (N_17652,N_17555,N_17512);
and U17653 (N_17653,N_17538,N_17577);
and U17654 (N_17654,N_17466,N_17553);
nor U17655 (N_17655,N_17444,N_17459);
or U17656 (N_17656,N_17441,N_17455);
or U17657 (N_17657,N_17502,N_17589);
nor U17658 (N_17658,N_17549,N_17458);
nand U17659 (N_17659,N_17487,N_17513);
nor U17660 (N_17660,N_17499,N_17488);
or U17661 (N_17661,N_17473,N_17535);
or U17662 (N_17662,N_17471,N_17529);
or U17663 (N_17663,N_17566,N_17451);
nor U17664 (N_17664,N_17503,N_17521);
and U17665 (N_17665,N_17562,N_17530);
nand U17666 (N_17666,N_17508,N_17563);
or U17667 (N_17667,N_17480,N_17454);
nor U17668 (N_17668,N_17541,N_17593);
nand U17669 (N_17669,N_17544,N_17448);
nand U17670 (N_17670,N_17559,N_17561);
and U17671 (N_17671,N_17485,N_17582);
and U17672 (N_17672,N_17585,N_17520);
xnor U17673 (N_17673,N_17560,N_17588);
nand U17674 (N_17674,N_17525,N_17498);
nor U17675 (N_17675,N_17514,N_17545);
and U17676 (N_17676,N_17586,N_17443);
and U17677 (N_17677,N_17495,N_17532);
nor U17678 (N_17678,N_17492,N_17472);
or U17679 (N_17679,N_17442,N_17531);
nand U17680 (N_17680,N_17558,N_17561);
xor U17681 (N_17681,N_17576,N_17442);
or U17682 (N_17682,N_17502,N_17512);
nor U17683 (N_17683,N_17451,N_17469);
or U17684 (N_17684,N_17560,N_17494);
and U17685 (N_17685,N_17535,N_17511);
nor U17686 (N_17686,N_17569,N_17510);
and U17687 (N_17687,N_17572,N_17461);
or U17688 (N_17688,N_17586,N_17560);
nand U17689 (N_17689,N_17545,N_17503);
nor U17690 (N_17690,N_17480,N_17477);
nand U17691 (N_17691,N_17440,N_17451);
nand U17692 (N_17692,N_17545,N_17491);
nor U17693 (N_17693,N_17554,N_17566);
nor U17694 (N_17694,N_17482,N_17440);
nor U17695 (N_17695,N_17585,N_17515);
xnor U17696 (N_17696,N_17475,N_17491);
and U17697 (N_17697,N_17443,N_17446);
xor U17698 (N_17698,N_17456,N_17560);
xnor U17699 (N_17699,N_17514,N_17533);
and U17700 (N_17700,N_17550,N_17570);
and U17701 (N_17701,N_17508,N_17516);
and U17702 (N_17702,N_17564,N_17464);
and U17703 (N_17703,N_17598,N_17562);
or U17704 (N_17704,N_17440,N_17525);
or U17705 (N_17705,N_17572,N_17441);
nand U17706 (N_17706,N_17516,N_17519);
xnor U17707 (N_17707,N_17544,N_17562);
xor U17708 (N_17708,N_17482,N_17529);
xnor U17709 (N_17709,N_17526,N_17578);
nand U17710 (N_17710,N_17534,N_17553);
or U17711 (N_17711,N_17500,N_17588);
nor U17712 (N_17712,N_17554,N_17521);
nor U17713 (N_17713,N_17598,N_17492);
and U17714 (N_17714,N_17521,N_17526);
nor U17715 (N_17715,N_17527,N_17444);
xnor U17716 (N_17716,N_17493,N_17538);
or U17717 (N_17717,N_17529,N_17492);
or U17718 (N_17718,N_17469,N_17446);
and U17719 (N_17719,N_17444,N_17464);
nor U17720 (N_17720,N_17495,N_17471);
nor U17721 (N_17721,N_17555,N_17584);
xor U17722 (N_17722,N_17513,N_17570);
nor U17723 (N_17723,N_17470,N_17482);
and U17724 (N_17724,N_17504,N_17559);
nor U17725 (N_17725,N_17467,N_17526);
and U17726 (N_17726,N_17592,N_17455);
and U17727 (N_17727,N_17588,N_17533);
xnor U17728 (N_17728,N_17483,N_17564);
and U17729 (N_17729,N_17463,N_17595);
or U17730 (N_17730,N_17495,N_17507);
or U17731 (N_17731,N_17443,N_17507);
nand U17732 (N_17732,N_17507,N_17540);
nor U17733 (N_17733,N_17581,N_17473);
or U17734 (N_17734,N_17491,N_17457);
nand U17735 (N_17735,N_17453,N_17537);
or U17736 (N_17736,N_17572,N_17478);
nand U17737 (N_17737,N_17584,N_17592);
nand U17738 (N_17738,N_17538,N_17506);
or U17739 (N_17739,N_17470,N_17471);
and U17740 (N_17740,N_17505,N_17461);
xor U17741 (N_17741,N_17571,N_17545);
nand U17742 (N_17742,N_17543,N_17532);
nor U17743 (N_17743,N_17521,N_17518);
xnor U17744 (N_17744,N_17558,N_17465);
and U17745 (N_17745,N_17569,N_17506);
xnor U17746 (N_17746,N_17513,N_17470);
xnor U17747 (N_17747,N_17582,N_17492);
or U17748 (N_17748,N_17522,N_17510);
and U17749 (N_17749,N_17464,N_17474);
nand U17750 (N_17750,N_17503,N_17575);
nand U17751 (N_17751,N_17464,N_17584);
and U17752 (N_17752,N_17576,N_17548);
xor U17753 (N_17753,N_17457,N_17549);
nand U17754 (N_17754,N_17469,N_17528);
and U17755 (N_17755,N_17518,N_17563);
nor U17756 (N_17756,N_17526,N_17520);
nor U17757 (N_17757,N_17462,N_17445);
nand U17758 (N_17758,N_17536,N_17465);
or U17759 (N_17759,N_17447,N_17440);
or U17760 (N_17760,N_17653,N_17672);
nand U17761 (N_17761,N_17688,N_17693);
or U17762 (N_17762,N_17746,N_17670);
nor U17763 (N_17763,N_17735,N_17610);
or U17764 (N_17764,N_17682,N_17627);
nand U17765 (N_17765,N_17754,N_17758);
xnor U17766 (N_17766,N_17676,N_17622);
nand U17767 (N_17767,N_17647,N_17628);
or U17768 (N_17768,N_17717,N_17685);
nand U17769 (N_17769,N_17711,N_17741);
xnor U17770 (N_17770,N_17749,N_17751);
and U17771 (N_17771,N_17620,N_17675);
nor U17772 (N_17772,N_17652,N_17637);
and U17773 (N_17773,N_17655,N_17624);
xnor U17774 (N_17774,N_17696,N_17737);
nand U17775 (N_17775,N_17612,N_17736);
nand U17776 (N_17776,N_17643,N_17738);
nand U17777 (N_17777,N_17690,N_17601);
and U17778 (N_17778,N_17740,N_17646);
nand U17779 (N_17779,N_17635,N_17634);
or U17780 (N_17780,N_17704,N_17694);
xnor U17781 (N_17781,N_17753,N_17720);
and U17782 (N_17782,N_17708,N_17718);
and U17783 (N_17783,N_17695,N_17650);
and U17784 (N_17784,N_17605,N_17698);
xor U17785 (N_17785,N_17661,N_17644);
or U17786 (N_17786,N_17631,N_17702);
xnor U17787 (N_17787,N_17629,N_17674);
xnor U17788 (N_17788,N_17617,N_17719);
xor U17789 (N_17789,N_17728,N_17671);
nor U17790 (N_17790,N_17656,N_17697);
nand U17791 (N_17791,N_17734,N_17700);
nand U17792 (N_17792,N_17616,N_17667);
nand U17793 (N_17793,N_17621,N_17649);
and U17794 (N_17794,N_17713,N_17680);
and U17795 (N_17795,N_17614,N_17721);
nor U17796 (N_17796,N_17733,N_17744);
nor U17797 (N_17797,N_17683,N_17714);
and U17798 (N_17798,N_17684,N_17677);
or U17799 (N_17799,N_17665,N_17750);
xor U17800 (N_17800,N_17663,N_17701);
and U17801 (N_17801,N_17633,N_17630);
xnor U17802 (N_17802,N_17613,N_17757);
xor U17803 (N_17803,N_17664,N_17623);
or U17804 (N_17804,N_17619,N_17759);
nand U17805 (N_17805,N_17747,N_17729);
or U17806 (N_17806,N_17658,N_17712);
nor U17807 (N_17807,N_17699,N_17681);
or U17808 (N_17808,N_17615,N_17625);
nor U17809 (N_17809,N_17692,N_17668);
nor U17810 (N_17810,N_17611,N_17742);
and U17811 (N_17811,N_17705,N_17607);
nor U17812 (N_17812,N_17732,N_17756);
and U17813 (N_17813,N_17731,N_17745);
or U17814 (N_17814,N_17726,N_17748);
xnor U17815 (N_17815,N_17636,N_17618);
xnor U17816 (N_17816,N_17606,N_17642);
xnor U17817 (N_17817,N_17659,N_17716);
or U17818 (N_17818,N_17654,N_17722);
and U17819 (N_17819,N_17710,N_17730);
xor U17820 (N_17820,N_17673,N_17604);
nand U17821 (N_17821,N_17703,N_17727);
nor U17822 (N_17822,N_17666,N_17600);
and U17823 (N_17823,N_17755,N_17669);
nor U17824 (N_17824,N_17707,N_17626);
xnor U17825 (N_17825,N_17691,N_17662);
and U17826 (N_17826,N_17715,N_17752);
nor U17827 (N_17827,N_17640,N_17660);
and U17828 (N_17828,N_17645,N_17608);
or U17829 (N_17829,N_17724,N_17725);
or U17830 (N_17830,N_17678,N_17639);
xnor U17831 (N_17831,N_17706,N_17679);
xnor U17832 (N_17832,N_17632,N_17739);
nand U17833 (N_17833,N_17687,N_17602);
or U17834 (N_17834,N_17609,N_17709);
or U17835 (N_17835,N_17743,N_17603);
xor U17836 (N_17836,N_17651,N_17723);
nor U17837 (N_17837,N_17686,N_17648);
xor U17838 (N_17838,N_17657,N_17638);
nor U17839 (N_17839,N_17641,N_17689);
xnor U17840 (N_17840,N_17675,N_17682);
nand U17841 (N_17841,N_17642,N_17680);
xor U17842 (N_17842,N_17758,N_17620);
nand U17843 (N_17843,N_17751,N_17694);
nor U17844 (N_17844,N_17621,N_17643);
xor U17845 (N_17845,N_17694,N_17722);
xor U17846 (N_17846,N_17706,N_17654);
and U17847 (N_17847,N_17639,N_17602);
nand U17848 (N_17848,N_17650,N_17725);
nor U17849 (N_17849,N_17673,N_17602);
or U17850 (N_17850,N_17725,N_17607);
or U17851 (N_17851,N_17600,N_17606);
nand U17852 (N_17852,N_17687,N_17643);
nor U17853 (N_17853,N_17715,N_17753);
nor U17854 (N_17854,N_17644,N_17663);
xor U17855 (N_17855,N_17677,N_17676);
nor U17856 (N_17856,N_17667,N_17634);
nor U17857 (N_17857,N_17614,N_17640);
nor U17858 (N_17858,N_17674,N_17720);
nor U17859 (N_17859,N_17641,N_17733);
and U17860 (N_17860,N_17722,N_17738);
nor U17861 (N_17861,N_17714,N_17675);
nor U17862 (N_17862,N_17714,N_17688);
nor U17863 (N_17863,N_17600,N_17691);
or U17864 (N_17864,N_17637,N_17706);
nand U17865 (N_17865,N_17750,N_17639);
xor U17866 (N_17866,N_17647,N_17729);
or U17867 (N_17867,N_17737,N_17679);
or U17868 (N_17868,N_17618,N_17671);
nor U17869 (N_17869,N_17626,N_17630);
and U17870 (N_17870,N_17654,N_17648);
or U17871 (N_17871,N_17649,N_17604);
and U17872 (N_17872,N_17618,N_17612);
nand U17873 (N_17873,N_17626,N_17684);
nand U17874 (N_17874,N_17624,N_17668);
nand U17875 (N_17875,N_17755,N_17753);
nand U17876 (N_17876,N_17679,N_17629);
xor U17877 (N_17877,N_17678,N_17672);
nand U17878 (N_17878,N_17618,N_17680);
xor U17879 (N_17879,N_17724,N_17718);
nor U17880 (N_17880,N_17732,N_17749);
nor U17881 (N_17881,N_17757,N_17728);
nand U17882 (N_17882,N_17609,N_17695);
xor U17883 (N_17883,N_17727,N_17712);
nor U17884 (N_17884,N_17602,N_17650);
or U17885 (N_17885,N_17638,N_17675);
or U17886 (N_17886,N_17688,N_17684);
xor U17887 (N_17887,N_17644,N_17675);
and U17888 (N_17888,N_17711,N_17726);
and U17889 (N_17889,N_17639,N_17650);
xnor U17890 (N_17890,N_17698,N_17615);
nand U17891 (N_17891,N_17690,N_17722);
xnor U17892 (N_17892,N_17683,N_17618);
or U17893 (N_17893,N_17714,N_17695);
or U17894 (N_17894,N_17687,N_17600);
nand U17895 (N_17895,N_17712,N_17755);
or U17896 (N_17896,N_17660,N_17606);
or U17897 (N_17897,N_17637,N_17749);
and U17898 (N_17898,N_17666,N_17668);
nor U17899 (N_17899,N_17638,N_17758);
and U17900 (N_17900,N_17600,N_17721);
nand U17901 (N_17901,N_17728,N_17650);
nand U17902 (N_17902,N_17600,N_17653);
xor U17903 (N_17903,N_17622,N_17670);
xor U17904 (N_17904,N_17658,N_17675);
nand U17905 (N_17905,N_17670,N_17728);
xnor U17906 (N_17906,N_17661,N_17736);
or U17907 (N_17907,N_17605,N_17663);
nor U17908 (N_17908,N_17624,N_17630);
xnor U17909 (N_17909,N_17733,N_17677);
or U17910 (N_17910,N_17604,N_17678);
nor U17911 (N_17911,N_17644,N_17711);
xor U17912 (N_17912,N_17747,N_17616);
nor U17913 (N_17913,N_17667,N_17650);
xnor U17914 (N_17914,N_17725,N_17616);
nor U17915 (N_17915,N_17618,N_17656);
nor U17916 (N_17916,N_17742,N_17679);
and U17917 (N_17917,N_17663,N_17730);
and U17918 (N_17918,N_17612,N_17643);
nand U17919 (N_17919,N_17640,N_17627);
nand U17920 (N_17920,N_17907,N_17881);
nand U17921 (N_17921,N_17829,N_17904);
nor U17922 (N_17922,N_17898,N_17871);
or U17923 (N_17923,N_17833,N_17780);
nand U17924 (N_17924,N_17854,N_17783);
or U17925 (N_17925,N_17803,N_17787);
or U17926 (N_17926,N_17834,N_17797);
nor U17927 (N_17927,N_17918,N_17794);
or U17928 (N_17928,N_17855,N_17826);
nor U17929 (N_17929,N_17909,N_17913);
nor U17930 (N_17930,N_17838,N_17901);
xnor U17931 (N_17931,N_17874,N_17844);
or U17932 (N_17932,N_17813,N_17806);
xnor U17933 (N_17933,N_17786,N_17825);
nand U17934 (N_17934,N_17796,N_17877);
or U17935 (N_17935,N_17775,N_17872);
xnor U17936 (N_17936,N_17883,N_17908);
or U17937 (N_17937,N_17882,N_17763);
nor U17938 (N_17938,N_17795,N_17876);
xor U17939 (N_17939,N_17867,N_17764);
nor U17940 (N_17940,N_17802,N_17866);
nor U17941 (N_17941,N_17864,N_17820);
nand U17942 (N_17942,N_17886,N_17770);
nand U17943 (N_17943,N_17902,N_17879);
or U17944 (N_17944,N_17812,N_17809);
nor U17945 (N_17945,N_17800,N_17859);
xnor U17946 (N_17946,N_17817,N_17840);
and U17947 (N_17947,N_17816,N_17841);
xnor U17948 (N_17948,N_17889,N_17765);
nor U17949 (N_17949,N_17789,N_17822);
nor U17950 (N_17950,N_17818,N_17837);
nand U17951 (N_17951,N_17891,N_17848);
and U17952 (N_17952,N_17870,N_17823);
xor U17953 (N_17953,N_17836,N_17845);
or U17954 (N_17954,N_17776,N_17779);
xnor U17955 (N_17955,N_17914,N_17778);
xor U17956 (N_17956,N_17884,N_17856);
nor U17957 (N_17957,N_17861,N_17835);
xnor U17958 (N_17958,N_17828,N_17819);
nor U17959 (N_17959,N_17893,N_17852);
or U17960 (N_17960,N_17865,N_17810);
nor U17961 (N_17961,N_17896,N_17821);
xnor U17962 (N_17962,N_17824,N_17912);
nor U17963 (N_17963,N_17830,N_17788);
nor U17964 (N_17964,N_17769,N_17792);
or U17965 (N_17965,N_17842,N_17799);
or U17966 (N_17966,N_17808,N_17790);
or U17967 (N_17967,N_17862,N_17811);
and U17968 (N_17968,N_17804,N_17895);
nand U17969 (N_17969,N_17839,N_17777);
nand U17970 (N_17970,N_17911,N_17793);
xnor U17971 (N_17971,N_17869,N_17791);
nor U17972 (N_17972,N_17863,N_17760);
and U17973 (N_17973,N_17860,N_17885);
nor U17974 (N_17974,N_17875,N_17815);
nor U17975 (N_17975,N_17849,N_17903);
nand U17976 (N_17976,N_17857,N_17880);
or U17977 (N_17977,N_17846,N_17851);
xnor U17978 (N_17978,N_17919,N_17827);
and U17979 (N_17979,N_17772,N_17773);
nand U17980 (N_17980,N_17892,N_17847);
xor U17981 (N_17981,N_17897,N_17878);
and U17982 (N_17982,N_17853,N_17782);
xnor U17983 (N_17983,N_17767,N_17873);
or U17984 (N_17984,N_17805,N_17766);
or U17985 (N_17985,N_17894,N_17814);
nand U17986 (N_17986,N_17850,N_17801);
nand U17987 (N_17987,N_17784,N_17910);
xnor U17988 (N_17988,N_17785,N_17887);
or U17989 (N_17989,N_17888,N_17807);
or U17990 (N_17990,N_17900,N_17906);
or U17991 (N_17991,N_17858,N_17843);
or U17992 (N_17992,N_17868,N_17915);
and U17993 (N_17993,N_17832,N_17774);
or U17994 (N_17994,N_17762,N_17781);
and U17995 (N_17995,N_17768,N_17917);
xnor U17996 (N_17996,N_17916,N_17890);
nor U17997 (N_17997,N_17761,N_17771);
nand U17998 (N_17998,N_17798,N_17899);
nand U17999 (N_17999,N_17905,N_17831);
xnor U18000 (N_18000,N_17869,N_17877);
nand U18001 (N_18001,N_17896,N_17881);
or U18002 (N_18002,N_17765,N_17818);
nor U18003 (N_18003,N_17841,N_17818);
nand U18004 (N_18004,N_17917,N_17891);
xnor U18005 (N_18005,N_17882,N_17807);
and U18006 (N_18006,N_17889,N_17786);
xor U18007 (N_18007,N_17800,N_17850);
or U18008 (N_18008,N_17780,N_17876);
nand U18009 (N_18009,N_17796,N_17805);
and U18010 (N_18010,N_17910,N_17837);
xnor U18011 (N_18011,N_17916,N_17877);
nand U18012 (N_18012,N_17918,N_17816);
nand U18013 (N_18013,N_17812,N_17777);
nand U18014 (N_18014,N_17905,N_17885);
and U18015 (N_18015,N_17796,N_17847);
nand U18016 (N_18016,N_17877,N_17799);
nor U18017 (N_18017,N_17835,N_17867);
or U18018 (N_18018,N_17811,N_17804);
or U18019 (N_18019,N_17899,N_17818);
nand U18020 (N_18020,N_17787,N_17867);
nand U18021 (N_18021,N_17762,N_17805);
or U18022 (N_18022,N_17792,N_17858);
nor U18023 (N_18023,N_17875,N_17792);
and U18024 (N_18024,N_17775,N_17887);
nor U18025 (N_18025,N_17884,N_17771);
and U18026 (N_18026,N_17850,N_17837);
nor U18027 (N_18027,N_17896,N_17859);
nor U18028 (N_18028,N_17919,N_17803);
and U18029 (N_18029,N_17779,N_17831);
and U18030 (N_18030,N_17794,N_17790);
or U18031 (N_18031,N_17843,N_17763);
xor U18032 (N_18032,N_17865,N_17822);
xor U18033 (N_18033,N_17850,N_17784);
or U18034 (N_18034,N_17787,N_17771);
and U18035 (N_18035,N_17897,N_17901);
nand U18036 (N_18036,N_17851,N_17884);
and U18037 (N_18037,N_17913,N_17857);
nor U18038 (N_18038,N_17877,N_17792);
and U18039 (N_18039,N_17847,N_17844);
nor U18040 (N_18040,N_17836,N_17838);
and U18041 (N_18041,N_17828,N_17882);
xnor U18042 (N_18042,N_17880,N_17911);
xnor U18043 (N_18043,N_17761,N_17879);
and U18044 (N_18044,N_17871,N_17775);
xnor U18045 (N_18045,N_17788,N_17888);
nand U18046 (N_18046,N_17762,N_17827);
nand U18047 (N_18047,N_17806,N_17767);
nand U18048 (N_18048,N_17806,N_17874);
nor U18049 (N_18049,N_17892,N_17772);
and U18050 (N_18050,N_17854,N_17773);
nand U18051 (N_18051,N_17789,N_17896);
and U18052 (N_18052,N_17914,N_17812);
nand U18053 (N_18053,N_17789,N_17804);
or U18054 (N_18054,N_17834,N_17763);
or U18055 (N_18055,N_17887,N_17830);
nand U18056 (N_18056,N_17791,N_17772);
xor U18057 (N_18057,N_17893,N_17915);
xor U18058 (N_18058,N_17817,N_17858);
or U18059 (N_18059,N_17856,N_17839);
and U18060 (N_18060,N_17798,N_17794);
nand U18061 (N_18061,N_17885,N_17889);
and U18062 (N_18062,N_17809,N_17775);
xnor U18063 (N_18063,N_17838,N_17816);
nand U18064 (N_18064,N_17762,N_17824);
and U18065 (N_18065,N_17913,N_17862);
and U18066 (N_18066,N_17890,N_17777);
and U18067 (N_18067,N_17798,N_17894);
and U18068 (N_18068,N_17855,N_17891);
nor U18069 (N_18069,N_17910,N_17818);
and U18070 (N_18070,N_17914,N_17784);
nor U18071 (N_18071,N_17771,N_17909);
xnor U18072 (N_18072,N_17798,N_17797);
xnor U18073 (N_18073,N_17801,N_17840);
nor U18074 (N_18074,N_17798,N_17781);
nor U18075 (N_18075,N_17781,N_17877);
or U18076 (N_18076,N_17910,N_17905);
nand U18077 (N_18077,N_17837,N_17765);
nand U18078 (N_18078,N_17788,N_17822);
and U18079 (N_18079,N_17893,N_17903);
nand U18080 (N_18080,N_17975,N_17966);
or U18081 (N_18081,N_17967,N_18054);
xnor U18082 (N_18082,N_17928,N_18018);
or U18083 (N_18083,N_17920,N_17939);
nand U18084 (N_18084,N_18017,N_18042);
xor U18085 (N_18085,N_18068,N_18050);
and U18086 (N_18086,N_17971,N_18013);
nor U18087 (N_18087,N_17973,N_17964);
and U18088 (N_18088,N_18055,N_18064);
nand U18089 (N_18089,N_17969,N_17930);
nor U18090 (N_18090,N_18029,N_18075);
nand U18091 (N_18091,N_17929,N_17993);
nor U18092 (N_18092,N_18000,N_18051);
or U18093 (N_18093,N_17933,N_17996);
xor U18094 (N_18094,N_18030,N_17992);
nor U18095 (N_18095,N_17963,N_17995);
nand U18096 (N_18096,N_18070,N_18033);
xnor U18097 (N_18097,N_17994,N_17924);
nand U18098 (N_18098,N_17934,N_18052);
nor U18099 (N_18099,N_18015,N_17926);
nand U18100 (N_18100,N_17978,N_18048);
nor U18101 (N_18101,N_18006,N_18026);
xor U18102 (N_18102,N_17981,N_18061);
nand U18103 (N_18103,N_18002,N_18073);
nand U18104 (N_18104,N_18071,N_18022);
and U18105 (N_18105,N_17997,N_17958);
and U18106 (N_18106,N_17946,N_17940);
and U18107 (N_18107,N_18014,N_17947);
nor U18108 (N_18108,N_18041,N_17982);
nor U18109 (N_18109,N_18020,N_18045);
xor U18110 (N_18110,N_17941,N_17990);
or U18111 (N_18111,N_17972,N_18032);
nor U18112 (N_18112,N_17959,N_18076);
and U18113 (N_18113,N_17953,N_18058);
nor U18114 (N_18114,N_18039,N_17985);
or U18115 (N_18115,N_18005,N_17938);
and U18116 (N_18116,N_18024,N_17998);
or U18117 (N_18117,N_18062,N_18049);
or U18118 (N_18118,N_17991,N_17980);
nor U18119 (N_18119,N_17943,N_17944);
xnor U18120 (N_18120,N_17956,N_18046);
xor U18121 (N_18121,N_18031,N_18034);
nor U18122 (N_18122,N_18021,N_18057);
and U18123 (N_18123,N_18067,N_17925);
and U18124 (N_18124,N_18044,N_17983);
or U18125 (N_18125,N_18009,N_17921);
nand U18126 (N_18126,N_17988,N_18037);
nor U18127 (N_18127,N_18069,N_18028);
nor U18128 (N_18128,N_17935,N_18001);
and U18129 (N_18129,N_17976,N_18035);
or U18130 (N_18130,N_17962,N_17989);
nand U18131 (N_18131,N_17954,N_17987);
nand U18132 (N_18132,N_17999,N_17984);
or U18133 (N_18133,N_18008,N_17949);
xnor U18134 (N_18134,N_18025,N_17952);
nand U18135 (N_18135,N_17965,N_17951);
nand U18136 (N_18136,N_17977,N_17979);
or U18137 (N_18137,N_17945,N_18016);
nand U18138 (N_18138,N_18010,N_17942);
xor U18139 (N_18139,N_17974,N_18007);
and U18140 (N_18140,N_17957,N_18056);
nand U18141 (N_18141,N_17986,N_18059);
and U18142 (N_18142,N_17961,N_18065);
nand U18143 (N_18143,N_17948,N_17970);
nand U18144 (N_18144,N_18038,N_17931);
or U18145 (N_18145,N_17950,N_18074);
and U18146 (N_18146,N_18063,N_17968);
nand U18147 (N_18147,N_17932,N_18047);
and U18148 (N_18148,N_17927,N_18053);
or U18149 (N_18149,N_18023,N_18012);
xor U18150 (N_18150,N_18027,N_17960);
nand U18151 (N_18151,N_18079,N_18036);
nor U18152 (N_18152,N_18019,N_18003);
nor U18153 (N_18153,N_18011,N_18060);
nor U18154 (N_18154,N_18066,N_18072);
or U18155 (N_18155,N_18043,N_17936);
nand U18156 (N_18156,N_18004,N_17923);
or U18157 (N_18157,N_18077,N_17937);
or U18158 (N_18158,N_18078,N_18040);
or U18159 (N_18159,N_17922,N_17955);
or U18160 (N_18160,N_17935,N_17955);
xor U18161 (N_18161,N_17994,N_18039);
nor U18162 (N_18162,N_17931,N_17922);
xnor U18163 (N_18163,N_18071,N_17943);
or U18164 (N_18164,N_17997,N_18043);
nand U18165 (N_18165,N_18050,N_18037);
nor U18166 (N_18166,N_17978,N_17979);
xor U18167 (N_18167,N_18014,N_18022);
nand U18168 (N_18168,N_17926,N_18048);
or U18169 (N_18169,N_17940,N_18057);
nor U18170 (N_18170,N_17989,N_18012);
and U18171 (N_18171,N_17992,N_17999);
xnor U18172 (N_18172,N_18034,N_17976);
or U18173 (N_18173,N_17928,N_18047);
or U18174 (N_18174,N_17930,N_17979);
nand U18175 (N_18175,N_17924,N_18026);
nor U18176 (N_18176,N_17937,N_17931);
or U18177 (N_18177,N_17942,N_17976);
xor U18178 (N_18178,N_18004,N_18065);
nor U18179 (N_18179,N_17921,N_18058);
xor U18180 (N_18180,N_18029,N_18064);
or U18181 (N_18181,N_17932,N_18053);
nand U18182 (N_18182,N_17995,N_18063);
xnor U18183 (N_18183,N_18000,N_17945);
and U18184 (N_18184,N_18041,N_17924);
nand U18185 (N_18185,N_18042,N_17933);
or U18186 (N_18186,N_17993,N_18019);
nand U18187 (N_18187,N_17929,N_18059);
nand U18188 (N_18188,N_17923,N_18017);
and U18189 (N_18189,N_18034,N_17923);
or U18190 (N_18190,N_18055,N_17935);
nand U18191 (N_18191,N_18071,N_17973);
nor U18192 (N_18192,N_18017,N_18031);
nor U18193 (N_18193,N_18043,N_17973);
or U18194 (N_18194,N_18067,N_17980);
or U18195 (N_18195,N_18034,N_17933);
and U18196 (N_18196,N_18059,N_18040);
nand U18197 (N_18197,N_18027,N_18062);
and U18198 (N_18198,N_17982,N_18076);
or U18199 (N_18199,N_17947,N_18050);
or U18200 (N_18200,N_18021,N_17974);
xor U18201 (N_18201,N_18012,N_18013);
nor U18202 (N_18202,N_18072,N_17950);
xnor U18203 (N_18203,N_17932,N_18039);
nand U18204 (N_18204,N_17996,N_18067);
nand U18205 (N_18205,N_18024,N_18040);
nor U18206 (N_18206,N_18069,N_18008);
nand U18207 (N_18207,N_18009,N_17949);
or U18208 (N_18208,N_17937,N_17925);
nand U18209 (N_18209,N_17923,N_17987);
or U18210 (N_18210,N_17985,N_18037);
nor U18211 (N_18211,N_18073,N_17999);
and U18212 (N_18212,N_17998,N_17938);
nor U18213 (N_18213,N_17944,N_17995);
and U18214 (N_18214,N_18006,N_18040);
or U18215 (N_18215,N_17927,N_18054);
or U18216 (N_18216,N_18072,N_17995);
and U18217 (N_18217,N_18070,N_18046);
nor U18218 (N_18218,N_17935,N_18010);
or U18219 (N_18219,N_17945,N_17942);
nand U18220 (N_18220,N_17935,N_18077);
or U18221 (N_18221,N_18070,N_18057);
nor U18222 (N_18222,N_18039,N_18076);
nand U18223 (N_18223,N_18048,N_17952);
xor U18224 (N_18224,N_18068,N_17929);
nand U18225 (N_18225,N_18008,N_17920);
xor U18226 (N_18226,N_18049,N_18045);
nand U18227 (N_18227,N_17954,N_18059);
xor U18228 (N_18228,N_17931,N_18008);
and U18229 (N_18229,N_18042,N_18001);
and U18230 (N_18230,N_18040,N_17961);
nand U18231 (N_18231,N_17932,N_18052);
and U18232 (N_18232,N_17973,N_17978);
nor U18233 (N_18233,N_17944,N_17968);
nor U18234 (N_18234,N_18034,N_18027);
nand U18235 (N_18235,N_18004,N_18036);
nand U18236 (N_18236,N_18027,N_18017);
nand U18237 (N_18237,N_17996,N_18052);
nor U18238 (N_18238,N_18066,N_17938);
xnor U18239 (N_18239,N_17923,N_18007);
or U18240 (N_18240,N_18085,N_18230);
or U18241 (N_18241,N_18208,N_18180);
and U18242 (N_18242,N_18216,N_18092);
and U18243 (N_18243,N_18174,N_18162);
and U18244 (N_18244,N_18119,N_18235);
and U18245 (N_18245,N_18196,N_18219);
xnor U18246 (N_18246,N_18133,N_18194);
or U18247 (N_18247,N_18081,N_18086);
nor U18248 (N_18248,N_18125,N_18179);
xnor U18249 (N_18249,N_18239,N_18183);
nand U18250 (N_18250,N_18226,N_18134);
or U18251 (N_18251,N_18200,N_18093);
and U18252 (N_18252,N_18204,N_18189);
nor U18253 (N_18253,N_18181,N_18228);
nor U18254 (N_18254,N_18236,N_18090);
nor U18255 (N_18255,N_18206,N_18156);
nand U18256 (N_18256,N_18182,N_18148);
or U18257 (N_18257,N_18102,N_18215);
nor U18258 (N_18258,N_18229,N_18187);
nor U18259 (N_18259,N_18130,N_18198);
and U18260 (N_18260,N_18153,N_18186);
and U18261 (N_18261,N_18136,N_18225);
nor U18262 (N_18262,N_18161,N_18207);
and U18263 (N_18263,N_18110,N_18096);
nand U18264 (N_18264,N_18115,N_18087);
or U18265 (N_18265,N_18117,N_18105);
nand U18266 (N_18266,N_18201,N_18113);
or U18267 (N_18267,N_18160,N_18095);
and U18268 (N_18268,N_18137,N_18164);
nor U18269 (N_18269,N_18214,N_18172);
nor U18270 (N_18270,N_18151,N_18108);
or U18271 (N_18271,N_18231,N_18211);
nand U18272 (N_18272,N_18190,N_18112);
and U18273 (N_18273,N_18205,N_18222);
nand U18274 (N_18274,N_18238,N_18233);
and U18275 (N_18275,N_18171,N_18101);
xor U18276 (N_18276,N_18155,N_18122);
nor U18277 (N_18277,N_18146,N_18184);
nand U18278 (N_18278,N_18209,N_18109);
and U18279 (N_18279,N_18167,N_18188);
and U18280 (N_18280,N_18132,N_18131);
and U18281 (N_18281,N_18124,N_18121);
xnor U18282 (N_18282,N_18203,N_18145);
or U18283 (N_18283,N_18158,N_18232);
nor U18284 (N_18284,N_18199,N_18138);
nor U18285 (N_18285,N_18217,N_18170);
nand U18286 (N_18286,N_18106,N_18103);
or U18287 (N_18287,N_18213,N_18089);
nand U18288 (N_18288,N_18129,N_18192);
nor U18289 (N_18289,N_18154,N_18227);
or U18290 (N_18290,N_18177,N_18126);
nor U18291 (N_18291,N_18099,N_18100);
and U18292 (N_18292,N_18191,N_18127);
or U18293 (N_18293,N_18150,N_18135);
or U18294 (N_18294,N_18080,N_18223);
xor U18295 (N_18295,N_18224,N_18193);
and U18296 (N_18296,N_18143,N_18178);
xnor U18297 (N_18297,N_18166,N_18149);
xor U18298 (N_18298,N_18212,N_18091);
nand U18299 (N_18299,N_18176,N_18141);
and U18300 (N_18300,N_18107,N_18202);
nor U18301 (N_18301,N_18142,N_18197);
and U18302 (N_18302,N_18157,N_18175);
and U18303 (N_18303,N_18120,N_18140);
nand U18304 (N_18304,N_18118,N_18152);
nand U18305 (N_18305,N_18221,N_18185);
and U18306 (N_18306,N_18234,N_18163);
xnor U18307 (N_18307,N_18123,N_18195);
nand U18308 (N_18308,N_18098,N_18168);
nor U18309 (N_18309,N_18165,N_18116);
nor U18310 (N_18310,N_18159,N_18210);
xor U18311 (N_18311,N_18084,N_18139);
nor U18312 (N_18312,N_18111,N_18083);
nor U18313 (N_18313,N_18094,N_18173);
xnor U18314 (N_18314,N_18114,N_18218);
xnor U18315 (N_18315,N_18237,N_18088);
nor U18316 (N_18316,N_18104,N_18128);
xnor U18317 (N_18317,N_18144,N_18220);
nand U18318 (N_18318,N_18082,N_18097);
nor U18319 (N_18319,N_18169,N_18147);
and U18320 (N_18320,N_18151,N_18080);
xnor U18321 (N_18321,N_18101,N_18090);
and U18322 (N_18322,N_18150,N_18220);
and U18323 (N_18323,N_18228,N_18118);
and U18324 (N_18324,N_18118,N_18234);
xor U18325 (N_18325,N_18085,N_18198);
nand U18326 (N_18326,N_18105,N_18205);
nand U18327 (N_18327,N_18123,N_18118);
and U18328 (N_18328,N_18218,N_18188);
and U18329 (N_18329,N_18233,N_18095);
or U18330 (N_18330,N_18181,N_18164);
or U18331 (N_18331,N_18121,N_18128);
and U18332 (N_18332,N_18085,N_18181);
or U18333 (N_18333,N_18098,N_18156);
nand U18334 (N_18334,N_18103,N_18086);
xor U18335 (N_18335,N_18174,N_18164);
xnor U18336 (N_18336,N_18176,N_18194);
or U18337 (N_18337,N_18239,N_18111);
and U18338 (N_18338,N_18096,N_18137);
xor U18339 (N_18339,N_18138,N_18223);
or U18340 (N_18340,N_18235,N_18103);
nor U18341 (N_18341,N_18201,N_18153);
nand U18342 (N_18342,N_18186,N_18179);
nand U18343 (N_18343,N_18127,N_18198);
and U18344 (N_18344,N_18201,N_18114);
nor U18345 (N_18345,N_18207,N_18163);
nor U18346 (N_18346,N_18170,N_18196);
or U18347 (N_18347,N_18218,N_18143);
nand U18348 (N_18348,N_18133,N_18113);
and U18349 (N_18349,N_18234,N_18094);
or U18350 (N_18350,N_18164,N_18120);
nor U18351 (N_18351,N_18157,N_18235);
nand U18352 (N_18352,N_18137,N_18139);
xor U18353 (N_18353,N_18104,N_18175);
nand U18354 (N_18354,N_18139,N_18173);
nand U18355 (N_18355,N_18168,N_18162);
xor U18356 (N_18356,N_18132,N_18196);
nor U18357 (N_18357,N_18084,N_18140);
xor U18358 (N_18358,N_18158,N_18098);
nand U18359 (N_18359,N_18217,N_18134);
nor U18360 (N_18360,N_18146,N_18130);
xor U18361 (N_18361,N_18088,N_18205);
or U18362 (N_18362,N_18216,N_18103);
and U18363 (N_18363,N_18094,N_18207);
nor U18364 (N_18364,N_18233,N_18211);
or U18365 (N_18365,N_18232,N_18141);
nand U18366 (N_18366,N_18185,N_18199);
xnor U18367 (N_18367,N_18086,N_18119);
nand U18368 (N_18368,N_18190,N_18230);
nand U18369 (N_18369,N_18170,N_18235);
xor U18370 (N_18370,N_18234,N_18189);
xor U18371 (N_18371,N_18155,N_18139);
and U18372 (N_18372,N_18192,N_18150);
and U18373 (N_18373,N_18108,N_18134);
nand U18374 (N_18374,N_18171,N_18127);
nand U18375 (N_18375,N_18189,N_18093);
and U18376 (N_18376,N_18231,N_18229);
nand U18377 (N_18377,N_18183,N_18202);
nand U18378 (N_18378,N_18169,N_18115);
nor U18379 (N_18379,N_18142,N_18094);
xor U18380 (N_18380,N_18228,N_18184);
and U18381 (N_18381,N_18081,N_18202);
and U18382 (N_18382,N_18207,N_18170);
nor U18383 (N_18383,N_18174,N_18153);
or U18384 (N_18384,N_18210,N_18080);
and U18385 (N_18385,N_18158,N_18211);
nor U18386 (N_18386,N_18139,N_18129);
and U18387 (N_18387,N_18162,N_18122);
nand U18388 (N_18388,N_18130,N_18156);
and U18389 (N_18389,N_18110,N_18102);
and U18390 (N_18390,N_18092,N_18145);
xnor U18391 (N_18391,N_18211,N_18118);
xnor U18392 (N_18392,N_18101,N_18214);
or U18393 (N_18393,N_18181,N_18106);
and U18394 (N_18394,N_18104,N_18236);
xnor U18395 (N_18395,N_18217,N_18115);
nor U18396 (N_18396,N_18113,N_18179);
xor U18397 (N_18397,N_18128,N_18096);
or U18398 (N_18398,N_18112,N_18165);
xor U18399 (N_18399,N_18132,N_18187);
xor U18400 (N_18400,N_18261,N_18390);
nand U18401 (N_18401,N_18371,N_18285);
nand U18402 (N_18402,N_18255,N_18373);
nand U18403 (N_18403,N_18331,N_18351);
xnor U18404 (N_18404,N_18289,N_18358);
or U18405 (N_18405,N_18393,N_18372);
xor U18406 (N_18406,N_18320,N_18360);
xor U18407 (N_18407,N_18365,N_18353);
nand U18408 (N_18408,N_18333,N_18303);
or U18409 (N_18409,N_18319,N_18375);
nand U18410 (N_18410,N_18349,N_18348);
or U18411 (N_18411,N_18329,N_18296);
nor U18412 (N_18412,N_18381,N_18282);
or U18413 (N_18413,N_18369,N_18352);
and U18414 (N_18414,N_18315,N_18325);
and U18415 (N_18415,N_18362,N_18310);
and U18416 (N_18416,N_18277,N_18346);
xnor U18417 (N_18417,N_18392,N_18370);
or U18418 (N_18418,N_18355,N_18253);
or U18419 (N_18419,N_18245,N_18366);
nor U18420 (N_18420,N_18267,N_18397);
xor U18421 (N_18421,N_18269,N_18243);
nand U18422 (N_18422,N_18378,N_18260);
and U18423 (N_18423,N_18299,N_18300);
xor U18424 (N_18424,N_18385,N_18318);
or U18425 (N_18425,N_18241,N_18252);
nand U18426 (N_18426,N_18386,N_18399);
nand U18427 (N_18427,N_18270,N_18343);
and U18428 (N_18428,N_18344,N_18391);
nor U18429 (N_18429,N_18304,N_18291);
or U18430 (N_18430,N_18247,N_18395);
and U18431 (N_18431,N_18364,N_18307);
or U18432 (N_18432,N_18273,N_18271);
xor U18433 (N_18433,N_18394,N_18278);
nor U18434 (N_18434,N_18379,N_18286);
nand U18435 (N_18435,N_18264,N_18322);
nor U18436 (N_18436,N_18317,N_18292);
nor U18437 (N_18437,N_18306,N_18374);
or U18438 (N_18438,N_18330,N_18383);
xor U18439 (N_18439,N_18274,N_18313);
or U18440 (N_18440,N_18327,N_18384);
nand U18441 (N_18441,N_18335,N_18336);
or U18442 (N_18442,N_18248,N_18246);
xor U18443 (N_18443,N_18341,N_18284);
and U18444 (N_18444,N_18265,N_18263);
and U18445 (N_18445,N_18387,N_18380);
or U18446 (N_18446,N_18250,N_18262);
or U18447 (N_18447,N_18339,N_18240);
nor U18448 (N_18448,N_18398,N_18272);
nand U18449 (N_18449,N_18308,N_18316);
and U18450 (N_18450,N_18301,N_18328);
and U18451 (N_18451,N_18281,N_18279);
nor U18452 (N_18452,N_18294,N_18254);
or U18453 (N_18453,N_18314,N_18338);
nand U18454 (N_18454,N_18359,N_18361);
nor U18455 (N_18455,N_18321,N_18367);
or U18456 (N_18456,N_18340,N_18356);
xor U18457 (N_18457,N_18311,N_18244);
or U18458 (N_18458,N_18312,N_18297);
nor U18459 (N_18459,N_18287,N_18389);
xnor U18460 (N_18460,N_18293,N_18347);
nor U18461 (N_18461,N_18266,N_18376);
and U18462 (N_18462,N_18302,N_18324);
or U18463 (N_18463,N_18268,N_18332);
or U18464 (N_18464,N_18290,N_18354);
nor U18465 (N_18465,N_18257,N_18309);
nand U18466 (N_18466,N_18326,N_18345);
xnor U18467 (N_18467,N_18242,N_18334);
nand U18468 (N_18468,N_18357,N_18368);
and U18469 (N_18469,N_18288,N_18323);
and U18470 (N_18470,N_18283,N_18305);
xor U18471 (N_18471,N_18350,N_18337);
or U18472 (N_18472,N_18382,N_18258);
xor U18473 (N_18473,N_18280,N_18342);
xnor U18474 (N_18474,N_18249,N_18295);
nand U18475 (N_18475,N_18259,N_18256);
nand U18476 (N_18476,N_18363,N_18298);
and U18477 (N_18477,N_18396,N_18276);
nand U18478 (N_18478,N_18388,N_18251);
nand U18479 (N_18479,N_18275,N_18377);
or U18480 (N_18480,N_18296,N_18357);
nand U18481 (N_18481,N_18339,N_18269);
or U18482 (N_18482,N_18355,N_18270);
xnor U18483 (N_18483,N_18242,N_18349);
or U18484 (N_18484,N_18368,N_18302);
or U18485 (N_18485,N_18331,N_18327);
nor U18486 (N_18486,N_18347,N_18317);
or U18487 (N_18487,N_18344,N_18394);
xor U18488 (N_18488,N_18283,N_18370);
and U18489 (N_18489,N_18364,N_18270);
xnor U18490 (N_18490,N_18257,N_18370);
and U18491 (N_18491,N_18303,N_18251);
nor U18492 (N_18492,N_18281,N_18384);
nor U18493 (N_18493,N_18279,N_18327);
or U18494 (N_18494,N_18244,N_18363);
xnor U18495 (N_18495,N_18322,N_18245);
nand U18496 (N_18496,N_18372,N_18255);
nor U18497 (N_18497,N_18305,N_18359);
nor U18498 (N_18498,N_18244,N_18346);
nor U18499 (N_18499,N_18373,N_18396);
or U18500 (N_18500,N_18258,N_18313);
or U18501 (N_18501,N_18320,N_18283);
and U18502 (N_18502,N_18362,N_18267);
xnor U18503 (N_18503,N_18263,N_18277);
or U18504 (N_18504,N_18358,N_18335);
nor U18505 (N_18505,N_18346,N_18348);
and U18506 (N_18506,N_18384,N_18256);
or U18507 (N_18507,N_18342,N_18268);
or U18508 (N_18508,N_18373,N_18262);
or U18509 (N_18509,N_18332,N_18375);
nor U18510 (N_18510,N_18320,N_18324);
and U18511 (N_18511,N_18364,N_18295);
nand U18512 (N_18512,N_18263,N_18354);
nand U18513 (N_18513,N_18379,N_18268);
and U18514 (N_18514,N_18266,N_18287);
nor U18515 (N_18515,N_18337,N_18303);
nand U18516 (N_18516,N_18390,N_18359);
nand U18517 (N_18517,N_18312,N_18278);
nor U18518 (N_18518,N_18361,N_18267);
and U18519 (N_18519,N_18392,N_18360);
xnor U18520 (N_18520,N_18370,N_18338);
or U18521 (N_18521,N_18285,N_18311);
nor U18522 (N_18522,N_18380,N_18299);
nor U18523 (N_18523,N_18256,N_18353);
nand U18524 (N_18524,N_18256,N_18343);
and U18525 (N_18525,N_18366,N_18331);
nand U18526 (N_18526,N_18377,N_18356);
xnor U18527 (N_18527,N_18393,N_18305);
and U18528 (N_18528,N_18364,N_18396);
nand U18529 (N_18529,N_18339,N_18380);
and U18530 (N_18530,N_18393,N_18244);
or U18531 (N_18531,N_18264,N_18268);
xnor U18532 (N_18532,N_18311,N_18332);
nor U18533 (N_18533,N_18343,N_18297);
nor U18534 (N_18534,N_18242,N_18394);
nor U18535 (N_18535,N_18383,N_18276);
xor U18536 (N_18536,N_18317,N_18373);
or U18537 (N_18537,N_18324,N_18311);
xnor U18538 (N_18538,N_18390,N_18330);
and U18539 (N_18539,N_18297,N_18305);
or U18540 (N_18540,N_18343,N_18361);
and U18541 (N_18541,N_18260,N_18301);
and U18542 (N_18542,N_18367,N_18329);
nand U18543 (N_18543,N_18273,N_18329);
and U18544 (N_18544,N_18245,N_18364);
or U18545 (N_18545,N_18336,N_18359);
or U18546 (N_18546,N_18300,N_18252);
or U18547 (N_18547,N_18286,N_18251);
nand U18548 (N_18548,N_18261,N_18369);
nor U18549 (N_18549,N_18371,N_18302);
nor U18550 (N_18550,N_18249,N_18265);
nor U18551 (N_18551,N_18332,N_18286);
and U18552 (N_18552,N_18386,N_18344);
nor U18553 (N_18553,N_18345,N_18247);
xor U18554 (N_18554,N_18392,N_18256);
and U18555 (N_18555,N_18291,N_18385);
nor U18556 (N_18556,N_18321,N_18282);
and U18557 (N_18557,N_18247,N_18309);
nor U18558 (N_18558,N_18372,N_18379);
nor U18559 (N_18559,N_18328,N_18384);
xor U18560 (N_18560,N_18506,N_18541);
nor U18561 (N_18561,N_18535,N_18508);
nor U18562 (N_18562,N_18498,N_18459);
or U18563 (N_18563,N_18474,N_18478);
nor U18564 (N_18564,N_18457,N_18488);
xnor U18565 (N_18565,N_18452,N_18479);
nand U18566 (N_18566,N_18558,N_18543);
nand U18567 (N_18567,N_18511,N_18526);
nor U18568 (N_18568,N_18552,N_18524);
and U18569 (N_18569,N_18499,N_18428);
nor U18570 (N_18570,N_18418,N_18473);
nor U18571 (N_18571,N_18444,N_18548);
xor U18572 (N_18572,N_18416,N_18436);
nor U18573 (N_18573,N_18434,N_18512);
nand U18574 (N_18574,N_18469,N_18497);
nor U18575 (N_18575,N_18464,N_18447);
and U18576 (N_18576,N_18505,N_18553);
nor U18577 (N_18577,N_18441,N_18504);
xnor U18578 (N_18578,N_18432,N_18516);
nand U18579 (N_18579,N_18487,N_18521);
xnor U18580 (N_18580,N_18411,N_18422);
xnor U18581 (N_18581,N_18518,N_18491);
xnor U18582 (N_18582,N_18419,N_18415);
nand U18583 (N_18583,N_18492,N_18472);
nand U18584 (N_18584,N_18554,N_18480);
and U18585 (N_18585,N_18443,N_18510);
and U18586 (N_18586,N_18476,N_18407);
or U18587 (N_18587,N_18537,N_18470);
nand U18588 (N_18588,N_18465,N_18460);
and U18589 (N_18589,N_18523,N_18533);
or U18590 (N_18590,N_18410,N_18517);
nor U18591 (N_18591,N_18502,N_18431);
nand U18592 (N_18592,N_18536,N_18438);
and U18593 (N_18593,N_18530,N_18405);
or U18594 (N_18594,N_18453,N_18495);
and U18595 (N_18595,N_18527,N_18542);
nand U18596 (N_18596,N_18519,N_18555);
or U18597 (N_18597,N_18456,N_18556);
nor U18598 (N_18598,N_18448,N_18440);
or U18599 (N_18599,N_18403,N_18404);
nor U18600 (N_18600,N_18471,N_18449);
nor U18601 (N_18601,N_18496,N_18525);
and U18602 (N_18602,N_18461,N_18402);
nand U18603 (N_18603,N_18439,N_18509);
nand U18604 (N_18604,N_18520,N_18413);
and U18605 (N_18605,N_18489,N_18538);
or U18606 (N_18606,N_18433,N_18445);
or U18607 (N_18607,N_18514,N_18475);
or U18608 (N_18608,N_18482,N_18450);
or U18609 (N_18609,N_18559,N_18500);
xnor U18610 (N_18610,N_18545,N_18435);
nand U18611 (N_18611,N_18454,N_18484);
and U18612 (N_18612,N_18539,N_18528);
nand U18613 (N_18613,N_18406,N_18513);
nand U18614 (N_18614,N_18494,N_18425);
xnor U18615 (N_18615,N_18550,N_18507);
nand U18616 (N_18616,N_18421,N_18481);
nor U18617 (N_18617,N_18557,N_18424);
or U18618 (N_18618,N_18551,N_18451);
and U18619 (N_18619,N_18483,N_18458);
xnor U18620 (N_18620,N_18503,N_18430);
or U18621 (N_18621,N_18400,N_18544);
xnor U18622 (N_18622,N_18462,N_18463);
nand U18623 (N_18623,N_18547,N_18420);
or U18624 (N_18624,N_18515,N_18409);
and U18625 (N_18625,N_18414,N_18446);
or U18626 (N_18626,N_18546,N_18401);
xor U18627 (N_18627,N_18486,N_18417);
or U18628 (N_18628,N_18501,N_18437);
xnor U18629 (N_18629,N_18455,N_18532);
nor U18630 (N_18630,N_18426,N_18534);
nand U18631 (N_18631,N_18540,N_18493);
nor U18632 (N_18632,N_18467,N_18427);
or U18633 (N_18633,N_18477,N_18429);
nor U18634 (N_18634,N_18466,N_18468);
nand U18635 (N_18635,N_18485,N_18549);
nand U18636 (N_18636,N_18412,N_18408);
nor U18637 (N_18637,N_18529,N_18522);
or U18638 (N_18638,N_18531,N_18490);
xor U18639 (N_18639,N_18423,N_18442);
nand U18640 (N_18640,N_18456,N_18500);
nand U18641 (N_18641,N_18413,N_18465);
xor U18642 (N_18642,N_18483,N_18473);
nor U18643 (N_18643,N_18468,N_18516);
or U18644 (N_18644,N_18456,N_18416);
nand U18645 (N_18645,N_18528,N_18557);
nor U18646 (N_18646,N_18422,N_18506);
nand U18647 (N_18647,N_18506,N_18531);
xor U18648 (N_18648,N_18442,N_18448);
and U18649 (N_18649,N_18447,N_18467);
or U18650 (N_18650,N_18417,N_18497);
xnor U18651 (N_18651,N_18440,N_18519);
nor U18652 (N_18652,N_18519,N_18464);
or U18653 (N_18653,N_18533,N_18431);
xor U18654 (N_18654,N_18527,N_18457);
or U18655 (N_18655,N_18547,N_18427);
or U18656 (N_18656,N_18507,N_18527);
nor U18657 (N_18657,N_18460,N_18468);
or U18658 (N_18658,N_18484,N_18547);
xor U18659 (N_18659,N_18498,N_18441);
or U18660 (N_18660,N_18444,N_18532);
xnor U18661 (N_18661,N_18556,N_18531);
nor U18662 (N_18662,N_18431,N_18469);
nor U18663 (N_18663,N_18476,N_18485);
xor U18664 (N_18664,N_18401,N_18523);
nor U18665 (N_18665,N_18541,N_18403);
and U18666 (N_18666,N_18431,N_18549);
and U18667 (N_18667,N_18558,N_18490);
xnor U18668 (N_18668,N_18531,N_18502);
and U18669 (N_18669,N_18428,N_18464);
nand U18670 (N_18670,N_18457,N_18456);
or U18671 (N_18671,N_18438,N_18414);
nand U18672 (N_18672,N_18548,N_18482);
nor U18673 (N_18673,N_18525,N_18550);
or U18674 (N_18674,N_18470,N_18423);
and U18675 (N_18675,N_18438,N_18527);
and U18676 (N_18676,N_18455,N_18413);
nand U18677 (N_18677,N_18450,N_18447);
xnor U18678 (N_18678,N_18545,N_18412);
xnor U18679 (N_18679,N_18416,N_18547);
nor U18680 (N_18680,N_18400,N_18476);
nand U18681 (N_18681,N_18501,N_18559);
or U18682 (N_18682,N_18548,N_18484);
nand U18683 (N_18683,N_18449,N_18549);
and U18684 (N_18684,N_18433,N_18479);
xor U18685 (N_18685,N_18409,N_18483);
nor U18686 (N_18686,N_18401,N_18403);
and U18687 (N_18687,N_18458,N_18491);
nor U18688 (N_18688,N_18437,N_18486);
or U18689 (N_18689,N_18496,N_18517);
nor U18690 (N_18690,N_18524,N_18407);
and U18691 (N_18691,N_18477,N_18553);
nor U18692 (N_18692,N_18401,N_18429);
and U18693 (N_18693,N_18526,N_18457);
xnor U18694 (N_18694,N_18474,N_18443);
nand U18695 (N_18695,N_18416,N_18467);
nor U18696 (N_18696,N_18550,N_18501);
nand U18697 (N_18697,N_18436,N_18431);
xor U18698 (N_18698,N_18559,N_18558);
or U18699 (N_18699,N_18502,N_18407);
nand U18700 (N_18700,N_18434,N_18468);
nand U18701 (N_18701,N_18427,N_18506);
nor U18702 (N_18702,N_18492,N_18508);
nand U18703 (N_18703,N_18417,N_18509);
xnor U18704 (N_18704,N_18417,N_18540);
nand U18705 (N_18705,N_18480,N_18537);
and U18706 (N_18706,N_18461,N_18554);
nand U18707 (N_18707,N_18487,N_18479);
xor U18708 (N_18708,N_18520,N_18452);
xor U18709 (N_18709,N_18460,N_18413);
and U18710 (N_18710,N_18545,N_18496);
xor U18711 (N_18711,N_18456,N_18551);
xnor U18712 (N_18712,N_18411,N_18481);
nand U18713 (N_18713,N_18448,N_18432);
or U18714 (N_18714,N_18487,N_18543);
nand U18715 (N_18715,N_18481,N_18407);
nor U18716 (N_18716,N_18516,N_18520);
nand U18717 (N_18717,N_18480,N_18489);
or U18718 (N_18718,N_18434,N_18511);
or U18719 (N_18719,N_18444,N_18479);
xor U18720 (N_18720,N_18680,N_18684);
xor U18721 (N_18721,N_18631,N_18625);
nand U18722 (N_18722,N_18622,N_18705);
xnor U18723 (N_18723,N_18587,N_18706);
or U18724 (N_18724,N_18681,N_18669);
nand U18725 (N_18725,N_18651,N_18656);
nand U18726 (N_18726,N_18613,N_18593);
nand U18727 (N_18727,N_18702,N_18606);
nand U18728 (N_18728,N_18576,N_18650);
or U18729 (N_18729,N_18608,N_18621);
xor U18730 (N_18730,N_18575,N_18662);
and U18731 (N_18731,N_18670,N_18668);
nor U18732 (N_18732,N_18629,N_18619);
xnor U18733 (N_18733,N_18663,N_18682);
nand U18734 (N_18734,N_18607,N_18704);
or U18735 (N_18735,N_18646,N_18626);
nand U18736 (N_18736,N_18692,N_18661);
and U18737 (N_18737,N_18640,N_18644);
xor U18738 (N_18738,N_18584,N_18602);
nand U18739 (N_18739,N_18641,N_18591);
nor U18740 (N_18740,N_18636,N_18701);
nor U18741 (N_18741,N_18601,N_18717);
xnor U18742 (N_18742,N_18686,N_18620);
or U18743 (N_18743,N_18696,N_18594);
or U18744 (N_18744,N_18562,N_18719);
nor U18745 (N_18745,N_18715,N_18618);
nand U18746 (N_18746,N_18609,N_18655);
nand U18747 (N_18747,N_18694,N_18679);
and U18748 (N_18748,N_18707,N_18561);
and U18749 (N_18749,N_18647,N_18642);
or U18750 (N_18750,N_18718,N_18600);
xor U18751 (N_18751,N_18638,N_18590);
and U18752 (N_18752,N_18627,N_18634);
or U18753 (N_18753,N_18581,N_18676);
xor U18754 (N_18754,N_18599,N_18716);
and U18755 (N_18755,N_18699,N_18712);
or U18756 (N_18756,N_18632,N_18714);
and U18757 (N_18757,N_18643,N_18582);
xor U18758 (N_18758,N_18672,N_18691);
nor U18759 (N_18759,N_18586,N_18637);
nand U18760 (N_18760,N_18580,N_18579);
nand U18761 (N_18761,N_18614,N_18571);
xnor U18762 (N_18762,N_18578,N_18595);
nor U18763 (N_18763,N_18604,N_18567);
or U18764 (N_18764,N_18572,N_18658);
and U18765 (N_18765,N_18564,N_18583);
nand U18766 (N_18766,N_18711,N_18574);
or U18767 (N_18767,N_18566,N_18603);
or U18768 (N_18768,N_18703,N_18624);
nor U18769 (N_18769,N_18652,N_18563);
and U18770 (N_18770,N_18639,N_18673);
or U18771 (N_18771,N_18597,N_18685);
nor U18772 (N_18772,N_18577,N_18654);
or U18773 (N_18773,N_18596,N_18617);
xor U18774 (N_18774,N_18565,N_18630);
xor U18775 (N_18775,N_18678,N_18611);
or U18776 (N_18776,N_18615,N_18677);
nand U18777 (N_18777,N_18589,N_18687);
xor U18778 (N_18778,N_18612,N_18688);
nor U18779 (N_18779,N_18709,N_18695);
xnor U18780 (N_18780,N_18635,N_18648);
or U18781 (N_18781,N_18659,N_18623);
and U18782 (N_18782,N_18666,N_18698);
or U18783 (N_18783,N_18653,N_18660);
nand U18784 (N_18784,N_18675,N_18585);
and U18785 (N_18785,N_18697,N_18689);
or U18786 (N_18786,N_18610,N_18700);
nand U18787 (N_18787,N_18693,N_18560);
xor U18788 (N_18788,N_18573,N_18690);
nand U18789 (N_18789,N_18671,N_18633);
and U18790 (N_18790,N_18665,N_18569);
nand U18791 (N_18791,N_18649,N_18605);
and U18792 (N_18792,N_18568,N_18598);
nand U18793 (N_18793,N_18710,N_18570);
nand U18794 (N_18794,N_18667,N_18657);
nor U18795 (N_18795,N_18713,N_18616);
or U18796 (N_18796,N_18683,N_18708);
nor U18797 (N_18797,N_18664,N_18674);
nor U18798 (N_18798,N_18628,N_18588);
nand U18799 (N_18799,N_18645,N_18592);
or U18800 (N_18800,N_18700,N_18698);
nand U18801 (N_18801,N_18583,N_18619);
and U18802 (N_18802,N_18578,N_18679);
nand U18803 (N_18803,N_18719,N_18602);
xnor U18804 (N_18804,N_18705,N_18593);
xor U18805 (N_18805,N_18562,N_18570);
xnor U18806 (N_18806,N_18616,N_18597);
xnor U18807 (N_18807,N_18591,N_18633);
nand U18808 (N_18808,N_18596,N_18591);
nor U18809 (N_18809,N_18615,N_18675);
or U18810 (N_18810,N_18649,N_18716);
and U18811 (N_18811,N_18642,N_18704);
or U18812 (N_18812,N_18623,N_18597);
nor U18813 (N_18813,N_18606,N_18653);
nor U18814 (N_18814,N_18638,N_18674);
xnor U18815 (N_18815,N_18685,N_18699);
nand U18816 (N_18816,N_18624,N_18607);
nand U18817 (N_18817,N_18697,N_18674);
nand U18818 (N_18818,N_18695,N_18689);
or U18819 (N_18819,N_18605,N_18716);
xor U18820 (N_18820,N_18597,N_18665);
and U18821 (N_18821,N_18702,N_18716);
nor U18822 (N_18822,N_18574,N_18704);
nand U18823 (N_18823,N_18567,N_18575);
xnor U18824 (N_18824,N_18573,N_18654);
xor U18825 (N_18825,N_18583,N_18575);
nand U18826 (N_18826,N_18634,N_18621);
and U18827 (N_18827,N_18603,N_18576);
nand U18828 (N_18828,N_18632,N_18577);
or U18829 (N_18829,N_18594,N_18625);
and U18830 (N_18830,N_18703,N_18570);
or U18831 (N_18831,N_18629,N_18566);
nor U18832 (N_18832,N_18677,N_18578);
or U18833 (N_18833,N_18574,N_18644);
xnor U18834 (N_18834,N_18576,N_18679);
and U18835 (N_18835,N_18577,N_18663);
xnor U18836 (N_18836,N_18640,N_18695);
nand U18837 (N_18837,N_18637,N_18645);
or U18838 (N_18838,N_18696,N_18595);
and U18839 (N_18839,N_18717,N_18631);
nor U18840 (N_18840,N_18651,N_18684);
nand U18841 (N_18841,N_18623,N_18572);
nand U18842 (N_18842,N_18634,N_18563);
and U18843 (N_18843,N_18599,N_18589);
or U18844 (N_18844,N_18563,N_18660);
nand U18845 (N_18845,N_18585,N_18586);
and U18846 (N_18846,N_18682,N_18571);
nor U18847 (N_18847,N_18685,N_18586);
nor U18848 (N_18848,N_18615,N_18689);
and U18849 (N_18849,N_18577,N_18587);
nand U18850 (N_18850,N_18673,N_18667);
or U18851 (N_18851,N_18668,N_18661);
xor U18852 (N_18852,N_18604,N_18656);
nor U18853 (N_18853,N_18663,N_18701);
xnor U18854 (N_18854,N_18657,N_18578);
nor U18855 (N_18855,N_18691,N_18595);
nor U18856 (N_18856,N_18643,N_18661);
nor U18857 (N_18857,N_18670,N_18667);
or U18858 (N_18858,N_18646,N_18610);
and U18859 (N_18859,N_18633,N_18605);
xor U18860 (N_18860,N_18704,N_18584);
or U18861 (N_18861,N_18674,N_18651);
nand U18862 (N_18862,N_18563,N_18655);
or U18863 (N_18863,N_18561,N_18677);
xor U18864 (N_18864,N_18618,N_18565);
xor U18865 (N_18865,N_18688,N_18576);
and U18866 (N_18866,N_18624,N_18657);
nand U18867 (N_18867,N_18661,N_18575);
nor U18868 (N_18868,N_18700,N_18618);
xnor U18869 (N_18869,N_18697,N_18635);
nand U18870 (N_18870,N_18641,N_18701);
nand U18871 (N_18871,N_18593,N_18629);
or U18872 (N_18872,N_18700,N_18625);
nor U18873 (N_18873,N_18608,N_18579);
nor U18874 (N_18874,N_18701,N_18682);
xor U18875 (N_18875,N_18714,N_18605);
or U18876 (N_18876,N_18696,N_18713);
and U18877 (N_18877,N_18621,N_18638);
or U18878 (N_18878,N_18568,N_18713);
nand U18879 (N_18879,N_18694,N_18574);
or U18880 (N_18880,N_18773,N_18766);
nand U18881 (N_18881,N_18774,N_18803);
or U18882 (N_18882,N_18750,N_18762);
nand U18883 (N_18883,N_18844,N_18863);
nand U18884 (N_18884,N_18874,N_18813);
or U18885 (N_18885,N_18824,N_18816);
nor U18886 (N_18886,N_18833,N_18777);
xnor U18887 (N_18887,N_18806,N_18815);
or U18888 (N_18888,N_18879,N_18834);
nor U18889 (N_18889,N_18760,N_18842);
and U18890 (N_18890,N_18846,N_18753);
nor U18891 (N_18891,N_18723,N_18866);
or U18892 (N_18892,N_18862,N_18763);
and U18893 (N_18893,N_18852,N_18828);
nor U18894 (N_18894,N_18741,N_18822);
nand U18895 (N_18895,N_18821,N_18738);
nand U18896 (N_18896,N_18872,N_18758);
and U18897 (N_18897,N_18751,N_18857);
or U18898 (N_18898,N_18817,N_18840);
nand U18899 (N_18899,N_18726,N_18819);
xnor U18900 (N_18900,N_18870,N_18849);
xnor U18901 (N_18901,N_18848,N_18865);
nand U18902 (N_18902,N_18804,N_18827);
or U18903 (N_18903,N_18755,N_18838);
or U18904 (N_18904,N_18859,N_18791);
and U18905 (N_18905,N_18761,N_18858);
xor U18906 (N_18906,N_18798,N_18770);
nor U18907 (N_18907,N_18787,N_18783);
and U18908 (N_18908,N_18793,N_18797);
or U18909 (N_18909,N_18745,N_18794);
nand U18910 (N_18910,N_18802,N_18731);
and U18911 (N_18911,N_18744,N_18854);
and U18912 (N_18912,N_18811,N_18767);
nand U18913 (N_18913,N_18868,N_18748);
or U18914 (N_18914,N_18869,N_18876);
xor U18915 (N_18915,N_18784,N_18743);
and U18916 (N_18916,N_18847,N_18807);
and U18917 (N_18917,N_18836,N_18775);
nor U18918 (N_18918,N_18769,N_18855);
nand U18919 (N_18919,N_18864,N_18809);
and U18920 (N_18920,N_18764,N_18754);
and U18921 (N_18921,N_18837,N_18850);
and U18922 (N_18922,N_18782,N_18832);
and U18923 (N_18923,N_18779,N_18768);
or U18924 (N_18924,N_18856,N_18825);
or U18925 (N_18925,N_18877,N_18772);
nand U18926 (N_18926,N_18737,N_18800);
or U18927 (N_18927,N_18878,N_18722);
or U18928 (N_18928,N_18725,N_18788);
nand U18929 (N_18929,N_18795,N_18752);
or U18930 (N_18930,N_18786,N_18720);
xnor U18931 (N_18931,N_18746,N_18778);
or U18932 (N_18932,N_18873,N_18812);
xor U18933 (N_18933,N_18831,N_18867);
and U18934 (N_18934,N_18818,N_18721);
and U18935 (N_18935,N_18739,N_18823);
or U18936 (N_18936,N_18829,N_18727);
or U18937 (N_18937,N_18742,N_18771);
or U18938 (N_18938,N_18765,N_18853);
nand U18939 (N_18939,N_18736,N_18810);
and U18940 (N_18940,N_18756,N_18728);
xnor U18941 (N_18941,N_18814,N_18801);
and U18942 (N_18942,N_18733,N_18820);
and U18943 (N_18943,N_18860,N_18730);
xnor U18944 (N_18944,N_18759,N_18826);
xnor U18945 (N_18945,N_18796,N_18740);
nand U18946 (N_18946,N_18747,N_18749);
and U18947 (N_18947,N_18808,N_18789);
and U18948 (N_18948,N_18732,N_18781);
nor U18949 (N_18949,N_18792,N_18757);
and U18950 (N_18950,N_18871,N_18729);
nand U18951 (N_18951,N_18799,N_18839);
or U18952 (N_18952,N_18735,N_18785);
and U18953 (N_18953,N_18805,N_18790);
xnor U18954 (N_18954,N_18835,N_18845);
xor U18955 (N_18955,N_18734,N_18851);
and U18956 (N_18956,N_18724,N_18875);
nand U18957 (N_18957,N_18830,N_18861);
and U18958 (N_18958,N_18780,N_18776);
or U18959 (N_18959,N_18841,N_18843);
or U18960 (N_18960,N_18878,N_18773);
nor U18961 (N_18961,N_18850,N_18733);
nor U18962 (N_18962,N_18844,N_18736);
and U18963 (N_18963,N_18843,N_18824);
or U18964 (N_18964,N_18870,N_18802);
and U18965 (N_18965,N_18784,N_18773);
and U18966 (N_18966,N_18838,N_18776);
nor U18967 (N_18967,N_18736,N_18740);
and U18968 (N_18968,N_18820,N_18848);
nand U18969 (N_18969,N_18833,N_18850);
nand U18970 (N_18970,N_18835,N_18722);
nor U18971 (N_18971,N_18732,N_18794);
xor U18972 (N_18972,N_18809,N_18808);
and U18973 (N_18973,N_18772,N_18827);
xnor U18974 (N_18974,N_18851,N_18874);
nor U18975 (N_18975,N_18866,N_18804);
nor U18976 (N_18976,N_18796,N_18752);
nand U18977 (N_18977,N_18739,N_18786);
xnor U18978 (N_18978,N_18754,N_18770);
xnor U18979 (N_18979,N_18795,N_18824);
nor U18980 (N_18980,N_18825,N_18768);
or U18981 (N_18981,N_18723,N_18764);
or U18982 (N_18982,N_18786,N_18811);
and U18983 (N_18983,N_18823,N_18839);
nand U18984 (N_18984,N_18812,N_18805);
nand U18985 (N_18985,N_18821,N_18798);
xor U18986 (N_18986,N_18798,N_18759);
nor U18987 (N_18987,N_18767,N_18728);
nand U18988 (N_18988,N_18844,N_18826);
nor U18989 (N_18989,N_18829,N_18871);
nor U18990 (N_18990,N_18800,N_18837);
and U18991 (N_18991,N_18837,N_18844);
nor U18992 (N_18992,N_18730,N_18752);
or U18993 (N_18993,N_18831,N_18725);
or U18994 (N_18994,N_18869,N_18809);
or U18995 (N_18995,N_18759,N_18823);
nor U18996 (N_18996,N_18843,N_18779);
xor U18997 (N_18997,N_18854,N_18846);
xnor U18998 (N_18998,N_18751,N_18823);
or U18999 (N_18999,N_18757,N_18799);
nand U19000 (N_19000,N_18874,N_18763);
nand U19001 (N_19001,N_18840,N_18788);
nand U19002 (N_19002,N_18796,N_18721);
or U19003 (N_19003,N_18825,N_18817);
and U19004 (N_19004,N_18732,N_18782);
xnor U19005 (N_19005,N_18801,N_18749);
or U19006 (N_19006,N_18878,N_18801);
xor U19007 (N_19007,N_18867,N_18848);
or U19008 (N_19008,N_18809,N_18842);
and U19009 (N_19009,N_18813,N_18847);
xor U19010 (N_19010,N_18831,N_18726);
and U19011 (N_19011,N_18767,N_18731);
nand U19012 (N_19012,N_18759,N_18830);
or U19013 (N_19013,N_18764,N_18822);
nor U19014 (N_19014,N_18806,N_18822);
or U19015 (N_19015,N_18810,N_18850);
nor U19016 (N_19016,N_18759,N_18735);
nand U19017 (N_19017,N_18871,N_18727);
and U19018 (N_19018,N_18840,N_18874);
and U19019 (N_19019,N_18808,N_18735);
nand U19020 (N_19020,N_18859,N_18757);
xor U19021 (N_19021,N_18785,N_18813);
nand U19022 (N_19022,N_18808,N_18742);
or U19023 (N_19023,N_18741,N_18868);
xnor U19024 (N_19024,N_18785,N_18809);
and U19025 (N_19025,N_18848,N_18728);
or U19026 (N_19026,N_18739,N_18801);
nand U19027 (N_19027,N_18809,N_18833);
and U19028 (N_19028,N_18865,N_18777);
xor U19029 (N_19029,N_18825,N_18844);
xnor U19030 (N_19030,N_18730,N_18794);
xnor U19031 (N_19031,N_18723,N_18805);
or U19032 (N_19032,N_18736,N_18787);
and U19033 (N_19033,N_18761,N_18865);
and U19034 (N_19034,N_18855,N_18852);
nor U19035 (N_19035,N_18792,N_18827);
nand U19036 (N_19036,N_18752,N_18760);
or U19037 (N_19037,N_18860,N_18752);
or U19038 (N_19038,N_18775,N_18739);
xnor U19039 (N_19039,N_18828,N_18772);
and U19040 (N_19040,N_19002,N_18991);
xnor U19041 (N_19041,N_19013,N_18929);
xnor U19042 (N_19042,N_18919,N_18901);
nand U19043 (N_19043,N_19024,N_18926);
xor U19044 (N_19044,N_18943,N_18935);
nor U19045 (N_19045,N_18913,N_18882);
xor U19046 (N_19046,N_18976,N_19022);
xor U19047 (N_19047,N_18973,N_18980);
xor U19048 (N_19048,N_19027,N_18992);
nand U19049 (N_19049,N_18881,N_18938);
nand U19050 (N_19050,N_18995,N_18896);
and U19051 (N_19051,N_18887,N_18956);
and U19052 (N_19052,N_18888,N_18936);
or U19053 (N_19053,N_18978,N_18904);
and U19054 (N_19054,N_18898,N_18931);
nor U19055 (N_19055,N_18903,N_19011);
nor U19056 (N_19056,N_18955,N_18883);
xnor U19057 (N_19057,N_18967,N_18975);
nand U19058 (N_19058,N_18905,N_18994);
nand U19059 (N_19059,N_18968,N_19030);
nor U19060 (N_19060,N_18998,N_18884);
and U19061 (N_19061,N_19033,N_19001);
and U19062 (N_19062,N_19003,N_19004);
xor U19063 (N_19063,N_18963,N_18894);
or U19064 (N_19064,N_18969,N_18880);
xnor U19065 (N_19065,N_18974,N_18893);
nand U19066 (N_19066,N_18902,N_18939);
xnor U19067 (N_19067,N_19026,N_18910);
xor U19068 (N_19068,N_19007,N_18941);
xor U19069 (N_19069,N_19035,N_18915);
nor U19070 (N_19070,N_19029,N_18911);
nand U19071 (N_19071,N_18972,N_18927);
nor U19072 (N_19072,N_18920,N_18957);
or U19073 (N_19073,N_18890,N_18988);
nor U19074 (N_19074,N_18959,N_18908);
xor U19075 (N_19075,N_18899,N_18924);
and U19076 (N_19076,N_18989,N_18891);
nor U19077 (N_19077,N_18987,N_19038);
nand U19078 (N_19078,N_18949,N_18946);
xor U19079 (N_19079,N_19037,N_19018);
nor U19080 (N_19080,N_18934,N_18960);
nor U19081 (N_19081,N_18990,N_18909);
nor U19082 (N_19082,N_18951,N_18954);
nor U19083 (N_19083,N_19031,N_18886);
nor U19084 (N_19084,N_18921,N_18885);
and U19085 (N_19085,N_19010,N_18983);
and U19086 (N_19086,N_18982,N_18922);
and U19087 (N_19087,N_19014,N_18965);
nand U19088 (N_19088,N_18979,N_18952);
xor U19089 (N_19089,N_18916,N_18925);
nor U19090 (N_19090,N_19028,N_19017);
and U19091 (N_19091,N_18897,N_18977);
xnor U19092 (N_19092,N_18999,N_18942);
or U19093 (N_19093,N_19023,N_18970);
or U19094 (N_19094,N_19032,N_18907);
and U19095 (N_19095,N_19009,N_19015);
nor U19096 (N_19096,N_18906,N_19036);
xnor U19097 (N_19097,N_18997,N_18895);
nand U19098 (N_19098,N_18986,N_18950);
and U19099 (N_19099,N_19021,N_18964);
nand U19100 (N_19100,N_18917,N_18930);
or U19101 (N_19101,N_18996,N_19034);
or U19102 (N_19102,N_18914,N_18923);
or U19103 (N_19103,N_18944,N_19016);
nor U19104 (N_19104,N_18928,N_18984);
and U19105 (N_19105,N_18985,N_18892);
and U19106 (N_19106,N_18971,N_18961);
nor U19107 (N_19107,N_19008,N_19039);
or U19108 (N_19108,N_19012,N_18937);
nand U19109 (N_19109,N_18912,N_18889);
nor U19110 (N_19110,N_18958,N_19000);
nor U19111 (N_19111,N_18933,N_18948);
xnor U19112 (N_19112,N_18932,N_19025);
xnor U19113 (N_19113,N_18993,N_18953);
nor U19114 (N_19114,N_18981,N_18900);
and U19115 (N_19115,N_18966,N_18940);
nor U19116 (N_19116,N_18918,N_19020);
and U19117 (N_19117,N_18947,N_19005);
xnor U19118 (N_19118,N_19006,N_18962);
and U19119 (N_19119,N_19019,N_18945);
nand U19120 (N_19120,N_19036,N_18956);
nor U19121 (N_19121,N_19035,N_19013);
xnor U19122 (N_19122,N_18887,N_18919);
or U19123 (N_19123,N_18881,N_18894);
nand U19124 (N_19124,N_19039,N_18919);
and U19125 (N_19125,N_18991,N_18962);
and U19126 (N_19126,N_18977,N_18912);
nor U19127 (N_19127,N_18927,N_19017);
nand U19128 (N_19128,N_18945,N_18980);
or U19129 (N_19129,N_18931,N_18890);
xor U19130 (N_19130,N_19006,N_19032);
and U19131 (N_19131,N_18972,N_18978);
and U19132 (N_19132,N_18968,N_18910);
xnor U19133 (N_19133,N_18984,N_18890);
and U19134 (N_19134,N_19036,N_18957);
or U19135 (N_19135,N_18940,N_18882);
xnor U19136 (N_19136,N_18905,N_18961);
xor U19137 (N_19137,N_19020,N_19037);
or U19138 (N_19138,N_18925,N_18953);
nor U19139 (N_19139,N_18960,N_18963);
and U19140 (N_19140,N_18965,N_19039);
nor U19141 (N_19141,N_18896,N_18968);
nor U19142 (N_19142,N_18883,N_18936);
and U19143 (N_19143,N_19030,N_18896);
nand U19144 (N_19144,N_18914,N_18955);
nor U19145 (N_19145,N_18941,N_18991);
or U19146 (N_19146,N_18888,N_19033);
and U19147 (N_19147,N_18928,N_18995);
nor U19148 (N_19148,N_18892,N_18913);
or U19149 (N_19149,N_18999,N_18938);
xnor U19150 (N_19150,N_18906,N_19012);
xor U19151 (N_19151,N_18933,N_18955);
nand U19152 (N_19152,N_18955,N_19014);
or U19153 (N_19153,N_18886,N_19026);
and U19154 (N_19154,N_18924,N_19001);
or U19155 (N_19155,N_18921,N_18977);
or U19156 (N_19156,N_18880,N_19000);
nor U19157 (N_19157,N_18918,N_19038);
and U19158 (N_19158,N_18934,N_18905);
nand U19159 (N_19159,N_18998,N_18953);
and U19160 (N_19160,N_19024,N_18963);
xor U19161 (N_19161,N_18981,N_18957);
and U19162 (N_19162,N_18881,N_18961);
xor U19163 (N_19163,N_19015,N_19008);
or U19164 (N_19164,N_18944,N_19039);
xor U19165 (N_19165,N_18888,N_19000);
nor U19166 (N_19166,N_18998,N_18971);
and U19167 (N_19167,N_18959,N_18939);
or U19168 (N_19168,N_18991,N_18969);
nor U19169 (N_19169,N_18925,N_18917);
and U19170 (N_19170,N_18918,N_18983);
and U19171 (N_19171,N_18988,N_18973);
nand U19172 (N_19172,N_18923,N_18980);
or U19173 (N_19173,N_19027,N_18967);
nand U19174 (N_19174,N_18928,N_19029);
xor U19175 (N_19175,N_18963,N_18948);
nor U19176 (N_19176,N_18900,N_19023);
or U19177 (N_19177,N_18974,N_18982);
xnor U19178 (N_19178,N_18899,N_18967);
xor U19179 (N_19179,N_18959,N_18997);
nand U19180 (N_19180,N_18885,N_18926);
xor U19181 (N_19181,N_18903,N_18926);
and U19182 (N_19182,N_19030,N_18962);
nor U19183 (N_19183,N_18973,N_18923);
or U19184 (N_19184,N_18954,N_19034);
xnor U19185 (N_19185,N_18931,N_18954);
or U19186 (N_19186,N_18950,N_19036);
xor U19187 (N_19187,N_18976,N_18958);
xor U19188 (N_19188,N_18931,N_18996);
nor U19189 (N_19189,N_18943,N_18946);
nand U19190 (N_19190,N_18909,N_18985);
and U19191 (N_19191,N_18912,N_19026);
and U19192 (N_19192,N_19013,N_19032);
or U19193 (N_19193,N_18949,N_18882);
xor U19194 (N_19194,N_18960,N_19008);
xor U19195 (N_19195,N_18926,N_18893);
nand U19196 (N_19196,N_18902,N_19016);
nand U19197 (N_19197,N_18952,N_19009);
nor U19198 (N_19198,N_18994,N_18985);
xnor U19199 (N_19199,N_18977,N_18956);
xnor U19200 (N_19200,N_19181,N_19151);
xnor U19201 (N_19201,N_19103,N_19086);
and U19202 (N_19202,N_19043,N_19067);
nand U19203 (N_19203,N_19112,N_19114);
and U19204 (N_19204,N_19052,N_19196);
or U19205 (N_19205,N_19191,N_19141);
and U19206 (N_19206,N_19128,N_19069);
and U19207 (N_19207,N_19070,N_19131);
or U19208 (N_19208,N_19090,N_19146);
and U19209 (N_19209,N_19168,N_19138);
xnor U19210 (N_19210,N_19197,N_19136);
nand U19211 (N_19211,N_19099,N_19186);
nand U19212 (N_19212,N_19057,N_19192);
or U19213 (N_19213,N_19120,N_19174);
nand U19214 (N_19214,N_19078,N_19180);
xor U19215 (N_19215,N_19049,N_19132);
xor U19216 (N_19216,N_19088,N_19163);
xnor U19217 (N_19217,N_19087,N_19139);
and U19218 (N_19218,N_19188,N_19123);
nor U19219 (N_19219,N_19195,N_19056);
nor U19220 (N_19220,N_19071,N_19082);
nand U19221 (N_19221,N_19077,N_19104);
xor U19222 (N_19222,N_19142,N_19182);
and U19223 (N_19223,N_19170,N_19100);
xnor U19224 (N_19224,N_19059,N_19083);
or U19225 (N_19225,N_19045,N_19165);
xnor U19226 (N_19226,N_19084,N_19183);
nand U19227 (N_19227,N_19058,N_19064);
or U19228 (N_19228,N_19193,N_19137);
xor U19229 (N_19229,N_19166,N_19135);
nor U19230 (N_19230,N_19089,N_19042);
xnor U19231 (N_19231,N_19062,N_19060);
xor U19232 (N_19232,N_19092,N_19157);
and U19233 (N_19233,N_19143,N_19164);
nor U19234 (N_19234,N_19073,N_19096);
nand U19235 (N_19235,N_19079,N_19047);
xnor U19236 (N_19236,N_19050,N_19162);
xor U19237 (N_19237,N_19121,N_19097);
and U19238 (N_19238,N_19110,N_19179);
and U19239 (N_19239,N_19101,N_19172);
or U19240 (N_19240,N_19159,N_19115);
and U19241 (N_19241,N_19040,N_19080);
xnor U19242 (N_19242,N_19061,N_19148);
or U19243 (N_19243,N_19055,N_19178);
or U19244 (N_19244,N_19169,N_19154);
or U19245 (N_19245,N_19187,N_19065);
and U19246 (N_19246,N_19063,N_19108);
nand U19247 (N_19247,N_19130,N_19118);
nand U19248 (N_19248,N_19107,N_19152);
and U19249 (N_19249,N_19140,N_19167);
nor U19250 (N_19250,N_19176,N_19093);
and U19251 (N_19251,N_19075,N_19051);
nand U19252 (N_19252,N_19046,N_19113);
nor U19253 (N_19253,N_19158,N_19145);
nor U19254 (N_19254,N_19127,N_19124);
nand U19255 (N_19255,N_19129,N_19199);
xor U19256 (N_19256,N_19091,N_19044);
or U19257 (N_19257,N_19102,N_19161);
and U19258 (N_19258,N_19048,N_19122);
nand U19259 (N_19259,N_19076,N_19177);
nand U19260 (N_19260,N_19125,N_19153);
or U19261 (N_19261,N_19111,N_19119);
nand U19262 (N_19262,N_19150,N_19155);
or U19263 (N_19263,N_19149,N_19184);
xor U19264 (N_19264,N_19134,N_19185);
xor U19265 (N_19265,N_19106,N_19041);
nand U19266 (N_19266,N_19160,N_19081);
or U19267 (N_19267,N_19053,N_19173);
xor U19268 (N_19268,N_19094,N_19116);
and U19269 (N_19269,N_19171,N_19198);
xnor U19270 (N_19270,N_19109,N_19072);
and U19271 (N_19271,N_19117,N_19126);
nor U19272 (N_19272,N_19085,N_19066);
or U19273 (N_19273,N_19054,N_19105);
or U19274 (N_19274,N_19147,N_19095);
and U19275 (N_19275,N_19156,N_19144);
nor U19276 (N_19276,N_19189,N_19074);
xnor U19277 (N_19277,N_19194,N_19175);
xor U19278 (N_19278,N_19190,N_19133);
or U19279 (N_19279,N_19098,N_19068);
nand U19280 (N_19280,N_19049,N_19145);
nor U19281 (N_19281,N_19098,N_19074);
xor U19282 (N_19282,N_19119,N_19116);
and U19283 (N_19283,N_19161,N_19068);
nand U19284 (N_19284,N_19053,N_19179);
and U19285 (N_19285,N_19178,N_19070);
nand U19286 (N_19286,N_19194,N_19124);
nor U19287 (N_19287,N_19181,N_19124);
nor U19288 (N_19288,N_19143,N_19057);
or U19289 (N_19289,N_19041,N_19070);
xnor U19290 (N_19290,N_19116,N_19054);
nor U19291 (N_19291,N_19096,N_19049);
nor U19292 (N_19292,N_19049,N_19042);
nand U19293 (N_19293,N_19159,N_19117);
nor U19294 (N_19294,N_19088,N_19118);
xnor U19295 (N_19295,N_19045,N_19043);
and U19296 (N_19296,N_19164,N_19092);
nand U19297 (N_19297,N_19099,N_19095);
and U19298 (N_19298,N_19151,N_19166);
nand U19299 (N_19299,N_19110,N_19067);
nand U19300 (N_19300,N_19062,N_19116);
xnor U19301 (N_19301,N_19096,N_19192);
nand U19302 (N_19302,N_19169,N_19051);
or U19303 (N_19303,N_19073,N_19117);
nor U19304 (N_19304,N_19119,N_19042);
nor U19305 (N_19305,N_19141,N_19080);
or U19306 (N_19306,N_19110,N_19141);
xor U19307 (N_19307,N_19197,N_19123);
nand U19308 (N_19308,N_19128,N_19136);
nor U19309 (N_19309,N_19163,N_19135);
or U19310 (N_19310,N_19150,N_19071);
xor U19311 (N_19311,N_19177,N_19102);
or U19312 (N_19312,N_19148,N_19147);
or U19313 (N_19313,N_19145,N_19198);
nor U19314 (N_19314,N_19195,N_19147);
nand U19315 (N_19315,N_19151,N_19130);
nor U19316 (N_19316,N_19162,N_19078);
xor U19317 (N_19317,N_19152,N_19191);
or U19318 (N_19318,N_19054,N_19127);
nor U19319 (N_19319,N_19115,N_19095);
xor U19320 (N_19320,N_19193,N_19196);
and U19321 (N_19321,N_19171,N_19191);
nand U19322 (N_19322,N_19153,N_19170);
nor U19323 (N_19323,N_19055,N_19100);
xor U19324 (N_19324,N_19078,N_19097);
or U19325 (N_19325,N_19122,N_19110);
and U19326 (N_19326,N_19145,N_19056);
nor U19327 (N_19327,N_19166,N_19099);
nand U19328 (N_19328,N_19159,N_19089);
xnor U19329 (N_19329,N_19068,N_19191);
xnor U19330 (N_19330,N_19070,N_19094);
or U19331 (N_19331,N_19106,N_19162);
nand U19332 (N_19332,N_19150,N_19104);
and U19333 (N_19333,N_19067,N_19186);
or U19334 (N_19334,N_19189,N_19041);
xnor U19335 (N_19335,N_19158,N_19042);
or U19336 (N_19336,N_19090,N_19116);
or U19337 (N_19337,N_19072,N_19135);
xor U19338 (N_19338,N_19124,N_19147);
nand U19339 (N_19339,N_19130,N_19099);
and U19340 (N_19340,N_19176,N_19067);
and U19341 (N_19341,N_19139,N_19083);
and U19342 (N_19342,N_19135,N_19190);
nor U19343 (N_19343,N_19041,N_19085);
nand U19344 (N_19344,N_19128,N_19137);
or U19345 (N_19345,N_19083,N_19051);
nand U19346 (N_19346,N_19049,N_19118);
nor U19347 (N_19347,N_19156,N_19197);
and U19348 (N_19348,N_19133,N_19106);
xor U19349 (N_19349,N_19101,N_19115);
nor U19350 (N_19350,N_19151,N_19137);
nand U19351 (N_19351,N_19132,N_19097);
or U19352 (N_19352,N_19154,N_19182);
or U19353 (N_19353,N_19148,N_19082);
and U19354 (N_19354,N_19121,N_19115);
nand U19355 (N_19355,N_19066,N_19143);
nor U19356 (N_19356,N_19106,N_19125);
xor U19357 (N_19357,N_19197,N_19142);
xor U19358 (N_19358,N_19168,N_19131);
nor U19359 (N_19359,N_19067,N_19095);
xnor U19360 (N_19360,N_19234,N_19286);
xor U19361 (N_19361,N_19252,N_19248);
or U19362 (N_19362,N_19222,N_19262);
or U19363 (N_19363,N_19269,N_19202);
xnor U19364 (N_19364,N_19214,N_19245);
nor U19365 (N_19365,N_19275,N_19350);
nor U19366 (N_19366,N_19201,N_19358);
xor U19367 (N_19367,N_19221,N_19302);
and U19368 (N_19368,N_19355,N_19329);
nor U19369 (N_19369,N_19328,N_19227);
and U19370 (N_19370,N_19289,N_19232);
or U19371 (N_19371,N_19346,N_19265);
nor U19372 (N_19372,N_19313,N_19307);
and U19373 (N_19373,N_19247,N_19240);
xnor U19374 (N_19374,N_19334,N_19229);
nor U19375 (N_19375,N_19238,N_19354);
nand U19376 (N_19376,N_19284,N_19263);
nor U19377 (N_19377,N_19276,N_19320);
nor U19378 (N_19378,N_19339,N_19255);
and U19379 (N_19379,N_19306,N_19220);
and U19380 (N_19380,N_19359,N_19231);
or U19381 (N_19381,N_19314,N_19312);
xor U19382 (N_19382,N_19260,N_19213);
or U19383 (N_19383,N_19356,N_19283);
and U19384 (N_19384,N_19341,N_19315);
or U19385 (N_19385,N_19282,N_19218);
nor U19386 (N_19386,N_19310,N_19239);
xor U19387 (N_19387,N_19215,N_19281);
nor U19388 (N_19388,N_19223,N_19323);
nor U19389 (N_19389,N_19216,N_19249);
or U19390 (N_19390,N_19309,N_19298);
xnor U19391 (N_19391,N_19330,N_19204);
xnor U19392 (N_19392,N_19272,N_19219);
or U19393 (N_19393,N_19333,N_19287);
nor U19394 (N_19394,N_19321,N_19357);
or U19395 (N_19395,N_19319,N_19261);
and U19396 (N_19396,N_19268,N_19208);
or U19397 (N_19397,N_19226,N_19308);
nand U19398 (N_19398,N_19278,N_19300);
nor U19399 (N_19399,N_19203,N_19206);
nor U19400 (N_19400,N_19210,N_19311);
xor U19401 (N_19401,N_19285,N_19270);
or U19402 (N_19402,N_19342,N_19235);
and U19403 (N_19403,N_19207,N_19295);
xnor U19404 (N_19404,N_19301,N_19259);
nor U19405 (N_19405,N_19217,N_19332);
nor U19406 (N_19406,N_19297,N_19317);
or U19407 (N_19407,N_19347,N_19336);
and U19408 (N_19408,N_19209,N_19266);
or U19409 (N_19409,N_19296,N_19279);
nor U19410 (N_19410,N_19293,N_19324);
or U19411 (N_19411,N_19267,N_19254);
and U19412 (N_19412,N_19337,N_19304);
nand U19413 (N_19413,N_19340,N_19327);
nand U19414 (N_19414,N_19335,N_19305);
and U19415 (N_19415,N_19299,N_19352);
xor U19416 (N_19416,N_19257,N_19200);
and U19417 (N_19417,N_19224,N_19318);
xnor U19418 (N_19418,N_19250,N_19316);
xnor U19419 (N_19419,N_19303,N_19349);
and U19420 (N_19420,N_19225,N_19271);
nor U19421 (N_19421,N_19322,N_19291);
nor U19422 (N_19422,N_19253,N_19230);
nor U19423 (N_19423,N_19256,N_19345);
and U19424 (N_19424,N_19233,N_19236);
and U19425 (N_19425,N_19243,N_19353);
nand U19426 (N_19426,N_19351,N_19205);
nand U19427 (N_19427,N_19273,N_19325);
and U19428 (N_19428,N_19288,N_19294);
nor U19429 (N_19429,N_19326,N_19280);
or U19430 (N_19430,N_19228,N_19292);
nor U19431 (N_19431,N_19242,N_19274);
nand U19432 (N_19432,N_19258,N_19343);
or U19433 (N_19433,N_19237,N_19344);
and U19434 (N_19434,N_19244,N_19264);
nor U19435 (N_19435,N_19211,N_19331);
xor U19436 (N_19436,N_19251,N_19338);
or U19437 (N_19437,N_19277,N_19246);
nand U19438 (N_19438,N_19290,N_19241);
nor U19439 (N_19439,N_19348,N_19212);
nor U19440 (N_19440,N_19240,N_19233);
or U19441 (N_19441,N_19358,N_19343);
and U19442 (N_19442,N_19201,N_19214);
xnor U19443 (N_19443,N_19213,N_19273);
or U19444 (N_19444,N_19293,N_19345);
and U19445 (N_19445,N_19277,N_19323);
nor U19446 (N_19446,N_19351,N_19294);
xor U19447 (N_19447,N_19299,N_19272);
nand U19448 (N_19448,N_19316,N_19215);
nand U19449 (N_19449,N_19289,N_19336);
and U19450 (N_19450,N_19241,N_19222);
and U19451 (N_19451,N_19273,N_19245);
and U19452 (N_19452,N_19275,N_19210);
nand U19453 (N_19453,N_19355,N_19281);
nand U19454 (N_19454,N_19275,N_19218);
nor U19455 (N_19455,N_19304,N_19207);
nand U19456 (N_19456,N_19292,N_19282);
nor U19457 (N_19457,N_19214,N_19262);
nor U19458 (N_19458,N_19343,N_19283);
and U19459 (N_19459,N_19256,N_19263);
or U19460 (N_19460,N_19329,N_19248);
and U19461 (N_19461,N_19279,N_19349);
xor U19462 (N_19462,N_19325,N_19203);
nand U19463 (N_19463,N_19261,N_19264);
nand U19464 (N_19464,N_19291,N_19317);
nand U19465 (N_19465,N_19207,N_19205);
and U19466 (N_19466,N_19249,N_19211);
nand U19467 (N_19467,N_19253,N_19236);
and U19468 (N_19468,N_19272,N_19354);
xnor U19469 (N_19469,N_19200,N_19218);
and U19470 (N_19470,N_19216,N_19338);
or U19471 (N_19471,N_19272,N_19294);
nor U19472 (N_19472,N_19208,N_19269);
nor U19473 (N_19473,N_19263,N_19220);
and U19474 (N_19474,N_19329,N_19231);
xnor U19475 (N_19475,N_19262,N_19264);
and U19476 (N_19476,N_19329,N_19345);
xnor U19477 (N_19477,N_19276,N_19264);
nand U19478 (N_19478,N_19346,N_19332);
and U19479 (N_19479,N_19247,N_19297);
or U19480 (N_19480,N_19215,N_19267);
and U19481 (N_19481,N_19306,N_19223);
nand U19482 (N_19482,N_19207,N_19291);
nand U19483 (N_19483,N_19268,N_19359);
and U19484 (N_19484,N_19249,N_19291);
nor U19485 (N_19485,N_19325,N_19222);
or U19486 (N_19486,N_19248,N_19337);
nand U19487 (N_19487,N_19237,N_19246);
and U19488 (N_19488,N_19358,N_19248);
nand U19489 (N_19489,N_19291,N_19340);
and U19490 (N_19490,N_19342,N_19297);
xnor U19491 (N_19491,N_19244,N_19226);
xnor U19492 (N_19492,N_19283,N_19270);
and U19493 (N_19493,N_19348,N_19262);
and U19494 (N_19494,N_19355,N_19306);
nand U19495 (N_19495,N_19344,N_19316);
and U19496 (N_19496,N_19250,N_19202);
and U19497 (N_19497,N_19290,N_19266);
xor U19498 (N_19498,N_19279,N_19343);
xnor U19499 (N_19499,N_19211,N_19250);
nor U19500 (N_19500,N_19290,N_19339);
or U19501 (N_19501,N_19221,N_19333);
nor U19502 (N_19502,N_19302,N_19289);
nor U19503 (N_19503,N_19224,N_19226);
nand U19504 (N_19504,N_19313,N_19204);
xor U19505 (N_19505,N_19275,N_19274);
and U19506 (N_19506,N_19235,N_19270);
and U19507 (N_19507,N_19354,N_19334);
xor U19508 (N_19508,N_19259,N_19203);
and U19509 (N_19509,N_19306,N_19333);
or U19510 (N_19510,N_19345,N_19274);
nand U19511 (N_19511,N_19226,N_19274);
xor U19512 (N_19512,N_19293,N_19348);
and U19513 (N_19513,N_19312,N_19317);
nand U19514 (N_19514,N_19293,N_19252);
nor U19515 (N_19515,N_19312,N_19300);
nand U19516 (N_19516,N_19269,N_19346);
and U19517 (N_19517,N_19284,N_19228);
xor U19518 (N_19518,N_19317,N_19214);
or U19519 (N_19519,N_19318,N_19304);
nor U19520 (N_19520,N_19457,N_19448);
or U19521 (N_19521,N_19445,N_19390);
nor U19522 (N_19522,N_19504,N_19456);
and U19523 (N_19523,N_19389,N_19486);
and U19524 (N_19524,N_19382,N_19380);
xor U19525 (N_19525,N_19452,N_19377);
or U19526 (N_19526,N_19519,N_19498);
nand U19527 (N_19527,N_19410,N_19502);
xnor U19528 (N_19528,N_19371,N_19416);
xor U19529 (N_19529,N_19372,N_19487);
xnor U19530 (N_19530,N_19387,N_19460);
nor U19531 (N_19531,N_19506,N_19399);
xnor U19532 (N_19532,N_19476,N_19364);
nand U19533 (N_19533,N_19493,N_19459);
xor U19534 (N_19534,N_19438,N_19407);
and U19535 (N_19535,N_19474,N_19484);
nand U19536 (N_19536,N_19458,N_19505);
and U19537 (N_19537,N_19411,N_19497);
or U19538 (N_19538,N_19501,N_19369);
nand U19539 (N_19539,N_19385,N_19499);
or U19540 (N_19540,N_19464,N_19404);
xor U19541 (N_19541,N_19494,N_19455);
nor U19542 (N_19542,N_19397,N_19509);
or U19543 (N_19543,N_19405,N_19413);
nand U19544 (N_19544,N_19518,N_19403);
xnor U19545 (N_19545,N_19480,N_19489);
xnor U19546 (N_19546,N_19415,N_19362);
nand U19547 (N_19547,N_19418,N_19450);
or U19548 (N_19548,N_19421,N_19447);
or U19549 (N_19549,N_19409,N_19378);
or U19550 (N_19550,N_19386,N_19492);
or U19551 (N_19551,N_19495,N_19483);
nand U19552 (N_19552,N_19436,N_19488);
and U19553 (N_19553,N_19425,N_19402);
and U19554 (N_19554,N_19444,N_19395);
or U19555 (N_19555,N_19414,N_19469);
nor U19556 (N_19556,N_19500,N_19510);
or U19557 (N_19557,N_19420,N_19485);
xnor U19558 (N_19558,N_19412,N_19496);
and U19559 (N_19559,N_19441,N_19431);
or U19560 (N_19560,N_19381,N_19401);
xnor U19561 (N_19561,N_19453,N_19426);
xor U19562 (N_19562,N_19408,N_19422);
nor U19563 (N_19563,N_19406,N_19514);
xor U19564 (N_19564,N_19437,N_19516);
xnor U19565 (N_19565,N_19461,N_19424);
xnor U19566 (N_19566,N_19434,N_19491);
nor U19567 (N_19567,N_19393,N_19490);
nor U19568 (N_19568,N_19507,N_19417);
nor U19569 (N_19569,N_19374,N_19433);
nor U19570 (N_19570,N_19472,N_19440);
xnor U19571 (N_19571,N_19370,N_19508);
nor U19572 (N_19572,N_19512,N_19379);
or U19573 (N_19573,N_19400,N_19468);
nand U19574 (N_19574,N_19376,N_19511);
nor U19575 (N_19575,N_19449,N_19481);
and U19576 (N_19576,N_19398,N_19503);
nor U19577 (N_19577,N_19428,N_19432);
xnor U19578 (N_19578,N_19454,N_19363);
xor U19579 (N_19579,N_19423,N_19479);
nand U19580 (N_19580,N_19471,N_19443);
and U19581 (N_19581,N_19478,N_19366);
xor U19582 (N_19582,N_19465,N_19427);
or U19583 (N_19583,N_19517,N_19361);
xnor U19584 (N_19584,N_19419,N_19373);
nor U19585 (N_19585,N_19467,N_19482);
or U19586 (N_19586,N_19475,N_19384);
nand U19587 (N_19587,N_19466,N_19375);
nor U19588 (N_19588,N_19513,N_19394);
nand U19589 (N_19589,N_19388,N_19360);
xnor U19590 (N_19590,N_19462,N_19430);
or U19591 (N_19591,N_19392,N_19477);
xor U19592 (N_19592,N_19365,N_19473);
or U19593 (N_19593,N_19391,N_19451);
nand U19594 (N_19594,N_19368,N_19463);
and U19595 (N_19595,N_19435,N_19439);
xnor U19596 (N_19596,N_19429,N_19470);
and U19597 (N_19597,N_19383,N_19396);
nor U19598 (N_19598,N_19515,N_19446);
nand U19599 (N_19599,N_19367,N_19442);
nor U19600 (N_19600,N_19376,N_19507);
or U19601 (N_19601,N_19427,N_19462);
or U19602 (N_19602,N_19501,N_19493);
nand U19603 (N_19603,N_19466,N_19518);
nand U19604 (N_19604,N_19515,N_19396);
xor U19605 (N_19605,N_19445,N_19483);
xnor U19606 (N_19606,N_19502,N_19433);
xnor U19607 (N_19607,N_19518,N_19437);
and U19608 (N_19608,N_19456,N_19442);
or U19609 (N_19609,N_19428,N_19409);
and U19610 (N_19610,N_19491,N_19462);
and U19611 (N_19611,N_19503,N_19455);
or U19612 (N_19612,N_19375,N_19409);
xnor U19613 (N_19613,N_19496,N_19386);
and U19614 (N_19614,N_19435,N_19447);
and U19615 (N_19615,N_19504,N_19430);
nand U19616 (N_19616,N_19444,N_19500);
or U19617 (N_19617,N_19399,N_19393);
and U19618 (N_19618,N_19498,N_19480);
nor U19619 (N_19619,N_19463,N_19492);
or U19620 (N_19620,N_19487,N_19461);
nor U19621 (N_19621,N_19381,N_19479);
nand U19622 (N_19622,N_19381,N_19412);
nand U19623 (N_19623,N_19382,N_19436);
and U19624 (N_19624,N_19489,N_19488);
nand U19625 (N_19625,N_19387,N_19471);
xnor U19626 (N_19626,N_19462,N_19484);
nor U19627 (N_19627,N_19461,N_19501);
nor U19628 (N_19628,N_19498,N_19417);
or U19629 (N_19629,N_19462,N_19382);
or U19630 (N_19630,N_19391,N_19470);
nor U19631 (N_19631,N_19370,N_19423);
and U19632 (N_19632,N_19478,N_19425);
nand U19633 (N_19633,N_19492,N_19363);
xnor U19634 (N_19634,N_19407,N_19429);
nand U19635 (N_19635,N_19514,N_19360);
or U19636 (N_19636,N_19504,N_19508);
xor U19637 (N_19637,N_19390,N_19470);
and U19638 (N_19638,N_19512,N_19389);
and U19639 (N_19639,N_19479,N_19474);
nor U19640 (N_19640,N_19510,N_19367);
or U19641 (N_19641,N_19411,N_19508);
and U19642 (N_19642,N_19499,N_19390);
and U19643 (N_19643,N_19418,N_19499);
xnor U19644 (N_19644,N_19474,N_19378);
or U19645 (N_19645,N_19420,N_19363);
or U19646 (N_19646,N_19463,N_19421);
nor U19647 (N_19647,N_19398,N_19498);
nor U19648 (N_19648,N_19507,N_19496);
nor U19649 (N_19649,N_19484,N_19446);
xnor U19650 (N_19650,N_19463,N_19436);
nor U19651 (N_19651,N_19467,N_19460);
or U19652 (N_19652,N_19404,N_19484);
or U19653 (N_19653,N_19361,N_19393);
and U19654 (N_19654,N_19437,N_19493);
nor U19655 (N_19655,N_19506,N_19472);
nor U19656 (N_19656,N_19456,N_19507);
nor U19657 (N_19657,N_19436,N_19448);
nor U19658 (N_19658,N_19509,N_19444);
xor U19659 (N_19659,N_19375,N_19496);
and U19660 (N_19660,N_19420,N_19488);
and U19661 (N_19661,N_19415,N_19444);
nand U19662 (N_19662,N_19484,N_19453);
nor U19663 (N_19663,N_19476,N_19367);
nand U19664 (N_19664,N_19384,N_19400);
and U19665 (N_19665,N_19361,N_19478);
xnor U19666 (N_19666,N_19414,N_19407);
nand U19667 (N_19667,N_19491,N_19476);
nor U19668 (N_19668,N_19448,N_19400);
nor U19669 (N_19669,N_19386,N_19425);
or U19670 (N_19670,N_19423,N_19407);
and U19671 (N_19671,N_19462,N_19452);
nand U19672 (N_19672,N_19515,N_19447);
nor U19673 (N_19673,N_19386,N_19472);
or U19674 (N_19674,N_19415,N_19416);
nor U19675 (N_19675,N_19518,N_19486);
nor U19676 (N_19676,N_19426,N_19512);
nor U19677 (N_19677,N_19376,N_19479);
xor U19678 (N_19678,N_19419,N_19475);
xnor U19679 (N_19679,N_19429,N_19519);
xnor U19680 (N_19680,N_19679,N_19606);
nand U19681 (N_19681,N_19632,N_19570);
nor U19682 (N_19682,N_19543,N_19669);
nor U19683 (N_19683,N_19622,N_19620);
and U19684 (N_19684,N_19646,N_19554);
nand U19685 (N_19685,N_19642,N_19582);
nand U19686 (N_19686,N_19578,N_19562);
xnor U19687 (N_19687,N_19590,N_19566);
and U19688 (N_19688,N_19636,N_19548);
nor U19689 (N_19689,N_19652,N_19569);
xnor U19690 (N_19690,N_19631,N_19637);
and U19691 (N_19691,N_19580,N_19648);
nand U19692 (N_19692,N_19593,N_19536);
xnor U19693 (N_19693,N_19533,N_19545);
xor U19694 (N_19694,N_19635,N_19623);
nor U19695 (N_19695,N_19535,N_19673);
or U19696 (N_19696,N_19576,N_19586);
nand U19697 (N_19697,N_19564,N_19575);
nand U19698 (N_19698,N_19573,N_19602);
nor U19699 (N_19699,N_19527,N_19655);
xnor U19700 (N_19700,N_19556,N_19539);
or U19701 (N_19701,N_19532,N_19670);
nor U19702 (N_19702,N_19625,N_19672);
nand U19703 (N_19703,N_19592,N_19547);
and U19704 (N_19704,N_19537,N_19540);
or U19705 (N_19705,N_19561,N_19563);
nand U19706 (N_19706,N_19671,N_19613);
xnor U19707 (N_19707,N_19608,N_19555);
xnor U19708 (N_19708,N_19601,N_19565);
and U19709 (N_19709,N_19571,N_19552);
nand U19710 (N_19710,N_19616,N_19583);
or U19711 (N_19711,N_19657,N_19597);
and U19712 (N_19712,N_19656,N_19675);
xnor U19713 (N_19713,N_19612,N_19574);
nand U19714 (N_19714,N_19660,N_19595);
or U19715 (N_19715,N_19530,N_19629);
or U19716 (N_19716,N_19619,N_19523);
and U19717 (N_19717,N_19529,N_19607);
nor U19718 (N_19718,N_19542,N_19643);
nand U19719 (N_19719,N_19638,N_19615);
and U19720 (N_19720,N_19653,N_19634);
or U19721 (N_19721,N_19665,N_19579);
or U19722 (N_19722,N_19538,N_19526);
xnor U19723 (N_19723,N_19645,N_19605);
xor U19724 (N_19724,N_19559,N_19621);
xor U19725 (N_19725,N_19603,N_19676);
xor U19726 (N_19726,N_19525,N_19534);
nor U19727 (N_19727,N_19528,N_19585);
or U19728 (N_19728,N_19522,N_19568);
or U19729 (N_19729,N_19549,N_19666);
xnor U19730 (N_19730,N_19520,N_19663);
nor U19731 (N_19731,N_19541,N_19584);
nand U19732 (N_19732,N_19618,N_19544);
xor U19733 (N_19733,N_19674,N_19598);
and U19734 (N_19734,N_19667,N_19604);
and U19735 (N_19735,N_19557,N_19600);
or U19736 (N_19736,N_19558,N_19531);
xnor U19737 (N_19737,N_19551,N_19659);
xor U19738 (N_19738,N_19611,N_19641);
and U19739 (N_19739,N_19572,N_19644);
nor U19740 (N_19740,N_19633,N_19591);
or U19741 (N_19741,N_19649,N_19668);
and U19742 (N_19742,N_19609,N_19550);
or U19743 (N_19743,N_19521,N_19588);
nor U19744 (N_19744,N_19627,N_19560);
xnor U19745 (N_19745,N_19664,N_19647);
xor U19746 (N_19746,N_19587,N_19594);
nand U19747 (N_19747,N_19651,N_19614);
and U19748 (N_19748,N_19661,N_19626);
xor U19749 (N_19749,N_19662,N_19524);
and U19750 (N_19750,N_19677,N_19678);
and U19751 (N_19751,N_19577,N_19658);
and U19752 (N_19752,N_19639,N_19617);
and U19753 (N_19753,N_19567,N_19640);
xor U19754 (N_19754,N_19553,N_19654);
and U19755 (N_19755,N_19581,N_19599);
xnor U19756 (N_19756,N_19624,N_19596);
xor U19757 (N_19757,N_19630,N_19610);
and U19758 (N_19758,N_19546,N_19650);
and U19759 (N_19759,N_19589,N_19628);
xor U19760 (N_19760,N_19622,N_19674);
and U19761 (N_19761,N_19635,N_19624);
nor U19762 (N_19762,N_19584,N_19624);
xnor U19763 (N_19763,N_19673,N_19566);
nand U19764 (N_19764,N_19574,N_19668);
nand U19765 (N_19765,N_19627,N_19608);
xor U19766 (N_19766,N_19673,N_19546);
nand U19767 (N_19767,N_19522,N_19625);
and U19768 (N_19768,N_19635,N_19646);
and U19769 (N_19769,N_19622,N_19540);
xor U19770 (N_19770,N_19664,N_19581);
nor U19771 (N_19771,N_19590,N_19612);
or U19772 (N_19772,N_19649,N_19559);
and U19773 (N_19773,N_19559,N_19666);
xor U19774 (N_19774,N_19523,N_19642);
nor U19775 (N_19775,N_19522,N_19641);
xnor U19776 (N_19776,N_19582,N_19551);
xor U19777 (N_19777,N_19677,N_19556);
nor U19778 (N_19778,N_19632,N_19587);
or U19779 (N_19779,N_19625,N_19635);
nor U19780 (N_19780,N_19601,N_19563);
nand U19781 (N_19781,N_19603,N_19630);
and U19782 (N_19782,N_19613,N_19665);
nand U19783 (N_19783,N_19581,N_19662);
nand U19784 (N_19784,N_19626,N_19658);
and U19785 (N_19785,N_19620,N_19578);
or U19786 (N_19786,N_19659,N_19657);
nand U19787 (N_19787,N_19581,N_19576);
or U19788 (N_19788,N_19605,N_19625);
or U19789 (N_19789,N_19678,N_19588);
or U19790 (N_19790,N_19576,N_19667);
nand U19791 (N_19791,N_19591,N_19578);
and U19792 (N_19792,N_19594,N_19602);
or U19793 (N_19793,N_19624,N_19588);
nand U19794 (N_19794,N_19658,N_19523);
or U19795 (N_19795,N_19655,N_19599);
or U19796 (N_19796,N_19541,N_19631);
xnor U19797 (N_19797,N_19643,N_19658);
nor U19798 (N_19798,N_19569,N_19549);
nor U19799 (N_19799,N_19598,N_19636);
xnor U19800 (N_19800,N_19609,N_19613);
nand U19801 (N_19801,N_19539,N_19534);
xor U19802 (N_19802,N_19624,N_19587);
nor U19803 (N_19803,N_19612,N_19576);
or U19804 (N_19804,N_19534,N_19581);
nand U19805 (N_19805,N_19666,N_19597);
nand U19806 (N_19806,N_19671,N_19609);
nand U19807 (N_19807,N_19526,N_19626);
nor U19808 (N_19808,N_19635,N_19664);
or U19809 (N_19809,N_19524,N_19581);
or U19810 (N_19810,N_19646,N_19634);
and U19811 (N_19811,N_19605,N_19556);
or U19812 (N_19812,N_19646,N_19537);
nor U19813 (N_19813,N_19615,N_19596);
or U19814 (N_19814,N_19602,N_19547);
xnor U19815 (N_19815,N_19626,N_19568);
or U19816 (N_19816,N_19595,N_19613);
and U19817 (N_19817,N_19637,N_19528);
or U19818 (N_19818,N_19534,N_19612);
nor U19819 (N_19819,N_19593,N_19546);
or U19820 (N_19820,N_19637,N_19561);
or U19821 (N_19821,N_19552,N_19650);
nor U19822 (N_19822,N_19522,N_19612);
nor U19823 (N_19823,N_19534,N_19662);
nand U19824 (N_19824,N_19596,N_19656);
or U19825 (N_19825,N_19520,N_19550);
nor U19826 (N_19826,N_19620,N_19564);
and U19827 (N_19827,N_19590,N_19653);
and U19828 (N_19828,N_19607,N_19592);
or U19829 (N_19829,N_19645,N_19531);
and U19830 (N_19830,N_19598,N_19630);
and U19831 (N_19831,N_19663,N_19644);
xor U19832 (N_19832,N_19591,N_19537);
nor U19833 (N_19833,N_19548,N_19663);
and U19834 (N_19834,N_19620,N_19558);
nand U19835 (N_19835,N_19644,N_19648);
xor U19836 (N_19836,N_19548,N_19554);
xnor U19837 (N_19837,N_19612,N_19609);
nand U19838 (N_19838,N_19570,N_19521);
nand U19839 (N_19839,N_19634,N_19667);
nor U19840 (N_19840,N_19757,N_19777);
or U19841 (N_19841,N_19684,N_19764);
or U19842 (N_19842,N_19748,N_19790);
or U19843 (N_19843,N_19767,N_19707);
and U19844 (N_19844,N_19789,N_19687);
nor U19845 (N_19845,N_19696,N_19690);
xor U19846 (N_19846,N_19727,N_19766);
or U19847 (N_19847,N_19752,N_19786);
nand U19848 (N_19848,N_19806,N_19762);
xnor U19849 (N_19849,N_19769,N_19787);
nand U19850 (N_19850,N_19710,N_19801);
nor U19851 (N_19851,N_19768,N_19740);
xnor U19852 (N_19852,N_19798,N_19830);
or U19853 (N_19853,N_19681,N_19820);
nand U19854 (N_19854,N_19708,N_19719);
and U19855 (N_19855,N_19728,N_19738);
nand U19856 (N_19856,N_19746,N_19754);
nand U19857 (N_19857,N_19826,N_19717);
nand U19858 (N_19858,N_19691,N_19739);
nor U19859 (N_19859,N_19760,N_19701);
and U19860 (N_19860,N_19814,N_19791);
and U19861 (N_19861,N_19810,N_19699);
or U19862 (N_19862,N_19750,N_19809);
and U19863 (N_19863,N_19712,N_19744);
xnor U19864 (N_19864,N_19730,N_19765);
xor U19865 (N_19865,N_19695,N_19822);
and U19866 (N_19866,N_19736,N_19733);
or U19867 (N_19867,N_19698,N_19702);
nand U19868 (N_19868,N_19759,N_19774);
or U19869 (N_19869,N_19795,N_19705);
xor U19870 (N_19870,N_19817,N_19823);
and U19871 (N_19871,N_19782,N_19689);
nand U19872 (N_19872,N_19753,N_19819);
or U19873 (N_19873,N_19731,N_19737);
nand U19874 (N_19874,N_19709,N_19703);
or U19875 (N_19875,N_19778,N_19706);
xnor U19876 (N_19876,N_19793,N_19811);
xnor U19877 (N_19877,N_19805,N_19725);
nor U19878 (N_19878,N_19682,N_19781);
nand U19879 (N_19879,N_19694,N_19756);
xor U19880 (N_19880,N_19761,N_19772);
and U19881 (N_19881,N_19838,N_19680);
and U19882 (N_19882,N_19718,N_19807);
xor U19883 (N_19883,N_19692,N_19815);
nor U19884 (N_19884,N_19683,N_19723);
or U19885 (N_19885,N_19779,N_19800);
and U19886 (N_19886,N_19755,N_19788);
nand U19887 (N_19887,N_19726,N_19808);
and U19888 (N_19888,N_19775,N_19776);
and U19889 (N_19889,N_19735,N_19688);
and U19890 (N_19890,N_19821,N_19796);
and U19891 (N_19891,N_19839,N_19785);
and U19892 (N_19892,N_19713,N_19802);
xor U19893 (N_19893,N_19721,N_19720);
xor U19894 (N_19894,N_19797,N_19751);
nand U19895 (N_19895,N_19784,N_19742);
or U19896 (N_19896,N_19700,N_19715);
and U19897 (N_19897,N_19816,N_19741);
nor U19898 (N_19898,N_19745,N_19771);
or U19899 (N_19899,N_19734,N_19732);
or U19900 (N_19900,N_19812,N_19835);
xnor U19901 (N_19901,N_19828,N_19716);
and U19902 (N_19902,N_19827,N_19722);
nand U19903 (N_19903,N_19832,N_19773);
and U19904 (N_19904,N_19833,N_19749);
and U19905 (N_19905,N_19685,N_19831);
xor U19906 (N_19906,N_19834,N_19704);
nand U19907 (N_19907,N_19829,N_19804);
nand U19908 (N_19908,N_19799,N_19693);
or U19909 (N_19909,N_19824,N_19758);
or U19910 (N_19910,N_19697,N_19825);
nand U19911 (N_19911,N_19836,N_19747);
xnor U19912 (N_19912,N_19714,N_19763);
or U19913 (N_19913,N_19813,N_19818);
or U19914 (N_19914,N_19783,N_19729);
nor U19915 (N_19915,N_19837,N_19686);
nand U19916 (N_19916,N_19711,N_19770);
nor U19917 (N_19917,N_19792,N_19803);
nor U19918 (N_19918,N_19780,N_19794);
nor U19919 (N_19919,N_19743,N_19724);
nand U19920 (N_19920,N_19699,N_19680);
xor U19921 (N_19921,N_19769,N_19728);
xor U19922 (N_19922,N_19815,N_19768);
or U19923 (N_19923,N_19829,N_19699);
xor U19924 (N_19924,N_19735,N_19782);
and U19925 (N_19925,N_19819,N_19836);
xnor U19926 (N_19926,N_19706,N_19715);
and U19927 (N_19927,N_19729,N_19771);
nand U19928 (N_19928,N_19808,N_19817);
or U19929 (N_19929,N_19705,N_19808);
nand U19930 (N_19930,N_19836,N_19796);
nand U19931 (N_19931,N_19803,N_19783);
and U19932 (N_19932,N_19785,N_19781);
nand U19933 (N_19933,N_19824,N_19763);
xor U19934 (N_19934,N_19804,N_19837);
and U19935 (N_19935,N_19711,N_19707);
or U19936 (N_19936,N_19833,N_19730);
nor U19937 (N_19937,N_19761,N_19766);
nor U19938 (N_19938,N_19681,N_19762);
nor U19939 (N_19939,N_19680,N_19711);
and U19940 (N_19940,N_19771,N_19780);
and U19941 (N_19941,N_19775,N_19707);
and U19942 (N_19942,N_19691,N_19703);
nand U19943 (N_19943,N_19713,N_19696);
nand U19944 (N_19944,N_19792,N_19736);
and U19945 (N_19945,N_19765,N_19737);
xor U19946 (N_19946,N_19810,N_19755);
xor U19947 (N_19947,N_19790,N_19814);
and U19948 (N_19948,N_19761,N_19812);
nor U19949 (N_19949,N_19795,N_19738);
nand U19950 (N_19950,N_19797,N_19702);
nand U19951 (N_19951,N_19782,N_19828);
xnor U19952 (N_19952,N_19696,N_19738);
or U19953 (N_19953,N_19776,N_19795);
or U19954 (N_19954,N_19763,N_19745);
nor U19955 (N_19955,N_19791,N_19695);
nor U19956 (N_19956,N_19708,N_19827);
or U19957 (N_19957,N_19728,N_19794);
xor U19958 (N_19958,N_19828,N_19704);
nand U19959 (N_19959,N_19715,N_19825);
and U19960 (N_19960,N_19778,N_19825);
nor U19961 (N_19961,N_19794,N_19756);
and U19962 (N_19962,N_19785,N_19838);
and U19963 (N_19963,N_19684,N_19786);
and U19964 (N_19964,N_19745,N_19708);
and U19965 (N_19965,N_19806,N_19724);
nand U19966 (N_19966,N_19759,N_19787);
xor U19967 (N_19967,N_19762,N_19820);
nand U19968 (N_19968,N_19748,N_19800);
xor U19969 (N_19969,N_19818,N_19732);
nor U19970 (N_19970,N_19750,N_19807);
and U19971 (N_19971,N_19792,N_19771);
nand U19972 (N_19972,N_19761,N_19749);
and U19973 (N_19973,N_19762,N_19807);
or U19974 (N_19974,N_19804,N_19710);
and U19975 (N_19975,N_19757,N_19721);
nor U19976 (N_19976,N_19748,N_19771);
nor U19977 (N_19977,N_19784,N_19785);
nor U19978 (N_19978,N_19769,N_19689);
and U19979 (N_19979,N_19791,N_19718);
nor U19980 (N_19980,N_19736,N_19707);
xnor U19981 (N_19981,N_19775,N_19729);
nor U19982 (N_19982,N_19717,N_19807);
nor U19983 (N_19983,N_19759,N_19813);
xor U19984 (N_19984,N_19711,N_19740);
nor U19985 (N_19985,N_19746,N_19684);
nand U19986 (N_19986,N_19714,N_19800);
and U19987 (N_19987,N_19800,N_19791);
or U19988 (N_19988,N_19737,N_19781);
nand U19989 (N_19989,N_19834,N_19753);
nand U19990 (N_19990,N_19722,N_19730);
nor U19991 (N_19991,N_19727,N_19713);
nand U19992 (N_19992,N_19773,N_19784);
nand U19993 (N_19993,N_19736,N_19751);
nand U19994 (N_19994,N_19726,N_19742);
or U19995 (N_19995,N_19764,N_19696);
or U19996 (N_19996,N_19801,N_19812);
xnor U19997 (N_19997,N_19703,N_19837);
nor U19998 (N_19998,N_19794,N_19696);
nand U19999 (N_19999,N_19713,N_19687);
xnor UO_0 (O_0,N_19896,N_19858);
or UO_1 (O_1,N_19870,N_19970);
and UO_2 (O_2,N_19921,N_19875);
nand UO_3 (O_3,N_19999,N_19846);
nor UO_4 (O_4,N_19990,N_19973);
nand UO_5 (O_5,N_19879,N_19862);
xnor UO_6 (O_6,N_19865,N_19908);
nand UO_7 (O_7,N_19893,N_19906);
and UO_8 (O_8,N_19867,N_19905);
nor UO_9 (O_9,N_19844,N_19956);
nand UO_10 (O_10,N_19866,N_19864);
and UO_11 (O_11,N_19929,N_19994);
nor UO_12 (O_12,N_19887,N_19901);
nor UO_13 (O_13,N_19903,N_19947);
xor UO_14 (O_14,N_19853,N_19876);
nor UO_15 (O_15,N_19873,N_19860);
nor UO_16 (O_16,N_19920,N_19911);
nand UO_17 (O_17,N_19933,N_19945);
xnor UO_18 (O_18,N_19847,N_19910);
and UO_19 (O_19,N_19951,N_19918);
and UO_20 (O_20,N_19952,N_19874);
and UO_21 (O_21,N_19872,N_19976);
xnor UO_22 (O_22,N_19968,N_19966);
or UO_23 (O_23,N_19924,N_19878);
and UO_24 (O_24,N_19871,N_19856);
or UO_25 (O_25,N_19961,N_19986);
and UO_26 (O_26,N_19937,N_19988);
nand UO_27 (O_27,N_19900,N_19941);
nand UO_28 (O_28,N_19996,N_19964);
or UO_29 (O_29,N_19979,N_19949);
nand UO_30 (O_30,N_19985,N_19975);
nor UO_31 (O_31,N_19957,N_19917);
or UO_32 (O_32,N_19895,N_19890);
and UO_33 (O_33,N_19977,N_19842);
xnor UO_34 (O_34,N_19938,N_19935);
or UO_35 (O_35,N_19885,N_19869);
nor UO_36 (O_36,N_19950,N_19904);
nand UO_37 (O_37,N_19926,N_19868);
nor UO_38 (O_38,N_19997,N_19927);
nor UO_39 (O_39,N_19897,N_19944);
nand UO_40 (O_40,N_19932,N_19978);
xor UO_41 (O_41,N_19991,N_19922);
or UO_42 (O_42,N_19959,N_19962);
or UO_43 (O_43,N_19851,N_19981);
or UO_44 (O_44,N_19849,N_19955);
and UO_45 (O_45,N_19850,N_19919);
nand UO_46 (O_46,N_19940,N_19845);
and UO_47 (O_47,N_19913,N_19914);
and UO_48 (O_48,N_19841,N_19861);
and UO_49 (O_49,N_19843,N_19972);
nand UO_50 (O_50,N_19995,N_19953);
nand UO_51 (O_51,N_19884,N_19930);
xor UO_52 (O_52,N_19923,N_19928);
and UO_53 (O_53,N_19971,N_19925);
nand UO_54 (O_54,N_19946,N_19931);
and UO_55 (O_55,N_19880,N_19894);
or UO_56 (O_56,N_19852,N_19983);
nand UO_57 (O_57,N_19943,N_19939);
and UO_58 (O_58,N_19980,N_19912);
or UO_59 (O_59,N_19855,N_19892);
nand UO_60 (O_60,N_19909,N_19859);
and UO_61 (O_61,N_19958,N_19987);
xor UO_62 (O_62,N_19982,N_19916);
and UO_63 (O_63,N_19888,N_19907);
nand UO_64 (O_64,N_19881,N_19967);
nand UO_65 (O_65,N_19863,N_19998);
and UO_66 (O_66,N_19848,N_19942);
nand UO_67 (O_67,N_19854,N_19965);
or UO_68 (O_68,N_19877,N_19902);
and UO_69 (O_69,N_19936,N_19840);
nor UO_70 (O_70,N_19857,N_19948);
or UO_71 (O_71,N_19898,N_19934);
xnor UO_72 (O_72,N_19899,N_19969);
or UO_73 (O_73,N_19889,N_19915);
or UO_74 (O_74,N_19886,N_19883);
nand UO_75 (O_75,N_19954,N_19992);
and UO_76 (O_76,N_19984,N_19974);
or UO_77 (O_77,N_19960,N_19891);
and UO_78 (O_78,N_19993,N_19963);
nor UO_79 (O_79,N_19989,N_19882);
nand UO_80 (O_80,N_19859,N_19864);
nand UO_81 (O_81,N_19874,N_19891);
xor UO_82 (O_82,N_19855,N_19926);
nor UO_83 (O_83,N_19974,N_19855);
or UO_84 (O_84,N_19841,N_19941);
and UO_85 (O_85,N_19896,N_19859);
nand UO_86 (O_86,N_19872,N_19971);
or UO_87 (O_87,N_19990,N_19904);
nand UO_88 (O_88,N_19935,N_19911);
nand UO_89 (O_89,N_19962,N_19898);
xnor UO_90 (O_90,N_19892,N_19925);
and UO_91 (O_91,N_19914,N_19841);
or UO_92 (O_92,N_19955,N_19861);
and UO_93 (O_93,N_19890,N_19868);
nand UO_94 (O_94,N_19938,N_19971);
and UO_95 (O_95,N_19973,N_19999);
nor UO_96 (O_96,N_19914,N_19861);
nand UO_97 (O_97,N_19903,N_19884);
or UO_98 (O_98,N_19886,N_19863);
nand UO_99 (O_99,N_19911,N_19969);
and UO_100 (O_100,N_19961,N_19966);
xnor UO_101 (O_101,N_19966,N_19844);
nor UO_102 (O_102,N_19989,N_19877);
nand UO_103 (O_103,N_19849,N_19934);
and UO_104 (O_104,N_19922,N_19930);
nor UO_105 (O_105,N_19901,N_19921);
nand UO_106 (O_106,N_19956,N_19927);
nor UO_107 (O_107,N_19864,N_19940);
and UO_108 (O_108,N_19929,N_19904);
or UO_109 (O_109,N_19890,N_19881);
nand UO_110 (O_110,N_19851,N_19928);
and UO_111 (O_111,N_19869,N_19968);
or UO_112 (O_112,N_19899,N_19880);
nor UO_113 (O_113,N_19875,N_19930);
nor UO_114 (O_114,N_19969,N_19895);
or UO_115 (O_115,N_19876,N_19955);
and UO_116 (O_116,N_19980,N_19926);
nand UO_117 (O_117,N_19961,N_19913);
xnor UO_118 (O_118,N_19840,N_19987);
nor UO_119 (O_119,N_19841,N_19948);
or UO_120 (O_120,N_19885,N_19937);
nor UO_121 (O_121,N_19976,N_19886);
xor UO_122 (O_122,N_19851,N_19976);
nand UO_123 (O_123,N_19984,N_19882);
nor UO_124 (O_124,N_19866,N_19907);
and UO_125 (O_125,N_19928,N_19976);
nor UO_126 (O_126,N_19950,N_19997);
nor UO_127 (O_127,N_19899,N_19999);
nor UO_128 (O_128,N_19950,N_19877);
nand UO_129 (O_129,N_19965,N_19890);
or UO_130 (O_130,N_19879,N_19869);
or UO_131 (O_131,N_19987,N_19929);
or UO_132 (O_132,N_19997,N_19940);
nor UO_133 (O_133,N_19847,N_19869);
or UO_134 (O_134,N_19988,N_19957);
nand UO_135 (O_135,N_19861,N_19911);
xor UO_136 (O_136,N_19966,N_19929);
nor UO_137 (O_137,N_19879,N_19897);
and UO_138 (O_138,N_19963,N_19852);
or UO_139 (O_139,N_19989,N_19904);
nor UO_140 (O_140,N_19939,N_19923);
nand UO_141 (O_141,N_19999,N_19929);
nor UO_142 (O_142,N_19895,N_19900);
nand UO_143 (O_143,N_19947,N_19958);
and UO_144 (O_144,N_19852,N_19946);
or UO_145 (O_145,N_19862,N_19850);
xnor UO_146 (O_146,N_19942,N_19951);
xnor UO_147 (O_147,N_19995,N_19961);
and UO_148 (O_148,N_19954,N_19967);
nor UO_149 (O_149,N_19877,N_19841);
nor UO_150 (O_150,N_19959,N_19866);
xor UO_151 (O_151,N_19960,N_19989);
or UO_152 (O_152,N_19882,N_19851);
nand UO_153 (O_153,N_19877,N_19948);
or UO_154 (O_154,N_19942,N_19867);
xnor UO_155 (O_155,N_19899,N_19872);
or UO_156 (O_156,N_19942,N_19915);
and UO_157 (O_157,N_19896,N_19893);
or UO_158 (O_158,N_19979,N_19983);
nand UO_159 (O_159,N_19954,N_19908);
xor UO_160 (O_160,N_19872,N_19857);
nor UO_161 (O_161,N_19970,N_19900);
nand UO_162 (O_162,N_19960,N_19850);
nor UO_163 (O_163,N_19847,N_19959);
or UO_164 (O_164,N_19855,N_19866);
or UO_165 (O_165,N_19912,N_19962);
nor UO_166 (O_166,N_19859,N_19955);
or UO_167 (O_167,N_19977,N_19946);
nor UO_168 (O_168,N_19941,N_19879);
or UO_169 (O_169,N_19938,N_19929);
or UO_170 (O_170,N_19973,N_19904);
or UO_171 (O_171,N_19871,N_19985);
and UO_172 (O_172,N_19897,N_19906);
nand UO_173 (O_173,N_19862,N_19962);
nor UO_174 (O_174,N_19844,N_19846);
xor UO_175 (O_175,N_19966,N_19854);
and UO_176 (O_176,N_19958,N_19986);
nor UO_177 (O_177,N_19945,N_19845);
xor UO_178 (O_178,N_19962,N_19941);
or UO_179 (O_179,N_19889,N_19914);
or UO_180 (O_180,N_19920,N_19903);
nor UO_181 (O_181,N_19982,N_19977);
xnor UO_182 (O_182,N_19971,N_19972);
nand UO_183 (O_183,N_19885,N_19905);
nand UO_184 (O_184,N_19911,N_19877);
nand UO_185 (O_185,N_19872,N_19897);
and UO_186 (O_186,N_19905,N_19845);
xnor UO_187 (O_187,N_19845,N_19927);
or UO_188 (O_188,N_19993,N_19990);
nand UO_189 (O_189,N_19982,N_19975);
xor UO_190 (O_190,N_19963,N_19916);
nor UO_191 (O_191,N_19852,N_19842);
and UO_192 (O_192,N_19937,N_19940);
and UO_193 (O_193,N_19968,N_19932);
or UO_194 (O_194,N_19860,N_19929);
xnor UO_195 (O_195,N_19858,N_19956);
nor UO_196 (O_196,N_19990,N_19881);
or UO_197 (O_197,N_19938,N_19983);
or UO_198 (O_198,N_19856,N_19967);
nand UO_199 (O_199,N_19941,N_19859);
nor UO_200 (O_200,N_19923,N_19845);
nand UO_201 (O_201,N_19996,N_19871);
or UO_202 (O_202,N_19924,N_19858);
xor UO_203 (O_203,N_19978,N_19973);
and UO_204 (O_204,N_19981,N_19899);
nor UO_205 (O_205,N_19904,N_19930);
nand UO_206 (O_206,N_19918,N_19883);
nand UO_207 (O_207,N_19919,N_19961);
or UO_208 (O_208,N_19964,N_19865);
nand UO_209 (O_209,N_19924,N_19850);
and UO_210 (O_210,N_19986,N_19906);
nand UO_211 (O_211,N_19926,N_19916);
xnor UO_212 (O_212,N_19859,N_19875);
nand UO_213 (O_213,N_19850,N_19955);
and UO_214 (O_214,N_19987,N_19878);
or UO_215 (O_215,N_19860,N_19877);
and UO_216 (O_216,N_19892,N_19968);
or UO_217 (O_217,N_19933,N_19973);
xor UO_218 (O_218,N_19868,N_19853);
xnor UO_219 (O_219,N_19987,N_19842);
xor UO_220 (O_220,N_19941,N_19975);
nor UO_221 (O_221,N_19871,N_19921);
or UO_222 (O_222,N_19872,N_19856);
nand UO_223 (O_223,N_19875,N_19869);
and UO_224 (O_224,N_19876,N_19966);
nor UO_225 (O_225,N_19958,N_19882);
nand UO_226 (O_226,N_19982,N_19941);
nand UO_227 (O_227,N_19919,N_19900);
xnor UO_228 (O_228,N_19843,N_19944);
nor UO_229 (O_229,N_19904,N_19985);
nand UO_230 (O_230,N_19944,N_19988);
nor UO_231 (O_231,N_19887,N_19905);
nand UO_232 (O_232,N_19988,N_19857);
or UO_233 (O_233,N_19892,N_19998);
or UO_234 (O_234,N_19924,N_19844);
nand UO_235 (O_235,N_19988,N_19853);
nor UO_236 (O_236,N_19859,N_19912);
xnor UO_237 (O_237,N_19857,N_19950);
or UO_238 (O_238,N_19919,N_19882);
nor UO_239 (O_239,N_19841,N_19951);
and UO_240 (O_240,N_19929,N_19906);
or UO_241 (O_241,N_19896,N_19996);
nor UO_242 (O_242,N_19980,N_19977);
or UO_243 (O_243,N_19914,N_19846);
and UO_244 (O_244,N_19996,N_19899);
and UO_245 (O_245,N_19984,N_19938);
or UO_246 (O_246,N_19968,N_19907);
and UO_247 (O_247,N_19991,N_19965);
and UO_248 (O_248,N_19897,N_19954);
and UO_249 (O_249,N_19879,N_19988);
nand UO_250 (O_250,N_19979,N_19851);
nand UO_251 (O_251,N_19956,N_19903);
nor UO_252 (O_252,N_19895,N_19851);
nand UO_253 (O_253,N_19873,N_19969);
xnor UO_254 (O_254,N_19950,N_19964);
or UO_255 (O_255,N_19955,N_19917);
nor UO_256 (O_256,N_19952,N_19997);
nor UO_257 (O_257,N_19914,N_19899);
or UO_258 (O_258,N_19866,N_19942);
xor UO_259 (O_259,N_19964,N_19913);
nor UO_260 (O_260,N_19853,N_19881);
nand UO_261 (O_261,N_19900,N_19855);
or UO_262 (O_262,N_19913,N_19925);
xnor UO_263 (O_263,N_19844,N_19864);
nand UO_264 (O_264,N_19940,N_19904);
nor UO_265 (O_265,N_19982,N_19857);
xnor UO_266 (O_266,N_19919,N_19869);
nor UO_267 (O_267,N_19996,N_19854);
xor UO_268 (O_268,N_19918,N_19917);
nand UO_269 (O_269,N_19970,N_19873);
nand UO_270 (O_270,N_19846,N_19949);
and UO_271 (O_271,N_19897,N_19912);
nand UO_272 (O_272,N_19981,N_19895);
xnor UO_273 (O_273,N_19863,N_19960);
and UO_274 (O_274,N_19875,N_19971);
nand UO_275 (O_275,N_19859,N_19971);
nor UO_276 (O_276,N_19937,N_19895);
nor UO_277 (O_277,N_19942,N_19929);
or UO_278 (O_278,N_19967,N_19991);
xnor UO_279 (O_279,N_19876,N_19847);
and UO_280 (O_280,N_19849,N_19884);
nand UO_281 (O_281,N_19897,N_19951);
and UO_282 (O_282,N_19942,N_19989);
and UO_283 (O_283,N_19876,N_19926);
nor UO_284 (O_284,N_19963,N_19925);
and UO_285 (O_285,N_19894,N_19976);
or UO_286 (O_286,N_19914,N_19917);
xnor UO_287 (O_287,N_19958,N_19996);
and UO_288 (O_288,N_19919,N_19931);
nor UO_289 (O_289,N_19866,N_19891);
nor UO_290 (O_290,N_19999,N_19868);
or UO_291 (O_291,N_19897,N_19924);
and UO_292 (O_292,N_19929,N_19849);
and UO_293 (O_293,N_19950,N_19943);
or UO_294 (O_294,N_19982,N_19928);
nand UO_295 (O_295,N_19849,N_19904);
nor UO_296 (O_296,N_19844,N_19981);
and UO_297 (O_297,N_19863,N_19867);
nand UO_298 (O_298,N_19870,N_19881);
and UO_299 (O_299,N_19973,N_19959);
nor UO_300 (O_300,N_19991,N_19885);
xor UO_301 (O_301,N_19847,N_19893);
xnor UO_302 (O_302,N_19926,N_19874);
nand UO_303 (O_303,N_19962,N_19913);
nor UO_304 (O_304,N_19925,N_19872);
xnor UO_305 (O_305,N_19933,N_19895);
nor UO_306 (O_306,N_19886,N_19983);
nor UO_307 (O_307,N_19945,N_19869);
and UO_308 (O_308,N_19861,N_19876);
and UO_309 (O_309,N_19871,N_19853);
nor UO_310 (O_310,N_19906,N_19937);
and UO_311 (O_311,N_19901,N_19875);
and UO_312 (O_312,N_19924,N_19988);
nor UO_313 (O_313,N_19890,N_19864);
and UO_314 (O_314,N_19870,N_19987);
nand UO_315 (O_315,N_19867,N_19959);
nor UO_316 (O_316,N_19987,N_19967);
or UO_317 (O_317,N_19935,N_19894);
nor UO_318 (O_318,N_19918,N_19948);
nand UO_319 (O_319,N_19855,N_19979);
and UO_320 (O_320,N_19995,N_19868);
xor UO_321 (O_321,N_19932,N_19904);
or UO_322 (O_322,N_19949,N_19958);
nor UO_323 (O_323,N_19865,N_19943);
or UO_324 (O_324,N_19990,N_19975);
nor UO_325 (O_325,N_19895,N_19926);
xor UO_326 (O_326,N_19986,N_19954);
and UO_327 (O_327,N_19890,N_19939);
and UO_328 (O_328,N_19967,N_19849);
nand UO_329 (O_329,N_19922,N_19891);
or UO_330 (O_330,N_19919,N_19966);
and UO_331 (O_331,N_19989,N_19945);
or UO_332 (O_332,N_19887,N_19974);
nand UO_333 (O_333,N_19912,N_19888);
nor UO_334 (O_334,N_19863,N_19897);
xor UO_335 (O_335,N_19871,N_19882);
nor UO_336 (O_336,N_19961,N_19950);
nand UO_337 (O_337,N_19999,N_19869);
xor UO_338 (O_338,N_19959,N_19864);
or UO_339 (O_339,N_19915,N_19962);
or UO_340 (O_340,N_19891,N_19845);
xor UO_341 (O_341,N_19963,N_19841);
nor UO_342 (O_342,N_19869,N_19930);
nand UO_343 (O_343,N_19961,N_19973);
xnor UO_344 (O_344,N_19902,N_19880);
xor UO_345 (O_345,N_19933,N_19972);
nand UO_346 (O_346,N_19858,N_19840);
or UO_347 (O_347,N_19883,N_19859);
nor UO_348 (O_348,N_19932,N_19849);
and UO_349 (O_349,N_19944,N_19871);
or UO_350 (O_350,N_19964,N_19901);
xor UO_351 (O_351,N_19939,N_19900);
nand UO_352 (O_352,N_19952,N_19930);
nand UO_353 (O_353,N_19985,N_19890);
or UO_354 (O_354,N_19956,N_19939);
xnor UO_355 (O_355,N_19863,N_19938);
or UO_356 (O_356,N_19942,N_19924);
and UO_357 (O_357,N_19960,N_19895);
and UO_358 (O_358,N_19892,N_19918);
nand UO_359 (O_359,N_19883,N_19881);
and UO_360 (O_360,N_19841,N_19852);
and UO_361 (O_361,N_19853,N_19843);
xnor UO_362 (O_362,N_19867,N_19982);
xnor UO_363 (O_363,N_19861,N_19877);
xnor UO_364 (O_364,N_19964,N_19934);
and UO_365 (O_365,N_19878,N_19914);
xnor UO_366 (O_366,N_19866,N_19871);
xor UO_367 (O_367,N_19929,N_19873);
nor UO_368 (O_368,N_19867,N_19860);
xor UO_369 (O_369,N_19844,N_19866);
or UO_370 (O_370,N_19958,N_19995);
nand UO_371 (O_371,N_19993,N_19872);
or UO_372 (O_372,N_19967,N_19869);
nand UO_373 (O_373,N_19973,N_19897);
nand UO_374 (O_374,N_19996,N_19990);
nor UO_375 (O_375,N_19971,N_19898);
xnor UO_376 (O_376,N_19878,N_19964);
nand UO_377 (O_377,N_19918,N_19890);
or UO_378 (O_378,N_19873,N_19890);
nor UO_379 (O_379,N_19864,N_19854);
xnor UO_380 (O_380,N_19976,N_19884);
or UO_381 (O_381,N_19926,N_19924);
nand UO_382 (O_382,N_19928,N_19924);
or UO_383 (O_383,N_19984,N_19982);
nor UO_384 (O_384,N_19843,N_19856);
nand UO_385 (O_385,N_19963,N_19927);
or UO_386 (O_386,N_19875,N_19917);
or UO_387 (O_387,N_19977,N_19974);
nor UO_388 (O_388,N_19980,N_19902);
and UO_389 (O_389,N_19941,N_19851);
nor UO_390 (O_390,N_19859,N_19956);
nand UO_391 (O_391,N_19880,N_19892);
nor UO_392 (O_392,N_19857,N_19953);
nor UO_393 (O_393,N_19936,N_19871);
xor UO_394 (O_394,N_19898,N_19940);
or UO_395 (O_395,N_19861,N_19858);
nor UO_396 (O_396,N_19900,N_19971);
xnor UO_397 (O_397,N_19864,N_19994);
xor UO_398 (O_398,N_19950,N_19886);
xor UO_399 (O_399,N_19977,N_19886);
xnor UO_400 (O_400,N_19862,N_19919);
or UO_401 (O_401,N_19989,N_19939);
nand UO_402 (O_402,N_19906,N_19840);
and UO_403 (O_403,N_19917,N_19999);
or UO_404 (O_404,N_19848,N_19912);
nor UO_405 (O_405,N_19867,N_19994);
or UO_406 (O_406,N_19851,N_19944);
nor UO_407 (O_407,N_19891,N_19948);
xor UO_408 (O_408,N_19962,N_19994);
nor UO_409 (O_409,N_19961,N_19945);
nor UO_410 (O_410,N_19938,N_19852);
xnor UO_411 (O_411,N_19946,N_19876);
xnor UO_412 (O_412,N_19972,N_19979);
and UO_413 (O_413,N_19915,N_19952);
nand UO_414 (O_414,N_19863,N_19978);
and UO_415 (O_415,N_19977,N_19928);
nand UO_416 (O_416,N_19981,N_19842);
and UO_417 (O_417,N_19996,N_19855);
nand UO_418 (O_418,N_19956,N_19947);
nand UO_419 (O_419,N_19998,N_19994);
and UO_420 (O_420,N_19994,N_19959);
xor UO_421 (O_421,N_19845,N_19941);
nor UO_422 (O_422,N_19977,N_19922);
nand UO_423 (O_423,N_19913,N_19989);
or UO_424 (O_424,N_19944,N_19996);
xnor UO_425 (O_425,N_19954,N_19947);
or UO_426 (O_426,N_19872,N_19845);
nor UO_427 (O_427,N_19847,N_19930);
nor UO_428 (O_428,N_19969,N_19850);
or UO_429 (O_429,N_19949,N_19847);
nor UO_430 (O_430,N_19914,N_19842);
or UO_431 (O_431,N_19919,N_19968);
and UO_432 (O_432,N_19848,N_19890);
and UO_433 (O_433,N_19997,N_19938);
nand UO_434 (O_434,N_19950,N_19856);
or UO_435 (O_435,N_19850,N_19977);
or UO_436 (O_436,N_19927,N_19885);
nand UO_437 (O_437,N_19932,N_19885);
and UO_438 (O_438,N_19937,N_19873);
or UO_439 (O_439,N_19876,N_19932);
and UO_440 (O_440,N_19878,N_19877);
and UO_441 (O_441,N_19872,N_19892);
nand UO_442 (O_442,N_19863,N_19869);
nand UO_443 (O_443,N_19956,N_19981);
or UO_444 (O_444,N_19866,N_19947);
nor UO_445 (O_445,N_19911,N_19946);
xnor UO_446 (O_446,N_19848,N_19953);
and UO_447 (O_447,N_19857,N_19943);
or UO_448 (O_448,N_19959,N_19848);
nor UO_449 (O_449,N_19937,N_19905);
nand UO_450 (O_450,N_19889,N_19869);
xnor UO_451 (O_451,N_19923,N_19973);
nand UO_452 (O_452,N_19894,N_19852);
or UO_453 (O_453,N_19958,N_19902);
or UO_454 (O_454,N_19843,N_19924);
nand UO_455 (O_455,N_19930,N_19883);
xor UO_456 (O_456,N_19925,N_19869);
or UO_457 (O_457,N_19952,N_19913);
xor UO_458 (O_458,N_19931,N_19877);
xnor UO_459 (O_459,N_19942,N_19969);
nor UO_460 (O_460,N_19884,N_19861);
nand UO_461 (O_461,N_19978,N_19999);
nor UO_462 (O_462,N_19993,N_19950);
xnor UO_463 (O_463,N_19920,N_19866);
and UO_464 (O_464,N_19935,N_19926);
or UO_465 (O_465,N_19841,N_19998);
or UO_466 (O_466,N_19902,N_19979);
or UO_467 (O_467,N_19994,N_19845);
xnor UO_468 (O_468,N_19944,N_19934);
xor UO_469 (O_469,N_19919,N_19986);
nand UO_470 (O_470,N_19873,N_19988);
or UO_471 (O_471,N_19858,N_19882);
and UO_472 (O_472,N_19964,N_19907);
and UO_473 (O_473,N_19957,N_19932);
nand UO_474 (O_474,N_19952,N_19962);
and UO_475 (O_475,N_19952,N_19928);
xnor UO_476 (O_476,N_19984,N_19861);
nor UO_477 (O_477,N_19972,N_19841);
nand UO_478 (O_478,N_19972,N_19922);
or UO_479 (O_479,N_19916,N_19931);
nor UO_480 (O_480,N_19918,N_19990);
nor UO_481 (O_481,N_19993,N_19957);
xnor UO_482 (O_482,N_19965,N_19993);
nor UO_483 (O_483,N_19942,N_19945);
nor UO_484 (O_484,N_19995,N_19951);
nand UO_485 (O_485,N_19914,N_19864);
nand UO_486 (O_486,N_19982,N_19861);
and UO_487 (O_487,N_19890,N_19928);
and UO_488 (O_488,N_19858,N_19968);
or UO_489 (O_489,N_19876,N_19909);
nor UO_490 (O_490,N_19935,N_19854);
or UO_491 (O_491,N_19893,N_19956);
or UO_492 (O_492,N_19951,N_19962);
xor UO_493 (O_493,N_19996,N_19934);
nand UO_494 (O_494,N_19920,N_19995);
nand UO_495 (O_495,N_19913,N_19918);
and UO_496 (O_496,N_19988,N_19942);
or UO_497 (O_497,N_19949,N_19933);
and UO_498 (O_498,N_19883,N_19955);
nor UO_499 (O_499,N_19901,N_19937);
and UO_500 (O_500,N_19971,N_19878);
nand UO_501 (O_501,N_19954,N_19896);
nand UO_502 (O_502,N_19933,N_19976);
nor UO_503 (O_503,N_19934,N_19984);
nand UO_504 (O_504,N_19960,N_19965);
and UO_505 (O_505,N_19891,N_19852);
and UO_506 (O_506,N_19910,N_19851);
nand UO_507 (O_507,N_19958,N_19876);
nand UO_508 (O_508,N_19909,N_19845);
and UO_509 (O_509,N_19914,N_19946);
xnor UO_510 (O_510,N_19841,N_19858);
nor UO_511 (O_511,N_19912,N_19874);
nand UO_512 (O_512,N_19962,N_19986);
nor UO_513 (O_513,N_19871,N_19904);
xor UO_514 (O_514,N_19923,N_19971);
xnor UO_515 (O_515,N_19948,N_19928);
xnor UO_516 (O_516,N_19846,N_19939);
and UO_517 (O_517,N_19969,N_19955);
nor UO_518 (O_518,N_19866,N_19889);
or UO_519 (O_519,N_19852,N_19854);
xnor UO_520 (O_520,N_19899,N_19911);
xnor UO_521 (O_521,N_19944,N_19905);
nor UO_522 (O_522,N_19946,N_19861);
or UO_523 (O_523,N_19987,N_19989);
xnor UO_524 (O_524,N_19879,N_19850);
xnor UO_525 (O_525,N_19979,N_19913);
and UO_526 (O_526,N_19893,N_19912);
nor UO_527 (O_527,N_19844,N_19965);
nor UO_528 (O_528,N_19985,N_19937);
and UO_529 (O_529,N_19929,N_19855);
or UO_530 (O_530,N_19947,N_19997);
xnor UO_531 (O_531,N_19886,N_19894);
nand UO_532 (O_532,N_19840,N_19845);
or UO_533 (O_533,N_19865,N_19895);
nand UO_534 (O_534,N_19886,N_19989);
xnor UO_535 (O_535,N_19842,N_19923);
and UO_536 (O_536,N_19973,N_19907);
or UO_537 (O_537,N_19952,N_19929);
nand UO_538 (O_538,N_19896,N_19939);
nand UO_539 (O_539,N_19981,N_19845);
xnor UO_540 (O_540,N_19907,N_19938);
or UO_541 (O_541,N_19899,N_19855);
nand UO_542 (O_542,N_19864,N_19896);
xnor UO_543 (O_543,N_19937,N_19861);
nand UO_544 (O_544,N_19962,N_19891);
nor UO_545 (O_545,N_19957,N_19927);
nand UO_546 (O_546,N_19904,N_19982);
or UO_547 (O_547,N_19885,N_19894);
nor UO_548 (O_548,N_19930,N_19975);
and UO_549 (O_549,N_19863,N_19879);
and UO_550 (O_550,N_19943,N_19959);
nor UO_551 (O_551,N_19937,N_19887);
xnor UO_552 (O_552,N_19975,N_19932);
nand UO_553 (O_553,N_19916,N_19841);
nand UO_554 (O_554,N_19930,N_19966);
or UO_555 (O_555,N_19845,N_19861);
and UO_556 (O_556,N_19920,N_19892);
and UO_557 (O_557,N_19991,N_19977);
nor UO_558 (O_558,N_19978,N_19915);
nor UO_559 (O_559,N_19887,N_19949);
xor UO_560 (O_560,N_19986,N_19847);
or UO_561 (O_561,N_19987,N_19869);
nor UO_562 (O_562,N_19973,N_19882);
or UO_563 (O_563,N_19956,N_19986);
or UO_564 (O_564,N_19858,N_19907);
xor UO_565 (O_565,N_19875,N_19950);
nand UO_566 (O_566,N_19938,N_19933);
or UO_567 (O_567,N_19841,N_19866);
nand UO_568 (O_568,N_19990,N_19899);
xnor UO_569 (O_569,N_19931,N_19939);
or UO_570 (O_570,N_19960,N_19844);
or UO_571 (O_571,N_19936,N_19933);
nand UO_572 (O_572,N_19995,N_19918);
nor UO_573 (O_573,N_19972,N_19881);
nand UO_574 (O_574,N_19851,N_19987);
or UO_575 (O_575,N_19946,N_19841);
or UO_576 (O_576,N_19869,N_19886);
and UO_577 (O_577,N_19917,N_19992);
nor UO_578 (O_578,N_19938,N_19967);
nand UO_579 (O_579,N_19891,N_19974);
xor UO_580 (O_580,N_19954,N_19963);
nand UO_581 (O_581,N_19906,N_19915);
and UO_582 (O_582,N_19891,N_19862);
nand UO_583 (O_583,N_19866,N_19876);
nand UO_584 (O_584,N_19983,N_19915);
nor UO_585 (O_585,N_19994,N_19986);
xor UO_586 (O_586,N_19898,N_19951);
nor UO_587 (O_587,N_19930,N_19996);
and UO_588 (O_588,N_19945,N_19875);
nor UO_589 (O_589,N_19927,N_19980);
nand UO_590 (O_590,N_19855,N_19877);
and UO_591 (O_591,N_19986,N_19925);
or UO_592 (O_592,N_19971,N_19967);
nand UO_593 (O_593,N_19845,N_19925);
or UO_594 (O_594,N_19975,N_19886);
nand UO_595 (O_595,N_19963,N_19968);
xnor UO_596 (O_596,N_19932,N_19900);
or UO_597 (O_597,N_19943,N_19955);
xnor UO_598 (O_598,N_19883,N_19853);
and UO_599 (O_599,N_19963,N_19892);
xor UO_600 (O_600,N_19907,N_19958);
nand UO_601 (O_601,N_19899,N_19871);
or UO_602 (O_602,N_19933,N_19996);
nor UO_603 (O_603,N_19891,N_19959);
and UO_604 (O_604,N_19996,N_19891);
nand UO_605 (O_605,N_19917,N_19977);
nor UO_606 (O_606,N_19933,N_19947);
nor UO_607 (O_607,N_19966,N_19917);
xor UO_608 (O_608,N_19916,N_19903);
and UO_609 (O_609,N_19986,N_19854);
or UO_610 (O_610,N_19877,N_19899);
and UO_611 (O_611,N_19998,N_19937);
xnor UO_612 (O_612,N_19875,N_19895);
nor UO_613 (O_613,N_19943,N_19868);
nand UO_614 (O_614,N_19916,N_19978);
or UO_615 (O_615,N_19916,N_19904);
nand UO_616 (O_616,N_19896,N_19992);
and UO_617 (O_617,N_19974,N_19849);
nor UO_618 (O_618,N_19941,N_19887);
xor UO_619 (O_619,N_19841,N_19982);
nor UO_620 (O_620,N_19952,N_19925);
xnor UO_621 (O_621,N_19963,N_19856);
xor UO_622 (O_622,N_19878,N_19909);
or UO_623 (O_623,N_19918,N_19986);
xnor UO_624 (O_624,N_19990,N_19968);
xnor UO_625 (O_625,N_19910,N_19849);
nor UO_626 (O_626,N_19840,N_19944);
or UO_627 (O_627,N_19884,N_19853);
or UO_628 (O_628,N_19903,N_19980);
and UO_629 (O_629,N_19897,N_19885);
or UO_630 (O_630,N_19963,N_19876);
or UO_631 (O_631,N_19988,N_19956);
xor UO_632 (O_632,N_19914,N_19903);
nand UO_633 (O_633,N_19952,N_19943);
nor UO_634 (O_634,N_19979,N_19910);
xor UO_635 (O_635,N_19970,N_19915);
or UO_636 (O_636,N_19994,N_19896);
or UO_637 (O_637,N_19948,N_19983);
and UO_638 (O_638,N_19871,N_19902);
xnor UO_639 (O_639,N_19893,N_19916);
nand UO_640 (O_640,N_19981,N_19930);
xor UO_641 (O_641,N_19932,N_19953);
nor UO_642 (O_642,N_19840,N_19950);
xor UO_643 (O_643,N_19915,N_19875);
and UO_644 (O_644,N_19969,N_19913);
xnor UO_645 (O_645,N_19887,N_19854);
and UO_646 (O_646,N_19941,N_19953);
nand UO_647 (O_647,N_19855,N_19863);
nor UO_648 (O_648,N_19944,N_19954);
or UO_649 (O_649,N_19905,N_19967);
or UO_650 (O_650,N_19976,N_19983);
or UO_651 (O_651,N_19849,N_19978);
nand UO_652 (O_652,N_19922,N_19956);
nor UO_653 (O_653,N_19931,N_19996);
and UO_654 (O_654,N_19925,N_19854);
nor UO_655 (O_655,N_19944,N_19909);
nand UO_656 (O_656,N_19897,N_19974);
xnor UO_657 (O_657,N_19960,N_19941);
nand UO_658 (O_658,N_19900,N_19957);
and UO_659 (O_659,N_19871,N_19982);
or UO_660 (O_660,N_19909,N_19928);
and UO_661 (O_661,N_19852,N_19950);
nand UO_662 (O_662,N_19908,N_19966);
nor UO_663 (O_663,N_19937,N_19914);
or UO_664 (O_664,N_19990,N_19940);
or UO_665 (O_665,N_19919,N_19916);
nor UO_666 (O_666,N_19841,N_19996);
and UO_667 (O_667,N_19960,N_19897);
or UO_668 (O_668,N_19952,N_19908);
or UO_669 (O_669,N_19924,N_19906);
nor UO_670 (O_670,N_19916,N_19894);
and UO_671 (O_671,N_19947,N_19952);
xor UO_672 (O_672,N_19940,N_19869);
xor UO_673 (O_673,N_19904,N_19951);
and UO_674 (O_674,N_19885,N_19920);
nor UO_675 (O_675,N_19846,N_19941);
and UO_676 (O_676,N_19965,N_19964);
and UO_677 (O_677,N_19883,N_19899);
or UO_678 (O_678,N_19991,N_19862);
nand UO_679 (O_679,N_19869,N_19920);
xnor UO_680 (O_680,N_19943,N_19917);
nand UO_681 (O_681,N_19934,N_19973);
nand UO_682 (O_682,N_19904,N_19934);
nand UO_683 (O_683,N_19947,N_19873);
or UO_684 (O_684,N_19969,N_19908);
or UO_685 (O_685,N_19922,N_19898);
or UO_686 (O_686,N_19877,N_19927);
nand UO_687 (O_687,N_19869,N_19878);
and UO_688 (O_688,N_19864,N_19930);
nand UO_689 (O_689,N_19956,N_19948);
nor UO_690 (O_690,N_19948,N_19921);
nand UO_691 (O_691,N_19964,N_19940);
xor UO_692 (O_692,N_19919,N_19928);
xnor UO_693 (O_693,N_19991,N_19884);
xnor UO_694 (O_694,N_19950,N_19982);
nand UO_695 (O_695,N_19894,N_19892);
nor UO_696 (O_696,N_19901,N_19861);
nor UO_697 (O_697,N_19878,N_19946);
nor UO_698 (O_698,N_19857,N_19966);
nand UO_699 (O_699,N_19928,N_19849);
nor UO_700 (O_700,N_19982,N_19873);
nor UO_701 (O_701,N_19985,N_19850);
xor UO_702 (O_702,N_19915,N_19988);
and UO_703 (O_703,N_19935,N_19857);
nand UO_704 (O_704,N_19911,N_19984);
nor UO_705 (O_705,N_19903,N_19987);
and UO_706 (O_706,N_19973,N_19879);
xor UO_707 (O_707,N_19876,N_19989);
nor UO_708 (O_708,N_19925,N_19989);
nor UO_709 (O_709,N_19958,N_19878);
or UO_710 (O_710,N_19941,N_19944);
or UO_711 (O_711,N_19873,N_19887);
or UO_712 (O_712,N_19911,N_19965);
nand UO_713 (O_713,N_19973,N_19889);
or UO_714 (O_714,N_19874,N_19894);
xnor UO_715 (O_715,N_19936,N_19972);
and UO_716 (O_716,N_19937,N_19898);
nand UO_717 (O_717,N_19952,N_19901);
xnor UO_718 (O_718,N_19941,N_19917);
or UO_719 (O_719,N_19859,N_19852);
and UO_720 (O_720,N_19925,N_19975);
nor UO_721 (O_721,N_19995,N_19973);
xor UO_722 (O_722,N_19966,N_19898);
xnor UO_723 (O_723,N_19982,N_19951);
nand UO_724 (O_724,N_19844,N_19885);
and UO_725 (O_725,N_19879,N_19926);
nor UO_726 (O_726,N_19927,N_19867);
nor UO_727 (O_727,N_19978,N_19890);
or UO_728 (O_728,N_19913,N_19868);
xnor UO_729 (O_729,N_19859,N_19998);
xnor UO_730 (O_730,N_19988,N_19977);
xnor UO_731 (O_731,N_19927,N_19923);
nor UO_732 (O_732,N_19983,N_19992);
nand UO_733 (O_733,N_19957,N_19891);
nand UO_734 (O_734,N_19904,N_19991);
and UO_735 (O_735,N_19882,N_19960);
or UO_736 (O_736,N_19915,N_19995);
or UO_737 (O_737,N_19956,N_19957);
xor UO_738 (O_738,N_19894,N_19854);
or UO_739 (O_739,N_19877,N_19984);
xor UO_740 (O_740,N_19912,N_19940);
nor UO_741 (O_741,N_19858,N_19888);
and UO_742 (O_742,N_19852,N_19882);
and UO_743 (O_743,N_19884,N_19955);
or UO_744 (O_744,N_19900,N_19962);
nor UO_745 (O_745,N_19933,N_19860);
xor UO_746 (O_746,N_19901,N_19857);
xnor UO_747 (O_747,N_19885,N_19945);
nand UO_748 (O_748,N_19984,N_19920);
nor UO_749 (O_749,N_19897,N_19862);
and UO_750 (O_750,N_19881,N_19860);
xnor UO_751 (O_751,N_19951,N_19928);
nand UO_752 (O_752,N_19913,N_19851);
nor UO_753 (O_753,N_19930,N_19901);
and UO_754 (O_754,N_19933,N_19992);
nand UO_755 (O_755,N_19941,N_19965);
nand UO_756 (O_756,N_19941,N_19896);
and UO_757 (O_757,N_19919,N_19845);
nor UO_758 (O_758,N_19899,N_19843);
nand UO_759 (O_759,N_19950,N_19913);
nor UO_760 (O_760,N_19845,N_19955);
and UO_761 (O_761,N_19948,N_19988);
xnor UO_762 (O_762,N_19881,N_19856);
and UO_763 (O_763,N_19888,N_19942);
and UO_764 (O_764,N_19899,N_19859);
or UO_765 (O_765,N_19876,N_19943);
or UO_766 (O_766,N_19949,N_19940);
or UO_767 (O_767,N_19947,N_19953);
nor UO_768 (O_768,N_19980,N_19865);
and UO_769 (O_769,N_19844,N_19986);
and UO_770 (O_770,N_19926,N_19992);
and UO_771 (O_771,N_19903,N_19950);
nand UO_772 (O_772,N_19987,N_19874);
nor UO_773 (O_773,N_19964,N_19936);
or UO_774 (O_774,N_19942,N_19919);
nor UO_775 (O_775,N_19903,N_19913);
and UO_776 (O_776,N_19950,N_19992);
and UO_777 (O_777,N_19900,N_19949);
nor UO_778 (O_778,N_19869,N_19913);
xor UO_779 (O_779,N_19921,N_19979);
nand UO_780 (O_780,N_19878,N_19944);
xnor UO_781 (O_781,N_19916,N_19968);
or UO_782 (O_782,N_19992,N_19945);
nand UO_783 (O_783,N_19974,N_19878);
or UO_784 (O_784,N_19912,N_19866);
and UO_785 (O_785,N_19980,N_19870);
and UO_786 (O_786,N_19956,N_19864);
nand UO_787 (O_787,N_19939,N_19928);
xor UO_788 (O_788,N_19903,N_19897);
or UO_789 (O_789,N_19893,N_19946);
nand UO_790 (O_790,N_19942,N_19879);
or UO_791 (O_791,N_19955,N_19880);
and UO_792 (O_792,N_19844,N_19854);
or UO_793 (O_793,N_19996,N_19858);
and UO_794 (O_794,N_19883,N_19867);
xnor UO_795 (O_795,N_19917,N_19882);
or UO_796 (O_796,N_19962,N_19850);
nor UO_797 (O_797,N_19991,N_19896);
nand UO_798 (O_798,N_19995,N_19914);
and UO_799 (O_799,N_19997,N_19955);
and UO_800 (O_800,N_19914,N_19859);
or UO_801 (O_801,N_19924,N_19925);
and UO_802 (O_802,N_19981,N_19912);
xnor UO_803 (O_803,N_19846,N_19848);
nand UO_804 (O_804,N_19864,N_19913);
xor UO_805 (O_805,N_19859,N_19928);
and UO_806 (O_806,N_19938,N_19982);
xnor UO_807 (O_807,N_19999,N_19893);
xnor UO_808 (O_808,N_19883,N_19945);
or UO_809 (O_809,N_19955,N_19844);
xor UO_810 (O_810,N_19892,N_19905);
and UO_811 (O_811,N_19879,N_19875);
or UO_812 (O_812,N_19931,N_19930);
nor UO_813 (O_813,N_19866,N_19956);
and UO_814 (O_814,N_19987,N_19962);
nand UO_815 (O_815,N_19907,N_19975);
nand UO_816 (O_816,N_19982,N_19895);
nand UO_817 (O_817,N_19975,N_19911);
nor UO_818 (O_818,N_19919,N_19953);
xor UO_819 (O_819,N_19966,N_19993);
nand UO_820 (O_820,N_19959,N_19854);
xnor UO_821 (O_821,N_19918,N_19957);
and UO_822 (O_822,N_19860,N_19954);
nand UO_823 (O_823,N_19880,N_19990);
xor UO_824 (O_824,N_19889,N_19882);
and UO_825 (O_825,N_19997,N_19894);
and UO_826 (O_826,N_19931,N_19901);
nand UO_827 (O_827,N_19934,N_19926);
xor UO_828 (O_828,N_19990,N_19879);
nand UO_829 (O_829,N_19949,N_19878);
or UO_830 (O_830,N_19939,N_19848);
and UO_831 (O_831,N_19897,N_19854);
nand UO_832 (O_832,N_19886,N_19931);
and UO_833 (O_833,N_19850,N_19968);
xnor UO_834 (O_834,N_19992,N_19853);
or UO_835 (O_835,N_19967,N_19952);
xor UO_836 (O_836,N_19991,N_19950);
xnor UO_837 (O_837,N_19896,N_19972);
xnor UO_838 (O_838,N_19979,N_19977);
xor UO_839 (O_839,N_19896,N_19936);
nand UO_840 (O_840,N_19975,N_19895);
xor UO_841 (O_841,N_19840,N_19938);
or UO_842 (O_842,N_19979,N_19944);
nand UO_843 (O_843,N_19873,N_19995);
and UO_844 (O_844,N_19977,N_19899);
xor UO_845 (O_845,N_19954,N_19869);
or UO_846 (O_846,N_19856,N_19866);
nor UO_847 (O_847,N_19942,N_19890);
and UO_848 (O_848,N_19854,N_19971);
xor UO_849 (O_849,N_19923,N_19858);
or UO_850 (O_850,N_19913,N_19854);
nor UO_851 (O_851,N_19848,N_19956);
and UO_852 (O_852,N_19840,N_19954);
nor UO_853 (O_853,N_19978,N_19870);
or UO_854 (O_854,N_19888,N_19945);
nand UO_855 (O_855,N_19951,N_19974);
nor UO_856 (O_856,N_19992,N_19952);
and UO_857 (O_857,N_19953,N_19999);
and UO_858 (O_858,N_19915,N_19921);
nor UO_859 (O_859,N_19843,N_19895);
nand UO_860 (O_860,N_19871,N_19857);
or UO_861 (O_861,N_19869,N_19980);
and UO_862 (O_862,N_19998,N_19914);
nand UO_863 (O_863,N_19896,N_19915);
nand UO_864 (O_864,N_19841,N_19892);
nor UO_865 (O_865,N_19859,N_19884);
xnor UO_866 (O_866,N_19924,N_19842);
or UO_867 (O_867,N_19894,N_19897);
nand UO_868 (O_868,N_19887,N_19940);
xor UO_869 (O_869,N_19881,N_19978);
xor UO_870 (O_870,N_19894,N_19949);
or UO_871 (O_871,N_19847,N_19921);
or UO_872 (O_872,N_19929,N_19919);
nand UO_873 (O_873,N_19970,N_19999);
nand UO_874 (O_874,N_19940,N_19875);
nor UO_875 (O_875,N_19968,N_19908);
nand UO_876 (O_876,N_19911,N_19885);
or UO_877 (O_877,N_19894,N_19863);
or UO_878 (O_878,N_19893,N_19958);
or UO_879 (O_879,N_19946,N_19926);
and UO_880 (O_880,N_19993,N_19967);
and UO_881 (O_881,N_19996,N_19872);
nor UO_882 (O_882,N_19957,N_19912);
and UO_883 (O_883,N_19955,N_19847);
or UO_884 (O_884,N_19855,N_19849);
xnor UO_885 (O_885,N_19993,N_19869);
nor UO_886 (O_886,N_19969,N_19907);
and UO_887 (O_887,N_19840,N_19932);
nor UO_888 (O_888,N_19920,N_19863);
nor UO_889 (O_889,N_19962,N_19882);
and UO_890 (O_890,N_19906,N_19846);
nor UO_891 (O_891,N_19847,N_19918);
nor UO_892 (O_892,N_19992,N_19957);
nand UO_893 (O_893,N_19971,N_19989);
or UO_894 (O_894,N_19913,N_19945);
xnor UO_895 (O_895,N_19929,N_19944);
nor UO_896 (O_896,N_19945,N_19994);
xor UO_897 (O_897,N_19940,N_19895);
xnor UO_898 (O_898,N_19909,N_19912);
nor UO_899 (O_899,N_19840,N_19952);
and UO_900 (O_900,N_19881,N_19963);
xnor UO_901 (O_901,N_19937,N_19848);
nand UO_902 (O_902,N_19840,N_19847);
and UO_903 (O_903,N_19890,N_19994);
nand UO_904 (O_904,N_19915,N_19955);
and UO_905 (O_905,N_19965,N_19862);
or UO_906 (O_906,N_19916,N_19886);
nor UO_907 (O_907,N_19899,N_19850);
nand UO_908 (O_908,N_19908,N_19918);
or UO_909 (O_909,N_19849,N_19957);
nand UO_910 (O_910,N_19996,N_19982);
nor UO_911 (O_911,N_19844,N_19951);
nor UO_912 (O_912,N_19917,N_19892);
nor UO_913 (O_913,N_19990,N_19902);
or UO_914 (O_914,N_19842,N_19976);
nand UO_915 (O_915,N_19929,N_19945);
or UO_916 (O_916,N_19939,N_19977);
and UO_917 (O_917,N_19948,N_19990);
nand UO_918 (O_918,N_19889,N_19844);
xor UO_919 (O_919,N_19861,N_19926);
xor UO_920 (O_920,N_19985,N_19991);
nor UO_921 (O_921,N_19922,N_19960);
or UO_922 (O_922,N_19928,N_19846);
nor UO_923 (O_923,N_19928,N_19969);
and UO_924 (O_924,N_19904,N_19971);
nor UO_925 (O_925,N_19856,N_19858);
nand UO_926 (O_926,N_19991,N_19869);
or UO_927 (O_927,N_19968,N_19868);
xor UO_928 (O_928,N_19906,N_19972);
nand UO_929 (O_929,N_19951,N_19933);
or UO_930 (O_930,N_19991,N_19988);
nor UO_931 (O_931,N_19902,N_19864);
nor UO_932 (O_932,N_19943,N_19946);
nand UO_933 (O_933,N_19853,N_19890);
and UO_934 (O_934,N_19975,N_19971);
or UO_935 (O_935,N_19974,N_19943);
and UO_936 (O_936,N_19903,N_19993);
or UO_937 (O_937,N_19917,N_19993);
nor UO_938 (O_938,N_19999,N_19859);
and UO_939 (O_939,N_19971,N_19906);
nor UO_940 (O_940,N_19893,N_19915);
and UO_941 (O_941,N_19850,N_19848);
nand UO_942 (O_942,N_19875,N_19981);
or UO_943 (O_943,N_19872,N_19885);
nand UO_944 (O_944,N_19942,N_19851);
and UO_945 (O_945,N_19955,N_19882);
nor UO_946 (O_946,N_19991,N_19973);
and UO_947 (O_947,N_19866,N_19904);
and UO_948 (O_948,N_19890,N_19871);
and UO_949 (O_949,N_19914,N_19880);
or UO_950 (O_950,N_19863,N_19950);
nand UO_951 (O_951,N_19868,N_19962);
xor UO_952 (O_952,N_19879,N_19967);
and UO_953 (O_953,N_19940,N_19967);
and UO_954 (O_954,N_19840,N_19910);
nand UO_955 (O_955,N_19941,N_19893);
xor UO_956 (O_956,N_19922,N_19997);
nor UO_957 (O_957,N_19941,N_19898);
nand UO_958 (O_958,N_19926,N_19857);
nand UO_959 (O_959,N_19866,N_19986);
or UO_960 (O_960,N_19968,N_19875);
and UO_961 (O_961,N_19904,N_19988);
or UO_962 (O_962,N_19923,N_19949);
nand UO_963 (O_963,N_19852,N_19884);
xor UO_964 (O_964,N_19979,N_19904);
nand UO_965 (O_965,N_19893,N_19965);
nor UO_966 (O_966,N_19992,N_19918);
xnor UO_967 (O_967,N_19975,N_19989);
xnor UO_968 (O_968,N_19948,N_19912);
xnor UO_969 (O_969,N_19971,N_19952);
xor UO_970 (O_970,N_19977,N_19910);
nor UO_971 (O_971,N_19924,N_19880);
or UO_972 (O_972,N_19913,N_19955);
and UO_973 (O_973,N_19916,N_19957);
nand UO_974 (O_974,N_19906,N_19957);
and UO_975 (O_975,N_19970,N_19964);
or UO_976 (O_976,N_19979,N_19877);
or UO_977 (O_977,N_19847,N_19913);
and UO_978 (O_978,N_19850,N_19888);
nand UO_979 (O_979,N_19907,N_19936);
or UO_980 (O_980,N_19886,N_19891);
xnor UO_981 (O_981,N_19892,N_19914);
nor UO_982 (O_982,N_19859,N_19860);
nand UO_983 (O_983,N_19955,N_19895);
or UO_984 (O_984,N_19857,N_19846);
nand UO_985 (O_985,N_19985,N_19950);
xnor UO_986 (O_986,N_19865,N_19992);
nor UO_987 (O_987,N_19893,N_19938);
nand UO_988 (O_988,N_19964,N_19866);
and UO_989 (O_989,N_19995,N_19892);
nor UO_990 (O_990,N_19902,N_19900);
xor UO_991 (O_991,N_19848,N_19872);
and UO_992 (O_992,N_19947,N_19899);
nor UO_993 (O_993,N_19987,N_19982);
and UO_994 (O_994,N_19894,N_19913);
and UO_995 (O_995,N_19842,N_19995);
and UO_996 (O_996,N_19987,N_19868);
nand UO_997 (O_997,N_19990,N_19917);
xnor UO_998 (O_998,N_19909,N_19843);
xnor UO_999 (O_999,N_19870,N_19938);
or UO_1000 (O_1000,N_19943,N_19958);
nand UO_1001 (O_1001,N_19940,N_19933);
nand UO_1002 (O_1002,N_19932,N_19917);
or UO_1003 (O_1003,N_19942,N_19978);
nand UO_1004 (O_1004,N_19921,N_19956);
and UO_1005 (O_1005,N_19910,N_19988);
nor UO_1006 (O_1006,N_19859,N_19933);
xnor UO_1007 (O_1007,N_19993,N_19840);
or UO_1008 (O_1008,N_19844,N_19850);
nand UO_1009 (O_1009,N_19928,N_19971);
and UO_1010 (O_1010,N_19849,N_19942);
nand UO_1011 (O_1011,N_19866,N_19993);
xor UO_1012 (O_1012,N_19996,N_19867);
and UO_1013 (O_1013,N_19914,N_19938);
xnor UO_1014 (O_1014,N_19958,N_19942);
nand UO_1015 (O_1015,N_19922,N_19921);
nand UO_1016 (O_1016,N_19845,N_19982);
nand UO_1017 (O_1017,N_19931,N_19972);
or UO_1018 (O_1018,N_19886,N_19876);
and UO_1019 (O_1019,N_19845,N_19938);
nand UO_1020 (O_1020,N_19857,N_19896);
and UO_1021 (O_1021,N_19895,N_19860);
xor UO_1022 (O_1022,N_19904,N_19844);
nor UO_1023 (O_1023,N_19868,N_19907);
nand UO_1024 (O_1024,N_19882,N_19904);
nor UO_1025 (O_1025,N_19965,N_19989);
and UO_1026 (O_1026,N_19863,N_19971);
or UO_1027 (O_1027,N_19988,N_19912);
nand UO_1028 (O_1028,N_19845,N_19918);
or UO_1029 (O_1029,N_19978,N_19971);
xor UO_1030 (O_1030,N_19883,N_19900);
xor UO_1031 (O_1031,N_19897,N_19918);
nand UO_1032 (O_1032,N_19880,N_19860);
and UO_1033 (O_1033,N_19974,N_19948);
and UO_1034 (O_1034,N_19900,N_19873);
or UO_1035 (O_1035,N_19978,N_19968);
nand UO_1036 (O_1036,N_19846,N_19852);
xnor UO_1037 (O_1037,N_19980,N_19974);
or UO_1038 (O_1038,N_19908,N_19912);
nor UO_1039 (O_1039,N_19935,N_19913);
and UO_1040 (O_1040,N_19963,N_19846);
xnor UO_1041 (O_1041,N_19842,N_19913);
xor UO_1042 (O_1042,N_19986,N_19901);
and UO_1043 (O_1043,N_19905,N_19859);
and UO_1044 (O_1044,N_19873,N_19936);
or UO_1045 (O_1045,N_19908,N_19983);
or UO_1046 (O_1046,N_19989,N_19934);
or UO_1047 (O_1047,N_19921,N_19873);
or UO_1048 (O_1048,N_19904,N_19962);
and UO_1049 (O_1049,N_19898,N_19860);
nor UO_1050 (O_1050,N_19909,N_19978);
xnor UO_1051 (O_1051,N_19938,N_19868);
nand UO_1052 (O_1052,N_19967,N_19859);
and UO_1053 (O_1053,N_19988,N_19876);
nand UO_1054 (O_1054,N_19920,N_19857);
and UO_1055 (O_1055,N_19918,N_19929);
xnor UO_1056 (O_1056,N_19960,N_19876);
and UO_1057 (O_1057,N_19844,N_19862);
or UO_1058 (O_1058,N_19996,N_19991);
or UO_1059 (O_1059,N_19898,N_19955);
and UO_1060 (O_1060,N_19935,N_19987);
or UO_1061 (O_1061,N_19994,N_19876);
nor UO_1062 (O_1062,N_19927,N_19900);
and UO_1063 (O_1063,N_19885,N_19907);
xor UO_1064 (O_1064,N_19923,N_19946);
xnor UO_1065 (O_1065,N_19965,N_19851);
nand UO_1066 (O_1066,N_19927,N_19925);
and UO_1067 (O_1067,N_19899,N_19939);
or UO_1068 (O_1068,N_19872,N_19919);
nor UO_1069 (O_1069,N_19984,N_19936);
and UO_1070 (O_1070,N_19876,N_19951);
xor UO_1071 (O_1071,N_19937,N_19929);
nor UO_1072 (O_1072,N_19872,N_19904);
or UO_1073 (O_1073,N_19885,N_19982);
nor UO_1074 (O_1074,N_19950,N_19966);
or UO_1075 (O_1075,N_19865,N_19882);
or UO_1076 (O_1076,N_19877,N_19867);
and UO_1077 (O_1077,N_19848,N_19908);
nand UO_1078 (O_1078,N_19985,N_19963);
or UO_1079 (O_1079,N_19935,N_19925);
nor UO_1080 (O_1080,N_19927,N_19881);
xnor UO_1081 (O_1081,N_19899,N_19898);
and UO_1082 (O_1082,N_19890,N_19990);
xor UO_1083 (O_1083,N_19963,N_19844);
or UO_1084 (O_1084,N_19870,N_19890);
xnor UO_1085 (O_1085,N_19931,N_19869);
or UO_1086 (O_1086,N_19985,N_19943);
nand UO_1087 (O_1087,N_19915,N_19941);
and UO_1088 (O_1088,N_19869,N_19924);
nor UO_1089 (O_1089,N_19883,N_19889);
nor UO_1090 (O_1090,N_19921,N_19844);
nor UO_1091 (O_1091,N_19887,N_19880);
and UO_1092 (O_1092,N_19960,N_19867);
or UO_1093 (O_1093,N_19960,N_19995);
xnor UO_1094 (O_1094,N_19849,N_19851);
nor UO_1095 (O_1095,N_19840,N_19951);
and UO_1096 (O_1096,N_19953,N_19847);
xor UO_1097 (O_1097,N_19927,N_19976);
nor UO_1098 (O_1098,N_19881,N_19947);
or UO_1099 (O_1099,N_19866,N_19842);
nand UO_1100 (O_1100,N_19906,N_19939);
and UO_1101 (O_1101,N_19996,N_19952);
or UO_1102 (O_1102,N_19886,N_19926);
nand UO_1103 (O_1103,N_19907,N_19896);
xor UO_1104 (O_1104,N_19986,N_19963);
nand UO_1105 (O_1105,N_19959,N_19951);
or UO_1106 (O_1106,N_19899,N_19965);
or UO_1107 (O_1107,N_19930,N_19991);
nand UO_1108 (O_1108,N_19936,N_19877);
nand UO_1109 (O_1109,N_19880,N_19897);
nor UO_1110 (O_1110,N_19877,N_19903);
xnor UO_1111 (O_1111,N_19909,N_19923);
nand UO_1112 (O_1112,N_19962,N_19841);
or UO_1113 (O_1113,N_19986,N_19940);
nand UO_1114 (O_1114,N_19940,N_19910);
xor UO_1115 (O_1115,N_19910,N_19872);
xor UO_1116 (O_1116,N_19976,N_19877);
nor UO_1117 (O_1117,N_19981,N_19872);
nand UO_1118 (O_1118,N_19978,N_19894);
nand UO_1119 (O_1119,N_19946,N_19980);
and UO_1120 (O_1120,N_19900,N_19908);
xnor UO_1121 (O_1121,N_19898,N_19921);
xor UO_1122 (O_1122,N_19907,N_19909);
or UO_1123 (O_1123,N_19932,N_19857);
nor UO_1124 (O_1124,N_19946,N_19940);
nor UO_1125 (O_1125,N_19856,N_19909);
and UO_1126 (O_1126,N_19999,N_19987);
nand UO_1127 (O_1127,N_19896,N_19917);
nor UO_1128 (O_1128,N_19898,N_19995);
nor UO_1129 (O_1129,N_19908,N_19860);
and UO_1130 (O_1130,N_19961,N_19991);
nor UO_1131 (O_1131,N_19979,N_19856);
or UO_1132 (O_1132,N_19883,N_19961);
or UO_1133 (O_1133,N_19934,N_19890);
xnor UO_1134 (O_1134,N_19937,N_19888);
nor UO_1135 (O_1135,N_19869,N_19970);
xnor UO_1136 (O_1136,N_19863,N_19926);
xnor UO_1137 (O_1137,N_19975,N_19950);
nand UO_1138 (O_1138,N_19889,N_19900);
nor UO_1139 (O_1139,N_19912,N_19911);
nor UO_1140 (O_1140,N_19867,N_19987);
or UO_1141 (O_1141,N_19919,N_19846);
nand UO_1142 (O_1142,N_19864,N_19918);
nand UO_1143 (O_1143,N_19844,N_19914);
nand UO_1144 (O_1144,N_19910,N_19995);
or UO_1145 (O_1145,N_19933,N_19994);
or UO_1146 (O_1146,N_19989,N_19866);
nor UO_1147 (O_1147,N_19840,N_19890);
or UO_1148 (O_1148,N_19865,N_19958);
or UO_1149 (O_1149,N_19932,N_19958);
nand UO_1150 (O_1150,N_19954,N_19924);
nand UO_1151 (O_1151,N_19968,N_19840);
and UO_1152 (O_1152,N_19846,N_19951);
nand UO_1153 (O_1153,N_19909,N_19914);
or UO_1154 (O_1154,N_19987,N_19897);
nand UO_1155 (O_1155,N_19954,N_19945);
nor UO_1156 (O_1156,N_19901,N_19912);
nor UO_1157 (O_1157,N_19960,N_19918);
xnor UO_1158 (O_1158,N_19978,N_19887);
xnor UO_1159 (O_1159,N_19915,N_19923);
and UO_1160 (O_1160,N_19918,N_19950);
xnor UO_1161 (O_1161,N_19939,N_19942);
and UO_1162 (O_1162,N_19914,N_19873);
nor UO_1163 (O_1163,N_19889,N_19881);
xnor UO_1164 (O_1164,N_19915,N_19940);
or UO_1165 (O_1165,N_19891,N_19990);
and UO_1166 (O_1166,N_19849,N_19857);
or UO_1167 (O_1167,N_19925,N_19914);
nor UO_1168 (O_1168,N_19963,N_19874);
nor UO_1169 (O_1169,N_19941,N_19854);
xor UO_1170 (O_1170,N_19996,N_19962);
nor UO_1171 (O_1171,N_19982,N_19858);
or UO_1172 (O_1172,N_19944,N_19875);
nand UO_1173 (O_1173,N_19894,N_19972);
xor UO_1174 (O_1174,N_19852,N_19849);
or UO_1175 (O_1175,N_19998,N_19996);
or UO_1176 (O_1176,N_19871,N_19950);
nor UO_1177 (O_1177,N_19868,N_19967);
or UO_1178 (O_1178,N_19943,N_19851);
or UO_1179 (O_1179,N_19915,N_19945);
nor UO_1180 (O_1180,N_19915,N_19926);
or UO_1181 (O_1181,N_19878,N_19885);
and UO_1182 (O_1182,N_19953,N_19955);
nor UO_1183 (O_1183,N_19938,N_19885);
or UO_1184 (O_1184,N_19915,N_19918);
nand UO_1185 (O_1185,N_19955,N_19938);
and UO_1186 (O_1186,N_19849,N_19892);
xor UO_1187 (O_1187,N_19845,N_19886);
nand UO_1188 (O_1188,N_19871,N_19924);
or UO_1189 (O_1189,N_19931,N_19929);
or UO_1190 (O_1190,N_19891,N_19884);
nor UO_1191 (O_1191,N_19897,N_19904);
or UO_1192 (O_1192,N_19966,N_19935);
or UO_1193 (O_1193,N_19874,N_19853);
and UO_1194 (O_1194,N_19971,N_19873);
xor UO_1195 (O_1195,N_19927,N_19932);
nor UO_1196 (O_1196,N_19993,N_19920);
nand UO_1197 (O_1197,N_19868,N_19989);
nand UO_1198 (O_1198,N_19886,N_19991);
or UO_1199 (O_1199,N_19857,N_19986);
and UO_1200 (O_1200,N_19885,N_19845);
or UO_1201 (O_1201,N_19954,N_19903);
nand UO_1202 (O_1202,N_19941,N_19971);
or UO_1203 (O_1203,N_19901,N_19841);
and UO_1204 (O_1204,N_19840,N_19841);
nand UO_1205 (O_1205,N_19956,N_19968);
or UO_1206 (O_1206,N_19960,N_19968);
xnor UO_1207 (O_1207,N_19990,N_19885);
nor UO_1208 (O_1208,N_19991,N_19899);
nand UO_1209 (O_1209,N_19966,N_19909);
or UO_1210 (O_1210,N_19905,N_19951);
nor UO_1211 (O_1211,N_19932,N_19883);
or UO_1212 (O_1212,N_19956,N_19846);
or UO_1213 (O_1213,N_19928,N_19917);
nand UO_1214 (O_1214,N_19855,N_19842);
or UO_1215 (O_1215,N_19999,N_19981);
nand UO_1216 (O_1216,N_19953,N_19924);
xnor UO_1217 (O_1217,N_19926,N_19845);
and UO_1218 (O_1218,N_19899,N_19910);
or UO_1219 (O_1219,N_19971,N_19894);
nand UO_1220 (O_1220,N_19994,N_19854);
and UO_1221 (O_1221,N_19938,N_19897);
xor UO_1222 (O_1222,N_19854,N_19914);
or UO_1223 (O_1223,N_19941,N_19926);
nor UO_1224 (O_1224,N_19886,N_19857);
and UO_1225 (O_1225,N_19895,N_19943);
and UO_1226 (O_1226,N_19908,N_19990);
or UO_1227 (O_1227,N_19998,N_19962);
nand UO_1228 (O_1228,N_19874,N_19923);
or UO_1229 (O_1229,N_19949,N_19898);
nand UO_1230 (O_1230,N_19925,N_19933);
nor UO_1231 (O_1231,N_19885,N_19881);
or UO_1232 (O_1232,N_19878,N_19842);
and UO_1233 (O_1233,N_19908,N_19961);
or UO_1234 (O_1234,N_19854,N_19912);
or UO_1235 (O_1235,N_19908,N_19904);
and UO_1236 (O_1236,N_19866,N_19930);
and UO_1237 (O_1237,N_19889,N_19938);
or UO_1238 (O_1238,N_19979,N_19971);
or UO_1239 (O_1239,N_19908,N_19924);
or UO_1240 (O_1240,N_19911,N_19954);
nand UO_1241 (O_1241,N_19934,N_19905);
and UO_1242 (O_1242,N_19869,N_19948);
or UO_1243 (O_1243,N_19977,N_19848);
xnor UO_1244 (O_1244,N_19997,N_19880);
and UO_1245 (O_1245,N_19988,N_19883);
or UO_1246 (O_1246,N_19914,N_19978);
nor UO_1247 (O_1247,N_19854,N_19881);
xnor UO_1248 (O_1248,N_19873,N_19907);
nand UO_1249 (O_1249,N_19875,N_19873);
and UO_1250 (O_1250,N_19963,N_19987);
or UO_1251 (O_1251,N_19899,N_19862);
xor UO_1252 (O_1252,N_19871,N_19854);
or UO_1253 (O_1253,N_19923,N_19993);
and UO_1254 (O_1254,N_19959,N_19985);
or UO_1255 (O_1255,N_19944,N_19997);
and UO_1256 (O_1256,N_19939,N_19972);
xnor UO_1257 (O_1257,N_19891,N_19950);
or UO_1258 (O_1258,N_19893,N_19882);
or UO_1259 (O_1259,N_19930,N_19989);
and UO_1260 (O_1260,N_19915,N_19954);
or UO_1261 (O_1261,N_19954,N_19950);
nor UO_1262 (O_1262,N_19982,N_19992);
nand UO_1263 (O_1263,N_19893,N_19889);
nor UO_1264 (O_1264,N_19939,N_19887);
xor UO_1265 (O_1265,N_19992,N_19987);
or UO_1266 (O_1266,N_19939,N_19984);
or UO_1267 (O_1267,N_19942,N_19927);
nor UO_1268 (O_1268,N_19985,N_19911);
xnor UO_1269 (O_1269,N_19846,N_19922);
xnor UO_1270 (O_1270,N_19897,N_19961);
nand UO_1271 (O_1271,N_19932,N_19960);
nand UO_1272 (O_1272,N_19914,N_19955);
nor UO_1273 (O_1273,N_19902,N_19919);
or UO_1274 (O_1274,N_19887,N_19894);
nand UO_1275 (O_1275,N_19969,N_19859);
and UO_1276 (O_1276,N_19939,N_19908);
nand UO_1277 (O_1277,N_19857,N_19853);
or UO_1278 (O_1278,N_19891,N_19880);
or UO_1279 (O_1279,N_19993,N_19879);
xor UO_1280 (O_1280,N_19844,N_19972);
and UO_1281 (O_1281,N_19849,N_19880);
xor UO_1282 (O_1282,N_19960,N_19930);
nand UO_1283 (O_1283,N_19871,N_19978);
nand UO_1284 (O_1284,N_19860,N_19887);
xnor UO_1285 (O_1285,N_19933,N_19842);
xnor UO_1286 (O_1286,N_19879,N_19906);
nor UO_1287 (O_1287,N_19941,N_19923);
or UO_1288 (O_1288,N_19981,N_19870);
nand UO_1289 (O_1289,N_19885,N_19971);
nand UO_1290 (O_1290,N_19904,N_19970);
nor UO_1291 (O_1291,N_19945,N_19948);
xnor UO_1292 (O_1292,N_19912,N_19941);
nor UO_1293 (O_1293,N_19900,N_19862);
nand UO_1294 (O_1294,N_19985,N_19880);
and UO_1295 (O_1295,N_19984,N_19874);
and UO_1296 (O_1296,N_19982,N_19856);
nand UO_1297 (O_1297,N_19921,N_19980);
nand UO_1298 (O_1298,N_19966,N_19843);
xnor UO_1299 (O_1299,N_19881,N_19999);
xor UO_1300 (O_1300,N_19881,N_19864);
and UO_1301 (O_1301,N_19875,N_19937);
and UO_1302 (O_1302,N_19917,N_19905);
nor UO_1303 (O_1303,N_19941,N_19864);
or UO_1304 (O_1304,N_19961,N_19947);
xor UO_1305 (O_1305,N_19901,N_19883);
xor UO_1306 (O_1306,N_19987,N_19977);
xor UO_1307 (O_1307,N_19855,N_19856);
and UO_1308 (O_1308,N_19984,N_19904);
nand UO_1309 (O_1309,N_19896,N_19965);
or UO_1310 (O_1310,N_19993,N_19932);
or UO_1311 (O_1311,N_19849,N_19906);
nor UO_1312 (O_1312,N_19867,N_19864);
nor UO_1313 (O_1313,N_19899,N_19989);
and UO_1314 (O_1314,N_19887,N_19955);
nand UO_1315 (O_1315,N_19922,N_19936);
nand UO_1316 (O_1316,N_19877,N_19888);
nor UO_1317 (O_1317,N_19983,N_19952);
xnor UO_1318 (O_1318,N_19909,N_19938);
xnor UO_1319 (O_1319,N_19849,N_19886);
nand UO_1320 (O_1320,N_19973,N_19948);
or UO_1321 (O_1321,N_19863,N_19913);
or UO_1322 (O_1322,N_19966,N_19928);
or UO_1323 (O_1323,N_19957,N_19894);
nor UO_1324 (O_1324,N_19925,N_19860);
nor UO_1325 (O_1325,N_19979,N_19931);
or UO_1326 (O_1326,N_19933,N_19978);
and UO_1327 (O_1327,N_19850,N_19889);
or UO_1328 (O_1328,N_19861,N_19897);
and UO_1329 (O_1329,N_19878,N_19865);
and UO_1330 (O_1330,N_19913,N_19987);
nand UO_1331 (O_1331,N_19878,N_19857);
xnor UO_1332 (O_1332,N_19949,N_19901);
xnor UO_1333 (O_1333,N_19900,N_19854);
nor UO_1334 (O_1334,N_19980,N_19840);
nor UO_1335 (O_1335,N_19990,N_19974);
or UO_1336 (O_1336,N_19987,N_19849);
and UO_1337 (O_1337,N_19916,N_19940);
nor UO_1338 (O_1338,N_19926,N_19957);
and UO_1339 (O_1339,N_19852,N_19897);
xor UO_1340 (O_1340,N_19915,N_19975);
nand UO_1341 (O_1341,N_19973,N_19840);
nand UO_1342 (O_1342,N_19888,N_19994);
and UO_1343 (O_1343,N_19911,N_19889);
and UO_1344 (O_1344,N_19910,N_19936);
and UO_1345 (O_1345,N_19958,N_19952);
nand UO_1346 (O_1346,N_19907,N_19967);
xnor UO_1347 (O_1347,N_19863,N_19962);
xor UO_1348 (O_1348,N_19877,N_19925);
nand UO_1349 (O_1349,N_19951,N_19984);
nand UO_1350 (O_1350,N_19854,N_19988);
xor UO_1351 (O_1351,N_19963,N_19995);
or UO_1352 (O_1352,N_19941,N_19894);
nand UO_1353 (O_1353,N_19873,N_19964);
nand UO_1354 (O_1354,N_19944,N_19881);
xor UO_1355 (O_1355,N_19895,N_19998);
and UO_1356 (O_1356,N_19997,N_19976);
xnor UO_1357 (O_1357,N_19896,N_19910);
nor UO_1358 (O_1358,N_19990,N_19886);
xor UO_1359 (O_1359,N_19976,N_19991);
nand UO_1360 (O_1360,N_19982,N_19851);
or UO_1361 (O_1361,N_19855,N_19911);
or UO_1362 (O_1362,N_19939,N_19967);
and UO_1363 (O_1363,N_19905,N_19961);
or UO_1364 (O_1364,N_19933,N_19930);
nor UO_1365 (O_1365,N_19862,N_19887);
nand UO_1366 (O_1366,N_19939,N_19916);
nor UO_1367 (O_1367,N_19870,N_19854);
or UO_1368 (O_1368,N_19881,N_19909);
nor UO_1369 (O_1369,N_19955,N_19944);
nand UO_1370 (O_1370,N_19938,N_19928);
xor UO_1371 (O_1371,N_19900,N_19978);
or UO_1372 (O_1372,N_19947,N_19970);
or UO_1373 (O_1373,N_19906,N_19979);
and UO_1374 (O_1374,N_19999,N_19944);
nor UO_1375 (O_1375,N_19844,N_19912);
nor UO_1376 (O_1376,N_19940,N_19870);
xnor UO_1377 (O_1377,N_19942,N_19875);
and UO_1378 (O_1378,N_19878,N_19938);
xnor UO_1379 (O_1379,N_19977,N_19889);
nor UO_1380 (O_1380,N_19911,N_19945);
nor UO_1381 (O_1381,N_19985,N_19964);
nand UO_1382 (O_1382,N_19947,N_19878);
and UO_1383 (O_1383,N_19933,N_19873);
nand UO_1384 (O_1384,N_19941,N_19956);
xnor UO_1385 (O_1385,N_19946,N_19918);
nor UO_1386 (O_1386,N_19958,N_19918);
or UO_1387 (O_1387,N_19872,N_19997);
nand UO_1388 (O_1388,N_19882,N_19986);
nor UO_1389 (O_1389,N_19989,N_19892);
and UO_1390 (O_1390,N_19884,N_19942);
and UO_1391 (O_1391,N_19898,N_19918);
nand UO_1392 (O_1392,N_19848,N_19999);
nor UO_1393 (O_1393,N_19961,N_19987);
nor UO_1394 (O_1394,N_19910,N_19915);
nor UO_1395 (O_1395,N_19901,N_19958);
and UO_1396 (O_1396,N_19920,N_19867);
xnor UO_1397 (O_1397,N_19929,N_19842);
nor UO_1398 (O_1398,N_19989,N_19958);
or UO_1399 (O_1399,N_19998,N_19850);
nand UO_1400 (O_1400,N_19864,N_19962);
and UO_1401 (O_1401,N_19845,N_19962);
or UO_1402 (O_1402,N_19957,N_19952);
nand UO_1403 (O_1403,N_19948,N_19933);
and UO_1404 (O_1404,N_19933,N_19967);
nor UO_1405 (O_1405,N_19872,N_19953);
nor UO_1406 (O_1406,N_19939,N_19849);
nor UO_1407 (O_1407,N_19959,N_19879);
nand UO_1408 (O_1408,N_19940,N_19993);
xor UO_1409 (O_1409,N_19875,N_19868);
or UO_1410 (O_1410,N_19937,N_19919);
xor UO_1411 (O_1411,N_19973,N_19894);
and UO_1412 (O_1412,N_19877,N_19942);
nand UO_1413 (O_1413,N_19945,N_19925);
or UO_1414 (O_1414,N_19921,N_19962);
nand UO_1415 (O_1415,N_19901,N_19879);
and UO_1416 (O_1416,N_19884,N_19996);
and UO_1417 (O_1417,N_19892,N_19929);
nor UO_1418 (O_1418,N_19900,N_19996);
or UO_1419 (O_1419,N_19967,N_19981);
nor UO_1420 (O_1420,N_19859,N_19985);
or UO_1421 (O_1421,N_19849,N_19902);
or UO_1422 (O_1422,N_19881,N_19930);
and UO_1423 (O_1423,N_19920,N_19943);
and UO_1424 (O_1424,N_19845,N_19920);
xnor UO_1425 (O_1425,N_19956,N_19895);
or UO_1426 (O_1426,N_19990,N_19987);
nand UO_1427 (O_1427,N_19933,N_19956);
nand UO_1428 (O_1428,N_19975,N_19949);
and UO_1429 (O_1429,N_19898,N_19914);
and UO_1430 (O_1430,N_19960,N_19869);
xor UO_1431 (O_1431,N_19938,N_19959);
nor UO_1432 (O_1432,N_19923,N_19849);
xnor UO_1433 (O_1433,N_19986,N_19969);
or UO_1434 (O_1434,N_19950,N_19942);
xnor UO_1435 (O_1435,N_19917,N_19950);
and UO_1436 (O_1436,N_19960,N_19904);
xnor UO_1437 (O_1437,N_19864,N_19953);
or UO_1438 (O_1438,N_19932,N_19915);
xnor UO_1439 (O_1439,N_19896,N_19914);
or UO_1440 (O_1440,N_19914,N_19954);
xor UO_1441 (O_1441,N_19844,N_19948);
nor UO_1442 (O_1442,N_19860,N_19906);
or UO_1443 (O_1443,N_19859,N_19850);
or UO_1444 (O_1444,N_19976,N_19856);
nor UO_1445 (O_1445,N_19989,N_19903);
nor UO_1446 (O_1446,N_19906,N_19974);
and UO_1447 (O_1447,N_19898,N_19973);
nand UO_1448 (O_1448,N_19950,N_19851);
nand UO_1449 (O_1449,N_19941,N_19995);
or UO_1450 (O_1450,N_19859,N_19897);
xor UO_1451 (O_1451,N_19991,N_19984);
or UO_1452 (O_1452,N_19956,N_19966);
nand UO_1453 (O_1453,N_19903,N_19909);
or UO_1454 (O_1454,N_19962,N_19933);
nor UO_1455 (O_1455,N_19846,N_19841);
and UO_1456 (O_1456,N_19957,N_19901);
or UO_1457 (O_1457,N_19941,N_19865);
nand UO_1458 (O_1458,N_19965,N_19975);
and UO_1459 (O_1459,N_19994,N_19900);
nand UO_1460 (O_1460,N_19935,N_19994);
nor UO_1461 (O_1461,N_19994,N_19967);
nand UO_1462 (O_1462,N_19995,N_19909);
and UO_1463 (O_1463,N_19943,N_19960);
nor UO_1464 (O_1464,N_19999,N_19909);
nand UO_1465 (O_1465,N_19961,N_19941);
or UO_1466 (O_1466,N_19931,N_19949);
xor UO_1467 (O_1467,N_19860,N_19951);
nand UO_1468 (O_1468,N_19886,N_19953);
xnor UO_1469 (O_1469,N_19856,N_19991);
and UO_1470 (O_1470,N_19842,N_19992);
xor UO_1471 (O_1471,N_19867,N_19939);
and UO_1472 (O_1472,N_19992,N_19898);
nand UO_1473 (O_1473,N_19872,N_19867);
and UO_1474 (O_1474,N_19872,N_19863);
xor UO_1475 (O_1475,N_19976,N_19840);
xnor UO_1476 (O_1476,N_19897,N_19845);
nand UO_1477 (O_1477,N_19935,N_19873);
nand UO_1478 (O_1478,N_19945,N_19995);
nand UO_1479 (O_1479,N_19891,N_19909);
nand UO_1480 (O_1480,N_19894,N_19974);
nand UO_1481 (O_1481,N_19862,N_19896);
nand UO_1482 (O_1482,N_19909,N_19963);
nor UO_1483 (O_1483,N_19999,N_19847);
nor UO_1484 (O_1484,N_19951,N_19925);
nand UO_1485 (O_1485,N_19860,N_19967);
or UO_1486 (O_1486,N_19951,N_19966);
nor UO_1487 (O_1487,N_19992,N_19862);
xnor UO_1488 (O_1488,N_19876,N_19906);
or UO_1489 (O_1489,N_19848,N_19867);
and UO_1490 (O_1490,N_19909,N_19904);
and UO_1491 (O_1491,N_19962,N_19988);
nor UO_1492 (O_1492,N_19937,N_19974);
nor UO_1493 (O_1493,N_19944,N_19852);
or UO_1494 (O_1494,N_19866,N_19906);
nor UO_1495 (O_1495,N_19866,N_19940);
xor UO_1496 (O_1496,N_19847,N_19848);
nor UO_1497 (O_1497,N_19895,N_19978);
nand UO_1498 (O_1498,N_19898,N_19888);
or UO_1499 (O_1499,N_19921,N_19895);
and UO_1500 (O_1500,N_19903,N_19923);
nor UO_1501 (O_1501,N_19865,N_19862);
or UO_1502 (O_1502,N_19947,N_19929);
xnor UO_1503 (O_1503,N_19877,N_19891);
nand UO_1504 (O_1504,N_19933,N_19884);
and UO_1505 (O_1505,N_19928,N_19972);
or UO_1506 (O_1506,N_19920,N_19875);
nand UO_1507 (O_1507,N_19910,N_19878);
nor UO_1508 (O_1508,N_19921,N_19918);
and UO_1509 (O_1509,N_19875,N_19995);
nor UO_1510 (O_1510,N_19956,N_19841);
nand UO_1511 (O_1511,N_19887,N_19843);
nand UO_1512 (O_1512,N_19859,N_19876);
xnor UO_1513 (O_1513,N_19888,N_19901);
and UO_1514 (O_1514,N_19854,N_19856);
and UO_1515 (O_1515,N_19863,N_19939);
xnor UO_1516 (O_1516,N_19925,N_19881);
and UO_1517 (O_1517,N_19999,N_19985);
and UO_1518 (O_1518,N_19971,N_19929);
and UO_1519 (O_1519,N_19948,N_19876);
and UO_1520 (O_1520,N_19941,N_19901);
and UO_1521 (O_1521,N_19862,N_19973);
and UO_1522 (O_1522,N_19994,N_19995);
or UO_1523 (O_1523,N_19972,N_19985);
nor UO_1524 (O_1524,N_19982,N_19899);
nand UO_1525 (O_1525,N_19891,N_19986);
and UO_1526 (O_1526,N_19980,N_19893);
xor UO_1527 (O_1527,N_19884,N_19867);
and UO_1528 (O_1528,N_19858,N_19901);
and UO_1529 (O_1529,N_19847,N_19920);
nor UO_1530 (O_1530,N_19929,N_19981);
nor UO_1531 (O_1531,N_19872,N_19860);
and UO_1532 (O_1532,N_19858,N_19871);
xor UO_1533 (O_1533,N_19908,N_19988);
or UO_1534 (O_1534,N_19840,N_19905);
nand UO_1535 (O_1535,N_19862,N_19860);
nor UO_1536 (O_1536,N_19868,N_19945);
and UO_1537 (O_1537,N_19940,N_19897);
and UO_1538 (O_1538,N_19953,N_19934);
xnor UO_1539 (O_1539,N_19959,N_19945);
xnor UO_1540 (O_1540,N_19927,N_19853);
xor UO_1541 (O_1541,N_19908,N_19985);
or UO_1542 (O_1542,N_19876,N_19840);
or UO_1543 (O_1543,N_19943,N_19853);
nor UO_1544 (O_1544,N_19843,N_19977);
or UO_1545 (O_1545,N_19882,N_19934);
xnor UO_1546 (O_1546,N_19961,N_19967);
and UO_1547 (O_1547,N_19910,N_19869);
xor UO_1548 (O_1548,N_19918,N_19984);
xor UO_1549 (O_1549,N_19976,N_19875);
and UO_1550 (O_1550,N_19889,N_19901);
or UO_1551 (O_1551,N_19912,N_19970);
xor UO_1552 (O_1552,N_19895,N_19850);
xor UO_1553 (O_1553,N_19906,N_19954);
and UO_1554 (O_1554,N_19929,N_19930);
xor UO_1555 (O_1555,N_19880,N_19946);
or UO_1556 (O_1556,N_19975,N_19958);
nand UO_1557 (O_1557,N_19927,N_19862);
and UO_1558 (O_1558,N_19957,N_19881);
and UO_1559 (O_1559,N_19882,N_19877);
nand UO_1560 (O_1560,N_19873,N_19981);
nand UO_1561 (O_1561,N_19844,N_19869);
nor UO_1562 (O_1562,N_19969,N_19954);
and UO_1563 (O_1563,N_19867,N_19871);
xor UO_1564 (O_1564,N_19865,N_19973);
or UO_1565 (O_1565,N_19965,N_19923);
nor UO_1566 (O_1566,N_19897,N_19877);
nand UO_1567 (O_1567,N_19853,N_19928);
nand UO_1568 (O_1568,N_19869,N_19890);
or UO_1569 (O_1569,N_19952,N_19942);
nor UO_1570 (O_1570,N_19925,N_19907);
nand UO_1571 (O_1571,N_19871,N_19999);
nand UO_1572 (O_1572,N_19959,N_19849);
or UO_1573 (O_1573,N_19875,N_19973);
xnor UO_1574 (O_1574,N_19870,N_19916);
or UO_1575 (O_1575,N_19917,N_19865);
and UO_1576 (O_1576,N_19854,N_19978);
nand UO_1577 (O_1577,N_19842,N_19991);
nor UO_1578 (O_1578,N_19885,N_19890);
xor UO_1579 (O_1579,N_19992,N_19937);
or UO_1580 (O_1580,N_19943,N_19858);
xor UO_1581 (O_1581,N_19880,N_19925);
or UO_1582 (O_1582,N_19998,N_19911);
nand UO_1583 (O_1583,N_19963,N_19869);
xnor UO_1584 (O_1584,N_19935,N_19886);
nand UO_1585 (O_1585,N_19873,N_19874);
nor UO_1586 (O_1586,N_19841,N_19980);
nand UO_1587 (O_1587,N_19990,N_19941);
nand UO_1588 (O_1588,N_19875,N_19918);
and UO_1589 (O_1589,N_19905,N_19980);
nand UO_1590 (O_1590,N_19938,N_19944);
and UO_1591 (O_1591,N_19989,N_19861);
or UO_1592 (O_1592,N_19926,N_19888);
xnor UO_1593 (O_1593,N_19987,N_19895);
nor UO_1594 (O_1594,N_19995,N_19964);
xor UO_1595 (O_1595,N_19921,N_19989);
or UO_1596 (O_1596,N_19884,N_19912);
and UO_1597 (O_1597,N_19970,N_19892);
nand UO_1598 (O_1598,N_19970,N_19876);
or UO_1599 (O_1599,N_19985,N_19978);
or UO_1600 (O_1600,N_19988,N_19923);
nor UO_1601 (O_1601,N_19983,N_19901);
or UO_1602 (O_1602,N_19949,N_19902);
xnor UO_1603 (O_1603,N_19919,N_19979);
nand UO_1604 (O_1604,N_19947,N_19908);
xnor UO_1605 (O_1605,N_19951,N_19895);
and UO_1606 (O_1606,N_19947,N_19879);
nor UO_1607 (O_1607,N_19842,N_19874);
nand UO_1608 (O_1608,N_19850,N_19881);
xor UO_1609 (O_1609,N_19979,N_19893);
or UO_1610 (O_1610,N_19860,N_19920);
nand UO_1611 (O_1611,N_19870,N_19956);
and UO_1612 (O_1612,N_19885,N_19904);
nor UO_1613 (O_1613,N_19964,N_19933);
and UO_1614 (O_1614,N_19938,N_19974);
nor UO_1615 (O_1615,N_19855,N_19902);
and UO_1616 (O_1616,N_19902,N_19895);
xnor UO_1617 (O_1617,N_19985,N_19962);
nor UO_1618 (O_1618,N_19867,N_19984);
and UO_1619 (O_1619,N_19901,N_19870);
nand UO_1620 (O_1620,N_19912,N_19872);
xnor UO_1621 (O_1621,N_19896,N_19973);
and UO_1622 (O_1622,N_19957,N_19950);
nand UO_1623 (O_1623,N_19968,N_19998);
nor UO_1624 (O_1624,N_19948,N_19987);
nand UO_1625 (O_1625,N_19960,N_19958);
nand UO_1626 (O_1626,N_19901,N_19872);
or UO_1627 (O_1627,N_19946,N_19968);
or UO_1628 (O_1628,N_19877,N_19917);
nand UO_1629 (O_1629,N_19888,N_19873);
xnor UO_1630 (O_1630,N_19977,N_19881);
xor UO_1631 (O_1631,N_19897,N_19847);
xnor UO_1632 (O_1632,N_19950,N_19889);
nor UO_1633 (O_1633,N_19860,N_19964);
nand UO_1634 (O_1634,N_19906,N_19862);
or UO_1635 (O_1635,N_19982,N_19915);
nand UO_1636 (O_1636,N_19904,N_19850);
or UO_1637 (O_1637,N_19972,N_19891);
and UO_1638 (O_1638,N_19874,N_19871);
nor UO_1639 (O_1639,N_19950,N_19860);
nand UO_1640 (O_1640,N_19842,N_19891);
and UO_1641 (O_1641,N_19988,N_19867);
nand UO_1642 (O_1642,N_19994,N_19843);
nor UO_1643 (O_1643,N_19907,N_19983);
nand UO_1644 (O_1644,N_19928,N_19968);
or UO_1645 (O_1645,N_19847,N_19988);
nand UO_1646 (O_1646,N_19929,N_19843);
nor UO_1647 (O_1647,N_19907,N_19974);
or UO_1648 (O_1648,N_19851,N_19947);
nand UO_1649 (O_1649,N_19970,N_19859);
nor UO_1650 (O_1650,N_19914,N_19888);
nor UO_1651 (O_1651,N_19952,N_19940);
nor UO_1652 (O_1652,N_19897,N_19992);
xor UO_1653 (O_1653,N_19906,N_19920);
nor UO_1654 (O_1654,N_19915,N_19863);
or UO_1655 (O_1655,N_19888,N_19939);
and UO_1656 (O_1656,N_19930,N_19908);
or UO_1657 (O_1657,N_19967,N_19946);
nand UO_1658 (O_1658,N_19916,N_19895);
or UO_1659 (O_1659,N_19953,N_19859);
nor UO_1660 (O_1660,N_19916,N_19875);
nor UO_1661 (O_1661,N_19937,N_19946);
xor UO_1662 (O_1662,N_19958,N_19895);
nand UO_1663 (O_1663,N_19882,N_19905);
or UO_1664 (O_1664,N_19926,N_19953);
nor UO_1665 (O_1665,N_19981,N_19980);
xor UO_1666 (O_1666,N_19944,N_19841);
and UO_1667 (O_1667,N_19841,N_19855);
nor UO_1668 (O_1668,N_19935,N_19896);
nor UO_1669 (O_1669,N_19935,N_19967);
nor UO_1670 (O_1670,N_19936,N_19897);
and UO_1671 (O_1671,N_19886,N_19909);
xnor UO_1672 (O_1672,N_19961,N_19859);
or UO_1673 (O_1673,N_19915,N_19957);
xor UO_1674 (O_1674,N_19890,N_19926);
nand UO_1675 (O_1675,N_19916,N_19936);
nor UO_1676 (O_1676,N_19958,N_19884);
nor UO_1677 (O_1677,N_19991,N_19921);
or UO_1678 (O_1678,N_19937,N_19973);
nor UO_1679 (O_1679,N_19878,N_19846);
nor UO_1680 (O_1680,N_19963,N_19904);
and UO_1681 (O_1681,N_19842,N_19865);
nand UO_1682 (O_1682,N_19925,N_19961);
and UO_1683 (O_1683,N_19907,N_19860);
and UO_1684 (O_1684,N_19857,N_19888);
nor UO_1685 (O_1685,N_19872,N_19879);
and UO_1686 (O_1686,N_19936,N_19928);
and UO_1687 (O_1687,N_19923,N_19869);
nor UO_1688 (O_1688,N_19995,N_19986);
xor UO_1689 (O_1689,N_19997,N_19943);
or UO_1690 (O_1690,N_19884,N_19872);
or UO_1691 (O_1691,N_19973,N_19919);
nor UO_1692 (O_1692,N_19874,N_19976);
nand UO_1693 (O_1693,N_19995,N_19981);
or UO_1694 (O_1694,N_19970,N_19949);
and UO_1695 (O_1695,N_19869,N_19864);
nand UO_1696 (O_1696,N_19960,N_19977);
xor UO_1697 (O_1697,N_19997,N_19957);
nand UO_1698 (O_1698,N_19852,N_19856);
and UO_1699 (O_1699,N_19840,N_19941);
nand UO_1700 (O_1700,N_19905,N_19897);
nand UO_1701 (O_1701,N_19918,N_19962);
or UO_1702 (O_1702,N_19859,N_19935);
nor UO_1703 (O_1703,N_19859,N_19945);
nand UO_1704 (O_1704,N_19859,N_19986);
xor UO_1705 (O_1705,N_19982,N_19907);
or UO_1706 (O_1706,N_19949,N_19960);
nor UO_1707 (O_1707,N_19882,N_19959);
and UO_1708 (O_1708,N_19918,N_19976);
or UO_1709 (O_1709,N_19937,N_19987);
xnor UO_1710 (O_1710,N_19927,N_19857);
nor UO_1711 (O_1711,N_19852,N_19876);
and UO_1712 (O_1712,N_19912,N_19954);
and UO_1713 (O_1713,N_19947,N_19984);
xor UO_1714 (O_1714,N_19946,N_19865);
or UO_1715 (O_1715,N_19961,N_19878);
nand UO_1716 (O_1716,N_19863,N_19940);
nand UO_1717 (O_1717,N_19917,N_19947);
nand UO_1718 (O_1718,N_19996,N_19932);
nand UO_1719 (O_1719,N_19881,N_19905);
and UO_1720 (O_1720,N_19955,N_19921);
nor UO_1721 (O_1721,N_19930,N_19977);
or UO_1722 (O_1722,N_19942,N_19956);
nand UO_1723 (O_1723,N_19845,N_19934);
nand UO_1724 (O_1724,N_19927,N_19990);
nor UO_1725 (O_1725,N_19948,N_19872);
and UO_1726 (O_1726,N_19915,N_19996);
nor UO_1727 (O_1727,N_19998,N_19867);
nand UO_1728 (O_1728,N_19898,N_19856);
nor UO_1729 (O_1729,N_19961,N_19910);
nand UO_1730 (O_1730,N_19992,N_19888);
and UO_1731 (O_1731,N_19993,N_19961);
and UO_1732 (O_1732,N_19891,N_19895);
xnor UO_1733 (O_1733,N_19914,N_19958);
and UO_1734 (O_1734,N_19965,N_19880);
or UO_1735 (O_1735,N_19887,N_19896);
xor UO_1736 (O_1736,N_19972,N_19987);
nand UO_1737 (O_1737,N_19942,N_19984);
nand UO_1738 (O_1738,N_19923,N_19956);
or UO_1739 (O_1739,N_19841,N_19994);
or UO_1740 (O_1740,N_19901,N_19904);
and UO_1741 (O_1741,N_19943,N_19916);
nand UO_1742 (O_1742,N_19987,N_19984);
and UO_1743 (O_1743,N_19973,N_19901);
or UO_1744 (O_1744,N_19880,N_19885);
nand UO_1745 (O_1745,N_19888,N_19959);
nand UO_1746 (O_1746,N_19851,N_19917);
nor UO_1747 (O_1747,N_19991,N_19912);
nand UO_1748 (O_1748,N_19980,N_19844);
or UO_1749 (O_1749,N_19857,N_19942);
and UO_1750 (O_1750,N_19847,N_19865);
nor UO_1751 (O_1751,N_19950,N_19927);
and UO_1752 (O_1752,N_19845,N_19893);
nand UO_1753 (O_1753,N_19960,N_19920);
and UO_1754 (O_1754,N_19845,N_19864);
nor UO_1755 (O_1755,N_19851,N_19938);
or UO_1756 (O_1756,N_19924,N_19937);
nor UO_1757 (O_1757,N_19966,N_19890);
or UO_1758 (O_1758,N_19955,N_19949);
nand UO_1759 (O_1759,N_19923,N_19860);
and UO_1760 (O_1760,N_19937,N_19938);
and UO_1761 (O_1761,N_19984,N_19907);
nand UO_1762 (O_1762,N_19867,N_19885);
or UO_1763 (O_1763,N_19997,N_19954);
nand UO_1764 (O_1764,N_19944,N_19910);
xor UO_1765 (O_1765,N_19957,N_19934);
and UO_1766 (O_1766,N_19878,N_19953);
xnor UO_1767 (O_1767,N_19859,N_19843);
xnor UO_1768 (O_1768,N_19978,N_19920);
xor UO_1769 (O_1769,N_19868,N_19979);
nand UO_1770 (O_1770,N_19935,N_19942);
nor UO_1771 (O_1771,N_19984,N_19854);
nor UO_1772 (O_1772,N_19975,N_19874);
or UO_1773 (O_1773,N_19982,N_19939);
nor UO_1774 (O_1774,N_19901,N_19914);
or UO_1775 (O_1775,N_19938,N_19994);
or UO_1776 (O_1776,N_19979,N_19988);
or UO_1777 (O_1777,N_19974,N_19840);
or UO_1778 (O_1778,N_19964,N_19854);
and UO_1779 (O_1779,N_19873,N_19923);
and UO_1780 (O_1780,N_19980,N_19849);
nand UO_1781 (O_1781,N_19935,N_19888);
nand UO_1782 (O_1782,N_19895,N_19909);
or UO_1783 (O_1783,N_19849,N_19856);
nor UO_1784 (O_1784,N_19918,N_19859);
xor UO_1785 (O_1785,N_19999,N_19994);
and UO_1786 (O_1786,N_19886,N_19938);
xnor UO_1787 (O_1787,N_19988,N_19869);
or UO_1788 (O_1788,N_19849,N_19972);
xor UO_1789 (O_1789,N_19901,N_19859);
nor UO_1790 (O_1790,N_19897,N_19928);
xor UO_1791 (O_1791,N_19968,N_19901);
nor UO_1792 (O_1792,N_19903,N_19845);
nor UO_1793 (O_1793,N_19889,N_19856);
or UO_1794 (O_1794,N_19889,N_19933);
nor UO_1795 (O_1795,N_19900,N_19865);
and UO_1796 (O_1796,N_19849,N_19866);
or UO_1797 (O_1797,N_19874,N_19997);
or UO_1798 (O_1798,N_19993,N_19939);
and UO_1799 (O_1799,N_19961,N_19926);
nor UO_1800 (O_1800,N_19911,N_19922);
and UO_1801 (O_1801,N_19863,N_19947);
nor UO_1802 (O_1802,N_19943,N_19972);
nand UO_1803 (O_1803,N_19879,N_19877);
xnor UO_1804 (O_1804,N_19911,N_19987);
xor UO_1805 (O_1805,N_19967,N_19928);
and UO_1806 (O_1806,N_19847,N_19919);
or UO_1807 (O_1807,N_19915,N_19851);
nand UO_1808 (O_1808,N_19887,N_19846);
and UO_1809 (O_1809,N_19905,N_19928);
nand UO_1810 (O_1810,N_19879,N_19935);
and UO_1811 (O_1811,N_19902,N_19862);
nand UO_1812 (O_1812,N_19997,N_19912);
nand UO_1813 (O_1813,N_19918,N_19848);
and UO_1814 (O_1814,N_19932,N_19916);
and UO_1815 (O_1815,N_19854,N_19950);
nand UO_1816 (O_1816,N_19973,N_19888);
xor UO_1817 (O_1817,N_19907,N_19891);
and UO_1818 (O_1818,N_19950,N_19849);
or UO_1819 (O_1819,N_19993,N_19964);
nand UO_1820 (O_1820,N_19954,N_19888);
or UO_1821 (O_1821,N_19981,N_19947);
or UO_1822 (O_1822,N_19966,N_19858);
nand UO_1823 (O_1823,N_19901,N_19970);
nand UO_1824 (O_1824,N_19929,N_19867);
or UO_1825 (O_1825,N_19984,N_19859);
nand UO_1826 (O_1826,N_19865,N_19912);
nor UO_1827 (O_1827,N_19923,N_19894);
xnor UO_1828 (O_1828,N_19850,N_19880);
or UO_1829 (O_1829,N_19894,N_19907);
and UO_1830 (O_1830,N_19841,N_19909);
or UO_1831 (O_1831,N_19873,N_19961);
and UO_1832 (O_1832,N_19894,N_19959);
or UO_1833 (O_1833,N_19978,N_19859);
or UO_1834 (O_1834,N_19915,N_19907);
nor UO_1835 (O_1835,N_19892,N_19866);
nor UO_1836 (O_1836,N_19904,N_19937);
and UO_1837 (O_1837,N_19853,N_19877);
and UO_1838 (O_1838,N_19900,N_19856);
and UO_1839 (O_1839,N_19921,N_19860);
and UO_1840 (O_1840,N_19843,N_19883);
and UO_1841 (O_1841,N_19873,N_19998);
or UO_1842 (O_1842,N_19931,N_19971);
nor UO_1843 (O_1843,N_19957,N_19890);
and UO_1844 (O_1844,N_19914,N_19840);
or UO_1845 (O_1845,N_19985,N_19906);
and UO_1846 (O_1846,N_19922,N_19904);
xnor UO_1847 (O_1847,N_19909,N_19991);
nand UO_1848 (O_1848,N_19902,N_19963);
nand UO_1849 (O_1849,N_19936,N_19863);
nor UO_1850 (O_1850,N_19888,N_19943);
xor UO_1851 (O_1851,N_19969,N_19881);
nand UO_1852 (O_1852,N_19915,N_19900);
and UO_1853 (O_1853,N_19918,N_19842);
xnor UO_1854 (O_1854,N_19970,N_19980);
nand UO_1855 (O_1855,N_19859,N_19881);
or UO_1856 (O_1856,N_19963,N_19937);
nor UO_1857 (O_1857,N_19919,N_19853);
nand UO_1858 (O_1858,N_19876,N_19959);
xnor UO_1859 (O_1859,N_19860,N_19981);
nor UO_1860 (O_1860,N_19889,N_19865);
and UO_1861 (O_1861,N_19884,N_19913);
or UO_1862 (O_1862,N_19896,N_19861);
or UO_1863 (O_1863,N_19907,N_19861);
xnor UO_1864 (O_1864,N_19953,N_19922);
nand UO_1865 (O_1865,N_19905,N_19874);
nor UO_1866 (O_1866,N_19993,N_19844);
and UO_1867 (O_1867,N_19940,N_19958);
nor UO_1868 (O_1868,N_19905,N_19959);
nor UO_1869 (O_1869,N_19898,N_19913);
and UO_1870 (O_1870,N_19840,N_19956);
or UO_1871 (O_1871,N_19988,N_19971);
and UO_1872 (O_1872,N_19989,N_19964);
nand UO_1873 (O_1873,N_19968,N_19897);
and UO_1874 (O_1874,N_19858,N_19960);
nor UO_1875 (O_1875,N_19925,N_19931);
nand UO_1876 (O_1876,N_19983,N_19947);
and UO_1877 (O_1877,N_19983,N_19859);
and UO_1878 (O_1878,N_19947,N_19914);
nand UO_1879 (O_1879,N_19992,N_19922);
nor UO_1880 (O_1880,N_19849,N_19949);
nor UO_1881 (O_1881,N_19934,N_19912);
xnor UO_1882 (O_1882,N_19896,N_19953);
nor UO_1883 (O_1883,N_19941,N_19885);
xnor UO_1884 (O_1884,N_19951,N_19952);
nor UO_1885 (O_1885,N_19927,N_19914);
xor UO_1886 (O_1886,N_19969,N_19936);
nand UO_1887 (O_1887,N_19877,N_19901);
and UO_1888 (O_1888,N_19867,N_19973);
nand UO_1889 (O_1889,N_19885,N_19887);
or UO_1890 (O_1890,N_19962,N_19964);
nor UO_1891 (O_1891,N_19864,N_19901);
nand UO_1892 (O_1892,N_19941,N_19985);
and UO_1893 (O_1893,N_19964,N_19925);
or UO_1894 (O_1894,N_19977,N_19924);
nor UO_1895 (O_1895,N_19865,N_19974);
or UO_1896 (O_1896,N_19992,N_19963);
or UO_1897 (O_1897,N_19922,N_19883);
xnor UO_1898 (O_1898,N_19864,N_19886);
nand UO_1899 (O_1899,N_19869,N_19953);
nor UO_1900 (O_1900,N_19876,N_19846);
xnor UO_1901 (O_1901,N_19914,N_19885);
and UO_1902 (O_1902,N_19978,N_19882);
nand UO_1903 (O_1903,N_19906,N_19877);
and UO_1904 (O_1904,N_19884,N_19938);
nor UO_1905 (O_1905,N_19988,N_19938);
or UO_1906 (O_1906,N_19966,N_19998);
and UO_1907 (O_1907,N_19975,N_19903);
nor UO_1908 (O_1908,N_19899,N_19992);
or UO_1909 (O_1909,N_19948,N_19970);
xnor UO_1910 (O_1910,N_19956,N_19935);
nor UO_1911 (O_1911,N_19984,N_19988);
xor UO_1912 (O_1912,N_19952,N_19998);
nor UO_1913 (O_1913,N_19849,N_19986);
xnor UO_1914 (O_1914,N_19971,N_19966);
and UO_1915 (O_1915,N_19979,N_19918);
nor UO_1916 (O_1916,N_19944,N_19949);
or UO_1917 (O_1917,N_19940,N_19846);
nor UO_1918 (O_1918,N_19921,N_19896);
nor UO_1919 (O_1919,N_19964,N_19984);
nor UO_1920 (O_1920,N_19852,N_19877);
or UO_1921 (O_1921,N_19954,N_19978);
or UO_1922 (O_1922,N_19913,N_19978);
xor UO_1923 (O_1923,N_19872,N_19940);
or UO_1924 (O_1924,N_19895,N_19845);
and UO_1925 (O_1925,N_19936,N_19955);
or UO_1926 (O_1926,N_19913,N_19960);
nor UO_1927 (O_1927,N_19987,N_19985);
xor UO_1928 (O_1928,N_19984,N_19841);
and UO_1929 (O_1929,N_19908,N_19951);
nand UO_1930 (O_1930,N_19884,N_19881);
or UO_1931 (O_1931,N_19850,N_19841);
or UO_1932 (O_1932,N_19895,N_19870);
xnor UO_1933 (O_1933,N_19899,N_19994);
nor UO_1934 (O_1934,N_19878,N_19932);
and UO_1935 (O_1935,N_19864,N_19922);
or UO_1936 (O_1936,N_19980,N_19923);
and UO_1937 (O_1937,N_19940,N_19973);
xnor UO_1938 (O_1938,N_19905,N_19947);
xor UO_1939 (O_1939,N_19906,N_19895);
or UO_1940 (O_1940,N_19945,N_19974);
or UO_1941 (O_1941,N_19896,N_19872);
and UO_1942 (O_1942,N_19900,N_19923);
and UO_1943 (O_1943,N_19868,N_19966);
or UO_1944 (O_1944,N_19870,N_19944);
xor UO_1945 (O_1945,N_19970,N_19921);
nor UO_1946 (O_1946,N_19937,N_19922);
xnor UO_1947 (O_1947,N_19962,N_19916);
and UO_1948 (O_1948,N_19924,N_19967);
and UO_1949 (O_1949,N_19980,N_19955);
nor UO_1950 (O_1950,N_19884,N_19914);
nor UO_1951 (O_1951,N_19994,N_19908);
nor UO_1952 (O_1952,N_19923,N_19872);
xnor UO_1953 (O_1953,N_19938,N_19867);
and UO_1954 (O_1954,N_19911,N_19980);
nand UO_1955 (O_1955,N_19900,N_19937);
and UO_1956 (O_1956,N_19884,N_19918);
xnor UO_1957 (O_1957,N_19899,N_19988);
or UO_1958 (O_1958,N_19910,N_19916);
or UO_1959 (O_1959,N_19922,N_19844);
xnor UO_1960 (O_1960,N_19950,N_19902);
and UO_1961 (O_1961,N_19950,N_19862);
nand UO_1962 (O_1962,N_19962,N_19935);
xnor UO_1963 (O_1963,N_19863,N_19876);
or UO_1964 (O_1964,N_19870,N_19942);
nand UO_1965 (O_1965,N_19925,N_19955);
nor UO_1966 (O_1966,N_19847,N_19842);
or UO_1967 (O_1967,N_19929,N_19922);
xnor UO_1968 (O_1968,N_19906,N_19951);
nand UO_1969 (O_1969,N_19951,N_19877);
nand UO_1970 (O_1970,N_19891,N_19936);
nand UO_1971 (O_1971,N_19847,N_19883);
or UO_1972 (O_1972,N_19899,N_19973);
nand UO_1973 (O_1973,N_19842,N_19974);
xor UO_1974 (O_1974,N_19912,N_19927);
nor UO_1975 (O_1975,N_19993,N_19901);
nand UO_1976 (O_1976,N_19901,N_19944);
or UO_1977 (O_1977,N_19905,N_19964);
xnor UO_1978 (O_1978,N_19923,N_19892);
nor UO_1979 (O_1979,N_19882,N_19927);
xnor UO_1980 (O_1980,N_19910,N_19893);
nor UO_1981 (O_1981,N_19983,N_19925);
and UO_1982 (O_1982,N_19998,N_19874);
xnor UO_1983 (O_1983,N_19958,N_19976);
or UO_1984 (O_1984,N_19952,N_19955);
nand UO_1985 (O_1985,N_19992,N_19978);
and UO_1986 (O_1986,N_19989,N_19914);
xnor UO_1987 (O_1987,N_19992,N_19847);
or UO_1988 (O_1988,N_19859,N_19900);
nand UO_1989 (O_1989,N_19914,N_19936);
nor UO_1990 (O_1990,N_19936,N_19853);
nor UO_1991 (O_1991,N_19869,N_19900);
or UO_1992 (O_1992,N_19924,N_19861);
nor UO_1993 (O_1993,N_19998,N_19944);
nor UO_1994 (O_1994,N_19930,N_19982);
nor UO_1995 (O_1995,N_19980,N_19937);
nor UO_1996 (O_1996,N_19949,N_19978);
nor UO_1997 (O_1997,N_19935,N_19950);
nand UO_1998 (O_1998,N_19990,N_19932);
and UO_1999 (O_1999,N_19963,N_19890);
xor UO_2000 (O_2000,N_19949,N_19946);
or UO_2001 (O_2001,N_19997,N_19867);
or UO_2002 (O_2002,N_19896,N_19869);
nor UO_2003 (O_2003,N_19974,N_19991);
nand UO_2004 (O_2004,N_19894,N_19975);
nand UO_2005 (O_2005,N_19877,N_19995);
xnor UO_2006 (O_2006,N_19994,N_19863);
nand UO_2007 (O_2007,N_19988,N_19972);
xor UO_2008 (O_2008,N_19862,N_19967);
nor UO_2009 (O_2009,N_19923,N_19918);
nand UO_2010 (O_2010,N_19888,N_19934);
nor UO_2011 (O_2011,N_19897,N_19882);
xnor UO_2012 (O_2012,N_19881,N_19903);
nand UO_2013 (O_2013,N_19971,N_19868);
or UO_2014 (O_2014,N_19925,N_19953);
xnor UO_2015 (O_2015,N_19984,N_19941);
and UO_2016 (O_2016,N_19973,N_19932);
or UO_2017 (O_2017,N_19929,N_19943);
nand UO_2018 (O_2018,N_19955,N_19948);
and UO_2019 (O_2019,N_19857,N_19909);
nand UO_2020 (O_2020,N_19888,N_19854);
xnor UO_2021 (O_2021,N_19854,N_19896);
and UO_2022 (O_2022,N_19986,N_19943);
or UO_2023 (O_2023,N_19874,N_19936);
nor UO_2024 (O_2024,N_19850,N_19840);
nor UO_2025 (O_2025,N_19908,N_19960);
nor UO_2026 (O_2026,N_19878,N_19888);
and UO_2027 (O_2027,N_19915,N_19860);
nand UO_2028 (O_2028,N_19850,N_19966);
or UO_2029 (O_2029,N_19863,N_19997);
nor UO_2030 (O_2030,N_19936,N_19903);
nor UO_2031 (O_2031,N_19950,N_19988);
and UO_2032 (O_2032,N_19931,N_19870);
or UO_2033 (O_2033,N_19990,N_19895);
or UO_2034 (O_2034,N_19966,N_19978);
or UO_2035 (O_2035,N_19840,N_19891);
nor UO_2036 (O_2036,N_19969,N_19925);
and UO_2037 (O_2037,N_19845,N_19960);
xnor UO_2038 (O_2038,N_19934,N_19858);
nand UO_2039 (O_2039,N_19899,N_19950);
and UO_2040 (O_2040,N_19896,N_19985);
xnor UO_2041 (O_2041,N_19944,N_19898);
nand UO_2042 (O_2042,N_19879,N_19905);
xor UO_2043 (O_2043,N_19927,N_19936);
xor UO_2044 (O_2044,N_19974,N_19999);
and UO_2045 (O_2045,N_19844,N_19849);
xnor UO_2046 (O_2046,N_19984,N_19932);
xor UO_2047 (O_2047,N_19858,N_19951);
nand UO_2048 (O_2048,N_19951,N_19880);
xor UO_2049 (O_2049,N_19956,N_19849);
or UO_2050 (O_2050,N_19882,N_19939);
xnor UO_2051 (O_2051,N_19880,N_19895);
and UO_2052 (O_2052,N_19942,N_19864);
or UO_2053 (O_2053,N_19962,N_19906);
or UO_2054 (O_2054,N_19990,N_19922);
and UO_2055 (O_2055,N_19941,N_19883);
nor UO_2056 (O_2056,N_19973,N_19917);
and UO_2057 (O_2057,N_19994,N_19911);
nor UO_2058 (O_2058,N_19976,N_19844);
or UO_2059 (O_2059,N_19916,N_19907);
or UO_2060 (O_2060,N_19871,N_19901);
or UO_2061 (O_2061,N_19937,N_19868);
nor UO_2062 (O_2062,N_19857,N_19996);
nor UO_2063 (O_2063,N_19876,N_19993);
and UO_2064 (O_2064,N_19853,N_19844);
xnor UO_2065 (O_2065,N_19972,N_19956);
and UO_2066 (O_2066,N_19992,N_19980);
xnor UO_2067 (O_2067,N_19852,N_19929);
xnor UO_2068 (O_2068,N_19967,N_19885);
or UO_2069 (O_2069,N_19897,N_19910);
nand UO_2070 (O_2070,N_19999,N_19968);
nor UO_2071 (O_2071,N_19905,N_19903);
nor UO_2072 (O_2072,N_19979,N_19857);
xor UO_2073 (O_2073,N_19931,N_19958);
xor UO_2074 (O_2074,N_19996,N_19852);
xnor UO_2075 (O_2075,N_19910,N_19951);
and UO_2076 (O_2076,N_19916,N_19935);
nand UO_2077 (O_2077,N_19862,N_19911);
and UO_2078 (O_2078,N_19864,N_19851);
nor UO_2079 (O_2079,N_19970,N_19920);
and UO_2080 (O_2080,N_19856,N_19893);
xor UO_2081 (O_2081,N_19841,N_19847);
and UO_2082 (O_2082,N_19864,N_19852);
or UO_2083 (O_2083,N_19900,N_19946);
and UO_2084 (O_2084,N_19998,N_19875);
and UO_2085 (O_2085,N_19851,N_19974);
nor UO_2086 (O_2086,N_19907,N_19853);
or UO_2087 (O_2087,N_19984,N_19888);
and UO_2088 (O_2088,N_19855,N_19859);
xnor UO_2089 (O_2089,N_19915,N_19891);
or UO_2090 (O_2090,N_19993,N_19955);
nand UO_2091 (O_2091,N_19868,N_19969);
xor UO_2092 (O_2092,N_19953,N_19998);
xnor UO_2093 (O_2093,N_19949,N_19942);
and UO_2094 (O_2094,N_19863,N_19973);
or UO_2095 (O_2095,N_19958,N_19921);
nand UO_2096 (O_2096,N_19916,N_19917);
nand UO_2097 (O_2097,N_19906,N_19965);
or UO_2098 (O_2098,N_19902,N_19842);
nor UO_2099 (O_2099,N_19959,N_19913);
nor UO_2100 (O_2100,N_19841,N_19919);
nand UO_2101 (O_2101,N_19925,N_19926);
xor UO_2102 (O_2102,N_19842,N_19928);
or UO_2103 (O_2103,N_19881,N_19939);
nand UO_2104 (O_2104,N_19943,N_19873);
nor UO_2105 (O_2105,N_19914,N_19930);
and UO_2106 (O_2106,N_19981,N_19902);
and UO_2107 (O_2107,N_19990,N_19964);
and UO_2108 (O_2108,N_19848,N_19965);
or UO_2109 (O_2109,N_19854,N_19928);
nand UO_2110 (O_2110,N_19960,N_19945);
nand UO_2111 (O_2111,N_19841,N_19897);
and UO_2112 (O_2112,N_19930,N_19941);
nor UO_2113 (O_2113,N_19995,N_19947);
and UO_2114 (O_2114,N_19915,N_19935);
or UO_2115 (O_2115,N_19929,N_19923);
xnor UO_2116 (O_2116,N_19896,N_19956);
nand UO_2117 (O_2117,N_19977,N_19992);
or UO_2118 (O_2118,N_19880,N_19974);
xor UO_2119 (O_2119,N_19924,N_19935);
nand UO_2120 (O_2120,N_19930,N_19983);
and UO_2121 (O_2121,N_19864,N_19939);
and UO_2122 (O_2122,N_19913,N_19856);
xnor UO_2123 (O_2123,N_19938,N_19919);
and UO_2124 (O_2124,N_19911,N_19931);
nor UO_2125 (O_2125,N_19922,N_19919);
or UO_2126 (O_2126,N_19852,N_19949);
xor UO_2127 (O_2127,N_19975,N_19844);
xor UO_2128 (O_2128,N_19855,N_19881);
or UO_2129 (O_2129,N_19845,N_19991);
xor UO_2130 (O_2130,N_19843,N_19959);
xnor UO_2131 (O_2131,N_19876,N_19843);
xor UO_2132 (O_2132,N_19934,N_19897);
nand UO_2133 (O_2133,N_19885,N_19859);
nand UO_2134 (O_2134,N_19913,N_19852);
nand UO_2135 (O_2135,N_19886,N_19889);
nand UO_2136 (O_2136,N_19898,N_19984);
nor UO_2137 (O_2137,N_19892,N_19931);
or UO_2138 (O_2138,N_19955,N_19851);
nand UO_2139 (O_2139,N_19871,N_19976);
nand UO_2140 (O_2140,N_19967,N_19896);
xor UO_2141 (O_2141,N_19859,N_19975);
xnor UO_2142 (O_2142,N_19929,N_19968);
xnor UO_2143 (O_2143,N_19932,N_19868);
and UO_2144 (O_2144,N_19860,N_19855);
xor UO_2145 (O_2145,N_19868,N_19981);
xnor UO_2146 (O_2146,N_19871,N_19911);
and UO_2147 (O_2147,N_19864,N_19968);
xor UO_2148 (O_2148,N_19926,N_19997);
nor UO_2149 (O_2149,N_19842,N_19873);
or UO_2150 (O_2150,N_19910,N_19873);
nand UO_2151 (O_2151,N_19989,N_19940);
and UO_2152 (O_2152,N_19917,N_19924);
nor UO_2153 (O_2153,N_19916,N_19944);
or UO_2154 (O_2154,N_19863,N_19864);
and UO_2155 (O_2155,N_19876,N_19880);
xnor UO_2156 (O_2156,N_19880,N_19867);
or UO_2157 (O_2157,N_19902,N_19930);
nor UO_2158 (O_2158,N_19855,N_19965);
or UO_2159 (O_2159,N_19962,N_19940);
xor UO_2160 (O_2160,N_19876,N_19997);
nand UO_2161 (O_2161,N_19926,N_19964);
nand UO_2162 (O_2162,N_19909,N_19927);
xnor UO_2163 (O_2163,N_19944,N_19890);
and UO_2164 (O_2164,N_19944,N_19859);
xor UO_2165 (O_2165,N_19889,N_19984);
nand UO_2166 (O_2166,N_19907,N_19945);
nand UO_2167 (O_2167,N_19952,N_19873);
nor UO_2168 (O_2168,N_19958,N_19988);
or UO_2169 (O_2169,N_19950,N_19998);
or UO_2170 (O_2170,N_19879,N_19960);
and UO_2171 (O_2171,N_19864,N_19877);
or UO_2172 (O_2172,N_19963,N_19988);
and UO_2173 (O_2173,N_19936,N_19935);
nor UO_2174 (O_2174,N_19847,N_19941);
nor UO_2175 (O_2175,N_19911,N_19842);
or UO_2176 (O_2176,N_19963,N_19882);
and UO_2177 (O_2177,N_19933,N_19923);
or UO_2178 (O_2178,N_19997,N_19852);
xor UO_2179 (O_2179,N_19913,N_19934);
and UO_2180 (O_2180,N_19880,N_19910);
or UO_2181 (O_2181,N_19922,N_19872);
or UO_2182 (O_2182,N_19958,N_19969);
nand UO_2183 (O_2183,N_19957,N_19865);
or UO_2184 (O_2184,N_19923,N_19954);
nor UO_2185 (O_2185,N_19945,N_19964);
xor UO_2186 (O_2186,N_19907,N_19843);
nand UO_2187 (O_2187,N_19936,N_19923);
nand UO_2188 (O_2188,N_19932,N_19991);
nor UO_2189 (O_2189,N_19954,N_19861);
nor UO_2190 (O_2190,N_19876,N_19917);
or UO_2191 (O_2191,N_19841,N_19937);
nand UO_2192 (O_2192,N_19966,N_19923);
nand UO_2193 (O_2193,N_19860,N_19896);
nor UO_2194 (O_2194,N_19961,N_19923);
or UO_2195 (O_2195,N_19869,N_19973);
xnor UO_2196 (O_2196,N_19937,N_19913);
or UO_2197 (O_2197,N_19988,N_19841);
and UO_2198 (O_2198,N_19930,N_19899);
nand UO_2199 (O_2199,N_19857,N_19972);
xor UO_2200 (O_2200,N_19912,N_19876);
nor UO_2201 (O_2201,N_19900,N_19976);
nor UO_2202 (O_2202,N_19975,N_19962);
nand UO_2203 (O_2203,N_19964,N_19982);
and UO_2204 (O_2204,N_19984,N_19883);
or UO_2205 (O_2205,N_19932,N_19865);
and UO_2206 (O_2206,N_19995,N_19955);
nand UO_2207 (O_2207,N_19997,N_19878);
xor UO_2208 (O_2208,N_19916,N_19993);
or UO_2209 (O_2209,N_19999,N_19844);
nand UO_2210 (O_2210,N_19946,N_19894);
nor UO_2211 (O_2211,N_19871,N_19860);
nor UO_2212 (O_2212,N_19967,N_19947);
nand UO_2213 (O_2213,N_19989,N_19885);
nor UO_2214 (O_2214,N_19881,N_19956);
xor UO_2215 (O_2215,N_19946,N_19982);
and UO_2216 (O_2216,N_19952,N_19860);
or UO_2217 (O_2217,N_19904,N_19981);
nand UO_2218 (O_2218,N_19869,N_19893);
nor UO_2219 (O_2219,N_19934,N_19940);
or UO_2220 (O_2220,N_19840,N_19885);
and UO_2221 (O_2221,N_19884,N_19848);
xnor UO_2222 (O_2222,N_19970,N_19973);
and UO_2223 (O_2223,N_19980,N_19968);
or UO_2224 (O_2224,N_19955,N_19999);
and UO_2225 (O_2225,N_19988,N_19955);
nor UO_2226 (O_2226,N_19920,N_19983);
nand UO_2227 (O_2227,N_19974,N_19844);
or UO_2228 (O_2228,N_19970,N_19965);
nand UO_2229 (O_2229,N_19855,N_19984);
xnor UO_2230 (O_2230,N_19999,N_19923);
and UO_2231 (O_2231,N_19912,N_19979);
and UO_2232 (O_2232,N_19961,N_19921);
xnor UO_2233 (O_2233,N_19931,N_19915);
and UO_2234 (O_2234,N_19907,N_19941);
xnor UO_2235 (O_2235,N_19980,N_19906);
xnor UO_2236 (O_2236,N_19899,N_19943);
xor UO_2237 (O_2237,N_19948,N_19994);
and UO_2238 (O_2238,N_19958,N_19967);
nand UO_2239 (O_2239,N_19959,N_19956);
xnor UO_2240 (O_2240,N_19925,N_19915);
or UO_2241 (O_2241,N_19882,N_19999);
or UO_2242 (O_2242,N_19920,N_19913);
or UO_2243 (O_2243,N_19896,N_19865);
xnor UO_2244 (O_2244,N_19929,N_19864);
nand UO_2245 (O_2245,N_19973,N_19876);
or UO_2246 (O_2246,N_19855,N_19901);
or UO_2247 (O_2247,N_19898,N_19974);
or UO_2248 (O_2248,N_19840,N_19883);
nand UO_2249 (O_2249,N_19960,N_19866);
xnor UO_2250 (O_2250,N_19941,N_19963);
xnor UO_2251 (O_2251,N_19976,N_19885);
xnor UO_2252 (O_2252,N_19972,N_19864);
or UO_2253 (O_2253,N_19936,N_19906);
and UO_2254 (O_2254,N_19856,N_19970);
or UO_2255 (O_2255,N_19881,N_19975);
xnor UO_2256 (O_2256,N_19927,N_19982);
nor UO_2257 (O_2257,N_19909,N_19855);
nor UO_2258 (O_2258,N_19877,N_19883);
and UO_2259 (O_2259,N_19960,N_19963);
xor UO_2260 (O_2260,N_19885,N_19919);
xnor UO_2261 (O_2261,N_19882,N_19874);
nand UO_2262 (O_2262,N_19849,N_19879);
xnor UO_2263 (O_2263,N_19871,N_19997);
or UO_2264 (O_2264,N_19907,N_19956);
nand UO_2265 (O_2265,N_19981,N_19964);
or UO_2266 (O_2266,N_19939,N_19971);
nand UO_2267 (O_2267,N_19988,N_19997);
and UO_2268 (O_2268,N_19913,N_19905);
nor UO_2269 (O_2269,N_19911,N_19857);
nand UO_2270 (O_2270,N_19921,N_19856);
or UO_2271 (O_2271,N_19959,N_19877);
or UO_2272 (O_2272,N_19860,N_19982);
or UO_2273 (O_2273,N_19891,N_19991);
nor UO_2274 (O_2274,N_19865,N_19850);
and UO_2275 (O_2275,N_19964,N_19886);
nor UO_2276 (O_2276,N_19866,N_19916);
nor UO_2277 (O_2277,N_19969,N_19875);
xor UO_2278 (O_2278,N_19882,N_19870);
nor UO_2279 (O_2279,N_19885,N_19842);
xnor UO_2280 (O_2280,N_19948,N_19885);
nand UO_2281 (O_2281,N_19926,N_19846);
nor UO_2282 (O_2282,N_19950,N_19880);
xor UO_2283 (O_2283,N_19943,N_19938);
nor UO_2284 (O_2284,N_19949,N_19950);
or UO_2285 (O_2285,N_19925,N_19922);
or UO_2286 (O_2286,N_19980,N_19852);
and UO_2287 (O_2287,N_19876,N_19971);
and UO_2288 (O_2288,N_19913,N_19850);
nand UO_2289 (O_2289,N_19997,N_19953);
or UO_2290 (O_2290,N_19974,N_19870);
nor UO_2291 (O_2291,N_19896,N_19871);
xor UO_2292 (O_2292,N_19905,N_19997);
xor UO_2293 (O_2293,N_19966,N_19889);
and UO_2294 (O_2294,N_19972,N_19989);
or UO_2295 (O_2295,N_19870,N_19898);
nand UO_2296 (O_2296,N_19899,N_19932);
xor UO_2297 (O_2297,N_19908,N_19915);
or UO_2298 (O_2298,N_19953,N_19951);
nor UO_2299 (O_2299,N_19928,N_19912);
or UO_2300 (O_2300,N_19947,N_19862);
xnor UO_2301 (O_2301,N_19948,N_19853);
xor UO_2302 (O_2302,N_19942,N_19946);
and UO_2303 (O_2303,N_19876,N_19923);
and UO_2304 (O_2304,N_19872,N_19944);
nor UO_2305 (O_2305,N_19914,N_19977);
nand UO_2306 (O_2306,N_19982,N_19994);
or UO_2307 (O_2307,N_19967,N_19934);
or UO_2308 (O_2308,N_19931,N_19867);
and UO_2309 (O_2309,N_19903,N_19852);
nor UO_2310 (O_2310,N_19929,N_19885);
and UO_2311 (O_2311,N_19881,N_19950);
or UO_2312 (O_2312,N_19932,N_19905);
nand UO_2313 (O_2313,N_19863,N_19884);
or UO_2314 (O_2314,N_19996,N_19877);
or UO_2315 (O_2315,N_19903,N_19842);
or UO_2316 (O_2316,N_19996,N_19868);
and UO_2317 (O_2317,N_19844,N_19927);
and UO_2318 (O_2318,N_19912,N_19975);
or UO_2319 (O_2319,N_19970,N_19886);
xor UO_2320 (O_2320,N_19879,N_19873);
or UO_2321 (O_2321,N_19938,N_19902);
or UO_2322 (O_2322,N_19970,N_19905);
xnor UO_2323 (O_2323,N_19841,N_19842);
or UO_2324 (O_2324,N_19961,N_19952);
nand UO_2325 (O_2325,N_19842,N_19887);
or UO_2326 (O_2326,N_19908,N_19882);
nor UO_2327 (O_2327,N_19880,N_19898);
xnor UO_2328 (O_2328,N_19909,N_19958);
xor UO_2329 (O_2329,N_19872,N_19942);
or UO_2330 (O_2330,N_19917,N_19854);
or UO_2331 (O_2331,N_19922,N_19920);
and UO_2332 (O_2332,N_19886,N_19963);
nor UO_2333 (O_2333,N_19901,N_19906);
xnor UO_2334 (O_2334,N_19992,N_19948);
nand UO_2335 (O_2335,N_19965,N_19894);
nand UO_2336 (O_2336,N_19985,N_19897);
or UO_2337 (O_2337,N_19921,N_19893);
nor UO_2338 (O_2338,N_19939,N_19844);
xnor UO_2339 (O_2339,N_19980,N_19963);
and UO_2340 (O_2340,N_19944,N_19958);
or UO_2341 (O_2341,N_19956,N_19983);
nand UO_2342 (O_2342,N_19906,N_19932);
nand UO_2343 (O_2343,N_19971,N_19861);
and UO_2344 (O_2344,N_19892,N_19945);
or UO_2345 (O_2345,N_19983,N_19985);
and UO_2346 (O_2346,N_19965,N_19977);
or UO_2347 (O_2347,N_19855,N_19950);
nand UO_2348 (O_2348,N_19962,N_19923);
and UO_2349 (O_2349,N_19896,N_19852);
nor UO_2350 (O_2350,N_19909,N_19952);
and UO_2351 (O_2351,N_19948,N_19901);
or UO_2352 (O_2352,N_19882,N_19876);
nor UO_2353 (O_2353,N_19967,N_19880);
xor UO_2354 (O_2354,N_19844,N_19996);
nor UO_2355 (O_2355,N_19850,N_19846);
and UO_2356 (O_2356,N_19949,N_19850);
or UO_2357 (O_2357,N_19953,N_19898);
nor UO_2358 (O_2358,N_19929,N_19934);
nor UO_2359 (O_2359,N_19973,N_19878);
or UO_2360 (O_2360,N_19992,N_19882);
or UO_2361 (O_2361,N_19858,N_19950);
nor UO_2362 (O_2362,N_19923,N_19912);
xor UO_2363 (O_2363,N_19969,N_19884);
nor UO_2364 (O_2364,N_19871,N_19865);
or UO_2365 (O_2365,N_19871,N_19920);
nor UO_2366 (O_2366,N_19852,N_19995);
nor UO_2367 (O_2367,N_19941,N_19862);
xor UO_2368 (O_2368,N_19900,N_19945);
nand UO_2369 (O_2369,N_19887,N_19983);
xor UO_2370 (O_2370,N_19944,N_19906);
xnor UO_2371 (O_2371,N_19932,N_19858);
and UO_2372 (O_2372,N_19944,N_19873);
nand UO_2373 (O_2373,N_19843,N_19912);
or UO_2374 (O_2374,N_19904,N_19944);
xnor UO_2375 (O_2375,N_19941,N_19931);
or UO_2376 (O_2376,N_19876,N_19983);
nor UO_2377 (O_2377,N_19982,N_19971);
xnor UO_2378 (O_2378,N_19858,N_19864);
and UO_2379 (O_2379,N_19919,N_19895);
and UO_2380 (O_2380,N_19890,N_19872);
or UO_2381 (O_2381,N_19874,N_19875);
nor UO_2382 (O_2382,N_19917,N_19946);
xor UO_2383 (O_2383,N_19849,N_19948);
or UO_2384 (O_2384,N_19894,N_19926);
nor UO_2385 (O_2385,N_19847,N_19845);
nor UO_2386 (O_2386,N_19902,N_19869);
or UO_2387 (O_2387,N_19969,N_19989);
xnor UO_2388 (O_2388,N_19884,N_19897);
nor UO_2389 (O_2389,N_19917,N_19883);
nand UO_2390 (O_2390,N_19922,N_19909);
nor UO_2391 (O_2391,N_19979,N_19884);
nor UO_2392 (O_2392,N_19902,N_19892);
nand UO_2393 (O_2393,N_19946,N_19877);
xor UO_2394 (O_2394,N_19942,N_19986);
or UO_2395 (O_2395,N_19849,N_19918);
or UO_2396 (O_2396,N_19987,N_19941);
xor UO_2397 (O_2397,N_19903,N_19879);
xnor UO_2398 (O_2398,N_19995,N_19969);
xnor UO_2399 (O_2399,N_19986,N_19967);
xor UO_2400 (O_2400,N_19974,N_19901);
or UO_2401 (O_2401,N_19843,N_19844);
nand UO_2402 (O_2402,N_19886,N_19951);
or UO_2403 (O_2403,N_19969,N_19896);
xor UO_2404 (O_2404,N_19933,N_19912);
and UO_2405 (O_2405,N_19843,N_19943);
xnor UO_2406 (O_2406,N_19977,N_19866);
or UO_2407 (O_2407,N_19991,N_19854);
and UO_2408 (O_2408,N_19956,N_19960);
or UO_2409 (O_2409,N_19986,N_19941);
nand UO_2410 (O_2410,N_19963,N_19977);
and UO_2411 (O_2411,N_19970,N_19855);
nor UO_2412 (O_2412,N_19894,N_19922);
xor UO_2413 (O_2413,N_19874,N_19935);
or UO_2414 (O_2414,N_19927,N_19920);
and UO_2415 (O_2415,N_19981,N_19890);
nor UO_2416 (O_2416,N_19917,N_19978);
xnor UO_2417 (O_2417,N_19894,N_19992);
and UO_2418 (O_2418,N_19878,N_19943);
nor UO_2419 (O_2419,N_19907,N_19879);
and UO_2420 (O_2420,N_19852,N_19869);
nor UO_2421 (O_2421,N_19868,N_19873);
nor UO_2422 (O_2422,N_19843,N_19939);
nor UO_2423 (O_2423,N_19922,N_19863);
nand UO_2424 (O_2424,N_19965,N_19875);
and UO_2425 (O_2425,N_19908,N_19995);
xnor UO_2426 (O_2426,N_19927,N_19894);
nor UO_2427 (O_2427,N_19887,N_19933);
nand UO_2428 (O_2428,N_19864,N_19955);
and UO_2429 (O_2429,N_19964,N_19852);
nor UO_2430 (O_2430,N_19847,N_19892);
or UO_2431 (O_2431,N_19914,N_19950);
xor UO_2432 (O_2432,N_19884,N_19850);
and UO_2433 (O_2433,N_19917,N_19889);
xor UO_2434 (O_2434,N_19860,N_19882);
nor UO_2435 (O_2435,N_19870,N_19976);
nor UO_2436 (O_2436,N_19842,N_19938);
nor UO_2437 (O_2437,N_19903,N_19904);
or UO_2438 (O_2438,N_19945,N_19968);
or UO_2439 (O_2439,N_19870,N_19864);
and UO_2440 (O_2440,N_19961,N_19999);
and UO_2441 (O_2441,N_19999,N_19842);
nand UO_2442 (O_2442,N_19993,N_19960);
or UO_2443 (O_2443,N_19871,N_19928);
nor UO_2444 (O_2444,N_19840,N_19917);
or UO_2445 (O_2445,N_19941,N_19876);
nor UO_2446 (O_2446,N_19893,N_19984);
or UO_2447 (O_2447,N_19888,N_19924);
nor UO_2448 (O_2448,N_19919,N_19858);
and UO_2449 (O_2449,N_19929,N_19883);
xor UO_2450 (O_2450,N_19983,N_19906);
and UO_2451 (O_2451,N_19975,N_19942);
nand UO_2452 (O_2452,N_19930,N_19963);
xor UO_2453 (O_2453,N_19916,N_19925);
or UO_2454 (O_2454,N_19937,N_19915);
or UO_2455 (O_2455,N_19983,N_19911);
or UO_2456 (O_2456,N_19997,N_19933);
nor UO_2457 (O_2457,N_19848,N_19843);
xnor UO_2458 (O_2458,N_19904,N_19919);
or UO_2459 (O_2459,N_19944,N_19846);
nor UO_2460 (O_2460,N_19927,N_19917);
and UO_2461 (O_2461,N_19995,N_19977);
nor UO_2462 (O_2462,N_19990,N_19851);
xor UO_2463 (O_2463,N_19880,N_19883);
xor UO_2464 (O_2464,N_19902,N_19972);
nor UO_2465 (O_2465,N_19974,N_19900);
and UO_2466 (O_2466,N_19918,N_19978);
and UO_2467 (O_2467,N_19985,N_19887);
nand UO_2468 (O_2468,N_19969,N_19879);
nand UO_2469 (O_2469,N_19967,N_19863);
or UO_2470 (O_2470,N_19952,N_19933);
and UO_2471 (O_2471,N_19984,N_19915);
nand UO_2472 (O_2472,N_19867,N_19924);
or UO_2473 (O_2473,N_19883,N_19890);
xnor UO_2474 (O_2474,N_19867,N_19855);
and UO_2475 (O_2475,N_19920,N_19865);
or UO_2476 (O_2476,N_19988,N_19907);
xnor UO_2477 (O_2477,N_19965,N_19898);
and UO_2478 (O_2478,N_19869,N_19877);
or UO_2479 (O_2479,N_19874,N_19918);
nand UO_2480 (O_2480,N_19905,N_19906);
or UO_2481 (O_2481,N_19992,N_19995);
and UO_2482 (O_2482,N_19972,N_19992);
or UO_2483 (O_2483,N_19972,N_19991);
or UO_2484 (O_2484,N_19983,N_19960);
nor UO_2485 (O_2485,N_19858,N_19902);
nor UO_2486 (O_2486,N_19844,N_19938);
xnor UO_2487 (O_2487,N_19924,N_19841);
and UO_2488 (O_2488,N_19925,N_19944);
nand UO_2489 (O_2489,N_19861,N_19840);
xor UO_2490 (O_2490,N_19992,N_19857);
xor UO_2491 (O_2491,N_19858,N_19880);
or UO_2492 (O_2492,N_19965,N_19841);
and UO_2493 (O_2493,N_19857,N_19936);
nor UO_2494 (O_2494,N_19990,N_19920);
nor UO_2495 (O_2495,N_19985,N_19953);
and UO_2496 (O_2496,N_19993,N_19911);
and UO_2497 (O_2497,N_19987,N_19904);
nor UO_2498 (O_2498,N_19870,N_19967);
nor UO_2499 (O_2499,N_19944,N_19850);
endmodule